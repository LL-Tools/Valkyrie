

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9565, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9616, n9617, n9618,
         n9620, n9621, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,
         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,
         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,
         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
         n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,
         n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
         n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
         n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
         n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,
         n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
         n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,
         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
         n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,
         n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,
         n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,
         n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
         n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
         n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
         n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,
         n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,
         n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
         n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
         n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,
         n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
         n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
         n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,
         n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
         n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432,
         n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440,
         n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,
         n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
         n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
         n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
         n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,
         n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,
         n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
         n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504,
         n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,
         n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,
         n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528,
         n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536,
         n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544,
         n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,
         n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,
         n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568,
         n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576,
         n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,
         n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,
         n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600,
         n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608,
         n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616,
         n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624,
         n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632,
         n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640,
         n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648,
         n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656,
         n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664,
         n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672,
         n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680,
         n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688,
         n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,
         n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704,
         n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,
         n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720,
         n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,
         n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
         n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
         n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
         n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,
         n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
         n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,
         n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,
         n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,
         n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,
         n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,
         n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
         n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,
         n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,
         n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
         n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,
         n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
         n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,
         n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,
         n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,
         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
         n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,
         n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
         n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
         n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,
         n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
         n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,
         n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,
         n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,
         n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
         n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968,
         n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,
         n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
         n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992,
         n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
         n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
         n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016,
         n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024,
         n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,
         n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040,
         n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048,
         n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056,
         n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064,
         n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072,
         n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080,
         n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088,
         n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096,
         n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104,
         n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112,
         n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120,
         n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128,
         n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136,
         n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144,
         n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152,
         n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160,
         n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168,
         n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176,
         n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184,
         n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192,
         n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200,
         n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208,
         n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216,
         n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224,
         n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232,
         n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240,
         n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248,
         n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256,
         n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264,
         n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272,
         n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280,
         n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288,
         n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296,
         n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304,
         n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312,
         n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320,
         n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328,
         n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336,
         n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344,
         n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352,
         n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360,
         n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368,
         n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376,
         n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384,
         n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392,
         n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400,
         n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408,
         n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416,
         n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424,
         n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432,
         n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440,
         n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448,
         n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456,
         n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464,
         n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472,
         n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480,
         n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488,
         n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496,
         n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504,
         n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512,
         n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520,
         n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528,
         n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536,
         n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544,
         n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552,
         n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560,
         n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568,
         n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576,
         n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584,
         n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592,
         n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600,
         n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608,
         n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616,
         n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624,
         n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632,
         n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640,
         n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648,
         n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656,
         n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664,
         n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672,
         n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680,
         n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688,
         n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696,
         n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704,
         n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712,
         n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720,
         n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728,
         n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736,
         n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744,
         n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752,
         n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760,
         n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768,
         n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776,
         n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784,
         n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792,
         n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800,
         n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808,
         n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816,
         n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824,
         n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832,
         n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840,
         n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848,
         n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856,
         n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864,
         n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872,
         n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880,
         n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888,
         n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896,
         n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904,
         n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912,
         n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920,
         n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928,
         n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936,
         n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944,
         n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952,
         n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960,
         n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968,
         n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976,
         n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984,
         n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992,
         n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000,
         n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008,
         n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016,
         n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024,
         n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032,
         n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040,
         n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048,
         n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056,
         n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064,
         n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072,
         n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080,
         n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088,
         n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096,
         n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104,
         n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112,
         n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120,
         n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128,
         n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136,
         n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144,
         n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152,
         n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160,
         n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168,
         n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176,
         n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184,
         n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192,
         n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200,
         n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208,
         n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216,
         n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224,
         n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232,
         n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240,
         n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248,
         n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256,
         n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264,
         n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272,
         n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280,
         n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288,
         n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296,
         n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304,
         n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312,
         n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320,
         n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328,
         n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336,
         n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344,
         n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352,
         n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360,
         n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368,
         n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376,
         n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384,
         n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392,
         n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,
         n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408,
         n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416,
         n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,
         n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432,
         n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440,
         n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448,
         n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456,
         n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464,
         n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472,
         n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480,
         n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488,
         n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496,
         n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504,
         n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512,
         n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520,
         n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528,
         n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536,
         n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544,
         n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552,
         n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560,
         n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568,
         n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576,
         n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584,
         n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592,
         n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600,
         n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608,
         n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616,
         n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624,
         n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632,
         n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640,
         n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648,
         n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656,
         n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664,
         n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672,
         n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680,
         n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688,
         n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696,
         n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704,
         n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712,
         n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720,
         n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728,
         n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736,
         n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744,
         n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752,
         n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760,
         n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768,
         n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776,
         n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784,
         n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792,
         n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800,
         n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808,
         n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816,
         n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824,
         n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832,
         n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840,
         n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848,
         n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856,
         n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864,
         n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872,
         n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880,
         n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888,
         n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896,
         n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904,
         n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912,
         n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920,
         n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928,
         n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936,
         n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944,
         n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952,
         n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960,
         n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968,
         n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976,
         n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984,
         n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992,
         n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000,
         n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008,
         n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016,
         n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024,
         n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032,
         n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040,
         n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048,
         n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056,
         n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064,
         n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072,
         n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080,
         n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088,
         n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096,
         n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104,
         n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112,
         n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120,
         n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128,
         n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136,
         n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144,
         n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152,
         n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160,
         n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168,
         n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176,
         n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184,
         n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192,
         n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200,
         n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208,
         n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216,
         n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224,
         n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232,
         n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240,
         n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248,
         n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256,
         n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264,
         n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272,
         n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280,
         n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288,
         n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296,
         n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304,
         n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312,
         n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320,
         n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328,
         n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336,
         n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344,
         n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352,
         n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360,
         n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368,
         n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376,
         n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384,
         n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392,
         n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400,
         n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408,
         n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416,
         n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424,
         n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432,
         n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440,
         n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448,
         n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456,
         n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464,
         n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472,
         n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480,
         n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488,
         n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496,
         n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504,
         n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512,
         n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520,
         n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528,
         n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536,
         n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544,
         n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552,
         n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560,
         n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568,
         n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576,
         n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584,
         n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592,
         n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600,
         n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608,
         n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616,
         n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624,
         n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632,
         n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640,
         n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648,
         n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656,
         n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664,
         n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672,
         n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680,
         n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688,
         n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696,
         n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704,
         n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712,
         n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720,
         n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728,
         n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736,
         n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744,
         n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752,
         n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760,
         n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768,
         n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776,
         n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784,
         n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792,
         n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800,
         n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808,
         n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816,
         n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824,
         n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832,
         n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840,
         n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848,
         n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856,
         n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864,
         n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872,
         n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880,
         n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888,
         n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896,
         n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904,
         n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912,
         n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920,
         n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928,
         n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936,
         n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944,
         n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952,
         n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960,
         n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968,
         n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976,
         n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984,
         n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992,
         n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000,
         n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008,
         n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016,
         n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024,
         n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032,
         n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040,
         n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048,
         n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056,
         n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064,
         n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072,
         n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080,
         n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088,
         n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096,
         n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104,
         n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112,
         n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120,
         n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128,
         n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136,
         n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144,
         n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152,
         n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160,
         n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168,
         n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176,
         n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184,
         n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192,
         n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200,
         n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208,
         n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216,
         n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224,
         n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232,
         n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240,
         n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248,
         n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256,
         n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264,
         n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272,
         n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280,
         n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288,
         n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296,
         n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304,
         n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312,
         n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320,
         n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328,
         n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336,
         n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344,
         n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352,
         n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360,
         n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368,
         n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376,
         n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384,
         n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392,
         n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400,
         n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408,
         n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416,
         n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424,
         n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432,
         n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440,
         n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448,
         n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456,
         n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464,
         n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472,
         n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480,
         n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488,
         n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496,
         n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504,
         n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512,
         n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520,
         n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528,
         n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536,
         n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544,
         n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552,
         n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560,
         n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568,
         n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576,
         n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584,
         n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592,
         n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600,
         n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608,
         n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616,
         n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624,
         n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632,
         n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640,
         n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648,
         n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656,
         n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664,
         n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672,
         n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680,
         n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688,
         n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696,
         n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704,
         n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712,
         n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720,
         n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728,
         n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736,
         n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744,
         n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752,
         n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760,
         n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768,
         n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776,
         n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784,
         n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792,
         n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800,
         n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808,
         n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816,
         n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824,
         n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832,
         n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840,
         n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848,
         n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856,
         n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864,
         n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872,
         n20873, n20874, n20875, n20876, n20877, n20878, n20879, n20880,
         n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888,
         n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896,
         n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904,
         n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912,
         n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920,
         n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928,
         n20929, n20930, n20931, n20932, n20933, n20934, n20935, n20936,
         n20937, n20938, n20939, n20940, n20941, n20942, n20943, n20944,
         n20945, n20946, n20947, n20948, n20949, n20950, n20951, n20952,
         n20953, n20954, n20955, n20956, n20957, n20958, n20959, n20960,
         n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968,
         n20969, n20970, n20971, n20972, n20973, n20974, n20975, n20976,
         n20977, n20978, n20979, n20980, n20981, n20982, n20983, n20984,
         n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992,
         n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000,
         n21001, n21002, n21003, n21004, n21005, n21006, n21007, n21008,
         n21009, n21010, n21011, n21012, n21013, n21014, n21015, n21016,
         n21017, n21018, n21019, n21020, n21021, n21022, n21023, n21024,
         n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032,
         n21033, n21034, n21035, n21036, n21037, n21038, n21039, n21040,
         n21041, n21042, n21043, n21044, n21045, n21046, n21047, n21048,
         n21049, n21050, n21051, n21052, n21053, n21054, n21055, n21056,
         n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21064,
         n21065, n21066, n21067, n21068, n21069, n21070, n21071, n21072,
         n21073, n21074, n21075, n21076, n21077, n21078, n21079, n21080,
         n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088,
         n21089, n21090, n21091, n21092, n21093, n21094, n21095, n21096,
         n21097, n21098, n21099, n21100, n21101, n21102, n21103, n21104,
         n21105, n21106, n21107, n21108, n21109, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21124, n21125, n21126, n21127, n21128, n21129, n21130,
         n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138,
         n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21146,
         n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154,
         n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162,
         n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170,
         n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178,
         n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186,
         n21187, n21188, n21189, n21190, n21191, n21192, n21193, n21194,
         n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202,
         n21203, n21204, n21205, n21206, n21207, n21208, n21209, n21210,
         n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218,
         n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226,
         n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234,
         n21235, n21236, n21237, n21238, n21239, n21240, n21241, n21242,
         n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250,
         n21251, n21252, n21253, n21254, n21255, n21256, n21257, n21258,
         n21259, n21260, n21261, n21262, n21263, n21264, n21265, n21266,
         n21267, n21268, n21269, n21270, n21271, n21272, n21273, n21274,
         n21275, n21276, n21277, n21278, n21279, n21280, n21281, n21282,
         n21283, n21284, n21285, n21286, n21287, n21288, n21289, n21290,
         n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298,
         n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306,
         n21307, n21308, n21309, n21310, n21311, n21312, n21313, n21314,
         n21315, n21316, n21317, n21318, n21319, n21320, n21321, n21322,
         n21323, n21324, n21325, n21326, n21327, n21328, n21329, n21330,
         n21331, n21332, n21333, n21334, n21335, n21336, n21337, n21338,
         n21339, n21340, n21341, n21342, n21343, n21344, n21345, n21346,
         n21347, n21348, n21349, n21350, n21351, n21352, n21353, n21354,
         n21355, n21356, n21357, n21358, n21359, n21360, n21361, n21362,
         n21363, n21364, n21365, n21366, n21367, n21368, n21369, n21370,
         n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378,
         n21379, n21380, n21381, n21382, n21383, n21384, n21385, n21386,
         n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394;

  OR2_X1 U11008 ( .A1(n21219), .A2(n13309), .ZN(n20410) );
  BUF_X4 U11009 ( .A(n13202), .Z(n9569) );
  NAND2_X1 U11010 ( .A1(n16908), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16907) );
  XNOR2_X1 U11011 ( .A(n12010), .B(n12008), .ZN(n14157) );
  CLKBUF_X2 U11012 ( .A(n10994), .Z(n11400) );
  CLKBUF_X2 U11013 ( .A(n13658), .Z(n17967) );
  CLKBUF_X1 U11014 ( .A(n12585), .Z(n12953) );
  CLKBUF_X2 U11015 ( .A(n12382), .Z(n13016) );
  CLKBUF_X2 U11016 ( .A(n12451), .Z(n13510) );
  BUF_X2 U11017 ( .A(n12368), .Z(n13513) );
  CLKBUF_X2 U11018 ( .A(n12358), .Z(n13503) );
  INV_X2 U11019 ( .A(n17948), .ZN(n17844) );
  INV_X1 U11020 ( .A(n11921), .ZN(n17931) );
  NAND2_X1 U11021 ( .A1(n9798), .A2(n10341), .ZN(n10901) );
  BUF_X1 U11022 ( .A(n11980), .Z(n12136) );
  CLKBUF_X2 U11023 ( .A(n13741), .Z(n9574) );
  CLKBUF_X2 U11024 ( .A(n13741), .Z(n9573) );
  INV_X1 U11025 ( .A(n9579), .ZN(n9580) );
  INV_X1 U11026 ( .A(n9579), .ZN(n9582) );
  NAND2_X1 U11027 ( .A1(n9907), .A2(n9906), .ZN(n9909) );
  CLKBUF_X2 U11028 ( .A(n13741), .Z(n9572) );
  INV_X1 U11029 ( .A(n13685), .ZN(n12101) );
  AND4_X1 U11030 ( .A1(n12372), .A2(n12371), .A3(n12370), .A4(n12369), .ZN(
        n12378) );
  INV_X1 U11031 ( .A(n12109), .ZN(n9575) );
  CLKBUF_X1 U11032 ( .A(n17980), .Z(n9568) );
  INV_X1 U11033 ( .A(n13676), .ZN(n9579) );
  AND2_X1 U11035 ( .A1(n10832), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9601) );
  AND2_X1 U11036 ( .A1(n9787), .A2(n13968), .ZN(n12453) );
  AND2_X1 U11037 ( .A1(n12279), .A2(n12276), .ZN(n12452) );
  AND2_X1 U11038 ( .A1(n9787), .A2(n13967), .ZN(n12383) );
  AND2_X1 U11039 ( .A1(n14023), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12277) );
  INV_X4 U11040 ( .A(n18739), .ZN(n18693) );
  INV_X1 U11042 ( .A(n21393), .ZN(n9565) );
  INV_X1 U11044 ( .A(n21394), .ZN(n9567) );
  CLKBUF_X1 U11046 ( .A(n12585), .Z(n9591) );
  INV_X1 U11047 ( .A(n13106), .ZN(n12451) );
  BUF_X1 U11048 ( .A(n12484), .Z(n13512) );
  NOR2_X2 U11049 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10449) );
  NAND2_X1 U11050 ( .A1(n9909), .A2(n10901), .ZN(n10847) );
  INV_X1 U11051 ( .A(n14658), .ZN(n13310) );
  INV_X2 U11052 ( .A(n12101), .ZN(n17817) );
  AND2_X1 U11053 ( .A1(n14658), .A2(n13324), .ZN(n13395) );
  INV_X1 U11054 ( .A(n13526), .ZN(n13032) );
  AND4_X1 U11056 ( .A1(n10612), .A2(n10611), .A3(n10610), .A4(n10398), .ZN(
        n16378) );
  NOR2_X1 U11057 ( .A1(n11022), .A2(n10345), .ZN(n19740) );
  OAI22_X1 U11058 ( .A1(n12173), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n19188), .ZN(n12182) );
  INV_X1 U11059 ( .A(n9579), .ZN(n9581) );
  INV_X1 U11060 ( .A(n9579), .ZN(n9583) );
  AND2_X1 U11061 ( .A1(n13760), .A2(n11888), .ZN(n13658) );
  NAND2_X1 U11062 ( .A1(n18298), .A2(n12023), .ZN(n18331) );
  NOR2_X1 U11063 ( .A1(n10319), .A2(n11422), .ZN(n11446) );
  XNOR2_X1 U11064 ( .A(n11588), .B(n11586), .ZN(n14005) );
  INV_X1 U11065 ( .A(n9909), .ZN(n13904) );
  MUX2_X1 U11066 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n13439), .S(
        n13438), .Z(n16761) );
  AOI211_X1 U11067 ( .C1(n18593), .C2(n14156), .A(n14155), .B(n14154), .ZN(
        n14257) );
  INV_X1 U11068 ( .A(n20424), .ZN(n20405) );
  INV_X1 U11069 ( .A(n15957), .ZN(n19400) );
  INV_X1 U11070 ( .A(n19445), .ZN(n19476) );
  AND2_X1 U11071 ( .A1(n10878), .A2(n17236), .ZN(n11409) );
  INV_X1 U11072 ( .A(n19794), .ZN(n19756) );
  OR2_X1 U11073 ( .A1(n11894), .A2(n11893), .ZN(n12224) );
  INV_X1 U11074 ( .A(n20404), .ZN(n20432) );
  NAND2_X1 U11075 ( .A1(n20070), .A2(n19870), .ZN(n19947) );
  NAND2_X1 U11076 ( .A1(n20037), .A2(n20036), .ZN(n20122) );
  INV_X1 U11077 ( .A(n18426), .ZN(n18490) );
  INV_X1 U11078 ( .A(n19347), .ZN(n19261) );
  NAND3_X2 U11079 ( .A1(n10255), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11846) );
  INV_X2 U11080 ( .A(n11846), .ZN(n10821) );
  AND2_X1 U11081 ( .A1(n12277), .A2(n13968), .ZN(n13505) );
  INV_X1 U11082 ( .A(n12452), .ZN(n9589) );
  NAND2_X1 U11083 ( .A1(n13170), .A2(n13194), .ZN(n13202) );
  NOR2_X2 U11084 ( .A1(n16932), .A2(n18251), .ZN(n16908) );
  AND2_X2 U11085 ( .A1(n12405), .A2(n12439), .ZN(n13271) );
  MUX2_X2 U11086 ( .A(n18730), .B(n13787), .S(n14105), .Z(n19171) );
  XNOR2_X2 U11088 ( .A(n9884), .B(n9681), .ZN(n11524) );
  OR2_X2 U11089 ( .A1(n14532), .A2(n20583), .ZN(n9674) );
  NAND2_X2 U11090 ( .A1(n18554), .A2(n18730), .ZN(n18593) );
  OR2_X2 U11091 ( .A1(n14518), .A2(n14519), .ZN(n9657) );
  NAND2_X1 U11092 ( .A1(n10065), .A2(n10990), .ZN(n10321) );
  XNOR2_X2 U11093 ( .A(n11951), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n14115) );
  XNOR2_X2 U11094 ( .A(n11953), .B(n11950), .ZN(n11951) );
  NOR2_X2 U11095 ( .A1(n18197), .A2(n18050), .ZN(n18046) );
  NOR2_X2 U11097 ( .A1(n14266), .A2(n10305), .ZN(n14330) );
  AND2_X2 U11098 ( .A1(n15139), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10382) );
  NOR2_X2 U11099 ( .A1(n14044), .A2(n17945), .ZN(n17862) );
  NAND2_X1 U11100 ( .A1(n13760), .A2(n11879), .ZN(n17980) );
  INV_X1 U11101 ( .A(n19335), .ZN(n18178) );
  NOR2_X2 U11102 ( .A1(n14251), .A2(n18678), .ZN(n14250) );
  BUF_X4 U11104 ( .A(n16829), .Z(n9571) );
  INV_X1 U11105 ( .A(n11287), .ZN(n16829) );
  OAI21_X2 U11106 ( .B1(n14114), .B2(n14115), .A(n11952), .ZN(n11970) );
  NAND2_X2 U11107 ( .A1(n14312), .A2(n13166), .ZN(n14429) );
  NAND2_X2 U11108 ( .A1(n14313), .A2(n14314), .ZN(n14312) );
  BUF_X4 U11109 ( .A(n11297), .Z(n11399) );
  NAND3_X2 U11110 ( .A1(n9972), .A2(n10966), .A3(n9971), .ZN(n10979) );
  INV_X2 U11112 ( .A(n9575), .ZN(n9576) );
  INV_X2 U11113 ( .A(n9575), .ZN(n9577) );
  INV_X2 U11114 ( .A(n9575), .ZN(n9578) );
  AND2_X1 U11115 ( .A1(n11884), .A2(n13784), .ZN(n12109) );
  NOR2_X4 U11116 ( .A1(n10810), .A2(n10809), .ZN(n16846) );
  MUX2_X2 U11117 ( .A(n10833), .B(n10808), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n10810) );
  AND2_X2 U11118 ( .A1(n12400), .A2(n13539), .ZN(n14480) );
  OAI21_X4 U11119 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19340), .A(n17362), 
        .ZN(n18495) );
  AND2_X4 U11120 ( .A1(n12277), .A2(n10082), .ZN(n9607) );
  AND3_X2 U11121 ( .A1(n12283), .A2(n12282), .A3(n10422), .ZN(n12284) );
  AOI21_X2 U11122 ( .B1(n19175), .B2(n19192), .A(n19174), .ZN(n19176) );
  XNOR2_X2 U11123 ( .A(n13165), .B(n20548), .ZN(n14314) );
  AND2_X1 U11124 ( .A1(n13785), .A2(n11886), .ZN(n13676) );
  NOR2_X2 U11125 ( .A1(n17012), .A2(n18464), .ZN(n18456) );
  NAND2_X2 U11126 ( .A1(n15315), .A2(n13164), .ZN(n13165) );
  CLKBUF_X1 U11127 ( .A(n16295), .Z(n16299) );
  NAND2_X1 U11128 ( .A1(n9970), .A2(n9811), .ZN(n16405) );
  OAI21_X1 U11129 ( .B1(n19957), .B2(n19972), .A(n20133), .ZN(n19975) );
  MUX2_X1 U11130 ( .A(n14659), .B(n14658), .S(n9657), .Z(n14661) );
  AOI21_X1 U11131 ( .B1(n9896), .B2(n9736), .A(n9893), .ZN(n9892) );
  NAND2_X1 U11132 ( .A1(n20037), .A2(n20069), .ZN(n20187) );
  AND3_X1 U11133 ( .A1(n11029), .A2(n11009), .A3(n11019), .ZN(n10105) );
  INV_X2 U11134 ( .A(n9600), .ZN(n18381) );
  INV_X1 U11135 ( .A(n18407), .ZN(n18656) );
  AND4_X1 U11136 ( .A1(n11011), .A2(n11020), .A3(n11018), .A4(n11008), .ZN(
        n10106) );
  AOI22_X1 U11137 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19740), .B1(
        n19651), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11009) );
  NAND2_X1 U11138 ( .A1(n14004), .A2(n14007), .ZN(n20288) );
  AND2_X1 U11139 ( .A1(n11026), .A2(n11013), .ZN(n19605) );
  NAND2_X1 U11140 ( .A1(n12656), .A2(n12659), .ZN(n20662) );
  NAND2_X1 U11141 ( .A1(n11026), .A2(n11024), .ZN(n16811) );
  INV_X1 U11142 ( .A(n18361), .ZN(n9586) );
  NAND3_X1 U11143 ( .A1(n10048), .A2(n9788), .A3(n10047), .ZN(n12646) );
  NAND2_X1 U11144 ( .A1(n10093), .A2(n10092), .ZN(n18361) );
  AND2_X1 U11145 ( .A1(n15401), .A2(n20579), .ZN(n20545) );
  AND2_X1 U11146 ( .A1(n11014), .A2(n11013), .ZN(n19880) );
  NOR2_X1 U11147 ( .A1(n14009), .A2(n9954), .ZN(n18101) );
  CLKBUF_X2 U11148 ( .A(n11006), .Z(n9613) );
  NAND2_X1 U11149 ( .A1(n11409), .A2(n16847), .ZN(n16515) );
  OR2_X1 U11150 ( .A1(n12923), .A2(n15195), .ZN(n12924) );
  NAND2_X1 U11151 ( .A1(n14157), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12012) );
  INV_X2 U11152 ( .A(n19386), .ZN(n15967) );
  NAND2_X1 U11153 ( .A1(n11171), .A2(n11197), .ZN(n11195) );
  INV_X2 U11154 ( .A(n18680), .ZN(n18730) );
  NAND2_X1 U11155 ( .A1(n13754), .A2(n13606), .ZN(n18680) );
  AND2_X1 U11156 ( .A1(n17361), .A2(n9771), .ZN(n13722) );
  NAND2_X1 U11157 ( .A1(n12204), .A2(n18175), .ZN(n17361) );
  NAND2_X1 U11158 ( .A1(n10944), .A2(n13713), .ZN(n10966) );
  AOI21_X1 U11159 ( .B1(n14149), .B2(n14544), .A(n13316), .ZN(n14305) );
  CLKBUF_X2 U11160 ( .A(n10517), .Z(n10703) );
  CLKBUF_X3 U11161 ( .A(n13324), .Z(n14544) );
  NOR2_X1 U11162 ( .A1(n10847), .A2(n10890), .ZN(n10855) );
  AND2_X1 U11163 ( .A1(n15992), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10954) );
  CLKBUF_X1 U11164 ( .A(n12411), .Z(n20615) );
  INV_X1 U11165 ( .A(n11088), .ZN(n10356) );
  INV_X1 U11166 ( .A(n10730), .ZN(n10454) );
  INV_X4 U11167 ( .A(n11716), .ZN(n15992) );
  NAND2_X1 U11168 ( .A1(n20603), .A2(n14486), .ZN(n21216) );
  NAND2_X1 U11169 ( .A1(n12061), .A2(n12060), .ZN(n18755) );
  AND2_X2 U11170 ( .A1(n10884), .A2(n20306), .ZN(n10479) );
  INV_X4 U11171 ( .A(n10884), .ZN(n11716) );
  NOR2_X1 U11172 ( .A1(n10884), .A2(n20311), .ZN(n10945) );
  INV_X1 U11173 ( .A(n19619), .ZN(n10903) );
  INV_X2 U11174 ( .A(n12406), .ZN(n12411) );
  OAI21_X1 U11175 ( .B1(n10284), .B2(n10283), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10282) );
  AND4_X1 U11176 ( .A1(n12275), .A2(n12274), .A3(n12273), .A4(n12272), .ZN(
        n12285) );
  AND2_X1 U11177 ( .A1(n11900), .A2(n11903), .ZN(n10089) );
  AND4_X1 U11178 ( .A1(n12304), .A2(n12303), .A3(n12302), .A4(n12301), .ZN(
        n12316) );
  INV_X4 U11180 ( .A(n10404), .ZN(n12119) );
  CLKBUF_X2 U11181 ( .A(n13657), .Z(n17833) );
  CLKBUF_X2 U11182 ( .A(n10590), .Z(n11677) );
  CLKBUF_X2 U11183 ( .A(n10505), .Z(n11683) );
  AND2_X2 U11184 ( .A1(n11697), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10594) );
  AND2_X1 U11185 ( .A1(n12278), .A2(n13951), .ZN(n12331) );
  CLKBUF_X1 U11186 ( .A(n9614), .Z(n9584) );
  AND2_X2 U11187 ( .A1(n12279), .A2(n13949), .ZN(n12368) );
  CLKBUF_X2 U11188 ( .A(n11960), .Z(n14172) );
  INV_X1 U11189 ( .A(n13106), .ZN(n9585) );
  AND2_X2 U11190 ( .A1(n13968), .A2(n13949), .ZN(n12358) );
  NAND2_X1 U11191 ( .A1(n12276), .A2(n13967), .ZN(n13110) );
  INV_X2 U11192 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12171) );
  INV_X2 U11193 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10783) );
  INV_X1 U11195 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n19196) );
  AND2_X1 U11196 ( .A1(n11560), .A2(n10041), .ZN(n10040) );
  AOI21_X1 U11197 ( .B1(n16097), .B2(n19384), .A(n10122), .ZN(n10121) );
  NOR2_X1 U11198 ( .A1(n9806), .A2(n16325), .ZN(n16614) );
  OR2_X1 U11199 ( .A1(n15598), .A2(n15597), .ZN(n16430) );
  NAND2_X1 U11200 ( .A1(n9794), .A2(n10374), .ZN(n10141) );
  OR2_X1 U11201 ( .A1(n16532), .A2(n19574), .ZN(n9781) );
  AOI21_X1 U11202 ( .B1(n15111), .B2(n20518), .A(n15110), .ZN(n15112) );
  AOI21_X1 U11203 ( .B1(n11426), .B2(n15620), .A(n15596), .ZN(n16097) );
  AOI21_X1 U11204 ( .B1(n16324), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n9806) );
  AOI21_X1 U11205 ( .B1(n10417), .B2(n17224), .A(n16542), .ZN(n16543) );
  XNOR2_X1 U11206 ( .A(n10333), .B(n9737), .ZN(n10417) );
  AOI21_X1 U11207 ( .B1(n11512), .B2(n11419), .A(n11456), .ZN(n16433) );
  XNOR2_X1 U11208 ( .A(n11541), .B(n11540), .ZN(n11870) );
  AND2_X1 U11209 ( .A1(n9871), .A2(n9867), .ZN(n15148) );
  CLKBUF_X1 U11210 ( .A(n11425), .Z(n15620) );
  NAND2_X1 U11211 ( .A1(n9886), .A2(n9885), .ZN(n9884) );
  NAND2_X1 U11212 ( .A1(n11476), .A2(n9654), .ZN(n16235) );
  NAND2_X1 U11213 ( .A1(n11474), .A2(n10352), .ZN(n16280) );
  XNOR2_X1 U11214 ( .A(n9664), .B(n13534), .ZN(n14588) );
  NAND2_X1 U11215 ( .A1(n16264), .A2(n11466), .ZN(n10333) );
  AND2_X1 U11216 ( .A1(n15139), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15150) );
  AND2_X1 U11217 ( .A1(n11418), .A2(n10364), .ZN(n11456) );
  AND2_X1 U11218 ( .A1(n11861), .A2(n11862), .ZN(n9863) );
  AOI21_X1 U11219 ( .B1(n13295), .B2(n13294), .A(n14662), .ZN(n15118) );
  NAND2_X1 U11220 ( .A1(n9873), .A2(n9872), .ZN(n15145) );
  NAND2_X1 U11221 ( .A1(n11278), .A2(n11277), .ZN(n11450) );
  CLKBUF_X1 U11222 ( .A(n14675), .Z(n14676) );
  CLKBUF_X2 U11223 ( .A(n11475), .Z(n11476) );
  NAND2_X1 U11224 ( .A1(n16283), .A2(n11465), .ZN(n16264) );
  NAND2_X1 U11225 ( .A1(n10008), .A2(n9692), .ZN(n14537) );
  NAND2_X1 U11226 ( .A1(n10010), .A2(n13211), .ZN(n15185) );
  NAND2_X1 U11227 ( .A1(n11497), .A2(n11463), .ZN(n16283) );
  NAND2_X1 U11228 ( .A1(n9812), .A2(n10037), .ZN(n16351) );
  OR2_X1 U11229 ( .A1(n14706), .A2(n14707), .ZN(n9872) );
  XNOR2_X1 U11230 ( .A(n11479), .B(n11478), .ZN(n11859) );
  NAND3_X1 U11231 ( .A1(n16250), .A2(n9928), .A3(n10129), .ZN(n9926) );
  NOR2_X1 U11232 ( .A1(n11479), .A2(n11478), .ZN(n11405) );
  NAND2_X1 U11233 ( .A1(n10070), .A2(n10074), .ZN(n11495) );
  OAI21_X1 U11234 ( .B1(n9732), .B2(n9663), .A(n9631), .ZN(n15160) );
  NAND2_X1 U11235 ( .A1(n10007), .A2(n15203), .ZN(n10008) );
  CLKBUF_X1 U11236 ( .A(n14705), .Z(n14706) );
  NAND2_X1 U11237 ( .A1(n9945), .A2(n9792), .ZN(n15203) );
  OR2_X1 U11238 ( .A1(n16314), .A2(n10077), .ZN(n10070) );
  NAND2_X1 U11239 ( .A1(n9882), .A2(n11415), .ZN(n9881) );
  NAND2_X1 U11240 ( .A1(n10327), .A2(n9640), .ZN(n16314) );
  INV_X2 U11241 ( .A(n10405), .ZN(n9611) );
  INV_X2 U11242 ( .A(n10405), .ZN(n14969) );
  INV_X1 U11243 ( .A(n10038), .ZN(n10037) );
  NAND2_X1 U11244 ( .A1(n10384), .A2(n10383), .ZN(n15211) );
  NAND2_X1 U11245 ( .A1(n11170), .A2(n11169), .ZN(n11459) );
  NAND2_X1 U11246 ( .A1(n9986), .A2(n9987), .ZN(n9985) );
  NOR2_X1 U11247 ( .A1(n10235), .A2(n10176), .ZN(n10175) );
  NOR2_X1 U11248 ( .A1(n11263), .A2(n10133), .ZN(n10132) );
  AND2_X1 U11249 ( .A1(n10027), .A2(n16376), .ZN(n10347) );
  NAND2_X1 U11250 ( .A1(n9948), .A2(n13181), .ZN(n9947) );
  AND2_X1 U11251 ( .A1(n9944), .A2(n13208), .ZN(n9792) );
  NOR2_X1 U11252 ( .A1(n15323), .A2(n20575), .ZN(n10176) );
  AND2_X1 U11253 ( .A1(n9903), .A2(n9901), .ZN(n10128) );
  AND2_X1 U11254 ( .A1(n18263), .A2(n12030), .ZN(n9989) );
  AND2_X1 U11255 ( .A1(n13198), .A2(n13192), .ZN(n10383) );
  NAND2_X1 U11256 ( .A1(n11045), .A2(n11044), .ZN(n16724) );
  OR2_X1 U11257 ( .A1(n11067), .A2(n11066), .ZN(n16711) );
  AND2_X1 U11258 ( .A1(n11064), .A2(n11075), .ZN(n16379) );
  AND3_X1 U11259 ( .A1(n14436), .A2(n14445), .A3(n14462), .ZN(n12701) );
  XNOR2_X1 U11260 ( .A(n9862), .B(n9861), .ZN(n16012) );
  NAND2_X1 U11261 ( .A1(n16929), .A2(n12022), .ZN(n12026) );
  NOR2_X1 U11262 ( .A1(n15362), .A2(n10023), .ZN(n15320) );
  NAND2_X1 U11263 ( .A1(n14300), .A2(n12677), .ZN(n14294) );
  NAND2_X1 U11264 ( .A1(n13134), .A2(n13133), .ZN(n13168) );
  NAND2_X1 U11265 ( .A1(n12618), .A2(n12617), .ZN(n14436) );
  OR2_X1 U11266 ( .A1(n16022), .A2(n9965), .ZN(n9862) );
  NAND2_X1 U11267 ( .A1(n10066), .A2(n11062), .ZN(n11141) );
  NAND4_X1 U11268 ( .A1(n9676), .A2(n10067), .A3(n9636), .A4(n11054), .ZN(
        n10066) );
  NOR2_X2 U11269 ( .A1(n19910), .A2(n19914), .ZN(n19974) );
  NOR2_X2 U11270 ( .A1(n20131), .A2(n19804), .ZN(n19866) );
  NAND2_X1 U11271 ( .A1(n11291), .A2(n11254), .ZN(n15643) );
  XNOR2_X1 U11272 ( .A(n13170), .B(n12600), .ZN(n13182) );
  NOR2_X2 U11273 ( .A1(n19914), .A2(n19840), .ZN(n19708) );
  NAND3_X1 U11274 ( .A1(n12655), .A2(n9706), .A3(n14146), .ZN(n14300) );
  NAND2_X1 U11275 ( .A1(n16821), .A2(n19482), .ZN(n19840) );
  NAND2_X1 U11276 ( .A1(n12654), .A2(n12653), .ZN(n12655) );
  AND2_X2 U11277 ( .A1(n18455), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n18391) );
  CLKBUF_X1 U11278 ( .A(n13145), .Z(n20585) );
  NAND2_X1 U11279 ( .A1(n16821), .A2(n16820), .ZN(n19804) );
  OR2_X1 U11280 ( .A1(n16821), .A2(n19482), .ZN(n19948) );
  NAND2_X1 U11281 ( .A1(n10293), .A2(n10294), .ZN(n14240) );
  OR2_X1 U11282 ( .A1(n16821), .A2(n16820), .ZN(n19910) );
  NAND2_X1 U11283 ( .A1(n12664), .A2(n12663), .ZN(n14146) );
  NAND2_X1 U11284 ( .A1(n14109), .A2(n14110), .ZN(n10294) );
  NAND2_X1 U11285 ( .A1(n19598), .A2(n19597), .ZN(n20131) );
  AND3_X1 U11286 ( .A1(n11055), .A2(n10069), .A3(n10068), .ZN(n10067) );
  NAND2_X1 U11287 ( .A1(n13011), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13054) );
  INV_X1 U11288 ( .A(n18343), .ZN(n18525) );
  CLKBUF_X2 U11289 ( .A(n18493), .Z(n9600) );
  AND2_X1 U11290 ( .A1(n11571), .A2(n14341), .ZN(n14109) );
  NOR2_X1 U11291 ( .A1(n16811), .A2(n11027), .ZN(n11028) );
  AOI22_X1 U11292 ( .A1(n19846), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n11057), .ZN(n11011) );
  INV_X1 U11293 ( .A(n12646), .ZN(n12648) );
  AOI22_X1 U11294 ( .A1(n19980), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n16822), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11008) );
  OR2_X1 U11295 ( .A1(n20039), .A2(n11017), .ZN(n11018) );
  NOR2_X1 U11296 ( .A1(n11245), .A2(n10228), .ZN(n11253) );
  NOR2_X1 U11297 ( .A1(n11245), .A2(n11244), .ZN(n11246) );
  OR2_X1 U11298 ( .A1(n17232), .A2(n10931), .ZN(n17214) );
  NAND2_X1 U11299 ( .A1(n12658), .A2(n12657), .ZN(n12659) );
  AND2_X1 U11300 ( .A1(n14806), .A2(n14807), .ZN(n14788) );
  AND2_X1 U11301 ( .A1(n11188), .A2(n11203), .ZN(n15792) );
  AND2_X1 U11302 ( .A1(n13996), .A2(n14001), .ZN(n20275) );
  NAND2_X1 U11303 ( .A1(n12943), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13009) );
  INV_X1 U11304 ( .A(n20570), .ZN(n15515) );
  NAND2_X1 U11305 ( .A1(n14186), .A2(n9769), .ZN(n19186) );
  AND2_X1 U11306 ( .A1(n13996), .A2(n11580), .ZN(n14006) );
  NOR2_X2 U11307 ( .A1(n18734), .A2(n16880), .ZN(n18672) );
  AND2_X1 U11308 ( .A1(n10045), .A2(n10136), .ZN(n9788) );
  NAND2_X1 U11309 ( .A1(n10051), .A2(n9671), .ZN(n12647) );
  NAND2_X1 U11310 ( .A1(n12012), .A2(n9703), .ZN(n18437) );
  AND2_X1 U11311 ( .A1(n14502), .A2(n14648), .ZN(n20570) );
  AND2_X1 U11312 ( .A1(n14502), .A2(n14491), .ZN(n20571) );
  OR2_X2 U11313 ( .A1(n12924), .A2(n15187), .ZN(n12965) );
  AND2_X1 U11314 ( .A1(n16746), .A2(n11577), .ZN(n11023) );
  NAND2_X1 U11315 ( .A1(n12012), .A2(n12011), .ZN(n9914) );
  AOI21_X1 U11316 ( .B1(n16746), .B2(n11575), .A(n11574), .ZN(n13997) );
  NOR2_X2 U11317 ( .A1(n19431), .A2(n16809), .ZN(n19638) );
  NAND2_X1 U11318 ( .A1(n9950), .A2(n12521), .ZN(n12522) );
  OR2_X2 U11319 ( .A1(n16761), .A2(n19417), .ZN(n15957) );
  NOR2_X1 U11320 ( .A1(n13979), .A2(n14156), .ZN(n13978) );
  NAND2_X2 U11321 ( .A1(n9768), .A2(n12166), .ZN(n18658) );
  NOR2_X1 U11322 ( .A1(n13675), .A2(n14194), .ZN(n13835) );
  XNOR2_X1 U11323 ( .A(n10998), .B(n11296), .ZN(n10999) );
  CLKBUF_X1 U11324 ( .A(n10400), .Z(n19567) );
  NAND2_X1 U11325 ( .A1(n10982), .A2(n10981), .ZN(n11000) );
  NAND2_X1 U11326 ( .A1(n10988), .A2(n10987), .ZN(n11297) );
  NOR2_X2 U11327 ( .A1(n12150), .A2(n12149), .ZN(n13754) );
  AOI21_X1 U11328 ( .B1(n12164), .B2(n12163), .A(n12162), .ZN(n12168) );
  AND2_X1 U11329 ( .A1(n13330), .A2(n10244), .ZN(n10247) );
  AND3_X1 U11330 ( .A1(n9933), .A2(n9932), .A3(n11137), .ZN(n9930) );
  AND2_X1 U11331 ( .A1(n10950), .A2(n10949), .ZN(n10951) );
  INV_X2 U11332 ( .A(n14059), .ZN(n19566) );
  NOR2_X1 U11333 ( .A1(n12826), .A2(n12770), .ZN(n12805) );
  NAND2_X1 U11334 ( .A1(n14305), .A2(n14304), .ZN(n14296) );
  OR2_X1 U11335 ( .A1(n12428), .A2(n12544), .ZN(n12429) );
  NOR2_X1 U11336 ( .A1(n15540), .A2(n15004), .ZN(n10237) );
  CLKBUF_X1 U11337 ( .A(n10497), .Z(n14353) );
  AND2_X1 U11338 ( .A1(n13349), .A2(n13348), .ZN(n15004) );
  NAND2_X1 U11339 ( .A1(n10953), .A2(n10946), .ZN(n14214) );
  NOR2_X1 U11340 ( .A1(n13926), .A2(n12148), .ZN(n12149) );
  NAND2_X1 U11341 ( .A1(n12743), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12826) );
  NAND2_X1 U11342 ( .A1(n12502), .A2(n13193), .ZN(n12505) );
  NAND2_X2 U11343 ( .A1(n17039), .A2(n17042), .ZN(n18357) );
  OAI21_X1 U11344 ( .B1(n11935), .B2(n9913), .A(n9911), .ZN(n14114) );
  OR2_X1 U11345 ( .A1(n17863), .A2(n13665), .ZN(n12148) );
  AND3_X1 U11346 ( .A1(n12200), .A2(n13728), .A3(n12167), .ZN(n13667) );
  NAND3_X1 U11347 ( .A1(n12424), .A2(n12423), .A3(n12422), .ZN(n12436) );
  OR2_X1 U11348 ( .A1(n11096), .A2(n11095), .ZN(n11107) );
  AND2_X1 U11349 ( .A1(n13322), .A2(n13321), .ZN(n14304) );
  AND2_X1 U11350 ( .A1(n10881), .A2(n10880), .ZN(n10944) );
  AOI21_X1 U11351 ( .B1(n12193), .B2(n12192), .A(n12191), .ZN(n19180) );
  NAND2_X1 U11352 ( .A1(n12498), .A2(n12497), .ZN(n12675) );
  NOR2_X1 U11353 ( .A1(n12164), .A2(n12146), .ZN(n12169) );
  INV_X2 U11354 ( .A(n10688), .ZN(n10765) );
  NAND2_X1 U11355 ( .A1(n11087), .A2(n11086), .ZN(n11124) );
  NOR2_X1 U11356 ( .A1(n12151), .A2(n12100), .ZN(n12201) );
  NAND2_X1 U11357 ( .A1(n13312), .A2(n13311), .ZN(n13316) );
  INV_X1 U11358 ( .A(n10880), .ZN(n16864) );
  AND2_X1 U11359 ( .A1(n12381), .A2(n12380), .ZN(n13535) );
  NAND2_X1 U11360 ( .A1(n12544), .A2(n12543), .ZN(n13248) );
  OAI211_X1 U11361 ( .C1(n13243), .C2(n12501), .A(n12500), .B(n12499), .ZN(
        n12674) );
  NAND2_X1 U11362 ( .A1(n13900), .A2(n10947), .ZN(n10034) );
  CLKBUF_X1 U11363 ( .A(n13350), .Z(n14551) );
  OAI21_X1 U11364 ( .B1(n12189), .B2(n12185), .A(n12190), .ZN(n12196) );
  MUX2_X1 U11365 ( .A(n13317), .B(n14641), .S(P1_EBX_REG_1__SCAN_IN), .Z(
        n13312) );
  NAND2_X1 U11366 ( .A1(n12152), .A2(n18775), .ZN(n13930) );
  INV_X1 U11367 ( .A(n13485), .ZN(n9920) );
  AND2_X1 U11368 ( .A1(n18779), .A2(n18775), .ZN(n12158) );
  NAND2_X1 U11369 ( .A1(n12483), .A2(n13186), .ZN(n13193) );
  NAND2_X1 U11370 ( .A1(n10357), .A2(n10358), .ZN(n10912) );
  NAND2_X1 U11371 ( .A1(n13599), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16932) );
  AND2_X1 U11372 ( .A1(n11287), .A2(n10399), .ZN(n10947) );
  OR2_X1 U11373 ( .A1(n11936), .A2(n18122), .ZN(n11953) );
  OR2_X1 U11374 ( .A1(n12438), .A2(n12409), .ZN(n15582) );
  AND2_X1 U11375 ( .A1(n10358), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10355) );
  NOR2_X1 U11376 ( .A1(n13904), .A2(n10901), .ZN(n10883) );
  AND2_X1 U11378 ( .A1(n12142), .A2(n12141), .ZN(n12194) );
  AND2_X1 U11379 ( .A1(n12115), .A2(n12114), .ZN(n12154) );
  AND2_X1 U11380 ( .A1(n10902), .A2(n10901), .ZN(n10358) );
  AND2_X1 U11381 ( .A1(n13904), .A2(n10889), .ZN(n10357) );
  AND2_X1 U11382 ( .A1(n11932), .A2(n9683), .ZN(n18122) );
  INV_X1 U11383 ( .A(n10847), .ZN(n10849) );
  AND2_X1 U11384 ( .A1(n11949), .A2(n10411), .ZN(n18117) );
  AND2_X2 U11385 ( .A1(n14486), .A2(n12441), .ZN(n13324) );
  INV_X1 U11386 ( .A(n12543), .ZN(n12483) );
  OR2_X1 U11387 ( .A1(n12494), .A2(n12493), .ZN(n13158) );
  NOR2_X1 U11388 ( .A1(n12055), .A2(n12054), .ZN(n12061) );
  OR2_X1 U11389 ( .A1(n11915), .A2(n11914), .ZN(n13938) );
  XNOR2_X1 U11390 ( .A(n13934), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13885) );
  INV_X1 U11391 ( .A(n12408), .ZN(n12421) );
  OR2_X2 U11392 ( .A1(n12047), .A2(n12046), .ZN(n19335) );
  OR2_X1 U11393 ( .A1(n12482), .A2(n12481), .ZN(n13186) );
  CLKBUF_X3 U11394 ( .A(n12397), .Z(n14486) );
  AND2_X1 U11395 ( .A1(n20311), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13713) );
  INV_X2 U11396 ( .A(n12441), .ZN(n20603) );
  NAND4_X1 U11397 ( .A1(n12366), .A2(n12365), .A3(n12364), .A4(n12363), .ZN(
        n12397) );
  NAND3_X2 U11398 ( .A1(n12396), .A2(n12395), .A3(n12394), .ZN(n12441) );
  NAND2_X2 U11399 ( .A1(n10033), .A2(n10032), .ZN(n10838) );
  NAND2_X1 U11400 ( .A1(n9848), .A2(n9846), .ZN(n19619) );
  NAND2_X2 U11401 ( .A1(n12378), .A2(n12377), .ZN(n12408) );
  NAND4_X2 U11402 ( .A1(n12317), .A2(n12316), .A3(n12315), .A4(n12314), .ZN(
        n12406) );
  AND4_X1 U11403 ( .A1(n12376), .A2(n12375), .A3(n12374), .A4(n12373), .ZN(
        n12377) );
  AND4_X1 U11404 ( .A1(n12290), .A2(n12289), .A3(n12288), .A4(n12287), .ZN(
        n12296) );
  AND3_X1 U11405 ( .A1(n12338), .A2(n12337), .A3(n12336), .ZN(n12340) );
  OAI21_X1 U11406 ( .B1(n10281), .B2(n10280), .A(n10441), .ZN(n10279) );
  AND4_X1 U11407 ( .A1(n12313), .A2(n12312), .A3(n12311), .A4(n12310), .ZN(
        n12314) );
  NAND2_X1 U11408 ( .A1(n10031), .A2(n10441), .ZN(n10032) );
  AND3_X1 U11409 ( .A1(n12327), .A2(n12326), .A3(n12325), .ZN(n12328) );
  AND4_X1 U11410 ( .A1(n12113), .A2(n12112), .A3(n12111), .A4(n12110), .ZN(
        n12114) );
  AND4_X1 U11411 ( .A1(n12345), .A2(n12344), .A3(n12343), .A4(n12342), .ZN(
        n12366) );
  AND4_X1 U11412 ( .A1(n10091), .A2(n11904), .A3(n11898), .A4(n11901), .ZN(
        n10090) );
  AND3_X1 U11413 ( .A1(n12393), .A2(n12392), .A3(n12391), .ZN(n12394) );
  NAND2_X2 U11414 ( .A1(n19261), .A2(n21319), .ZN(n19311) );
  AND4_X1 U11415 ( .A1(n12294), .A2(n12293), .A3(n12292), .A4(n12291), .ZN(
        n12295) );
  AND4_X1 U11416 ( .A1(n12300), .A2(n12299), .A3(n12298), .A4(n12297), .ZN(
        n12317) );
  AND4_X1 U11417 ( .A1(n12387), .A2(n12386), .A3(n12385), .A4(n12384), .ZN(
        n12396) );
  INV_X2 U11418 ( .A(n10834), .ZN(n11675) );
  AND4_X1 U11419 ( .A1(n12323), .A2(n12322), .A3(n12321), .A4(n12320), .ZN(
        n12330) );
  AND4_X1 U11420 ( .A1(n12357), .A2(n12356), .A3(n12355), .A4(n12354), .ZN(
        n12364) );
  AND4_X1 U11421 ( .A1(n12308), .A2(n12307), .A3(n12306), .A4(n12305), .ZN(
        n12315) );
  CLKBUF_X3 U11422 ( .A(n12453), .Z(n13511) );
  CLKBUF_X3 U11423 ( .A(n12331), .Z(n13068) );
  CLKBUF_X2 U11424 ( .A(n13657), .Z(n17966) );
  AND2_X1 U11425 ( .A1(n11728), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n9777) );
  INV_X2 U11426 ( .A(n17348), .ZN(U215) );
  NAND2_X2 U11427 ( .A1(n20260), .A2(n20208), .ZN(n20258) );
  INV_X2 U11428 ( .A(n12117), .ZN(n17947) );
  AND2_X2 U11429 ( .A1(n14215), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10548) );
  AND2_X1 U11430 ( .A1(n11875), .A2(n19196), .ZN(n11921) );
  CLKBUF_X3 U11431 ( .A(n13110), .Z(n9604) );
  CLKBUF_X2 U11432 ( .A(n13658), .Z(n17834) );
  INV_X2 U11433 ( .A(n17350), .ZN(n17352) );
  NAND2_X2 U11434 ( .A1(n12279), .A2(n9787), .ZN(n13106) );
  BUF_X2 U11435 ( .A(n11960), .Z(n17953) );
  AND3_X1 U11436 ( .A1(n12170), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11875) );
  NOR4_X1 U11437 ( .A1(n16991), .A2(n18440), .A3(n18421), .A4(n18402), .ZN(
        n18352) );
  AND2_X1 U11438 ( .A1(n11877), .A2(n9689), .ZN(n11994) );
  AND2_X1 U11439 ( .A1(n13760), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n17094) );
  AND2_X1 U11440 ( .A1(n19196), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11884) );
  AND2_X2 U11441 ( .A1(n12271), .A2(n13951), .ZN(n13504) );
  INV_X1 U11442 ( .A(n9612), .ZN(n9590) );
  AND2_X2 U11443 ( .A1(n10234), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10082) );
  AND2_X1 U11444 ( .A1(n12269), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12279) );
  INV_X1 U11445 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14023) );
  INV_X1 U11446 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10234) );
  AND2_X1 U11447 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13784) );
  INV_X1 U11448 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13758) );
  NOR2_X2 U11449 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13785) );
  INV_X1 U11450 ( .A(n16351), .ZN(n11474) );
  NAND2_X1 U11451 ( .A1(n12402), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n9592) );
  INV_X1 U11452 ( .A(n10391), .ZN(n9593) );
  NOR2_X1 U11453 ( .A1(n14336), .A2(n14335), .ZN(n9594) );
  XNOR2_X1 U11454 ( .A(n14663), .B(n14662), .ZN(n9595) );
  XNOR2_X1 U11455 ( .A(n14663), .B(n14662), .ZN(n9596) );
  OAI211_X2 U11456 ( .C1(n13413), .C2(n13298), .A(n14480), .B(n14500), .ZN(
        n12402) );
  NAND2_X1 U11457 ( .A1(n14826), .A2(n14827), .ZN(n14812) );
  NOR2_X1 U11458 ( .A1(n14336), .A2(n14335), .ZN(n14437) );
  NAND2_X1 U11459 ( .A1(n14294), .A2(n14295), .ZN(n14336) );
  XNOR2_X1 U11460 ( .A(n12648), .B(n12647), .ZN(n13145) );
  XNOR2_X1 U11461 ( .A(n14663), .B(n14662), .ZN(n14664) );
  AND2_X1 U11462 ( .A1(n12520), .A2(n9722), .ZN(n9950) );
  AND2_X1 U11463 ( .A1(n12271), .A2(n13951), .ZN(n9597) );
  NOR2_X1 U11464 ( .A1(n12415), .A2(n12421), .ZN(n12381) );
  AND2_X2 U11465 ( .A1(n12270), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9787) );
  NOR2_X1 U11466 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12271) );
  NOR2_X1 U11467 ( .A1(n12681), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12278) );
  NOR2_X2 U11468 ( .A1(n12622), .A2(n12628), .ZN(n12623) );
  AND2_X2 U11469 ( .A1(n12277), .A2(n13968), .ZN(n9614) );
  AND2_X1 U11470 ( .A1(n12404), .A2(n12408), .ZN(n12439) );
  AND2_X1 U11471 ( .A1(n12408), .A2(n12417), .ZN(n13871) );
  NOR2_X2 U11472 ( .A1(n11772), .A2(n11771), .ZN(n15990) );
  NAND2_X2 U11473 ( .A1(n11049), .A2(n11048), .ZN(n16709) );
  CLKBUF_X1 U11476 ( .A(n9614), .Z(n9618) );
  CLKBUF_X1 U11477 ( .A(n9614), .Z(n9617) );
  CLKBUF_X1 U11478 ( .A(n9614), .Z(n9616) );
  AOI211_X2 U11479 ( .C1(P1_REIP_REG_4__SCAN_IN), .C2(n20436), .A(n20435), .B(
        n20434), .ZN(n20437) );
  AND2_X1 U11480 ( .A1(n10447), .A2(n16834), .ZN(n9598) );
  AND2_X1 U11481 ( .A1(n10447), .A2(n16834), .ZN(n9599) );
  NOR2_X2 U11482 ( .A1(n14503), .A2(n10236), .ZN(n14909) );
  NOR2_X1 U11483 ( .A1(n17362), .A2(n19335), .ZN(n18493) );
  AND2_X2 U11484 ( .A1(n10832), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14215) );
  NAND2_X1 U11485 ( .A1(n16961), .A2(n13595), .ZN(n16962) );
  NOR2_X2 U11486 ( .A1(n17632), .A2(n18367), .ZN(n16961) );
  OAI222_X1 U11487 ( .A1(n15011), .A2(n14664), .B1(n14976), .B2(n20447), .C1(
        n15323), .C2(n15013), .ZN(P1_U2842) );
  NOR2_X2 U11488 ( .A1(n14296), .A2(n10246), .ZN(n14449) );
  AND4_X1 U11489 ( .A1(n12335), .A2(n12334), .A3(n12333), .A4(n12332), .ZN(
        n12341) );
  XNOR2_X2 U11490 ( .A(n13297), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14583) );
  NOR2_X2 U11491 ( .A1(n13501), .A2(n15109), .ZN(n13297) );
  AND2_X4 U11492 ( .A1(n20635), .A2(n12521), .ZN(n10366) );
  NAND2_X2 U11493 ( .A1(n12449), .A2(n12450), .ZN(n20635) );
  AND2_X1 U11494 ( .A1(n10447), .A2(n16834), .ZN(n9602) );
  AND2_X1 U11495 ( .A1(n10447), .A2(n16834), .ZN(n9603) );
  AND2_X1 U11496 ( .A1(n11012), .A2(n11013), .ZN(n16822) );
  AND2_X1 U11497 ( .A1(n11012), .A2(n11024), .ZN(n20128) );
  NOR4_X2 U11498 ( .A1(n14193), .A2(n17604), .A3(n17995), .A4(n13670), .ZN(
        n13671) );
  BUF_X2 U11499 ( .A(n13110), .Z(n9605) );
  AOI22_X1 U11500 ( .A1(n12452), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9610), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12332) );
  AND2_X4 U11501 ( .A1(n10082), .A2(n9787), .ZN(n12720) );
  INV_X2 U11502 ( .A(n12407), .ZN(n12403) );
  XNOR2_X2 U11503 ( .A(n10978), .B(n10977), .ZN(n10277) );
  AND2_X1 U11504 ( .A1(n12277), .A2(n10082), .ZN(n9606) );
  NAND2_X2 U11505 ( .A1(n9898), .A2(n10951), .ZN(n10977) );
  AND2_X1 U11506 ( .A1(n11014), .A2(n11024), .ZN(n19980) );
  NOR2_X1 U11507 ( .A1(n12401), .A2(n12414), .ZN(n13950) );
  NAND2_X1 U11508 ( .A1(n10988), .A2(n10987), .ZN(n9608) );
  AND2_X1 U11509 ( .A1(n11014), .A2(n11015), .ZN(n19918) );
  AND3_X1 U11510 ( .A1(n14486), .A2(n12406), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n13260) );
  NAND2_X1 U11511 ( .A1(n12402), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n9866) );
  NAND2_X1 U11512 ( .A1(n13772), .A2(n10838), .ZN(n10730) );
  NAND2_X1 U11513 ( .A1(n10472), .A2(n10838), .ZN(n10906) );
  NAND2_X2 U11514 ( .A1(n14770), .A2(n14772), .ZN(n14749) );
  INV_X2 U11515 ( .A(n10838), .ZN(n10902) );
  OAI21_X1 U11516 ( .B1(n11567), .B2(n13712), .A(n11566), .ZN(n11591) );
  AND2_X1 U11517 ( .A1(n12278), .A2(n13951), .ZN(n9609) );
  AND2_X1 U11518 ( .A1(n12278), .A2(n13951), .ZN(n9610) );
  INV_X1 U11519 ( .A(n9589), .ZN(n9623) );
  NOR2_X2 U11521 ( .A1(n14830), .A2(n14814), .ZN(n14806) );
  NOR2_X2 U11522 ( .A1(n15810), .A2(n13585), .ZN(n13584) );
  AOI21_X2 U11523 ( .B1(n12437), .B2(n14937), .A(n20383), .ZN(n20433) );
  INV_X2 U11524 ( .A(n20393), .ZN(n20383) );
  AND2_X2 U11525 ( .A1(n10082), .A2(n12276), .ZN(n12469) );
  AND2_X1 U11526 ( .A1(n10832), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9612) );
  XNOR2_X1 U11527 ( .A(n10065), .B(n9924), .ZN(n11006) );
  NOR2_X2 U11528 ( .A1(n18478), .A2(n18368), .ZN(n18455) );
  INV_X4 U11529 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n16834) );
  CLKBUF_X1 U11530 ( .A(n13505), .Z(n9620) );
  CLKBUF_X1 U11531 ( .A(n13505), .Z(n9621) );
  INV_X1 U11532 ( .A(n9589), .ZN(n9624) );
  INV_X1 U11533 ( .A(n11846), .ZN(n9625) );
  INV_X1 U11534 ( .A(n11846), .ZN(n9626) );
  NOR2_X4 U11535 ( .A1(n14675), .A2(n10393), .ZN(n14662) );
  XNOR2_X1 U11536 ( .A(n13316), .B(n13909), .ZN(n14149) );
  NOR4_X2 U11537 ( .A1(n15220), .A2(n15233), .A3(n15231), .A4(n15234), .ZN(
        n15222) );
  NAND2_X4 U11538 ( .A1(n13310), .A2(n13324), .ZN(n13317) );
  AND2_X1 U11539 ( .A1(n11451), .A2(n10884), .ZN(n9627) );
  NAND2_X4 U11540 ( .A1(n10267), .A2(n10266), .ZN(n10884) );
  INV_X1 U11541 ( .A(n9853), .ZN(n9859) );
  AOI21_X1 U11542 ( .B1(n10076), .B2(n10078), .A(n10075), .ZN(n10074) );
  INV_X1 U11543 ( .A(n16290), .ZN(n10075) );
  INV_X1 U11544 ( .A(n10079), .ZN(n10076) );
  AND4_X1 U11545 ( .A1(n10603), .A2(n10602), .A3(n10601), .A4(n10600), .ZN(
        n10611) );
  NAND2_X1 U11546 ( .A1(n16864), .A2(n10952), .ZN(n10987) );
  NAND3_X1 U11547 ( .A1(n9921), .A2(n10849), .A3(n9668), .ZN(n13485) );
  AND2_X1 U11548 ( .A1(n10848), .A2(n20311), .ZN(n9921) );
  INV_X1 U11549 ( .A(n16970), .ZN(n12015) );
  NAND2_X1 U11550 ( .A1(n12407), .A2(n20607), .ZN(n13154) );
  NAND2_X1 U11551 ( .A1(n10882), .A2(n10903), .ZN(n10061) );
  AND4_X1 U11552 ( .A1(n10819), .A2(n10818), .A3(n10817), .A4(n10816), .ZN(
        n10820) );
  NAND2_X1 U11553 ( .A1(n11697), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n9802) );
  NAND2_X1 U11554 ( .A1(n13127), .A2(n10397), .ZN(n10396) );
  INV_X1 U11555 ( .A(n14677), .ZN(n10397) );
  NAND2_X1 U11556 ( .A1(n10386), .A2(n14721), .ZN(n10385) );
  INV_X1 U11557 ( .A(n10388), .ZN(n10386) );
  OAI21_X2 U11558 ( .B1(n10382), .B2(n9796), .A(n9793), .ZN(n9797) );
  INV_X1 U11559 ( .A(n15335), .ZN(n9796) );
  NAND2_X1 U11560 ( .A1(n14537), .A2(n9763), .ZN(n9793) );
  NAND2_X1 U11561 ( .A1(n10379), .A2(n10380), .ZN(n10142) );
  INV_X1 U11562 ( .A(n14881), .ZN(n10243) );
  INV_X1 U11563 ( .A(n20571), .ZN(n15401) );
  OAI211_X1 U11564 ( .C1(n13018), .C2(n13243), .A(n12504), .B(n12503), .ZN(
        n12506) );
  NAND2_X1 U11565 ( .A1(n9852), .A2(n11777), .ZN(n11778) );
  NAND2_X1 U11566 ( .A1(n10300), .A2(n9734), .ZN(n9853) );
  INV_X1 U11567 ( .A(n11775), .ZN(n14241) );
  INV_X1 U11568 ( .A(n9881), .ZN(n9879) );
  NAND2_X1 U11569 ( .A1(n9927), .A2(n9928), .ZN(n9925) );
  INV_X1 U11570 ( .A(n10132), .ZN(n9927) );
  INV_X1 U11571 ( .A(n11414), .ZN(n9928) );
  NAND2_X1 U11572 ( .A1(n9810), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9809) );
  NAND2_X1 U11573 ( .A1(n10472), .A2(n10901), .ZN(n9779) );
  AND2_X2 U11574 ( .A1(n14111), .A2(n9613), .ZN(n11026) );
  NAND2_X1 U11575 ( .A1(n17100), .A2(n13608), .ZN(n13721) );
  NOR2_X1 U11576 ( .A1(n17251), .A2(n17412), .ZN(n17250) );
  NAND2_X1 U11577 ( .A1(n16877), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17251) );
  AND2_X1 U11578 ( .A1(n11993), .A2(n11992), .ZN(n17039) );
  NAND2_X1 U11579 ( .A1(n14536), .A2(n10374), .ZN(n15130) );
  INV_X1 U11580 ( .A(n15185), .ZN(n10375) );
  NAND2_X1 U11581 ( .A1(n20662), .A2(n21384), .ZN(n20926) );
  OR2_X1 U11582 ( .A1(n20662), .A2(n21384), .ZN(n20959) );
  NOR2_X1 U11583 ( .A1(n16346), .A2(n10185), .ZN(n10184) );
  INV_X1 U11584 ( .A(n16359), .ZN(n10185) );
  AND2_X1 U11585 ( .A1(n9693), .A2(n11590), .ZN(n10293) );
  NOR2_X1 U11586 ( .A1(n10889), .A2(n13438), .ZN(n13770) );
  AND2_X1 U11587 ( .A1(n13486), .A2(n13630), .ZN(n13633) );
  NAND2_X1 U11588 ( .A1(n9714), .A2(n16301), .ZN(n10078) );
  INV_X1 U11589 ( .A(n16300), .ZN(n10080) );
  INV_X1 U11590 ( .A(n10354), .ZN(n10107) );
  INV_X1 U11591 ( .A(n11296), .ZN(n10320) );
  NAND2_X1 U11592 ( .A1(n11397), .A2(n9843), .ZN(n11398) );
  INV_X1 U11593 ( .A(n9844), .ZN(n9843) );
  NAND2_X1 U11594 ( .A1(n15632), .A2(n9740), .ZN(n11479) );
  NOR2_X1 U11595 ( .A1(n11422), .A2(n10318), .ZN(n10316) );
  INV_X1 U11596 ( .A(n11445), .ZN(n10318) );
  AND2_X1 U11597 ( .A1(n11276), .A2(n11417), .ZN(n11277) );
  NAND2_X1 U11598 ( .A1(n10134), .A2(n9977), .ZN(n11278) );
  NOR2_X1 U11599 ( .A1(n15626), .A2(n16378), .ZN(n11415) );
  AND2_X1 U11600 ( .A1(n9677), .A2(n16627), .ZN(n10126) );
  AND2_X1 U11601 ( .A1(n10353), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10352) );
  INV_X1 U11602 ( .A(n10337), .ZN(n10336) );
  NAND2_X1 U11603 ( .A1(n10432), .A2(n10441), .ZN(n10267) );
  INV_X1 U11604 ( .A(n12196), .ZN(n19185) );
  INV_X1 U11605 ( .A(n16880), .ZN(n17042) );
  NOR2_X1 U11606 ( .A1(n10098), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10097) );
  INV_X1 U11607 ( .A(n10415), .ZN(n10098) );
  NOR2_X1 U11608 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n12207), .ZN(n19214) );
  OR2_X1 U11609 ( .A1(n21134), .A2(n10368), .ZN(n20330) );
  OR2_X1 U11610 ( .A1(n13896), .A2(n13629), .ZN(n20309) );
  OAI21_X1 U11611 ( .B1(n11525), .B2(n15911), .A(n9742), .ZN(n10122) );
  NAND2_X1 U11612 ( .A1(n11434), .A2(n11433), .ZN(n11435) );
  NAND2_X1 U11613 ( .A1(n16097), .A2(n17215), .ZN(n11434) );
  OR2_X1 U11614 ( .A1(n9984), .A2(n9690), .ZN(n9981) );
  NOR2_X1 U11615 ( .A1(n17031), .A2(n13765), .ZN(n9917) );
  OR2_X1 U11616 ( .A1(n12535), .A2(n12534), .ZN(n12536) );
  AOI21_X1 U11617 ( .B1(n13043), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A(
        n10154), .ZN(n12562) );
  AND2_X1 U11618 ( .A1(n12353), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n10154) );
  NAND2_X1 U11619 ( .A1(n13240), .A2(n13221), .ZN(n13255) );
  AOI21_X1 U11620 ( .B1(n9607), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A(
        n10170), .ZN(n12915) );
  AND2_X1 U11621 ( .A1(n10147), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n10170) );
  AOI21_X1 U11622 ( .B1(n13043), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n10153), .ZN(n12889) );
  AND2_X1 U11623 ( .A1(n10147), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n10153) );
  AOI21_X1 U11624 ( .B1(n13068), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A(
        n10172), .ZN(n12837) );
  AND2_X1 U11625 ( .A1(n10147), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n10172) );
  NAND2_X1 U11626 ( .A1(n9632), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10006) );
  AOI21_X1 U11627 ( .B1(n9569), .B2(n10378), .A(n10373), .ZN(n10372) );
  INV_X1 U11628 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n10373) );
  NOR2_X1 U11629 ( .A1(n9952), .A2(n10143), .ZN(n9943) );
  AND2_X1 U11630 ( .A1(n12353), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10155) );
  AOI21_X1 U11631 ( .B1(n12461), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A(
        n10162), .ZN(n12580) );
  NAND2_X1 U11632 ( .A1(n12353), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12355) );
  INV_X1 U11633 ( .A(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12347) );
  AND2_X1 U11634 ( .A1(n12353), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n10160) );
  INV_X1 U11635 ( .A(n13260), .ZN(n13243) );
  AND2_X1 U11636 ( .A1(n10149), .A2(n10148), .ZN(n12455) );
  NAND2_X1 U11637 ( .A1(n12353), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10149) );
  NAND2_X1 U11638 ( .A1(n13068), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10148) );
  MUX2_X1 U11639 ( .A(n12504), .B(n13193), .S(n12495), .Z(n12498) );
  INV_X1 U11640 ( .A(n9592), .ZN(n10056) );
  AND2_X1 U11641 ( .A1(n13255), .A2(n13254), .ZN(n13257) );
  INV_X1 U11642 ( .A(n13300), .ZN(n13247) );
  INV_X1 U11643 ( .A(n13301), .ZN(n13237) );
  NAND2_X1 U11644 ( .A1(n12427), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12544) );
  OAI21_X1 U11645 ( .B1(n11390), .B2(n20226), .A(n11328), .ZN(n9830) );
  INV_X1 U11646 ( .A(n11165), .ZN(n10338) );
  OR2_X1 U11647 ( .A1(n10555), .A2(n10554), .ZN(n11093) );
  NAND2_X1 U11648 ( .A1(n13904), .A2(n20306), .ZN(n10526) );
  AND2_X1 U11649 ( .A1(n13905), .A2(n13772), .ZN(n10516) );
  NAND2_X1 U11650 ( .A1(n10906), .A2(n19619), .ZN(n10891) );
  AND4_X1 U11651 ( .A1(n9727), .A2(n9800), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A4(n10812), .ZN(n9799) );
  NOR2_X1 U11652 ( .A1(n10344), .A2(n9695), .ZN(n10343) );
  NAND2_X1 U11653 ( .A1(n11699), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10124) );
  AND3_X1 U11654 ( .A1(n9959), .A2(n9958), .A3(n9957), .ZN(n10342) );
  NAND2_X1 U11655 ( .A1(n11700), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n9959) );
  NAND2_X1 U11656 ( .A1(n11694), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n9958) );
  NAND2_X1 U11657 ( .A1(n11697), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n9957) );
  AND2_X1 U11658 ( .A1(n19682), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10782) );
  NAND2_X1 U11659 ( .A1(n10796), .A2(n10795), .ZN(n10801) );
  AND2_X1 U11660 ( .A1(n11973), .A2(n12218), .ZN(n11993) );
  NAND2_X1 U11661 ( .A1(n10390), .A2(n14786), .ZN(n10389) );
  INV_X1 U11662 ( .A(n10392), .ZN(n10390) );
  OR2_X1 U11663 ( .A1(n14800), .A2(n14813), .ZN(n10392) );
  INV_X1 U11664 ( .A(n13078), .ZN(n13528) );
  NAND2_X1 U11665 ( .A1(n14024), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13078) );
  XNOR2_X1 U11666 ( .A(n12611), .B(n12610), .ZN(n13130) );
  INV_X1 U11667 ( .A(n12609), .ZN(n12610) );
  NAND2_X1 U11668 ( .A1(n14537), .A2(n14563), .ZN(n14539) );
  INV_X1 U11669 ( .A(n20416), .ZN(n10244) );
  NAND2_X1 U11670 ( .A1(n12611), .A2(n12609), .ZN(n12621) );
  AND2_X1 U11671 ( .A1(n12609), .A2(n12619), .ZN(n9814) );
  NAND2_X1 U11672 ( .A1(n10139), .A2(n9739), .ZN(n10145) );
  NAND2_X1 U11673 ( .A1(n13135), .A2(n13858), .ZN(n10139) );
  NAND2_X1 U11674 ( .A1(n12419), .A2(n12418), .ZN(n12423) );
  AND2_X1 U11675 ( .A1(n13350), .A2(n12415), .ZN(n13864) );
  OAI21_X1 U11676 ( .B1(n17115), .B2(n14470), .A(n20607), .ZN(n10020) );
  NAND2_X1 U11677 ( .A1(n14474), .A2(n12401), .ZN(n10019) );
  OR2_X1 U11678 ( .A1(n12557), .A2(n12556), .ZN(n13140) );
  AND2_X1 U11679 ( .A1(n13880), .A2(n13879), .ZN(n17117) );
  NAND2_X1 U11680 ( .A1(n12542), .A2(n12541), .ZN(n20724) );
  XNOR2_X1 U11681 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10786) );
  NOR2_X1 U11682 ( .A1(n10225), .A2(n11287), .ZN(n9929) );
  OAI21_X1 U11683 ( .B1(n11390), .B2(n17201), .A(n10996), .ZN(n9828) );
  NOR2_X1 U11684 ( .A1(n15954), .A2(n16773), .ZN(n15939) );
  MUX2_X1 U11685 ( .A(n11084), .B(n15947), .S(n11287), .Z(n11114) );
  INV_X1 U11686 ( .A(n11083), .ZN(n11084) );
  NAND2_X1 U11687 ( .A1(n13770), .A2(n15992), .ZN(n11775) );
  NAND2_X1 U11688 ( .A1(n10750), .A2(n10259), .ZN(n10258) );
  INV_X1 U11689 ( .A(n15664), .ZN(n10259) );
  INV_X1 U11690 ( .A(n10420), .ZN(n10295) );
  NOR2_X1 U11691 ( .A1(n10298), .A2(n16041), .ZN(n10297) );
  INV_X1 U11692 ( .A(n16034), .ZN(n10298) );
  NAND2_X1 U11693 ( .A1(n10261), .A2(n10702), .ZN(n10260) );
  INV_X1 U11694 ( .A(n15795), .ZN(n10261) );
  AND2_X1 U11695 ( .A1(n10630), .A2(n13894), .ZN(n10254) );
  INV_X1 U11696 ( .A(n13943), .ZN(n10630) );
  OAI21_X1 U11697 ( .B1(n9820), .B2(n11386), .A(n11384), .ZN(n9840) );
  NOR2_X1 U11698 ( .A1(n13469), .A2(n15654), .ZN(n13472) );
  INV_X1 U11699 ( .A(n15745), .ZN(n11180) );
  NAND2_X1 U11700 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n10109) );
  AND2_X1 U11701 ( .A1(n10115), .A2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10113) );
  NOR2_X1 U11702 ( .A1(n17199), .A2(n10112), .ZN(n10115) );
  NOR2_X1 U11703 ( .A1(n10513), .A2(n10512), .ZN(n11038) );
  INV_X1 U11704 ( .A(n15622), .ZN(n10317) );
  NAND2_X1 U11705 ( .A1(n10276), .A2(n15595), .ZN(n10275) );
  INV_X1 U11706 ( .A(n11426), .ZN(n10276) );
  OAI21_X1 U11707 ( .B1(n9820), .B2(n11377), .A(n11375), .ZN(n9842) );
  NAND2_X1 U11708 ( .A1(n16250), .A2(n10129), .ZN(n10134) );
  AND2_X1 U11709 ( .A1(n15706), .A2(n15688), .ZN(n10324) );
  OAI21_X1 U11710 ( .B1(n9820), .B2(n20241), .A(n11356), .ZN(n9838) );
  OR2_X1 U11711 ( .A1(n10314), .A2(n10313), .ZN(n10312) );
  INV_X1 U11712 ( .A(n11503), .ZN(n10313) );
  OAI21_X1 U11713 ( .B1(n9820), .B2(n20233), .A(n11342), .ZN(n9836) );
  NAND2_X1 U11714 ( .A1(n10315), .A2(n11345), .ZN(n10314) );
  INV_X1 U11715 ( .A(n15783), .ZN(n11345) );
  INV_X1 U11716 ( .A(n16049), .ZN(n10315) );
  OAI21_X1 U11717 ( .B1(n9820), .B2(n11340), .A(n11338), .ZN(n9826) );
  NAND2_X1 U11718 ( .A1(n14282), .A2(n14284), .ZN(n13587) );
  OAI21_X1 U11719 ( .B1(n11390), .B2(n16343), .A(n11324), .ZN(n9824) );
  AOI21_X1 U11720 ( .B1(n10347), .B2(n10349), .A(n10039), .ZN(n9786) );
  NAND2_X1 U11721 ( .A1(n9785), .A2(n10347), .ZN(n9784) );
  AND2_X1 U11722 ( .A1(n9646), .A2(n9748), .ZN(n10028) );
  AND2_X1 U11723 ( .A1(n10862), .A2(n10861), .ZN(n10918) );
  INV_X1 U11724 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9969) );
  NAND2_X1 U11725 ( .A1(n10855), .A2(n10854), .ZN(n9780) );
  INV_X1 U11726 ( .A(n11013), .ZN(n10345) );
  AND2_X1 U11727 ( .A1(n11582), .A2(n11581), .ZN(n19738) );
  NAND2_X1 U11728 ( .A1(n10806), .A2(n10805), .ZN(n10827) );
  OR2_X1 U11729 ( .A1(n10804), .A2(n10803), .ZN(n10806) );
  INV_X1 U11730 ( .A(n18306), .ZN(n10204) );
  OAI21_X1 U11731 ( .B1(n12117), .B2(n13847), .A(n10096), .ZN(n11874) );
  NAND2_X1 U11732 ( .A1(n17948), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n10096) );
  NAND2_X1 U11733 ( .A1(n18456), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17632) );
  NOR2_X1 U11734 ( .A1(n13978), .A2(n12239), .ZN(n12243) );
  NOR2_X1 U11735 ( .A1(n18463), .A2(n18699), .ZN(n9995) );
  NAND2_X1 U11736 ( .A1(n12224), .A2(n13934), .ZN(n11936) );
  XNOR2_X1 U11737 ( .A(n12224), .B(n13934), .ZN(n11918) );
  AND2_X1 U11738 ( .A1(n12154), .A2(n12194), .ZN(n13753) );
  NAND2_X1 U11739 ( .A1(n12165), .A2(n12168), .ZN(n13751) );
  NAND2_X1 U11740 ( .A1(n17948), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n9968) );
  NOR2_X1 U11741 ( .A1(n9963), .A2(n9962), .ZN(n9961) );
  INV_X1 U11742 ( .A(n12066), .ZN(n9963) );
  INV_X1 U11743 ( .A(n12067), .ZN(n9962) );
  AND2_X1 U11744 ( .A1(n19168), .A2(n19167), .ZN(n19191) );
  XNOR2_X1 U11745 ( .A(n13881), .B(n20724), .ZN(n13962) );
  NOR2_X1 U11746 ( .A1(n14939), .A2(n12427), .ZN(n13424) );
  AND2_X1 U11747 ( .A1(n10250), .A2(n10249), .ZN(n10248) );
  INV_X1 U11748 ( .A(n14691), .ZN(n10249) );
  OR2_X1 U11749 ( .A1(n15076), .A2(n14468), .ZN(n14016) );
  INV_X1 U11750 ( .A(n20330), .ZN(n14077) );
  OR2_X1 U11751 ( .A1(n13296), .A2(n13427), .ZN(n13501) );
  INV_X1 U11752 ( .A(n10395), .ZN(n10393) );
  NAND2_X1 U11753 ( .A1(n13101), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13296) );
  NAND2_X1 U11754 ( .A1(n13056), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13099) );
  NAND2_X1 U11755 ( .A1(n12899), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12923) );
  INV_X1 U11756 ( .A(n15002), .ZN(n12719) );
  INV_X1 U11757 ( .A(n14849), .ZN(n14925) );
  NAND2_X1 U11758 ( .A1(n9874), .A2(n12688), .ZN(n14295) );
  NAND2_X1 U11759 ( .A1(n14146), .A2(n14145), .ZN(n14302) );
  OR2_X1 U11760 ( .A1(n17115), .A2(n14645), .ZN(n17128) );
  NAND2_X1 U11761 ( .A1(n9795), .A2(n9797), .ZN(n9794) );
  INV_X1 U11762 ( .A(n14536), .ZN(n9795) );
  INV_X1 U11763 ( .A(n10142), .ZN(n10140) );
  NAND2_X1 U11764 ( .A1(n10382), .A2(n14539), .ZN(n15120) );
  NAND2_X1 U11765 ( .A1(n13210), .A2(n10377), .ZN(n10371) );
  NAND2_X1 U11766 ( .A1(n13381), .A2(n15175), .ZN(n10376) );
  INV_X1 U11767 ( .A(n15203), .ZN(n10010) );
  INV_X1 U11768 ( .A(n15183), .ZN(n13210) );
  NAND2_X1 U11769 ( .A1(n15203), .A2(n15202), .ZN(n15183) );
  NOR2_X1 U11770 ( .A1(n10242), .A2(n9639), .ZN(n10239) );
  NAND2_X1 U11771 ( .A1(n14927), .A2(n10237), .ZN(n10236) );
  INV_X1 U11772 ( .A(n20526), .ZN(n15267) );
  INV_X1 U11773 ( .A(n10366), .ZN(n14959) );
  NOR2_X1 U11774 ( .A1(n14485), .A2(n13870), .ZN(n14022) );
  INV_X1 U11775 ( .A(n20585), .ZN(n20587) );
  NOR2_X1 U11776 ( .A1(n20729), .A2(n20590), .ZN(n20898) );
  NOR2_X1 U11777 ( .A1(n20730), .A2(n20729), .ZN(n21027) );
  INV_X1 U11778 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21069) );
  INV_X1 U11779 ( .A(n20893), .ZN(n21016) );
  AOI21_X1 U11780 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20988), .A(n20729), 
        .ZN(n21080) );
  OAI21_X1 U11781 ( .B1(n13477), .B2(n9645), .A(n10186), .ZN(n14603) );
  INV_X1 U11782 ( .A(n10187), .ZN(n10186) );
  OAI22_X1 U11783 ( .A1(n16761), .A2(n15600), .B1(n9645), .B2(n16761), .ZN(
        n10187) );
  NAND2_X1 U11784 ( .A1(n16210), .A2(n15615), .ZN(n10189) );
  NAND2_X1 U11785 ( .A1(n13477), .A2(n16761), .ZN(n15623) );
  NAND2_X1 U11786 ( .A1(n16761), .A2(n13465), .ZN(n15677) );
  NAND2_X1 U11787 ( .A1(n9936), .A2(n11260), .ZN(n11235) );
  NOR2_X1 U11788 ( .A1(n9658), .A2(n11504), .ZN(n13462) );
  NAND2_X1 U11789 ( .A1(n15846), .A2(n10184), .ZN(n15814) );
  NAND2_X1 U11790 ( .A1(n15939), .A2(n15941), .ZN(n15928) );
  NAND2_X1 U11791 ( .A1(n10940), .A2(n9701), .ZN(n9971) );
  NAND2_X1 U11792 ( .A1(n11368), .A2(n9831), .ZN(n11370) );
  INV_X1 U11793 ( .A(n9832), .ZN(n9831) );
  OR2_X1 U11794 ( .A1(n10641), .A2(n10640), .ZN(n11594) );
  AND3_X1 U11795 ( .A1(n10267), .A2(n10266), .A3(n20306), .ZN(n13772) );
  NOR2_X1 U11796 ( .A1(n10275), .A2(n9755), .ZN(n10274) );
  AND2_X1 U11797 ( .A1(n10274), .A2(n10272), .ZN(n10271) );
  INV_X1 U11798 ( .A(n10769), .ZN(n10272) );
  AOI21_X2 U11799 ( .B1(n15985), .B2(n11812), .A(n11830), .ZN(n15976) );
  INV_X1 U11800 ( .A(n16006), .ZN(n10303) );
  OR2_X1 U11801 ( .A1(n16006), .A2(n16014), .ZN(n10302) );
  INV_X1 U11802 ( .A(n11717), .ZN(n10301) );
  OR2_X1 U11803 ( .A1(n16012), .A2(n16014), .ZN(n10304) );
  INV_X1 U11804 ( .A(n16022), .ZN(n9964) );
  NAND2_X1 U11805 ( .A1(n11591), .A2(n11570), .ZN(n14341) );
  NOR2_X1 U11806 ( .A1(n11487), .A2(n10222), .ZN(n10221) );
  NAND2_X1 U11807 ( .A1(n13479), .A2(n9650), .ZN(n11526) );
  AND2_X1 U11808 ( .A1(n13479), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13478) );
  AND2_X1 U11809 ( .A1(n13472), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13479) );
  AND2_X1 U11810 ( .A1(n16301), .A2(n16312), .ZN(n10079) );
  NAND2_X1 U11811 ( .A1(n11311), .A2(n9833), .ZN(n11312) );
  INV_X1 U11812 ( .A(n9834), .ZN(n9833) );
  NOR2_X1 U11813 ( .A1(n13446), .A2(n16420), .ZN(n13448) );
  NAND2_X1 U11814 ( .A1(n11299), .A2(n9821), .ZN(n11301) );
  INV_X1 U11815 ( .A(n9822), .ZN(n9821) );
  NAND2_X1 U11816 ( .A1(n11392), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n9845) );
  NAND2_X1 U11817 ( .A1(n9881), .A2(n9883), .ZN(n9880) );
  NOR2_X1 U11818 ( .A1(n9879), .A2(n9670), .ZN(n9878) );
  INV_X1 U11819 ( .A(n16248), .ZN(n9891) );
  INV_X1 U11820 ( .A(n16253), .ZN(n9893) );
  INV_X1 U11821 ( .A(n11218), .ZN(n9895) );
  AOI21_X1 U11822 ( .B1(n15710), .B2(n11293), .A(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16270) );
  OAI21_X1 U11823 ( .B1(n11231), .B2(n16378), .A(n16548), .ZN(n11536) );
  NAND2_X1 U11824 ( .A1(n10072), .A2(n10071), .ZN(n11497) );
  AOI21_X1 U11825 ( .B1(n10074), .B2(n10077), .A(n9712), .ZN(n10071) );
  NAND2_X1 U11826 ( .A1(n16314), .A2(n16312), .ZN(n10081) );
  AND2_X1 U11827 ( .A1(n11331), .A2(n11327), .ZN(n10325) );
  NAND2_X1 U11828 ( .A1(n9902), .A2(n10339), .ZN(n9901) );
  OAI21_X1 U11829 ( .B1(n10347), .B2(n10039), .A(n11552), .ZN(n10038) );
  NAND3_X1 U11830 ( .A1(n10100), .A2(n10989), .A3(n10099), .ZN(n11001) );
  NAND2_X1 U11831 ( .A1(n11392), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n10100) );
  NAND2_X1 U11832 ( .A1(n10103), .A2(n10101), .ZN(n10065) );
  NAND2_X1 U11833 ( .A1(n10102), .A2(n10978), .ZN(n10101) );
  OAI21_X1 U11834 ( .B1(n11577), .B2(n13712), .A(n11576), .ZN(n11578) );
  INV_X1 U11835 ( .A(n11573), .ZN(n11574) );
  NAND2_X1 U11836 ( .A1(n14232), .A2(n14231), .ZN(n16836) );
  AND2_X1 U11837 ( .A1(n16821), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19845) );
  NOR2_X2 U11838 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20305) );
  NAND2_X1 U11839 ( .A1(n20288), .A2(n20275), .ZN(n19914) );
  NAND2_X1 U11840 ( .A1(n19598), .A2(n20275), .ZN(n20043) );
  NAND2_X1 U11841 ( .A1(n9773), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9772) );
  NAND2_X1 U11842 ( .A1(n9775), .A2(n9910), .ZN(n9774) );
  INV_X1 U11843 ( .A(n19910), .ZN(n20037) );
  AND2_X1 U11844 ( .A1(n17407), .A2(n17388), .ZN(n17399) );
  NAND2_X1 U11845 ( .A1(n10202), .A2(n18288), .ZN(n10201) );
  NAND2_X1 U11846 ( .A1(n10203), .A2(n10204), .ZN(n10202) );
  XNOR2_X1 U11847 ( .A(n13601), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16881) );
  NAND2_X1 U11848 ( .A1(n17250), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13601) );
  AND2_X1 U11849 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11887) );
  NAND2_X1 U11850 ( .A1(n13721), .A2(n9688), .ZN(n9956) );
  OR2_X1 U11851 ( .A1(n19335), .A2(n18755), .ZN(n13926) );
  NAND2_X1 U11852 ( .A1(n12201), .A2(n12145), .ZN(n18175) );
  AND2_X1 U11853 ( .A1(n12200), .A2(n12144), .ZN(n12145) );
  NOR2_X1 U11854 ( .A1(n16962), .A2(n10214), .ZN(n10213) );
  NAND2_X1 U11855 ( .A1(n10215), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10214) );
  INV_X1 U11856 ( .A(n10216), .ZN(n10215) );
  NOR2_X1 U11857 ( .A1(n16962), .A2(n10216), .ZN(n18301) );
  NOR2_X1 U11858 ( .A1(n16962), .A2(n16966), .ZN(n18338) );
  OR2_X1 U11859 ( .A1(n18373), .A2(n18354), .ZN(n16965) );
  NOR2_X1 U11860 ( .A1(n14250), .A2(n12248), .ZN(n18407) );
  XNOR2_X1 U11861 ( .A(n12249), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16883) );
  AND2_X1 U11862 ( .A1(n18365), .A2(n9764), .ZN(n10095) );
  NAND2_X1 U11863 ( .A1(n9992), .A2(n9990), .ZN(n16970) );
  AND2_X1 U11864 ( .A1(n16979), .A2(n9991), .ZN(n9990) );
  NAND2_X1 U11865 ( .A1(n18357), .A2(n9757), .ZN(n9991) );
  OR2_X1 U11866 ( .A1(n19183), .A2(n17042), .ZN(n18524) );
  AND2_X1 U11867 ( .A1(n12011), .A2(n18678), .ZN(n10212) );
  OR3_X1 U11868 ( .A1(n17115), .A2(n20330), .A3(n13298), .ZN(n14372) );
  NAND2_X1 U11869 ( .A1(n14372), .A2(n13637), .ZN(n21219) );
  NAND2_X1 U11870 ( .A1(n13294), .A2(n13128), .ZN(n14532) );
  OR2_X1 U11871 ( .A1(n13127), .A2(n13126), .ZN(n13128) );
  INV_X1 U11872 ( .A(n14689), .ZN(n9873) );
  NOR2_X1 U11873 ( .A1(n9870), .A2(n9869), .ZN(n9868) );
  INV_X1 U11874 ( .A(n15147), .ZN(n9870) );
  NAND2_X1 U11875 ( .A1(n13129), .A2(n21383), .ZN(n20583) );
  NAND2_X1 U11876 ( .A1(n10025), .A2(n10024), .ZN(n10023) );
  INV_X1 U11877 ( .A(n14575), .ZN(n10025) );
  NOR2_X1 U11878 ( .A1(n15325), .A2(n15328), .ZN(n10024) );
  XNOR2_X1 U11879 ( .A(n15106), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15324) );
  NAND2_X1 U11880 ( .A1(n15105), .A2(n15104), .ZN(n15106) );
  NAND2_X1 U11881 ( .A1(n9675), .A2(n15103), .ZN(n15104) );
  XNOR2_X1 U11882 ( .A(n10084), .B(n10083), .ZN(n15341) );
  INV_X1 U11883 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10083) );
  XNOR2_X1 U11884 ( .A(n9815), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15469) );
  NAND2_X1 U11885 ( .A1(n9819), .A2(n9816), .ZN(n9815) );
  NOR2_X1 U11886 ( .A1(n15252), .A2(n9817), .ZN(n9816) );
  NAND2_X1 U11887 ( .A1(n15250), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n9819) );
  AND2_X1 U11888 ( .A1(n15431), .A2(n15430), .ZN(n15483) );
  AND2_X1 U11889 ( .A1(n14502), .A2(n14501), .ZN(n20560) );
  INV_X1 U11890 ( .A(n15267), .ZN(n20577) );
  NAND2_X1 U11891 ( .A1(n10365), .A2(n12468), .ZN(n12658) );
  INV_X1 U11892 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21022) );
  CLKBUF_X1 U11893 ( .A(n14959), .Z(n14960) );
  NAND2_X1 U11894 ( .A1(n20585), .A2(n12679), .ZN(n21017) );
  INV_X1 U11895 ( .A(n21383), .ZN(n21075) );
  OAI21_X1 U11896 ( .B1(n11859), .B2(n15911), .A(n10179), .ZN(n10178) );
  INV_X1 U11897 ( .A(n10180), .ZN(n10179) );
  OAI21_X1 U11898 ( .B1(n14611), .B2(n19405), .A(n14610), .ZN(n10180) );
  AND2_X1 U11899 ( .A1(n15623), .A2(n16210), .ZN(n15612) );
  AND2_X1 U11900 ( .A1(n13484), .A2(n13777), .ZN(n15942) );
  AND2_X1 U11901 ( .A1(n10184), .A2(n16337), .ZN(n10183) );
  NAND2_X1 U11902 ( .A1(n20309), .A2(n13488), .ZN(n15958) );
  NAND2_X1 U11903 ( .A1(n16761), .A2(n15942), .ZN(n19386) );
  INV_X1 U11904 ( .A(n19407), .ZN(n19384) );
  INV_X1 U11905 ( .A(n19403), .ZN(n19392) );
  INV_X1 U11906 ( .A(n19404), .ZN(n19389) );
  NAND2_X1 U11907 ( .A1(n13628), .A2(n16865), .ZN(n19407) );
  AND2_X1 U11908 ( .A1(n15958), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19404) );
  OR2_X1 U11909 ( .A1(n13581), .A2(n13580), .ZN(n19403) );
  INV_X1 U11910 ( .A(n15911), .ZN(n19413) );
  INV_X1 U11911 ( .A(n11859), .ZN(n11860) );
  XNOR2_X1 U11912 ( .A(n15598), .B(n9755), .ZN(n14612) );
  NAND2_X1 U11913 ( .A1(n9864), .A2(n10287), .ZN(n16079) );
  NAND2_X1 U11914 ( .A1(n15976), .A2(n10288), .ZN(n10287) );
  INV_X1 U11915 ( .A(n9865), .ZN(n9864) );
  NOR2_X1 U11916 ( .A1(n10289), .A2(n11856), .ZN(n10288) );
  INV_X1 U11917 ( .A(n16430), .ZN(n16088) );
  OR2_X1 U11918 ( .A1(n14636), .A2(n19431), .ZN(n16200) );
  INV_X1 U11919 ( .A(n10912), .ZN(n13899) );
  NOR2_X1 U11920 ( .A1(n11448), .A2(n9975), .ZN(n9974) );
  INV_X1 U11921 ( .A(n11455), .ZN(n9975) );
  NAND2_X1 U11922 ( .A1(n16295), .A2(n16571), .ZN(n16558) );
  INV_X1 U11923 ( .A(n19586), .ZN(n19574) );
  AND2_X1 U11924 ( .A1(n11451), .A2(n10884), .ZN(n19586) );
  NAND2_X1 U11925 ( .A1(n17198), .A2(n16755), .ZN(n19573) );
  INV_X1 U11926 ( .A(n19573), .ZN(n19592) );
  XNOR2_X1 U11927 ( .A(n11450), .B(n9678), .ZN(n16436) );
  INV_X1 U11928 ( .A(n11531), .ZN(n11420) );
  OAI211_X1 U11929 ( .C1(n9926), .C2(n9883), .A(n9881), .B(n9877), .ZN(n16208)
         );
  NAND2_X1 U11930 ( .A1(n9926), .A2(n9670), .ZN(n9877) );
  NAND2_X1 U11931 ( .A1(n16250), .A2(n11242), .ZN(n16238) );
  NAND2_X1 U11932 ( .A1(n10042), .A2(n17224), .ZN(n10041) );
  INV_X1 U11933 ( .A(n11870), .ZN(n10042) );
  AND2_X1 U11934 ( .A1(n10330), .A2(n10331), .ZN(n16323) );
  NAND2_X1 U11935 ( .A1(n11409), .A2(n10888), .ZN(n17203) );
  NAND2_X1 U11936 ( .A1(n11409), .A2(n11408), .ZN(n17227) );
  INV_X1 U11937 ( .A(n17203), .ZN(n17215) );
  INV_X2 U11938 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20306) );
  AND2_X1 U11939 ( .A1(n13626), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n17236) );
  NAND2_X1 U11940 ( .A1(n19214), .A2(n19185), .ZN(n18173) );
  XNOR2_X1 U11941 ( .A(n17399), .B(n10209), .ZN(n10208) );
  INV_X1 U11942 ( .A(n17400), .ZN(n10209) );
  INV_X1 U11943 ( .A(n17706), .ZN(n17725) );
  NAND2_X1 U11944 ( .A1(n9753), .A2(n9651), .ZN(n9954) );
  AND2_X1 U11945 ( .A1(n12006), .A2(n12005), .ZN(n16880) );
  OR2_X1 U11946 ( .A1(n14009), .A2(n13930), .ZN(n18123) );
  OR2_X1 U11947 ( .A1(n14009), .A2(n17863), .ZN(n18120) );
  NAND2_X1 U11948 ( .A1(n10088), .A2(n9765), .ZN(n10087) );
  INV_X1 U11949 ( .A(n16896), .ZN(n10088) );
  AND2_X1 U11950 ( .A1(n18473), .A2(n17042), .ZN(n18428) );
  NOR2_X1 U11951 ( .A1(n9980), .A2(n9981), .ZN(n16878) );
  AOI21_X1 U11952 ( .B1(n16883), .B2(n18728), .A(n10000), .ZN(n12256) );
  NAND2_X1 U11953 ( .A1(n10002), .A2(n10001), .ZN(n10000) );
  AOI21_X1 U11954 ( .B1(n17026), .B2(n12251), .A(n16882), .ZN(n10001) );
  OR2_X1 U11955 ( .A1(n12250), .A2(n13765), .ZN(n10002) );
  AND2_X1 U11956 ( .A1(n12208), .A2(n19214), .ZN(n18724) );
  AND2_X1 U11957 ( .A1(n19178), .A2(n18724), .ZN(n18728) );
  AOI21_X1 U11958 ( .B1(n9607), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n10168), .ZN(n13072) );
  AND2_X1 U11959 ( .A1(n10147), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n10168) );
  AOI21_X1 U11960 ( .B1(n9607), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n10163), .ZN(n12989) );
  AND2_X1 U11961 ( .A1(n12353), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10163) );
  AND2_X1 U11962 ( .A1(n12353), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10162) );
  INV_X1 U11963 ( .A(n13504), .ZN(n13108) );
  NAND2_X1 U11964 ( .A1(n11698), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n10125) );
  OR3_X1 U11965 ( .A1(n12151), .A2(n13752), .A3(n18762), .ZN(n12161) );
  NAND2_X1 U11966 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20988), .ZN(
        n13227) );
  OR2_X1 U11967 ( .A1(n13224), .A2(n13227), .ZN(n13226) );
  AND2_X1 U11968 ( .A1(n13226), .A2(n13217), .ZN(n13239) );
  AND2_X1 U11969 ( .A1(n10151), .A2(n10150), .ZN(n13514) );
  NAND2_X1 U11970 ( .A1(n13068), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10150) );
  NAND2_X1 U11971 ( .A1(n10147), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10151) );
  AOI21_X1 U11972 ( .B1(n13043), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A(
        n10156), .ZN(n12633) );
  AND2_X1 U11973 ( .A1(n10147), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10156) );
  AOI21_X1 U11974 ( .B1(n13503), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A(
        n10171), .ZN(n13040) );
  AND2_X1 U11975 ( .A1(n10147), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n10171) );
  AOI21_X1 U11976 ( .B1(n9607), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A(
        n10164), .ZN(n13027) );
  AND2_X1 U11977 ( .A1(n10147), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10164) );
  AOI21_X1 U11978 ( .B1(n13068), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n10173), .ZN(n12954) );
  AND2_X1 U11979 ( .A1(n10147), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n10173) );
  AOI21_X1 U11980 ( .B1(n13513), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A(
        n10161), .ZN(n12967) );
  AND2_X1 U11981 ( .A1(n10147), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10161) );
  AOI21_X1 U11982 ( .B1(n13016), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n10174), .ZN(n12933) );
  AND2_X1 U11983 ( .A1(n10147), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n10174) );
  AOI21_X1 U11984 ( .B1(n9606), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A(
        n10167), .ZN(n12872) );
  AND2_X1 U11985 ( .A1(n10147), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10167) );
  AOI21_X1 U11986 ( .B1(n13043), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A(
        n10159), .ZN(n12767) );
  AND2_X1 U11987 ( .A1(n10147), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10159) );
  AOI21_X1 U11988 ( .B1(n13043), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A(
        n10152), .ZN(n12794) );
  AND2_X1 U11989 ( .A1(n10147), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n10152) );
  AOI21_X1 U11990 ( .B1(n9607), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n10166), .ZN(n12814) );
  AND2_X1 U11991 ( .A1(n10147), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n10166) );
  AOI21_X1 U11992 ( .B1(n13043), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A(
        n10157), .ZN(n12778) );
  AND2_X1 U11993 ( .A1(n10147), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10157) );
  AOI21_X1 U11994 ( .B1(n9607), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A(
        n10169), .ZN(n12723) );
  AND2_X1 U11995 ( .A1(n10147), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n10169) );
  AOI21_X1 U11996 ( .B1(n13043), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A(
        n10158), .ZN(n12711) );
  AND2_X1 U11997 ( .A1(n10147), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10158) );
  INV_X1 U11998 ( .A(n12536), .ZN(n13146) );
  AOI21_X1 U11999 ( .B1(n10372), .B2(n10374), .A(n9710), .ZN(n10370) );
  OR2_X1 U12000 ( .A1(n12569), .A2(n12568), .ZN(n13136) );
  NAND2_X1 U12001 ( .A1(n13154), .A2(n12417), .ZN(n12419) );
  OAI22_X1 U12002 ( .A1(n10138), .A2(n9662), .B1(n12538), .B2(n10137), .ZN(
        n10136) );
  INV_X1 U12003 ( .A(n12538), .ZN(n10138) );
  NOR2_X1 U12004 ( .A1(n9662), .A2(n10368), .ZN(n10137) );
  NOR2_X1 U12005 ( .A1(n12538), .A2(n9662), .ZN(n10135) );
  AND2_X1 U12006 ( .A1(n12522), .A2(n9684), .ZN(n10044) );
  AOI21_X1 U12007 ( .B1(n12484), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n12286), .ZN(n12288) );
  OAI21_X1 U12008 ( .B1(n12544), .B2(n20603), .A(n10012), .ZN(n13234) );
  AND2_X1 U12009 ( .A1(n13222), .A2(n10013), .ZN(n10012) );
  NAND2_X1 U12010 ( .A1(n12483), .A2(n17135), .ZN(n10013) );
  INV_X1 U12011 ( .A(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12389) );
  NOR2_X1 U12012 ( .A1(n11175), .A2(n10233), .ZN(n10232) );
  NAND2_X1 U12013 ( .A1(n10408), .A2(n9697), .ZN(n10233) );
  NOR2_X1 U12014 ( .A1(n11107), .A2(n11109), .ZN(n9932) );
  CLKBUF_X1 U12015 ( .A(n11694), .Z(n11842) );
  CLKBUF_X1 U12016 ( .A(n11728), .Z(n11702) );
  CLKBUF_X1 U12017 ( .A(n11699), .Z(n11848) );
  CLKBUF_X1 U12018 ( .A(n11697), .Z(n11849) );
  AOI22_X1 U12019 ( .A1(n10821), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11700), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10436) );
  INV_X1 U12020 ( .A(n16236), .ZN(n10133) );
  NAND2_X1 U12021 ( .A1(n11262), .A2(n9937), .ZN(n11263) );
  AND2_X1 U12022 ( .A1(n9646), .A2(n11142), .ZN(n10332) );
  INV_X1 U12023 ( .A(n11073), .ZN(n9785) );
  INV_X1 U12024 ( .A(n16379), .ZN(n11065) );
  NAND2_X1 U12025 ( .A1(n10889), .A2(n10838), .ZN(n10890) );
  NOR2_X1 U12026 ( .A1(n10403), .A2(n9777), .ZN(n9776) );
  XNOR2_X1 U12027 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10799) );
  OR2_X1 U12028 ( .A1(n18175), .A2(n18178), .ZN(n13608) );
  NOR2_X1 U12029 ( .A1(n11953), .A2(n18117), .ZN(n11973) );
  INV_X1 U12030 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12170) );
  AOI21_X1 U12031 ( .B1(n12171), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n12179), .ZN(n12177) );
  NAND2_X1 U12032 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21323), .ZN(
        n12180) );
  NOR2_X1 U12033 ( .A1(n12188), .A2(n12180), .ZN(n12179) );
  AND2_X1 U12034 ( .A1(n12143), .A2(n18779), .ZN(n12151) );
  OR2_X1 U12035 ( .A1(n13257), .A2(n13256), .ZN(n13299) );
  NOR2_X1 U12036 ( .A1(n10396), .A2(n13295), .ZN(n10395) );
  NAND2_X1 U12037 ( .A1(n10401), .A2(n9732), .ZN(n10388) );
  AOI21_X1 U12038 ( .B1(n12461), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A(
        n10165), .ZN(n12750) );
  AND2_X1 U12039 ( .A1(n10147), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n10165) );
  AND2_X1 U12040 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n12602), .ZN(
        n12682) );
  NAND2_X1 U12041 ( .A1(n10004), .A2(n10005), .ZN(n13163) );
  AND2_X1 U12042 ( .A1(n13156), .A2(n10006), .ZN(n10005) );
  NAND2_X1 U12043 ( .A1(n14535), .A2(n14534), .ZN(n14536) );
  AND2_X1 U12044 ( .A1(n10252), .A2(n10251), .ZN(n10250) );
  INV_X1 U12045 ( .A(n14708), .ZN(n10251) );
  NOR2_X1 U12046 ( .A1(n14723), .A2(n10253), .ZN(n10252) );
  INV_X1 U12047 ( .A(n14734), .ZN(n10253) );
  NAND2_X1 U12048 ( .A1(n10060), .A2(n10372), .ZN(n14538) );
  AND2_X1 U12049 ( .A1(n9942), .A2(n9941), .ZN(n10060) );
  NAND2_X1 U12050 ( .A1(n15291), .A2(n15251), .ZN(n15249) );
  INV_X1 U12051 ( .A(n14503), .ZN(n10238) );
  AOI21_X1 U12052 ( .B1(n13043), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A(
        n10155), .ZN(n12592) );
  NAND2_X1 U12053 ( .A1(n13130), .A2(n13858), .ZN(n13134) );
  NOR2_X1 U12054 ( .A1(n12352), .A2(n12351), .ZN(n12365) );
  AOI21_X1 U12055 ( .B1(n9591), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A(n10160), .ZN(n12491) );
  INV_X1 U12056 ( .A(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n21252) );
  OR2_X1 U12057 ( .A1(n12467), .A2(n12466), .ZN(n13152) );
  NAND2_X1 U12058 ( .A1(n10366), .A2(n9694), .ZN(n10051) );
  INV_X1 U12059 ( .A(n12509), .ZN(n10050) );
  NAND2_X1 U12060 ( .A1(n12646), .A2(n12647), .ZN(n12678) );
  XNOR2_X1 U12061 ( .A(n12675), .B(n12674), .ZN(n20661) );
  NAND2_X1 U12062 ( .A1(n10056), .A2(n9711), .ZN(n10055) );
  NAND2_X1 U12063 ( .A1(n10054), .A2(n10053), .ZN(n10052) );
  AOI22_X1 U12064 ( .A1(n12324), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13504), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12329) );
  AOI21_X1 U12065 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n20589), .A(
        n13257), .ZN(n13252) );
  INV_X1 U12066 ( .A(n13299), .ZN(n13262) );
  NAND2_X1 U12067 ( .A1(n13251), .A2(n13250), .ZN(n13263) );
  OR2_X1 U12068 ( .A1(n15557), .A2(n15556), .ZN(n17129) );
  AND2_X1 U12069 ( .A1(n15562), .A2(n15561), .ZN(n17130) );
  OR2_X1 U12070 ( .A1(n11244), .A2(n9762), .ZN(n10228) );
  INV_X1 U12071 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n10229) );
  INV_X1 U12072 ( .A(n15767), .ZN(n10191) );
  AND2_X1 U12073 ( .A1(n21360), .A2(n11320), .ZN(n10227) );
  NAND2_X1 U12074 ( .A1(n9571), .A2(n10356), .ZN(n11116) );
  OAI21_X1 U12075 ( .B1(n9820), .B2(n11369), .A(n11367), .ZN(n9832) );
  AND2_X1 U12076 ( .A1(n10299), .A2(n11771), .ZN(n9856) );
  INV_X1 U12077 ( .A(n16589), .ZN(n10262) );
  NOR2_X1 U12078 ( .A1(n10586), .A2(n10585), .ZN(n11098) );
  OR2_X1 U12079 ( .A1(n10584), .A2(n10583), .ZN(n10585) );
  NOR2_X1 U12080 ( .A1(n13466), .A2(n11452), .ZN(n13467) );
  NOR2_X1 U12081 ( .A1(n15737), .A2(n10118), .ZN(n10117) );
  NAND2_X1 U12082 ( .A1(n13462), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13461) );
  NOR2_X1 U12083 ( .A1(n11554), .A2(n10127), .ZN(n10354) );
  NOR2_X1 U12084 ( .A1(n13455), .A2(n16328), .ZN(n13457) );
  OAI21_X1 U12085 ( .B1(n11390), .B2(n20217), .A(n11310), .ZN(n9834) );
  OAI21_X1 U12086 ( .B1(n11390), .B2(n11300), .A(n11298), .ZN(n9822) );
  NOR2_X1 U12087 ( .A1(n10363), .A2(n11484), .ZN(n10362) );
  INV_X1 U12088 ( .A(n10364), .ZN(n10363) );
  OAI21_X1 U12089 ( .B1(n9820), .B2(n11480), .A(n11396), .ZN(n9844) );
  AND2_X1 U12090 ( .A1(n10132), .A2(n11269), .ZN(n9977) );
  AND2_X1 U12091 ( .A1(n11416), .A2(n10414), .ZN(n11269) );
  OR2_X1 U12092 ( .A1(n11415), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10414) );
  NOR2_X1 U12093 ( .A1(n11512), .A2(n11274), .ZN(n10364) );
  INV_X1 U12094 ( .A(n11242), .ZN(n10130) );
  INV_X1 U12095 ( .A(n9691), .ZN(n10131) );
  INV_X1 U12096 ( .A(n15648), .ZN(n10256) );
  NAND2_X1 U12097 ( .A1(n9938), .A2(n11293), .ZN(n11270) );
  INV_X1 U12098 ( .A(n15655), .ZN(n9938) );
  NAND2_X1 U12099 ( .A1(n10264), .A2(n15721), .ZN(n10263) );
  INV_X1 U12100 ( .A(n10078), .ZN(n10077) );
  NOR2_X1 U12101 ( .A1(n16333), .A2(n10329), .ZN(n10328) );
  INV_X1 U12102 ( .A(n16320), .ZN(n10329) );
  NAND2_X1 U12103 ( .A1(n11329), .A2(n9829), .ZN(n11330) );
  INV_X1 U12104 ( .A(n9830), .ZN(n9829) );
  OAI21_X1 U12105 ( .B1(n10339), .B2(n10338), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10337) );
  NOR2_X1 U12106 ( .A1(n10338), .A2(n9902), .ZN(n10335) );
  NOR2_X1 U12107 ( .A1(n16354), .A2(n10340), .ZN(n10339) );
  INV_X1 U12108 ( .A(n16365), .ZN(n10340) );
  INV_X1 U12109 ( .A(n10994), .ZN(n11380) );
  NAND2_X1 U12110 ( .A1(n9808), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9807) );
  INV_X1 U12111 ( .A(n9811), .ZN(n9808) );
  NAND2_X1 U12112 ( .A1(n10348), .A2(n10350), .ZN(n10027) );
  INV_X1 U12113 ( .A(n10351), .ZN(n10348) );
  NAND2_X1 U12114 ( .A1(n9919), .A2(n16379), .ZN(n11073) );
  NAND2_X1 U12115 ( .A1(n11072), .A2(n16711), .ZN(n9919) );
  AND2_X1 U12116 ( .A1(n16711), .A2(n16379), .ZN(n11068) );
  NAND2_X1 U12117 ( .A1(n10979), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n9898) );
  AOI21_X1 U12118 ( .B1(n10994), .B2(P2_EBX_REG_0__SCAN_IN), .A(n10965), .ZN(
        n10967) );
  AND3_X1 U12119 ( .A1(n10541), .A2(n10540), .A3(n10539), .ZN(n14357) );
  NAND2_X1 U12120 ( .A1(n11561), .A2(n20306), .ZN(n11583) );
  NOR2_X2 U12121 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16786) );
  OR2_X1 U12122 ( .A1(n11775), .A2(n11585), .ZN(n11586) );
  INV_X1 U12123 ( .A(n10946), .ZN(n10911) );
  AND2_X1 U12124 ( .A1(n11572), .A2(n11577), .ZN(n11013) );
  INV_X1 U12125 ( .A(n10773), .ZN(n10284) );
  INV_X1 U12126 ( .A(n10777), .ZN(n10280) );
  NAND2_X1 U12127 ( .A1(n10820), .A2(n10441), .ZN(n9851) );
  INV_X1 U12128 ( .A(n20288), .ZN(n19598) );
  NAND3_X1 U12129 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n20305), .A3(n20133), 
        .ZN(n16809) );
  XNOR2_X1 U12130 ( .A(n10980), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10793) );
  NAND2_X1 U12131 ( .A1(n10779), .A2(n10778), .ZN(n10794) );
  OR3_X1 U12132 ( .A1(n10804), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(
        n17156), .ZN(n11094) );
  INV_X1 U12133 ( .A(n17464), .ZN(n10197) );
  AND2_X1 U12134 ( .A1(n11884), .A2(n13785), .ZN(n11980) );
  AND2_X1 U12135 ( .A1(n13758), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11885) );
  NOR2_X2 U12136 ( .A1(n13596), .A2(n18277), .ZN(n13599) );
  OR2_X1 U12137 ( .A1(n10217), .A2(n18316), .ZN(n10216) );
  NAND2_X1 U12138 ( .A1(n10218), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10217) );
  INV_X1 U12139 ( .A(n16966), .ZN(n10218) );
  NAND2_X1 U12140 ( .A1(n17040), .A2(n9916), .ZN(n9915) );
  AND2_X1 U12141 ( .A1(n10095), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9916) );
  AOI21_X1 U12142 ( .B1(n12026), .B2(n18357), .A(n12025), .ZN(n12027) );
  NAND2_X1 U12143 ( .A1(n18258), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9923) );
  AOI21_X1 U12144 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n19188), .A(
        n12184), .ZN(n12190) );
  AND2_X1 U12145 ( .A1(n18766), .A2(n18783), .ZN(n12200) );
  INV_X1 U12146 ( .A(n13930), .ZN(n13728) );
  INV_X1 U12147 ( .A(n20420), .ZN(n20376) );
  INV_X1 U12148 ( .A(n10247), .ZN(n10245) );
  AOI21_X1 U12149 ( .B1(n15107), .B2(n13531), .A(n13530), .ZN(n14663) );
  INV_X1 U12150 ( .A(n20584), .ZN(n20582) );
  NAND2_X1 U12151 ( .A1(n14663), .A2(n10395), .ZN(n10394) );
  AND2_X1 U12152 ( .A1(n13100), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13101) );
  OAI21_X1 U12153 ( .B1(n15125), .B2(n13524), .A(n13098), .ZN(n14677) );
  AND2_X1 U12154 ( .A1(n13055), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13056) );
  AND2_X1 U12155 ( .A1(n13081), .A2(n13080), .ZN(n14690) );
  OR2_X1 U12156 ( .A1(n15134), .A2(n13524), .ZN(n13081) );
  INV_X1 U12157 ( .A(n13009), .ZN(n13010) );
  AND2_X1 U12158 ( .A1(n13036), .A2(n13035), .ZN(n14721) );
  OR2_X1 U12159 ( .A1(n15153), .A2(n13524), .ZN(n13036) );
  NOR2_X2 U12160 ( .A1(n12965), .A2(n15179), .ZN(n12943) );
  INV_X1 U12161 ( .A(n10401), .ZN(n10387) );
  AND2_X1 U12162 ( .A1(n12922), .A2(n12921), .ZN(n14786) );
  CLKBUF_X1 U12163 ( .A(n14770), .Z(n14771) );
  AND2_X1 U12164 ( .A1(n12898), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12899) );
  OR2_X1 U12165 ( .A1(n15206), .A2(n13524), .ZN(n12903) );
  INV_X1 U12166 ( .A(n14812), .ZN(n10391) );
  AND2_X1 U12167 ( .A1(n12855), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12856) );
  AND2_X1 U12168 ( .A1(n12861), .A2(n12860), .ZN(n14827) );
  NAND2_X1 U12169 ( .A1(n12805), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12854) );
  NOR2_X1 U12170 ( .A1(n12836), .A2(n14926), .ZN(n9875) );
  OR2_X1 U12171 ( .A1(n12835), .A2(n12834), .ZN(n12836) );
  AND3_X1 U12172 ( .A1(n14850), .A2(n14877), .A3(n14893), .ZN(n14878) );
  AND2_X1 U12173 ( .A1(n12742), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12743) );
  INV_X1 U12174 ( .A(n12741), .ZN(n12742) );
  NAND2_X1 U12175 ( .A1(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n12734), .ZN(
        n12741) );
  AND2_X1 U12176 ( .A1(n12715), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12734) );
  INV_X1 U12177 ( .A(n12642), .ZN(n12715) );
  NAND2_X1 U12178 ( .A1(n12623), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12642) );
  NAND2_X1 U12179 ( .A1(n12603), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12622) );
  INV_X1 U12180 ( .A(n12698), .ZN(n12603) );
  NAND2_X1 U12181 ( .A1(n12682), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12698) );
  NAND2_X1 U12182 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12683) );
  NAND2_X1 U12183 ( .A1(n10086), .A2(n13404), .ZN(n10085) );
  INV_X1 U12184 ( .A(n13214), .ZN(n10086) );
  NAND2_X1 U12185 ( .A1(n14746), .A2(n10250), .ZN(n14710) );
  NAND2_X1 U12186 ( .A1(n14746), .A2(n10252), .ZN(n14725) );
  NAND2_X1 U12187 ( .A1(n14746), .A2(n14734), .ZN(n14736) );
  NOR2_X1 U12188 ( .A1(n15396), .A2(n14573), .ZN(n15377) );
  AND2_X1 U12189 ( .A1(n13389), .A2(n13388), .ZN(n14748) );
  AND2_X1 U12190 ( .A1(n13387), .A2(n13386), .ZN(n14762) );
  NOR2_X2 U12191 ( .A1(n14774), .A2(n14762), .ZN(n14761) );
  XNOR2_X1 U12192 ( .A(n9569), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15202) );
  AND2_X1 U12193 ( .A1(n9569), .A2(n15218), .ZN(n15233) );
  AOI21_X1 U12194 ( .B1(n14569), .B2(n10017), .A(n10016), .ZN(n10015) );
  INV_X1 U12195 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n10016) );
  INV_X1 U12196 ( .A(n15426), .ZN(n10017) );
  OR2_X1 U12197 ( .A1(n20549), .A2(n10018), .ZN(n10014) );
  INV_X1 U12198 ( .A(n14569), .ZN(n10018) );
  AND2_X1 U12199 ( .A1(n13368), .A2(n13367), .ZN(n14853) );
  NAND2_X1 U12200 ( .A1(n9818), .A2(n15264), .ZN(n9817) );
  NAND2_X1 U12201 ( .A1(n9569), .A2(n15482), .ZN(n9818) );
  AND2_X1 U12202 ( .A1(n13361), .A2(n13360), .ZN(n14881) );
  NOR2_X1 U12203 ( .A1(n14897), .A2(n14881), .ZN(n14880) );
  NAND2_X1 U12204 ( .A1(n10247), .A2(n13339), .ZN(n10246) );
  NAND2_X1 U12205 ( .A1(n9791), .A2(n10057), .ZN(n9790) );
  XNOR2_X1 U12206 ( .A(n13168), .B(n14495), .ZN(n17162) );
  NAND2_X1 U12207 ( .A1(n17163), .A2(n17162), .ZN(n17165) );
  AND2_X1 U12208 ( .A1(n15586), .A2(n10368), .ZN(n13275) );
  OR2_X1 U12209 ( .A1(n14296), .A2(n14297), .ZN(n20417) );
  NAND2_X1 U12210 ( .A1(n14658), .A2(n13860), .ZN(n14487) );
  AOI21_X1 U12211 ( .B1(n14479), .B2(n14478), .A(n20330), .ZN(n14502) );
  NAND2_X1 U12212 ( .A1(n10020), .A2(n10019), .ZN(n14479) );
  INV_X1 U12213 ( .A(n20661), .ZN(n21384) );
  NAND2_X1 U12214 ( .A1(n10366), .A2(n10368), .ZN(n10365) );
  NAND2_X1 U12215 ( .A1(n13962), .A2(n10368), .ZN(n9789) );
  NAND2_X1 U12216 ( .A1(n12559), .A2(n12679), .ZN(n12690) );
  NOR2_X1 U12217 ( .A1(n20662), .A2(n20661), .ZN(n20872) );
  NOR2_X2 U12218 ( .A1(n20584), .A2(n20583), .ZN(n20628) );
  OR2_X1 U12219 ( .A1(n21017), .A2(n20926), .ZN(n20591) );
  NAND3_X1 U12220 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n10368), .A3(n20588), 
        .ZN(n20627) );
  INV_X1 U12221 ( .A(n17185), .ZN(n17141) );
  XNOR2_X1 U12222 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n13413) );
  INV_X1 U12223 ( .A(n17236), .ZN(n13629) );
  NAND2_X1 U12224 ( .A1(n10869), .A2(n10868), .ZN(n11083) );
  NAND2_X1 U12225 ( .A1(n11038), .A2(n10356), .ZN(n10869) );
  INV_X1 U12226 ( .A(n10879), .ZN(n16854) );
  INV_X1 U12227 ( .A(n20297), .ZN(n11440) );
  AND2_X1 U12228 ( .A1(n19404), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10123) );
  NAND2_X1 U12229 ( .A1(n15652), .A2(n16228), .ZN(n15637) );
  OAI21_X1 U12230 ( .B1(n15668), .B2(n16239), .A(n16761), .ZN(n15652) );
  NAND2_X1 U12231 ( .A1(n13459), .A2(n9672), .ZN(n15765) );
  NOR2_X1 U12232 ( .A1(n11175), .A2(n10231), .ZN(n10230) );
  INV_X1 U12233 ( .A(n10408), .ZN(n10231) );
  NAND2_X1 U12234 ( .A1(n11158), .A2(n10226), .ZN(n11199) );
  AND2_X1 U12235 ( .A1(n10227), .A2(n16064), .ZN(n10226) );
  INV_X1 U12236 ( .A(n15814), .ZN(n15813) );
  NAND2_X1 U12237 ( .A1(n15846), .A2(n16359), .ZN(n15836) );
  NAND2_X1 U12238 ( .A1(n11158), .A2(n21360), .ZN(n11160) );
  NAND2_X1 U12239 ( .A1(n15875), .A2(n16387), .ZN(n15861) );
  INV_X1 U12240 ( .A(n15875), .ZN(n15872) );
  NOR2_X1 U12241 ( .A1(n15887), .A2(n16401), .ZN(n15875) );
  NAND2_X1 U12242 ( .A1(n9680), .A2(n9934), .ZN(n11104) );
  INV_X1 U12243 ( .A(n11107), .ZN(n9934) );
  NAND2_X1 U12244 ( .A1(n10995), .A2(n9827), .ZN(n10997) );
  INV_X1 U12245 ( .A(n9828), .ZN(n9827) );
  INV_X1 U12246 ( .A(n14229), .ZN(n16848) );
  INV_X1 U12247 ( .A(n15975), .ZN(n10289) );
  OAI21_X1 U12248 ( .B1(n15976), .B2(n10290), .A(n10286), .ZN(n9865) );
  INV_X1 U12249 ( .A(n10291), .ZN(n10290) );
  AOI21_X1 U12250 ( .B1(n10291), .B2(n10289), .A(n9648), .ZN(n10286) );
  NOR2_X1 U12251 ( .A1(n10292), .A2(n11834), .ZN(n10291) );
  AND2_X1 U12252 ( .A1(n10762), .A2(n10761), .ZN(n11426) );
  XNOR2_X1 U12253 ( .A(n11778), .B(n11796), .ZN(n15987) );
  NOR2_X1 U12254 ( .A1(n9854), .A2(n9853), .ZN(n11772) );
  NAND2_X1 U12255 ( .A1(n9857), .A2(n9855), .ZN(n16001) );
  AND2_X1 U12256 ( .A1(n10752), .A2(n10751), .ZN(n15664) );
  AND2_X1 U12257 ( .A1(n9750), .A2(n11612), .ZN(n9860) );
  OR2_X1 U12258 ( .A1(n11632), .A2(n11631), .ZN(n16034) );
  AND2_X1 U12259 ( .A1(n10734), .A2(n10733), .ZN(n15775) );
  CLKBUF_X1 U12260 ( .A(n15778), .Z(n15779) );
  AND3_X1 U12261 ( .A1(n10717), .A2(n10716), .A3(n10715), .ZN(n15795) );
  AND3_X1 U12262 ( .A1(n10661), .A2(n10660), .A3(n10659), .ZN(n14201) );
  AND3_X1 U12263 ( .A1(n10644), .A2(n10643), .A3(n10642), .ZN(n15856) );
  CLKBUF_X1 U12264 ( .A(n14200), .Z(n15859) );
  AND3_X1 U12265 ( .A1(n10558), .A2(n10557), .A3(n10556), .ZN(n14362) );
  CLKBUF_X1 U12266 ( .A(n14360), .Z(n14361) );
  AND2_X1 U12267 ( .A1(n10946), .A2(n10945), .ZN(n13900) );
  AND2_X1 U12268 ( .A1(n19445), .A2(n10399), .ZN(n14635) );
  AND2_X1 U12269 ( .A1(n19445), .A2(n13905), .ZN(n16197) );
  AND2_X1 U12270 ( .A1(n13633), .A2(n13498), .ZN(n19538) );
  INV_X1 U12271 ( .A(n19430), .ZN(n19431) );
  NAND2_X1 U12272 ( .A1(n11385), .A2(n9839), .ZN(n11387) );
  INV_X1 U12273 ( .A(n9840), .ZN(n9839) );
  AND2_X1 U12274 ( .A1(n13462), .A2(n10116), .ZN(n13464) );
  AND2_X1 U12275 ( .A1(n9647), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10116) );
  NAND2_X1 U12276 ( .A1(n13462), .A2(n9647), .ZN(n13463) );
  AND2_X1 U12277 ( .A1(n10354), .A2(n11555), .ZN(n10353) );
  NOR3_X1 U12278 ( .A1(n13455), .A2(n10109), .A3(n10110), .ZN(n13460) );
  NAND2_X1 U12279 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10108) );
  AND2_X1 U12280 ( .A1(n13454), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13452) );
  NAND2_X1 U12281 ( .A1(n9713), .A2(n10114), .ZN(n13450) );
  NOR2_X1 U12282 ( .A1(n16368), .A2(n13450), .ZN(n13454) );
  INV_X1 U12283 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16368) );
  AND2_X1 U12284 ( .A1(n10114), .A2(n10113), .ZN(n13451) );
  NAND2_X1 U12285 ( .A1(n10114), .A2(n10115), .ZN(n13445) );
  NOR2_X1 U12286 ( .A1(n13447), .A2(n17199), .ZN(n13449) );
  CLKBUF_X1 U12287 ( .A(n14244), .Z(n14245) );
  INV_X1 U12288 ( .A(n16731), .ZN(n11302) );
  INV_X1 U12289 ( .A(n16732), .ZN(n11303) );
  INV_X1 U12290 ( .A(n10362), .ZN(n10361) );
  OR2_X1 U12291 ( .A1(n11275), .A2(n11274), .ZN(n11417) );
  AND2_X1 U12292 ( .A1(n16465), .A2(n16451), .ZN(n16439) );
  INV_X1 U12293 ( .A(n11415), .ZN(n9883) );
  INV_X1 U12294 ( .A(n9925), .ZN(n9882) );
  NAND2_X1 U12295 ( .A1(n11376), .A2(n9841), .ZN(n11378) );
  INV_X1 U12296 ( .A(n9842), .ZN(n9841) );
  NOR2_X1 U12297 ( .A1(n15675), .A2(n10323), .ZN(n10322) );
  INV_X1 U12298 ( .A(n10324), .ZN(n10323) );
  INV_X1 U12299 ( .A(n15683), .ZN(n10257) );
  CLKBUF_X1 U12300 ( .A(n15690), .Z(n15691) );
  NAND2_X1 U12301 ( .A1(n11476), .A2(n10933), .ZN(n16258) );
  AND2_X1 U12302 ( .A1(n10739), .A2(n9752), .ZN(n10264) );
  INV_X1 U12303 ( .A(n15760), .ZN(n10265) );
  NAND2_X1 U12304 ( .A1(n11357), .A2(n9837), .ZN(n11358) );
  INV_X1 U12305 ( .A(n9838), .ZN(n9837) );
  CLKBUF_X1 U12306 ( .A(n11468), .Z(n11469) );
  AND2_X1 U12307 ( .A1(n10738), .A2(n10737), .ZN(n15761) );
  NOR2_X1 U12308 ( .A1(n10312), .A2(n10311), .ZN(n10310) );
  INV_X1 U12309 ( .A(n15749), .ZN(n10311) );
  NAND2_X1 U12310 ( .A1(n11343), .A2(n9835), .ZN(n11344) );
  INV_X1 U12311 ( .A(n9836), .ZN(n9835) );
  NAND2_X1 U12312 ( .A1(n11339), .A2(n9825), .ZN(n11341) );
  INV_X1 U12313 ( .A(n9826), .ZN(n9825) );
  AND3_X1 U12314 ( .A1(n10675), .A2(n10674), .A3(n10673), .ZN(n15829) );
  CLKBUF_X1 U12315 ( .A(n14282), .Z(n15827) );
  NAND2_X1 U12316 ( .A1(n11325), .A2(n9823), .ZN(n11326) );
  INV_X1 U12317 ( .A(n9824), .ZN(n9823) );
  NAND2_X1 U12318 ( .A1(n16367), .A2(n16365), .ZN(n16353) );
  NAND2_X1 U12319 ( .A1(n10308), .A2(n14331), .ZN(n10305) );
  INV_X1 U12320 ( .A(n14266), .ZN(n10306) );
  NAND2_X1 U12321 ( .A1(n16392), .A2(n11074), .ZN(n10351) );
  OR2_X1 U12322 ( .A1(n16392), .A2(n11074), .ZN(n10350) );
  XNOR2_X1 U12323 ( .A(n11075), .B(n16378), .ZN(n16392) );
  NAND2_X1 U12324 ( .A1(n16406), .A2(n11073), .ZN(n16394) );
  NAND2_X1 U12325 ( .A1(n16405), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16406) );
  AND2_X1 U12326 ( .A1(n11037), .A2(n11092), .ZN(n10104) );
  NAND2_X1 U12327 ( .A1(n10035), .A2(n11037), .ZN(n11050) );
  AND2_X1 U12328 ( .A1(n10918), .A2(n10917), .ZN(n16847) );
  OAI22_X1 U12329 ( .A1(n10979), .A2(n10973), .B1(n10994), .B2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10976) );
  NAND2_X1 U12330 ( .A1(n11003), .A2(n11002), .ZN(n11005) );
  XNOR2_X1 U12331 ( .A(n12259), .B(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13439) );
  AND2_X1 U12332 ( .A1(n13713), .A2(n10872), .ZN(n10809) );
  INV_X1 U12333 ( .A(n9780), .ZN(n10856) );
  CLKBUF_X1 U12334 ( .A(n10832), .Z(n16785) );
  INV_X1 U12335 ( .A(n11023), .ZN(n11021) );
  INV_X1 U12336 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19911) );
  INV_X1 U12337 ( .A(n19914), .ZN(n19870) );
  NOR2_X1 U12338 ( .A1(n19948), .A2(n20271), .ZN(n19952) );
  NAND2_X1 U12339 ( .A1(n20288), .A2(n19597), .ZN(n20271) );
  INV_X1 U12340 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19682) );
  NAND2_X1 U12341 ( .A1(n9849), .A2(n10441), .ZN(n9848) );
  NAND2_X1 U12342 ( .A1(n9847), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9846) );
  INV_X1 U12343 ( .A(n10901), .ZN(n19624) );
  INV_X1 U12344 ( .A(n19948), .ZN(n20070) );
  INV_X1 U12345 ( .A(n20131), .ZN(n20069) );
  NAND2_X1 U12346 ( .A1(n10464), .A2(n9910), .ZN(n9907) );
  NAND2_X1 U12347 ( .A1(n10463), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9906) );
  AND2_X1 U12348 ( .A1(n20133), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19644) );
  NOR2_X2 U12349 ( .A1(n19430), .A2(n16809), .ZN(n19639) );
  XNOR2_X1 U12350 ( .A(n10794), .B(n10780), .ZN(n10829) );
  INV_X1 U12351 ( .A(n10793), .ZN(n10780) );
  NOR2_X1 U12352 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n20307) );
  NAND2_X1 U12353 ( .A1(n10211), .A2(n10210), .ZN(n17407) );
  INV_X1 U12354 ( .A(n17410), .ZN(n10210) );
  OAI21_X1 U12355 ( .B1(n17473), .B2(n10195), .A(n10194), .ZN(n17463) );
  NAND2_X1 U12356 ( .A1(n10197), .A2(n10196), .ZN(n10195) );
  NAND2_X1 U12357 ( .A1(n17695), .A2(n10197), .ZN(n10194) );
  INV_X1 U12358 ( .A(n17474), .ZN(n10196) );
  NOR2_X1 U12359 ( .A1(n17473), .A2(n17474), .ZN(n17472) );
  NOR2_X1 U12360 ( .A1(n17695), .A2(n13602), .ZN(n17494) );
  NAND2_X1 U12361 ( .A1(n10205), .A2(n10204), .ZN(n10206) );
  INV_X1 U12362 ( .A(n17494), .ZN(n10205) );
  NOR4_X1 U12363 ( .A1(n19269), .A2(n17630), .A3(n19267), .A4(n19265), .ZN(
        n17591) );
  INV_X1 U12364 ( .A(n17673), .ZN(n17645) );
  OR2_X1 U12365 ( .A1(n19351), .A2(n13609), .ZN(n17644) );
  NAND2_X1 U12366 ( .A1(n19351), .A2(n18755), .ZN(n13614) );
  INV_X1 U12367 ( .A(n14042), .ZN(n14043) );
  NAND2_X1 U12368 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(P3_EAX_REG_28__SCAN_IN), 
        .ZN(n9960) );
  INV_X1 U12369 ( .A(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13686) );
  OR2_X1 U12370 ( .A1(n11966), .A2(n11965), .ZN(n12218) );
  AND3_X1 U12371 ( .A1(n11897), .A2(n11902), .A3(n11899), .ZN(n10091) );
  AND2_X1 U12372 ( .A1(n11885), .A2(n13785), .ZN(n13741) );
  NAND2_X1 U12373 ( .A1(n17948), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10219) );
  INV_X1 U12374 ( .A(n17251), .ZN(n16910) );
  CLKBUF_X1 U12375 ( .A(n13599), .Z(n16949) );
  INV_X1 U12376 ( .A(n18272), .ZN(n18329) );
  INV_X1 U12377 ( .A(n16965), .ZN(n13595) );
  INV_X1 U12378 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n18440) );
  NAND2_X1 U12379 ( .A1(n9922), .A2(n9923), .ZN(n17077) );
  AND2_X1 U12380 ( .A1(n12027), .A2(n12028), .ZN(n9922) );
  INV_X1 U12381 ( .A(n12026), .ZN(n18257) );
  AND2_X1 U12382 ( .A1(n18284), .A2(n18286), .ZN(n18269) );
  OR2_X1 U12383 ( .A1(n18437), .A2(n9652), .ZN(n18358) );
  INV_X1 U12384 ( .A(n18590), .ZN(n10092) );
  INV_X1 U12385 ( .A(n18652), .ZN(n10093) );
  NOR2_X1 U12386 ( .A1(n18437), .A2(n12013), .ZN(n18392) );
  INV_X1 U12387 ( .A(n13751), .ZN(n9768) );
  NAND2_X1 U12388 ( .A1(n12243), .A2(n12244), .ZN(n14151) );
  NAND2_X1 U12389 ( .A1(n9994), .A2(n9993), .ZN(n18462) );
  NAND2_X1 U12390 ( .A1(n9997), .A2(n9995), .ZN(n9993) );
  INV_X1 U12391 ( .A(n18463), .ZN(n9996) );
  INV_X1 U12392 ( .A(n9997), .ZN(n14121) );
  NAND2_X1 U12393 ( .A1(n9912), .A2(n21349), .ZN(n9911) );
  AND2_X1 U12394 ( .A1(n11934), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9913) );
  INV_X1 U12395 ( .A(n11934), .ZN(n9912) );
  AOI21_X1 U12396 ( .B1(n18485), .B2(n9998), .A(n12229), .ZN(n18476) );
  INV_X1 U12397 ( .A(n18484), .ZN(n9998) );
  XNOR2_X1 U12398 ( .A(n11918), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n18487) );
  NOR2_X1 U12399 ( .A1(n12229), .A2(n9999), .ZN(n18485) );
  AND2_X1 U12400 ( .A1(n12225), .A2(n18727), .ZN(n9999) );
  NAND2_X1 U12401 ( .A1(n13754), .A2(n13607), .ZN(n17100) );
  INV_X1 U12402 ( .A(n9956), .ZN(n13929) );
  NOR2_X1 U12403 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18754), .ZN(n19087) );
  INV_X1 U12404 ( .A(n12194), .ZN(n18762) );
  AND2_X1 U12405 ( .A1(n12099), .A2(n12098), .ZN(n18770) );
  AND4_X1 U12406 ( .A1(n12097), .A2(n12096), .A3(n12095), .A4(n12094), .ZN(
        n12098) );
  OAI21_X1 U12407 ( .B1(n12117), .B2(n12063), .A(n9968), .ZN(n12065) );
  INV_X2 U12408 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n21070) );
  CLKBUF_X1 U12409 ( .A(n13962), .Z(n20839) );
  OR2_X1 U12410 ( .A1(n20577), .A2(n13308), .ZN(n13309) );
  INV_X1 U12411 ( .A(n20427), .ZN(n20407) );
  AND2_X1 U12412 ( .A1(n13424), .A2(n13412), .ZN(n20404) );
  INV_X1 U12413 ( .A(n15013), .ZN(n20439) );
  AND2_X2 U12414 ( .A1(n13916), .A2(n14077), .ZN(n20447) );
  NAND2_X1 U12415 ( .A1(n15098), .A2(n14015), .ZN(n15070) );
  NOR2_X2 U12416 ( .A1(n14016), .A2(n20584), .ZN(n15082) );
  OAI21_X1 U12417 ( .B1(n17115), .B2(n13542), .A(n13541), .ZN(n13543) );
  AND2_X1 U12418 ( .A1(n14646), .A2(n13537), .ZN(n13542) );
  INV_X2 U12419 ( .A(n15076), .ZN(n15098) );
  AND2_X1 U12420 ( .A1(n15070), .A2(n14016), .ZN(n15100) );
  NAND2_X1 U12421 ( .A1(n20475), .A2(n20449), .ZN(n17155) );
  AND2_X1 U12422 ( .A1(n14079), .A2(n14466), .ZN(n20453) );
  INV_X2 U12423 ( .A(n17155), .ZN(n20472) );
  AND2_X1 U12424 ( .A1(n21216), .A2(n21142), .ZN(n14371) );
  INV_X1 U12425 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15179) );
  INV_X1 U12426 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15187) );
  INV_X1 U12427 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15195) );
  CLKBUF_X1 U12428 ( .A(n14923), .Z(n14924) );
  OR2_X1 U12429 ( .A1(n15010), .A2(n15009), .ZN(n20382) );
  NAND2_X1 U12430 ( .A1(n12655), .A2(n12677), .ZN(n14303) );
  INV_X1 U12431 ( .A(n17161), .ZN(n20511) );
  INV_X1 U12432 ( .A(n20338), .ZN(n20519) );
  XNOR2_X1 U12433 ( .A(n14554), .B(n14553), .ZN(n14587) );
  INV_X1 U12434 ( .A(n14549), .ZN(n14554) );
  XNOR2_X1 U12435 ( .A(n10003), .B(n9682), .ZN(n15333) );
  NAND2_X1 U12436 ( .A1(n10141), .A2(n10140), .ZN(n10003) );
  NAND2_X1 U12437 ( .A1(n9953), .A2(n9951), .ZN(n15122) );
  NAND2_X1 U12438 ( .A1(n15121), .A2(n9569), .ZN(n9953) );
  NAND2_X1 U12439 ( .A1(n15120), .A2(n9699), .ZN(n9951) );
  NAND2_X1 U12440 ( .A1(n15377), .A2(n14574), .ZN(n15362) );
  OAI21_X1 U12441 ( .B1(n15185), .B2(n10376), .A(n10374), .ZN(n15166) );
  NAND2_X1 U12442 ( .A1(n10371), .A2(n9569), .ZN(n15165) );
  OR2_X1 U12443 ( .A1(n15421), .A2(n14571), .ZN(n15396) );
  NAND2_X1 U12444 ( .A1(n13210), .A2(n13209), .ZN(n15173) );
  NAND2_X1 U12445 ( .A1(n10375), .A2(n13381), .ZN(n15174) );
  NAND2_X1 U12446 ( .A1(n10014), .A2(n10015), .ZN(n15462) );
  NAND2_X1 U12447 ( .A1(n10384), .A2(n13192), .ZN(n15307) );
  NOR2_X1 U12448 ( .A1(n20545), .A2(n20561), .ZN(n20549) );
  OR2_X1 U12449 ( .A1(n20586), .A2(n20585), .ZN(n20934) );
  INV_X1 U12450 ( .A(n15591), .ZN(n15566) );
  NOR2_X1 U12451 ( .A1(n17115), .A2(n20963), .ZN(n15591) );
  OAI22_X1 U12452 ( .A1(n20600), .A2(n20599), .B1(n20902), .B2(n20726), .ZN(
        n20631) );
  OAI211_X1 U12453 ( .C1(n10413), .C2(n20963), .A(n20898), .B(n20594), .ZN(
        n20632) );
  OAI22_X1 U12454 ( .A1(n20671), .A2(n20670), .B1(n20783), .B2(n20902), .ZN(
        n20688) );
  OAI21_X1 U12455 ( .B1(n20687), .B2(n20963), .A(n20667), .ZN(n20689) );
  OAI22_X1 U12456 ( .A1(n20702), .A2(n20701), .B1(n21070), .B2(n20700), .ZN(
        n20719) );
  INV_X1 U12457 ( .A(n20751), .ZN(n20742) );
  OAI21_X1 U12458 ( .B1(n10419), .B2(n20731), .A(n21027), .ZN(n20748) );
  INV_X1 U12459 ( .A(n20777), .ZN(n20767) );
  OAI21_X1 U12460 ( .B1(n20756), .B2(n20755), .A(n21080), .ZN(n20774) );
  OAI211_X1 U12461 ( .C1(n20802), .C2(n20963), .A(n21027), .B(n20781), .ZN(
        n20804) );
  OAI22_X1 U12462 ( .A1(n20785), .A2(n20784), .B1(n21019), .B2(n20783), .ZN(
        n20803) );
  INV_X1 U12463 ( .A(n20798), .ZN(n20801) );
  OR2_X1 U12464 ( .A1(n20807), .A2(n21016), .ZN(n20837) );
  OAI221_X1 U12465 ( .B1(n21383), .B2(n20815), .C1(n21075), .C2(n20814), .A(
        n21080), .ZN(n20834) );
  OAI211_X1 U12466 ( .C1(n10412), .C2(n20963), .A(n20898), .B(n20846), .ZN(
        n20863) );
  INV_X1 U12467 ( .A(n20900), .ZN(n20923) );
  INV_X1 U12468 ( .A(n20919), .ZN(n20921) );
  INV_X1 U12469 ( .A(n20957), .ZN(n20946) );
  OAI211_X1 U12470 ( .C1(n10418), .C2(n20963), .A(n21027), .B(n20962), .ZN(
        n20984) );
  OAI22_X1 U12471 ( .A1(n20967), .A2(n20966), .B1(n21019), .B2(n20965), .ZN(
        n20983) );
  INV_X1 U12472 ( .A(n21015), .ZN(n20982) );
  OAI221_X1 U12473 ( .B1(n21383), .B2(n20994), .C1(n21075), .C2(n20993), .A(
        n21080), .ZN(n21012) );
  OAI211_X1 U12474 ( .C1(n21057), .C2(n21028), .A(n21027), .B(n21026), .ZN(
        n21061) );
  NOR2_X2 U12475 ( .A1(n21017), .A2(n20995), .ZN(n21060) );
  OAI211_X1 U12476 ( .C1(n21383), .C2(n21081), .A(n21080), .B(n21079), .ZN(
        n21128) );
  INV_X1 U12477 ( .A(n20591), .ZN(n21127) );
  INV_X1 U12478 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20963) );
  AND2_X1 U12479 ( .A1(n16854), .A2(n13436), .ZN(n20299) );
  NOR2_X1 U12480 ( .A1(n10188), .A2(n19416), .ZN(n15601) );
  NOR2_X1 U12481 ( .A1(n10190), .A2(n10189), .ZN(n10188) );
  INV_X1 U12482 ( .A(n15623), .ZN(n10190) );
  INV_X1 U12483 ( .A(n15668), .ZN(n15665) );
  AND2_X1 U12484 ( .A1(n11214), .A2(n11213), .ZN(n15710) );
  NAND2_X1 U12485 ( .A1(n11173), .A2(n9637), .ZN(n11212) );
  NAND2_X1 U12486 ( .A1(n11179), .A2(n9630), .ZN(n15745) );
  AND2_X1 U12487 ( .A1(n13459), .A2(n16304), .ZN(n19387) );
  NOR2_X1 U12488 ( .A1(n15928), .A2(n15927), .ZN(n19415) );
  INV_X1 U12489 ( .A(n11594), .ZN(n16055) );
  OR2_X1 U12490 ( .A1(n10625), .A2(n10624), .ZN(n14326) );
  NAND2_X1 U12491 ( .A1(n16768), .A2(n13773), .ZN(n16820) );
  OAI21_X1 U12492 ( .B1(n11425), .B2(n10273), .A(n10769), .ZN(n10270) );
  NAND2_X1 U12493 ( .A1(n10269), .A2(n10271), .ZN(n10268) );
  INV_X1 U12494 ( .A(n10274), .ZN(n10273) );
  AND2_X1 U12495 ( .A1(n10301), .A2(n10304), .ZN(n16007) );
  NAND2_X1 U12496 ( .A1(n10300), .A2(n10299), .ZN(n16005) );
  AND2_X1 U12497 ( .A1(n14635), .A2(n19431), .ZN(n16193) );
  NAND2_X1 U12498 ( .A1(n13892), .A2(n13894), .ZN(n13942) );
  INV_X1 U12499 ( .A(n19451), .ZN(n19441) );
  OR2_X1 U12500 ( .A1(n19479), .A2(n19477), .ZN(n19451) );
  NAND2_X1 U12501 ( .A1(n10294), .A2(n11590), .ZN(n14344) );
  OR2_X1 U12502 ( .A1(n16197), .A2(n14635), .ZN(n19434) );
  INV_X1 U12503 ( .A(n19434), .ZN(n19485) );
  INV_X1 U12504 ( .A(n13794), .ZN(n19489) );
  NAND2_X1 U12505 ( .A1(n19523), .A2(n20310), .ZN(n19492) );
  INV_X1 U12506 ( .A(n19492), .ZN(n19521) );
  XNOR2_X1 U12507 ( .A(n10223), .B(n11295), .ZN(n12264) );
  NAND2_X1 U12508 ( .A1(n10220), .A2(n9696), .ZN(n10223) );
  NAND2_X1 U12509 ( .A1(n11537), .A2(n11536), .ZN(n11541) );
  NAND2_X1 U12510 ( .A1(n10073), .A2(n10078), .ZN(n16291) );
  NAND2_X1 U12511 ( .A1(n16314), .A2(n10079), .ZN(n10073) );
  INV_X1 U12512 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17199) );
  INV_X1 U12513 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16420) );
  NAND2_X1 U12514 ( .A1(n13624), .A2(n11444), .ZN(n17198) );
  INV_X1 U12515 ( .A(n17192), .ZN(n19582) );
  AND2_X1 U12516 ( .A1(n17198), .A2(n19583), .ZN(n17192) );
  INV_X1 U12517 ( .A(n11577), .ZN(n19593) );
  INV_X1 U12518 ( .A(n17198), .ZN(n19584) );
  NAND2_X1 U12519 ( .A1(n10361), .A2(n11081), .ZN(n10360) );
  XNOR2_X1 U12520 ( .A(n11405), .B(n11404), .ZN(n14600) );
  NAND2_X1 U12521 ( .A1(n11402), .A2(n9754), .ZN(n11404) );
  OAI21_X1 U12522 ( .B1(n9897), .B2(n9888), .A(n9890), .ZN(n9887) );
  OR2_X1 U12523 ( .A1(n9892), .A2(n9891), .ZN(n9890) );
  OAI21_X1 U12524 ( .B1(n9897), .B2(n9889), .A(n9892), .ZN(n16249) );
  NAND2_X1 U12525 ( .A1(n11218), .A2(n9736), .ZN(n9889) );
  INV_X1 U12526 ( .A(n9894), .ZN(n16255) );
  OAI21_X1 U12527 ( .B1(n9897), .B2(n9895), .A(n11234), .ZN(n9894) );
  AND2_X1 U12528 ( .A1(n10081), .A2(n16311), .ZN(n16302) );
  NAND2_X1 U12529 ( .A1(n10128), .A2(n11165), .ZN(n16342) );
  INV_X1 U12530 ( .A(n11476), .ZN(n16350) );
  CLKBUF_X1 U12531 ( .A(n13892), .Z(n13893) );
  CLKBUF_X1 U12532 ( .A(n14111), .Z(n17207) );
  XNOR2_X1 U12533 ( .A(n11001), .B(n11000), .ZN(n9924) );
  INV_X1 U12534 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20317) );
  INV_X1 U12535 ( .A(n16820), .ZN(n19482) );
  INV_X1 U12536 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20293) );
  INV_X1 U12537 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17156) );
  AND2_X1 U12538 ( .A1(n16775), .A2(n16774), .ZN(n16797) );
  NOR2_X1 U12539 ( .A1(n16846), .A2(n20306), .ZN(n17239) );
  CLKBUF_X1 U12540 ( .A(n10948), .Z(n10857) );
  AOI21_X1 U12541 ( .B1(n16836), .B2(n17236), .A(n14233), .ZN(n16802) );
  OAI211_X1 U12542 ( .C1(n19732), .C2(n16815), .A(n16814), .B(n20133), .ZN(
        n19735) );
  OAI21_X1 U12543 ( .B1(n19761), .B2(n20306), .A(n19745), .ZN(n19764) );
  OAI21_X1 U12544 ( .B1(n19776), .B2(n19771), .A(n19770), .ZN(n19801) );
  OAI211_X1 U12545 ( .C1(n19921), .C2(n19917), .A(n20133), .B(n19916), .ZN(
        n19944) );
  OAI22_X1 U12546 ( .A1(n16142), .A2(n19640), .B1(n19632), .B2(n19642), .ZN(
        n20025) );
  AND2_X1 U12547 ( .A1(n16827), .A2(n16826), .ZN(n20030) );
  AND2_X1 U12548 ( .A1(n20045), .A2(n20041), .ZN(n20064) );
  INV_X1 U12549 ( .A(n20071), .ZN(n20126) );
  INV_X1 U12550 ( .A(n20085), .ZN(n20140) );
  AND2_X1 U12551 ( .A1(n20133), .A2(n19611), .ZN(n20141) );
  INV_X1 U12552 ( .A(n20090), .ZN(n20146) );
  AND2_X1 U12553 ( .A1(n20133), .A2(n19616), .ZN(n20147) );
  INV_X1 U12554 ( .A(n20095), .ZN(n20152) );
  AND2_X1 U12555 ( .A1(n20133), .A2(n19621), .ZN(n20153) );
  AND2_X1 U12556 ( .A1(n20133), .A2(n19626), .ZN(n20159) );
  AND2_X1 U12557 ( .A1(n19644), .A2(n9571), .ZN(n20164) );
  AND2_X1 U12558 ( .A1(n20133), .A2(n16828), .ZN(n20165) );
  AND2_X1 U12559 ( .A1(n20133), .A2(n19635), .ZN(n20173) );
  INV_X1 U12560 ( .A(n20025), .ZN(n20177) );
  OAI22_X1 U12561 ( .A1(n19643), .A2(n19642), .B1(n19641), .B2(n19640), .ZN(
        n20182) );
  INV_X1 U12562 ( .A(n15942), .ZN(n19417) );
  NOR2_X1 U12563 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n20319) );
  OR2_X1 U12564 ( .A1(n20190), .A2(P2_STATE_REG_0__SCAN_IN), .ZN(n20326) );
  NOR2_X1 U12565 ( .A1(n19184), .A2(n18173), .ZN(n19351) );
  NOR2_X1 U12566 ( .A1(n17455), .A2(n17380), .ZN(n17420) );
  NAND2_X1 U12567 ( .A1(n10200), .A2(n10198), .ZN(n17485) );
  OR2_X1 U12568 ( .A1(n10202), .A2(n10199), .ZN(n10198) );
  INV_X1 U12569 ( .A(n13602), .ZN(n10199) );
  AND2_X1 U12570 ( .A1(n10206), .A2(n17388), .ZN(n17486) );
  NOR2_X2 U12571 ( .A1(n19211), .A2(n13614), .ZN(n17658) );
  INV_X1 U12572 ( .A(n17658), .ZN(n17729) );
  INV_X1 U12573 ( .A(n17644), .ZN(n17721) );
  NOR2_X1 U12574 ( .A1(n17865), .A2(n17885), .ZN(n17890) );
  INV_X1 U12575 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17604) );
  INV_X1 U12576 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n21250) );
  INV_X2 U12577 ( .A(n18016), .ZN(n18013) );
  NOR2_X1 U12578 ( .A1(n18041), .A2(n9960), .ZN(n18029) );
  NOR2_X1 U12579 ( .A1(n18041), .A2(n18201), .ZN(n18037) );
  NOR2_X1 U12580 ( .A1(n18783), .A2(n18056), .ZN(n18051) );
  NAND2_X1 U12581 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n18051), .ZN(n18050) );
  NOR2_X1 U12582 ( .A1(n18019), .A2(n9967), .ZN(n18057) );
  NAND2_X1 U12583 ( .A1(n18057), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n18056) );
  NOR2_X1 U12584 ( .A1(n18188), .A2(n18071), .ZN(n18067) );
  NOR2_X1 U12585 ( .A1(n18184), .A2(n18078), .ZN(n18077) );
  NOR2_X1 U12586 ( .A1(n18085), .A2(n18238), .ZN(n14164) );
  NAND2_X1 U12587 ( .A1(n14164), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n18019) );
  INV_X1 U12588 ( .A(n18120), .ZN(n18102) );
  AND2_X1 U12589 ( .A1(n11986), .A2(n11985), .ZN(n18110) );
  AND4_X1 U12590 ( .A1(n11984), .A2(n11983), .A3(n11982), .A4(n11981), .ZN(
        n11985) );
  INV_X1 U12591 ( .A(n12218), .ZN(n18113) );
  NOR3_X1 U12592 ( .A1(n18211), .A2(n18209), .A3(n18020), .ZN(n18121) );
  NAND2_X1 U12593 ( .A1(n9955), .A2(n19214), .ZN(n14009) );
  NAND2_X1 U12594 ( .A1(n9956), .A2(n9700), .ZN(n9955) );
  INV_X1 U12595 ( .A(n18123), .ZN(n18104) );
  NOR2_X1 U12596 ( .A1(n18173), .A2(n18127), .ZN(n18164) );
  INV_X1 U12597 ( .A(n18164), .ZN(n18172) );
  NOR2_X1 U12598 ( .A1(n18173), .A2(n19212), .ZN(n18228) );
  NAND2_X2 U12599 ( .A1(n18177), .A2(n18176), .ZN(n18234) );
  INV_X1 U12600 ( .A(n18230), .ZN(n18235) );
  INV_X1 U12601 ( .A(n18228), .ZN(n18237) );
  INV_X1 U12602 ( .A(n16877), .ZN(n17255) );
  CLKBUF_X1 U12603 ( .A(n16908), .Z(n18239) );
  INV_X1 U12604 ( .A(n18391), .ZN(n18377) );
  OAI21_X1 U12605 ( .B1(n18350), .B2(n18573), .A(n18329), .ZN(n18347) );
  INV_X1 U12606 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n18402) );
  NAND2_X1 U12607 ( .A1(n16894), .A2(n16893), .ZN(n18438) );
  OR2_X1 U12608 ( .A1(n16990), .A2(n18391), .ZN(n18426) );
  INV_X2 U12609 ( .A(n18495), .ZN(n18478) );
  INV_X1 U12610 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18477) );
  INV_X1 U12611 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18496) );
  INV_X1 U12612 ( .A(n16992), .ZN(n18857) );
  NAND2_X1 U12613 ( .A1(n17104), .A2(n10094), .ZN(n17105) );
  NAND2_X1 U12614 ( .A1(n17040), .A2(n10095), .ZN(n10094) );
  INV_X1 U12615 ( .A(n18593), .ZN(n17088) );
  AND2_X1 U12616 ( .A1(n17056), .A2(n18500), .ZN(n18532) );
  NAND2_X1 U12617 ( .A1(n12015), .A2(n10415), .ZN(n18344) );
  INV_X1 U12618 ( .A(n18672), .ZN(n18689) );
  NAND2_X1 U12619 ( .A1(n12012), .A2(n10212), .ZN(n14253) );
  INV_X1 U12620 ( .A(n18728), .ZN(n18629) );
  NAND2_X1 U12621 ( .A1(n11935), .A2(n11934), .ZN(n18470) );
  OR2_X1 U12622 ( .A1(n11935), .A2(n11934), .ZN(n18471) );
  INV_X1 U12623 ( .A(n18729), .ZN(n18701) );
  INV_X1 U12624 ( .A(n18712), .ZN(n19179) );
  INV_X1 U12625 ( .A(n12186), .ZN(n9770) );
  INV_X1 U12626 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21323) );
  INV_X1 U12627 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n19188) );
  INV_X1 U12628 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14105) );
  NOR2_X1 U12629 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19322), .ZN(
        n19209) );
  INV_X1 U12630 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n19322) );
  AND2_X2 U12631 ( .A1(n13555), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20584)
         );
  OAI211_X1 U12633 ( .C1(n15341), .C2(n20338), .A(n9674), .B(n13277), .ZN(
        P1_U2971) );
  NOR2_X1 U12634 ( .A1(n15146), .A2(n9868), .ZN(n9867) );
  OAI21_X1 U12635 ( .B1(n15324), .B2(n20573), .A(n10175), .ZN(P1_U3001) );
  NAND2_X1 U12636 ( .A1(n15321), .A2(n15322), .ZN(n10235) );
  NAND2_X1 U12637 ( .A1(n15469), .A2(n20563), .ZN(n15475) );
  NAND2_X1 U12638 ( .A1(n10181), .A2(n10177), .ZN(P2_U2825) );
  INV_X1 U12639 ( .A(n14607), .ZN(n10181) );
  NOR2_X1 U12640 ( .A1(n9687), .A2(n10178), .ZN(n10177) );
  OAI211_X1 U12641 ( .C1(n15616), .C2(n15615), .A(n9733), .B(n10121), .ZN(
        P2_U2827) );
  OR4_X1 U12642 ( .A1(n13594), .A2(n13593), .A3(n13592), .A4(n13591), .ZN(
        P2_U2842) );
  AOI21_X1 U12643 ( .B1(n19413), .B2(n9973), .A(n15936), .ZN(n15937) );
  INV_X1 U12644 ( .A(n11567), .ZN(n9973) );
  OAI21_X1 U12645 ( .B1(n16079), .B2(n16066), .A(n9863), .ZN(P2_U2857) );
  NAND2_X1 U12646 ( .A1(n11860), .A2(n19429), .ZN(n11861) );
  AOI21_X1 U12647 ( .B1(n16088), .B2(n19477), .A(n16087), .ZN(n16089) );
  NAND2_X1 U12648 ( .A1(n11520), .A2(n9627), .ZN(n11492) );
  NAND2_X1 U12649 ( .A1(n11519), .A2(n19577), .ZN(n11493) );
  NAND2_X1 U12650 ( .A1(n11457), .A2(n9702), .ZN(P2_U2985) );
  OR2_X1 U12651 ( .A1(n11510), .A2(n11509), .ZN(P2_U2997) );
  AOI21_X1 U12652 ( .B1(n16568), .B2(n9627), .A(n11507), .ZN(n11508) );
  INV_X1 U12653 ( .A(n9804), .ZN(n9803) );
  OAI21_X1 U12654 ( .B1(n16624), .B2(n19574), .A(n16330), .ZN(n9804) );
  NAND2_X1 U12655 ( .A1(n11420), .A2(n17209), .ZN(n11438) );
  NAND2_X1 U12656 ( .A1(n11863), .A2(n17209), .ZN(n10043) );
  INV_X1 U12657 ( .A(n17361), .ZN(n17355) );
  OR2_X1 U12658 ( .A1(n17402), .A2(n17403), .ZN(n10207) );
  AND2_X1 U12659 ( .A1(n16889), .A2(n10087), .ZN(n9982) );
  INV_X1 U12660 ( .A(n9981), .ZN(n9979) );
  AND2_X1 U12661 ( .A1(n12256), .A2(n12255), .ZN(n12257) );
  NAND2_X1 U12662 ( .A1(n10326), .A2(n11327), .ZN(n15809) );
  AND4_X1 U12663 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n9628)
         );
  AND2_X1 U12664 ( .A1(n9654), .A2(n16451), .ZN(n9629) );
  INV_X2 U12665 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n10368) );
  INV_X1 U12666 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n10955) );
  CLKBUF_X3 U12667 ( .A(n11994), .Z(n17973) );
  NAND2_X1 U12668 ( .A1(n10241), .A2(n10240), .ZN(n14828) );
  NAND2_X1 U12669 ( .A1(n11173), .A2(n9679), .ZN(n9630) );
  INV_X1 U12670 ( .A(n13319), .ZN(n13396) );
  OR2_X1 U12671 ( .A1(n14749), .A2(n10388), .ZN(n9631) );
  AND2_X1 U12672 ( .A1(n12468), .A2(n17135), .ZN(n9632) );
  NAND2_X1 U12673 ( .A1(n10128), .A2(n9677), .ZN(n9633) );
  INV_X1 U12674 ( .A(n10884), .ZN(n20314) );
  NAND2_X1 U12675 ( .A1(n11005), .A2(n11004), .ZN(n11577) );
  CLKBUF_X3 U12676 ( .A(n12383), .Z(n13088) );
  AND2_X1 U12677 ( .A1(n13452), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13443) );
  NAND2_X1 U12678 ( .A1(n14240), .A2(n11612), .ZN(n16040) );
  NAND2_X1 U12679 ( .A1(n10296), .A2(n10297), .ZN(n16030) );
  NAND2_X1 U12680 ( .A1(n11475), .A2(n9629), .ZN(n16212) );
  AND2_X1 U12681 ( .A1(n11158), .A2(n10227), .ZN(n11166) );
  NOR2_X1 U12682 ( .A1(n14422), .A2(n10312), .ZN(n11501) );
  NOR2_X1 U12683 ( .A1(n14422), .A2(n10314), .ZN(n11500) );
  NOR2_X1 U12684 ( .A1(n15683), .A2(n10258), .ZN(n15646) );
  NAND2_X1 U12685 ( .A1(n11468), .A2(n15706), .ZN(n9634) );
  AND2_X1 U12686 ( .A1(n10391), .A2(n12879), .ZN(n9635) );
  INV_X1 U12687 ( .A(n10029), .ZN(n16256) );
  NAND2_X1 U12688 ( .A1(n11476), .A2(n9655), .ZN(n10029) );
  AND2_X1 U12689 ( .A1(n11059), .A2(n11058), .ZN(n9636) );
  NAND2_X1 U12690 ( .A1(n9964), .A2(n11663), .ZN(n16017) );
  NAND2_X2 U12691 ( .A1(n9774), .A2(n9772), .ZN(n10889) );
  OR2_X1 U12692 ( .A1(n13587), .A2(n13588), .ZN(n13586) );
  AND2_X1 U12693 ( .A1(n9679), .A2(n11211), .ZN(n9637) );
  NAND2_X1 U12694 ( .A1(n11475), .A2(n9756), .ZN(n11419) );
  NAND2_X1 U12695 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13446) );
  AND3_X1 U12696 ( .A1(n9708), .A2(n12068), .A3(n9961), .ZN(n9638) );
  OR2_X1 U12697 ( .A1(n9569), .A2(n13207), .ZN(n13208) );
  NOR2_X1 U12698 ( .A1(n10131), .A2(n10130), .ZN(n10129) );
  OR2_X1 U12699 ( .A1(n14829), .A2(n14853), .ZN(n9639) );
  OR2_X1 U12700 ( .A1(n10328), .A2(n11460), .ZN(n9640) );
  NAND2_X1 U12701 ( .A1(n11105), .A2(n11100), .ZN(n10225) );
  AND2_X1 U12702 ( .A1(n16248), .A2(n9736), .ZN(n9641) );
  INV_X1 U12703 ( .A(n10319), .ZN(n11421) );
  AND3_X1 U12704 ( .A1(n10883), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n10891), 
        .ZN(n9642) );
  AND2_X1 U12705 ( .A1(n10015), .A2(n14570), .ZN(n9643) );
  AND2_X1 U12706 ( .A1(n10374), .A2(n10381), .ZN(n9644) );
  INV_X1 U12707 ( .A(n9569), .ZN(n9952) );
  OR2_X1 U12708 ( .A1(n15600), .A2(n10189), .ZN(n9645) );
  NAND2_X1 U12709 ( .A1(n10306), .A2(n11313), .ZN(n14288) );
  AND2_X1 U12710 ( .A1(n11037), .A2(n9741), .ZN(n9646) );
  AND2_X1 U12711 ( .A1(n10117), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9647) );
  NOR2_X1 U12712 ( .A1(n11835), .A2(n11856), .ZN(n9648) );
  AND2_X1 U12713 ( .A1(n10297), .A2(n10295), .ZN(n9649) );
  AND2_X1 U12714 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n9650) );
  AND4_X1 U12715 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .A3(P3_EAX_REG_1__SCAN_IN), .A4(P3_EAX_REG_0__SCAN_IN), .ZN(n9651) );
  OR2_X1 U12716 ( .A1(n12013), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n9652) );
  AND2_X1 U12717 ( .A1(n9650), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9653) );
  AND2_X1 U12718 ( .A1(n11080), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9654) );
  AND2_X1 U12719 ( .A1(n10933), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9655) );
  AND2_X1 U12720 ( .A1(n9629), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9656) );
  AND2_X4 U12721 ( .A1(n12277), .A2(n10082), .ZN(n12461) );
  AND2_X2 U12722 ( .A1(n10446), .A2(n11692), .ZN(n10507) );
  NAND2_X1 U12723 ( .A1(n13761), .A2(n11876), .ZN(n10404) );
  NOR2_X1 U12724 ( .A1(n12601), .A2(n21070), .ZN(n12668) );
  OR3_X1 U12725 ( .A1(n13455), .A2(n10109), .A3(n10108), .ZN(n9658) );
  NAND2_X1 U12726 ( .A1(n13881), .A2(n12522), .ZN(n13947) );
  INV_X1 U12727 ( .A(n12417), .ZN(n20622) );
  INV_X1 U12728 ( .A(n11937), .ZN(n14037) );
  INV_X2 U12729 ( .A(n12101), .ZN(n17972) );
  AND2_X2 U12730 ( .A1(n14215), .A2(n10441), .ZN(n10482) );
  AND2_X2 U12731 ( .A1(n11694), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10578) );
  NOR2_X1 U12732 ( .A1(n18407), .A2(n18630), .ZN(n9659) );
  AND2_X1 U12733 ( .A1(n10367), .A2(n12468), .ZN(n9660) );
  OR3_X1 U12734 ( .A1(n18041), .A2(n9960), .A3(n18205), .ZN(n9661) );
  BUF_X4 U12735 ( .A(n10902), .Z(n11287) );
  AND2_X1 U12736 ( .A1(n11014), .A2(n11023), .ZN(n11052) );
  NAND2_X1 U12737 ( .A1(n12740), .A2(n12739), .ZN(n14849) );
  NOR2_X1 U12738 ( .A1(n13146), .A2(n12543), .ZN(n9662) );
  INV_X1 U12739 ( .A(n13447), .ZN(n10114) );
  NOR2_X1 U12740 ( .A1(n14749), .A2(n10387), .ZN(n9663) );
  NAND2_X1 U12741 ( .A1(n10265), .A2(n10739), .ZN(n11542) );
  OR2_X1 U12742 ( .A1(n11104), .A2(n10225), .ZN(n11135) );
  OR2_X1 U12743 ( .A1(n14675), .A2(n10394), .ZN(n9664) );
  NAND2_X1 U12744 ( .A1(n12611), .A2(n9814), .ZN(n13170) );
  NOR2_X1 U12745 ( .A1(n9593), .A2(n10392), .ZN(n14785) );
  NOR2_X1 U12746 ( .A1(n13587), .A2(n10260), .ZN(n9665) );
  AND2_X1 U12747 ( .A1(n15649), .A2(n11379), .ZN(n15632) );
  AND2_X1 U12748 ( .A1(n11778), .A2(n10285), .ZN(n9666) );
  AND2_X1 U12749 ( .A1(n11468), .A2(n10324), .ZN(n9667) );
  NOR2_X1 U12750 ( .A1(n11543), .A2(n11544), .ZN(n11467) );
  NOR2_X1 U12751 ( .A1(n10889), .A2(n10838), .ZN(n9668) );
  OR2_X1 U12752 ( .A1(n11104), .A2(n11097), .ZN(n9669) );
  AND2_X1 U12753 ( .A1(n9925), .A2(n9883), .ZN(n9670) );
  OR2_X1 U12754 ( .A1(n9660), .A2(n10050), .ZN(n9671) );
  INV_X1 U12755 ( .A(n12679), .ZN(n15572) );
  NOR3_X1 U12756 ( .A1(n13455), .A2(n10110), .A3(n16328), .ZN(n13440) );
  AND2_X1 U12757 ( .A1(n16304), .A2(n16293), .ZN(n9672) );
  AND2_X1 U12758 ( .A1(n9672), .A2(n10191), .ZN(n9673) );
  AND2_X1 U12759 ( .A1(n14746), .A2(n10248), .ZN(n14683) );
  XNOR2_X1 U12760 ( .A(n11005), .B(n11007), .ZN(n11572) );
  AND2_X1 U12761 ( .A1(n15130), .A2(n9797), .ZN(n9675) );
  AND3_X1 U12762 ( .A1(n11053), .A2(n11060), .A3(n11061), .ZN(n9676) );
  AND2_X1 U12763 ( .A1(n11165), .A2(n10127), .ZN(n9677) );
  NAND2_X1 U12764 ( .A1(n10346), .A2(n10350), .ZN(n16375) );
  AND2_X1 U12765 ( .A1(n11449), .A2(n11485), .ZN(n9678) );
  AND2_X1 U12766 ( .A1(n10232), .A2(n10409), .ZN(n9679) );
  OR2_X1 U12767 ( .A1(n14675), .A2(n10396), .ZN(n13294) );
  NOR2_X1 U12768 ( .A1(n11110), .A2(n11109), .ZN(n9680) );
  NAND2_X1 U12769 ( .A1(n10884), .A2(n20311), .ZN(n11088) );
  NAND2_X1 U12770 ( .A1(n10134), .A2(n16236), .ZN(n16215) );
  NAND2_X1 U12771 ( .A1(n11417), .A2(n11416), .ZN(n9681) );
  NAND2_X1 U12772 ( .A1(n15114), .A2(n15113), .ZN(n9682) );
  NAND2_X1 U12773 ( .A1(n10365), .A2(n9660), .ZN(n12656) );
  AND4_X1 U12774 ( .A1(n11931), .A2(n11930), .A3(n11929), .A4(n11928), .ZN(
        n9683) );
  AND2_X1 U12775 ( .A1(n12538), .A2(n10368), .ZN(n9684) );
  NAND2_X1 U12776 ( .A1(n10885), .A2(n11088), .ZN(n10895) );
  NAND2_X1 U12777 ( .A1(n12680), .A2(n12690), .ZN(n20586) );
  OR2_X1 U12778 ( .A1(n15861), .A2(n16370), .ZN(n9685) );
  INV_X1 U12779 ( .A(n16333), .ZN(n10331) );
  INV_X1 U12780 ( .A(n18357), .ZN(n18365) );
  NAND2_X1 U12781 ( .A1(n10270), .A2(n10268), .ZN(n14634) );
  INV_X1 U12782 ( .A(n10277), .ZN(n11007) );
  AND2_X1 U12783 ( .A1(n11010), .A2(n11030), .ZN(n9686) );
  INV_X1 U12784 ( .A(n9569), .ZN(n10374) );
  AND2_X1 U12785 ( .A1(n14612), .A2(n19384), .ZN(n9687) );
  NAND2_X1 U12786 ( .A1(n14004), .A2(n11589), .ZN(n14110) );
  AND2_X1 U12787 ( .A1(n19185), .A2(n19222), .ZN(n9688) );
  AND2_X1 U12788 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9689) );
  AND2_X1 U12789 ( .A1(n9918), .A2(n9917), .ZN(n9690) );
  OR2_X1 U12790 ( .A1(n11251), .A2(n16480), .ZN(n9691) );
  INV_X1 U12791 ( .A(n11078), .ZN(n10039) );
  AND2_X1 U12792 ( .A1(n10370), .A2(n10009), .ZN(n9692) );
  NAND2_X1 U12793 ( .A1(n11591), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n9693) );
  AND2_X1 U12794 ( .A1(n12509), .A2(n10368), .ZN(n9694) );
  INV_X1 U12795 ( .A(n9988), .ZN(n17040) );
  AND2_X1 U12796 ( .A1(n10821), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n9695) );
  AND2_X1 U12797 ( .A1(n11488), .A2(n11485), .ZN(n9696) );
  OR2_X1 U12798 ( .A1(n9571), .A2(n11176), .ZN(n9697) );
  AND2_X1 U12799 ( .A1(n10265), .A2(n10264), .ZN(n9698) );
  AND2_X1 U12800 ( .A1(n15130), .A2(n9952), .ZN(n9699) );
  NAND2_X1 U12801 ( .A1(n13928), .A2(n13927), .ZN(n9700) );
  NAND2_X1 U12802 ( .A1(n11476), .A2(n11080), .ZN(n16233) );
  XNOR2_X1 U12804 ( .A(n11032), .B(n11031), .ZN(n16725) );
  INV_X1 U12805 ( .A(n10350), .ZN(n10349) );
  AND2_X1 U12806 ( .A1(n10356), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9701) );
  AND2_X1 U12807 ( .A1(n9976), .A2(n9974), .ZN(n9702) );
  AND2_X1 U12808 ( .A1(n10212), .A2(n18357), .ZN(n9703) );
  AND2_X1 U12809 ( .A1(n9637), .A2(n9935), .ZN(n9704) );
  AND2_X1 U12810 ( .A1(n9926), .A2(n9925), .ZN(n9705) );
  AND2_X1 U12811 ( .A1(n19593), .A2(n10277), .ZN(n11024) );
  AND2_X1 U12812 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11879) );
  AND2_X1 U12813 ( .A1(n14145), .A2(n12677), .ZN(n9706) );
  NAND2_X1 U12814 ( .A1(n15896), .A2(n11142), .ZN(n9707) );
  AND4_X1 U12815 ( .A1(n12073), .A2(n12072), .A3(n12071), .A4(n12070), .ZN(
        n9708) );
  INV_X1 U12816 ( .A(n10242), .ZN(n10240) );
  NAND2_X1 U12817 ( .A1(n14862), .A2(n10243), .ZN(n10242) );
  BUF_X1 U12818 ( .A(n12441), .Z(n17135) );
  INV_X1 U12819 ( .A(n11152), .ZN(n9902) );
  OR2_X1 U12820 ( .A1(n14430), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9709) );
  NOR2_X1 U12821 ( .A1(n11233), .A2(n11464), .ZN(n11234) );
  AND2_X1 U12822 ( .A1(n10374), .A2(n10376), .ZN(n9710) );
  OR2_X1 U12823 ( .A1(n12406), .A2(n10368), .ZN(n12543) );
  INV_X1 U12824 ( .A(n10022), .ZN(n15342) );
  NOR2_X1 U12825 ( .A1(n15362), .A2(n14575), .ZN(n10022) );
  NAND2_X1 U12826 ( .A1(n11173), .A2(n9704), .ZN(n9936) );
  AND2_X1 U12827 ( .A1(n12431), .A2(n13215), .ZN(n9711) );
  NAND2_X1 U12828 ( .A1(n11498), .A2(n11496), .ZN(n9712) );
  NAND2_X1 U12829 ( .A1(n10257), .A2(n10750), .ZN(n15663) );
  INV_X1 U12830 ( .A(n10308), .ZN(n10307) );
  NOR2_X1 U12831 ( .A1(n14321), .A2(n14289), .ZN(n10308) );
  AND2_X1 U12832 ( .A1(n10113), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9713) );
  NAND2_X1 U12833 ( .A1(n10905), .A2(n10904), .ZN(n10940) );
  OR2_X1 U12834 ( .A1(n11461), .A2(n10080), .ZN(n9714) );
  AND2_X1 U12835 ( .A1(n13352), .A2(n13351), .ZN(n14927) );
  NAND2_X1 U12836 ( .A1(n11155), .A2(n11260), .ZN(n11158) );
  AND3_X1 U12837 ( .A1(n10813), .A2(n9801), .A3(n9802), .ZN(n9715) );
  AND2_X1 U12838 ( .A1(n9633), .A2(n11459), .ZN(n9716) );
  AND2_X1 U12839 ( .A1(n15202), .A2(n10372), .ZN(n9717) );
  AND2_X1 U12840 ( .A1(n10943), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9718) );
  AND2_X1 U12841 ( .A1(n10892), .A2(n10890), .ZN(n9719) );
  XNOR2_X1 U12842 ( .A(n10889), .B(n10902), .ZN(n10863) );
  AOI21_X1 U12843 ( .B1(n11297), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n10997), .ZN(n11296) );
  AND2_X1 U12844 ( .A1(n11144), .A2(n10339), .ZN(n9720) );
  AND2_X1 U12845 ( .A1(n10883), .A2(n10891), .ZN(n9721) );
  AND2_X1 U12846 ( .A1(n12518), .A2(n12519), .ZN(n9722) );
  AND2_X1 U12847 ( .A1(n9908), .A2(n20306), .ZN(n9723) );
  AND2_X1 U12848 ( .A1(n16321), .A2(n16331), .ZN(n9724) );
  AOI21_X1 U12849 ( .B1(n15734), .B2(n17215), .A(n11559), .ZN(n11560) );
  AND2_X1 U12850 ( .A1(n19593), .A2(n11007), .ZN(n11015) );
  AND2_X1 U12851 ( .A1(n9673), .A2(n16285), .ZN(n9725) );
  AND2_X1 U12852 ( .A1(n10350), .A2(n11078), .ZN(n9726) );
  AND2_X1 U12853 ( .A1(n11077), .A2(n11078), .ZN(n16376) );
  INV_X1 U12854 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16399) );
  NAND2_X1 U12855 ( .A1(n11698), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n9727) );
  INV_X1 U12856 ( .A(n9983), .ZN(n9980) );
  NAND2_X1 U12857 ( .A1(n12036), .A2(n12037), .ZN(n9983) );
  NAND3_X1 U12858 ( .A1(n14430), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n9728) );
  BUF_X2 U12859 ( .A(n12720), .Z(n13502) );
  INV_X1 U12860 ( .A(n19426), .ZN(n16066) );
  NOR2_X1 U12861 ( .A1(n14296), .A2(n10245), .ZN(n14441) );
  NAND4_X1 U12862 ( .A1(n10356), .A2(n10358), .A3(n10357), .A4(n10946), .ZN(
        n9729) );
  INV_X1 U12863 ( .A(n17226), .ZN(n17209) );
  NAND2_X1 U12864 ( .A1(n11409), .A2(n20299), .ZN(n17226) );
  BUF_X1 U12865 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n10980) );
  NOR2_X1 U12866 ( .A1(n16040), .A2(n16041), .ZN(n16033) );
  AND2_X1 U12867 ( .A1(n10296), .A2(n9649), .ZN(n9730) );
  NAND2_X1 U12868 ( .A1(n11303), .A2(n11302), .ZN(n14243) );
  OR2_X1 U12869 ( .A1(n14422), .A2(n16049), .ZN(n9731) );
  INV_X2 U12870 ( .A(n19429), .ZN(n16073) );
  AND2_X1 U12871 ( .A1(n11858), .A2(n17236), .ZN(n19429) );
  INV_X1 U12872 ( .A(n12689), .ZN(n10369) );
  INV_X1 U12873 ( .A(n11736), .ZN(n9861) );
  NOR2_X1 U12874 ( .A1(n14266), .A2(n10307), .ZN(n14322) );
  NAND2_X1 U12875 ( .A1(n10238), .A2(n13346), .ZN(n15003) );
  AND2_X1 U12876 ( .A1(n13008), .A2(n13007), .ZN(n9732) );
  AND2_X2 U12877 ( .A1(n11409), .A2(n20298), .ZN(n17224) );
  OR3_X1 U12878 ( .A1(n15612), .A2(n15611), .A3(n19386), .ZN(n9733) );
  OR3_X1 U12879 ( .A1(n9861), .A2(n11738), .A3(n16009), .ZN(n9734) );
  INV_X1 U12880 ( .A(n15675), .ZN(n11371) );
  AND2_X1 U12881 ( .A1(n15633), .A2(n10317), .ZN(n9735) );
  OR2_X1 U12882 ( .A1(n11239), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9736) );
  AND2_X1 U12883 ( .A1(n16265), .A2(n11458), .ZN(n9737) );
  AND3_X1 U12884 ( .A1(n10061), .A2(n9721), .A3(n10895), .ZN(n10953) );
  NAND2_X1 U12885 ( .A1(n14502), .A2(n14482), .ZN(n20573) );
  INV_X1 U12886 ( .A(n20573), .ZN(n20563) );
  INV_X1 U12887 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17709) );
  OR2_X1 U12888 ( .A1(n14896), .A2(n14898), .ZN(n14897) );
  INV_X1 U12889 ( .A(n14897), .ZN(n10241) );
  INV_X1 U12890 ( .A(n15825), .ZN(n10326) );
  NOR2_X1 U12891 ( .A1(n15613), .A2(n10123), .ZN(n9738) );
  AND2_X1 U12892 ( .A1(n13139), .A2(n14494), .ZN(n9739) );
  AND2_X1 U12893 ( .A1(n17161), .A2(n13920), .ZN(n15200) );
  INV_X1 U12894 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13215) );
  AND2_X1 U12895 ( .A1(n9735), .A2(n10316), .ZN(n9740) );
  INV_X1 U12896 ( .A(n11142), .ZN(n11063) );
  OR2_X1 U12897 ( .A1(n10568), .A2(n10567), .ZN(n11142) );
  BUF_X1 U12898 ( .A(n12416), .Z(n20607) );
  AND2_X1 U12899 ( .A1(n11093), .A2(n11092), .ZN(n9741) );
  OR2_X1 U12900 ( .A1(n11652), .A2(n11651), .ZN(n16026) );
  AND3_X1 U12901 ( .A1(n12738), .A2(n12737), .A3(n12736), .ZN(n14926) );
  AND2_X1 U12902 ( .A1(n15614), .A2(n9738), .ZN(n9742) );
  OR2_X1 U12903 ( .A1(n10258), .A2(n10256), .ZN(n9743) );
  INV_X1 U12904 ( .A(n9937), .ZN(n16224) );
  NAND2_X1 U12905 ( .A1(n11270), .A2(n16468), .ZN(n9937) );
  OR2_X1 U12906 ( .A1(n10260), .A2(n10262), .ZN(n9744) );
  NAND2_X1 U12907 ( .A1(n14240), .A2(n9860), .ZN(n16022) );
  NOR2_X2 U12908 ( .A1(n12417), .A2(n21070), .ZN(n12823) );
  INV_X1 U12909 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16328) );
  AND2_X1 U12910 ( .A1(n12407), .A2(n17135), .ZN(n13858) );
  AND2_X1 U12911 ( .A1(n13479), .A2(n9653), .ZN(n9745) );
  AND2_X1 U12912 ( .A1(n10238), .A2(n10237), .ZN(n9746) );
  NOR2_X1 U12913 ( .A1(n17472), .A2(n17695), .ZN(n9747) );
  AND2_X1 U12914 ( .A1(n11062), .A2(n11142), .ZN(n9748) );
  NAND2_X1 U12915 ( .A1(n13462), .A2(n10117), .ZN(n10120) );
  OR2_X1 U12916 ( .A1(n10537), .A2(n10536), .ZN(n11092) );
  NAND2_X1 U12917 ( .A1(n12511), .A2(n13215), .ZN(n9749) );
  AND3_X1 U12918 ( .A1(n12878), .A2(n12877), .A3(n12876), .ZN(n14813) );
  AND2_X1 U12919 ( .A1(n9649), .A2(n16026), .ZN(n9750) );
  INV_X1 U12920 ( .A(n18288), .ZN(n10203) );
  INV_X1 U12921 ( .A(n16285), .ZN(n10192) );
  INV_X1 U12922 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10112) );
  OR2_X1 U12923 ( .A1(n16962), .A2(n10217), .ZN(n9751) );
  INV_X1 U12924 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n13438) );
  INV_X1 U12925 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12681) );
  NAND2_X1 U12926 ( .A1(n10741), .A2(n10740), .ZN(n9752) );
  INV_X1 U12927 ( .A(n16378), .ZN(n11293) );
  AND4_X1 U12928 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n9753) );
  AND2_X1 U12929 ( .A1(n11401), .A2(n9845), .ZN(n9754) );
  AND2_X1 U12930 ( .A1(n10767), .A2(n10766), .ZN(n9755) );
  AND2_X1 U12931 ( .A1(n9656), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9756) );
  INV_X1 U12932 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10110) );
  INV_X1 U12933 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10118) );
  OR2_X1 U12934 ( .A1(n9652), .A2(n12014), .ZN(n9757) );
  INV_X1 U12935 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18384) );
  NAND2_X1 U12936 ( .A1(n13459), .A2(n9673), .ZN(n10193) );
  AND2_X1 U12937 ( .A1(n9997), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n9758) );
  NOR2_X1 U12938 ( .A1(n16000), .A2(n15991), .ZN(n9759) );
  NOR2_X1 U12939 ( .A1(n14120), .A2(n9758), .ZN(n9760) );
  AND3_X1 U12940 ( .A1(n10701), .A2(n10700), .A3(n10699), .ZN(n13588) );
  AND2_X1 U12941 ( .A1(n9653), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9761) );
  NAND2_X1 U12942 ( .A1(n16010), .A2(n10229), .ZN(n9762) );
  INV_X1 U12943 ( .A(n19308), .ZN(n19347) );
  NOR2_X2 U12944 ( .A1(n17353), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n19308) );
  INV_X1 U12945 ( .A(n15927), .ZN(n10182) );
  NAND2_X1 U12946 ( .A1(n13926), .A2(n12062), .ZN(n19333) );
  INV_X1 U12947 ( .A(n19333), .ZN(n9771) );
  AND2_X1 U12948 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14272) );
  AND2_X1 U12949 ( .A1(n14563), .A2(n15335), .ZN(n9763) );
  INV_X1 U12950 ( .A(n10378), .ZN(n10377) );
  NAND2_X1 U12951 ( .A1(n13209), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10378) );
  INV_X1 U12952 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n9935) );
  INV_X1 U12953 ( .A(n13211), .ZN(n10011) );
  AND2_X1 U12954 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9764) );
  INV_X1 U12955 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10255) );
  INV_X1 U12956 ( .A(n15325), .ZN(n10381) );
  XOR2_X1 U12957 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(n9765) );
  INV_X1 U12958 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10127) );
  INV_X1 U12959 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10119) );
  AND2_X1 U12960 ( .A1(n10362), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9766) );
  NAND4_X1 U12961 ( .A1(n19349), .A2(n19338), .A3(n21312), .A4(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n9767) );
  INV_X1 U12962 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n19349) );
  INV_X1 U12963 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n19338) );
  AOI22_X2 U12964 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n20629), .B1(DATAI_31_), 
        .B2(n20628), .ZN(n21132) );
  AOI22_X2 U12965 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20629), .B1(DATAI_30_), 
        .B2(n20628), .ZN(n21121) );
  NOR2_X2 U12966 ( .A1(n18658), .A2(n19179), .ZN(n18554) );
  OR2_X2 U12967 ( .A1(n19183), .A2(n19177), .ZN(n9769) );
  OR2_X2 U12968 ( .A1(n18593), .A2(n9770), .ZN(n19183) );
  OR2_X2 U12969 ( .A1(n12147), .A2(n13722), .ZN(n12150) );
  NAND2_X4 U12970 ( .A1(n17094), .A2(n14105), .ZN(n12117) );
  AND2_X2 U12971 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13760) );
  NAND2_X1 U12972 ( .A1(n16414), .A2(n16415), .ZN(n11045) );
  XNOR2_X2 U12973 ( .A(n11050), .B(n11092), .ZN(n16414) );
  NAND4_X1 U12974 ( .A1(n10469), .A2(n10471), .A3(n10468), .A4(n10470), .ZN(
        n9773) );
  NAND4_X1 U12975 ( .A1(n9776), .A2(n10465), .A3(n10467), .A4(n10466), .ZN(
        n9775) );
  NAND2_X1 U12976 ( .A1(n9778), .A2(n9780), .ZN(n10942) );
  NAND4_X1 U12977 ( .A1(n9719), .A2(n9909), .A3(n9779), .A4(n10891), .ZN(n9778) );
  NAND2_X1 U12978 ( .A1(n16279), .A2(n9781), .ZN(P2_U2993) );
  AND2_X1 U12979 ( .A1(n9782), .A2(n16258), .ZN(n16530) );
  NAND2_X1 U12980 ( .A1(n16273), .A2(n16523), .ZN(n9782) );
  NAND3_X1 U12981 ( .A1(n9786), .A2(n9784), .A3(n9783), .ZN(n11475) );
  NAND3_X1 U12982 ( .A1(n16405), .A2(n10347), .A3(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n9783) );
  NAND2_X2 U12983 ( .A1(n9789), .A2(n12558), .ZN(n12679) );
  NAND2_X1 U12984 ( .A1(n15572), .A2(n12678), .ZN(n12680) );
  NAND3_X1 U12985 ( .A1(n9728), .A2(n10144), .A3(n9790), .ZN(n17163) );
  INV_X1 U12986 ( .A(n13167), .ZN(n9791) );
  NAND2_X1 U12987 ( .A1(n9799), .A2(n9715), .ZN(n9798) );
  NAND2_X1 U12988 ( .A1(n11699), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n9800) );
  NAND2_X1 U12989 ( .A1(n11694), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n9801) );
  NAND2_X1 U12990 ( .A1(n9805), .A2(n9803), .ZN(P2_U3001) );
  NAND2_X1 U12991 ( .A1(n16614), .A2(n19577), .ZN(n9805) );
  NOR2_X1 U12992 ( .A1(n16309), .A2(n16602), .ZN(n16325) );
  NAND4_X1 U12993 ( .A1(n9809), .A2(n9807), .A3(n9726), .A4(n11073), .ZN(n9812) );
  INV_X1 U12994 ( .A(n9970), .ZN(n9810) );
  AND2_X2 U12995 ( .A1(n11070), .A2(n11071), .ZN(n9811) );
  NAND2_X1 U12996 ( .A1(n11143), .A2(n9813), .ZN(n9904) );
  NOR2_X1 U12997 ( .A1(n11051), .A2(n9707), .ZN(n9813) );
  NAND2_X1 U12998 ( .A1(n10035), .A2(n9646), .ZN(n11051) );
  NAND2_X2 U12999 ( .A1(n15281), .A2(n15214), .ZN(n15291) );
  NAND2_X2 U13000 ( .A1(n15302), .A2(n15213), .ZN(n15281) );
  NAND2_X1 U13001 ( .A1(n15211), .A2(n15210), .ZN(n15302) );
  CLKBUF_X1 U13002 ( .A(n11390), .Z(n9820) );
  INV_X2 U13003 ( .A(n11390), .ZN(n11392) );
  OAI21_X2 U13004 ( .B1(n9613), .B2(n13712), .A(n11584), .ZN(n11588) );
  NAND2_X1 U13005 ( .A1(n14006), .A2(n14005), .ZN(n14004) );
  AND2_X2 U13006 ( .A1(n10892), .A2(n19619), .ZN(n10848) );
  NAND4_X1 U13007 ( .A1(n10844), .A2(n10845), .A3(n10843), .A4(n10846), .ZN(
        n9847) );
  NAND4_X1 U13008 ( .A1(n10842), .A2(n10841), .A3(n10839), .A4(n10840), .ZN(
        n9849) );
  NAND2_X2 U13009 ( .A1(n9851), .A2(n9850), .ZN(n10892) );
  NAND3_X1 U13010 ( .A1(n10410), .A2(n10825), .A3(n10824), .ZN(n9850) );
  NAND3_X1 U13011 ( .A1(n9857), .A2(n9855), .A3(n9759), .ZN(n9852) );
  INV_X1 U13012 ( .A(n10299), .ZN(n9854) );
  NAND2_X1 U13013 ( .A1(n9859), .A2(n9856), .ZN(n9855) );
  INV_X1 U13014 ( .A(n9858), .ZN(n9857) );
  AOI21_X1 U13015 ( .B1(n9859), .B2(n10299), .A(n11771), .ZN(n9858) );
  INV_X1 U13016 ( .A(n9862), .ZN(n16018) );
  NAND3_X1 U13017 ( .A1(n12430), .A2(n12429), .A3(n9866), .ZN(n12512) );
  NAND2_X1 U13018 ( .A1(n10056), .A2(n9749), .ZN(n12518) );
  NOR2_X1 U13019 ( .A1(n10056), .A2(n9711), .ZN(n10054) );
  NAND4_X1 U13020 ( .A1(n12430), .A2(n9592), .A3(n12429), .A4(n12431), .ZN(
        n10053) );
  INV_X2 U13021 ( .A(n15200), .ZN(n9869) );
  OR2_X1 U13022 ( .A1(n15145), .A2(n20583), .ZN(n9871) );
  NAND3_X1 U13023 ( .A1(n12680), .A2(n12690), .A3(n12823), .ZN(n9874) );
  AND2_X2 U13024 ( .A1(n12740), .A2(n9875), .ZN(n14826) );
  NOR2_X2 U13025 ( .A1(n14812), .A2(n10389), .ZN(n14770) );
  NAND2_X2 U13026 ( .A1(n12448), .A2(n20694), .ZN(n12521) );
  NAND2_X1 U13027 ( .A1(n9926), .A2(n9878), .ZN(n9876) );
  OAI211_X1 U13028 ( .C1(n9926), .C2(n9880), .A(n9876), .B(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9886) );
  NAND2_X1 U13029 ( .A1(n9705), .A2(n11415), .ZN(n9885) );
  NAND2_X1 U13030 ( .A1(n11218), .A2(n9641), .ZN(n9888) );
  INV_X1 U13031 ( .A(n9887), .ZN(n16250) );
  INV_X1 U13032 ( .A(n11234), .ZN(n9896) );
  NAND2_X1 U13033 ( .A1(n11459), .A2(n11217), .ZN(n9897) );
  AND2_X2 U13034 ( .A1(n9900), .A2(n9899), .ZN(n10978) );
  NAND2_X1 U13035 ( .A1(n10970), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9899) );
  INV_X1 U13036 ( .A(n10959), .ZN(n9900) );
  NAND3_X1 U13037 ( .A1(n10064), .A2(n10063), .A3(n10062), .ZN(n10970) );
  NAND3_X1 U13038 ( .A1(n9904), .A2(n11144), .A3(n9905), .ZN(n11153) );
  NAND3_X1 U13039 ( .A1(n11103), .A2(n15896), .A3(n11141), .ZN(n9905) );
  NAND3_X1 U13040 ( .A1(n9904), .A2(n9905), .A3(n9720), .ZN(n9903) );
  NAND2_X1 U13041 ( .A1(n11153), .A2(n11152), .ZN(n16367) );
  INV_X1 U13042 ( .A(n12657), .ZN(n10367) );
  NOR2_X2 U13043 ( .A1(n14356), .A2(n14362), .ZN(n14360) );
  NOR2_X2 U13044 ( .A1(n11425), .A2(n11426), .ZN(n15596) );
  NAND2_X1 U13045 ( .A1(n16709), .A2(n16710), .ZN(n11072) );
  NAND4_X1 U13046 ( .A1(n10474), .A2(n10526), .A3(n10514), .A4(n10473), .ZN(
        n14355) );
  NAND2_X1 U13047 ( .A1(n14346), .A2(n14345), .ZN(n14348) );
  INV_X1 U13048 ( .A(n10906), .ZN(n13903) );
  NAND2_X1 U13049 ( .A1(n15912), .A2(n10587), .ZN(n15907) );
  NOR2_X1 U13050 ( .A1(n11436), .A2(n11435), .ZN(n11437) );
  NOR2_X1 U13051 ( .A1(n14200), .A2(n14201), .ZN(n10662) );
  NAND2_X2 U13052 ( .A1(n10760), .A2(n10759), .ZN(n11425) );
  NAND2_X2 U13053 ( .A1(n15690), .A2(n15692), .ZN(n15683) );
  NAND2_X1 U13054 ( .A1(n10942), .A2(n10941), .ZN(n10036) );
  NAND2_X1 U13055 ( .A1(n10036), .A2(n9718), .ZN(n9972) );
  NAND2_X2 U13056 ( .A1(n19186), .A2(n19214), .ZN(n17362) );
  OR2_X1 U13057 ( .A1(n19396), .A2(n16378), .ZN(n11194) );
  NAND2_X1 U13058 ( .A1(n9930), .A2(n9931), .ZN(n11154) );
  INV_X2 U13059 ( .A(n11195), .ZN(n11173) );
  AOI22_X1 U13060 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19773), .B1(
        n19918), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11019) );
  NAND2_X1 U13061 ( .A1(n12432), .A2(n12496), .ZN(n12667) );
  OR2_X1 U13062 ( .A1(n9717), .A2(n10374), .ZN(n10007) );
  NAND2_X1 U13063 ( .A1(n10059), .A2(n14542), .ZN(n10058) );
  XNOR2_X1 U13064 ( .A(n10058), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14586) );
  NOR2_X2 U13065 ( .A1(n16595), .A2(n11551), .ZN(n16549) );
  NAND2_X1 U13066 ( .A1(n10043), .A2(n10040), .ZN(P2_U3027) );
  AOI211_X2 U13067 ( .C1(n16518), .C2(n10920), .A(n17216), .B(n10919), .ZN(
        n17212) );
  OAI211_X1 U13068 ( .C1(n11531), .C2(n19590), .A(n11532), .B(n11533), .ZN(
        P2_U2986) );
  NAND2_X2 U13069 ( .A1(n14689), .A2(n14690), .ZN(n14675) );
  NAND2_X1 U13070 ( .A1(n13904), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n9908) );
  AND2_X1 U13071 ( .A1(n10902), .A2(n9909), .ZN(n13905) );
  AND2_X1 U13072 ( .A1(n10889), .A2(n9909), .ZN(n10399) );
  NAND2_X1 U13073 ( .A1(n10906), .A2(n9909), .ZN(n10493) );
  NAND3_X1 U13074 ( .A1(n10894), .A2(n10893), .A3(n9909), .ZN(n10900) );
  NAND2_X1 U13075 ( .A1(n10859), .A2(n9909), .ZN(n10860) );
  AND2_X1 U13076 ( .A1(n19429), .A2(n9909), .ZN(n19426) );
  AND2_X1 U13077 ( .A1(n19644), .A2(n9909), .ZN(n20178) );
  INV_X1 U13078 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9910) );
  NAND2_X2 U13079 ( .A1(n9914), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18652) );
  INV_X1 U13080 ( .A(n9915), .ZN(n16890) );
  NAND2_X1 U13081 ( .A1(n9915), .A2(n12210), .ZN(n9918) );
  INV_X1 U13082 ( .A(n9918), .ZN(n12035) );
  NAND2_X4 U13083 ( .A1(n9920), .A2(n10954), .ZN(n11390) );
  NAND2_X1 U13084 ( .A1(n9989), .A2(n17077), .ZN(n9988) );
  NAND2_X1 U13085 ( .A1(n9923), .A2(n12027), .ZN(n17079) );
  AND2_X2 U13086 ( .A1(n11475), .A2(n9656), .ZN(n11418) );
  INV_X1 U13087 ( .A(n10225), .ZN(n9931) );
  NAND2_X1 U13088 ( .A1(n9930), .A2(n9929), .ZN(n11260) );
  INV_X1 U13089 ( .A(n11110), .ZN(n9933) );
  NAND2_X1 U13090 ( .A1(n11258), .A2(n9939), .ZN(n11259) );
  AND2_X1 U13091 ( .A1(n11287), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n9939) );
  NAND2_X1 U13092 ( .A1(n11246), .A2(n16010), .ZN(n11258) );
  NAND2_X1 U13093 ( .A1(n9940), .A2(n9569), .ZN(n9941) );
  INV_X1 U13094 ( .A(n15202), .ZN(n9940) );
  NAND3_X1 U13095 ( .A1(n9944), .A2(n9945), .A3(n9943), .ZN(n9942) );
  NAND2_X1 U13096 ( .A1(n13205), .A2(n15212), .ZN(n9944) );
  NAND2_X1 U13097 ( .A1(n15211), .A2(n13205), .ZN(n9945) );
  NAND2_X1 U13098 ( .A1(n9946), .A2(n13181), .ZN(n14484) );
  NAND2_X1 U13099 ( .A1(n14456), .A2(n13180), .ZN(n9946) );
  OAI211_X2 U13100 ( .C1(n14456), .C2(n9949), .A(n9947), .B(n14483), .ZN(
        n10384) );
  INV_X1 U13101 ( .A(n13180), .ZN(n9948) );
  INV_X1 U13102 ( .A(n13181), .ZN(n9949) );
  NAND2_X2 U13103 ( .A1(n17165), .A2(n13169), .ZN(n14456) );
  AND2_X2 U13104 ( .A1(n12667), .A2(n12665), .ZN(n12448) );
  AOI21_X2 U13105 ( .B1(n12513), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12515), .ZN(n12520) );
  INV_X1 U13106 ( .A(n10057), .ZN(n20513) );
  NAND2_X1 U13107 ( .A1(n10139), .A2(n13139), .ZN(n10057) );
  XNOR2_X1 U13108 ( .A(n12690), .B(n10369), .ZN(n13135) );
  AND2_X4 U13109 ( .A1(n16786), .A2(n10783), .ZN(n11697) );
  AND2_X4 U13110 ( .A1(n10449), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11694) );
  INV_X1 U13111 ( .A(n18029), .ZN(n18032) );
  NAND2_X2 U13112 ( .A1(n12069), .A2(n9638), .ZN(n18775) );
  NAND2_X1 U13113 ( .A1(n11663), .A2(n9966), .ZN(n9965) );
  INV_X1 U13114 ( .A(n16019), .ZN(n9966) );
  NAND3_X1 U13115 ( .A1(n9628), .A2(P3_EAX_REG_22__SCAN_IN), .A3(
        P3_EAX_REG_21__SCAN_IN), .ZN(n9967) );
  AND2_X4 U13116 ( .A1(n10446), .A2(n16834), .ZN(n11728) );
  AND2_X2 U13117 ( .A1(n9969), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10446) );
  NAND2_X1 U13118 ( .A1(n11072), .A2(n11068), .ZN(n9970) );
  NAND2_X1 U13119 ( .A1(n10863), .A2(n10901), .ZN(n10894) );
  NAND2_X1 U13120 ( .A1(n11012), .A2(n11015), .ZN(n20039) );
  NOR2_X1 U13121 ( .A1(n9613), .A2(n11567), .ZN(n11012) );
  NOR2_X2 U13122 ( .A1(n16235), .A2(n16468), .ZN(n16230) );
  AND2_X4 U13123 ( .A1(n10832), .A2(n10783), .ZN(n11700) );
  AND2_X2 U13124 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10832) );
  NOR2_X1 U13125 ( .A1(n15952), .A2(n11567), .ZN(n11014) );
  OR2_X1 U13126 ( .A1(n16436), .A2(n19574), .ZN(n9976) );
  NAND3_X1 U13127 ( .A1(n10848), .A2(n9668), .A3(n10849), .ZN(n10880) );
  NAND2_X2 U13128 ( .A1(n18345), .A2(n18357), .ZN(n18298) );
  NAND3_X1 U13129 ( .A1(n12016), .A2(n12015), .A3(n10097), .ZN(n18345) );
  NAND2_X1 U13130 ( .A1(n9978), .A2(n9982), .ZN(P3_U2799) );
  NAND3_X1 U13131 ( .A1(n9983), .A2(n18428), .A3(n9979), .ZN(n9978) );
  AOI21_X1 U13132 ( .B1(n16891), .B2(n12035), .A(n12034), .ZN(n9984) );
  OAI21_X2 U13133 ( .B1(n9989), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n9985), .ZN(n17053) );
  INV_X1 U13134 ( .A(n17079), .ZN(n9986) );
  AND2_X1 U13135 ( .A1(n12028), .A2(n17070), .ZN(n9987) );
  NAND2_X1 U13136 ( .A1(n18258), .A2(n18365), .ZN(n18263) );
  NAND2_X1 U13137 ( .A1(n18437), .A2(n18357), .ZN(n9992) );
  NAND2_X1 U13138 ( .A1(n12233), .A2(n12234), .ZN(n9997) );
  NAND2_X1 U13139 ( .A1(n14120), .A2(n9996), .ZN(n9994) );
  XNOR2_X1 U13140 ( .A(n12237), .B(n12238), .ZN(n13979) );
  NOR2_X2 U13141 ( .A1(n18609), .A2(n17027), .ZN(n17044) );
  NAND2_X2 U13142 ( .A1(n18656), .A2(n18568), .ZN(n18609) );
  NAND2_X1 U13143 ( .A1(n14959), .A2(n9632), .ZN(n10004) );
  NAND2_X1 U13144 ( .A1(n10374), .A2(n10011), .ZN(n10009) );
  INV_X1 U13145 ( .A(n13234), .ZN(n13223) );
  NAND2_X1 U13146 ( .A1(n9643), .A2(n10014), .ZN(n15421) );
  AND2_X2 U13147 ( .A1(n10021), .A2(n13270), .ZN(n17115) );
  NAND4_X1 U13148 ( .A1(n13266), .A2(n13264), .A3(n13265), .A4(n13267), .ZN(
        n10021) );
  NAND3_X1 U13149 ( .A1(n15320), .A2(n14576), .A3(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14577) );
  INV_X1 U13150 ( .A(n10026), .ZN(n10985) );
  NAND2_X1 U13151 ( .A1(n10026), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10064) );
  NAND2_X1 U13152 ( .A1(n10034), .A2(n10948), .ZN(n10026) );
  NOR2_X2 U13153 ( .A1(n11022), .A2(n11016), .ZN(n19773) );
  NAND3_X2 U13154 ( .A1(n10106), .A2(n10105), .A3(n9686), .ZN(n10035) );
  NAND3_X1 U13155 ( .A1(n10035), .A2(n10066), .A3(n10028), .ZN(n11075) );
  NAND4_X1 U13156 ( .A1(n10435), .A2(n10434), .A3(n10436), .A4(n10433), .ZN(
        n10031) );
  NAND2_X1 U13157 ( .A1(n10030), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10033) );
  NAND4_X1 U13158 ( .A1(n10440), .A2(n10438), .A3(n10437), .A4(n10439), .ZN(
        n10030) );
  NAND3_X1 U13159 ( .A1(n16709), .A2(n16710), .A3(n11065), .ZN(n11071) );
  NAND2_X1 U13160 ( .A1(n10856), .A2(n10943), .ZN(n10948) );
  NAND3_X1 U13161 ( .A1(n10034), .A2(n10948), .A3(n13485), .ZN(n11406) );
  NAND2_X1 U13162 ( .A1(n10035), .A2(n10104), .ZN(n11032) );
  NAND2_X1 U13163 ( .A1(n10035), .A2(n10332), .ZN(n11103) );
  NAND2_X1 U13164 ( .A1(n10036), .A2(n10943), .ZN(n10961) );
  NAND2_X1 U13165 ( .A1(n10044), .A2(n13881), .ZN(n10047) );
  NAND2_X1 U13166 ( .A1(n10046), .A2(n10135), .ZN(n10045) );
  INV_X1 U13167 ( .A(n12522), .ZN(n10046) );
  NAND2_X1 U13168 ( .A1(n10049), .A2(n10135), .ZN(n10048) );
  INV_X1 U13169 ( .A(n13881), .ZN(n10049) );
  NAND2_X2 U13170 ( .A1(n10052), .A2(n10055), .ZN(n20694) );
  NAND3_X1 U13171 ( .A1(n10141), .A2(n10140), .A3(n14541), .ZN(n10059) );
  NAND4_X1 U13172 ( .A1(n9642), .A2(n10946), .A3(n10895), .A4(n10061), .ZN(
        n10062) );
  NAND3_X1 U13173 ( .A1(n16864), .A2(n10952), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n10063) );
  NAND2_X1 U13174 ( .A1(n19773), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n10068) );
  NAND2_X1 U13175 ( .A1(n19880), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n10069) );
  NAND2_X1 U13176 ( .A1(n16314), .A2(n10074), .ZN(n10072) );
  AND2_X4 U13177 ( .A1(n10082), .A2(n13949), .ZN(n12353) );
  NAND2_X2 U13178 ( .A1(n12517), .A2(n12516), .ZN(n13881) );
  NAND3_X1 U13179 ( .A1(n13213), .A2(n10085), .A3(n13212), .ZN(n10084) );
  NAND2_X1 U13180 ( .A1(n13182), .A2(n13858), .ZN(n13190) );
  AND3_X2 U13181 ( .A1(n12559), .A2(n10369), .A3(n12679), .ZN(n12611) );
  NAND2_X4 U13182 ( .A1(n10090), .A2(n10089), .ZN(n13934) );
  NAND2_X2 U13183 ( .A1(n9586), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18343) );
  AND2_X2 U13184 ( .A1(n12021), .A2(n18298), .ZN(n16929) );
  INV_X1 U13185 ( .A(n10984), .ZN(n10099) );
  INV_X1 U13186 ( .A(n10977), .ZN(n10102) );
  NAND2_X1 U13187 ( .A1(n10277), .A2(n11005), .ZN(n10103) );
  NAND2_X1 U13188 ( .A1(n16394), .A2(n10351), .ZN(n10346) );
  NOR2_X2 U13189 ( .A1(n16351), .A2(n10107), .ZN(n16295) );
  NAND2_X1 U13190 ( .A1(n13479), .A2(n9761), .ZN(n12259) );
  INV_X1 U13191 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10111) );
  INV_X1 U13192 ( .A(n10120), .ZN(n11864) );
  NAND3_X1 U13193 ( .A1(n10125), .A2(n10124), .A3(n9910), .ZN(n10344) );
  AND3_X4 U13194 ( .A1(n10783), .A2(n16834), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11699) );
  AND2_X4 U13195 ( .A1(n10447), .A2(n16834), .ZN(n11698) );
  AND2_X2 U13196 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10447) );
  NAND2_X1 U13197 ( .A1(n10128), .A2(n10126), .ZN(n11218) );
  AND2_X2 U13198 ( .A1(n10142), .A2(n14540), .ZN(n15102) );
  INV_X1 U13199 ( .A(n13208), .ZN(n10143) );
  NAND3_X1 U13200 ( .A1(n9709), .A2(n14429), .A3(n10145), .ZN(n10144) );
  NAND3_X1 U13201 ( .A1(n12680), .A2(n12690), .A3(n13858), .ZN(n10146) );
  NAND2_X1 U13202 ( .A1(n10146), .A2(n13144), .ZN(n14430) );
  CLKBUF_X1 U13203 ( .A(n12353), .Z(n10147) );
  NAND4_X1 U13204 ( .A1(n10182), .A2(n15939), .A3(n15941), .A4(n19581), .ZN(
        n15914) );
  NAND2_X1 U13205 ( .A1(n15846), .A2(n10183), .ZN(n13577) );
  NAND2_X1 U13206 ( .A1(n13459), .A2(n9725), .ZN(n15741) );
  INV_X1 U13207 ( .A(n10193), .ZN(n15750) );
  NOR2_X2 U13208 ( .A1(n17431), .A2(n17695), .ZN(n17423) );
  NOR2_X1 U13209 ( .A1(n17432), .A2(n17433), .ZN(n17431) );
  NOR2_X2 U13210 ( .A1(n17382), .A2(n17695), .ZN(n17473) );
  NAND3_X1 U13211 ( .A1(n16941), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n12026), .ZN(n18258) );
  NAND2_X1 U13212 ( .A1(n17695), .A2(n10201), .ZN(n10200) );
  INV_X1 U13213 ( .A(n10206), .ZN(n17493) );
  AOI21_X1 U13214 ( .B1(n10208), .B2(n19228), .A(n10207), .ZN(n17406) );
  INV_X1 U13215 ( .A(n17409), .ZN(n10211) );
  INV_X1 U13216 ( .A(n10213), .ZN(n13596) );
  NOR2_X2 U13217 ( .A1(n16907), .A2(n13600), .ZN(n16877) );
  OAI21_X1 U13218 ( .B1(n12117), .B2(n12053), .A(n10219), .ZN(n11905) );
  NAND3_X1 U13219 ( .A1(n12267), .A2(n12266), .A3(n12268), .ZN(P2_U2983) );
  NAND2_X1 U13220 ( .A1(n11450), .A2(n11449), .ZN(n11486) );
  NAND2_X1 U13221 ( .A1(n11450), .A2(n10221), .ZN(n10220) );
  INV_X1 U13222 ( .A(n11449), .ZN(n10222) );
  NAND2_X1 U13223 ( .A1(n14601), .A2(n10224), .ZN(n11488) );
  NOR2_X1 U13224 ( .A1(n16378), .A2(n11484), .ZN(n10224) );
  AND2_X1 U13225 ( .A1(n11173), .A2(n10232), .ZN(n11181) );
  NAND2_X1 U13226 ( .A1(n11173), .A2(n10408), .ZN(n11190) );
  NAND2_X1 U13227 ( .A1(n11173), .A2(n10230), .ZN(n11192) );
  XNOR2_X2 U13228 ( .A(n14661), .B(n14660), .ZN(n15323) );
  NAND2_X1 U13229 ( .A1(n10241), .A2(n10239), .ZN(n14830) );
  NAND2_X1 U13230 ( .A1(n13892), .A2(n10254), .ZN(n13940) );
  INV_X1 U13231 ( .A(n13940), .ZN(n10646) );
  NOR2_X2 U13232 ( .A1(n15683), .A2(n9743), .ZN(n15634) );
  NOR2_X2 U13233 ( .A1(n13587), .A2(n9744), .ZN(n15778) );
  NOR2_X2 U13234 ( .A1(n15760), .A2(n10263), .ZN(n15708) );
  NAND2_X1 U13235 ( .A1(n10427), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10266) );
  INV_X1 U13236 ( .A(n11425), .ZN(n10269) );
  NOR2_X1 U13237 ( .A1(n11425), .A2(n10275), .ZN(n15598) );
  XNOR2_X2 U13238 ( .A(n10278), .B(n10999), .ZN(n11567) );
  NAND2_X2 U13239 ( .A1(n10321), .A2(n10993), .ZN(n10278) );
  NAND2_X2 U13240 ( .A1(n10282), .A2(n10279), .ZN(n20311) );
  NAND3_X1 U13241 ( .A1(n10774), .A2(n10776), .A3(n10775), .ZN(n10281) );
  NAND3_X1 U13242 ( .A1(n10772), .A2(n10770), .A3(n10771), .ZN(n10283) );
  NAND2_X1 U13243 ( .A1(n15987), .A2(n15986), .ZN(n15985) );
  INV_X1 U13244 ( .A(n11796), .ZN(n10285) );
  NAND2_X1 U13245 ( .A1(n15976), .A2(n15975), .ZN(n15977) );
  INV_X1 U13246 ( .A(n11856), .ZN(n10292) );
  INV_X1 U13247 ( .A(n16040), .ZN(n10296) );
  NAND2_X1 U13248 ( .A1(n11717), .A2(n10303), .ZN(n10300) );
  OR2_X2 U13249 ( .A1(n16012), .A2(n10302), .ZN(n10299) );
  INV_X1 U13250 ( .A(n10304), .ZN(n16013) );
  INV_X1 U13251 ( .A(n14422), .ZN(n10309) );
  NAND2_X1 U13252 ( .A1(n10309), .A2(n10310), .ZN(n11543) );
  NAND2_X1 U13253 ( .A1(n15632), .A2(n9735), .ZN(n10319) );
  NAND2_X1 U13254 ( .A1(n15632), .A2(n15633), .ZN(n15621) );
  NAND3_X1 U13255 ( .A1(n10321), .A2(n10993), .A3(n10320), .ZN(n16732) );
  NAND2_X1 U13256 ( .A1(n11468), .A2(n10322), .ZN(n15676) );
  NAND2_X1 U13257 ( .A1(n10326), .A2(n10325), .ZN(n15810) );
  NAND3_X1 U13258 ( .A1(n9633), .A2(n11459), .A3(n16331), .ZN(n10330) );
  NAND3_X1 U13259 ( .A1(n9633), .A2(n11459), .A3(n9724), .ZN(n10327) );
  NAND2_X1 U13260 ( .A1(n11153), .A2(n10335), .ZN(n10334) );
  NAND2_X1 U13261 ( .A1(n10334), .A2(n10336), .ZN(n11170) );
  NAND3_X1 U13262 ( .A1(n10343), .A2(n10342), .A3(n10811), .ZN(n10341) );
  NOR2_X2 U13263 ( .A1(n11022), .A2(n11025), .ZN(n19846) );
  AND2_X1 U13264 ( .A1(n11474), .A2(n10353), .ZN(n16281) );
  NAND2_X1 U13265 ( .A1(n11474), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16309) );
  AND4_X2 U13266 ( .A1(n10355), .A2(n10356), .A3(n10357), .A4(n10946), .ZN(
        n10994) );
  NAND2_X1 U13267 ( .A1(n11418), .A2(n9766), .ZN(n10359) );
  OAI211_X1 U13268 ( .C1(n11418), .C2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n10360), .B(n10359), .ZN(n12265) );
  NAND2_X1 U13269 ( .A1(n14536), .A2(n9644), .ZN(n10379) );
  NAND3_X1 U13270 ( .A1(n10382), .A2(n14539), .A3(n10381), .ZN(n10380) );
  NOR2_X2 U13271 ( .A1(n14749), .A2(n10385), .ZN(n14705) );
  INV_X1 U13272 ( .A(n14923), .ZN(n12740) );
  NAND4_X1 U13273 ( .A1(n14460), .A2(n12719), .A3(n14437), .A4(n12701), .ZN(
        n14923) );
  NAND3_X1 U13274 ( .A1(n14460), .A2(n12701), .A3(n9594), .ZN(n14461) );
  NOR2_X1 U13275 ( .A1(n14675), .A2(n14677), .ZN(n13126) );
  CLKBUF_X1 U13276 ( .A(n14503), .Z(n15539) );
  NAND2_X1 U13277 ( .A1(n13179), .A2(n13178), .ZN(n13180) );
  AND3_X1 U13278 ( .A1(n12426), .A2(n12401), .A3(n12407), .ZN(n12398) );
  INV_X1 U13279 ( .A(n12401), .ZN(n12416) );
  OR2_X1 U13280 ( .A1(n13110), .A2(n12309), .ZN(n12311) );
  INV_X1 U13281 ( .A(n11253), .ZN(n11261) );
  CLKBUF_X1 U13282 ( .A(n14422), .Z(n16050) );
  INV_X1 U13283 ( .A(n15617), .ZN(n10760) );
  NAND2_X1 U13284 ( .A1(n15634), .A2(n15635), .ZN(n15617) );
  NAND2_X1 U13285 ( .A1(n14214), .A2(n10985), .ZN(n10986) );
  NAND2_X1 U13286 ( .A1(n11235), .A2(n11236), .ZN(n11245) );
  CLKBUF_X1 U13287 ( .A(n13940), .Z(n15857) );
  CLKBUF_X1 U13288 ( .A(n15774), .Z(n15782) );
  NAND2_X1 U13289 ( .A1(n16283), .A2(n16282), .ZN(n11537) );
  CLKBUF_X1 U13290 ( .A(n15683), .Z(n15694) );
  OR2_X1 U13291 ( .A1(n16544), .A2(n19590), .ZN(n10421) );
  CLKBUF_X1 U13292 ( .A(n13587), .Z(n14283) );
  INV_X1 U13293 ( .A(n11006), .ZN(n15952) );
  CLKBUF_X1 U13294 ( .A(n14199), .Z(n15828) );
  XNOR2_X1 U13295 ( .A(n9657), .B(n14546), .ZN(n15331) );
  NAND2_X1 U13296 ( .A1(n10912), .A2(n10903), .ZN(n10904) );
  NAND2_X1 U13297 ( .A1(n14355), .A2(n14354), .ZN(n10497) );
  OR2_X1 U13298 ( .A1(n11003), .A2(n11002), .ZN(n11004) );
  NAND2_X1 U13299 ( .A1(n11253), .A2(n11252), .ZN(n11265) );
  NAND2_X1 U13300 ( .A1(n11479), .A2(n11447), .ZN(n15599) );
  OAI21_X1 U13301 ( .B1(n14634), .B2(n17203), .A(n10938), .ZN(n10939) );
  AOI22_X1 U13302 ( .A1(n12368), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12585), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12387) );
  NAND2_X1 U13303 ( .A1(n20840), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13221) );
  OR2_X1 U13304 ( .A1(n14600), .A2(n19573), .ZN(n12268) );
  OR2_X1 U13305 ( .A1(n14600), .A2(n17227), .ZN(n11410) );
  AOI21_X1 U13306 ( .B1(n14588), .B2(n20518), .A(n14584), .ZN(n14585) );
  NAND2_X1 U13307 ( .A1(n15572), .A2(n20585), .ZN(n20807) );
  INV_X1 U13308 ( .A(n12420), .ZN(n13860) );
  INV_X1 U13309 ( .A(n11297), .ZN(n11395) );
  AND4_X1 U13310 ( .A1(n10609), .A2(n10608), .A3(n10607), .A4(n10606), .ZN(
        n10398) );
  NOR2_X2 U13311 ( .A1(n19566), .A2(n19538), .ZN(n10400) );
  AND2_X1 U13312 ( .A1(n19445), .A2(n13904), .ZN(n19477) );
  NOR2_X1 U13313 ( .A1(n14750), .A2(n14760), .ZN(n10401) );
  OR2_X1 U13314 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n13524) );
  AND3_X1 U13315 ( .A1(n10452), .A2(n10451), .A3(n10450), .ZN(n10402) );
  AND2_X1 U13316 ( .A1(n14215), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n10403) );
  INV_X1 U13317 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n10833) );
  AND2_X2 U13318 ( .A1(n14583), .A2(n13426), .ZN(n10405) );
  AND4_X1 U13319 ( .A1(n16290), .A2(n11210), .A3(n11463), .A4(n16312), .ZN(
        n10406) );
  NAND2_X2 U13320 ( .A1(n15098), .A2(n14014), .ZN(n15101) );
  INV_X1 U13321 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n13636) );
  OR2_X1 U13322 ( .A1(n14977), .A2(n20432), .ZN(n10407) );
  NAND2_X1 U13323 ( .A1(n11424), .A2(n11423), .ZN(n11525) );
  OR2_X1 U13324 ( .A1(n9571), .A2(n11172), .ZN(n10408) );
  OR2_X1 U13325 ( .A1(n9571), .A2(n11178), .ZN(n10409) );
  INV_X1 U13326 ( .A(n21198), .ZN(n21214) );
  AND3_X1 U13327 ( .A1(n10823), .A2(n10822), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10410) );
  INV_X1 U13328 ( .A(n11105), .ZN(n11097) );
  AND4_X1 U13329 ( .A1(n11948), .A2(n11947), .A3(n11946), .A4(n11945), .ZN(
        n10411) );
  INV_X1 U13330 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n11252) );
  INV_X1 U13331 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12172) );
  INV_X1 U13332 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12028) );
  INV_X2 U13333 ( .A(n18166), .ZN(n18169) );
  NAND3_X2 U13334 ( .A1(n12330), .A2(n12329), .A3(n12328), .ZN(n12414) );
  INV_X1 U13335 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11484) );
  NOR2_X1 U13336 ( .A1(n20958), .A2(n20929), .ZN(n10412) );
  NOR2_X1 U13337 ( .A1(n20958), .A2(n20693), .ZN(n10413) );
  OR2_X1 U13338 ( .A1(n18357), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10415) );
  AND4_X1 U13339 ( .A1(n10445), .A2(n10444), .A3(n10443), .A4(n10442), .ZN(
        n10416) );
  NOR2_X1 U13340 ( .A1(n20958), .A2(n21068), .ZN(n10418) );
  NOR2_X1 U13341 ( .A1(n20958), .A2(n20778), .ZN(n10419) );
  INV_X1 U13342 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12649) );
  NOR2_X1 U13343 ( .A1(n18313), .A2(n18478), .ZN(n16990) );
  NAND2_X1 U13344 ( .A1(n20611), .A2(n14486), .ZN(n13323) );
  NOR2_X1 U13345 ( .A1(n11642), .A2(n11641), .ZN(n10420) );
  AND2_X1 U13346 ( .A1(n20447), .A2(n12408), .ZN(n20440) );
  INV_X2 U13347 ( .A(n20440), .ZN(n15011) );
  NAND2_X1 U13348 ( .A1(n20447), .A2(n20626), .ZN(n15013) );
  INV_X1 U13349 ( .A(n20505), .ZN(n14381) );
  AND2_X1 U13350 ( .A1(n13779), .A2(n13778), .ZN(n19808) );
  INV_X1 U13351 ( .A(n19590), .ZN(n19577) );
  INV_X1 U13352 ( .A(n19718), .ZN(n19763) );
  OR2_X1 U13353 ( .A1(n19840), .A2(n20271), .ZN(n19718) );
  INV_X1 U13354 ( .A(n19726), .ZN(n19733) );
  INV_X1 U13355 ( .A(n10516), .ZN(n10688) );
  NAND2_X2 U13356 ( .A1(n12296), .A2(n12295), .ZN(n12417) );
  AND2_X1 U13357 ( .A1(n12281), .A2(n12280), .ZN(n10422) );
  NAND2_X1 U13358 ( .A1(n12403), .A2(n12417), .ZN(n12404) );
  NAND2_X1 U13359 ( .A1(n12406), .A2(n20622), .ZN(n12418) );
  INV_X1 U13360 ( .A(n13239), .ZN(n13220) );
  INV_X1 U13361 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12269) );
  OR2_X1 U13362 ( .A1(n12582), .A2(n12581), .ZN(n13173) );
  INV_X1 U13363 ( .A(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12388) );
  AND2_X1 U13364 ( .A1(n21134), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12510) );
  AND2_X1 U13365 ( .A1(n13713), .A2(n11716), .ZN(n10952) );
  NAND2_X1 U13366 ( .A1(n13220), .A2(n13219), .ZN(n13240) );
  NAND2_X1 U13367 ( .A1(n12414), .A2(n12416), .ZN(n12415) );
  INV_X1 U13368 ( .A(n9604), .ZN(n12484) );
  AOI22_X1 U13369 ( .A1(n12451), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12324), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12283) );
  NAND2_X1 U13370 ( .A1(n11088), .A2(n10867), .ZN(n10868) );
  NAND2_X1 U13371 ( .A1(n19624), .A2(n10906), .ZN(n10893) );
  AOI22_X1 U13372 ( .A1(n11728), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10821), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10431) );
  AOI22_X1 U13373 ( .A1(n12368), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12358), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12321) );
  INV_X1 U13374 ( .A(n14813), .ZN(n12879) );
  INV_X1 U13375 ( .A(n12854), .ZN(n12855) );
  INV_X1 U13376 ( .A(n14926), .ZN(n12739) );
  OR2_X1 U13377 ( .A1(n12595), .A2(n12594), .ZN(n13184) );
  AND2_X1 U13378 ( .A1(n12411), .A2(n12417), .ZN(n13538) );
  INV_X1 U13379 ( .A(n12448), .ZN(n12449) );
  OR2_X1 U13380 ( .A1(n11691), .A2(n11690), .ZN(n11719) );
  INV_X1 U13381 ( .A(n16023), .ZN(n11663) );
  AOI22_X1 U13382 ( .A1(n10517), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n10479), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10480) );
  NAND2_X1 U13383 ( .A1(n11180), .A2(n11293), .ZN(n11230) );
  INV_X1 U13384 ( .A(n20626), .ZN(n12601) );
  INV_X1 U13385 ( .A(n15540), .ZN(n13346) );
  OAI22_X1 U13386 ( .A1(n9605), .A2(n12350), .B1(n12349), .B2(n12348), .ZN(
        n12351) );
  INV_X1 U13387 ( .A(n12897), .ZN(n12898) );
  INV_X1 U13388 ( .A(n12668), .ZN(n13526) );
  NAND2_X1 U13389 ( .A1(n13310), .A2(n13323), .ZN(n13350) );
  NAND2_X1 U13390 ( .A1(n12411), .A2(n12407), .ZN(n12420) );
  INV_X1 U13391 ( .A(n13858), .ZN(n13258) );
  INV_X1 U13392 ( .A(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n21286) );
  XNOR2_X1 U13393 ( .A(n12505), .B(n12506), .ZN(n12657) );
  INV_X1 U13394 ( .A(n15826), .ZN(n11327) );
  OR2_X1 U13395 ( .A1(n11775), .A2(n10635), .ZN(n11579) );
  OR2_X1 U13396 ( .A1(n11793), .A2(n11797), .ZN(n11829) );
  INV_X1 U13397 ( .A(n15685), .ZN(n10750) );
  AND2_X1 U13398 ( .A1(n14241), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n11570) );
  INV_X1 U13399 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15737) );
  OR2_X1 U13400 ( .A1(n10492), .A2(n10491), .ZN(n11033) );
  AND2_X1 U13401 ( .A1(n11140), .A2(n16384), .ZN(n11144) );
  AND2_X1 U13402 ( .A1(n10605), .A2(n10604), .ZN(n10610) );
  INV_X1 U13403 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11066) );
  INV_X1 U13404 ( .A(n10827), .ZN(n10872) );
  AND2_X1 U13405 ( .A1(n10785), .A2(n10784), .ZN(n11117) );
  AND2_X1 U13406 ( .A1(n18357), .A2(n18577), .ZN(n18330) );
  NOR2_X1 U13407 ( .A1(n18117), .A2(n12232), .ZN(n12221) );
  AND4_X1 U13408 ( .A1(n12362), .A2(n12361), .A3(n12360), .A4(n12359), .ZN(
        n12363) );
  OR2_X1 U13409 ( .A1(n15169), .A2(n13524), .ZN(n12964) );
  NAND2_X1 U13410 ( .A1(n12856), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12897) );
  INV_X1 U13411 ( .A(n12627), .ZN(n13532) );
  INV_X1 U13412 ( .A(n14571), .ZN(n13209) );
  AND2_X1 U13413 ( .A1(n13374), .A2(n13373), .ZN(n14814) );
  INV_X1 U13414 ( .A(n15306), .ZN(n13198) );
  AND2_X1 U13415 ( .A1(n13271), .A2(n13272), .ZN(n13876) );
  INV_X1 U13416 ( .A(n14297), .ZN(n13330) );
  INV_X1 U13417 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20589) );
  INV_X1 U13418 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20840) );
  AND2_X1 U13419 ( .A1(n20958), .A2(n21065), .ZN(n20897) );
  AOI21_X1 U13420 ( .B1(n15957), .B2(n14606), .A(n14605), .ZN(n14607) );
  INV_X1 U13421 ( .A(n15761), .ZN(n10739) );
  INV_X1 U13422 ( .A(n15856), .ZN(n10645) );
  INV_X1 U13423 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16083) );
  INV_X1 U13424 ( .A(n13588), .ZN(n10702) );
  NAND2_X1 U13425 ( .A1(n11241), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11242) );
  AND3_X1 U13426 ( .A1(n11216), .A2(n10406), .A3(n11215), .ZN(n11217) );
  INV_X1 U13427 ( .A(n15812), .ZN(n11331) );
  AND2_X1 U13428 ( .A1(n11293), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11146) );
  INV_X1 U13429 ( .A(n10482), .ZN(n14220) );
  NAND2_X1 U13430 ( .A1(n17239), .A2(n13438), .ZN(n13779) );
  AND2_X1 U13431 ( .A1(n18273), .A2(n17728), .ZN(n13602) );
  INV_X1 U13432 ( .A(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13847) );
  AND2_X1 U13433 ( .A1(n18331), .A2(n12024), .ZN(n16941) );
  NOR2_X1 U13434 ( .A1(n12236), .A2(n18462), .ZN(n12237) );
  AND4_X1 U13435 ( .A1(n12140), .A2(n12139), .A3(n12138), .A4(n12137), .ZN(
        n12141) );
  INV_X1 U13436 ( .A(n19243), .ZN(n19334) );
  OR2_X1 U13437 ( .A1(n14682), .A2(n13431), .ZN(n14667) );
  INV_X1 U13438 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12628) );
  NAND2_X1 U13439 ( .A1(n20410), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14939) );
  AND2_X1 U13440 ( .A1(n13376), .A2(n13375), .ZN(n14807) );
  INV_X1 U13441 ( .A(n13395), .ZN(n13408) );
  AOI22_X1 U13442 ( .A1(n14523), .A2(n13531), .B1(n13125), .B2(n13124), .ZN(
        n13127) );
  OR2_X1 U13443 ( .A1(n14016), .A2(n20582), .ZN(n15080) );
  AOI21_X1 U13444 ( .B1(n13135), .B2(n12823), .A(n12700), .ZN(n14335) );
  NAND2_X1 U13445 ( .A1(n14925), .A2(n14874), .ZN(n14875) );
  AND3_X1 U13446 ( .A1(n12718), .A2(n12717), .A3(n12716), .ZN(n15002) );
  INV_X1 U13447 ( .A(n14552), .ZN(n14553) );
  AND2_X1 U13448 ( .A1(n13363), .A2(n13362), .ZN(n14862) );
  AND2_X1 U13449 ( .A1(n14022), .A2(n13872), .ZN(n14648) );
  OAI21_X1 U13450 ( .B1(n21218), .B2(n17141), .A(n15566), .ZN(n20588) );
  INV_X1 U13451 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20988) );
  AND2_X1 U13452 ( .A1(n13493), .A2(n15968), .ZN(n13494) );
  AND2_X1 U13453 ( .A1(n20313), .A2(n20191), .ZN(n14228) );
  INV_X1 U13454 ( .A(n15968), .ZN(n19405) );
  AND3_X1 U13455 ( .A1(n10629), .A2(n10628), .A3(n10627), .ZN(n13943) );
  AOI21_X1 U13456 ( .B1(n15600), .B2(n17192), .A(n11454), .ZN(n11455) );
  OR2_X1 U13457 ( .A1(n16649), .A2(n10934), .ZN(n16494) );
  NAND2_X1 U13458 ( .A1(n11076), .A2(n11146), .ZN(n11078) );
  AND3_X1 U13459 ( .A1(n10910), .A2(n10909), .A3(n10908), .ZN(n16795) );
  OR2_X1 U13460 ( .A1(n19804), .A2(n20271), .ZN(n19726) );
  OR2_X1 U13461 ( .A1(n19804), .A2(n20043), .ZN(n19794) );
  INV_X1 U13462 ( .A(n20275), .ZN(n19597) );
  OR3_X1 U13463 ( .A1(n19980), .A2(n20001), .A3(n20317), .ZN(n19984) );
  OR3_X1 U13464 ( .A1(n16822), .A2(n20029), .A3(n20317), .ZN(n16827) );
  AND2_X1 U13465 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17591), .ZN(n17572) );
  OR2_X1 U13466 ( .A1(n13614), .A2(n13612), .ZN(n17706) );
  NAND2_X1 U13467 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n13836), .ZN(n14042) );
  INV_X1 U13468 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18354) );
  NOR2_X1 U13469 ( .A1(n18567), .A2(n18601), .ZN(n18642) );
  NAND2_X1 U13470 ( .A1(n13667), .A2(n19333), .ZN(n18712) );
  NOR2_X2 U13471 ( .A1(n18593), .A2(n19335), .ZN(n19178) );
  AND4_X1 U13472 ( .A1(n12059), .A2(n12058), .A3(n12057), .A4(n12056), .ZN(
        n12060) );
  AOI21_X1 U13473 ( .B1(n18741), .B2(n19337), .A(n19209), .ZN(n18754) );
  INV_X1 U13474 ( .A(n19341), .ZN(n12207) );
  AND2_X1 U13475 ( .A1(n13432), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n13433) );
  AND2_X1 U13476 ( .A1(n20410), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20427) );
  INV_X1 U13477 ( .A(n20447), .ZN(n14996) );
  AND2_X1 U13478 ( .A1(n15098), .A2(n20626), .ZN(n13544) );
  INV_X1 U13479 ( .A(n15080), .ZN(n15072) );
  NAND2_X1 U13480 ( .A1(n13543), .A2(n14077), .ZN(n15076) );
  INV_X2 U13481 ( .A(n14379), .ZN(n20508) );
  AND2_X1 U13482 ( .A1(n13296), .A2(n13103), .ZN(n14523) );
  OR2_X1 U13483 ( .A1(n14447), .A2(n14446), .ZN(n15008) );
  INV_X1 U13484 ( .A(n20583), .ZN(n20518) );
  OR2_X1 U13485 ( .A1(n15232), .A2(n15233), .ZN(n15242) );
  AND2_X1 U13486 ( .A1(n13275), .A2(n21070), .ZN(n20526) );
  NAND2_X1 U13487 ( .A1(n10368), .A2(n20588), .ZN(n20729) );
  NOR2_X1 U13488 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n15586) );
  OAI21_X1 U13489 ( .B1(n20639), .B2(n20638), .A(n21080), .ZN(n20657) );
  INV_X1 U13490 ( .A(n20692), .ZN(n20682) );
  INV_X1 U13491 ( .A(n20723), .ZN(n20713) );
  NAND2_X1 U13492 ( .A1(n20587), .A2(n20586), .ZN(n20697) );
  INV_X1 U13493 ( .A(n20872), .ZN(n20995) );
  INV_X1 U13494 ( .A(n20837), .ZN(n20828) );
  INV_X1 U13495 ( .A(n20831), .ZN(n20862) );
  OAI21_X1 U13496 ( .B1(n20871), .B2(n20870), .A(n21080), .ZN(n20889) );
  OAI22_X1 U13497 ( .A1(n20904), .A2(n20903), .B1(n20902), .B2(n21018), .ZN(
        n20922) );
  AND2_X1 U13498 ( .A1(n20662), .A2(n20661), .ZN(n20893) );
  INV_X1 U13499 ( .A(n20934), .ZN(n20928) );
  INV_X1 U13500 ( .A(n21115), .ZN(n21049) );
  NOR2_X2 U13501 ( .A1(n20583), .A2(n20582), .ZN(n20629) );
  INV_X1 U13502 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n21137) );
  INV_X1 U13503 ( .A(n21221), .ZN(n21142) );
  INV_X1 U13504 ( .A(n21182), .ZN(n21193) );
  AND2_X1 U13505 ( .A1(n10955), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13626) );
  OR2_X1 U13506 ( .A1(n13495), .A2(n13494), .ZN(n13496) );
  AND2_X1 U13507 ( .A1(n13579), .A2(n13492), .ZN(n15968) );
  INV_X1 U13508 ( .A(n15958), .ZN(n19410) );
  INV_X1 U13509 ( .A(n16851), .ZN(n13630) );
  OR2_X1 U13510 ( .A1(n10713), .A2(n10712), .ZN(n14425) );
  OR2_X1 U13511 ( .A1(n10657), .A2(n10656), .ZN(n16069) );
  NOR2_X1 U13512 ( .A1(n14242), .A2(n14340), .ZN(n14383) );
  OR2_X1 U13513 ( .A1(n14006), .A2(n14005), .ZN(n14007) );
  INV_X1 U13514 ( .A(n16030), .ZN(n16036) );
  INV_X1 U13515 ( .A(n19472), .ZN(n19479) );
  INV_X1 U13516 ( .A(n17227), .ZN(n16745) );
  NAND2_X1 U13517 ( .A1(n19607), .A2(n19606), .ZN(n19647) );
  OAI21_X1 U13518 ( .B1(n16807), .B2(n16812), .A(n16806), .ZN(n19734) );
  OAI21_X1 U13519 ( .B1(n19776), .B2(n19775), .A(n19774), .ZN(n19800) );
  INV_X1 U13520 ( .A(n19821), .ZN(n19836) );
  NAND2_X1 U13521 ( .A1(n19882), .A2(n19881), .ZN(n19905) );
  OAI21_X1 U13522 ( .B1(n19921), .B2(n19920), .A(n19919), .ZN(n19943) );
  AND2_X1 U13523 ( .A1(n19984), .A2(n19982), .ZN(n20002) );
  NOR2_X2 U13524 ( .A1(n19910), .A2(n20271), .ZN(n20031) );
  NOR2_X2 U13525 ( .A1(n19948), .A2(n20043), .ZN(n20065) );
  NAND2_X1 U13526 ( .A1(n20081), .A2(n20080), .ZN(n20118) );
  AND2_X1 U13527 ( .A1(n20133), .A2(n16808), .ZN(n20127) );
  INV_X1 U13528 ( .A(n20100), .ZN(n20158) );
  AND2_X1 U13529 ( .A1(n20133), .A2(n19646), .ZN(n20180) );
  AND3_X1 U13530 ( .A1(n20195), .A2(n20259), .A3(n20202), .ZN(n20313) );
  INV_X1 U13531 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20208) );
  INV_X1 U13532 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n20190) );
  NOR2_X1 U13533 ( .A1(n13722), .A2(n13721), .ZN(n19184) );
  NOR2_X1 U13534 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17438), .ZN(n17421) );
  NOR2_X1 U13535 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17480), .ZN(n17462) );
  INV_X1 U13536 ( .A(n17724), .ZN(n17687) );
  NAND2_X1 U13537 ( .A1(n17519), .A2(n17510), .ZN(n17509) );
  NOR2_X1 U13538 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17557), .ZN(n17542) );
  NOR2_X1 U13539 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17603), .ZN(n17587) );
  NOR2_X1 U13540 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17652), .ZN(n17631) );
  INV_X1 U13541 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17653) );
  NOR3_X1 U13542 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17708) );
  NOR2_X2 U13543 ( .A1(n19322), .A2(n17721), .ZN(n17700) );
  NOR2_X1 U13544 ( .A1(n17927), .A2(n17926), .ZN(n17902) );
  AND2_X1 U13545 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n13835), .ZN(n13836) );
  INV_X1 U13546 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17992) );
  AND2_X1 U13547 ( .A1(n13928), .A2(n13669), .ZN(n18007) );
  NAND2_X1 U13548 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n18046), .ZN(n18041) );
  INV_X1 U13549 ( .A(n18061), .ZN(n18075) );
  INV_X1 U13550 ( .A(n18783), .ZN(n17863) );
  AND4_X1 U13551 ( .A1(n12004), .A2(n12003), .A3(n12002), .A4(n12001), .ZN(
        n12005) );
  AOI21_X1 U13552 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16990), .A(
        n16992), .ZN(n18315) );
  AND2_X1 U13553 ( .A1(n18526), .A2(n18538), .ZN(n18522) );
  OR2_X1 U13554 ( .A1(n16983), .A2(n16985), .ZN(n18272) );
  AND2_X1 U13555 ( .A1(n18473), .A2(n16880), .ZN(n18405) );
  INV_X1 U13556 ( .A(n18524), .ZN(n18653) );
  NOR2_X1 U13557 ( .A1(n18532), .A2(n18616), .ZN(n18560) );
  NOR2_X1 U13558 ( .A1(n18642), .A2(n18616), .ZN(n18677) );
  INV_X1 U13559 ( .A(n18713), .ZN(n18576) );
  INV_X1 U13560 ( .A(n19087), .ZN(n18856) );
  NOR2_X1 U13561 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19350) );
  INV_X1 U13562 ( .A(n19108), .ZN(n19088) );
  INV_X1 U13563 ( .A(n19165), .ZN(n18829) );
  INV_X1 U13564 ( .A(n18790), .ZN(n18851) );
  INV_X1 U13565 ( .A(n18811), .ZN(n18875) );
  INV_X1 U13566 ( .A(n18833), .ZN(n18897) );
  INV_X1 U13567 ( .A(n18879), .ZN(n18944) );
  INV_X1 U13568 ( .A(n18902), .ZN(n18965) );
  NOR2_X1 U13569 ( .A1(n19189), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19016) );
  INV_X1 U13570 ( .A(n18969), .ZN(n19032) );
  INV_X1 U13571 ( .A(n18992), .ZN(n19054) );
  INV_X1 U13572 ( .A(n19014), .ZN(n19078) );
  AND2_X1 U13573 ( .A1(n16992), .A2(BUF2_REG_21__SCAN_IN), .ZN(n19144) );
  OR2_X2 U13574 ( .A1(n12129), .A2(n12128), .ZN(n18783) );
  NOR2_X1 U13575 ( .A1(n19338), .A2(n19349), .ZN(n19341) );
  INV_X1 U13576 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n19235) );
  INV_X1 U13577 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n17353) );
  NAND2_X2 U13578 ( .A1(n13574), .A2(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19430)
         );
  INV_X1 U13579 ( .A(U212), .ZN(n17313) );
  NOR2_X1 U13580 ( .A1(n13434), .A2(n13433), .ZN(n13435) );
  INV_X1 U13581 ( .A(n15331), .ZN(n14977) );
  OAI21_X1 U13582 ( .B1(n14802), .B2(n9635), .A(n14801), .ZN(n15204) );
  AND2_X1 U13583 ( .A1(n14404), .A2(n14403), .ZN(n20630) );
  AND2_X1 U13584 ( .A1(n14398), .A2(n14397), .ZN(n20619) );
  INV_X1 U13585 ( .A(n20453), .ZN(n20475) );
  NOR2_X1 U13586 ( .A1(n14372), .A2(n14371), .ZN(n14379) );
  NAND2_X1 U13587 ( .A1(n20338), .A2(n13273), .ZN(n17161) );
  OR2_X2 U13588 ( .A1(n17128), .A2(n20330), .ZN(n20338) );
  INV_X1 U13589 ( .A(n20560), .ZN(n20575) );
  AND2_X1 U13590 ( .A1(n15567), .A2(n20729), .ZN(n21382) );
  OR2_X1 U13591 ( .A1(n20697), .A2(n20959), .ZN(n20660) );
  OR2_X1 U13592 ( .A1(n20697), .A2(n20995), .ZN(n20692) );
  OR2_X1 U13593 ( .A1(n20697), .A2(n21016), .ZN(n20723) );
  OR2_X1 U13594 ( .A1(n20697), .A2(n20926), .ZN(n20751) );
  OR2_X1 U13595 ( .A1(n20807), .A2(n20959), .ZN(n20777) );
  OR2_X1 U13596 ( .A1(n20807), .A2(n20995), .ZN(n20798) );
  OR2_X1 U13597 ( .A1(n20807), .A2(n20926), .ZN(n20831) );
  NAND2_X1 U13598 ( .A1(n20928), .A2(n20838), .ZN(n20892) );
  NAND2_X1 U13599 ( .A1(n20928), .A2(n20893), .ZN(n20957) );
  NAND2_X1 U13600 ( .A1(n20928), .A2(n20927), .ZN(n20987) );
  OR2_X1 U13601 ( .A1(n21017), .A2(n20959), .ZN(n21015) );
  OR2_X1 U13602 ( .A1(n21017), .A2(n21016), .ZN(n21131) );
  NAND2_X1 U13603 ( .A1(n13636), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21134) );
  INV_X1 U13604 ( .A(n21136), .ZN(n21204) );
  OR2_X1 U13605 ( .A1(n21151), .A2(n21198), .ZN(n21179) );
  INV_X1 U13606 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n20272) );
  NAND2_X1 U13607 ( .A1(n11443), .A2(n17236), .ZN(n13624) );
  OR2_X1 U13608 ( .A1(n14600), .A2(n15911), .ZN(n13499) );
  NAND2_X1 U13609 ( .A1(n19538), .A2(n20272), .ZN(n15911) );
  INV_X1 U13610 ( .A(n19477), .ZN(n16191) );
  AND2_X1 U13611 ( .A1(n13902), .A2(n17236), .ZN(n19445) );
  NAND2_X1 U13612 ( .A1(n19445), .A2(n13903), .ZN(n19472) );
  OR2_X1 U13613 ( .A1(n19523), .A2(n20312), .ZN(n13794) );
  OR2_X1 U13614 ( .A1(n13712), .A2(n10955), .ZN(n20310) );
  NAND2_X1 U13615 ( .A1(n13711), .A2(n20313), .ZN(n19523) );
  NAND2_X1 U13616 ( .A1(n13633), .A2(n11716), .ZN(n14059) );
  INV_X1 U13617 ( .A(n19538), .ZN(n19569) );
  INV_X1 U13618 ( .A(n11871), .ZN(n11872) );
  OR2_X1 U13619 ( .A1(n13624), .A2(n15992), .ZN(n19590) );
  NAND2_X1 U13620 ( .A1(n11519), .A2(n17209), .ZN(n11522) );
  INV_X1 U13621 ( .A(n17224), .ZN(n16737) );
  INV_X1 U13622 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20284) );
  OR2_X1 U13623 ( .A1(n19914), .A2(n19804), .ZN(n19680) );
  AND2_X1 U13624 ( .A1(n19812), .A2(n19811), .ZN(n19821) );
  OR2_X1 U13625 ( .A1(n19840), .A2(n20043), .ZN(n19839) );
  OR2_X1 U13626 ( .A1(n19840), .A2(n20131), .ZN(n19909) );
  INV_X1 U13627 ( .A(n19952), .ZN(n20006) );
  AOI21_X1 U13628 ( .B1(n16824), .B2(n16825), .A(n16823), .ZN(n20035) );
  INV_X1 U13629 ( .A(n20182), .ZN(n20123) );
  NAND2_X1 U13630 ( .A1(n20070), .A2(n20069), .ZN(n20170) );
  AND2_X1 U13631 ( .A1(n10837), .A2(n13774), .ZN(n20297) );
  INV_X1 U13632 ( .A(n20267), .ZN(n20189) );
  AOI211_X1 U13633 ( .C1(n17404), .C2(n17742), .A(n17394), .B(n17393), .ZN(
        n17395) );
  INV_X1 U13634 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18464) );
  INV_X1 U13635 ( .A(n17700), .ZN(n17726) );
  AND2_X1 U13636 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17890), .ZN(n17884) );
  NOR2_X1 U13637 ( .A1(n17864), .A2(n17895), .ZN(n17901) );
  AND2_X1 U13638 ( .A1(n18007), .A2(n18783), .ZN(n18016) );
  AND2_X1 U13639 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n14183), .ZN(n14236) );
  INV_X1 U13640 ( .A(n18099), .ZN(n14182) );
  NAND2_X1 U13641 ( .A1(n19342), .A2(n18172), .ZN(n18166) );
  OR2_X1 U13642 ( .A1(n18234), .A2(n18178), .ZN(n18230) );
  INV_X1 U13643 ( .A(n18405), .ZN(n18380) );
  INV_X1 U13644 ( .A(n18320), .ZN(n18350) );
  INV_X1 U13645 ( .A(n18428), .ZN(n18451) );
  INV_X1 U13646 ( .A(n18724), .ZN(n18616) );
  OR2_X1 U13647 ( .A1(n18724), .A2(n18693), .ZN(n18729) );
  OR2_X1 U13648 ( .A1(n19183), .A2(n18616), .ZN(n18734) );
  INV_X1 U13649 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19189) );
  INV_X1 U13650 ( .A(n19104), .ZN(n19036) );
  NOR2_X1 U13651 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19232) );
  INV_X1 U13652 ( .A(n19319), .ZN(n19233) );
  INV_X1 U13653 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n21313) );
  NOR2_X1 U13654 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13575), .ZN(n17349)
         );
  INV_X1 U13655 ( .A(n17317), .ZN(n17316) );
  OAI211_X1 U13656 ( .C1(n15025), .C2(n20393), .A(n10407), .B(n13435), .ZN(
        P1_U2811) );
  AOI22_X1 U13657 ( .A1(n10821), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9601), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10426) );
  AOI22_X1 U13658 ( .A1(n11697), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11694), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10425) );
  AOI22_X1 U13659 ( .A1(n11728), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11700), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10424) );
  AOI22_X1 U13660 ( .A1(n11699), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9602), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10423) );
  NAND4_X1 U13661 ( .A1(n10426), .A2(n10425), .A3(n10424), .A4(n10423), .ZN(
        n10427) );
  AOI22_X1 U13662 ( .A1(n11697), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11694), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10430) );
  AOI22_X1 U13663 ( .A1(n11699), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11698), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10429) );
  AOI22_X1 U13664 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11700), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10428) );
  NAND4_X1 U13665 ( .A1(n10431), .A2(n10430), .A3(n10429), .A4(n10428), .ZN(
        n10432) );
  AOI22_X1 U13666 ( .A1(n11728), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n14215), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10435) );
  AOI22_X1 U13667 ( .A1(n11697), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11694), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10434) );
  AOI22_X1 U13668 ( .A1(n11699), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9598), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10433) );
  AOI22_X1 U13669 ( .A1(n11728), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11700), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10440) );
  AOI22_X1 U13670 ( .A1(n10821), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14215), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10439) );
  AOI22_X1 U13671 ( .A1(n11697), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11694), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10438) );
  AOI22_X1 U13672 ( .A1(n11699), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9599), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10437) );
  AND2_X2 U13673 ( .A1(n11699), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11676) );
  AOI22_X1 U13674 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10445) );
  NAND2_X1 U13675 ( .A1(n10821), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10834) );
  AND2_X1 U13676 ( .A1(n11698), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10590) );
  AOI22_X1 U13677 ( .A1(n11675), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10590), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10444) );
  AOI22_X1 U13678 ( .A1(n10548), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10443) );
  AND2_X2 U13679 ( .A1(n11700), .A2(n9910), .ZN(n10506) );
  AND2_X2 U13680 ( .A1(n11700), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10549) );
  AOI22_X1 U13681 ( .A1(n10506), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10549), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10442) );
  AND2_X2 U13682 ( .A1(n11728), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10651) );
  AND2_X2 U13683 ( .A1(n9625), .A2(n10441), .ZN(n11678) );
  AOI22_X1 U13684 ( .A1(n10651), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11678), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10453) );
  AND2_X1 U13685 ( .A1(n11694), .A2(n10441), .ZN(n10505) );
  AOI22_X1 U13686 ( .A1(n10505), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10578), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10452) );
  NOR2_X2 U13687 ( .A1(n10980), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11692) );
  INV_X1 U13688 ( .A(n10447), .ZN(n14211) );
  AND2_X2 U13689 ( .A1(n11692), .A2(n10447), .ZN(n11664) );
  AOI22_X1 U13690 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11664), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10451) );
  NAND2_X1 U13691 ( .A1(n10783), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n16776) );
  INV_X1 U13692 ( .A(n16776), .ZN(n10448) );
  AND2_X2 U13693 ( .A1(n10448), .A2(n11692), .ZN(n11685) );
  AND2_X2 U13694 ( .A1(n11692), .A2(n10449), .ZN(n11684) );
  AOI22_X1 U13695 ( .A1(n11685), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11684), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10450) );
  NAND3_X1 U13696 ( .A1(n10416), .A2(n10453), .A3(n10402), .ZN(n17218) );
  NAND2_X1 U13697 ( .A1(n10454), .A2(n17218), .ZN(n10474) );
  AOI22_X1 U13698 ( .A1(n11728), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14215), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10458) );
  AOI22_X1 U13699 ( .A1(n11697), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11694), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10457) );
  AOI22_X1 U13700 ( .A1(n10821), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11700), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10456) );
  AOI22_X1 U13701 ( .A1(n11699), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11698), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10455) );
  NAND4_X1 U13702 ( .A1(n10458), .A2(n10457), .A3(n10456), .A4(n10455), .ZN(
        n10464) );
  AOI22_X1 U13703 ( .A1(n11728), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14215), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10462) );
  AOI22_X1 U13704 ( .A1(n11697), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11694), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10461) );
  AOI22_X1 U13705 ( .A1(n9625), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11700), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10460) );
  AOI22_X1 U13706 ( .A1(n11699), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9603), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10459) );
  NAND4_X1 U13707 ( .A1(n10462), .A2(n10461), .A3(n10460), .A4(n10459), .ZN(
        n10463) );
  AOI22_X1 U13708 ( .A1(n11697), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11694), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10466) );
  AOI22_X1 U13709 ( .A1(n11699), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9602), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10465) );
  AOI22_X1 U13710 ( .A1(n9625), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11700), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10467) );
  AOI22_X1 U13711 ( .A1(n11697), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11694), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10469) );
  AOI22_X1 U13712 ( .A1(n11699), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9602), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10468) );
  AOI22_X1 U13713 ( .A1(n11728), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14215), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10471) );
  AOI22_X1 U13714 ( .A1(n10821), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11700), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10470) );
  INV_X1 U13715 ( .A(n10889), .ZN(n10472) );
  NAND2_X1 U13716 ( .A1(n13903), .A2(n10479), .ZN(n10514) );
  NAND2_X1 U13717 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10473) );
  NAND2_X1 U13718 ( .A1(n10516), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10478) );
  NAND2_X1 U13719 ( .A1(n15992), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10476) );
  INV_X1 U13720 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n10475) );
  AND2_X1 U13721 ( .A1(n10476), .A2(n9723), .ZN(n10477) );
  NAND2_X1 U13722 ( .A1(n10478), .A2(n10477), .ZN(n14354) );
  NAND2_X1 U13723 ( .A1(n10516), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n10481) );
  INV_X1 U13724 ( .A(n10526), .ZN(n10517) );
  NAND2_X1 U13725 ( .A1(n10481), .A2(n10480), .ZN(n10498) );
  XNOR2_X1 U13726 ( .A(n10497), .B(n10498), .ZN(n14350) );
  AOI22_X1 U13727 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n11678), .B1(
        n10651), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10486) );
  AOI22_X1 U13728 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10485) );
  AOI22_X1 U13729 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n10506), .B1(
        n11677), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10484) );
  AOI22_X1 U13730 ( .A1(n11675), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10483) );
  NAND4_X1 U13731 ( .A1(n10486), .A2(n10485), .A3(n10484), .A4(n10483), .ZN(
        n10492) );
  AOI22_X1 U13732 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n11683), .B1(
        n10578), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10490) );
  AOI22_X1 U13733 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10548), .B1(
        n10549), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10489) );
  AOI22_X1 U13734 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n11685), .B1(
        n11684), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10488) );
  AOI22_X1 U13735 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10507), .B1(
        n11664), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10487) );
  NAND4_X1 U13736 ( .A1(n10490), .A2(n10489), .A3(n10488), .A4(n10487), .ZN(
        n10491) );
  NAND2_X1 U13737 ( .A1(n11033), .A2(n9571), .ZN(n11087) );
  INV_X1 U13738 ( .A(n13772), .ZN(n10495) );
  MUX2_X1 U13739 ( .A(n10493), .B(n19911), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n10494) );
  OAI21_X1 U13740 ( .B1(n11087), .B2(n10495), .A(n10494), .ZN(n10496) );
  INV_X1 U13741 ( .A(n10496), .ZN(n14349) );
  NAND2_X1 U13742 ( .A1(n14350), .A2(n14349), .ZN(n14352) );
  INV_X1 U13743 ( .A(n10498), .ZN(n10499) );
  NAND2_X1 U13744 ( .A1(n14353), .A2(n10499), .ZN(n10500) );
  NAND2_X1 U13745 ( .A1(n14352), .A2(n10500), .ZN(n10522) );
  AOI22_X1 U13746 ( .A1(n11675), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10504) );
  AOI22_X1 U13747 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10503) );
  AOI22_X1 U13748 ( .A1(n10651), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10549), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10502) );
  AOI22_X1 U13749 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10548), .B1(
        n10590), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10501) );
  NAND4_X1 U13750 ( .A1(n10504), .A2(n10503), .A3(n10502), .A4(n10501), .ZN(
        n10513) );
  AOI22_X1 U13751 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n10505), .B1(
        n10578), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10511) );
  AOI22_X1 U13752 ( .A1(n11678), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10506), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10510) );
  AOI22_X1 U13753 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n11685), .B1(
        n11684), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10509) );
  AOI22_X1 U13754 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10507), .B1(
        n11664), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10508) );
  NAND4_X1 U13755 ( .A1(n10511), .A2(n10510), .A3(n10509), .A4(n10508), .ZN(
        n10512) );
  OR2_X1 U13756 ( .A1(n10730), .A2(n11038), .ZN(n10515) );
  OAI211_X1 U13757 ( .C1(n20306), .C2(n20293), .A(n10515), .B(n10514), .ZN(
        n10520) );
  XNOR2_X1 U13758 ( .A(n10522), .B(n10520), .ZN(n14346) );
  NAND2_X1 U13759 ( .A1(n10765), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n10519) );
  AOI22_X1 U13760 ( .A1(n10703), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n10768), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10518) );
  AND2_X1 U13761 ( .A1(n10519), .A2(n10518), .ZN(n14345) );
  INV_X1 U13762 ( .A(n10520), .ZN(n10521) );
  NAND2_X1 U13763 ( .A1(n10522), .A2(n10521), .ZN(n10523) );
  NAND2_X1 U13764 ( .A1(n14348), .A2(n10523), .ZN(n14358) );
  INV_X1 U13765 ( .A(n14358), .ZN(n10543) );
  NAND2_X1 U13766 ( .A1(n10765), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n10541) );
  INV_X1 U13767 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19515) );
  NAND2_X1 U13768 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10525) );
  NAND2_X1 U13769 ( .A1(n10479), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10524) );
  OAI211_X1 U13770 ( .C1(n10526), .C2(n19515), .A(n10525), .B(n10524), .ZN(
        n10527) );
  INV_X1 U13771 ( .A(n10527), .ZN(n10540) );
  AOI22_X1 U13772 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n11675), .B1(
        n11676), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10531) );
  AOI22_X1 U13773 ( .A1(n10594), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11677), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10530) );
  AOI22_X1 U13774 ( .A1(n11678), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10529) );
  AOI22_X1 U13775 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10548), .B1(
        n10549), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10528) );
  NAND4_X1 U13776 ( .A1(n10531), .A2(n10530), .A3(n10529), .A4(n10528), .ZN(
        n10537) );
  AOI22_X1 U13777 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n11683), .B1(
        n10578), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10535) );
  AOI22_X1 U13778 ( .A1(n10651), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10506), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10534) );
  AOI22_X1 U13779 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n11685), .B1(
        n11684), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10533) );
  AOI22_X1 U13780 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10507), .B1(
        n11664), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10532) );
  NAND4_X1 U13781 ( .A1(n10535), .A2(n10534), .A3(n10533), .A4(n10532), .ZN(
        n10536) );
  INV_X1 U13782 ( .A(n11092), .ZN(n10538) );
  OR2_X1 U13783 ( .A1(n10730), .A2(n10538), .ZN(n10539) );
  INV_X1 U13784 ( .A(n14357), .ZN(n10542) );
  NAND2_X1 U13785 ( .A1(n10543), .A2(n10542), .ZN(n14356) );
  NAND2_X1 U13786 ( .A1(n10765), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n10558) );
  AOI22_X1 U13787 ( .A1(n10703), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n10768), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10557) );
  AOI22_X1 U13788 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n11678), .B1(
        n10651), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10547) );
  AOI22_X1 U13789 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n11683), .B1(
        n10578), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10546) );
  AOI22_X1 U13790 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n11685), .B1(
        n11684), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10545) );
  AOI22_X1 U13791 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10507), .B1(
        n11664), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10544) );
  NAND4_X1 U13792 ( .A1(n10547), .A2(n10546), .A3(n10545), .A4(n10544), .ZN(
        n10555) );
  AOI22_X1 U13793 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10553) );
  AOI22_X1 U13794 ( .A1(n11675), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11677), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10552) );
  AOI22_X1 U13795 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10548), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10551) );
  AOI22_X1 U13796 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10506), .B1(
        n10549), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10550) );
  NAND4_X1 U13797 ( .A1(n10553), .A2(n10552), .A3(n10551), .A4(n10550), .ZN(
        n10554) );
  INV_X1 U13798 ( .A(n11093), .ZN(n11031) );
  OR2_X1 U13799 ( .A1(n10730), .A2(n11031), .ZN(n10556) );
  AOI22_X1 U13800 ( .A1(n10651), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11678), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10562) );
  AOI22_X1 U13801 ( .A1(n11683), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10578), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10561) );
  AOI22_X1 U13802 ( .A1(n11685), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11684), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10560) );
  AOI22_X1 U13803 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11664), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10559) );
  NAND4_X1 U13804 ( .A1(n10562), .A2(n10561), .A3(n10560), .A4(n10559), .ZN(
        n10568) );
  AOI22_X1 U13805 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10566) );
  AOI22_X1 U13806 ( .A1(n11675), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11677), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10565) );
  AOI22_X1 U13807 ( .A1(n10548), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10564) );
  AOI22_X1 U13808 ( .A1(n10506), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10549), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10563) );
  NAND4_X1 U13809 ( .A1(n10566), .A2(n10565), .A3(n10564), .A4(n10563), .ZN(
        n10567) );
  NAND2_X1 U13810 ( .A1(n10765), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n10570) );
  AOI22_X1 U13811 ( .A1(n10703), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n10768), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10569) );
  OAI211_X1 U13812 ( .C1(n10730), .C2(n11063), .A(n10570), .B(n10569), .ZN(
        n15913) );
  NAND2_X1 U13813 ( .A1(n14360), .A2(n15913), .ZN(n15912) );
  AOI22_X1 U13814 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10574) );
  AOI22_X1 U13815 ( .A1(n11675), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11677), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10573) );
  AOI22_X1 U13816 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10548), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10572) );
  AOI22_X1 U13817 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10506), .B1(
        n10549), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10571) );
  NAND4_X1 U13818 ( .A1(n10574), .A2(n10573), .A3(n10572), .A4(n10571), .ZN(
        n10586) );
  INV_X1 U13819 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11815) );
  INV_X1 U13820 ( .A(n11678), .ZN(n10577) );
  INV_X1 U13821 ( .A(n10651), .ZN(n10576) );
  INV_X1 U13822 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10575) );
  OAI22_X1 U13823 ( .A1(n11815), .A2(n10577), .B1(n10576), .B2(n10575), .ZN(
        n10584) );
  AOI22_X1 U13824 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n11685), .B1(
        n11684), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10582) );
  AOI22_X1 U13825 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10507), .B1(
        n11664), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10581) );
  NAND2_X1 U13826 ( .A1(n10578), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n10580) );
  NAND2_X1 U13827 ( .A1(n11683), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n10579) );
  NAND4_X1 U13828 ( .A1(n10582), .A2(n10581), .A3(n10580), .A4(n10579), .ZN(
        n10583) );
  OR2_X1 U13829 ( .A1(n10730), .A2(n11098), .ZN(n10587) );
  NAND2_X1 U13830 ( .A1(n10765), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n10589) );
  AOI22_X1 U13831 ( .A1(n10703), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n10768), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n10588) );
  NAND2_X1 U13832 ( .A1(n10589), .A2(n10588), .ZN(n15906) );
  NAND2_X1 U13833 ( .A1(n15907), .A2(n15906), .ZN(n15905) );
  INV_X1 U13834 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10593) );
  INV_X1 U13835 ( .A(n10590), .ZN(n10592) );
  INV_X1 U13836 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10591) );
  OAI22_X1 U13837 ( .A1(n10834), .A2(n10593), .B1(n10592), .B2(n10591), .ZN(
        n10599) );
  INV_X1 U13838 ( .A(n11676), .ZN(n10597) );
  INV_X1 U13839 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10596) );
  INV_X1 U13840 ( .A(n10594), .ZN(n10595) );
  INV_X1 U13841 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11845) );
  OAI22_X1 U13842 ( .A1(n10597), .A2(n10596), .B1(n10595), .B2(n11845), .ZN(
        n10598) );
  NOR2_X1 U13843 ( .A1(n10599), .A2(n10598), .ZN(n10612) );
  AOI22_X1 U13844 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n11685), .B1(
        n11684), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10603) );
  AOI22_X1 U13845 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n10507), .B1(
        n11664), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10602) );
  NAND2_X1 U13846 ( .A1(n10578), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10601) );
  NAND2_X1 U13847 ( .A1(n11683), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10600) );
  NAND2_X1 U13848 ( .A1(n11678), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10605) );
  NAND2_X1 U13849 ( .A1(n10651), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10604) );
  NAND2_X1 U13850 ( .A1(n10482), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10609) );
  NAND2_X1 U13851 ( .A1(n10548), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10608) );
  NAND2_X1 U13852 ( .A1(n10549), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10607) );
  NAND2_X1 U13853 ( .A1(n10506), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10606) );
  OR2_X1 U13854 ( .A1(n10730), .A2(n16378), .ZN(n10613) );
  NAND2_X1 U13855 ( .A1(n15905), .A2(n10613), .ZN(n13892) );
  NAND2_X1 U13856 ( .A1(n10765), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n10615) );
  AOI22_X1 U13857 ( .A1(n10703), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n10768), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n10614) );
  NAND2_X1 U13858 ( .A1(n10615), .A2(n10614), .ZN(n13894) );
  NAND2_X1 U13859 ( .A1(n10765), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n10629) );
  AOI22_X1 U13860 ( .A1(n10703), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n10768), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10628) );
  AOI22_X1 U13861 ( .A1(n11675), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10619) );
  AOI22_X1 U13862 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10618) );
  AOI22_X1 U13863 ( .A1(n10506), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11677), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10617) );
  AOI22_X1 U13864 ( .A1(n11678), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10549), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10616) );
  NAND4_X1 U13865 ( .A1(n10619), .A2(n10618), .A3(n10617), .A4(n10616), .ZN(
        n10625) );
  AOI22_X1 U13866 ( .A1(n11683), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10578), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10623) );
  AOI22_X1 U13867 ( .A1(n10651), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10548), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10622) );
  AOI22_X1 U13868 ( .A1(n11685), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11684), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10621) );
  AOI22_X1 U13869 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11664), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10620) );
  NAND4_X1 U13870 ( .A1(n10623), .A2(n10622), .A3(n10621), .A4(n10620), .ZN(
        n10624) );
  INV_X1 U13871 ( .A(n14326), .ZN(n10626) );
  OR2_X1 U13872 ( .A1(n10730), .A2(n10626), .ZN(n10627) );
  NAND2_X1 U13873 ( .A1(n10765), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n10644) );
  AOI22_X1 U13874 ( .A1(n10703), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n10768), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10643) );
  AOI22_X1 U13875 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11678), .B1(
        n10651), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10634) );
  AOI22_X1 U13876 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n11683), .B1(
        n10578), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10633) );
  AOI22_X1 U13877 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n11685), .B1(
        n11684), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10632) );
  AOI22_X1 U13878 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10507), .B1(
        n11664), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10631) );
  NAND4_X1 U13879 ( .A1(n10634), .A2(n10633), .A3(n10632), .A4(n10631), .ZN(
        n10641) );
  AOI22_X1 U13880 ( .A1(n11675), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n11677), .ZN(n10639) );
  AOI22_X1 U13881 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10638) );
  AOI22_X1 U13882 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10548), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10637) );
  INV_X1 U13883 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10635) );
  AOI22_X1 U13884 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n10506), .B1(
        n10549), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10636) );
  NAND4_X1 U13885 ( .A1(n10639), .A2(n10638), .A3(n10637), .A4(n10636), .ZN(
        n10640) );
  OR2_X1 U13886 ( .A1(n10730), .A2(n16055), .ZN(n10642) );
  NAND2_X1 U13887 ( .A1(n10646), .A2(n10645), .ZN(n14200) );
  NAND2_X1 U13888 ( .A1(n10765), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n10661) );
  AOI22_X1 U13889 ( .A1(n10703), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n10768), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n10660) );
  AOI22_X1 U13890 ( .A1(n11675), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_9__2__SCAN_IN), .B2(n10482), .ZN(n10650) );
  AOI22_X1 U13891 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10649) );
  AOI22_X1 U13892 ( .A1(n11678), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11677), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10648) );
  AOI22_X1 U13893 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10548), .B1(
        n10549), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10647) );
  NAND4_X1 U13894 ( .A1(n10650), .A2(n10649), .A3(n10648), .A4(n10647), .ZN(
        n10657) );
  AOI22_X1 U13895 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n11683), .B1(
        n10578), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10655) );
  AOI22_X1 U13896 ( .A1(n10651), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10506), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10654) );
  AOI22_X1 U13897 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n11685), .B1(
        n11684), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10653) );
  AOI22_X1 U13898 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10507), .B1(
        n11664), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10652) );
  NAND4_X1 U13899 ( .A1(n10655), .A2(n10654), .A3(n10653), .A4(n10652), .ZN(
        n10656) );
  INV_X1 U13900 ( .A(n16069), .ZN(n10658) );
  OR2_X1 U13901 ( .A1(n10730), .A2(n10658), .ZN(n10659) );
  INV_X1 U13902 ( .A(n10662), .ZN(n14199) );
  NAND2_X1 U13903 ( .A1(n10765), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n10675) );
  AOI22_X1 U13904 ( .A1(n10703), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n10768), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10674) );
  AOI22_X1 U13905 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n11678), .B1(
        n10651), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10666) );
  AOI22_X1 U13906 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n11683), .B1(
        n10578), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10665) );
  AOI22_X1 U13907 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n11685), .B1(
        n11684), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10664) );
  AOI22_X1 U13908 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10507), .B1(
        n11664), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10663) );
  NAND4_X1 U13909 ( .A1(n10666), .A2(n10665), .A3(n10664), .A4(n10663), .ZN(
        n10672) );
  AOI22_X1 U13910 ( .A1(n11675), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__3__SCAN_IN), .B2(n10590), .ZN(n10670) );
  AOI22_X1 U13911 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10669) );
  AOI22_X1 U13912 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n10548), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10668) );
  AOI22_X1 U13913 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n10506), .B1(
        n10549), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10667) );
  NAND4_X1 U13914 ( .A1(n10670), .A2(n10669), .A3(n10668), .A4(n10667), .ZN(
        n10671) );
  OR2_X1 U13915 ( .A1(n10672), .A2(n10671), .ZN(n11593) );
  INV_X1 U13916 ( .A(n11593), .ZN(n16063) );
  OR2_X1 U13917 ( .A1(n10730), .A2(n16063), .ZN(n10673) );
  NOR2_X2 U13918 ( .A1(n14199), .A2(n15829), .ZN(n14282) );
  INV_X1 U13919 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n20226) );
  AOI22_X1 U13920 ( .A1(n10703), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n10768), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n10687) );
  AOI22_X1 U13921 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n11678), .B1(
        n10651), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10679) );
  AOI22_X1 U13922 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n11683), .B1(
        n10578), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10678) );
  AOI22_X1 U13923 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n11685), .B1(
        n11684), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10677) );
  AOI22_X1 U13924 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10507), .B1(
        n11664), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10676) );
  NAND4_X1 U13925 ( .A1(n10679), .A2(n10678), .A3(n10677), .A4(n10676), .ZN(
        n10685) );
  AOI22_X1 U13926 ( .A1(n11675), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_8__4__SCAN_IN), .B2(n10506), .ZN(n10683) );
  AOI22_X1 U13927 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10682) );
  AOI22_X1 U13928 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n10482), .B1(
        n11677), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10681) );
  AOI22_X1 U13929 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10548), .B1(
        n10549), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10680) );
  NAND4_X1 U13930 ( .A1(n10683), .A2(n10682), .A3(n10681), .A4(n10680), .ZN(
        n10684) );
  OR2_X1 U13931 ( .A1(n10685), .A2(n10684), .ZN(n16058) );
  NAND2_X1 U13932 ( .A1(n10454), .A2(n16058), .ZN(n10686) );
  OAI211_X1 U13933 ( .C1(n10688), .C2(n20226), .A(n10687), .B(n10686), .ZN(
        n14284) );
  NAND2_X1 U13934 ( .A1(n10765), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n10701) );
  AOI22_X1 U13935 ( .A1(n10703), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n10768), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10700) );
  AOI22_X1 U13936 ( .A1(n10651), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11678), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10692) );
  AOI22_X1 U13937 ( .A1(n11683), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10578), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10691) );
  AOI22_X1 U13938 ( .A1(n11685), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11684), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10690) );
  AOI22_X1 U13939 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11664), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10689) );
  NAND4_X1 U13940 ( .A1(n10692), .A2(n10691), .A3(n10690), .A4(n10689), .ZN(
        n10698) );
  AOI22_X1 U13941 ( .A1(n11675), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10590), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10696) );
  AOI22_X1 U13942 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10695) );
  AOI22_X1 U13943 ( .A1(n10548), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10694) );
  AOI22_X1 U13944 ( .A1(n10506), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10549), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10693) );
  NAND4_X1 U13945 ( .A1(n10696), .A2(n10695), .A3(n10694), .A4(n10693), .ZN(
        n10697) );
  OR2_X1 U13946 ( .A1(n10698), .A2(n10697), .ZN(n11607) );
  INV_X1 U13947 ( .A(n11607), .ZN(n14424) );
  OR2_X1 U13948 ( .A1(n10730), .A2(n14424), .ZN(n10699) );
  NAND2_X1 U13949 ( .A1(n10765), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n10717) );
  AOI22_X1 U13950 ( .A1(n10703), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n10768), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n10716) );
  AOI22_X1 U13951 ( .A1(n11675), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11678), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10707) );
  AOI22_X1 U13952 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n10651), .B1(
        n11676), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10706) );
  AOI22_X1 U13953 ( .A1(n10594), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10590), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10705) );
  AOI22_X1 U13954 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10548), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10704) );
  NAND4_X1 U13955 ( .A1(n10707), .A2(n10706), .A3(n10705), .A4(n10704), .ZN(
        n10713) );
  AOI22_X1 U13956 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n10578), .B1(
        n11683), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10711) );
  AOI22_X1 U13957 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10549), .B1(
        n10506), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10710) );
  AOI22_X1 U13958 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n11685), .B1(
        n11684), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10709) );
  AOI22_X1 U13959 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n10507), .B1(
        n11664), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10708) );
  NAND4_X1 U13960 ( .A1(n10711), .A2(n10710), .A3(n10709), .A4(n10708), .ZN(
        n10712) );
  INV_X1 U13961 ( .A(n14425), .ZN(n10714) );
  OR2_X1 U13962 ( .A1(n10730), .A2(n10714), .ZN(n10715) );
  AOI22_X1 U13963 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n11678), .B1(
        n10651), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10721) );
  AOI22_X1 U13964 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n11683), .B1(
        n10578), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10720) );
  AOI22_X1 U13965 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n11685), .B1(
        n11684), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10719) );
  AOI22_X1 U13966 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10507), .B1(
        n11664), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10718) );
  NAND4_X1 U13967 ( .A1(n10721), .A2(n10720), .A3(n10719), .A4(n10718), .ZN(
        n10727) );
  AOI22_X1 U13968 ( .A1(n11675), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__7__SCAN_IN), .B2(n10590), .ZN(n10725) );
  AOI22_X1 U13969 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10724) );
  AOI22_X1 U13970 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10548), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10723) );
  AOI22_X1 U13971 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n10506), .B1(
        n10549), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10722) );
  NAND4_X1 U13972 ( .A1(n10725), .A2(n10724), .A3(n10723), .A4(n10722), .ZN(
        n10726) );
  OR2_X1 U13973 ( .A1(n10727), .A2(n10726), .ZN(n11608) );
  INV_X1 U13974 ( .A(n11608), .ZN(n16047) );
  NAND2_X1 U13975 ( .A1(n10765), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n10729) );
  AOI22_X1 U13976 ( .A1(n10703), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n10768), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n10728) );
  OAI211_X1 U13977 ( .C1(n10730), .C2(n16047), .A(n10729), .B(n10728), .ZN(
        n16589) );
  NAND2_X1 U13978 ( .A1(n10765), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n10732) );
  AOI22_X1 U13979 ( .A1(n10703), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n10768), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10731) );
  NAND2_X1 U13980 ( .A1(n10732), .A2(n10731), .ZN(n15780) );
  NAND2_X1 U13981 ( .A1(n15778), .A2(n15780), .ZN(n15774) );
  INV_X1 U13982 ( .A(n15774), .ZN(n10736) );
  NAND2_X1 U13983 ( .A1(n10765), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n10734) );
  AOI22_X1 U13984 ( .A1(n10703), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n10768), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10733) );
  INV_X1 U13985 ( .A(n15775), .ZN(n10735) );
  NAND2_X1 U13986 ( .A1(n10736), .A2(n10735), .ZN(n15760) );
  NAND2_X1 U13987 ( .A1(n10765), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n10738) );
  AOI22_X1 U13988 ( .A1(n10703), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n10768), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n10737) );
  NAND2_X1 U13989 ( .A1(n10765), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n10741) );
  AOI22_X1 U13990 ( .A1(n10703), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n10768), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n10740) );
  NAND2_X1 U13991 ( .A1(n10765), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n10743) );
  AOI22_X1 U13992 ( .A1(n10703), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n10479), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n10742) );
  NAND2_X1 U13993 ( .A1(n10743), .A2(n10742), .ZN(n15721) );
  NAND2_X1 U13994 ( .A1(n10765), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n10745) );
  AOI22_X1 U13995 ( .A1(n10703), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n10479), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10744) );
  NAND2_X1 U13996 ( .A1(n10745), .A2(n10744), .ZN(n15707) );
  AND2_X2 U13997 ( .A1(n15708), .A2(n15707), .ZN(n15690) );
  NAND2_X1 U13998 ( .A1(n10765), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n10747) );
  AOI22_X1 U13999 ( .A1(n10703), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n10479), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n10746) );
  NAND2_X1 U14000 ( .A1(n10747), .A2(n10746), .ZN(n15692) );
  NAND2_X1 U14001 ( .A1(n10765), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n10749) );
  AOI22_X1 U14002 ( .A1(n10703), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n10768), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n10748) );
  AND2_X1 U14003 ( .A1(n10749), .A2(n10748), .ZN(n15685) );
  NAND2_X1 U14004 ( .A1(n10765), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n10752) );
  AOI22_X1 U14005 ( .A1(n10703), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n10479), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10751) );
  NAND2_X1 U14006 ( .A1(n10765), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n10754) );
  AOI22_X1 U14007 ( .A1(n10703), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n10479), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n10753) );
  NAND2_X1 U14008 ( .A1(n10754), .A2(n10753), .ZN(n15648) );
  NAND2_X1 U14009 ( .A1(n10765), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n10756) );
  AOI22_X1 U14010 ( .A1(n10703), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n10479), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10755) );
  NAND2_X1 U14011 ( .A1(n10756), .A2(n10755), .ZN(n15635) );
  NAND2_X1 U14012 ( .A1(n10765), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n10758) );
  AOI22_X1 U14013 ( .A1(n10703), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n10479), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10757) );
  AND2_X1 U14014 ( .A1(n10758), .A2(n10757), .ZN(n15618) );
  INV_X1 U14015 ( .A(n15618), .ZN(n10759) );
  NAND2_X1 U14016 ( .A1(n10765), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n10762) );
  AOI22_X1 U14017 ( .A1(n10703), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n10479), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10761) );
  NAND2_X1 U14018 ( .A1(n10765), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n10764) );
  AOI22_X1 U14019 ( .A1(n10703), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n10479), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n10763) );
  NAND2_X1 U14020 ( .A1(n10764), .A2(n10763), .ZN(n15595) );
  NAND2_X1 U14021 ( .A1(n10765), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n10767) );
  AOI22_X1 U14022 ( .A1(n10703), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n10479), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10766) );
  AOI222_X1 U14023 ( .A1(n10765), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n10703), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n10768), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n10769) );
  AOI22_X1 U14024 ( .A1(n11728), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9625), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10773) );
  AOI22_X1 U14025 ( .A1(n11697), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11694), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10772) );
  AOI22_X1 U14026 ( .A1(n11699), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11698), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10771) );
  AOI22_X1 U14027 ( .A1(n11700), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9601), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10770) );
  AOI22_X1 U14028 ( .A1(n11728), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11700), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10774) );
  AOI22_X1 U14029 ( .A1(n9625), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14215), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10777) );
  AOI22_X1 U14030 ( .A1(n11699), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11698), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10776) );
  AOI22_X1 U14031 ( .A1(n11697), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11694), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10775) );
  NOR2_X1 U14032 ( .A1(n13713), .A2(n11716), .ZN(n10781) );
  NAND2_X1 U14033 ( .A1(n10786), .A2(n10782), .ZN(n10779) );
  NAND2_X1 U14034 ( .A1(n19911), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10778) );
  MUX2_X1 U14035 ( .A(n10781), .B(n10356), .S(n10829), .Z(n10792) );
  INV_X1 U14036 ( .A(n10782), .ZN(n10785) );
  NAND2_X1 U14037 ( .A1(n10783), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10784) );
  NAND2_X1 U14038 ( .A1(n11117), .A2(n10786), .ZN(n10870) );
  NAND2_X1 U14039 ( .A1(n10356), .A2(n10870), .ZN(n10790) );
  INV_X1 U14040 ( .A(n10829), .ZN(n10867) );
  XNOR2_X1 U14041 ( .A(n10786), .B(n10785), .ZN(n10826) );
  INV_X1 U14042 ( .A(n10826), .ZN(n10787) );
  OAI21_X1 U14043 ( .B1(n15992), .B2(n10867), .A(n10787), .ZN(n10788) );
  INV_X1 U14044 ( .A(n20311), .ZN(n10943) );
  OAI211_X1 U14045 ( .C1(n10829), .C2(n11117), .A(n10788), .B(n10943), .ZN(
        n10789) );
  AND2_X1 U14046 ( .A1(n10790), .A2(n10789), .ZN(n10791) );
  NOR2_X1 U14047 ( .A1(n10792), .A2(n10791), .ZN(n10802) );
  NAND2_X1 U14048 ( .A1(n10794), .A2(n10793), .ZN(n10796) );
  NAND2_X1 U14049 ( .A1(n20293), .A2(n10980), .ZN(n10795) );
  NAND2_X1 U14050 ( .A1(n10801), .A2(n10799), .ZN(n10798) );
  NAND2_X1 U14051 ( .A1(n20284), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10797) );
  NAND2_X1 U14052 ( .A1(n10798), .A2(n10797), .ZN(n10804) );
  INV_X1 U14053 ( .A(n10799), .ZN(n10800) );
  XNOR2_X1 U14054 ( .A(n10801), .B(n10800), .ZN(n11089) );
  NAND2_X1 U14055 ( .A1(n11094), .A2(n11089), .ZN(n10871) );
  MUX2_X1 U14056 ( .A(n10802), .B(n10356), .S(n10871), .Z(n10807) );
  NOR2_X1 U14057 ( .A1(n10833), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n10803) );
  NAND2_X1 U14058 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n10833), .ZN(
        n10805) );
  NOR2_X1 U14059 ( .A1(n10807), .A2(n10872), .ZN(n10808) );
  INV_X1 U14060 ( .A(n16846), .ZN(n13898) );
  NAND2_X1 U14061 ( .A1(n13898), .A2(n15992), .ZN(n13710) );
  NOR2_X1 U14062 ( .A1(n10810), .A2(n20311), .ZN(n10814) );
  AOI22_X1 U14063 ( .A1(n11728), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9601), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10811) );
  AOI22_X1 U14064 ( .A1(n11728), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9601), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10813) );
  AOI22_X1 U14065 ( .A1(n11700), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__4__SCAN_IN), .B2(n10821), .ZN(n10812) );
  NOR2_X1 U14066 ( .A1(n10814), .A2(n10901), .ZN(n10815) );
  NAND2_X1 U14067 ( .A1(n13710), .A2(n10815), .ZN(n10877) );
  INV_X1 U14068 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n20195) );
  NAND2_X2 U14069 ( .A1(n20260), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n20259) );
  NAND2_X1 U14070 ( .A1(n20190), .A2(n20208), .ZN(n20202) );
  NAND2_X1 U14071 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n20191) );
  AOI22_X1 U14072 ( .A1(n11728), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9601), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10819) );
  AOI22_X1 U14073 ( .A1(n11697), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11694), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10818) );
  AOI22_X1 U14074 ( .A1(n9625), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11700), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10817) );
  AOI22_X1 U14075 ( .A1(n11699), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9603), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10816) );
  AOI22_X1 U14076 ( .A1(n9625), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11700), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10825) );
  AOI22_X1 U14077 ( .A1(n11728), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9601), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10824) );
  AOI22_X1 U14078 ( .A1(n11697), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11694), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10823) );
  AOI22_X1 U14079 ( .A1(n11699), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11698), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10822) );
  INV_X1 U14080 ( .A(n10892), .ZN(n19614) );
  NAND2_X1 U14081 ( .A1(n14228), .A2(n19614), .ZN(n10852) );
  NAND2_X1 U14082 ( .A1(n10829), .A2(n10826), .ZN(n10828) );
  OAI21_X1 U14083 ( .B1(n10871), .B2(n10828), .A(n10827), .ZN(n16851) );
  NAND2_X1 U14084 ( .A1(n10829), .A2(n11117), .ZN(n10830) );
  OAI21_X1 U14085 ( .B1(n10871), .B2(n10830), .A(n10955), .ZN(n10831) );
  OR2_X1 U14086 ( .A1(n16851), .A2(n10831), .ZN(n10837) );
  AOI21_X1 U14087 ( .B1(n16785), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16852) );
  NAND2_X1 U14088 ( .A1(n10834), .A2(n16852), .ZN(n10835) );
  INV_X1 U14089 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n13625) );
  NAND2_X1 U14090 ( .A1(n10835), .A2(n13625), .ZN(n10836) );
  NAND2_X1 U14091 ( .A1(n10836), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13774) );
  AOI22_X1 U14092 ( .A1(n11697), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11694), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10842) );
  AOI22_X1 U14093 ( .A1(n11728), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n14215), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10841) );
  AOI22_X1 U14094 ( .A1(n10821), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11700), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10840) );
  AOI22_X1 U14095 ( .A1(n11699), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9603), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10839) );
  AOI22_X1 U14096 ( .A1(n10821), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11700), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10846) );
  AOI22_X1 U14097 ( .A1(n11728), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9601), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10845) );
  AOI22_X1 U14098 ( .A1(n11697), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11694), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10844) );
  AOI22_X1 U14099 ( .A1(n11699), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11698), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10843) );
  NAND2_X1 U14100 ( .A1(n10855), .A2(n10848), .ZN(n10879) );
  NAND2_X1 U14101 ( .A1(n11440), .A2(n16854), .ZN(n10851) );
  NAND2_X1 U14102 ( .A1(n10880), .A2(n15992), .ZN(n10850) );
  NAND3_X1 U14103 ( .A1(n10850), .A2(n20191), .A3(n13630), .ZN(n10865) );
  OAI211_X1 U14104 ( .C1(n16846), .C2(n10852), .A(n10851), .B(n10865), .ZN(
        n10853) );
  NAND2_X1 U14105 ( .A1(n10853), .A2(n10884), .ZN(n10876) );
  AND2_X1 U14106 ( .A1(n19614), .A2(n10903), .ZN(n10854) );
  NAND2_X1 U14107 ( .A1(n10893), .A2(n10892), .ZN(n10858) );
  NAND2_X1 U14108 ( .A1(n10857), .A2(n10858), .ZN(n10862) );
  NAND2_X1 U14109 ( .A1(n19624), .A2(n11716), .ZN(n10914) );
  NAND2_X1 U14110 ( .A1(n10914), .A2(n10943), .ZN(n10859) );
  AND2_X2 U14111 ( .A1(n10903), .A2(n10892), .ZN(n10946) );
  AOI21_X1 U14112 ( .B1(n10860), .B2(n10892), .A(n10946), .ZN(n10861) );
  AND2_X1 U14113 ( .A1(n11716), .A2(n20311), .ZN(n13436) );
  OAI21_X1 U14114 ( .B1(n10863), .B2(n13904), .A(n13436), .ZN(n10916) );
  NAND3_X1 U14115 ( .A1(n16864), .A2(n13630), .A3(n14228), .ZN(n10864) );
  NAND4_X1 U14116 ( .A1(n10894), .A2(n10918), .A3(n10916), .A4(n10864), .ZN(
        n14224) );
  NOR2_X1 U14117 ( .A1(n10865), .A2(n10892), .ZN(n10866) );
  NOR2_X1 U14118 ( .A1(n14224), .A2(n10866), .ZN(n10875) );
  NAND2_X1 U14119 ( .A1(n11083), .A2(n10870), .ZN(n10874) );
  INV_X1 U14120 ( .A(n10871), .ZN(n10873) );
  AOI21_X1 U14121 ( .B1(n10874), .B2(n10873), .A(n10872), .ZN(n20296) );
  NAND2_X1 U14122 ( .A1(n20296), .A2(n20299), .ZN(n11442) );
  NAND4_X1 U14123 ( .A1(n10877), .A2(n10876), .A3(n10875), .A4(n11442), .ZN(
        n10878) );
  NAND3_X1 U14124 ( .A1(n10879), .A2(n10892), .A3(n15992), .ZN(n10881) );
  INV_X1 U14125 ( .A(n10944), .ZN(n10886) );
  NAND2_X1 U14126 ( .A1(n9668), .A2(n20314), .ZN(n10882) );
  INV_X1 U14127 ( .A(n10945), .ZN(n10885) );
  NAND2_X1 U14128 ( .A1(n10886), .A2(n10953), .ZN(n14229) );
  NAND2_X1 U14129 ( .A1(n10857), .A2(n13485), .ZN(n16850) );
  NAND2_X1 U14130 ( .A1(n16850), .A2(n15992), .ZN(n10887) );
  NAND2_X1 U14131 ( .A1(n14229), .A2(n10887), .ZN(n10888) );
  MUX2_X1 U14132 ( .A(n10942), .B(n10892), .S(n20311), .Z(n10910) );
  NAND2_X1 U14133 ( .A1(n10900), .A2(n15992), .ZN(n16763) );
  NAND2_X1 U14134 ( .A1(n16763), .A2(n10916), .ZN(n10899) );
  INV_X1 U14135 ( .A(n10895), .ZN(n10896) );
  OAI21_X1 U14136 ( .B1(n10946), .B2(n19624), .A(n10896), .ZN(n10897) );
  INV_X1 U14137 ( .A(n10897), .ZN(n10898) );
  AOI21_X1 U14138 ( .B1(n10899), .B2(n19619), .A(n10898), .ZN(n10909) );
  NAND2_X1 U14139 ( .A1(n10900), .A2(n19619), .ZN(n10905) );
  AND2_X1 U14140 ( .A1(n10906), .A2(n11716), .ZN(n10941) );
  NOR2_X1 U14141 ( .A1(n10941), .A2(n10911), .ZN(n10907) );
  NAND2_X1 U14142 ( .A1(n10940), .A2(n10907), .ZN(n10908) );
  NAND2_X1 U14143 ( .A1(n16795), .A2(n9729), .ZN(n10913) );
  NAND2_X1 U14144 ( .A1(n11409), .A2(n10913), .ZN(n16562) );
  INV_X1 U14145 ( .A(n10914), .ZN(n10915) );
  AND2_X1 U14146 ( .A1(n10916), .A2(n10915), .ZN(n10917) );
  AND2_X2 U14147 ( .A1(n16562), .A2(n16515), .ZN(n17232) );
  INV_X1 U14148 ( .A(n16562), .ZN(n16518) );
  INV_X1 U14149 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11127) );
  NAND2_X1 U14150 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n16749) );
  NOR2_X1 U14151 ( .A1(n11127), .A2(n16749), .ZN(n10929) );
  INV_X1 U14152 ( .A(n10929), .ZN(n10920) );
  AND2_X2 U14153 ( .A1(n20305), .A2(n20307), .ZN(n19571) );
  NOR2_X1 U14154 ( .A1(n11409), .A2(n19571), .ZN(n17216) );
  INV_X1 U14155 ( .A(n16749), .ZN(n14616) );
  NOR3_X1 U14156 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n14616), .A3(
        n16515), .ZN(n10919) );
  INV_X1 U14157 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n21322) );
  NAND3_X1 U14158 ( .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16699) );
  NOR2_X1 U14159 ( .A1(n21322), .A2(n16699), .ZN(n16673) );
  NAND2_X1 U14160 ( .A1(n17212), .A2(n16673), .ZN(n16672) );
  NAND2_X1 U14161 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16674) );
  INV_X1 U14162 ( .A(n17216), .ZN(n10921) );
  AND2_X1 U14163 ( .A1(n10921), .A2(n17232), .ZN(n16713) );
  INV_X1 U14164 ( .A(n16713), .ZN(n16671) );
  OAI21_X1 U14165 ( .B1(n16672), .B2(n16674), .A(n16671), .ZN(n16666) );
  INV_X1 U14166 ( .A(n17232), .ZN(n16750) );
  AND2_X1 U14167 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16310) );
  AND2_X1 U14168 ( .A1(n16310), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11549) );
  AND2_X1 U14169 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16571) );
  AND2_X1 U14170 ( .A1(n16571), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11555) );
  NAND4_X1 U14171 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A4(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10922) );
  NAND2_X1 U14172 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16637) );
  NOR2_X1 U14173 ( .A1(n10922), .A2(n16637), .ZN(n10923) );
  AND3_X1 U14174 ( .A1(n11549), .A2(n11555), .A3(n10923), .ZN(n16519) );
  NAND2_X1 U14175 ( .A1(n16519), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16517) );
  NAND2_X1 U14176 ( .A1(n16750), .A2(n16517), .ZN(n10924) );
  NAND2_X1 U14177 ( .A1(n16666), .A2(n10924), .ZN(n16507) );
  NAND2_X1 U14178 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11079) );
  INV_X1 U14179 ( .A(n11079), .ZN(n10925) );
  OAI21_X1 U14180 ( .B1(n17232), .B2(n10925), .A(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10926) );
  OR2_X1 U14181 ( .A1(n16507), .A2(n10926), .ZN(n16484) );
  NAND2_X1 U14182 ( .A1(n16484), .A2(n16671), .ZN(n16469) );
  AND2_X1 U14183 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16451) );
  OR2_X1 U14184 ( .A1(n16713), .A2(n16451), .ZN(n10927) );
  NAND2_X1 U14185 ( .A1(n16469), .A2(n10927), .ZN(n16443) );
  AND2_X1 U14186 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11427) );
  AOI21_X1 U14187 ( .B1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n11427), .A(
        n17232), .ZN(n10928) );
  NOR2_X1 U14188 ( .A1(n16443), .A2(n10928), .ZN(n11511) );
  OAI21_X1 U14189 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n17232), .A(
        n11511), .ZN(n10937) );
  INV_X2 U14190 ( .A(n19571), .ZN(n17200) );
  INV_X1 U14191 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n11403) );
  NOR2_X1 U14192 ( .A1(n17200), .A2(n11403), .ZN(n12260) );
  INV_X1 U14193 ( .A(n16515), .ZN(n16559) );
  NAND2_X1 U14194 ( .A1(n11127), .A2(n16749), .ZN(n10930) );
  AOI21_X1 U14195 ( .B1(n16559), .B2(n10930), .A(n10929), .ZN(n10931) );
  INV_X1 U14196 ( .A(n16673), .ZN(n10932) );
  NOR2_X1 U14197 ( .A1(n17214), .A2(n10932), .ZN(n16688) );
  AND2_X1 U14198 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11147) );
  NAND2_X1 U14199 ( .A1(n16688), .A2(n11147), .ZN(n16649) );
  INV_X1 U14200 ( .A(n16517), .ZN(n10933) );
  NAND2_X1 U14201 ( .A1(n10933), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10934) );
  NAND2_X1 U14202 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n10935) );
  NOR2_X1 U14203 ( .A1(n16494), .A2(n10935), .ZN(n16465) );
  NAND2_X1 U14204 ( .A1(n16439), .A2(n11427), .ZN(n16426) );
  INV_X1 U14205 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11512) );
  NOR4_X1 U14206 ( .A1(n16426), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n11512), .A4(n11484), .ZN(n10936) );
  AOI211_X1 U14207 ( .C1(n10937), .C2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n12260), .B(n10936), .ZN(n10938) );
  INV_X1 U14208 ( .A(n10939), .ZN(n11413) );
  NAND2_X1 U14209 ( .A1(n11406), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10950) );
  NAND2_X1 U14210 ( .A1(n20307), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10949) );
  INV_X1 U14211 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n10958) );
  NAND2_X1 U14212 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10957) );
  NAND2_X1 U14213 ( .A1(n10994), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n10956) );
  OAI211_X1 U14214 ( .C1(n11390), .C2(n10958), .A(n10957), .B(n10956), .ZN(
        n10959) );
  INV_X1 U14215 ( .A(n10941), .ZN(n10960) );
  NAND2_X1 U14216 ( .A1(n10940), .A2(n10960), .ZN(n10962) );
  AOI21_X1 U14217 ( .B1(n10962), .B2(n10961), .A(n13438), .ZN(n10969) );
  INV_X1 U14218 ( .A(n20307), .ZN(n10964) );
  NAND2_X1 U14219 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10963) );
  NAND2_X1 U14220 ( .A1(n10964), .A2(n10963), .ZN(n10965) );
  OAI211_X1 U14221 ( .C1(n11390), .C2(n19375), .A(n10967), .B(n10966), .ZN(
        n10968) );
  NOR2_X1 U14222 ( .A1(n10969), .A2(n10968), .ZN(n10972) );
  NAND2_X1 U14223 ( .A1(n10970), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10971) );
  NAND2_X1 U14224 ( .A1(n10972), .A2(n10971), .ZN(n11002) );
  AND3_X1 U14225 ( .A1(n10946), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n10356), 
        .ZN(n10973) );
  INV_X1 U14226 ( .A(n14214), .ZN(n10974) );
  AOI22_X1 U14227 ( .A1(n10974), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n20307), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n10975) );
  NAND2_X1 U14228 ( .A1(n10976), .A2(n10975), .ZN(n11003) );
  NAND2_X1 U14229 ( .A1(n10979), .A2(n10980), .ZN(n10982) );
  AOI21_X1 U14230 ( .B1(n13438), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10981) );
  INV_X1 U14231 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n15947) );
  INV_X1 U14232 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10983) );
  OAI22_X1 U14233 ( .A1(n11380), .A2(n15947), .B1(n10955), .B2(n10983), .ZN(
        n10984) );
  NAND2_X1 U14234 ( .A1(n10986), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10988) );
  NAND2_X1 U14235 ( .A1(n9608), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10989) );
  NAND2_X1 U14236 ( .A1(n11000), .A2(n11001), .ZN(n10990) );
  INV_X1 U14237 ( .A(n11000), .ZN(n10992) );
  INV_X1 U14238 ( .A(n11001), .ZN(n10991) );
  NAND2_X1 U14239 ( .A1(n10992), .A2(n10991), .ZN(n10993) );
  AOI22_X1 U14240 ( .A1(n10979), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n20307), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10998) );
  INV_X1 U14241 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n17201) );
  NAND2_X1 U14242 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10996) );
  NAND2_X1 U14243 ( .A1(n11400), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10995) );
  BUF_X2 U14244 ( .A(n11567), .Z(n14111) );
  NAND2_X2 U14245 ( .A1(n14111), .A2(n15952), .ZN(n11022) );
  INV_X1 U14246 ( .A(n11572), .ZN(n16746) );
  AND2_X2 U14247 ( .A1(n11012), .A2(n11023), .ZN(n11057) );
  AOI22_X1 U14248 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19605), .B1(
        n11052), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11010) );
  AND2_X2 U14249 ( .A1(n11026), .A2(n11015), .ZN(n19651) );
  AOI22_X1 U14250 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20128), .B1(
        n19880), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11020) );
  INV_X1 U14251 ( .A(n11015), .ZN(n11016) );
  INV_X1 U14252 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11017) );
  NOR2_X2 U14253 ( .A1(n11022), .A2(n11021), .ZN(n19814) );
  AND2_X2 U14254 ( .A1(n11026), .A2(n11023), .ZN(n19687) );
  AOI22_X1 U14255 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19814), .B1(
        n19687), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11030) );
  INV_X1 U14256 ( .A(n11024), .ZN(n11025) );
  INV_X1 U14257 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11027) );
  NOR2_X1 U14258 ( .A1(n11028), .A2(n11716), .ZN(n11029) );
  NAND3_X1 U14259 ( .A1(n11716), .A2(n17218), .A3(n11033), .ZN(n11039) );
  NAND2_X1 U14260 ( .A1(n11039), .A2(n11038), .ZN(n11037) );
  INV_X1 U14261 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n16726) );
  NAND2_X1 U14262 ( .A1(n16725), .A2(n16726), .ZN(n11046) );
  XNOR2_X1 U14263 ( .A(n17218), .B(n11033), .ZN(n11035) );
  INV_X1 U14264 ( .A(n11035), .ZN(n11034) );
  INV_X1 U14265 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n17217) );
  AOI21_X1 U14266 ( .B1(n11716), .B2(n17218), .A(n17217), .ZN(n17219) );
  NAND2_X1 U14267 ( .A1(n11034), .A2(n17219), .ZN(n11036) );
  XNOR2_X1 U14268 ( .A(n17219), .B(n11035), .ZN(n13640) );
  NAND2_X1 U14269 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13640), .ZN(
        n13639) );
  NAND2_X1 U14270 ( .A1(n11036), .A2(n13639), .ZN(n11040) );
  XOR2_X1 U14271 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n11040), .Z(
        n14614) );
  OAI21_X1 U14272 ( .B1(n11039), .B2(n11038), .A(n11037), .ZN(n14615) );
  NAND2_X1 U14273 ( .A1(n14614), .A2(n14615), .ZN(n11042) );
  NAND2_X1 U14274 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11040), .ZN(
        n11041) );
  NAND2_X1 U14275 ( .A1(n11042), .A2(n11041), .ZN(n11043) );
  INV_X1 U14276 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n17213) );
  XNOR2_X1 U14277 ( .A(n11043), .B(n17213), .ZN(n16415) );
  NAND2_X1 U14278 ( .A1(n11043), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11044) );
  NAND2_X1 U14279 ( .A1(n11046), .A2(n16724), .ZN(n11049) );
  INV_X1 U14280 ( .A(n16725), .ZN(n11047) );
  NAND2_X1 U14281 ( .A1(n11047), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11048) );
  XNOR2_X1 U14282 ( .A(n11051), .B(n11063), .ZN(n11067) );
  NAND2_X1 U14283 ( .A1(n11067), .A2(n11066), .ZN(n16710) );
  AOI22_X1 U14284 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19846), .B1(
        n19687), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11055) );
  AOI22_X1 U14285 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20128), .B1(
        n11052), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11054) );
  INV_X1 U14286 ( .A(n16811), .ZN(n16805) );
  AOI22_X1 U14287 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n16805), .B1(
        n19814), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11053) );
  INV_X1 U14288 ( .A(n20039), .ZN(n11056) );
  AOI22_X1 U14289 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19651), .B1(
        n11056), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11061) );
  AOI22_X1 U14290 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n16822), .B1(
        n19980), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11060) );
  AOI22_X1 U14291 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19605), .B1(
        n19918), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11059) );
  AOI22_X1 U14292 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n11057), .B1(
        n19740), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11058) );
  NAND2_X1 U14293 ( .A1(n11098), .A2(n11716), .ZN(n11062) );
  NAND2_X1 U14294 ( .A1(n11103), .A2(n11141), .ZN(n11064) );
  INV_X1 U14295 ( .A(n16711), .ZN(n11069) );
  NAND2_X1 U14296 ( .A1(n11069), .A2(n11141), .ZN(n11070) );
  INV_X1 U14297 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11074) );
  INV_X1 U14298 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11139) );
  OAI21_X1 U14299 ( .B1(n11075), .B2(n16378), .A(n11139), .ZN(n11077) );
  INV_X1 U14300 ( .A(n11075), .ZN(n11076) );
  NOR2_X1 U14301 ( .A1(n16517), .A2(n11079), .ZN(n11080) );
  INV_X1 U14302 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16438) );
  INV_X1 U14303 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11081) );
  INV_X1 U14304 ( .A(n12265), .ZN(n11082) );
  NAND2_X1 U14305 ( .A1(n11082), .A2(n17209), .ZN(n11412) );
  NOR2_X1 U14306 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n11085) );
  NAND2_X1 U14307 ( .A1(n11287), .A2(n11085), .ZN(n11086) );
  NAND2_X1 U14308 ( .A1(n11114), .A2(n11124), .ZN(n11110) );
  NAND2_X1 U14309 ( .A1(n11088), .A2(n9570), .ZN(n11119) );
  OR2_X1 U14310 ( .A1(n11119), .A2(n11089), .ZN(n11091) );
  NAND2_X1 U14311 ( .A1(n11287), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n11090) );
  OAI211_X1 U14312 ( .C1(n11116), .C2(n11092), .A(n11091), .B(n11090), .ZN(
        n11109) );
  NOR2_X1 U14313 ( .A1(n11116), .A2(n11093), .ZN(n11096) );
  INV_X1 U14314 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n19428) );
  OAI22_X1 U14315 ( .A1(n11119), .A2(n11094), .B1(n9571), .B2(n19428), .ZN(
        n11095) );
  INV_X1 U14316 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n14247) );
  MUX2_X1 U14317 ( .A(n14247), .B(n11142), .S(n9571), .Z(n11105) );
  INV_X1 U14318 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n14268) );
  INV_X1 U14319 ( .A(n11098), .ZN(n11099) );
  MUX2_X1 U14320 ( .A(n14268), .B(n11099), .S(n9571), .Z(n11100) );
  INV_X1 U14321 ( .A(n11100), .ZN(n11101) );
  NAND2_X1 U14322 ( .A1(n9669), .A2(n11101), .ZN(n11102) );
  NAND2_X1 U14323 ( .A1(n11135), .A2(n11102), .ZN(n15896) );
  NAND2_X1 U14324 ( .A1(n11104), .A2(n11097), .ZN(n11106) );
  NAND2_X1 U14325 ( .A1(n9669), .A2(n11106), .ZN(n15921) );
  XNOR2_X1 U14326 ( .A(n15921), .B(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16714) );
  INV_X1 U14327 ( .A(n9680), .ZN(n11112) );
  NAND2_X1 U14328 ( .A1(n11112), .A2(n11107), .ZN(n11108) );
  NAND2_X1 U14329 ( .A1(n11104), .A2(n11108), .ZN(n19406) );
  XNOR2_X1 U14330 ( .A(n19406), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n16729) );
  NAND2_X1 U14331 ( .A1(n11110), .A2(n11109), .ZN(n11111) );
  NAND2_X1 U14332 ( .A1(n11112), .A2(n11111), .ZN(n15935) );
  INV_X1 U14333 ( .A(n15935), .ZN(n11113) );
  NOR2_X1 U14334 ( .A1(n11113), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n16416) );
  XNOR2_X1 U14335 ( .A(n11114), .B(n11124), .ZN(n15938) );
  NOR2_X1 U14336 ( .A1(n15938), .A2(n11127), .ZN(n11128) );
  INV_X1 U14337 ( .A(n17218), .ZN(n11115) );
  NOR2_X1 U14338 ( .A1(n11116), .A2(n11115), .ZN(n11121) );
  INV_X1 U14339 ( .A(n11117), .ZN(n11118) );
  INV_X1 U14340 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n13994) );
  OAI22_X1 U14341 ( .A1(n11119), .A2(n11118), .B1(n13994), .B2(n9571), .ZN(
        n11120) );
  OR2_X1 U14342 ( .A1(n11121), .A2(n11120), .ZN(n17221) );
  AND2_X1 U14343 ( .A1(n17221), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17223) );
  NAND2_X1 U14344 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n11122) );
  NOR2_X1 U14345 ( .A1(n9571), .A2(n11122), .ZN(n11123) );
  NOR2_X1 U14346 ( .A1(n11124), .A2(n11123), .ZN(n15961) );
  AND2_X1 U14347 ( .A1(n17223), .A2(n15961), .ZN(n13641) );
  INV_X1 U14348 ( .A(n17223), .ZN(n11126) );
  INV_X1 U14349 ( .A(n15961), .ZN(n11125) );
  NAND2_X1 U14350 ( .A1(n11126), .A2(n11125), .ZN(n13642) );
  OAI21_X1 U14351 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13641), .A(
        n13642), .ZN(n14619) );
  XNOR2_X1 U14352 ( .A(n15938), .B(n11127), .ZN(n14620) );
  NOR2_X1 U14353 ( .A1(n14619), .A2(n14620), .ZN(n14618) );
  NOR2_X1 U14354 ( .A1(n11128), .A2(n14618), .ZN(n16419) );
  NOR2_X1 U14355 ( .A1(n15935), .A2(n17213), .ZN(n16417) );
  INV_X1 U14356 ( .A(n16417), .ZN(n11129) );
  OAI21_X1 U14357 ( .B1(n16416), .B2(n16419), .A(n11129), .ZN(n16730) );
  NAND2_X1 U14358 ( .A1(n16729), .A2(n16730), .ZN(n16728) );
  OAI21_X1 U14359 ( .B1(n19406), .B2(n16726), .A(n16728), .ZN(n16715) );
  NAND2_X1 U14360 ( .A1(n16714), .A2(n16715), .ZN(n11132) );
  INV_X1 U14361 ( .A(n15921), .ZN(n11130) );
  NAND2_X1 U14362 ( .A1(n11130), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11131) );
  NAND2_X1 U14363 ( .A1(n11132), .A2(n11131), .ZN(n16408) );
  MUX2_X1 U14364 ( .A(P2_EBX_REG_7__SCAN_IN), .B(n16378), .S(n9571), .Z(n11136) );
  XNOR2_X1 U14365 ( .A(n11135), .B(n11136), .ZN(n15884) );
  NAND2_X1 U14366 ( .A1(n15884), .A2(n11074), .ZN(n16396) );
  NAND2_X1 U14367 ( .A1(n15896), .A2(n11293), .ZN(n11133) );
  OAI211_X1 U14368 ( .C1(n16408), .C2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n16396), .B(n11133), .ZN(n11134) );
  INV_X1 U14369 ( .A(n11134), .ZN(n11140) );
  INV_X1 U14370 ( .A(n11136), .ZN(n11137) );
  NAND2_X1 U14371 ( .A1(n11287), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11138) );
  XNOR2_X1 U14372 ( .A(n11154), .B(n11138), .ZN(n15873) );
  NAND2_X1 U14373 ( .A1(n15873), .A2(n11293), .ZN(n11145) );
  NAND2_X1 U14374 ( .A1(n11145), .A2(n11139), .ZN(n16384) );
  INV_X1 U14375 ( .A(n11141), .ZN(n11143) );
  NAND4_X1 U14376 ( .A1(n16384), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        n16408), .A4(n16396), .ZN(n11151) );
  INV_X1 U14377 ( .A(n15884), .ZN(n11148) );
  NAND2_X1 U14378 ( .A1(n11148), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16395) );
  OR2_X1 U14379 ( .A1(n11145), .A2(n16395), .ZN(n11150) );
  NAND2_X1 U14380 ( .A1(n15873), .A2(n11146), .ZN(n16383) );
  NAND2_X1 U14381 ( .A1(n11148), .A2(n11147), .ZN(n11149) );
  AND4_X1 U14382 ( .A1(n11151), .A2(n11150), .A3(n16383), .A4(n11149), .ZN(
        n11152) );
  OR2_X1 U14383 ( .A1(n11154), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11155) );
  INV_X1 U14384 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n21360) );
  NOR2_X1 U14385 ( .A1(n9571), .A2(n21360), .ZN(n11156) );
  XNOR2_X1 U14386 ( .A(n11158), .B(n11156), .ZN(n15863) );
  NAND2_X1 U14387 ( .A1(n15863), .A2(n11293), .ZN(n11157) );
  INV_X1 U14388 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16665) );
  NAND2_X1 U14389 ( .A1(n11157), .A2(n16665), .ZN(n16365) );
  INV_X1 U14390 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n11320) );
  NOR2_X1 U14391 ( .A1(n9571), .A2(n11320), .ZN(n11159) );
  INV_X1 U14392 ( .A(n11260), .ZN(n11247) );
  AOI21_X1 U14393 ( .B1(n11160), .B2(n11159), .A(n11247), .ZN(n11162) );
  INV_X1 U14394 ( .A(n11166), .ZN(n11161) );
  AND2_X1 U14395 ( .A1(n11162), .A2(n11161), .ZN(n15845) );
  AOI21_X1 U14396 ( .B1(n15845), .B2(n11293), .A(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16354) );
  AND2_X1 U14397 ( .A1(n11293), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11163) );
  NAND2_X1 U14398 ( .A1(n15845), .A2(n11163), .ZN(n16355) );
  AND2_X1 U14399 ( .A1(n11293), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11164) );
  NAND2_X1 U14400 ( .A1(n15863), .A2(n11164), .ZN(n16364) );
  AND2_X1 U14401 ( .A1(n16355), .A2(n16364), .ZN(n11165) );
  INV_X1 U14402 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16627) );
  NAND2_X1 U14403 ( .A1(n11287), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n11168) );
  INV_X1 U14404 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n16064) );
  NAND2_X1 U14405 ( .A1(n11199), .A2(n11260), .ZN(n11171) );
  INV_X1 U14406 ( .A(n11171), .ZN(n11167) );
  OAI21_X1 U14407 ( .B1(n11166), .B2(n11168), .A(n11167), .ZN(n15831) );
  NOR2_X1 U14408 ( .A1(n15831), .A2(n16378), .ZN(n16340) );
  INV_X1 U14409 ( .A(n16340), .ZN(n11169) );
  NAND2_X1 U14410 ( .A1(n11287), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11197) );
  INV_X1 U14411 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n11172) );
  NOR2_X1 U14412 ( .A1(P2_EBX_REG_15__SCAN_IN), .A2(P2_EBX_REG_14__SCAN_IN), 
        .ZN(n11174) );
  NOR2_X1 U14413 ( .A1(n9571), .A2(n11174), .ZN(n11175) );
  NOR2_X1 U14414 ( .A1(P2_EBX_REG_17__SCAN_IN), .A2(P2_EBX_REG_16__SCAN_IN), 
        .ZN(n11176) );
  INV_X1 U14415 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n16037) );
  NAND2_X1 U14416 ( .A1(n11181), .A2(n16037), .ZN(n11183) );
  AND2_X1 U14417 ( .A1(n11287), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n11177) );
  NAND2_X1 U14418 ( .A1(n11183), .A2(n11177), .ZN(n11179) );
  NOR2_X1 U14419 ( .A1(P2_EBX_REG_19__SCAN_IN), .A2(P2_EBX_REG_18__SCAN_IN), 
        .ZN(n11178) );
  INV_X1 U14420 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11535) );
  NAND2_X1 U14421 ( .A1(n11230), .A2(n11535), .ZN(n11538) );
  OR2_X1 U14422 ( .A1(n11181), .A2(n16037), .ZN(n11182) );
  INV_X1 U14423 ( .A(n11181), .ZN(n11204) );
  MUX2_X1 U14424 ( .A(n11182), .B(n11204), .S(n9571), .Z(n11184) );
  NAND2_X1 U14425 ( .A1(n11184), .A2(n11183), .ZN(n11231) );
  INV_X1 U14426 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16548) );
  AND2_X1 U14427 ( .A1(n11538), .A2(n11536), .ZN(n11466) );
  NAND2_X1 U14428 ( .A1(n11287), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11185) );
  XNOR2_X1 U14429 ( .A(n9630), .B(n11185), .ZN(n15731) );
  NAND2_X1 U14430 ( .A1(n15731), .A2(n11293), .ZN(n11227) );
  INV_X1 U14431 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11226) );
  NAND2_X1 U14432 ( .A1(n11227), .A2(n11226), .ZN(n11458) );
  NAND2_X1 U14433 ( .A1(n11466), .A2(n11458), .ZN(n16266) );
  INV_X1 U14434 ( .A(n16266), .ZN(n11216) );
  INV_X1 U14435 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n11186) );
  NOR2_X1 U14436 ( .A1(n9571), .A2(n11186), .ZN(n11187) );
  AOI21_X1 U14437 ( .B1(n11192), .B2(n11187), .A(n11247), .ZN(n11188) );
  OR2_X1 U14438 ( .A1(n11192), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11203) );
  NAND2_X1 U14439 ( .A1(n15792), .A2(n11293), .ZN(n11189) );
  XNOR2_X1 U14440 ( .A(n11189), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16290) );
  OR2_X1 U14441 ( .A1(n11190), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11207) );
  INV_X1 U14442 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n19391) );
  NOR2_X1 U14443 ( .A1(n9571), .A2(n19391), .ZN(n11191) );
  NAND2_X1 U14444 ( .A1(n11207), .A2(n11191), .ZN(n11193) );
  NAND2_X1 U14445 ( .A1(n11193), .A2(n11192), .ZN(n19396) );
  INV_X1 U14446 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16590) );
  NAND2_X1 U14447 ( .A1(n11194), .A2(n16590), .ZN(n16301) );
  XNOR2_X1 U14448 ( .A(n11195), .B(n10408), .ZN(n13582) );
  NAND2_X1 U14449 ( .A1(n13582), .A2(n11293), .ZN(n11196) );
  INV_X1 U14450 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11224) );
  NAND2_X1 U14451 ( .A1(n11196), .A2(n11224), .ZN(n16321) );
  INV_X1 U14452 ( .A(n11197), .ZN(n11198) );
  NAND2_X1 U14453 ( .A1(n11199), .A2(n11198), .ZN(n11200) );
  NAND2_X1 U14454 ( .A1(n11195), .A2(n11200), .ZN(n15821) );
  OR2_X1 U14455 ( .A1(n15821), .A2(n16378), .ZN(n11201) );
  NAND2_X1 U14456 ( .A1(n11201), .A2(n16627), .ZN(n16331) );
  AND3_X1 U14457 ( .A1(n16301), .A2(n16321), .A3(n16331), .ZN(n11210) );
  INV_X1 U14458 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n11346) );
  NOR2_X1 U14459 ( .A1(n10838), .A2(n11346), .ZN(n11202) );
  NAND2_X1 U14460 ( .A1(n11203), .A2(n11202), .ZN(n11205) );
  NAND2_X1 U14461 ( .A1(n11205), .A2(n11204), .ZN(n11220) );
  INV_X1 U14462 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16574) );
  OAI21_X1 U14463 ( .B1(n11220), .B2(n16378), .A(n16574), .ZN(n11463) );
  NAND2_X1 U14464 ( .A1(n11190), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11206) );
  MUX2_X1 U14465 ( .A(n11190), .B(n11206), .S(n11287), .Z(n11208) );
  NAND2_X1 U14466 ( .A1(n11208), .A2(n11207), .ZN(n15806) );
  OR2_X1 U14467 ( .A1(n15806), .A2(n16378), .ZN(n11209) );
  INV_X1 U14468 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16601) );
  NAND2_X1 U14469 ( .A1(n11209), .A2(n16601), .ZN(n16312) );
  INV_X1 U14470 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n11211) );
  INV_X1 U14471 ( .A(n11235), .ZN(n11214) );
  NAND3_X1 U14472 ( .A1(n11212), .A2(P2_EBX_REG_21__SCAN_IN), .A3(n11287), 
        .ZN(n11213) );
  INV_X1 U14473 ( .A(n16270), .ZN(n11215) );
  AND2_X1 U14474 ( .A1(n11293), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11219) );
  NAND2_X1 U14475 ( .A1(n15710), .A2(n11219), .ZN(n16268) );
  INV_X1 U14476 ( .A(n11220), .ZN(n15773) );
  AND2_X1 U14477 ( .A1(n11293), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11221) );
  NAND2_X1 U14478 ( .A1(n15773), .A2(n11221), .ZN(n11462) );
  AND2_X1 U14479 ( .A1(n11293), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11222) );
  NAND2_X1 U14480 ( .A1(n15792), .A2(n11222), .ZN(n11496) );
  NAND2_X1 U14481 ( .A1(n11293), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11223) );
  OR2_X1 U14482 ( .A1(n19396), .A2(n11223), .ZN(n16300) );
  INV_X1 U14483 ( .A(n13582), .ZN(n11225) );
  OR3_X1 U14484 ( .A1(n11225), .A2(n16378), .A3(n11224), .ZN(n16320) );
  AND4_X1 U14485 ( .A1(n11462), .A2(n11496), .A3(n16300), .A4(n16320), .ZN(
        n11229) );
  OR2_X1 U14486 ( .A1(n11227), .A2(n11226), .ZN(n16265) );
  NAND2_X1 U14487 ( .A1(n11293), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11228) );
  OR2_X1 U14488 ( .A1(n15806), .A2(n11228), .ZN(n16311) );
  NAND4_X1 U14489 ( .A1(n16268), .A2(n11229), .A3(n16265), .A4(n16311), .ZN(
        n11233) );
  OR2_X1 U14490 ( .A1(n11230), .A2(n11535), .ZN(n11539) );
  INV_X1 U14491 ( .A(n11231), .ZN(n15758) );
  AND2_X1 U14492 ( .A1(n11293), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11232) );
  NAND2_X1 U14493 ( .A1(n15758), .A2(n11232), .ZN(n16282) );
  NAND2_X1 U14494 ( .A1(n11539), .A2(n16282), .ZN(n11464) );
  NAND2_X1 U14495 ( .A1(n11287), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11236) );
  INV_X1 U14496 ( .A(n11236), .ZN(n11237) );
  NAND2_X1 U14497 ( .A1(n9936), .A2(n11237), .ZN(n11238) );
  NAND2_X1 U14498 ( .A1(n11245), .A2(n11238), .ZN(n15695) );
  NOR2_X1 U14499 ( .A1(n15695), .A2(n16378), .ZN(n11239) );
  NAND2_X1 U14500 ( .A1(n11239), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16253) );
  NAND2_X1 U14501 ( .A1(n11287), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11243) );
  XNOR2_X1 U14502 ( .A(n11245), .B(n11243), .ZN(n15682) );
  NAND2_X1 U14503 ( .A1(n15682), .A2(n11293), .ZN(n11240) );
  XNOR2_X1 U14504 ( .A(n11240), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16248) );
  INV_X1 U14505 ( .A(n11240), .ZN(n11241) );
  INV_X1 U14506 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16481) );
  INV_X1 U14507 ( .A(n11243), .ZN(n11244) );
  INV_X1 U14508 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n16010) );
  INV_X1 U14509 ( .A(n11246), .ZN(n11249) );
  NOR2_X1 U14510 ( .A1(n9571), .A2(n16010), .ZN(n11248) );
  AOI21_X1 U14511 ( .B1(n11249), .B2(n11248), .A(n11247), .ZN(n11250) );
  NAND2_X1 U14512 ( .A1(n11258), .A2(n11250), .ZN(n15672) );
  OR2_X1 U14513 ( .A1(n15672), .A2(n16378), .ZN(n11251) );
  INV_X1 U14514 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16480) );
  NAND2_X1 U14515 ( .A1(n11251), .A2(n16480), .ZN(n16236) );
  NAND2_X1 U14516 ( .A1(n11265), .A2(n11260), .ZN(n11264) );
  INV_X1 U14517 ( .A(n11264), .ZN(n11291) );
  NAND3_X1 U14518 ( .A1(n11261), .A2(P2_EBX_REG_26__SCAN_IN), .A3(n11287), 
        .ZN(n11254) );
  INV_X1 U14519 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16456) );
  OAI21_X1 U14520 ( .B1(n15643), .B2(n16378), .A(n16456), .ZN(n11257) );
  INV_X1 U14521 ( .A(n15643), .ZN(n11256) );
  AND2_X1 U14522 ( .A1(n11293), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11255) );
  NAND2_X1 U14523 ( .A1(n11256), .A2(n11255), .ZN(n11272) );
  NAND2_X1 U14524 ( .A1(n11257), .A2(n11272), .ZN(n16216) );
  INV_X1 U14525 ( .A(n16216), .ZN(n11262) );
  NAND3_X1 U14526 ( .A1(n11261), .A2(n11260), .A3(n11259), .ZN(n15655) );
  INV_X1 U14527 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16468) );
  NAND2_X1 U14528 ( .A1(n11287), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11266) );
  NAND2_X1 U14529 ( .A1(n11264), .A2(n11266), .ZN(n11279) );
  NAND2_X1 U14530 ( .A1(n11287), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11280) );
  XNOR2_X1 U14531 ( .A(n11279), .B(n11280), .ZN(n15609) );
  NAND2_X1 U14532 ( .A1(n15609), .A2(n11293), .ZN(n11275) );
  INV_X1 U14533 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11274) );
  NAND2_X1 U14534 ( .A1(n11275), .A2(n11274), .ZN(n11416) );
  INV_X1 U14535 ( .A(n11266), .ZN(n11267) );
  NAND2_X1 U14536 ( .A1(n11265), .A2(n11267), .ZN(n11268) );
  NAND2_X1 U14537 ( .A1(n11279), .A2(n11268), .ZN(n15626) );
  INV_X1 U14538 ( .A(n11275), .ZN(n11273) );
  INV_X1 U14539 ( .A(n11270), .ZN(n11271) );
  NAND2_X1 U14540 ( .A1(n11271), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16225) );
  NAND2_X1 U14541 ( .A1(n11272), .A2(n16225), .ZN(n11414) );
  AOI21_X1 U14542 ( .B1(n11273), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n11414), .ZN(n11276) );
  INV_X1 U14543 ( .A(n11279), .ZN(n11281) );
  NAND2_X1 U14544 ( .A1(n11281), .A2(n11280), .ZN(n11283) );
  INV_X1 U14545 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n11282) );
  NOR2_X1 U14546 ( .A1(n9571), .A2(n11282), .ZN(n11284) );
  XNOR2_X1 U14547 ( .A(n11283), .B(n11284), .ZN(n11289) );
  OAI21_X1 U14548 ( .B1(n11289), .B2(n16378), .A(n11512), .ZN(n11449) );
  INV_X1 U14549 ( .A(n11283), .ZN(n11286) );
  INV_X1 U14550 ( .A(n11284), .ZN(n11285) );
  NAND2_X1 U14551 ( .A1(n11286), .A2(n11285), .ZN(n11290) );
  NAND2_X1 U14552 ( .A1(n11287), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11288) );
  XNOR2_X1 U14553 ( .A(n11290), .B(n11288), .ZN(n14601) );
  AOI21_X1 U14554 ( .B1(n14601), .B2(n11293), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11487) );
  INV_X1 U14555 ( .A(n11289), .ZN(n15606) );
  NAND3_X1 U14556 ( .A1(n15606), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n11293), .ZN(n11485) );
  NOR2_X1 U14557 ( .A1(n11290), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11292) );
  MUX2_X1 U14558 ( .A(n11292), .B(n11291), .S(n10838), .Z(n13493) );
  NAND2_X1 U14559 ( .A1(n13493), .A2(n11293), .ZN(n11294) );
  XOR2_X1 U14560 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n11294), .Z(
        n11295) );
  AND2_X1 U14561 ( .A1(n16854), .A2(n10356), .ZN(n20298) );
  NAND2_X1 U14562 ( .A1(n12264), .A2(n17224), .ZN(n11411) );
  INV_X1 U14563 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n11300) );
  NAND2_X1 U14564 ( .A1(n11400), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n11299) );
  NAND2_X1 U14565 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11298) );
  AOI21_X1 U14566 ( .B1(n11399), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n11301), .ZN(n16731) );
  INV_X1 U14567 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n15920) );
  NAND2_X1 U14568 ( .A1(n11400), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n11305) );
  NAND2_X1 U14569 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11304) );
  OAI211_X1 U14570 ( .C1(n11390), .C2(n15920), .A(n11305), .B(n11304), .ZN(
        n11306) );
  AOI21_X1 U14571 ( .B1(n11399), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n11306), .ZN(n14246) );
  NOR2_X2 U14572 ( .A1(n14243), .A2(n14246), .ZN(n14244) );
  NAND2_X1 U14573 ( .A1(n11399), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11309) );
  OAI22_X1 U14574 ( .A1(n11380), .A2(n14268), .B1(n10955), .B2(n10112), .ZN(
        n11307) );
  AOI21_X1 U14575 ( .B1(n11392), .B2(P2_REIP_REG_6__SCAN_IN), .A(n11307), .ZN(
        n11308) );
  NAND2_X1 U14576 ( .A1(n11309), .A2(n11308), .ZN(n14267) );
  NAND2_X1 U14577 ( .A1(n14244), .A2(n14267), .ZN(n14266) );
  INV_X1 U14578 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n20217) );
  NAND2_X1 U14579 ( .A1(n11400), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n11311) );
  NAND2_X1 U14580 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11310) );
  AOI21_X1 U14581 ( .B1(n11399), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n11312), .ZN(n14289) );
  INV_X1 U14582 ( .A(n14289), .ZN(n11313) );
  INV_X1 U14583 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n20219) );
  NAND2_X1 U14584 ( .A1(n11400), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11315) );
  NAND2_X1 U14585 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11314) );
  OAI211_X1 U14586 ( .C1(n11390), .C2(n20219), .A(n11315), .B(n11314), .ZN(
        n11316) );
  AOI21_X1 U14587 ( .B1(n11399), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n11316), .ZN(n14321) );
  NAND2_X1 U14588 ( .A1(n11399), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11319) );
  OAI22_X1 U14589 ( .A1(n11380), .A2(n21360), .B1(n10955), .B2(n16368), .ZN(
        n11317) );
  AOI21_X1 U14590 ( .B1(n11392), .B2(P2_REIP_REG_9__SCAN_IN), .A(n11317), .ZN(
        n11318) );
  NAND2_X1 U14591 ( .A1(n11319), .A2(n11318), .ZN(n14331) );
  NAND2_X1 U14592 ( .A1(n11399), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11323) );
  INV_X1 U14593 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n15853) );
  OAI22_X1 U14594 ( .A1(n11380), .A2(n11320), .B1(n10955), .B2(n15853), .ZN(
        n11321) );
  AOI21_X1 U14595 ( .B1(n11392), .B2(P2_REIP_REG_10__SCAN_IN), .A(n11321), 
        .ZN(n11322) );
  NAND2_X1 U14596 ( .A1(n11323), .A2(n11322), .ZN(n15842) );
  NAND2_X1 U14597 ( .A1(n14330), .A2(n15842), .ZN(n15825) );
  INV_X1 U14598 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n16343) );
  NAND2_X1 U14599 ( .A1(n11400), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n11325) );
  NAND2_X1 U14600 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11324) );
  AOI21_X1 U14601 ( .B1(n11399), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n11326), .ZN(n15826) );
  NAND2_X1 U14602 ( .A1(n11400), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11329) );
  NAND2_X1 U14603 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11328) );
  AOI21_X1 U14604 ( .B1(n11399), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n11330), .ZN(n15812) );
  INV_X1 U14605 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n20228) );
  NAND2_X1 U14606 ( .A1(n11400), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11333) );
  NAND2_X1 U14607 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11332) );
  OAI211_X1 U14608 ( .C1(n11390), .C2(n20228), .A(n11333), .B(n11332), .ZN(
        n11334) );
  AOI21_X1 U14609 ( .B1(n11399), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n11334), .ZN(n13585) );
  NAND2_X1 U14610 ( .A1(n11399), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11337) );
  INV_X1 U14611 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n15803) );
  OAI22_X1 U14612 ( .A1(n11380), .A2(n15803), .B1(n10955), .B2(n10110), .ZN(
        n11335) );
  AOI21_X1 U14613 ( .B1(n11392), .B2(P2_REIP_REG_14__SCAN_IN), .A(n11335), 
        .ZN(n11336) );
  NAND2_X1 U14614 ( .A1(n11337), .A2(n11336), .ZN(n14423) );
  NAND2_X1 U14615 ( .A1(n13584), .A2(n14423), .ZN(n14422) );
  INV_X1 U14616 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n11340) );
  NAND2_X1 U14617 ( .A1(n11400), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11339) );
  NAND2_X1 U14618 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11338) );
  AOI21_X1 U14619 ( .B1(n11399), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n11341), .ZN(n16049) );
  INV_X1 U14620 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n20233) );
  NAND2_X1 U14621 ( .A1(n11400), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11343) );
  NAND2_X1 U14622 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11342) );
  AOI21_X1 U14623 ( .B1(n11399), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n11344), .ZN(n15783) );
  NAND2_X1 U14624 ( .A1(n11399), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11349) );
  INV_X1 U14625 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11504) );
  OAI22_X1 U14626 ( .A1(n11380), .A2(n11346), .B1(n10955), .B2(n11504), .ZN(
        n11347) );
  AOI21_X1 U14627 ( .B1(n11392), .B2(P2_REIP_REG_17__SCAN_IN), .A(n11347), 
        .ZN(n11348) );
  NAND2_X1 U14628 ( .A1(n11349), .A2(n11348), .ZN(n11503) );
  NAND2_X1 U14629 ( .A1(n11399), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11352) );
  OAI22_X1 U14630 ( .A1(n11380), .A2(n16037), .B1(n10955), .B2(n10118), .ZN(
        n11350) );
  AOI21_X1 U14631 ( .B1(n11392), .B2(P2_REIP_REG_18__SCAN_IN), .A(n11350), 
        .ZN(n11351) );
  NAND2_X1 U14632 ( .A1(n11352), .A2(n11351), .ZN(n15749) );
  INV_X1 U14633 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n20239) );
  NAND2_X1 U14634 ( .A1(n11400), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n11354) );
  NAND2_X1 U14635 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n11353) );
  OAI211_X1 U14636 ( .C1(n11390), .C2(n20239), .A(n11354), .B(n11353), .ZN(
        n11355) );
  AOI21_X1 U14637 ( .B1(n11399), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n11355), .ZN(n11544) );
  INV_X1 U14638 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n20241) );
  NAND2_X1 U14639 ( .A1(n11400), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11357) );
  NAND2_X1 U14640 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11356) );
  AOI21_X1 U14641 ( .B1(n11399), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n11358), .ZN(n11470) );
  INV_X1 U14642 ( .A(n11470), .ZN(n11359) );
  AND2_X2 U14643 ( .A1(n11467), .A2(n11359), .ZN(n11468) );
  NAND2_X1 U14644 ( .A1(n11399), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11362) );
  INV_X1 U14645 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n16274) );
  OAI22_X1 U14646 ( .A1(n11380), .A2(n9935), .B1(n10955), .B2(n16274), .ZN(
        n11360) );
  AOI21_X1 U14647 ( .B1(n11392), .B2(P2_REIP_REG_21__SCAN_IN), .A(n11360), 
        .ZN(n11361) );
  NAND2_X1 U14648 ( .A1(n11362), .A2(n11361), .ZN(n15706) );
  NAND2_X1 U14649 ( .A1(n11399), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11366) );
  INV_X1 U14650 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n15696) );
  INV_X1 U14651 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11363) );
  OAI22_X1 U14652 ( .A1(n11380), .A2(n15696), .B1(n10955), .B2(n11363), .ZN(
        n11364) );
  AOI21_X1 U14653 ( .B1(n11392), .B2(P2_REIP_REG_22__SCAN_IN), .A(n11364), 
        .ZN(n11365) );
  NAND2_X1 U14654 ( .A1(n11366), .A2(n11365), .ZN(n15688) );
  INV_X1 U14655 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n11369) );
  NAND2_X1 U14656 ( .A1(n11400), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11368) );
  NAND2_X1 U14657 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n11367) );
  AOI21_X1 U14658 ( .B1(n11399), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n11370), .ZN(n15675) );
  INV_X1 U14659 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n20248) );
  NAND2_X1 U14660 ( .A1(n11400), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n11373) );
  NAND2_X1 U14661 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n11372) );
  OAI211_X1 U14662 ( .C1(n11390), .C2(n20248), .A(n11373), .B(n11372), .ZN(
        n11374) );
  AOI21_X1 U14663 ( .B1(n11399), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n11374), .ZN(n15661) );
  NOR2_X2 U14664 ( .A1(n15676), .A2(n15661), .ZN(n15649) );
  INV_X1 U14665 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n11377) );
  NAND2_X1 U14666 ( .A1(n11400), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n11376) );
  NAND2_X1 U14667 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11375) );
  AOI21_X1 U14668 ( .B1(n11399), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n11378), .ZN(n15651) );
  INV_X1 U14669 ( .A(n15651), .ZN(n11379) );
  NAND2_X1 U14670 ( .A1(n11399), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11383) );
  INV_X1 U14671 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16218) );
  OAI22_X1 U14672 ( .A1(n11380), .A2(n11252), .B1(n10955), .B2(n16218), .ZN(
        n11381) );
  AOI21_X1 U14673 ( .B1(n11392), .B2(P2_REIP_REG_26__SCAN_IN), .A(n11381), 
        .ZN(n11382) );
  NAND2_X1 U14674 ( .A1(n11383), .A2(n11382), .ZN(n15633) );
  INV_X1 U14675 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n11386) );
  NAND2_X1 U14676 ( .A1(n11400), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11385) );
  NAND2_X1 U14677 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n11384) );
  AOI21_X1 U14678 ( .B1(n11399), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n11387), .ZN(n15622) );
  INV_X1 U14679 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n20254) );
  NAND2_X1 U14680 ( .A1(n11400), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11389) );
  NAND2_X1 U14681 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11388) );
  OAI211_X1 U14682 ( .C1(n11390), .C2(n20254), .A(n11389), .B(n11388), .ZN(
        n11391) );
  AOI21_X1 U14683 ( .B1(n11399), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n11391), .ZN(n11422) );
  AOI22_X1 U14684 ( .A1(n11400), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n11394) );
  NAND2_X1 U14685 ( .A1(n11392), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11393) );
  OAI211_X1 U14686 ( .C1(n11395), .C2(n11512), .A(n11394), .B(n11393), .ZN(
        n11445) );
  INV_X1 U14687 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n11480) );
  NAND2_X1 U14688 ( .A1(n11400), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11397) );
  NAND2_X1 U14689 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n11396) );
  AOI21_X1 U14690 ( .B1(n11399), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n11398), .ZN(n11478) );
  NAND2_X1 U14691 ( .A1(n11399), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11402) );
  AOI22_X1 U14692 ( .A1(n11400), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n11401) );
  INV_X1 U14693 ( .A(n11406), .ZN(n16765) );
  INV_X1 U14694 ( .A(n16765), .ZN(n16787) );
  NAND2_X1 U14695 ( .A1(n16787), .A2(n11716), .ZN(n11407) );
  NAND2_X1 U14696 ( .A1(n11407), .A2(n14214), .ZN(n11408) );
  NAND4_X1 U14697 ( .A1(n11413), .A2(n11412), .A3(n11411), .A4(n11410), .ZN(
        P2_U3015) );
  NAND2_X1 U14698 ( .A1(n11524), .A2(n17224), .ZN(n11439) );
  OAI21_X1 U14699 ( .B1(n11418), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n11419), .ZN(n11531) );
  NAND2_X1 U14700 ( .A1(n10319), .A2(n11422), .ZN(n11424) );
  INV_X1 U14701 ( .A(n11446), .ZN(n11423) );
  NOR2_X1 U14702 ( .A1(n11525), .A2(n17227), .ZN(n11436) );
  INV_X1 U14703 ( .A(n11427), .ZN(n11428) );
  AND2_X1 U14704 ( .A1(n16439), .A2(n11428), .ZN(n11429) );
  OR2_X1 U14705 ( .A1(n16443), .A2(n11429), .ZN(n16428) );
  INV_X1 U14706 ( .A(n16428), .ZN(n11431) );
  AOI21_X1 U14707 ( .B1(n16439), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11430) );
  NAND2_X1 U14708 ( .A1(n19571), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11528) );
  OAI21_X1 U14709 ( .B1(n11431), .B2(n11430), .A(n11528), .ZN(n11432) );
  INV_X1 U14710 ( .A(n11432), .ZN(n11433) );
  NAND3_X1 U14711 ( .A1(n11439), .A2(n11438), .A3(n11437), .ZN(P2_U3018) );
  NAND2_X1 U14712 ( .A1(n20298), .A2(n11440), .ZN(n11441) );
  NAND2_X1 U14713 ( .A1(n11442), .A2(n11441), .ZN(n11443) );
  NOR2_X1 U14714 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20273) );
  OR2_X1 U14715 ( .A1(n20305), .A2(n20273), .ZN(n20276) );
  NAND2_X1 U14716 ( .A1(n20276), .A2(n13438), .ZN(n11444) );
  AND2_X1 U14717 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n16755) );
  OR2_X1 U14718 ( .A1(n11446), .A2(n11445), .ZN(n11447) );
  NOR2_X1 U14719 ( .A1(n19573), .A2(n15599), .ZN(n11448) );
  INV_X1 U14720 ( .A(n13624), .ZN(n11451) );
  NAND2_X1 U14721 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n13448), .ZN(
        n13447) );
  NAND2_X1 U14722 ( .A1(n13443), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13455) );
  NAND2_X1 U14723 ( .A1(n13464), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13466) );
  INV_X1 U14724 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n11452) );
  NAND2_X1 U14725 ( .A1(n13467), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13469) );
  INV_X1 U14726 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15654) );
  INV_X1 U14727 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n21293) );
  AND2_X1 U14728 ( .A1(n11526), .A2(n21293), .ZN(n11453) );
  NOR2_X1 U14729 ( .A1(n9745), .A2(n11453), .ZN(n15600) );
  NAND2_X1 U14730 ( .A1(n13438), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13712) );
  NAND2_X1 U14731 ( .A1(n20272), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13483) );
  NAND2_X1 U14732 ( .A1(n13712), .A2(n13483), .ZN(n19583) );
  NAND2_X1 U14733 ( .A1(n19571), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n16425) );
  OAI21_X1 U14734 ( .B1(n17198), .B2(n21293), .A(n16425), .ZN(n11454) );
  NAND2_X1 U14735 ( .A1(n16433), .A2(n19577), .ZN(n11457) );
  NOR3_X1 U14736 ( .A1(n15821), .A2(n16378), .A3(n16627), .ZN(n16333) );
  INV_X1 U14737 ( .A(n16321), .ZN(n11460) );
  INV_X1 U14738 ( .A(n16311), .ZN(n11461) );
  AND2_X1 U14739 ( .A1(n11463), .A2(n11462), .ZN(n11498) );
  INV_X1 U14740 ( .A(n11464), .ZN(n11465) );
  OAI21_X1 U14741 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n11864), .A(
        n13463), .ZN(n15725) );
  INV_X1 U14742 ( .A(n11467), .ZN(n11546) );
  AOI21_X1 U14743 ( .B1(n11470), .B2(n11546), .A(n11469), .ZN(n16533) );
  NAND2_X1 U14744 ( .A1(n16533), .A2(n19592), .ZN(n11472) );
  NOR2_X1 U14745 ( .A1(n17200), .A2(n20241), .ZN(n16537) );
  AOI21_X1 U14746 ( .B1(n19584), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16537), .ZN(n11471) );
  OAI211_X1 U14747 ( .C1(n15725), .C2(n19582), .A(n11472), .B(n11471), .ZN(
        n11473) );
  AOI21_X1 U14748 ( .B1(n10417), .B2(n9627), .A(n11473), .ZN(n11477) );
  INV_X1 U14749 ( .A(n16637), .ZN(n11552) );
  INV_X1 U14750 ( .A(n11549), .ZN(n11554) );
  NOR2_X2 U14751 ( .A1(n16280), .A2(n11535), .ZN(n11534) );
  NAND2_X1 U14752 ( .A1(n11476), .A2(n16519), .ZN(n16273) );
  OAI21_X1 U14753 ( .B1(n11534), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n16273), .ZN(n16544) );
  NAND2_X1 U14754 ( .A1(n11477), .A2(n10421), .ZN(P2_U2994) );
  NOR2_X1 U14755 ( .A1(n17200), .A2(n11480), .ZN(n11514) );
  XNOR2_X1 U14756 ( .A(n9745), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14602) );
  NOR2_X1 U14757 ( .A1(n19582), .A2(n14602), .ZN(n11481) );
  AOI211_X1 U14758 ( .C1(n19584), .C2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n11514), .B(n11481), .ZN(n11482) );
  OAI21_X1 U14759 ( .B1(n11859), .B2(n19573), .A(n11482), .ZN(n11483) );
  INV_X1 U14760 ( .A(n11483), .ZN(n11494) );
  XNOR2_X1 U14761 ( .A(n11456), .B(n11484), .ZN(n11519) );
  NAND2_X1 U14762 ( .A1(n11486), .A2(n11485), .ZN(n11491) );
  INV_X1 U14763 ( .A(n11487), .ZN(n11489) );
  NAND2_X1 U14764 ( .A1(n11489), .A2(n11488), .ZN(n11490) );
  XNOR2_X1 U14765 ( .A(n11491), .B(n11490), .ZN(n11520) );
  NAND3_X1 U14766 ( .A1(n11494), .A2(n11493), .A3(n11492), .ZN(P2_U2984) );
  AOI211_X1 U14767 ( .C1(n16574), .C2(n16558), .A(n19590), .B(n16281), .ZN(
        n11510) );
  AND2_X1 U14768 ( .A1(n11495), .A2(n11496), .ZN(n11499) );
  OAI21_X1 U14769 ( .B1(n11499), .B2(n11498), .A(n11497), .ZN(n16568) );
  INV_X1 U14770 ( .A(n11501), .ZN(n11502) );
  OAI21_X1 U14771 ( .B1(n11500), .B2(n11503), .A(n11502), .ZN(n16566) );
  AOI21_X1 U14772 ( .B1(n11504), .B2(n9658), .A(n13462), .ZN(n15767) );
  NAND2_X1 U14773 ( .A1(n19571), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n16565) );
  OAI21_X1 U14774 ( .B1(n17198), .B2(n11504), .A(n16565), .ZN(n11505) );
  AOI21_X1 U14775 ( .B1(n15767), .B2(n17192), .A(n11505), .ZN(n11506) );
  OAI21_X1 U14776 ( .B1(n16566), .B2(n19573), .A(n11506), .ZN(n11507) );
  INV_X1 U14777 ( .A(n11508), .ZN(n11509) );
  INV_X1 U14778 ( .A(n11511), .ZN(n11515) );
  NOR3_X1 U14779 ( .A1(n16426), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n11512), .ZN(n11513) );
  AOI211_X1 U14780 ( .C1(n11515), .C2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n11514), .B(n11513), .ZN(n11517) );
  NAND2_X1 U14781 ( .A1(n14612), .A2(n17215), .ZN(n11516) );
  OAI211_X1 U14782 ( .C1(n11859), .C2(n17227), .A(n11517), .B(n11516), .ZN(
        n11518) );
  INV_X1 U14783 ( .A(n11518), .ZN(n11523) );
  NAND2_X1 U14784 ( .A1(n11520), .A2(n17224), .ZN(n11521) );
  NAND3_X1 U14785 ( .A1(n11523), .A2(n11522), .A3(n11521), .ZN(P2_U3016) );
  NAND2_X1 U14786 ( .A1(n11524), .A2(n9627), .ZN(n11533) );
  INV_X1 U14787 ( .A(n11525), .ZN(n11530) );
  OAI21_X1 U14788 ( .B1(n13478), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n11526), .ZN(n15615) );
  NAND2_X1 U14789 ( .A1(n19584), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11527) );
  OAI211_X1 U14790 ( .C1(n19582), .C2(n15615), .A(n11528), .B(n11527), .ZN(
        n11529) );
  AOI21_X1 U14791 ( .B1(n11530), .B2(n19592), .A(n11529), .ZN(n11532) );
  AOI21_X1 U14792 ( .B1(n11535), .B2(n16280), .A(n11534), .ZN(n11863) );
  NAND2_X1 U14793 ( .A1(n11539), .A2(n11538), .ZN(n11540) );
  XNOR2_X1 U14794 ( .A(n11542), .B(n9752), .ZN(n15734) );
  NAND2_X1 U14795 ( .A1(n11543), .A2(n11544), .ZN(n11545) );
  NAND2_X1 U14796 ( .A1(n11546), .A2(n11545), .ZN(n16032) );
  OR2_X1 U14797 ( .A1(n16649), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16661) );
  NAND2_X1 U14798 ( .A1(n16666), .A2(n16661), .ZN(n16648) );
  AND2_X1 U14799 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11547) );
  NOR2_X1 U14800 ( .A1(n16649), .A2(n11547), .ZN(n11548) );
  OR2_X2 U14801 ( .A1(n16648), .A2(n11548), .ZN(n16638) );
  NOR2_X1 U14802 ( .A1(n17232), .A2(n11549), .ZN(n11550) );
  OR2_X1 U14803 ( .A1(n16638), .A2(n11550), .ZN(n16595) );
  NOR2_X1 U14804 ( .A1(n17232), .A2(n11555), .ZN(n11551) );
  NAND2_X1 U14805 ( .A1(n11552), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11553) );
  OR2_X1 U14806 ( .A1(n16649), .A2(n11553), .ZN(n16603) );
  NOR2_X1 U14807 ( .A1(n16603), .A2(n11554), .ZN(n16591) );
  AND2_X1 U14808 ( .A1(n16591), .A2(n11555), .ZN(n11556) );
  NAND2_X1 U14809 ( .A1(n11556), .A2(n16548), .ZN(n16547) );
  NAND2_X1 U14810 ( .A1(n16549), .A2(n16547), .ZN(n16538) );
  NAND2_X1 U14811 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n11556), .ZN(
        n16534) );
  NAND2_X1 U14812 ( .A1(n19571), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11866) );
  OAI21_X1 U14813 ( .B1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n16534), .A(
        n11866), .ZN(n11557) );
  AOI21_X1 U14814 ( .B1(n16538), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n11557), .ZN(n11558) );
  OAI21_X1 U14815 ( .B1(n17227), .B2(n16032), .A(n11558), .ZN(n11559) );
  NAND2_X1 U14816 ( .A1(n10889), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11561) );
  NAND2_X1 U14817 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20130) );
  INV_X1 U14818 ( .A(n20130), .ZN(n11562) );
  NAND2_X1 U14819 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n11562), .ZN(
        n11581) );
  INV_X1 U14820 ( .A(n11581), .ZN(n11563) );
  NAND2_X1 U14821 ( .A1(n11563), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19603) );
  NAND2_X1 U14822 ( .A1(n20284), .A2(n11581), .ZN(n11564) );
  AND3_X1 U14823 ( .A1(n19603), .A2(n20305), .A3(n11564), .ZN(n11565) );
  AOI21_X1 U14824 ( .B1(n11583), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n11565), .ZN(n11566) );
  INV_X1 U14825 ( .A(n11591), .ZN(n11569) );
  INV_X1 U14826 ( .A(n11570), .ZN(n11568) );
  NAND2_X1 U14827 ( .A1(n11569), .A2(n11568), .ZN(n11571) );
  INV_X1 U14828 ( .A(n13712), .ZN(n11575) );
  NAND2_X1 U14829 ( .A1(n19911), .A2(n19682), .ZN(n19871) );
  NAND2_X1 U14830 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19978) );
  AND2_X1 U14831 ( .A1(n19871), .A2(n19978), .ZN(n19805) );
  AND2_X1 U14832 ( .A1(n19805), .A2(n20305), .ZN(n19813) );
  AOI21_X1 U14833 ( .B1(n11583), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n19813), .ZN(n11573) );
  AOI22_X1 U14834 ( .A1(n11583), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20305), .B2(n19682), .ZN(n11576) );
  XNOR2_X1 U14835 ( .A(n11578), .B(n11579), .ZN(n13998) );
  NAND2_X1 U14836 ( .A1(n13997), .A2(n13998), .ZN(n13996) );
  INV_X1 U14837 ( .A(n11578), .ZN(n16768) );
  NAND2_X1 U14838 ( .A1(n16768), .A2(n11579), .ZN(n11580) );
  NAND2_X1 U14839 ( .A1(n19978), .A2(n20293), .ZN(n11582) );
  AOI22_X1 U14840 ( .A1(n11583), .A2(n10980), .B1(n20305), .B2(n19738), .ZN(
        n11584) );
  INV_X1 U14841 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11585) );
  INV_X1 U14842 ( .A(n11586), .ZN(n11587) );
  NAND2_X1 U14843 ( .A1(n11588), .A2(n11587), .ZN(n11589) );
  NAND2_X1 U14844 ( .A1(n10889), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11590) );
  NAND2_X1 U14845 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14264) );
  INV_X1 U14846 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14324) );
  NOR2_X1 U14847 ( .A1(n14264), .A2(n14324), .ZN(n11592) );
  NAND4_X1 U14848 ( .A1(n11593), .A2(n16058), .A3(n16069), .A4(n11592), .ZN(
        n11596) );
  NAND2_X1 U14849 ( .A1(n11594), .A2(n14326), .ZN(n11595) );
  NOR2_X1 U14850 ( .A1(n11596), .A2(n11595), .ZN(n14382) );
  AOI22_X1 U14851 ( .A1(n10651), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11678), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11600) );
  AOI22_X1 U14852 ( .A1(n11683), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10578), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11599) );
  AOI22_X1 U14853 ( .A1(n11685), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11684), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11598) );
  AOI22_X1 U14854 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11664), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11597) );
  NAND4_X1 U14855 ( .A1(n11600), .A2(n11599), .A3(n11598), .A4(n11597), .ZN(
        n11606) );
  AOI22_X1 U14856 ( .A1(n11675), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11677), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11604) );
  AOI22_X1 U14857 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11603) );
  AOI22_X1 U14858 ( .A1(n10548), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11602) );
  AOI22_X1 U14859 ( .A1(n10506), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10549), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11601) );
  NAND4_X1 U14860 ( .A1(n11604), .A2(n11603), .A3(n11602), .A4(n11601), .ZN(
        n11605) );
  OR2_X1 U14861 ( .A1(n11606), .A2(n11605), .ZN(n16043) );
  NAND3_X1 U14862 ( .A1(n11607), .A2(n16043), .A3(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11610) );
  NAND2_X1 U14863 ( .A1(n14425), .A2(n11608), .ZN(n11609) );
  NOR2_X1 U14864 ( .A1(n11610), .A2(n11609), .ZN(n11611) );
  AND3_X1 U14865 ( .A1(n14382), .A2(n14241), .A3(n11611), .ZN(n11612) );
  AOI22_X1 U14866 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n10651), .B1(
        n11678), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11616) );
  AOI22_X1 U14867 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11683), .B1(
        n10578), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11615) );
  AOI22_X1 U14868 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n11685), .B1(
        n11684), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11614) );
  AOI22_X1 U14869 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10507), .B1(
        n11664), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11613) );
  NAND4_X1 U14870 ( .A1(n11616), .A2(n11615), .A3(n11614), .A4(n11613), .ZN(
        n11622) );
  AOI22_X1 U14871 ( .A1(n11675), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n11677), .ZN(n11620) );
  AOI22_X1 U14872 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11619) );
  AOI22_X1 U14873 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10548), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11618) );
  AOI22_X1 U14874 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10549), .B1(
        n10506), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11617) );
  NAND4_X1 U14875 ( .A1(n11620), .A2(n11619), .A3(n11618), .A4(n11617), .ZN(
        n11621) );
  NOR2_X1 U14876 ( .A1(n11622), .A2(n11621), .ZN(n16041) );
  AOI22_X1 U14877 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n10651), .B1(
        n11678), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11626) );
  AOI22_X1 U14878 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n11683), .B1(
        n10578), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11625) );
  AOI22_X1 U14879 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n11685), .B1(
        n11684), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11624) );
  AOI22_X1 U14880 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10507), .B1(
        n11664), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11623) );
  NAND4_X1 U14881 ( .A1(n11626), .A2(n11625), .A3(n11624), .A4(n11623), .ZN(
        n11632) );
  AOI22_X1 U14882 ( .A1(n11675), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_14__2__SCAN_IN), .B2(n11677), .ZN(n11630) );
  AOI22_X1 U14883 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11629) );
  AOI22_X1 U14884 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10548), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11628) );
  AOI22_X1 U14885 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10549), .B1(
        n10506), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11627) );
  NAND4_X1 U14886 ( .A1(n11630), .A2(n11629), .A3(n11628), .A4(n11627), .ZN(
        n11631) );
  AOI22_X1 U14887 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n10651), .B1(
        n11678), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11636) );
  AOI22_X1 U14888 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n11683), .B1(
        n10578), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11635) );
  AOI22_X1 U14889 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n11685), .B1(
        n11684), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11634) );
  AOI22_X1 U14890 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10507), .B1(
        n11664), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11633) );
  NAND4_X1 U14891 ( .A1(n11636), .A2(n11635), .A3(n11634), .A4(n11633), .ZN(
        n11642) );
  AOI22_X1 U14892 ( .A1(n11675), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_14__3__SCAN_IN), .B2(n11677), .ZN(n11640) );
  AOI22_X1 U14893 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11639) );
  AOI22_X1 U14894 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10548), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11638) );
  AOI22_X1 U14895 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n10549), .B1(
        n10506), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11637) );
  NAND4_X1 U14896 ( .A1(n11640), .A2(n11639), .A3(n11638), .A4(n11637), .ZN(
        n11641) );
  AOI22_X1 U14897 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n10651), .B1(
        n11678), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11646) );
  AOI22_X1 U14898 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n11683), .B1(
        n10578), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11645) );
  AOI22_X1 U14899 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n11685), .B1(
        n11684), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11644) );
  AOI22_X1 U14900 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10507), .B1(
        n11664), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11643) );
  NAND4_X1 U14901 ( .A1(n11646), .A2(n11645), .A3(n11644), .A4(n11643), .ZN(
        n11652) );
  AOI22_X1 U14902 ( .A1(n11675), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_14__4__SCAN_IN), .B2(n10590), .ZN(n11650) );
  AOI22_X1 U14903 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11649) );
  AOI22_X1 U14904 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10548), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11648) );
  AOI22_X1 U14905 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10549), .B1(
        n10506), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11647) );
  NAND4_X1 U14906 ( .A1(n11650), .A2(n11649), .A3(n11648), .A4(n11647), .ZN(
        n11651) );
  AOI22_X1 U14907 ( .A1(n10651), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11678), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11656) );
  AOI22_X1 U14908 ( .A1(n11683), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10578), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11655) );
  AOI22_X1 U14909 ( .A1(n11685), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11684), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11654) );
  AOI22_X1 U14910 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11664), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11653) );
  NAND4_X1 U14911 ( .A1(n11656), .A2(n11655), .A3(n11654), .A4(n11653), .ZN(
        n11662) );
  AOI22_X1 U14912 ( .A1(n11675), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10590), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11660) );
  AOI22_X1 U14913 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11659) );
  AOI22_X1 U14914 ( .A1(n10548), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11658) );
  AOI22_X1 U14915 ( .A1(n10506), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10549), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11657) );
  NAND4_X1 U14916 ( .A1(n11660), .A2(n11659), .A3(n11658), .A4(n11657), .ZN(
        n11661) );
  NOR2_X1 U14917 ( .A1(n11662), .A2(n11661), .ZN(n16023) );
  AOI22_X1 U14918 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n10651), .B1(
        n11678), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11668) );
  AOI22_X1 U14919 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n11683), .B1(
        n10578), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11667) );
  AOI22_X1 U14920 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n11685), .B1(
        n11684), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11666) );
  AOI22_X1 U14921 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10507), .B1(
        n11664), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11665) );
  NAND4_X1 U14922 ( .A1(n11668), .A2(n11667), .A3(n11666), .A4(n11665), .ZN(
        n11674) );
  AOI22_X1 U14923 ( .A1(n11675), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_14__6__SCAN_IN), .B2(n10590), .ZN(n11672) );
  AOI22_X1 U14924 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11671) );
  AOI22_X1 U14925 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10548), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11670) );
  AOI22_X1 U14926 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10549), .B1(
        n10506), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11669) );
  NAND4_X1 U14927 ( .A1(n11672), .A2(n11671), .A3(n11670), .A4(n11669), .ZN(
        n11673) );
  NOR2_X1 U14928 ( .A1(n11674), .A2(n11673), .ZN(n16019) );
  AOI22_X1 U14929 ( .A1(n11675), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n10549), .ZN(n11682) );
  AOI22_X1 U14930 ( .A1(n11676), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10594), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11681) );
  AOI22_X1 U14931 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n10548), .B1(
        n11677), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11680) );
  AOI22_X1 U14932 ( .A1(n11678), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11679) );
  NAND4_X1 U14933 ( .A1(n11682), .A2(n11681), .A3(n11680), .A4(n11679), .ZN(
        n11691) );
  AOI22_X1 U14934 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n11683), .B1(
        n10578), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11689) );
  AOI22_X1 U14935 ( .A1(n10651), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10506), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11688) );
  AOI22_X1 U14936 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n11685), .B1(
        n11684), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11687) );
  AOI22_X1 U14937 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10507), .B1(
        n11664), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11686) );
  NAND4_X1 U14938 ( .A1(n11689), .A2(n11688), .A3(n11687), .A4(n11686), .ZN(
        n11690) );
  NAND2_X1 U14939 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11696) );
  AND2_X1 U14940 ( .A1(n10980), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11693) );
  OR2_X1 U14941 ( .A1(n11693), .A2(n11692), .ZN(n11841) );
  NAND2_X1 U14942 ( .A1(n11842), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11695) );
  AND3_X1 U14943 ( .A1(n11696), .A2(n11841), .A3(n11695), .ZN(n11706) );
  AOI22_X1 U14944 ( .A1(n11849), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11698), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11705) );
  AOI22_X1 U14945 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9612), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11704) );
  INV_X1 U14946 ( .A(n11700), .ZN(n11701) );
  INV_X1 U14947 ( .A(n11701), .ZN(n11847) );
  AOI22_X1 U14948 ( .A1(n11702), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11847), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11703) );
  NAND4_X1 U14949 ( .A1(n11706), .A2(n11705), .A3(n11704), .A4(n11703), .ZN(
        n11714) );
  NAND2_X1 U14950 ( .A1(n11702), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11708) );
  INV_X1 U14951 ( .A(n11841), .ZN(n11822) );
  NAND2_X1 U14952 ( .A1(n11842), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11707) );
  AND3_X1 U14953 ( .A1(n11708), .A2(n11822), .A3(n11707), .ZN(n11712) );
  AOI22_X1 U14954 ( .A1(n11849), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11698), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11711) );
  AOI22_X1 U14955 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9612), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11710) );
  AOI22_X1 U14956 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11847), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11709) );
  NAND4_X1 U14957 ( .A1(n11712), .A2(n11711), .A3(n11710), .A4(n11709), .ZN(
        n11713) );
  NAND2_X1 U14958 ( .A1(n11714), .A2(n11713), .ZN(n11738) );
  NOR2_X1 U14959 ( .A1(n11716), .A2(n11738), .ZN(n11715) );
  XOR2_X1 U14960 ( .A(n11719), .B(n11715), .Z(n11736) );
  INV_X1 U14961 ( .A(n11738), .ZN(n11718) );
  NAND2_X1 U14962 ( .A1(n11716), .A2(n11718), .ZN(n16014) );
  AND2_X1 U14963 ( .A1(n16018), .A2(n11736), .ZN(n11717) );
  NAND2_X1 U14964 ( .A1(n11719), .A2(n11718), .ZN(n11740) );
  NAND2_X1 U14965 ( .A1(n11842), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11721) );
  NAND2_X1 U14966 ( .A1(n11847), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11720) );
  AND3_X1 U14967 ( .A1(n11822), .A2(n11721), .A3(n11720), .ZN(n11725) );
  AOI22_X1 U14968 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11849), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11724) );
  AOI22_X1 U14969 ( .A1(n11702), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9602), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11723) );
  AOI22_X1 U14970 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(n9612), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11722) );
  NAND4_X1 U14971 ( .A1(n11725), .A2(n11724), .A3(n11723), .A4(n11722), .ZN(
        n11734) );
  AOI22_X1 U14972 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11849), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11732) );
  NAND2_X1 U14973 ( .A1(n11842), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11727) );
  NAND2_X1 U14974 ( .A1(n11847), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11726) );
  AND3_X1 U14975 ( .A1(n11727), .A2(n11841), .A3(n11726), .ZN(n11731) );
  AOI22_X1 U14976 ( .A1(n11702), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9603), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11730) );
  AOI22_X1 U14977 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(n9612), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11729) );
  NAND4_X1 U14978 ( .A1(n11732), .A2(n11731), .A3(n11730), .A4(n11729), .ZN(
        n11733) );
  NAND2_X1 U14979 ( .A1(n11734), .A2(n11733), .ZN(n11739) );
  XOR2_X1 U14980 ( .A(n11740), .B(n11739), .Z(n11735) );
  NAND2_X1 U14981 ( .A1(n11735), .A2(n14241), .ZN(n16006) );
  INV_X1 U14982 ( .A(n11739), .ZN(n11737) );
  NAND2_X1 U14983 ( .A1(n20314), .A2(n11737), .ZN(n16009) );
  NOR2_X1 U14984 ( .A1(n11740), .A2(n11739), .ZN(n11755) );
  NAND2_X1 U14985 ( .A1(n11842), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n11742) );
  NAND2_X1 U14986 ( .A1(n11847), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11741) );
  AND3_X1 U14987 ( .A1(n11822), .A2(n11742), .A3(n11741), .ZN(n11746) );
  AOI22_X1 U14988 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11849), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11745) );
  AOI22_X1 U14989 ( .A1(n11702), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11698), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11744) );
  AOI22_X1 U14990 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(n9612), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11743) );
  NAND4_X1 U14991 ( .A1(n11746), .A2(n11745), .A3(n11744), .A4(n11743), .ZN(
        n11754) );
  AOI22_X1 U14992 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11849), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11752) );
  NAND2_X1 U14993 ( .A1(n11842), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11748) );
  NAND2_X1 U14994 ( .A1(n11847), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11747) );
  AND3_X1 U14995 ( .A1(n11748), .A2(n11841), .A3(n11747), .ZN(n11751) );
  AOI22_X1 U14996 ( .A1(n11702), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11698), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11750) );
  AOI22_X1 U14997 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(n9612), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11749) );
  NAND4_X1 U14998 ( .A1(n11752), .A2(n11751), .A3(n11750), .A4(n11749), .ZN(
        n11753) );
  AND2_X1 U14999 ( .A1(n11754), .A2(n11753), .ZN(n11756) );
  NAND2_X1 U15000 ( .A1(n11755), .A2(n11756), .ZN(n11776) );
  OAI211_X1 U15001 ( .C1(n11755), .C2(n11756), .A(n14241), .B(n11776), .ZN(
        n11771) );
  NAND2_X1 U15002 ( .A1(n20314), .A2(n11756), .ZN(n16000) );
  NAND2_X1 U15003 ( .A1(n11842), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n11758) );
  NAND2_X1 U15004 ( .A1(n11847), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11757) );
  AND3_X1 U15005 ( .A1(n11822), .A2(n11758), .A3(n11757), .ZN(n11762) );
  AOI22_X1 U15006 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11849), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11761) );
  AOI22_X1 U15007 ( .A1(n11702), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9602), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11760) );
  AOI22_X1 U15008 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(n9612), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11759) );
  NAND4_X1 U15009 ( .A1(n11762), .A2(n11761), .A3(n11760), .A4(n11759), .ZN(
        n11770) );
  AOI22_X1 U15010 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11849), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11768) );
  NAND2_X1 U15011 ( .A1(n11842), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n11764) );
  NAND2_X1 U15012 ( .A1(n11847), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11763) );
  AND3_X1 U15013 ( .A1(n11764), .A2(n11841), .A3(n11763), .ZN(n11767) );
  AOI22_X1 U15014 ( .A1(n11702), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9603), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11766) );
  AOI22_X1 U15015 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(n9612), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11765) );
  NAND4_X1 U15016 ( .A1(n11768), .A2(n11767), .A3(n11766), .A4(n11765), .ZN(
        n11769) );
  NAND2_X1 U15017 ( .A1(n11770), .A2(n11769), .ZN(n15991) );
  INV_X1 U15018 ( .A(n11776), .ZN(n11774) );
  INV_X1 U15019 ( .A(n15991), .ZN(n11773) );
  AND2_X1 U15020 ( .A1(n11774), .A2(n11773), .ZN(n11794) );
  AOI211_X1 U15021 ( .C1(n15991), .C2(n11776), .A(n11775), .B(n11794), .ZN(
        n15994) );
  NAND2_X1 U15022 ( .A1(n15990), .A2(n15994), .ZN(n11777) );
  NAND2_X1 U15023 ( .A1(n11842), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11780) );
  NAND2_X1 U15024 ( .A1(n11847), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11779) );
  AND3_X1 U15025 ( .A1(n11822), .A2(n11780), .A3(n11779), .ZN(n11784) );
  AOI22_X1 U15026 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11849), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11783) );
  AOI22_X1 U15027 ( .A1(n11702), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9599), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11782) );
  AOI22_X1 U15028 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(n9612), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11781) );
  NAND4_X1 U15029 ( .A1(n11784), .A2(n11783), .A3(n11782), .A4(n11781), .ZN(
        n11792) );
  AOI22_X1 U15030 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11849), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11790) );
  NAND2_X1 U15031 ( .A1(n11842), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11786) );
  NAND2_X1 U15032 ( .A1(n11847), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11785) );
  AND3_X1 U15033 ( .A1(n11786), .A2(n11841), .A3(n11785), .ZN(n11789) );
  AOI22_X1 U15034 ( .A1(n11702), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11698), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11788) );
  AOI22_X1 U15035 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(n9612), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11787) );
  NAND4_X1 U15036 ( .A1(n11790), .A2(n11789), .A3(n11788), .A4(n11787), .ZN(
        n11791) );
  NAND2_X1 U15037 ( .A1(n11792), .A2(n11791), .ZN(n11797) );
  INV_X1 U15038 ( .A(n11797), .ZN(n11795) );
  INV_X1 U15039 ( .A(n11794), .ZN(n11793) );
  OAI211_X1 U15040 ( .C1(n11795), .C2(n11794), .A(n11829), .B(n14241), .ZN(
        n11796) );
  NOR2_X1 U15041 ( .A1(n15992), .A2(n11797), .ZN(n15986) );
  INV_X1 U15042 ( .A(n9666), .ZN(n11812) );
  NAND2_X1 U15043 ( .A1(n11842), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11799) );
  NAND2_X1 U15044 ( .A1(n11847), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11798) );
  AND3_X1 U15045 ( .A1(n11822), .A2(n11799), .A3(n11798), .ZN(n11803) );
  AOI22_X1 U15046 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11849), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11802) );
  AOI22_X1 U15047 ( .A1(n11702), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9603), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11801) );
  AOI22_X1 U15048 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(n9612), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11800) );
  NAND4_X1 U15049 ( .A1(n11803), .A2(n11802), .A3(n11801), .A4(n11800), .ZN(
        n11811) );
  AOI22_X1 U15050 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11849), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11809) );
  NAND2_X1 U15051 ( .A1(n11842), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11805) );
  NAND2_X1 U15052 ( .A1(n11847), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11804) );
  AND3_X1 U15053 ( .A1(n11805), .A2(n11841), .A3(n11804), .ZN(n11808) );
  AOI22_X1 U15054 ( .A1(n11702), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11698), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11807) );
  AOI22_X1 U15055 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(n9612), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11806) );
  NAND4_X1 U15056 ( .A1(n11809), .A2(n11808), .A3(n11807), .A4(n11806), .ZN(
        n11810) );
  NAND2_X1 U15057 ( .A1(n11811), .A2(n11810), .ZN(n11830) );
  NAND2_X1 U15058 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11814) );
  NAND2_X1 U15059 ( .A1(n11842), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11813) );
  AND3_X1 U15060 ( .A1(n11814), .A2(n11841), .A3(n11813), .ZN(n11819) );
  AOI22_X1 U15061 ( .A1(n11849), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9602), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11818) );
  AOI22_X1 U15062 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9612), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11817) );
  AOI22_X1 U15063 ( .A1(n11702), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11847), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11816) );
  NAND4_X1 U15064 ( .A1(n11819), .A2(n11818), .A3(n11817), .A4(n11816), .ZN(
        n11828) );
  NAND2_X1 U15065 ( .A1(n11842), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11821) );
  NAND2_X1 U15066 ( .A1(n9612), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11820) );
  AND3_X1 U15067 ( .A1(n11822), .A2(n11821), .A3(n11820), .ZN(n11826) );
  AOI22_X1 U15068 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11849), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11825) );
  AOI22_X1 U15069 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11698), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11824) );
  AOI22_X1 U15070 ( .A1(n11702), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11847), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11823) );
  NAND4_X1 U15071 ( .A1(n11826), .A2(n11825), .A3(n11824), .A4(n11823), .ZN(
        n11827) );
  NAND2_X1 U15072 ( .A1(n11828), .A2(n11827), .ZN(n11833) );
  INV_X1 U15073 ( .A(n11829), .ZN(n15980) );
  INV_X1 U15074 ( .A(n11830), .ZN(n15981) );
  AND2_X1 U15075 ( .A1(n10884), .A2(n15981), .ZN(n11831) );
  NAND2_X1 U15076 ( .A1(n15980), .A2(n11831), .ZN(n11832) );
  NOR2_X1 U15077 ( .A1(n11832), .A2(n11833), .ZN(n11834) );
  AOI21_X1 U15078 ( .B1(n11833), .B2(n11832), .A(n11834), .ZN(n15975) );
  INV_X1 U15079 ( .A(n11834), .ZN(n11835) );
  AOI22_X1 U15080 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11849), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11837) );
  AOI22_X1 U15081 ( .A1(n11847), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11698), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11836) );
  NAND2_X1 U15082 ( .A1(n11837), .A2(n11836), .ZN(n11855) );
  AOI22_X1 U15083 ( .A1(n11702), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9612), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11840) );
  NAND2_X1 U15084 ( .A1(n11842), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11839) );
  NAND2_X1 U15085 ( .A1(n9626), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11838) );
  NAND4_X1 U15086 ( .A1(n11840), .A2(n11839), .A3(n11838), .A4(n11841), .ZN(
        n11854) );
  AOI22_X1 U15087 ( .A1(n11702), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9612), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11844) );
  AOI21_X1 U15088 ( .B1(n11842), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n11841), .ZN(n11843) );
  OAI211_X1 U15089 ( .C1(n11846), .C2(n11845), .A(n11844), .B(n11843), .ZN(
        n11853) );
  AOI22_X1 U15090 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11847), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11851) );
  AOI22_X1 U15091 ( .A1(n11849), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9598), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11850) );
  NAND2_X1 U15092 ( .A1(n11851), .A2(n11850), .ZN(n11852) );
  OAI22_X1 U15093 ( .A1(n11855), .A2(n11854), .B1(n11853), .B2(n11852), .ZN(
        n11856) );
  NAND2_X1 U15094 ( .A1(n16846), .A2(n16848), .ZN(n11857) );
  NAND2_X1 U15095 ( .A1(n11857), .A2(n9729), .ZN(n11858) );
  NAND2_X1 U15096 ( .A1(n16073), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11862) );
  NAND2_X1 U15097 ( .A1(n11863), .A2(n19577), .ZN(n11873) );
  NAND2_X1 U15098 ( .A1(n13461), .A2(n15737), .ZN(n11865) );
  AND2_X1 U15099 ( .A1(n11865), .A2(n10120), .ZN(n15740) );
  OAI21_X1 U15100 ( .B1(n17198), .B2(n15737), .A(n11866), .ZN(n11868) );
  NOR2_X1 U15101 ( .A1(n16032), .A2(n19573), .ZN(n11867) );
  AOI211_X1 U15102 ( .C1(n17192), .C2(n15740), .A(n11868), .B(n11867), .ZN(
        n11869) );
  OAI21_X1 U15103 ( .B1(n11870), .B2(n19574), .A(n11869), .ZN(n11871) );
  NAND2_X1 U15104 ( .A1(n11873), .A2(n11872), .ZN(P2_U2995) );
  INV_X1 U15105 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18009) );
  INV_X1 U15106 ( .A(n11874), .ZN(n11883) );
  AND2_X2 U15107 ( .A1(n11875), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13685) );
  AOI22_X1 U15108 ( .A1(n13685), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11921), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11882) );
  NOR2_X2 U15109 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13761) );
  AND2_X1 U15110 ( .A1(n19196), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11876) );
  NOR2_X1 U15111 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11877) );
  AOI22_X1 U15112 ( .A1(n12119), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11994), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11881) );
  NOR2_X2 U15113 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11886) );
  NOR2_X1 U15114 ( .A1(n12170), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11878) );
  AND2_X2 U15115 ( .A1(n11886), .A2(n11878), .ZN(n11937) );
  AND2_X2 U15116 ( .A1(n13761), .A2(n11879), .ZN(n17767) );
  AOI22_X1 U15117 ( .A1(n11937), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17767), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11880) );
  NAND4_X1 U15118 ( .A1(n11883), .A2(n11882), .A3(n11881), .A4(n11880), .ZN(
        n11894) );
  AOI22_X1 U15119 ( .A1(n9578), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12136), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11892) );
  AND2_X2 U15120 ( .A1(n11885), .A2(n13784), .ZN(n13657) );
  AOI22_X1 U15121 ( .A1(n13657), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9573), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11891) );
  AND2_X2 U15122 ( .A1(n11886), .A2(n13784), .ZN(n11944) );
  AOI22_X1 U15123 ( .A1(n9581), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11944), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11890) );
  AND2_X2 U15124 ( .A1(n13785), .A2(n11887), .ZN(n11960) );
  NOR2_X1 U15125 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11888) );
  AOI22_X1 U15126 ( .A1(n11960), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13658), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11889) );
  NAND4_X1 U15127 ( .A1(n11892), .A2(n11891), .A3(n11890), .A4(n11889), .ZN(
        n11893) );
  INV_X1 U15128 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18014) );
  INV_X1 U15129 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11895) );
  OAI22_X1 U15130 ( .A1(n9568), .A2(n18014), .B1(n12117), .B2(n11895), .ZN(
        n11896) );
  INV_X1 U15131 ( .A(n11896), .ZN(n11900) );
  AOI22_X1 U15132 ( .A1(n13685), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11921), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11899) );
  AOI22_X1 U15133 ( .A1(n17903), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11994), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11898) );
  AOI22_X1 U15134 ( .A1(n11937), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17767), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11897) );
  AOI22_X1 U15135 ( .A1(n13657), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12136), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11904) );
  AOI22_X1 U15136 ( .A1(n9576), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(n9580), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11903) );
  AOI22_X1 U15137 ( .A1(n11960), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11944), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11902) );
  AOI22_X1 U15138 ( .A1(n9572), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13658), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11901) );
  INV_X1 U15139 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13702) );
  INV_X1 U15140 ( .A(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12053) );
  INV_X1 U15141 ( .A(n11905), .ZN(n11909) );
  AOI22_X1 U15142 ( .A1(n13685), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11921), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11908) );
  INV_X1 U15143 ( .A(n10404), .ZN(n17903) );
  AOI22_X1 U15144 ( .A1(n12119), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11994), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11907) );
  AOI22_X1 U15145 ( .A1(n11937), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17767), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11906) );
  NAND4_X1 U15146 ( .A1(n11909), .A2(n11908), .A3(n11907), .A4(n11906), .ZN(
        n11915) );
  AOI22_X1 U15147 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17954), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11913) );
  AOI22_X1 U15148 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17953), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11912) );
  AOI22_X1 U15149 ( .A1(n9577), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11911) );
  AOI22_X1 U15150 ( .A1(n9582), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17834), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11910) );
  NAND4_X1 U15151 ( .A1(n11913), .A2(n11912), .A3(n11911), .A4(n11910), .ZN(
        n11914) );
  AND2_X1 U15152 ( .A1(n13938), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14188) );
  NAND2_X1 U15153 ( .A1(n13885), .A2(n14188), .ZN(n11917) );
  INV_X1 U15154 ( .A(n13934), .ZN(n12226) );
  NAND2_X1 U15155 ( .A1(n12226), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11916) );
  NAND2_X1 U15156 ( .A1(n11917), .A2(n11916), .ZN(n18486) );
  NAND2_X1 U15157 ( .A1(n18487), .A2(n18486), .ZN(n11920) );
  INV_X1 U15158 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18727) );
  OR2_X1 U15159 ( .A1(n11918), .A2(n18727), .ZN(n11919) );
  NAND2_X1 U15160 ( .A1(n11920), .A2(n11919), .ZN(n11935) );
  INV_X1 U15161 ( .A(n11936), .ZN(n11933) );
  AOI22_X1 U15162 ( .A1(n11937), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17767), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11925) );
  AOI22_X1 U15163 ( .A1(n12119), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11994), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11924) );
  NAND2_X1 U15164 ( .A1(n17817), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n11923) );
  NAND2_X1 U15165 ( .A1(n11921), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11922) );
  NAND4_X1 U15166 ( .A1(n11925), .A2(n11924), .A3(n11923), .A4(n11922), .ZN(
        n11927) );
  INV_X1 U15167 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18002) );
  OAI22_X1 U15168 ( .A1(n18002), .A2(n9568), .B1(n12117), .B2(n14060), .ZN(
        n11926) );
  NOR2_X1 U15169 ( .A1(n11927), .A2(n11926), .ZN(n11932) );
  AOI22_X1 U15170 ( .A1(n13657), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12136), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11931) );
  AOI22_X1 U15171 ( .A1(n9572), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(n9580), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11930) );
  AOI22_X1 U15172 ( .A1(n14172), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11929) );
  AOI22_X1 U15173 ( .A1(n9577), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13658), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11928) );
  XNOR2_X1 U15174 ( .A(n11933), .B(n18122), .ZN(n11934) );
  INV_X1 U15175 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21349) );
  AOI22_X1 U15176 ( .A1(n17975), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17974), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11941) );
  AOI22_X1 U15177 ( .A1(n12119), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11994), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11940) );
  NAND2_X1 U15178 ( .A1(n17817), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11939) );
  INV_X4 U15179 ( .A(n17931), .ZN(n17818) );
  NAND2_X1 U15180 ( .A1(n17818), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11938) );
  NAND4_X1 U15181 ( .A1(n11941), .A2(n11940), .A3(n11939), .A4(n11938), .ZN(
        n11943) );
  INV_X1 U15182 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17997) );
  INV_X1 U15183 ( .A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12091) );
  OAI22_X1 U15184 ( .A1(n17997), .A2(n17844), .B1(n12117), .B2(n12091), .ZN(
        n11942) );
  NOR2_X1 U15185 ( .A1(n11943), .A2(n11942), .ZN(n11949) );
  AOI22_X1 U15186 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12136), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11948) );
  AOI22_X1 U15187 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(n9582), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11947) );
  AOI22_X1 U15188 ( .A1(n9578), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17953), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11946) );
  BUF_X4 U15189 ( .A(n11944), .Z(n17932) );
  AOI22_X1 U15190 ( .A1(n17932), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17834), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11945) );
  INV_X1 U15191 ( .A(n18117), .ZN(n11950) );
  NAND2_X1 U15192 ( .A1(n11951), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11952) );
  INV_X1 U15193 ( .A(n11973), .ZN(n11967) );
  INV_X1 U15194 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11954) );
  INV_X1 U15195 ( .A(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12064) );
  OAI22_X1 U15196 ( .A1(n17844), .A2(n11954), .B1(n12117), .B2(n12064), .ZN(
        n11955) );
  INV_X1 U15197 ( .A(n11955), .ZN(n11959) );
  AOI22_X1 U15198 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17818), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11958) );
  AOI22_X1 U15199 ( .A1(n12119), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17973), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11957) );
  AOI22_X1 U15200 ( .A1(n11937), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17767), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11956) );
  NAND4_X1 U15201 ( .A1(n11959), .A2(n11958), .A3(n11957), .A4(n11956), .ZN(
        n11966) );
  AOI22_X1 U15202 ( .A1(n13657), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12136), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11964) );
  AOI22_X1 U15203 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(n9581), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11963) );
  AOI22_X1 U15204 ( .A1(n14172), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11962) );
  AOI22_X1 U15205 ( .A1(n9577), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13658), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11961) );
  NAND4_X1 U15206 ( .A1(n11964), .A2(n11963), .A3(n11962), .A4(n11961), .ZN(
        n11965) );
  XNOR2_X1 U15207 ( .A(n11967), .B(n18113), .ZN(n11968) );
  XNOR2_X1 U15208 ( .A(n11970), .B(n11968), .ZN(n18461) );
  NAND2_X1 U15209 ( .A1(n18461), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11972) );
  INV_X1 U15210 ( .A(n11968), .ZN(n11969) );
  NAND2_X1 U15211 ( .A1(n11970), .A2(n11969), .ZN(n11971) );
  NAND2_X1 U15212 ( .A1(n11972), .A2(n11971), .ZN(n13986) );
  INV_X1 U15213 ( .A(n11993), .ZN(n11987) );
  INV_X2 U15214 ( .A(n14037), .ZN(n17975) );
  AOI22_X1 U15215 ( .A1(n17975), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17767), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11977) );
  AOI22_X1 U15216 ( .A1(n12119), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17973), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11976) );
  NAND2_X1 U15217 ( .A1(n17817), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11975) );
  NAND2_X1 U15218 ( .A1(n17818), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n11974) );
  NAND4_X1 U15219 ( .A1(n11977), .A2(n11976), .A3(n11975), .A4(n11974), .ZN(
        n11979) );
  INV_X1 U15220 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17982) );
  INV_X1 U15221 ( .A(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12075) );
  OAI22_X1 U15222 ( .A1(n17982), .A2(n17844), .B1(n12117), .B2(n12075), .ZN(
        n11978) );
  NOR2_X1 U15223 ( .A1(n11979), .A2(n11978), .ZN(n11986) );
  CLKBUF_X3 U15224 ( .A(n11980), .Z(n17954) );
  AOI22_X1 U15225 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17954), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11984) );
  AOI22_X1 U15226 ( .A1(n9577), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(n9582), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11983) );
  AOI22_X1 U15227 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17953), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11982) );
  AOI22_X1 U15228 ( .A1(n17932), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17834), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11981) );
  XNOR2_X1 U15229 ( .A(n11987), .B(n18110), .ZN(n11988) );
  XNOR2_X1 U15230 ( .A(n11988), .B(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13985) );
  NAND2_X1 U15231 ( .A1(n13986), .A2(n13985), .ZN(n11991) );
  INV_X1 U15232 ( .A(n11988), .ZN(n11989) );
  NAND2_X1 U15233 ( .A1(n11989), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11990) );
  NAND2_X1 U15234 ( .A1(n11991), .A2(n11990), .ZN(n12010) );
  INV_X1 U15235 ( .A(n18110), .ZN(n11992) );
  INV_X1 U15236 ( .A(n17767), .ZN(n13684) );
  INV_X2 U15237 ( .A(n13684), .ZN(n17974) );
  AOI22_X1 U15238 ( .A1(n17974), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12119), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11998) );
  AOI22_X1 U15239 ( .A1(n17975), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17973), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11997) );
  NAND2_X1 U15240 ( .A1(n17817), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11996) );
  NAND2_X1 U15241 ( .A1(n17818), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11995) );
  NAND4_X1 U15242 ( .A1(n11998), .A2(n11997), .A3(n11996), .A4(n11995), .ZN(
        n12000) );
  INV_X1 U15243 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13688) );
  OAI22_X1 U15244 ( .A1(n13688), .A2(n17844), .B1(n12117), .B2(n13686), .ZN(
        n11999) );
  NOR2_X1 U15245 ( .A1(n12000), .A2(n11999), .ZN(n12006) );
  AOI22_X1 U15246 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17954), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12004) );
  AOI22_X1 U15247 ( .A1(n9572), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(n9583), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12003) );
  AOI22_X1 U15248 ( .A1(n17953), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12002) );
  AOI22_X1 U15249 ( .A1(n9578), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17834), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12001) );
  INV_X1 U15250 ( .A(n17039), .ZN(n17050) );
  NAND2_X1 U15251 ( .A1(n17050), .A2(n16880), .ZN(n12007) );
  NAND2_X1 U15252 ( .A1(n18357), .A2(n12007), .ZN(n12008) );
  INV_X1 U15253 ( .A(n12008), .ZN(n12009) );
  NAND2_X1 U15254 ( .A1(n12010), .A2(n12009), .ZN(n12011) );
  INV_X1 U15255 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18415) );
  INV_X1 U15256 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18409) );
  INV_X1 U15257 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18676) );
  NAND3_X1 U15258 ( .A1(n18415), .A2(n18409), .A3(n18676), .ZN(n12013) );
  INV_X1 U15259 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18619) );
  INV_X1 U15260 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16978) );
  NAND2_X1 U15261 ( .A1(n18619), .A2(n16978), .ZN(n12014) );
  NAND2_X1 U15262 ( .A1(n18357), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16979) );
  NAND2_X1 U15263 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18649) );
  NOR2_X1 U15264 ( .A1(n18649), .A2(n18415), .ZN(n18664) );
  NAND2_X1 U15265 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18664), .ZN(
        n18630) );
  NOR2_X1 U15266 ( .A1(n18630), .A2(n18384), .ZN(n18600) );
  NAND2_X1 U15267 ( .A1(n18600), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n18590) );
  NAND2_X1 U15268 ( .A1(n18343), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12016) );
  INV_X1 U15269 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18583) );
  NAND2_X1 U15270 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18293) );
  INV_X1 U15271 ( .A(n18293), .ZN(n18542) );
  AND2_X1 U15272 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18542), .ZN(
        n18526) );
  AND2_X1 U15273 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18573) );
  NAND2_X1 U15274 ( .A1(n18573), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18519) );
  INV_X1 U15275 ( .A(n18519), .ZN(n18538) );
  AND2_X1 U15276 ( .A1(n18522), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16946) );
  NAND2_X1 U15277 ( .A1(n16946), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16931) );
  INV_X1 U15278 ( .A(n16931), .ZN(n12017) );
  NAND2_X1 U15279 ( .A1(n18525), .A2(n12017), .ZN(n16943) );
  INV_X1 U15280 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18299) );
  NAND2_X1 U15281 ( .A1(n18330), .A2(n18299), .ZN(n12018) );
  NOR2_X1 U15282 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n12018), .ZN(
        n18284) );
  INV_X1 U15283 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18286) );
  NOR2_X1 U15284 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12019) );
  NAND2_X1 U15285 ( .A1(n18269), .A2(n12019), .ZN(n12020) );
  NAND2_X1 U15286 ( .A1(n16943), .A2(n12020), .ZN(n12021) );
  INV_X1 U15287 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12022) );
  NAND2_X1 U15288 ( .A1(n18525), .A2(n18573), .ZN(n12023) );
  AND3_X1 U15289 ( .A1(n18526), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12024) );
  NOR2_X1 U15290 ( .A1(n18357), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12025) );
  NAND2_X1 U15291 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17063) );
  INV_X1 U15292 ( .A(n17063), .ZN(n12029) );
  OR2_X1 U15293 ( .A1(n18357), .A2(n12029), .ZN(n12030) );
  INV_X1 U15294 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17248) );
  INV_X1 U15295 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13765) );
  NAND2_X1 U15296 ( .A1(n18357), .A2(n13765), .ZN(n12034) );
  INV_X1 U15297 ( .A(n12034), .ZN(n12032) );
  INV_X1 U15298 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n17031) );
  AOI21_X1 U15299 ( .B1(n18357), .B2(n17031), .A(n13765), .ZN(n12031) );
  AOI211_X1 U15300 ( .C1(n16890), .C2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n12032), .B(n12031), .ZN(n12037) );
  INV_X1 U15301 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17106) );
  NAND3_X1 U15302 ( .A1(n17053), .A2(n18357), .A3(n17106), .ZN(n17104) );
  NOR2_X2 U15303 ( .A1(n17104), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16891) );
  INV_X1 U15304 ( .A(n16891), .ZN(n12033) );
  NAND2_X1 U15305 ( .A1(n12033), .A2(n18357), .ZN(n12036) );
  AND2_X1 U15306 ( .A1(n13765), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12253) );
  AOI22_X1 U15307 ( .A1(n17948), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17947), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12041) );
  AOI22_X1 U15308 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17818), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12040) );
  AOI22_X1 U15309 ( .A1(n12119), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17973), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12039) );
  AOI22_X1 U15310 ( .A1(n11937), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17767), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12038) );
  NAND4_X1 U15311 ( .A1(n12041), .A2(n12040), .A3(n12039), .A4(n12038), .ZN(
        n12047) );
  AOI22_X1 U15312 ( .A1(n9578), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(n9572), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12045) );
  AOI22_X1 U15313 ( .A1(n17954), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9583), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12044) );
  AOI22_X1 U15314 ( .A1(n17953), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12043) );
  AOI22_X1 U15315 ( .A1(n17966), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17967), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12042) );
  NAND4_X1 U15316 ( .A1(n12045), .A2(n12044), .A3(n12043), .A4(n12042), .ZN(
        n12046) );
  AOI22_X1 U15317 ( .A1(n11937), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17767), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12051) );
  AOI22_X1 U15318 ( .A1(n12119), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17973), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12050) );
  NAND2_X1 U15319 ( .A1(n17817), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12049) );
  NAND2_X1 U15320 ( .A1(n17818), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12048) );
  NAND4_X1 U15321 ( .A1(n12051), .A2(n12050), .A3(n12049), .A4(n12048), .ZN(
        n12055) );
  INV_X1 U15322 ( .A(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12052) );
  OAI22_X1 U15323 ( .A1(n17844), .A2(n12053), .B1(n12117), .B2(n12052), .ZN(
        n12054) );
  AOI22_X1 U15324 ( .A1(n13657), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12136), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12059) );
  AOI22_X1 U15325 ( .A1(n9572), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(n9580), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12058) );
  AOI22_X1 U15326 ( .A1(n14172), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12057) );
  AOI22_X1 U15327 ( .A1(n9576), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17967), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12056) );
  NAND2_X1 U15328 ( .A1(n18755), .A2(n19335), .ZN(n12062) );
  INV_X1 U15329 ( .A(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12063) );
  INV_X1 U15330 ( .A(n12065), .ZN(n12069) );
  AOI22_X1 U15331 ( .A1(n17817), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17818), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12068) );
  AOI22_X1 U15332 ( .A1(n12119), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11994), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12067) );
  AOI22_X1 U15333 ( .A1(n11937), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17767), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12066) );
  AOI22_X1 U15334 ( .A1(n9576), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(n9573), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12073) );
  AOI22_X1 U15335 ( .A1(n13657), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12136), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12072) );
  AOI22_X1 U15336 ( .A1(n9581), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12071) );
  AOI22_X1 U15337 ( .A1(n14172), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13658), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12070) );
  INV_X1 U15338 ( .A(n18775), .ZN(n12143) );
  INV_X1 U15339 ( .A(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12074) );
  OAI22_X1 U15340 ( .A1(n17844), .A2(n12075), .B1(n17981), .B2(n12074), .ZN(
        n12076) );
  INV_X1 U15341 ( .A(n12076), .ZN(n12080) );
  AOI22_X1 U15342 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17818), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12079) );
  AOI22_X1 U15343 ( .A1(n12119), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17973), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12078) );
  AOI22_X1 U15344 ( .A1(n11937), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17767), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12077) );
  NAND4_X1 U15345 ( .A1(n12080), .A2(n12079), .A3(n12078), .A4(n12077), .ZN(
        n12086) );
  AOI22_X1 U15346 ( .A1(n17954), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9574), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12084) );
  AOI22_X1 U15347 ( .A1(n9577), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17953), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12083) );
  AOI22_X1 U15348 ( .A1(n9582), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12082) );
  AOI22_X1 U15349 ( .A1(n13657), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17967), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12081) );
  NAND4_X1 U15350 ( .A1(n12084), .A2(n12083), .A3(n12082), .A4(n12081), .ZN(
        n12085) );
  OR2_X2 U15351 ( .A1(n12086), .A2(n12085), .ZN(n18779) );
  AOI22_X1 U15352 ( .A1(n11937), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17767), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12090) );
  AOI22_X1 U15353 ( .A1(n12119), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17973), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12089) );
  NAND2_X1 U15354 ( .A1(n17817), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n12088) );
  NAND2_X1 U15355 ( .A1(n17818), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n12087) );
  NAND4_X1 U15356 ( .A1(n12090), .A2(n12089), .A3(n12088), .A4(n12087), .ZN(
        n12093) );
  INV_X4 U15357 ( .A(n17947), .ZN(n17981) );
  OAI22_X1 U15358 ( .A1(n21286), .A2(n17981), .B1(n9568), .B2(n12091), .ZN(
        n12092) );
  NOR2_X1 U15359 ( .A1(n12093), .A2(n12092), .ZN(n12099) );
  AOI22_X1 U15360 ( .A1(n13657), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12136), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12097) );
  AOI22_X1 U15361 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(n9581), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12096) );
  AOI22_X1 U15362 ( .A1(n17953), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12095) );
  AOI22_X1 U15363 ( .A1(n9577), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13658), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12094) );
  NAND2_X1 U15364 ( .A1(n18770), .A2(n18755), .ZN(n12100) );
  INV_X1 U15365 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n21266) );
  AOI22_X1 U15366 ( .A1(n17975), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17974), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12105) );
  AOI22_X1 U15367 ( .A1(n12119), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17973), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12104) );
  NAND2_X1 U15368 ( .A1(n17817), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n12103) );
  NAND2_X1 U15369 ( .A1(n17818), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n12102) );
  NAND4_X1 U15370 ( .A1(n12105), .A2(n12104), .A3(n12103), .A4(n12102), .ZN(
        n12108) );
  INV_X1 U15371 ( .A(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14060) );
  INV_X1 U15372 ( .A(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12106) );
  OAI22_X1 U15373 ( .A1(n14060), .A2(n17844), .B1(n17981), .B2(n12106), .ZN(
        n12107) );
  NOR2_X1 U15374 ( .A1(n12108), .A2(n12107), .ZN(n12115) );
  AOI22_X1 U15375 ( .A1(n13657), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17954), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12113) );
  AOI22_X1 U15376 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(n9580), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12112) );
  AOI22_X1 U15377 ( .A1(n14172), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12111) );
  AOI22_X1 U15378 ( .A1(n9577), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13658), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12110) );
  INV_X1 U15379 ( .A(n12154), .ZN(n18766) );
  INV_X1 U15380 ( .A(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12116) );
  OAI22_X1 U15381 ( .A1(n17844), .A2(n13686), .B1(n12117), .B2(n12116), .ZN(
        n12118) );
  INV_X1 U15382 ( .A(n12118), .ZN(n12123) );
  AOI22_X1 U15383 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n17818), .B1(
        n17972), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12122) );
  AOI22_X1 U15384 ( .A1(n12119), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17973), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12121) );
  AOI22_X1 U15385 ( .A1(n11937), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17767), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12120) );
  NAND4_X1 U15386 ( .A1(n12123), .A2(n12122), .A3(n12121), .A4(n12120), .ZN(
        n12129) );
  AOI22_X1 U15387 ( .A1(n17966), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12136), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12127) );
  AOI22_X1 U15388 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(n9583), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12126) );
  AOI22_X1 U15389 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n14172), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12125) );
  AOI22_X1 U15390 ( .A1(n9578), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17967), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12124) );
  NAND4_X1 U15391 ( .A1(n12127), .A2(n12126), .A3(n12125), .A4(n12124), .ZN(
        n12128) );
  AOI22_X1 U15392 ( .A1(n11937), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17974), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12133) );
  AOI22_X1 U15393 ( .A1(n12119), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17973), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12132) );
  NAND2_X1 U15394 ( .A1(n17817), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n12131) );
  NAND2_X1 U15395 ( .A1(n17818), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n12130) );
  NAND4_X1 U15396 ( .A1(n12133), .A2(n12132), .A3(n12131), .A4(n12130), .ZN(
        n12135) );
  OAI22_X1 U15397 ( .A1(n17844), .A2(n13847), .B1(n17981), .B2(n21252), .ZN(
        n12134) );
  NOR2_X1 U15398 ( .A1(n12135), .A2(n12134), .ZN(n12142) );
  AOI22_X1 U15399 ( .A1(n13657), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12136), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12140) );
  AOI22_X1 U15400 ( .A1(n9572), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(n9583), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12139) );
  AOI22_X1 U15401 ( .A1(n17953), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12138) );
  AOI22_X1 U15402 ( .A1(n9576), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13658), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12137) );
  AND2_X1 U15403 ( .A1(n12143), .A2(n12194), .ZN(n12144) );
  INV_X1 U15404 ( .A(n18755), .ZN(n14103) );
  NAND3_X1 U15405 ( .A1(n14103), .A2(n12154), .A3(n18783), .ZN(n12164) );
  NAND2_X1 U15406 ( .A1(n12158), .A2(n18770), .ZN(n12146) );
  NAND2_X1 U15407 ( .A1(n12169), .A2(n18762), .ZN(n12204) );
  INV_X1 U15408 ( .A(n13608), .ZN(n12147) );
  NAND2_X1 U15409 ( .A1(n13753), .A2(n12151), .ZN(n13665) );
  NAND2_X1 U15410 ( .A1(n13754), .A2(n13753), .ZN(n12166) );
  OR3_X1 U15411 ( .A1(n12150), .A2(n18178), .A3(n12200), .ZN(n12165) );
  NOR2_X1 U15412 ( .A1(n18779), .A2(n18770), .ZN(n13752) );
  NAND2_X1 U15413 ( .A1(n12194), .A2(n18775), .ZN(n12198) );
  INV_X1 U15414 ( .A(n18779), .ZN(n12152) );
  NAND2_X1 U15415 ( .A1(n18178), .A2(n18755), .ZN(n12153) );
  AOI21_X1 U15416 ( .B1(n18783), .B2(n13930), .A(n12153), .ZN(n12202) );
  AOI211_X1 U15417 ( .C1(n12161), .C2(n12198), .A(n12154), .B(n12202), .ZN(
        n12155) );
  INV_X1 U15418 ( .A(n12155), .ZN(n12163) );
  OAI21_X1 U15419 ( .B1(n18178), .B2(n18755), .A(n12194), .ZN(n12156) );
  AOI21_X1 U15420 ( .B1(n18770), .B2(n13728), .A(n12156), .ZN(n12199) );
  NOR2_X1 U15421 ( .A1(n12158), .A2(n17863), .ZN(n12157) );
  OAI22_X1 U15422 ( .A1(n12199), .A2(n12158), .B1(n18770), .B2(n12157), .ZN(
        n12159) );
  INV_X1 U15423 ( .A(n12159), .ZN(n12160) );
  OAI21_X1 U15424 ( .B1(n18755), .B2(n12161), .A(n12160), .ZN(n12162) );
  NOR2_X1 U15425 ( .A1(n18762), .A2(n18770), .ZN(n12167) );
  NAND2_X1 U15426 ( .A1(n12169), .A2(n12168), .ZN(n13606) );
  AND2_X1 U15427 ( .A1(n12194), .A2(n19335), .ZN(n12186) );
  MUX2_X1 U15428 ( .A(n12171), .B(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        n12170), .Z(n12188) );
  MUX2_X1 U15429 ( .A(n12172), .B(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        n13758), .Z(n12175) );
  OAI22_X1 U15430 ( .A1(n12177), .A2(n12175), .B1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n13758), .ZN(n12173) );
  NOR2_X1 U15431 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19188), .ZN(
        n12174) );
  NAND2_X1 U15432 ( .A1(n12173), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12183) );
  AOI22_X1 U15433 ( .A1(n12182), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B1(
        n12174), .B2(n12183), .ZN(n12192) );
  INV_X1 U15434 ( .A(n12175), .ZN(n12176) );
  XNOR2_X1 U15435 ( .A(n12177), .B(n12176), .ZN(n12178) );
  NAND2_X1 U15436 ( .A1(n12192), .A2(n12178), .ZN(n12189) );
  OAI21_X1 U15437 ( .B1(n21323), .B2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n12180), .ZN(n12187) );
  AOI21_X1 U15438 ( .B1(n12180), .B2(n12188), .A(n12179), .ZN(n12181) );
  INV_X1 U15439 ( .A(n12181), .ZN(n12185) );
  AOI21_X1 U15440 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n12183), .A(
        n12182), .ZN(n12184) );
  OAI21_X1 U15441 ( .B1(n12189), .B2(n12187), .A(n19185), .ZN(n19177) );
  NAND2_X1 U15442 ( .A1(n12186), .A2(n18779), .ZN(n12206) );
  NOR2_X1 U15443 ( .A1(n12188), .A2(n12187), .ZN(n12193) );
  NAND2_X1 U15444 ( .A1(n12190), .A2(n12189), .ZN(n12191) );
  NAND2_X2 U15445 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n19261), .ZN(n19306) );
  INV_X1 U15446 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n21319) );
  NAND2_X1 U15447 ( .A1(n21319), .A2(n17353), .ZN(n19234) );
  NAND3_X1 U15448 ( .A1(n19235), .A2(n19306), .A3(n19234), .ZN(n19243) );
  XNOR2_X1 U15449 ( .A(n12194), .B(n19335), .ZN(n12195) );
  NAND2_X1 U15450 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n19222) );
  OAI21_X1 U15451 ( .B1(n19334), .B2(n12195), .A(n19222), .ZN(n17360) );
  OAI21_X1 U15452 ( .B1(n17360), .B2(n12196), .A(n12198), .ZN(n12197) );
  OAI21_X1 U15453 ( .B1(n19180), .B2(n12198), .A(n12197), .ZN(n12205) );
  OAI211_X1 U15454 ( .C1(n12201), .C2(n13728), .A(n12200), .B(n12199), .ZN(
        n12203) );
  AOI21_X1 U15455 ( .B1(n12204), .B2(n12203), .A(n12202), .ZN(n13724) );
  OAI211_X1 U15456 ( .C1(n19177), .C2(n12206), .A(n12205), .B(n13724), .ZN(
        n12208) );
  NAND2_X1 U15457 ( .A1(n16878), .A2(n18672), .ZN(n12258) );
  NOR2_X1 U15458 ( .A1(n18590), .A2(n16978), .ZN(n18568) );
  NAND3_X1 U15459 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12209) );
  INV_X1 U15460 ( .A(n12209), .ZN(n13989) );
  AOI21_X1 U15461 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18718) );
  INV_X1 U15462 ( .A(n18718), .ZN(n14116) );
  NAND2_X1 U15463 ( .A1(n13989), .A2(n14116), .ZN(n13981) );
  NAND3_X1 U15464 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18566) );
  NOR2_X1 U15465 ( .A1(n13981), .A2(n18566), .ZN(n18650) );
  NAND2_X1 U15466 ( .A1(n18568), .A2(n18650), .ZN(n18571) );
  INV_X1 U15467 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18678) );
  NAND2_X1 U15468 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14118) );
  NOR2_X1 U15469 ( .A1(n12209), .A2(n14118), .ZN(n13983) );
  NAND3_X1 U15470 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n13983), .ZN(n18679) );
  NOR2_X1 U15471 ( .A1(n18678), .A2(n18679), .ZN(n12212) );
  NAND2_X1 U15472 ( .A1(n18568), .A2(n12212), .ZN(n12213) );
  INV_X1 U15473 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13980) );
  NAND2_X1 U15474 ( .A1(n18730), .A2(n13980), .ZN(n13887) );
  NOR2_X1 U15475 ( .A1(n18658), .A2(n18680), .ZN(n18713) );
  NAND2_X1 U15476 ( .A1(n13887), .A2(n18576), .ZN(n18709) );
  OAI22_X1 U15477 ( .A1(n18712), .A2(n18571), .B1(n12213), .B2(n18709), .ZN(
        n17026) );
  NAND2_X1 U15478 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18501) );
  INV_X1 U15479 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18509) );
  NOR3_X1 U15480 ( .A1(n18501), .A2(n18509), .A3(n12028), .ZN(n17073) );
  NAND2_X1 U15481 ( .A1(n16946), .A2(n17073), .ZN(n17027) );
  INV_X1 U15482 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17070) );
  NOR2_X1 U15483 ( .A1(n17106), .A2(n17070), .ZN(n17112) );
  NAND2_X1 U15484 ( .A1(n17112), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16895) );
  INV_X1 U15485 ( .A(n12253), .ZN(n12210) );
  NOR4_X1 U15486 ( .A1(n18616), .A2(n17027), .A3(n16895), .A4(n12210), .ZN(
        n12251) );
  AND2_X1 U15487 ( .A1(n18593), .A2(n18724), .ZN(n14119) );
  NOR2_X1 U15488 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n12211) );
  NAND2_X2 U15489 ( .A1(n19350), .A2(n12211), .ZN(n18739) );
  INV_X1 U15490 ( .A(n18658), .ZN(n18683) );
  INV_X1 U15491 ( .A(n17073), .ZN(n12214) );
  NAND2_X1 U15492 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n12212), .ZN(
        n18657) );
  INV_X1 U15493 ( .A(n18657), .ZN(n18684) );
  AND2_X1 U15494 ( .A1(n18568), .A2(n18684), .ZN(n18592) );
  NAND2_X1 U15495 ( .A1(n16946), .A2(n18592), .ZN(n18528) );
  NOR3_X1 U15496 ( .A1(n12214), .A2(n17070), .A3(n18528), .ZN(n12216) );
  OAI21_X1 U15497 ( .B1(n17027), .B2(n18571), .A(n19179), .ZN(n17067) );
  INV_X1 U15498 ( .A(n12213), .ZN(n18570) );
  NAND2_X1 U15499 ( .A1(n16946), .A2(n18570), .ZN(n17066) );
  OAI21_X1 U15500 ( .B1(n12214), .B2(n17066), .A(n18680), .ZN(n12215) );
  OAI211_X1 U15501 ( .C1(n18683), .C2(n12216), .A(n17067), .B(n12215), .ZN(
        n17045) );
  AOI22_X1 U15502 ( .A1(n14119), .A2(n16895), .B1(n17045), .B2(n18724), .ZN(
        n17032) );
  INV_X1 U15503 ( .A(n17032), .ZN(n12217) );
  AOI211_X1 U15504 ( .C1(n14119), .C2(n17031), .A(n18701), .B(n12217), .ZN(
        n12250) );
  NAND2_X1 U15505 ( .A1(n13934), .A2(n13938), .ZN(n12227) );
  INV_X1 U15506 ( .A(n12224), .ZN(n14021) );
  NAND2_X1 U15507 ( .A1(n12227), .A2(n14021), .ZN(n12223) );
  INV_X1 U15508 ( .A(n18122), .ZN(n12222) );
  NAND2_X1 U15509 ( .A1(n12223), .A2(n12222), .ZN(n12232) );
  NAND2_X1 U15510 ( .A1(n12221), .A2(n12218), .ZN(n12240) );
  INV_X1 U15511 ( .A(n12240), .ZN(n12220) );
  NOR2_X1 U15512 ( .A1(n18110), .A2(n16880), .ZN(n12219) );
  NAND2_X1 U15513 ( .A1(n12220), .A2(n12219), .ZN(n12242) );
  XNOR2_X1 U15514 ( .A(n18113), .B(n12221), .ZN(n12235) );
  AND2_X1 U15515 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n12235), .ZN(
        n12236) );
  OAI21_X1 U15516 ( .B1(n12223), .B2(n12222), .A(n12232), .ZN(n12230) );
  NOR2_X1 U15517 ( .A1(n21349), .A2(n12230), .ZN(n12231) );
  XNOR2_X1 U15518 ( .A(n12227), .B(n12224), .ZN(n12225) );
  NOR2_X1 U15519 ( .A1(n12225), .A2(n18727), .ZN(n12229) );
  NOR2_X1 U15520 ( .A1(n13938), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14187) );
  INV_X1 U15521 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18710) );
  OAI21_X1 U15522 ( .B1(n14187), .B2(n18710), .A(n12226), .ZN(n12228) );
  OAI211_X1 U15523 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n12228), .B(n12227), .ZN(n18484) );
  XOR2_X1 U15524 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n12230), .Z(
        n18475) );
  NOR2_X1 U15525 ( .A1(n18476), .A2(n18475), .ZN(n18474) );
  NOR2_X1 U15526 ( .A1(n12231), .A2(n18474), .ZN(n12233) );
  XNOR2_X1 U15527 ( .A(n18117), .B(n12232), .ZN(n12234) );
  NOR2_X1 U15528 ( .A1(n12233), .A2(n12234), .ZN(n14120) );
  INV_X1 U15529 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18699) );
  INV_X1 U15530 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18691) );
  XOR2_X1 U15531 ( .A(n18691), .B(n12235), .Z(n18463) );
  XNOR2_X1 U15532 ( .A(n18110), .B(n12240), .ZN(n12238) );
  NOR2_X1 U15533 ( .A1(n12237), .A2(n12238), .ZN(n12239) );
  INV_X1 U15534 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14156) );
  OAI21_X1 U15535 ( .B1(n12240), .B2(n18110), .A(n16880), .ZN(n12241) );
  NAND2_X1 U15536 ( .A1(n12242), .A2(n12241), .ZN(n12244) );
  NAND2_X1 U15537 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n14151), .ZN(
        n12246) );
  NOR2_X1 U15538 ( .A1(n12242), .A2(n12246), .ZN(n12248) );
  INV_X1 U15539 ( .A(n12242), .ZN(n12247) );
  OR2_X1 U15540 ( .A1(n12244), .A2(n12243), .ZN(n14152) );
  OAI21_X1 U15541 ( .B1(n12247), .B2(n12246), .A(n14152), .ZN(n12245) );
  AOI21_X1 U15542 ( .B1(n12247), .B2(n12246), .A(n12245), .ZN(n14251) );
  INV_X1 U15543 ( .A(n17044), .ZN(n17064) );
  NOR2_X1 U15544 ( .A1(n17064), .A2(n16895), .ZN(n17247) );
  NAND2_X1 U15545 ( .A1(n17247), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12249) );
  INV_X1 U15546 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n19310) );
  NOR2_X1 U15547 ( .A1(n18739), .A2(n19310), .ZN(n16882) );
  INV_X1 U15548 ( .A(n17027), .ZN(n12252) );
  NAND2_X1 U15549 ( .A1(n18525), .A2(n12252), .ZN(n17065) );
  NOR2_X1 U15550 ( .A1(n17065), .A2(n16895), .ZN(n17260) );
  NAND2_X1 U15551 ( .A1(n17260), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12254) );
  AOI22_X1 U15552 ( .A1(n12254), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        n17260), .B2(n12253), .ZN(n16886) );
  NAND2_X1 U15553 ( .A1(n18653), .A2(n18724), .ZN(n18622) );
  OR2_X1 U15554 ( .A1(n16886), .A2(n18622), .ZN(n12255) );
  NAND2_X1 U15555 ( .A1(n12258), .A2(n12257), .ZN(P3_U2831) );
  NAND2_X1 U15556 ( .A1(n17192), .A2(n13439), .ZN(n12262) );
  AOI21_X1 U15557 ( .B1(n19584), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n12260), .ZN(n12261) );
  NAND2_X1 U15558 ( .A1(n12262), .A2(n12261), .ZN(n12263) );
  AOI21_X1 U15559 ( .B1(n12264), .B2(n9627), .A(n12263), .ZN(n12267) );
  NAND2_X1 U15560 ( .A1(n11082), .A2(n19577), .ZN(n12266) );
  NOR2_X4 U15561 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12276) );
  AOI22_X1 U15562 ( .A1(n12452), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9606), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12275) );
  INV_X1 U15563 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12270) );
  NOR2_X4 U15564 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13968) );
  AOI22_X1 U15565 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12453), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12274) );
  AOI22_X1 U15567 ( .A1(n12469), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12585), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12273) );
  AND2_X2 U15568 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13967) );
  AND2_X4 U15569 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13949) );
  AND2_X2 U15570 ( .A1(n13967), .A2(n13949), .ZN(n12382) );
  AND2_X2 U15571 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13951) );
  AOI22_X1 U15572 ( .A1(n12382), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13504), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12272) );
  AOI22_X1 U15573 ( .A1(n13505), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12383), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12282) );
  AOI22_X1 U15574 ( .A1(n12353), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9609), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12281) );
  AOI22_X1 U15575 ( .A1(n12368), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12358), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12280) );
  INV_X1 U15577 ( .A(n12407), .ZN(n12319) );
  AOI22_X1 U15578 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12453), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12290) );
  AOI22_X1 U15579 ( .A1(n13505), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12383), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12289) );
  AND2_X1 U15580 ( .A1(n9597), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12286) );
  AOI22_X1 U15581 ( .A1(n12451), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12382), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12287) );
  AOI22_X1 U15582 ( .A1(n12461), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12353), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12294) );
  AOI22_X1 U15583 ( .A1(n12469), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12585), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12293) );
  AOI22_X1 U15584 ( .A1(n12368), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12358), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12292) );
  AOI22_X1 U15585 ( .A1(n12452), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12331), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12291) );
  INV_X1 U15586 ( .A(n12417), .ZN(n12318) );
  NAND2_X1 U15587 ( .A1(n12452), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n12300) );
  NAND2_X1 U15588 ( .A1(n12461), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n12299) );
  NAND2_X1 U15589 ( .A1(n12353), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n12298) );
  NAND2_X1 U15590 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12297) );
  NAND2_X1 U15591 ( .A1(n12453), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12304) );
  NAND2_X1 U15592 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n12303) );
  NAND2_X1 U15593 ( .A1(n9614), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n12302) );
  NAND2_X1 U15594 ( .A1(n12383), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n12301) );
  NAND2_X1 U15595 ( .A1(n12368), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n12308) );
  NAND2_X1 U15596 ( .A1(n12469), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n12307) );
  NAND2_X1 U15597 ( .A1(n12585), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12306) );
  NAND2_X1 U15598 ( .A1(n12358), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n12305) );
  NAND2_X1 U15599 ( .A1(n9585), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n12313) );
  NAND2_X1 U15600 ( .A1(n9597), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n12312) );
  INV_X1 U15601 ( .A(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12309) );
  NAND2_X1 U15602 ( .A1(n12382), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n12310) );
  AOI22_X1 U15604 ( .A1(n12461), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12353), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12323) );
  AOI22_X1 U15605 ( .A1(n12469), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12585), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12322) );
  AOI22_X1 U15606 ( .A1(n12452), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12331), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12320) );
  INV_X1 U15607 ( .A(n9604), .ZN(n12324) );
  AOI22_X1 U15608 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12453), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12327) );
  AOI22_X1 U15609 ( .A1(n12451), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12382), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12326) );
  AOI22_X1 U15610 ( .A1(n9614), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12383), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12325) );
  AOI22_X1 U15611 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12353), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12335) );
  AOI22_X1 U15612 ( .A1(n12469), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12585), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12334) );
  AOI22_X1 U15613 ( .A1(n12368), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12358), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12333) );
  AOI22_X1 U15614 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12453), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12338) );
  AOI22_X1 U15615 ( .A1(n9585), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12382), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12337) );
  AOI22_X1 U15616 ( .A1(n13505), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12383), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12336) );
  AOI22_X1 U15617 ( .A1(n12484), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13504), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12339) );
  NAND3_X2 U15618 ( .A1(n12341), .A2(n12340), .A3(n12339), .ZN(n12401) );
  INV_X1 U15619 ( .A(n12415), .ZN(n12367) );
  NAND2_X1 U15620 ( .A1(n12453), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12345) );
  NAND2_X1 U15621 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12344) );
  NAND2_X1 U15622 ( .A1(n9614), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12343) );
  NAND2_X1 U15623 ( .A1(n12383), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12342) );
  NAND2_X1 U15624 ( .A1(n12382), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12346) );
  OAI21_X1 U15625 ( .B1(n13106), .B2(n12347), .A(n12346), .ZN(n12352) );
  INV_X1 U15626 ( .A(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12350) );
  INV_X1 U15627 ( .A(n13504), .ZN(n12349) );
  INV_X1 U15628 ( .A(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12348) );
  NAND2_X1 U15629 ( .A1(n12452), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12357) );
  NAND2_X1 U15630 ( .A1(n12461), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12356) );
  NAND2_X1 U15631 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12354) );
  NAND2_X1 U15632 ( .A1(n12368), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12362) );
  NAND2_X1 U15633 ( .A1(n12469), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12361) );
  NAND2_X1 U15634 ( .A1(n12585), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12360) );
  NAND2_X1 U15635 ( .A1(n12358), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12359) );
  NAND3_X1 U15636 ( .A1(n12380), .A2(n12367), .A3(n14486), .ZN(n14644) );
  INV_X1 U15637 ( .A(n14644), .ZN(n12379) );
  AOI22_X1 U15638 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12453), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12372) );
  AOI22_X1 U15639 ( .A1(n12461), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12353), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12371) );
  AOI22_X1 U15640 ( .A1(n12484), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12331), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12370) );
  AOI22_X1 U15641 ( .A1(n12368), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12358), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12369) );
  AOI22_X1 U15642 ( .A1(n13505), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12383), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12376) );
  AOI22_X1 U15643 ( .A1(n12469), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12585), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12375) );
  AOI22_X1 U15644 ( .A1(n12451), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13504), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12374) );
  AOI22_X1 U15645 ( .A1(n12452), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12382), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12373) );
  NAND2_X1 U15646 ( .A1(n12379), .A2(n12601), .ZN(n13298) );
  AOI22_X1 U15647 ( .A1(n13504), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12382), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12386) );
  AOI22_X1 U15648 ( .A1(n12452), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12331), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12385) );
  AOI22_X1 U15649 ( .A1(n9614), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12383), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12384) );
  AOI22_X1 U15650 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12353), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12395) );
  AOI22_X1 U15651 ( .A1(n12453), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12720), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12393) );
  AOI22_X1 U15652 ( .A1(n12469), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12358), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12392) );
  OAI22_X1 U15653 ( .A1(n13106), .A2(n12389), .B1(n9605), .B2(n12388), .ZN(
        n12390) );
  INV_X1 U15654 ( .A(n12390), .ZN(n12391) );
  NAND2_X1 U15655 ( .A1(n13535), .A2(n13324), .ZN(n12400) );
  NOR2_X1 U15656 ( .A1(n12421), .A2(n12414), .ZN(n12399) );
  INV_X1 U15657 ( .A(n12397), .ZN(n12426) );
  AND3_X2 U15658 ( .A1(n12399), .A2(n12398), .A3(n13538), .ZN(n13305) );
  NAND2_X1 U15659 ( .A1(n13305), .A2(n20603), .ZN(n13539) );
  NOR2_X2 U15660 ( .A1(n14486), .A2(n12441), .ZN(n12437) );
  NAND4_X1 U15661 ( .A1(n12437), .A2(n12403), .A3(n13871), .A4(n13950), .ZN(
        n14500) );
  NAND2_X1 U15662 ( .A1(n13860), .A2(n20622), .ZN(n12405) );
  NAND2_X1 U15663 ( .A1(n13271), .A2(n20615), .ZN(n13857) );
  NAND2_X1 U15664 ( .A1(n12318), .A2(n12407), .ZN(n12438) );
  NAND2_X1 U15665 ( .A1(n12406), .A2(n12408), .ZN(n12409) );
  NAND2_X1 U15666 ( .A1(n13857), .A2(n15582), .ZN(n12413) );
  AND2_X4 U15667 ( .A1(n12414), .A2(n12441), .ZN(n14658) );
  NAND2_X1 U15668 ( .A1(n12401), .A2(n14486), .ZN(n12410) );
  NAND2_X1 U15669 ( .A1(n14487), .A2(n12410), .ZN(n13868) );
  NOR2_X1 U15670 ( .A1(n21216), .A2(n20615), .ZN(n12412) );
  NOR2_X2 U15671 ( .A1(n13868), .A2(n12412), .ZN(n12434) );
  NAND2_X1 U15672 ( .A1(n12413), .A2(n12434), .ZN(n12433) );
  INV_X1 U15673 ( .A(n12414), .ZN(n20611) );
  OAI21_X2 U15674 ( .B1(n12433), .B2(n13864), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n12430) );
  NAND2_X1 U15675 ( .A1(n15582), .A2(n12414), .ZN(n12424) );
  AOI21_X1 U15676 ( .B1(n12420), .B2(n12401), .A(n12421), .ZN(n12422) );
  INV_X1 U15677 ( .A(n13950), .ZN(n13861) );
  NAND2_X1 U15678 ( .A1(n13861), .A2(n20603), .ZN(n12425) );
  NOR2_X1 U15679 ( .A1(n12436), .A2(n12425), .ZN(n12428) );
  NAND2_X1 U15681 ( .A1(n21069), .A2(n20988), .ZN(n20958) );
  NAND2_X1 U15682 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21065) );
  AOI21_X1 U15683 ( .B1(n13275), .B2(n20897), .A(n12510), .ZN(n12431) );
  NAND2_X1 U15684 ( .A1(n12512), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12432) );
  INV_X1 U15685 ( .A(n21134), .ZN(n17146) );
  INV_X1 U15686 ( .A(n13275), .ZN(n12514) );
  MUX2_X1 U15687 ( .A(n17146), .B(n12514), .S(n20988), .Z(n12496) );
  NAND2_X1 U15688 ( .A1(n12434), .A2(n20603), .ZN(n12435) );
  NAND2_X1 U15689 ( .A1(n12433), .A2(n12435), .ZN(n12447) );
  INV_X1 U15690 ( .A(n12437), .ZN(n14640) );
  NAND3_X1 U15691 ( .A1(n14640), .A2(n12438), .A3(n12414), .ZN(n12445) );
  INV_X1 U15692 ( .A(n12439), .ZN(n12440) );
  INV_X1 U15693 ( .A(n21216), .ZN(n13187) );
  NAND2_X1 U15694 ( .A1(n12440), .A2(n13187), .ZN(n12443) );
  NAND2_X1 U15695 ( .A1(n13950), .A2(n20622), .ZN(n14489) );
  AND2_X1 U15696 ( .A1(n15586), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12442) );
  NAND2_X1 U15697 ( .A1(n12427), .A2(n17135), .ZN(n14938) );
  NAND4_X1 U15698 ( .A1(n12443), .A2(n14489), .A3(n12442), .A4(n14938), .ZN(
        n12444) );
  AOI21_X1 U15699 ( .B1(n12436), .B2(n12445), .A(n12444), .ZN(n12446) );
  NAND2_X1 U15700 ( .A1(n12447), .A2(n12446), .ZN(n12665) );
  INV_X1 U15701 ( .A(n20694), .ZN(n12450) );
  AOI22_X1 U15702 ( .A1(n13510), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9623), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12457) );
  AOI22_X1 U15703 ( .A1(n9616), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13511), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12456) );
  AOI22_X1 U15704 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13503), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12454) );
  NAND4_X1 U15705 ( .A1(n12457), .A2(n12456), .A3(n12455), .A4(n12454), .ZN(
        n12467) );
  AOI22_X1 U15706 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13088), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12465) );
  AOI22_X1 U15707 ( .A1(n13043), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9591), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12464) );
  INV_X1 U15708 ( .A(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12459) );
  INV_X1 U15709 ( .A(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12458) );
  OAI22_X1 U15710 ( .A1(n9604), .A2(n12459), .B1(n13108), .B2(n12458), .ZN(
        n12460) );
  INV_X1 U15711 ( .A(n12460), .ZN(n12463) );
  AOI22_X1 U15712 ( .A1(n12461), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12382), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12462) );
  NAND4_X1 U15713 ( .A1(n12465), .A2(n12464), .A3(n12463), .A4(n12462), .ZN(
        n12466) );
  NAND2_X1 U15714 ( .A1(n12483), .A2(n13152), .ZN(n12468) );
  AOI22_X1 U15715 ( .A1(n9617), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n13088), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12476) );
  AOI22_X1 U15716 ( .A1(n12461), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12353), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12475) );
  AOI22_X1 U15717 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12469), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12474) );
  INV_X1 U15718 ( .A(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12471) );
  INV_X1 U15719 ( .A(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12470) );
  OAI22_X1 U15720 ( .A1(n13106), .A2(n12471), .B1(n9605), .B2(n12470), .ZN(
        n12472) );
  INV_X1 U15721 ( .A(n12472), .ZN(n12473) );
  NAND4_X1 U15722 ( .A1(n12476), .A2(n12475), .A3(n12474), .A4(n12473), .ZN(
        n12482) );
  AOI22_X1 U15723 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13511), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12480) );
  AOI22_X1 U15724 ( .A1(n12585), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13503), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12479) );
  AOI22_X1 U15725 ( .A1(n9623), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13068), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12478) );
  AOI22_X1 U15726 ( .A1(n13504), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12382), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12477) );
  NAND4_X1 U15727 ( .A1(n12480), .A2(n12479), .A3(n12478), .A4(n12477), .ZN(
        n12481) );
  INV_X1 U15728 ( .A(n13186), .ZN(n13195) );
  NAND2_X1 U15729 ( .A1(n12483), .A2(n13195), .ZN(n12504) );
  AOI22_X1 U15730 ( .A1(n13511), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13088), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12488) );
  AOI22_X1 U15731 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n13512), .B1(
        n9617), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12487) );
  AOI22_X1 U15732 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n9623), .B1(
        n13043), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12486) );
  AOI22_X1 U15733 ( .A1(n13504), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13016), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12485) );
  NAND4_X1 U15734 ( .A1(n12488), .A2(n12487), .A3(n12486), .A4(n12485), .ZN(
        n12494) );
  AOI22_X1 U15735 ( .A1(n13510), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13502), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12492) );
  AOI22_X1 U15736 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n13513), .B1(
        n13503), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12490) );
  AOI22_X1 U15737 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13068), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12489) );
  NAND4_X1 U15738 ( .A1(n12492), .A2(n12491), .A3(n12490), .A4(n12489), .ZN(
        n12493) );
  INV_X1 U15739 ( .A(n13158), .ZN(n12495) );
  NAND2_X1 U15740 ( .A1(n12496), .A2(n10368), .ZN(n12497) );
  INV_X1 U15741 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12501) );
  AOI21_X1 U15742 ( .B1(n20615), .B2(n13186), .A(n10368), .ZN(n12500) );
  NAND2_X1 U15743 ( .A1(n12427), .A2(n13158), .ZN(n12499) );
  NAND2_X1 U15744 ( .A1(n12675), .A2(n12674), .ZN(n12502) );
  INV_X1 U15745 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13018) );
  INV_X1 U15746 ( .A(n12544), .ZN(n12537) );
  NAND2_X1 U15747 ( .A1(n12537), .A2(n13152), .ZN(n12503) );
  INV_X1 U15748 ( .A(n12505), .ZN(n12508) );
  INV_X1 U15749 ( .A(n12506), .ZN(n12507) );
  NAND2_X1 U15750 ( .A1(n12508), .A2(n12507), .ZN(n12509) );
  INV_X1 U15751 ( .A(n12510), .ZN(n12511) );
  NAND2_X1 U15752 ( .A1(n12521), .A2(n12518), .ZN(n12517) );
  BUF_X1 U15753 ( .A(n12512), .Z(n12513) );
  XNOR2_X1 U15754 ( .A(n21065), .B(n20840), .ZN(n20597) );
  NOR2_X1 U15755 ( .A1(n20597), .A2(n12514), .ZN(n12515) );
  NAND2_X1 U15756 ( .A1(n21134), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12519) );
  NAND2_X1 U15757 ( .A1(n12520), .A2(n12519), .ZN(n12516) );
  AOI22_X1 U15758 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13511), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12529) );
  AOI22_X1 U15759 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13088), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12528) );
  AOI22_X1 U15760 ( .A1(n13510), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12382), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12527) );
  INV_X1 U15761 ( .A(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12524) );
  INV_X1 U15762 ( .A(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12523) );
  OAI22_X1 U15763 ( .A1(n9605), .A2(n12524), .B1(n13108), .B2(n12523), .ZN(
        n12525) );
  INV_X1 U15764 ( .A(n12525), .ZN(n12526) );
  NAND4_X1 U15765 ( .A1(n12529), .A2(n12528), .A3(n12527), .A4(n12526), .ZN(
        n12535) );
  AOI22_X1 U15766 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10147), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12533) );
  AOI22_X1 U15767 ( .A1(n13043), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12953), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12532) );
  AOI22_X1 U15768 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13503), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12531) );
  AOI22_X1 U15769 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13068), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12530) );
  NAND4_X1 U15770 ( .A1(n12533), .A2(n12532), .A3(n12531), .A4(n12530), .ZN(
        n12534) );
  AOI22_X1 U15771 ( .A1(n12537), .A2(n12536), .B1(n13260), .B2(
        P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12538) );
  INV_X1 U15772 ( .A(n12678), .ZN(n12559) );
  NAND2_X1 U15773 ( .A1(n12513), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12542) );
  OAI21_X1 U15774 ( .B1(n21065), .B2(n20840), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12540) );
  INV_X1 U15775 ( .A(n21065), .ZN(n17118) );
  NAND2_X1 U15776 ( .A1(n20589), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20778) );
  INV_X1 U15777 ( .A(n20778), .ZN(n12539) );
  NAND2_X1 U15778 ( .A1(n17118), .A2(n12539), .ZN(n20808) );
  NAND2_X1 U15779 ( .A1(n12540), .A2(n20808), .ZN(n20841) );
  AOI22_X1 U15780 ( .A1(n13275), .A2(n20841), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n21134), .ZN(n12541) );
  AOI22_X1 U15781 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13511), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12551) );
  AOI22_X1 U15782 ( .A1(n9584), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13088), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12550) );
  AOI22_X1 U15783 ( .A1(n13510), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13016), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12549) );
  INV_X1 U15784 ( .A(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12546) );
  INV_X1 U15785 ( .A(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12545) );
  OAI22_X1 U15786 ( .A1(n9604), .A2(n12546), .B1(n13108), .B2(n12545), .ZN(
        n12547) );
  INV_X1 U15787 ( .A(n12547), .ZN(n12548) );
  NAND4_X1 U15788 ( .A1(n12551), .A2(n12550), .A3(n12549), .A4(n12548), .ZN(
        n12557) );
  AOI22_X1 U15789 ( .A1(n12461), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10147), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12555) );
  AOI22_X1 U15790 ( .A1(n13043), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12953), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12554) );
  AOI22_X1 U15791 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13503), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12553) );
  AOI22_X1 U15792 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13068), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12552) );
  NAND4_X1 U15793 ( .A1(n12555), .A2(n12554), .A3(n12553), .A4(n12552), .ZN(
        n12556) );
  AOI22_X1 U15794 ( .A1(n13248), .A2(n13140), .B1(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n13260), .ZN(n12558) );
  AOI22_X1 U15795 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13088), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12563) );
  AOI22_X1 U15796 ( .A1(n13510), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13016), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12561) );
  AOI22_X1 U15797 ( .A1(n9584), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13504), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12560) );
  NAND4_X1 U15798 ( .A1(n12563), .A2(n12562), .A3(n12561), .A4(n12560), .ZN(
        n12569) );
  AOI22_X1 U15799 ( .A1(n13512), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13511), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12567) );
  AOI22_X1 U15800 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12953), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12566) );
  AOI22_X1 U15801 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13503), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12565) );
  AOI22_X1 U15802 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13068), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12564) );
  NAND4_X1 U15803 ( .A1(n12567), .A2(n12566), .A3(n12565), .A4(n12564), .ZN(
        n12568) );
  AOI22_X1 U15804 ( .A1(n13248), .A2(n13136), .B1(
        P1_INSTQUEUE_REG_0__4__SCAN_IN), .B2(n13260), .ZN(n12689) );
  AOI22_X1 U15805 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13511), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12576) );
  AOI22_X1 U15806 ( .A1(n9618), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13088), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12575) );
  INV_X1 U15807 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13109) );
  AOI22_X1 U15808 ( .A1(n13510), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13016), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12574) );
  INV_X1 U15809 ( .A(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12571) );
  INV_X1 U15810 ( .A(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12570) );
  OAI22_X1 U15811 ( .A1(n9605), .A2(n12571), .B1(n13108), .B2(n12570), .ZN(
        n12572) );
  INV_X1 U15812 ( .A(n12572), .ZN(n12573) );
  NAND4_X1 U15813 ( .A1(n12576), .A2(n12575), .A3(n12574), .A4(n12573), .ZN(
        n12582) );
  AOI22_X1 U15814 ( .A1(n13043), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12953), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12579) );
  AOI22_X1 U15815 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13503), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12578) );
  AOI22_X1 U15816 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13068), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12577) );
  NAND4_X1 U15817 ( .A1(n12580), .A2(n12579), .A3(n12578), .A4(n12577), .ZN(
        n12581) );
  NAND2_X1 U15818 ( .A1(n13248), .A2(n13173), .ZN(n12584) );
  NAND2_X1 U15819 ( .A1(n13260), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12583) );
  NAND2_X1 U15820 ( .A1(n12584), .A2(n12583), .ZN(n12609) );
  AOI22_X1 U15821 ( .A1(n13510), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9620), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12589) );
  AOI22_X1 U15822 ( .A1(n13511), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13088), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12588) );
  AOI22_X1 U15823 ( .A1(n12461), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12953), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12587) );
  AOI22_X1 U15824 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13503), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12586) );
  NAND4_X1 U15825 ( .A1(n12589), .A2(n12588), .A3(n12587), .A4(n12586), .ZN(
        n12595) );
  AOI22_X1 U15826 ( .A1(n13512), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12720), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12593) );
  AOI22_X1 U15827 ( .A1(n13504), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13016), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12591) );
  AOI22_X1 U15828 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13068), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12590) );
  NAND4_X1 U15829 ( .A1(n12593), .A2(n12592), .A3(n12591), .A4(n12590), .ZN(
        n12594) );
  NAND2_X1 U15830 ( .A1(n13248), .A2(n13184), .ZN(n12597) );
  NAND2_X1 U15831 ( .A1(n13260), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12596) );
  NAND2_X1 U15832 ( .A1(n12597), .A2(n12596), .ZN(n12619) );
  INV_X1 U15833 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12599) );
  NAND2_X1 U15834 ( .A1(n13248), .A2(n13186), .ZN(n12598) );
  OAI21_X1 U15835 ( .B1(n12599), .B2(n13243), .A(n12598), .ZN(n12600) );
  NAND2_X1 U15836 ( .A1(n13182), .A2(n12823), .ZN(n12608) );
  INV_X1 U15837 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12605) );
  NAND2_X1 U15838 ( .A1(n21070), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12627) );
  INV_X1 U15839 ( .A(n12683), .ZN(n12602) );
  OAI21_X1 U15840 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n12623), .A(
        n12642), .ZN(n20387) );
  INV_X2 U15841 ( .A(n13524), .ZN(n13531) );
  NAND2_X1 U15842 ( .A1(n20387), .A2(n13531), .ZN(n12604) );
  OAI21_X1 U15843 ( .B1(n12605), .B2(n12627), .A(n12604), .ZN(n12606) );
  AOI21_X1 U15844 ( .B1(n13032), .B2(P1_EAX_REG_7__SCAN_IN), .A(n12606), .ZN(
        n12607) );
  NAND2_X1 U15845 ( .A1(n12608), .A2(n12607), .ZN(n14460) );
  NAND2_X1 U15846 ( .A1(n13130), .A2(n12823), .ZN(n12618) );
  INV_X1 U15847 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12612) );
  NAND2_X1 U15848 ( .A1(n12698), .A2(n12612), .ZN(n12613) );
  NAND2_X1 U15849 ( .A1(n12622), .A2(n12613), .ZN(n20415) );
  NAND2_X1 U15850 ( .A1(n20415), .A2(n13531), .ZN(n12615) );
  NAND2_X1 U15851 ( .A1(n13532), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12614) );
  NAND2_X1 U15852 ( .A1(n12615), .A2(n12614), .ZN(n12616) );
  AOI21_X1 U15853 ( .B1(n13032), .B2(P1_EAX_REG_5__SCAN_IN), .A(n12616), .ZN(
        n12617) );
  INV_X1 U15854 ( .A(n12619), .ZN(n12620) );
  NAND2_X1 U15855 ( .A1(n12621), .A2(n12620), .ZN(n13171) );
  NAND2_X1 U15856 ( .A1(n13171), .A2(n12823), .ZN(n12631) );
  NAND2_X1 U15857 ( .A1(n12622), .A2(n12628), .ZN(n12625) );
  INV_X1 U15858 ( .A(n12623), .ZN(n12624) );
  NAND2_X1 U15859 ( .A1(n12625), .A2(n12624), .ZN(n20402) );
  NAND2_X1 U15860 ( .A1(n20402), .A2(n13531), .ZN(n12626) );
  OAI21_X1 U15861 ( .B1(n12628), .B2(n12627), .A(n12626), .ZN(n12629) );
  AOI21_X1 U15862 ( .B1(n13032), .B2(P1_EAX_REG_6__SCAN_IN), .A(n12629), .ZN(
        n12630) );
  NAND2_X1 U15863 ( .A1(n12631), .A2(n12630), .ZN(n14445) );
  AOI22_X1 U15864 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13088), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12635) );
  AOI22_X1 U15865 ( .A1(n13512), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9621), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12634) );
  AOI22_X1 U15866 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n12953), .B1(
        n13503), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12632) );
  NAND4_X1 U15867 ( .A1(n12635), .A2(n12634), .A3(n12633), .A4(n12632), .ZN(
        n12641) );
  AOI22_X1 U15868 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n13513), .B1(
        n9607), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12639) );
  AOI22_X1 U15869 ( .A1(n13510), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        P1_INSTQUEUE_REG_1__0__SCAN_IN), .B2(n13016), .ZN(n12638) );
  AOI22_X1 U15870 ( .A1(n13511), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13504), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12637) );
  AOI22_X1 U15871 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13068), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12636) );
  NAND4_X1 U15872 ( .A1(n12639), .A2(n12638), .A3(n12637), .A4(n12636), .ZN(
        n12640) );
  NOR2_X1 U15873 ( .A1(n12641), .A2(n12640), .ZN(n12645) );
  INV_X1 U15874 ( .A(n12823), .ZN(n12791) );
  NAND2_X1 U15875 ( .A1(n13032), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n12644) );
  XNOR2_X1 U15876 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n12715), .ZN(
        n20369) );
  AOI22_X1 U15877 ( .A1(n13531), .A2(n20369), .B1(n13532), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12643) );
  OAI211_X1 U15878 ( .C1(n12645), .C2(n12791), .A(n12644), .B(n12643), .ZN(
        n14462) );
  NAND2_X1 U15879 ( .A1(n13145), .A2(n12823), .ZN(n12654) );
  NAND2_X1 U15880 ( .A1(n13871), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12694) );
  XNOR2_X1 U15881 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14951) );
  AOI21_X1 U15882 ( .B1(n13531), .B2(n14951), .A(n13532), .ZN(n12651) );
  NAND2_X1 U15883 ( .A1(n13032), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n12650) );
  OAI211_X1 U15884 ( .C1(n12694), .C2(n12649), .A(n12651), .B(n12650), .ZN(
        n12652) );
  INV_X1 U15885 ( .A(n12652), .ZN(n12653) );
  NAND2_X1 U15886 ( .A1(n13532), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12677) );
  NAND2_X1 U15887 ( .A1(n20662), .A2(n12823), .ZN(n12664) );
  NAND2_X1 U15888 ( .A1(n13032), .A2(P1_EAX_REG_1__SCAN_IN), .ZN(n12661) );
  NAND2_X1 U15889 ( .A1(n21070), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12660) );
  OAI211_X1 U15890 ( .C1(n12694), .C2(n13215), .A(n12661), .B(n12660), .ZN(
        n12662) );
  INV_X1 U15891 ( .A(n12662), .ZN(n12663) );
  INV_X1 U15892 ( .A(n12665), .ZN(n12666) );
  XNOR2_X1 U15893 ( .A(n12667), .B(n12666), .ZN(n21386) );
  NAND2_X1 U15894 ( .A1(n21386), .A2(n12823), .ZN(n12673) );
  AOI22_X1 U15895 ( .A1(n12668), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n21070), .ZN(n12671) );
  INV_X1 U15896 ( .A(n12694), .ZN(n12669) );
  NAND2_X1 U15897 ( .A1(n12669), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12670) );
  AND2_X1 U15898 ( .A1(n12671), .A2(n12670), .ZN(n12672) );
  NAND2_X1 U15899 ( .A1(n12673), .A2(n12672), .ZN(n13919) );
  AOI21_X1 U15900 ( .B1(n20661), .B2(n20622), .A(n21070), .ZN(n13918) );
  NAND2_X1 U15901 ( .A1(n13919), .A2(n13918), .ZN(n13917) );
  OR2_X1 U15902 ( .A1(n13919), .A2(n13524), .ZN(n12676) );
  NAND2_X1 U15903 ( .A1(n13917), .A2(n12676), .ZN(n14145) );
  INV_X1 U15904 ( .A(n12682), .ZN(n12695) );
  INV_X1 U15905 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n21271) );
  NAND2_X1 U15906 ( .A1(n21271), .A2(n12683), .ZN(n12684) );
  NAND2_X1 U15907 ( .A1(n12695), .A2(n12684), .ZN(n14942) );
  AOI22_X1 U15908 ( .A1(n14942), .A2(n13531), .B1(n13532), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12686) );
  NAND2_X1 U15909 ( .A1(n13032), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n12685) );
  OAI211_X1 U15910 ( .C1(n12694), .C2(n12681), .A(n12686), .B(n12685), .ZN(
        n12687) );
  INV_X1 U15911 ( .A(n12687), .ZN(n12688) );
  INV_X1 U15912 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n12693) );
  NAND2_X1 U15913 ( .A1(n21070), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12692) );
  NAND2_X1 U15914 ( .A1(n13032), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n12691) );
  OAI211_X1 U15915 ( .C1(n12694), .C2(n12693), .A(n12692), .B(n12691), .ZN(
        n12699) );
  INV_X1 U15916 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n12696) );
  NAND2_X1 U15917 ( .A1(n12696), .A2(n12695), .ZN(n12697) );
  NAND2_X1 U15918 ( .A1(n12698), .A2(n12697), .ZN(n20522) );
  MUX2_X1 U15919 ( .A(n12699), .B(n20522), .S(n13531), .Z(n12700) );
  AOI22_X1 U15920 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13088), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12705) );
  AOI22_X1 U15921 ( .A1(n13510), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13068), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12704) );
  AOI22_X1 U15922 ( .A1(n12461), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12953), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12703) );
  AOI22_X1 U15923 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13503), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12702) );
  NAND4_X1 U15924 ( .A1(n12705), .A2(n12704), .A3(n12703), .A4(n12702), .ZN(
        n12714) );
  AOI22_X1 U15925 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13511), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12712) );
  INV_X1 U15926 ( .A(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12707) );
  INV_X1 U15927 ( .A(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12706) );
  OAI22_X1 U15928 ( .A1(n9605), .A2(n12707), .B1(n13108), .B2(n12706), .ZN(
        n12708) );
  INV_X1 U15929 ( .A(n12708), .ZN(n12710) );
  AOI22_X1 U15930 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13016), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12709) );
  NAND4_X1 U15931 ( .A1(n12712), .A2(n12711), .A3(n12710), .A4(n12709), .ZN(
        n12713) );
  OAI21_X1 U15932 ( .B1(n12714), .B2(n12713), .A(n12823), .ZN(n12718) );
  NAND2_X1 U15933 ( .A1(n13032), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n12717) );
  XNOR2_X1 U15934 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n12734), .ZN(
        n20359) );
  AOI22_X1 U15935 ( .A1(n13531), .A2(n20359), .B1(n13532), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12716) );
  AOI22_X1 U15936 ( .A1(n13502), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13088), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12724) );
  AOI22_X1 U15937 ( .A1(n13510), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13068), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12722) );
  AOI22_X1 U15938 ( .A1(n13043), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13503), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12721) );
  NAND4_X1 U15939 ( .A1(n12724), .A2(n12723), .A3(n12722), .A4(n12721), .ZN(
        n12733) );
  AOI22_X1 U15940 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13511), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12731) );
  AOI22_X1 U15941 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12953), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12730) );
  INV_X1 U15942 ( .A(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12726) );
  INV_X1 U15943 ( .A(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12725) );
  OAI22_X1 U15944 ( .A1(n9604), .A2(n12726), .B1(n13108), .B2(n12725), .ZN(
        n12727) );
  INV_X1 U15945 ( .A(n12727), .ZN(n12729) );
  AOI22_X1 U15946 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13016), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12728) );
  NAND4_X1 U15947 ( .A1(n12731), .A2(n12730), .A3(n12729), .A4(n12728), .ZN(
        n12732) );
  OAI21_X1 U15948 ( .B1(n12733), .B2(n12732), .A(n12823), .ZN(n12738) );
  NAND2_X1 U15949 ( .A1(n12668), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n12737) );
  INV_X1 U15950 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12735) );
  XNOR2_X1 U15951 ( .A(n12741), .B(n12735), .ZN(n15297) );
  AOI22_X1 U15952 ( .A1(n15297), .A2(n13531), .B1(n13532), .B2(
        P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12736) );
  NAND2_X1 U15953 ( .A1(n13032), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n12748) );
  INV_X1 U15954 ( .A(n12743), .ZN(n12745) );
  INV_X1 U15955 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12744) );
  NAND2_X1 U15956 ( .A1(n12745), .A2(n12744), .ZN(n12746) );
  NAND2_X1 U15957 ( .A1(n12826), .A2(n12746), .ZN(n15285) );
  AOI22_X1 U15958 ( .A1(n15285), .A2(n13531), .B1(n13532), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12747) );
  NAND2_X1 U15959 ( .A1(n12748), .A2(n12747), .ZN(n14874) );
  AOI22_X1 U15960 ( .A1(n13502), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13511), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12752) );
  AOI22_X1 U15961 ( .A1(n13510), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9616), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12751) );
  AOI22_X1 U15962 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13043), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12749) );
  NAND4_X1 U15963 ( .A1(n12752), .A2(n12751), .A3(n12750), .A4(n12749), .ZN(
        n12758) );
  AOI22_X1 U15964 ( .A1(n13512), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13088), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12756) );
  AOI22_X1 U15965 ( .A1(n12953), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13503), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12755) );
  AOI22_X1 U15966 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13068), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12754) );
  AOI22_X1 U15967 ( .A1(n13504), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13016), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12753) );
  NAND4_X1 U15968 ( .A1(n12756), .A2(n12755), .A3(n12754), .A4(n12753), .ZN(
        n12757) );
  NOR2_X1 U15969 ( .A1(n12758), .A2(n12757), .ZN(n12759) );
  NOR2_X1 U15970 ( .A1(n12791), .A2(n12759), .ZN(n14918) );
  AOI22_X1 U15971 ( .A1(n13502), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13511), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12763) );
  AOI22_X1 U15972 ( .A1(n13512), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13088), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12762) );
  AOI22_X1 U15973 ( .A1(n13510), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13068), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12761) );
  AOI22_X1 U15974 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12953), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12760) );
  NAND4_X1 U15975 ( .A1(n12763), .A2(n12762), .A3(n12761), .A4(n12760), .ZN(
        n12769) );
  AOI22_X1 U15976 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13503), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12766) );
  AOI22_X1 U15977 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13504), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12765) );
  AOI22_X1 U15978 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13016), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12764) );
  NAND4_X1 U15979 ( .A1(n12767), .A2(n12766), .A3(n12765), .A4(n12764), .ZN(
        n12768) );
  OAI21_X1 U15980 ( .B1(n12769), .B2(n12768), .A(n12823), .ZN(n12775) );
  NAND2_X1 U15981 ( .A1(n13032), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n12774) );
  NAND2_X1 U15982 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12770) );
  INV_X1 U15983 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12771) );
  XNOR2_X1 U15984 ( .A(n12854), .B(n12771), .ZN(n15245) );
  NAND2_X1 U15985 ( .A1(n15245), .A2(n13531), .ZN(n12773) );
  NAND2_X1 U15986 ( .A1(n13532), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12772) );
  NAND4_X1 U15987 ( .A1(n12775), .A2(n12774), .A3(n12773), .A4(n12772), .ZN(
        n14851) );
  AOI22_X1 U15988 ( .A1(n9584), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13088), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12779) );
  AOI22_X1 U15989 ( .A1(n13510), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13068), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12777) );
  AOI22_X1 U15990 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12953), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12776) );
  NAND4_X1 U15991 ( .A1(n12779), .A2(n12778), .A3(n12777), .A4(n12776), .ZN(
        n12787) );
  AOI22_X1 U15992 ( .A1(n13502), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13511), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12785) );
  AOI22_X1 U15993 ( .A1(n12461), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13503), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12784) );
  INV_X1 U15994 ( .A(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12780) );
  INV_X1 U15995 ( .A(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12931) );
  OAI22_X1 U15996 ( .A1(n9605), .A2(n12780), .B1(n13108), .B2(n12931), .ZN(
        n12781) );
  INV_X1 U15997 ( .A(n12781), .ZN(n12783) );
  AOI22_X1 U15998 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13016), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12782) );
  NAND4_X1 U15999 ( .A1(n12785), .A2(n12784), .A3(n12783), .A4(n12782), .ZN(
        n12786) );
  NOR2_X1 U16000 ( .A1(n12787), .A2(n12786), .ZN(n12792) );
  NAND2_X1 U16001 ( .A1(n13032), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n12790) );
  INV_X1 U16002 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12788) );
  XNOR2_X1 U16003 ( .A(n12826), .B(n12788), .ZN(n15276) );
  AOI22_X1 U16004 ( .A1(n15276), .A2(n13531), .B1(n13532), .B2(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12789) );
  OAI211_X1 U16005 ( .C1(n12792), .C2(n12791), .A(n12790), .B(n12789), .ZN(
        n14893) );
  OAI211_X1 U16006 ( .C1(n14874), .C2(n14918), .A(n14851), .B(n14893), .ZN(
        n12835) );
  AOI22_X1 U16007 ( .A1(n13502), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9620), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12796) );
  AOI22_X1 U16008 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12461), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12795) );
  AOI22_X1 U16009 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12953), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12793) );
  NAND4_X1 U16010 ( .A1(n12796), .A2(n12795), .A3(n12794), .A4(n12793), .ZN(
        n12804) );
  AOI22_X1 U16011 ( .A1(n13511), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13088), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12802) );
  AOI22_X1 U16012 ( .A1(n13510), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13016), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12801) );
  INV_X1 U16013 ( .A(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12797) );
  INV_X1 U16014 ( .A(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12951) );
  OAI22_X1 U16015 ( .A1(n9604), .A2(n12797), .B1(n13108), .B2(n12951), .ZN(
        n12798) );
  INV_X1 U16016 ( .A(n12798), .ZN(n12800) );
  AOI22_X1 U16017 ( .A1(n13503), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13068), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12799) );
  NAND4_X1 U16018 ( .A1(n12802), .A2(n12801), .A3(n12800), .A4(n12799), .ZN(
        n12803) );
  OAI21_X1 U16019 ( .B1(n12804), .B2(n12803), .A(n12823), .ZN(n12811) );
  NAND2_X1 U16020 ( .A1(n13032), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n12810) );
  INV_X1 U16021 ( .A(n12805), .ZN(n12807) );
  INV_X1 U16022 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12806) );
  XNOR2_X1 U16023 ( .A(n12807), .B(n12806), .ZN(n15254) );
  NAND2_X1 U16024 ( .A1(n15254), .A2(n13531), .ZN(n12809) );
  NAND2_X1 U16025 ( .A1(n13532), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12808) );
  NAND4_X1 U16026 ( .A1(n12811), .A2(n12810), .A3(n12809), .A4(n12808), .ZN(
        n14865) );
  AOI22_X1 U16027 ( .A1(n13502), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13511), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12815) );
  AOI22_X1 U16028 ( .A1(n13043), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12953), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12813) );
  AOI22_X1 U16029 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13068), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12812) );
  NAND4_X1 U16030 ( .A1(n12815), .A2(n12814), .A3(n12813), .A4(n12812), .ZN(
        n12825) );
  AOI22_X1 U16031 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13088), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12822) );
  AOI22_X1 U16032 ( .A1(n13510), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13016), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12821) );
  AOI22_X1 U16033 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13503), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12820) );
  INV_X1 U16034 ( .A(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12817) );
  INV_X1 U16035 ( .A(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12816) );
  OAI22_X1 U16036 ( .A1(n9605), .A2(n12817), .B1(n13108), .B2(n12816), .ZN(
        n12818) );
  INV_X1 U16037 ( .A(n12818), .ZN(n12819) );
  NAND4_X1 U16038 ( .A1(n12822), .A2(n12821), .A3(n12820), .A4(n12819), .ZN(
        n12824) );
  OAI21_X1 U16039 ( .B1(n12825), .B2(n12824), .A(n12823), .ZN(n12833) );
  NAND2_X1 U16040 ( .A1(n13032), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n12832) );
  NAND2_X1 U16041 ( .A1(n13532), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12831) );
  INV_X1 U16042 ( .A(n12826), .ZN(n12827) );
  NAND2_X1 U16043 ( .A1(n12827), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12829) );
  INV_X1 U16044 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12828) );
  XNOR2_X1 U16045 ( .A(n12829), .B(n12828), .ZN(n15269) );
  NAND2_X1 U16046 ( .A1(n15269), .A2(n13531), .ZN(n12830) );
  NAND4_X1 U16047 ( .A1(n12833), .A2(n12832), .A3(n12831), .A4(n12830), .ZN(
        n14877) );
  NAND2_X1 U16048 ( .A1(n14865), .A2(n14877), .ZN(n12834) );
  INV_X1 U16049 ( .A(n15582), .ZN(n14024) );
  AOI22_X1 U16050 ( .A1(n13512), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9623), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12840) );
  AOI22_X1 U16051 ( .A1(n13511), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13088), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12839) );
  AOI22_X1 U16052 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n13513), .B1(
        n9591), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12838) );
  NAND4_X1 U16053 ( .A1(n12840), .A2(n12839), .A3(n12838), .A4(n12837), .ZN(
        n12849) );
  AOI22_X1 U16054 ( .A1(n13502), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9620), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12847) );
  INV_X1 U16055 ( .A(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12842) );
  INV_X1 U16056 ( .A(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12841) );
  OAI22_X1 U16057 ( .A1(n13106), .A2(n12842), .B1(n13108), .B2(n12841), .ZN(
        n12843) );
  INV_X1 U16058 ( .A(n12843), .ZN(n12846) );
  AOI22_X1 U16059 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n13043), .B1(
        n13503), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12845) );
  AOI22_X1 U16060 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13016), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12844) );
  NAND4_X1 U16061 ( .A1(n12847), .A2(n12846), .A3(n12845), .A4(n12844), .ZN(
        n12848) );
  NOR2_X1 U16062 ( .A1(n12849), .A2(n12848), .ZN(n12853) );
  NAND2_X1 U16063 ( .A1(n21070), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12850) );
  NAND2_X1 U16064 ( .A1(n13524), .A2(n12850), .ZN(n12851) );
  AOI21_X1 U16065 ( .B1(n13032), .B2(P1_EAX_REG_16__SCAN_IN), .A(n12851), .ZN(
        n12852) );
  OAI21_X1 U16066 ( .B1(n13078), .B2(n12853), .A(n12852), .ZN(n12861) );
  INV_X1 U16067 ( .A(n12856), .ZN(n12858) );
  INV_X1 U16068 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n12857) );
  NAND2_X1 U16069 ( .A1(n12858), .A2(n12857), .ZN(n12859) );
  NAND2_X1 U16070 ( .A1(n12897), .A2(n12859), .ZN(n15236) );
  OR2_X1 U16071 ( .A1(n15236), .A2(n13524), .ZN(n12860) );
  AOI22_X1 U16072 ( .A1(n13502), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13511), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12865) );
  AOI22_X1 U16073 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13088), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12864) );
  AOI22_X1 U16074 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13068), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12863) );
  AOI22_X1 U16075 ( .A1(n12953), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13503), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12862) );
  NAND4_X1 U16076 ( .A1(n12865), .A2(n12864), .A3(n12863), .A4(n12862), .ZN(
        n12874) );
  AOI22_X1 U16077 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13043), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12871) );
  AOI22_X1 U16078 ( .A1(n13510), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13016), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12870) );
  INV_X1 U16079 ( .A(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12867) );
  INV_X1 U16080 ( .A(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12866) );
  OAI22_X1 U16081 ( .A1(n9605), .A2(n12867), .B1(n13108), .B2(n12866), .ZN(
        n12868) );
  INV_X1 U16082 ( .A(n12868), .ZN(n12869) );
  NAND4_X1 U16083 ( .A1(n12872), .A2(n12871), .A3(n12870), .A4(n12869), .ZN(
        n12873) );
  OAI21_X1 U16084 ( .B1(n12874), .B2(n12873), .A(n13528), .ZN(n12878) );
  AOI22_X1 U16085 ( .A1(n13032), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n13532), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12877) );
  INV_X1 U16086 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12875) );
  XNOR2_X1 U16087 ( .A(n12897), .B(n12875), .ZN(n15225) );
  NAND2_X1 U16088 ( .A1(n15225), .A2(n13531), .ZN(n12876) );
  AOI22_X1 U16089 ( .A1(n13510), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9624), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12883) );
  AOI22_X1 U16090 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13511), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12882) );
  AOI22_X1 U16091 ( .A1(n12953), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13068), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12881) );
  AOI22_X1 U16092 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13503), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12880) );
  NAND4_X1 U16093 ( .A1(n12883), .A2(n12882), .A3(n12881), .A4(n12880), .ZN(
        n12892) );
  AOI22_X1 U16094 ( .A1(n13502), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13088), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12890) );
  INV_X1 U16095 ( .A(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12885) );
  INV_X1 U16096 ( .A(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12884) );
  OAI22_X1 U16097 ( .A1(n9605), .A2(n12885), .B1(n13108), .B2(n12884), .ZN(
        n12886) );
  INV_X1 U16098 ( .A(n12886), .ZN(n12888) );
  AOI22_X1 U16099 ( .A1(n12461), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13016), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12887) );
  NAND4_X1 U16100 ( .A1(n12890), .A2(n12889), .A3(n12888), .A4(n12887), .ZN(
        n12891) );
  NOR2_X1 U16101 ( .A1(n12892), .A2(n12891), .ZN(n12896) );
  OAI21_X1 U16102 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n21022), .A(
        n21070), .ZN(n12893) );
  INV_X1 U16103 ( .A(n12893), .ZN(n12894) );
  AOI21_X1 U16104 ( .B1(n13032), .B2(P1_EAX_REG_18__SCAN_IN), .A(n12894), .ZN(
        n12895) );
  OAI21_X1 U16105 ( .B1(n13078), .B2(n12896), .A(n12895), .ZN(n12904) );
  INV_X1 U16106 ( .A(n12899), .ZN(n12901) );
  INV_X1 U16107 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n12900) );
  NAND2_X1 U16108 ( .A1(n12901), .A2(n12900), .ZN(n12902) );
  NAND2_X1 U16109 ( .A1(n12923), .A2(n12902), .ZN(n15206) );
  NAND2_X1 U16110 ( .A1(n12904), .A2(n12903), .ZN(n14800) );
  XNOR2_X1 U16111 ( .A(n12923), .B(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15199) );
  NAND2_X1 U16112 ( .A1(n15199), .A2(n13531), .ZN(n12922) );
  AOI22_X1 U16113 ( .A1(n13502), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13511), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12911) );
  AOI22_X1 U16114 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13088), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12910) );
  AOI22_X1 U16115 ( .A1(n13510), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13016), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12909) );
  INV_X1 U16116 ( .A(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12906) );
  INV_X1 U16117 ( .A(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12905) );
  OAI22_X1 U16118 ( .A1(n9604), .A2(n12906), .B1(n13108), .B2(n12905), .ZN(
        n12907) );
  INV_X1 U16119 ( .A(n12907), .ZN(n12908) );
  NAND4_X1 U16120 ( .A1(n12911), .A2(n12910), .A3(n12909), .A4(n12908), .ZN(
        n12917) );
  AOI22_X1 U16121 ( .A1(n13043), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9591), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12914) );
  AOI22_X1 U16122 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13503), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12913) );
  AOI22_X1 U16123 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13068), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12912) );
  NAND4_X1 U16124 ( .A1(n12915), .A2(n12914), .A3(n12913), .A4(n12912), .ZN(
        n12916) );
  NOR2_X1 U16125 ( .A1(n12917), .A2(n12916), .ZN(n12920) );
  AOI21_X1 U16126 ( .B1(n15195), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12918) );
  AOI21_X1 U16127 ( .B1(n12668), .B2(P1_EAX_REG_19__SCAN_IN), .A(n12918), .ZN(
        n12919) );
  OAI21_X1 U16128 ( .B1(n13078), .B2(n12920), .A(n12919), .ZN(n12921) );
  NAND2_X1 U16129 ( .A1(n12924), .A2(n15187), .ZN(n12925) );
  AND2_X1 U16130 ( .A1(n12965), .A2(n12925), .ZN(n15191) );
  AOI22_X1 U16131 ( .A1(n9623), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(n9621), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12929) );
  AOI22_X1 U16132 ( .A1(n13511), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13088), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12928) );
  AOI22_X1 U16133 ( .A1(n9606), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13068), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12927) );
  AOI22_X1 U16134 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13503), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12926) );
  NAND4_X1 U16135 ( .A1(n12929), .A2(n12928), .A3(n12927), .A4(n12926), .ZN(
        n12938) );
  AOI22_X1 U16136 ( .A1(n13512), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12720), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12936) );
  AOI22_X1 U16137 ( .A1(n13043), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12953), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12935) );
  INV_X1 U16138 ( .A(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12930) );
  OAI22_X1 U16139 ( .A1(n13106), .A2(n12931), .B1(n13108), .B2(n12930), .ZN(
        n12932) );
  INV_X1 U16140 ( .A(n12932), .ZN(n12934) );
  NAND4_X1 U16141 ( .A1(n12936), .A2(n12935), .A3(n12934), .A4(n12933), .ZN(
        n12937) );
  OR2_X1 U16142 ( .A1(n12938), .A2(n12937), .ZN(n12941) );
  INV_X1 U16143 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n14102) );
  OAI21_X1 U16144 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n21022), .A(
        n21070), .ZN(n12939) );
  OAI21_X1 U16145 ( .B1(n13526), .B2(n14102), .A(n12939), .ZN(n12940) );
  AOI21_X1 U16146 ( .B1(n13528), .B2(n12941), .A(n12940), .ZN(n12942) );
  AOI21_X1 U16147 ( .B1(n15191), .B2(n13531), .A(n12942), .ZN(n14772) );
  INV_X1 U16148 ( .A(n12943), .ZN(n12944) );
  INV_X1 U16149 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n21302) );
  NAND2_X1 U16150 ( .A1(n12944), .A2(n21302), .ZN(n12945) );
  NAND2_X1 U16151 ( .A1(n13009), .A2(n12945), .ZN(n15169) );
  AOI22_X1 U16152 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12461), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12949) );
  AOI22_X1 U16153 ( .A1(n12720), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13088), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12948) );
  AOI22_X1 U16154 ( .A1(n9597), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13016), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12947) );
  AOI22_X1 U16155 ( .A1(n13043), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13503), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12946) );
  NAND4_X1 U16156 ( .A1(n12949), .A2(n12948), .A3(n12947), .A4(n12946), .ZN(
        n12959) );
  AOI22_X1 U16157 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13511), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12957) );
  INV_X1 U16158 ( .A(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12950) );
  OAI22_X1 U16159 ( .A1(n13106), .A2(n12951), .B1(n9605), .B2(n12950), .ZN(
        n12952) );
  INV_X1 U16160 ( .A(n12952), .ZN(n12956) );
  AOI22_X1 U16161 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12953), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12955) );
  NAND4_X1 U16162 ( .A1(n12957), .A2(n12956), .A3(n12955), .A4(n12954), .ZN(
        n12958) );
  NOR2_X1 U16163 ( .A1(n12959), .A2(n12958), .ZN(n12962) );
  OAI21_X1 U16164 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n21022), .A(
        n21070), .ZN(n12961) );
  NAND2_X1 U16165 ( .A1(n12668), .A2(P1_EAX_REG_22__SCAN_IN), .ZN(n12960) );
  OAI211_X1 U16166 ( .C1(n13078), .C2(n12962), .A(n12961), .B(n12960), .ZN(
        n12963) );
  NAND2_X1 U16167 ( .A1(n12964), .A2(n12963), .ZN(n14750) );
  XNOR2_X1 U16168 ( .A(n12965), .B(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15177) );
  NAND2_X1 U16169 ( .A1(n15177), .A2(n13531), .ZN(n12981) );
  AOI22_X1 U16170 ( .A1(n13502), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13088), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12969) );
  AOI22_X1 U16171 ( .A1(n13510), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9621), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12968) );
  AOI22_X1 U16172 ( .A1(n12461), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13068), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12966) );
  NAND4_X1 U16173 ( .A1(n12969), .A2(n12968), .A3(n12967), .A4(n12966), .ZN(
        n12975) );
  AOI22_X1 U16174 ( .A1(n13512), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13511), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12973) );
  AOI22_X1 U16175 ( .A1(n9623), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13043), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12972) );
  AOI22_X1 U16176 ( .A1(n9597), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13016), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12971) );
  AOI22_X1 U16177 ( .A1(n9591), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13503), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12970) );
  NAND4_X1 U16178 ( .A1(n12973), .A2(n12972), .A3(n12971), .A4(n12970), .ZN(
        n12974) );
  NOR2_X1 U16179 ( .A1(n12975), .A2(n12974), .ZN(n12979) );
  NAND2_X1 U16180 ( .A1(n21070), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12976) );
  NAND2_X1 U16181 ( .A1(n13524), .A2(n12976), .ZN(n12977) );
  AOI21_X1 U16182 ( .B1(n13032), .B2(P1_EAX_REG_21__SCAN_IN), .A(n12977), .ZN(
        n12978) );
  OAI21_X1 U16183 ( .B1(n13078), .B2(n12979), .A(n12978), .ZN(n12980) );
  NAND2_X1 U16184 ( .A1(n12981), .A2(n12980), .ZN(n14760) );
  XNOR2_X1 U16185 ( .A(n13009), .B(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15163) );
  NAND2_X1 U16186 ( .A1(n15163), .A2(n13531), .ZN(n13008) );
  AOI22_X1 U16187 ( .A1(n13502), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13511), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12985) );
  AOI22_X1 U16188 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13088), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12984) );
  AOI22_X1 U16189 ( .A1(n13510), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13016), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12983) );
  AOI22_X1 U16190 ( .A1(n13512), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13504), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12982) );
  NAND4_X1 U16191 ( .A1(n12985), .A2(n12984), .A3(n12983), .A4(n12982), .ZN(
        n12991) );
  AOI22_X1 U16192 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n13043), .B1(
        n12953), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12988) );
  AOI22_X1 U16193 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n13513), .B1(
        n13503), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12987) );
  AOI22_X1 U16194 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13068), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12986) );
  NAND4_X1 U16195 ( .A1(n12989), .A2(n12988), .A3(n12987), .A4(n12986), .ZN(
        n12990) );
  NOR2_X1 U16196 ( .A1(n12991), .A2(n12990), .ZN(n13014) );
  AOI22_X1 U16197 ( .A1(n13502), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13511), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12995) );
  AOI22_X1 U16198 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12953), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12994) );
  AOI22_X1 U16199 ( .A1(n13088), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n13504), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12993) );
  AOI22_X1 U16200 ( .A1(n10147), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13016), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12992) );
  NAND4_X1 U16201 ( .A1(n12995), .A2(n12994), .A3(n12993), .A4(n12992), .ZN(
        n13001) );
  AOI22_X1 U16202 ( .A1(n13510), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9624), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12999) );
  AOI22_X1 U16203 ( .A1(n13512), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9617), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12998) );
  AOI22_X1 U16204 ( .A1(n12461), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13068), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12997) );
  AOI22_X1 U16205 ( .A1(n13043), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13503), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12996) );
  NAND4_X1 U16206 ( .A1(n12999), .A2(n12998), .A3(n12997), .A4(n12996), .ZN(
        n13000) );
  NOR2_X1 U16207 ( .A1(n13001), .A2(n13000), .ZN(n13015) );
  XOR2_X1 U16208 ( .A(n13014), .B(n13015), .Z(n13002) );
  NAND2_X1 U16209 ( .A1(n13002), .A2(n13528), .ZN(n13006) );
  NAND2_X1 U16210 ( .A1(n21070), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13003) );
  NAND2_X1 U16211 ( .A1(n13524), .A2(n13003), .ZN(n13004) );
  AOI21_X1 U16212 ( .B1(n13032), .B2(P1_EAX_REG_23__SCAN_IN), .A(n13004), .ZN(
        n13005) );
  NAND2_X1 U16213 ( .A1(n13006), .A2(n13005), .ZN(n13007) );
  AND2_X2 U16214 ( .A1(n13010), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13011) );
  INV_X1 U16215 ( .A(n13011), .ZN(n13012) );
  INV_X1 U16216 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14727) );
  NAND2_X1 U16217 ( .A1(n13012), .A2(n14727), .ZN(n13013) );
  NAND2_X1 U16218 ( .A1(n13054), .A2(n13013), .ZN(n15153) );
  NOR2_X1 U16219 ( .A1(n13015), .A2(n13014), .ZN(n13038) );
  AOI22_X1 U16220 ( .A1(n13502), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13511), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13023) );
  AOI22_X1 U16221 ( .A1(n9584), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13088), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13022) );
  AOI22_X1 U16222 ( .A1(n13510), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13016), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13021) );
  INV_X1 U16223 ( .A(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13017) );
  OAI22_X1 U16224 ( .A1(n9604), .A2(n13018), .B1(n13108), .B2(n13017), .ZN(
        n13019) );
  INV_X1 U16225 ( .A(n13019), .ZN(n13020) );
  NAND4_X1 U16226 ( .A1(n13023), .A2(n13022), .A3(n13021), .A4(n13020), .ZN(
        n13029) );
  INV_X1 U16227 ( .A(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n21253) );
  AOI22_X1 U16228 ( .A1(n13043), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12953), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13026) );
  AOI22_X1 U16229 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13503), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13025) );
  AOI22_X1 U16230 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13068), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13024) );
  NAND4_X1 U16231 ( .A1(n13027), .A2(n13026), .A3(n13025), .A4(n13024), .ZN(
        n13028) );
  OR2_X1 U16232 ( .A1(n13029), .A2(n13028), .ZN(n13037) );
  XNOR2_X1 U16233 ( .A(n13038), .B(n13037), .ZN(n13034) );
  NAND2_X1 U16234 ( .A1(n21070), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13030) );
  NAND2_X1 U16235 ( .A1(n13524), .A2(n13030), .ZN(n13031) );
  AOI21_X1 U16236 ( .B1(n13032), .B2(P1_EAX_REG_24__SCAN_IN), .A(n13031), .ZN(
        n13033) );
  OAI21_X1 U16237 ( .B1(n13034), .B2(n13078), .A(n13033), .ZN(n13035) );
  XNOR2_X1 U16238 ( .A(n13054), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15147) );
  NAND2_X1 U16239 ( .A1(n13038), .A2(n13037), .ZN(n13059) );
  AOI22_X1 U16240 ( .A1(n13512), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13088), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13042) );
  AOI22_X1 U16241 ( .A1(n13510), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9597), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13041) );
  AOI22_X1 U16242 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12382), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13039) );
  NAND4_X1 U16243 ( .A1(n13042), .A2(n13041), .A3(n13040), .A4(n13039), .ZN(
        n13049) );
  AOI22_X1 U16244 ( .A1(n13502), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13511), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13047) );
  AOI22_X1 U16245 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13043), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13046) );
  AOI22_X1 U16246 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12953), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13045) );
  AOI22_X1 U16247 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13068), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13044) );
  NAND4_X1 U16248 ( .A1(n13047), .A2(n13046), .A3(n13045), .A4(n13044), .ZN(
        n13048) );
  NOR2_X1 U16249 ( .A1(n13049), .A2(n13048), .ZN(n13060) );
  XOR2_X1 U16250 ( .A(n13059), .B(n13060), .Z(n13052) );
  INV_X1 U16251 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n15038) );
  OAI21_X1 U16252 ( .B1(n21022), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n21070), .ZN(n13050) );
  OAI21_X1 U16253 ( .B1(n13526), .B2(n15038), .A(n13050), .ZN(n13051) );
  AOI21_X1 U16254 ( .B1(n13052), .B2(n13528), .A(n13051), .ZN(n13053) );
  AOI21_X1 U16255 ( .B1(n15147), .B2(n13531), .A(n13053), .ZN(n14707) );
  AND2_X2 U16256 ( .A1(n14705), .A2(n14707), .ZN(n14689) );
  INV_X1 U16257 ( .A(n13054), .ZN(n13055) );
  INV_X1 U16258 ( .A(n13056), .ZN(n13057) );
  INV_X1 U16259 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n13075) );
  NAND2_X1 U16260 ( .A1(n13057), .A2(n13075), .ZN(n13058) );
  NAND2_X1 U16261 ( .A1(n13099), .A2(n13058), .ZN(n15134) );
  NOR2_X1 U16262 ( .A1(n13060), .A2(n13059), .ZN(n13083) );
  AOI22_X1 U16263 ( .A1(n13502), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13511), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13067) );
  AOI22_X1 U16264 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13088), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13066) );
  AOI22_X1 U16265 ( .A1(n13510), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12382), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13065) );
  INV_X1 U16266 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13062) );
  INV_X1 U16267 ( .A(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13061) );
  OAI22_X1 U16268 ( .A1(n9604), .A2(n13062), .B1(n13108), .B2(n13061), .ZN(
        n13063) );
  INV_X1 U16269 ( .A(n13063), .ZN(n13064) );
  NAND4_X1 U16270 ( .A1(n13067), .A2(n13066), .A3(n13065), .A4(n13064), .ZN(
        n13074) );
  AOI22_X1 U16271 ( .A1(n13043), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12953), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13071) );
  AOI22_X1 U16272 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13503), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13070) );
  AOI22_X1 U16273 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13068), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13069) );
  NAND4_X1 U16274 ( .A1(n13072), .A2(n13071), .A3(n13070), .A4(n13069), .ZN(
        n13073) );
  OR2_X1 U16275 ( .A1(n13074), .A2(n13073), .ZN(n13082) );
  XNOR2_X1 U16276 ( .A(n13083), .B(n13082), .ZN(n13079) );
  AOI21_X1 U16277 ( .B1(n13075), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13076) );
  AOI21_X1 U16278 ( .B1(n12668), .B2(P1_EAX_REG_26__SCAN_IN), .A(n13076), .ZN(
        n13077) );
  OAI21_X1 U16279 ( .B1(n13079), .B2(n13078), .A(n13077), .ZN(n13080) );
  INV_X1 U16280 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14679) );
  XNOR2_X1 U16281 ( .A(n13099), .B(n14679), .ZN(n15125) );
  INV_X1 U16282 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n15028) );
  NAND2_X1 U16283 ( .A1(n13083), .A2(n13082), .ZN(n13121) );
  AOI22_X1 U16284 ( .A1(n13502), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9621), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13087) );
  AOI22_X1 U16285 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10147), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13086) );
  AOI22_X1 U16286 ( .A1(n13043), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12953), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13085) );
  AOI22_X1 U16287 ( .A1(n9597), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12382), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13084) );
  NAND4_X1 U16288 ( .A1(n13087), .A2(n13086), .A3(n13085), .A4(n13084), .ZN(
        n13094) );
  AOI22_X1 U16289 ( .A1(n13510), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13512), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13092) );
  AOI22_X1 U16290 ( .A1(n13511), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13088), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13091) );
  AOI22_X1 U16291 ( .A1(n9606), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13068), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13090) );
  AOI22_X1 U16292 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13503), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13089) );
  NAND4_X1 U16293 ( .A1(n13092), .A2(n13091), .A3(n13090), .A4(n13089), .ZN(
        n13093) );
  NOR2_X1 U16294 ( .A1(n13094), .A2(n13093), .ZN(n13122) );
  XOR2_X1 U16295 ( .A(n13121), .B(n13122), .Z(n13095) );
  NAND2_X1 U16296 ( .A1(n13095), .A2(n13528), .ZN(n13097) );
  AOI21_X1 U16297 ( .B1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n21070), .A(
        n13531), .ZN(n13096) );
  OAI211_X1 U16298 ( .C1(n13526), .C2(n15028), .A(n13097), .B(n13096), .ZN(
        n13098) );
  INV_X1 U16299 ( .A(n13099), .ZN(n13100) );
  INV_X1 U16300 ( .A(n13101), .ZN(n13102) );
  INV_X1 U16301 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14524) );
  NAND2_X1 U16302 ( .A1(n13102), .A2(n14524), .ZN(n13103) );
  NOR2_X1 U16303 ( .A1(n14524), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13104) );
  AOI211_X1 U16304 ( .C1(n12668), .C2(P1_EAX_REG_28__SCAN_IN), .A(n13531), .B(
        n13104), .ZN(n13125) );
  INV_X1 U16305 ( .A(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13105) );
  NOR2_X1 U16306 ( .A1(n13106), .A2(n13105), .ZN(n13112) );
  INV_X1 U16307 ( .A(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13107) );
  OAI22_X1 U16308 ( .A1(n9604), .A2(n13109), .B1(n13108), .B2(n13107), .ZN(
        n13111) );
  AOI211_X1 U16309 ( .C1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .C2(n13016), .A(
        n13112), .B(n13111), .ZN(n13120) );
  AOI22_X1 U16310 ( .A1(n13502), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13511), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13119) );
  AOI22_X1 U16311 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13088), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13118) );
  AOI22_X1 U16312 ( .A1(n12461), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12353), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13116) );
  AOI22_X1 U16313 ( .A1(n13043), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12953), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13115) );
  AOI22_X1 U16314 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13503), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13114) );
  AOI22_X1 U16315 ( .A1(n9623), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13068), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13113) );
  AND4_X1 U16316 ( .A1(n13116), .A2(n13115), .A3(n13114), .A4(n13113), .ZN(
        n13117) );
  NAND4_X1 U16317 ( .A1(n13120), .A2(n13119), .A3(n13118), .A4(n13117), .ZN(
        n13278) );
  NOR2_X1 U16318 ( .A1(n13122), .A2(n13121), .ZN(n13279) );
  XOR2_X1 U16319 ( .A(n13278), .B(n13279), .Z(n13123) );
  NAND2_X1 U16320 ( .A1(n13123), .A2(n13528), .ZN(n13124) );
  NAND3_X1 U16321 ( .A1(n10368), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n17183) );
  INV_X1 U16322 ( .A(n17183), .ZN(n13129) );
  NOR2_X2 U16323 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21383) );
  NAND2_X1 U16324 ( .A1(n13158), .A2(n13152), .ZN(n13151) );
  NAND2_X1 U16325 ( .A1(n13151), .A2(n13146), .ZN(n13142) );
  AND2_X1 U16326 ( .A1(n13140), .A2(n13136), .ZN(n13131) );
  NAND2_X1 U16327 ( .A1(n13142), .A2(n13131), .ZN(n13172) );
  XNOR2_X1 U16328 ( .A(n13172), .B(n13173), .ZN(n13132) );
  NAND2_X1 U16329 ( .A1(n13132), .A2(n13187), .ZN(n13133) );
  INV_X1 U16330 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n14495) );
  NAND2_X1 U16331 ( .A1(n13142), .A2(n13140), .ZN(n13137) );
  XNOR2_X1 U16332 ( .A(n13137), .B(n13136), .ZN(n13138) );
  NAND2_X1 U16333 ( .A1(n13138), .A2(n13187), .ZN(n13139) );
  INV_X1 U16334 ( .A(n13140), .ZN(n13141) );
  XNOR2_X1 U16335 ( .A(n13142), .B(n13141), .ZN(n13143) );
  NAND2_X1 U16336 ( .A1(n13143), .A2(n13187), .ZN(n13144) );
  AOI21_X1 U16337 ( .B1(n14430), .B2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13167) );
  NAND2_X1 U16338 ( .A1(n13145), .A2(n13858), .ZN(n13150) );
  XNOR2_X1 U16339 ( .A(n13151), .B(n13146), .ZN(n13148) );
  NAND2_X1 U16340 ( .A1(n12427), .A2(n12414), .ZN(n13157) );
  INV_X1 U16341 ( .A(n13157), .ZN(n13147) );
  AOI21_X1 U16342 ( .B1(n13148), .B2(n13187), .A(n13147), .ZN(n13149) );
  NAND2_X1 U16343 ( .A1(n13150), .A2(n13149), .ZN(n14313) );
  OAI21_X1 U16344 ( .B1(n13152), .B2(n13158), .A(n13151), .ZN(n13153) );
  INV_X1 U16345 ( .A(n13153), .ZN(n13155) );
  AOI21_X1 U16346 ( .B1(n13187), .B2(n13155), .A(n13154), .ZN(n13156) );
  OR2_X1 U16347 ( .A1(n20661), .A2(n13258), .ZN(n13161) );
  OAI21_X1 U16348 ( .B1(n21216), .B2(n13158), .A(n13157), .ZN(n13159) );
  INV_X1 U16349 ( .A(n13159), .ZN(n13160) );
  NAND2_X1 U16350 ( .A1(n13161), .A2(n13160), .ZN(n13922) );
  NAND2_X1 U16351 ( .A1(n13922), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13921) );
  XNOR2_X1 U16352 ( .A(n13163), .B(n13921), .ZN(n15314) );
  NAND2_X1 U16353 ( .A1(n15314), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15315) );
  INV_X1 U16354 ( .A(n13921), .ZN(n13162) );
  NAND2_X1 U16355 ( .A1(n13163), .A2(n13162), .ZN(n13164) );
  INV_X1 U16356 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20548) );
  NAND2_X1 U16357 ( .A1(n13165), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13166) );
  NAND2_X1 U16358 ( .A1(n13168), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13169) );
  NAND3_X1 U16359 ( .A1(n13170), .A2(n13858), .A3(n13171), .ZN(n13177) );
  INV_X1 U16360 ( .A(n13172), .ZN(n13174) );
  NAND2_X1 U16361 ( .A1(n13174), .A2(n13173), .ZN(n13183) );
  XNOR2_X1 U16362 ( .A(n13183), .B(n13184), .ZN(n13175) );
  NAND2_X1 U16363 ( .A1(n13175), .A2(n13187), .ZN(n13176) );
  NAND2_X1 U16364 ( .A1(n13177), .A2(n13176), .ZN(n14454) );
  INV_X1 U16365 ( .A(n14454), .ZN(n13179) );
  INV_X1 U16366 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13178) );
  NAND2_X1 U16367 ( .A1(n14454), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13181) );
  INV_X1 U16368 ( .A(n13183), .ZN(n13185) );
  NAND2_X1 U16369 ( .A1(n13185), .A2(n13184), .ZN(n13196) );
  XNOR2_X1 U16370 ( .A(n13196), .B(n13186), .ZN(n13188) );
  NAND2_X1 U16371 ( .A1(n13188), .A2(n13187), .ZN(n13189) );
  NAND2_X1 U16372 ( .A1(n13190), .A2(n13189), .ZN(n13191) );
  INV_X1 U16373 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n14506) );
  XNOR2_X1 U16374 ( .A(n13191), .B(n14506), .ZN(n14483) );
  NAND2_X1 U16375 ( .A1(n13191), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13192) );
  NOR2_X1 U16376 ( .A1(n13193), .A2(n13258), .ZN(n13194) );
  OR3_X1 U16377 ( .A1(n13196), .A2(n13195), .A3(n21216), .ZN(n13197) );
  NAND2_X1 U16378 ( .A1(n13202), .A2(n13197), .ZN(n13199) );
  XNOR2_X1 U16379 ( .A(n13199), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15306) );
  INV_X1 U16380 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15530) );
  NOR2_X1 U16381 ( .A1(n9569), .A2(n15530), .ZN(n15212) );
  AND2_X1 U16382 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15454) );
  AND2_X1 U16383 ( .A1(n15454), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15435) );
  OR2_X1 U16384 ( .A1(n13199), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15210) );
  NAND2_X1 U16385 ( .A1(n9569), .A2(n15530), .ZN(n15214) );
  OAI211_X1 U16386 ( .C1(n9952), .C2(n15435), .A(n15210), .B(n15214), .ZN(
        n13204) );
  INV_X1 U16387 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15502) );
  NAND2_X1 U16388 ( .A1(n13202), .A2(n15502), .ZN(n15264) );
  NAND2_X1 U16389 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n13200) );
  NAND2_X1 U16390 ( .A1(n13202), .A2(n13200), .ZN(n15261) );
  AND2_X1 U16391 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14556) );
  INV_X1 U16392 ( .A(n14556), .ZN(n13201) );
  NAND2_X1 U16393 ( .A1(n9569), .A2(n13201), .ZN(n13203) );
  NAND3_X1 U16394 ( .A1(n15264), .A2(n15261), .A3(n13203), .ZN(n15231) );
  NOR2_X1 U16395 ( .A1(n13204), .A2(n15231), .ZN(n13205) );
  NOR2_X1 U16396 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15259) );
  NAND2_X1 U16397 ( .A1(n15259), .A2(n15502), .ZN(n15215) );
  NOR2_X1 U16398 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15217) );
  NOR2_X1 U16399 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15455) );
  INV_X1 U16400 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n13369) );
  NAND3_X1 U16401 ( .A1(n15217), .A2(n15455), .A3(n13369), .ZN(n13206) );
  NOR2_X1 U16402 ( .A1(n15215), .A2(n13206), .ZN(n13207) );
  NAND2_X1 U16403 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14571) );
  INV_X1 U16404 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15175) );
  NOR2_X1 U16405 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n13211) );
  AND2_X1 U16406 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14574) );
  NAND2_X1 U16407 ( .A1(n14574), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14563) );
  NAND2_X1 U16408 ( .A1(n9569), .A2(n14563), .ZN(n15129) );
  NAND2_X1 U16409 ( .A1(n15158), .A2(n15129), .ZN(n13214) );
  NOR2_X1 U16410 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15138) );
  INV_X1 U16411 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15142) );
  NAND2_X1 U16412 ( .A1(n15138), .A2(n15142), .ZN(n14533) );
  OAI21_X1 U16413 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n14533), .A(
        n13214), .ZN(n13213) );
  INV_X1 U16414 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13404) );
  MUX2_X1 U16415 ( .A(n13404), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n9569), .Z(n13212) );
  NAND2_X1 U16416 ( .A1(n21069), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13217) );
  NAND2_X1 U16417 ( .A1(n13215), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n13216) );
  NAND2_X1 U16418 ( .A1(n13217), .A2(n13216), .ZN(n13224) );
  NAND2_X1 U16419 ( .A1(n12649), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n13218) );
  NAND2_X1 U16420 ( .A1(n13221), .A2(n13218), .ZN(n13238) );
  INV_X1 U16421 ( .A(n13238), .ZN(n13219) );
  MUX2_X1 U16422 ( .A(n20589), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n13254) );
  AOI222_X1 U16423 ( .A1(n13252), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .B1(n13252), .B2(n12693), .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .C2(n12693), .ZN(n13303) );
  NAND2_X1 U16424 ( .A1(n13303), .A2(n13248), .ZN(n13267) );
  NAND2_X1 U16425 ( .A1(n12403), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13222) );
  NAND2_X1 U16426 ( .A1(n13223), .A2(n17135), .ZN(n13259) );
  NAND2_X1 U16427 ( .A1(n13224), .A2(n13227), .ZN(n13225) );
  NAND2_X1 U16428 ( .A1(n13226), .A2(n13225), .ZN(n13301) );
  NAND2_X1 U16429 ( .A1(n13234), .A2(n13237), .ZN(n13236) );
  OAI21_X1 U16430 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20988), .A(
        n13227), .ZN(n13228) );
  INV_X1 U16431 ( .A(n13228), .ZN(n13231) );
  NAND2_X1 U16432 ( .A1(n13248), .A2(n13231), .ZN(n13229) );
  NAND2_X1 U16433 ( .A1(n13260), .A2(n13858), .ZN(n13268) );
  NAND2_X1 U16434 ( .A1(n13229), .A2(n13268), .ZN(n13233) );
  NAND2_X1 U16435 ( .A1(n12403), .A2(n14486), .ZN(n13230) );
  NAND2_X1 U16436 ( .A1(n13230), .A2(n20603), .ZN(n13246) );
  OAI211_X1 U16437 ( .C1(n12420), .C2(n12427), .A(n13246), .B(n13231), .ZN(
        n13232) );
  OAI211_X1 U16438 ( .C1(n13234), .C2(n13237), .A(n13233), .B(n13232), .ZN(
        n13235) );
  OAI211_X1 U16439 ( .C1(n13259), .C2(n13237), .A(n13236), .B(n13235), .ZN(
        n13245) );
  NAND2_X1 U16440 ( .A1(n13239), .A2(n13238), .ZN(n13241) );
  NAND2_X1 U16441 ( .A1(n13241), .A2(n13240), .ZN(n13300) );
  NAND2_X1 U16442 ( .A1(n13248), .A2(n13247), .ZN(n13242) );
  OAI211_X1 U16443 ( .C1(n13247), .C2(n13243), .A(n13242), .B(n13246), .ZN(
        n13244) );
  NAND2_X1 U16444 ( .A1(n13245), .A2(n13244), .ZN(n13251) );
  INV_X1 U16445 ( .A(n13246), .ZN(n13249) );
  NAND3_X1 U16446 ( .A1(n13249), .A2(n13248), .A3(n13247), .ZN(n13250) );
  AND2_X1 U16447 ( .A1(n12693), .A2(n13252), .ZN(n13253) );
  NAND2_X1 U16448 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n13253), .ZN(
        n13302) );
  NOR2_X1 U16449 ( .A1(n13255), .A2(n13254), .ZN(n13256) );
  OAI22_X1 U16450 ( .A1(n13259), .A2(n13302), .B1(n13262), .B2(n13258), .ZN(
        n13261) );
  OAI21_X1 U16451 ( .B1(n13263), .B2(n13261), .A(n13260), .ZN(n13266) );
  NAND2_X1 U16452 ( .A1(n10368), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13265) );
  NAND3_X1 U16453 ( .A1(n13263), .A2(n13262), .A3(n13302), .ZN(n13264) );
  INV_X1 U16454 ( .A(n13268), .ZN(n13269) );
  NAND2_X1 U16455 ( .A1(n13303), .A2(n13269), .ZN(n13270) );
  AOI21_X1 U16456 ( .B1(n15582), .B2(n12427), .A(n12415), .ZN(n13272) );
  NAND2_X1 U16457 ( .A1(n13876), .A2(n13860), .ZN(n14645) );
  OR2_X1 U16458 ( .A1(n13275), .A2(n21383), .ZN(n21220) );
  NAND2_X1 U16459 ( .A1(n21220), .A2(n10368), .ZN(n13273) );
  NAND2_X1 U16460 ( .A1(n10368), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21133) );
  NAND2_X1 U16461 ( .A1(n21022), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13274) );
  NAND2_X1 U16462 ( .A1(n21133), .A2(n13274), .ZN(n13920) );
  NAND2_X1 U16463 ( .A1(n20577), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n15334) );
  OAI21_X1 U16464 ( .B1(n17161), .B2(n14524), .A(n15334), .ZN(n13276) );
  AOI21_X1 U16465 ( .B1(n14523), .B2(n15200), .A(n13276), .ZN(n13277) );
  INV_X1 U16466 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n13427) );
  XNOR2_X1 U16467 ( .A(n13296), .B(n13427), .ZN(n15116) );
  INV_X1 U16468 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n15021) );
  NAND2_X1 U16469 ( .A1(n13279), .A2(n13278), .ZN(n13520) );
  AOI22_X1 U16470 ( .A1(n13512), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13511), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13283) );
  AOI22_X1 U16471 ( .A1(n13510), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13504), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13282) );
  AOI22_X1 U16472 ( .A1(n12953), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13503), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13281) );
  AOI22_X1 U16473 ( .A1(n9606), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12382), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13280) );
  NAND4_X1 U16474 ( .A1(n13283), .A2(n13282), .A3(n13281), .A4(n13280), .ZN(
        n13289) );
  AOI22_X1 U16475 ( .A1(n13502), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13088), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13287) );
  AOI22_X1 U16476 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(n9621), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13286) );
  AOI22_X1 U16477 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13043), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13285) );
  AOI22_X1 U16478 ( .A1(n12353), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13068), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13284) );
  NAND4_X1 U16479 ( .A1(n13287), .A2(n13286), .A3(n13285), .A4(n13284), .ZN(
        n13288) );
  NOR2_X1 U16480 ( .A1(n13289), .A2(n13288), .ZN(n13521) );
  XOR2_X1 U16481 ( .A(n13520), .B(n13521), .Z(n13290) );
  NAND2_X1 U16482 ( .A1(n13290), .A2(n13528), .ZN(n13292) );
  AOI21_X1 U16483 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n21070), .A(
        n13531), .ZN(n13291) );
  OAI211_X1 U16484 ( .C1(n13526), .C2(n15021), .A(n13292), .B(n13291), .ZN(
        n13293) );
  OAI21_X1 U16485 ( .B1(n15116), .B2(n13524), .A(n13293), .ZN(n13295) );
  INV_X1 U16486 ( .A(n15118), .ZN(n15025) );
  INV_X1 U16487 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n15109) );
  NOR3_X1 U16488 ( .A1(n13301), .A2(n13300), .A3(n13299), .ZN(n13304) );
  OAI21_X1 U16489 ( .B1(n13304), .B2(n13303), .A(n13302), .ZN(n14650) );
  AND2_X1 U16490 ( .A1(n14650), .A2(n13305), .ZN(n14654) );
  NAND2_X1 U16491 ( .A1(n14654), .A2(n14077), .ZN(n13637) );
  NOR2_X1 U16492 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21218) );
  NAND2_X1 U16493 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21218), .ZN(n17143) );
  AND2_X1 U16494 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n10368), .ZN(n13306) );
  NAND2_X1 U16495 ( .A1(n13531), .A2(n13306), .ZN(n13307) );
  OAI21_X1 U16496 ( .B1(n17143), .B2(n10368), .A(n13307), .ZN(n13308) );
  NAND2_X1 U16497 ( .A1(n20410), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13425) );
  OR2_X4 U16498 ( .A1(n14583), .A2(n13425), .ZN(n20393) );
  INV_X2 U16499 ( .A(n14658), .ZN(n14641) );
  OR2_X1 U16500 ( .A1(n13350), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13311) );
  INV_X1 U16501 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13313) );
  OR2_X1 U16502 ( .A1(n13323), .A2(n13313), .ZN(n13315) );
  NAND2_X1 U16503 ( .A1(n14658), .A2(n13313), .ZN(n13314) );
  NAND2_X1 U16504 ( .A1(n13315), .A2(n13314), .ZN(n13909) );
  INV_X1 U16505 ( .A(n13317), .ZN(n13318) );
  INV_X1 U16506 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n14952) );
  NAND2_X1 U16507 ( .A1(n13318), .A2(n14952), .ZN(n13322) );
  NAND2_X1 U16508 ( .A1(n14544), .A2(n14952), .ZN(n13320) );
  INV_X1 U16509 ( .A(n13323), .ZN(n13319) );
  OAI211_X1 U16510 ( .C1(n14658), .C2(n20548), .A(n13320), .B(n13396), .ZN(
        n13321) );
  INV_X1 U16511 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13325) );
  NAND2_X1 U16512 ( .A1(n13395), .A2(n13325), .ZN(n13329) );
  INV_X1 U16513 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14493) );
  NAND2_X1 U16514 ( .A1(n13396), .A2(n14493), .ZN(n13327) );
  NAND2_X1 U16515 ( .A1(n14544), .A2(n13325), .ZN(n13326) );
  NAND3_X1 U16516 ( .A1(n13327), .A2(n14641), .A3(n13326), .ZN(n13328) );
  AND2_X1 U16517 ( .A1(n13329), .A2(n13328), .ZN(n14297) );
  INV_X1 U16518 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n14494) );
  INV_X1 U16519 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n20446) );
  NAND2_X1 U16520 ( .A1(n14544), .A2(n20446), .ZN(n13331) );
  OAI211_X1 U16521 ( .C1(n14658), .C2(n14494), .A(n13331), .B(n13396), .ZN(
        n13332) );
  OAI21_X1 U16522 ( .B1(n13317), .B2(P1_EBX_REG_4__SCAN_IN), .A(n13332), .ZN(
        n20416) );
  INV_X1 U16523 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n20391) );
  NAND2_X1 U16524 ( .A1(n14544), .A2(n20391), .ZN(n13333) );
  OAI211_X1 U16525 ( .C1(n14658), .C2(n13178), .A(n13333), .B(n13396), .ZN(
        n13334) );
  OAI21_X1 U16526 ( .B1(n13317), .B2(P1_EBX_REG_6__SCAN_IN), .A(n13334), .ZN(
        n14450) );
  OAI21_X1 U16527 ( .B1(n14658), .B2(n14495), .A(n13396), .ZN(n13336) );
  INV_X1 U16528 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n14443) );
  NAND2_X1 U16529 ( .A1(n14544), .A2(n14443), .ZN(n13335) );
  NAND2_X1 U16530 ( .A1(n13336), .A2(n13335), .ZN(n13338) );
  NAND2_X1 U16531 ( .A1(n13395), .A2(n14443), .ZN(n13337) );
  AND2_X1 U16532 ( .A1(n13338), .A2(n13337), .ZN(n14442) );
  NOR2_X1 U16533 ( .A1(n14450), .A2(n14442), .ZN(n13339) );
  OAI21_X1 U16534 ( .B1(n14658), .B2(n14506), .A(n13396), .ZN(n13341) );
  INV_X1 U16535 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n15012) );
  NAND2_X1 U16536 ( .A1(n14544), .A2(n15012), .ZN(n13340) );
  NAND2_X1 U16537 ( .A1(n13341), .A2(n13340), .ZN(n13342) );
  OAI21_X1 U16538 ( .B1(P1_EBX_REG_7__SCAN_IN), .B2(n13408), .A(n13342), .ZN(
        n14504) );
  NAND2_X1 U16539 ( .A1(n14449), .A2(n14504), .ZN(n14503) );
  INV_X1 U16540 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n13344) );
  INV_X1 U16541 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n20443) );
  NAND2_X1 U16542 ( .A1(n14544), .A2(n20443), .ZN(n13343) );
  OAI211_X1 U16543 ( .C1(n14658), .C2(n13344), .A(n13343), .B(n13396), .ZN(
        n13345) );
  OAI21_X1 U16544 ( .B1(n13317), .B2(P1_EBX_REG_8__SCAN_IN), .A(n13345), .ZN(
        n15540) );
  INV_X1 U16545 ( .A(n14544), .ZN(n14550) );
  OAI21_X1 U16546 ( .B1(n14658), .B2(n15530), .A(n13396), .ZN(n13347) );
  OAI21_X1 U16547 ( .B1(P1_EBX_REG_9__SCAN_IN), .B2(n14550), .A(n13347), .ZN(
        n13349) );
  INV_X1 U16548 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n15006) );
  NAND2_X1 U16549 ( .A1(n13395), .A2(n15006), .ZN(n13348) );
  MUX2_X1 U16550 ( .A(n13317), .B(n14641), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n13352) );
  OR2_X1 U16551 ( .A1(n14551), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13351) );
  INV_X1 U16552 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15493) );
  NAND2_X1 U16553 ( .A1(n13396), .A2(n15493), .ZN(n13354) );
  INV_X1 U16554 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n14998) );
  NAND2_X1 U16555 ( .A1(n14544), .A2(n14998), .ZN(n13353) );
  NAND3_X1 U16556 ( .A1(n13354), .A2(n14641), .A3(n13353), .ZN(n13355) );
  OAI21_X1 U16557 ( .B1(n13408), .B2(P1_EBX_REG_11__SCAN_IN), .A(n13355), .ZN(
        n14910) );
  NAND2_X1 U16558 ( .A1(n14909), .A2(n14910), .ZN(n14896) );
  MUX2_X1 U16559 ( .A(n13317), .B(n14641), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n13356) );
  OAI21_X1 U16560 ( .B1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n14551), .A(
        n13356), .ZN(n14898) );
  INV_X1 U16561 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n13357) );
  NAND2_X1 U16562 ( .A1(n13395), .A2(n13357), .ZN(n13361) );
  INV_X1 U16563 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15482) );
  NAND2_X1 U16564 ( .A1(n13396), .A2(n15482), .ZN(n13359) );
  NAND2_X1 U16565 ( .A1(n14544), .A2(n13357), .ZN(n13358) );
  NAND3_X1 U16566 ( .A1(n13359), .A2(n14641), .A3(n13358), .ZN(n13360) );
  MUX2_X1 U16567 ( .A(n13317), .B(n14641), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n13363) );
  OR2_X1 U16568 ( .A1(n14551), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13362) );
  MUX2_X1 U16569 ( .A(n13317), .B(n14641), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n13364) );
  OAI21_X1 U16570 ( .B1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n14551), .A(
        n13364), .ZN(n14829) );
  INV_X1 U16571 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14993) );
  NAND2_X1 U16572 ( .A1(n13395), .A2(n14993), .ZN(n13368) );
  INV_X1 U16573 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15218) );
  NAND2_X1 U16574 ( .A1(n13396), .A2(n15218), .ZN(n13366) );
  NAND2_X1 U16575 ( .A1(n14544), .A2(n14993), .ZN(n13365) );
  NAND3_X1 U16576 ( .A1(n13366), .A2(n14641), .A3(n13365), .ZN(n13367) );
  INV_X1 U16577 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n13370) );
  NAND2_X1 U16578 ( .A1(n13395), .A2(n13370), .ZN(n13374) );
  NAND2_X1 U16579 ( .A1(n13396), .A2(n13369), .ZN(n13372) );
  NAND2_X1 U16580 ( .A1(n14544), .A2(n13370), .ZN(n13371) );
  NAND3_X1 U16581 ( .A1(n13372), .A2(n14641), .A3(n13371), .ZN(n13373) );
  MUX2_X1 U16582 ( .A(n13317), .B(n14641), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n13376) );
  OR2_X1 U16583 ( .A1(n14551), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13375) );
  INV_X1 U16584 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15409) );
  OAI21_X1 U16585 ( .B1(n14658), .B2(n15409), .A(n13323), .ZN(n13378) );
  INV_X1 U16586 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14989) );
  NAND2_X1 U16587 ( .A1(n14544), .A2(n14989), .ZN(n13377) );
  NAND2_X1 U16588 ( .A1(n13378), .A2(n13377), .ZN(n13379) );
  OAI21_X1 U16589 ( .B1(P1_EBX_REG_19__SCAN_IN), .B2(n13408), .A(n13379), .ZN(
        n14789) );
  NAND2_X1 U16590 ( .A1(n14788), .A2(n14789), .ZN(n14773) );
  INV_X1 U16591 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n13381) );
  INV_X1 U16592 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14782) );
  NAND2_X1 U16593 ( .A1(n14544), .A2(n14782), .ZN(n13380) );
  OAI211_X1 U16594 ( .C1(n14658), .C2(n13381), .A(n13380), .B(n13396), .ZN(
        n13382) );
  OAI21_X1 U16595 ( .B1(n13317), .B2(P1_EBX_REG_20__SCAN_IN), .A(n13382), .ZN(
        n14776) );
  OR2_X2 U16596 ( .A1(n14773), .A2(n14776), .ZN(n14774) );
  INV_X1 U16597 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n13383) );
  NAND2_X1 U16598 ( .A1(n13395), .A2(n13383), .ZN(n13387) );
  NAND2_X1 U16599 ( .A1(n13396), .A2(n15175), .ZN(n13385) );
  NAND2_X1 U16600 ( .A1(n14544), .A2(n13383), .ZN(n13384) );
  NAND3_X1 U16601 ( .A1(n13385), .A2(n14641), .A3(n13384), .ZN(n13386) );
  MUX2_X1 U16602 ( .A(n13317), .B(n14641), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n13389) );
  OR2_X1 U16603 ( .A1(n14551), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13388) );
  AND2_X2 U16604 ( .A1(n14761), .A2(n14748), .ZN(n14746) );
  INV_X1 U16605 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n13390) );
  OAI21_X1 U16606 ( .B1(n14658), .B2(n13390), .A(n13323), .ZN(n13392) );
  INV_X1 U16607 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14985) );
  NAND2_X1 U16608 ( .A1(n14544), .A2(n14985), .ZN(n13391) );
  NAND2_X1 U16609 ( .A1(n13392), .A2(n13391), .ZN(n13393) );
  OAI21_X1 U16610 ( .B1(P1_EBX_REG_23__SCAN_IN), .B2(n13408), .A(n13393), .ZN(
        n14734) );
  MUX2_X1 U16611 ( .A(n13317), .B(n14641), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n13394) );
  OAI21_X1 U16612 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n14551), .A(
        n13394), .ZN(n14723) );
  INV_X1 U16613 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n13397) );
  NAND2_X1 U16614 ( .A1(n13395), .A2(n13397), .ZN(n13401) );
  NAND2_X1 U16615 ( .A1(n13396), .A2(n15142), .ZN(n13399) );
  NAND2_X1 U16616 ( .A1(n14544), .A2(n13397), .ZN(n13398) );
  NAND3_X1 U16617 ( .A1(n13399), .A2(n14641), .A3(n13398), .ZN(n13400) );
  AND2_X1 U16618 ( .A1(n13401), .A2(n13400), .ZN(n14708) );
  INV_X1 U16619 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14565) );
  INV_X1 U16620 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14981) );
  NAND2_X1 U16621 ( .A1(n14544), .A2(n14981), .ZN(n13402) );
  OAI211_X1 U16622 ( .C1(n14658), .C2(n14565), .A(n13402), .B(n13396), .ZN(
        n13403) );
  OAI21_X1 U16623 ( .B1(n13317), .B2(P1_EBX_REG_26__SCAN_IN), .A(n13403), .ZN(
        n14691) );
  NAND2_X1 U16624 ( .A1(n13396), .A2(n13404), .ZN(n13406) );
  INV_X1 U16625 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14979) );
  NAND2_X1 U16626 ( .A1(n14544), .A2(n14979), .ZN(n13405) );
  NAND3_X1 U16627 ( .A1(n13406), .A2(n14641), .A3(n13405), .ZN(n13407) );
  OAI21_X1 U16628 ( .B1(n13408), .B2(P1_EBX_REG_27__SCAN_IN), .A(n13407), .ZN(
        n14684) );
  NAND2_X1 U16629 ( .A1(n14683), .A2(n14684), .ZN(n14518) );
  MUX2_X1 U16630 ( .A(n13317), .B(n14641), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n13409) );
  OAI21_X1 U16631 ( .B1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n14551), .A(
        n13409), .ZN(n14519) );
  NAND2_X1 U16632 ( .A1(n14551), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n13411) );
  NAND2_X1 U16633 ( .A1(n14550), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13410) );
  NAND2_X1 U16634 ( .A1(n13411), .A2(n13410), .ZN(n14659) );
  XNOR2_X1 U16635 ( .A(n14659), .B(n14641), .ZN(n14546) );
  NAND2_X1 U16636 ( .A1(n17135), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13420) );
  NAND2_X1 U16637 ( .A1(READY11_REG_SCAN_IN), .A2(READY1), .ZN(n21221) );
  AND2_X1 U16638 ( .A1(n21221), .A2(n21022), .ZN(n17137) );
  NOR2_X1 U16639 ( .A1(n13420), .A2(n17137), .ZN(n13412) );
  INV_X1 U16640 ( .A(n13413), .ZN(n13414) );
  NAND2_X1 U16641 ( .A1(n13414), .A2(n21137), .ZN(n17153) );
  INV_X1 U16642 ( .A(n17137), .ZN(n13415) );
  AOI21_X1 U16643 ( .B1(n20603), .B2(n17153), .A(n13415), .ZN(n13422) );
  NAND2_X2 U16644 ( .A1(n13424), .A2(n13422), .ZN(n20420) );
  INV_X1 U16645 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n14695) );
  INV_X1 U16646 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n14718) );
  INV_X1 U16647 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n21162) );
  INV_X1 U16648 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n21160) );
  INV_X1 U16649 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21157) );
  NAND3_X1 U16650 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n20422) );
  NOR2_X1 U16651 ( .A1(n21157), .A2(n20422), .ZN(n20419) );
  NAND2_X1 U16652 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n20419), .ZN(n20395) );
  NOR2_X1 U16653 ( .A1(n21160), .A2(n20395), .ZN(n20396) );
  NAND2_X1 U16654 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20396), .ZN(n20366) );
  NOR2_X1 U16655 ( .A1(n21162), .A2(n20366), .ZN(n14837) );
  NAND2_X1 U16656 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n14832) );
  NAND4_X1 U16657 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .A3(P1_REIP_REG_12__SCAN_IN), .A4(P1_REIP_REG_11__SCAN_IN), .ZN(n14855) );
  NAND2_X1 U16658 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n14841) );
  NOR3_X1 U16659 ( .A1(n14832), .A2(n14855), .A3(n14841), .ZN(n14818) );
  AND2_X1 U16660 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n14818), .ZN(n13416) );
  NAND2_X1 U16661 ( .A1(n14837), .A2(n13416), .ZN(n14795) );
  NAND2_X1 U16662 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n13417) );
  OR2_X1 U16663 ( .A1(n14795), .A2(n13417), .ZN(n14777) );
  INV_X1 U16664 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n13418) );
  NOR2_X1 U16665 ( .A1(n14777), .A2(n13418), .ZN(n14751) );
  AND2_X1 U16666 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n13419) );
  AND2_X1 U16667 ( .A1(n14751), .A2(n13419), .ZN(n14738) );
  NAND2_X1 U16668 ( .A1(n14738), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n14726) );
  INV_X1 U16669 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n14731) );
  OR2_X1 U16670 ( .A1(n14726), .A2(n14731), .ZN(n14694) );
  NOR3_X1 U16671 ( .A1(n14695), .A2(n14718), .A3(n14694), .ZN(n13430) );
  NAND2_X1 U16672 ( .A1(n20376), .A2(n13430), .ZN(n14682) );
  NAND2_X1 U16673 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(P1_REIP_REG_27__SCAN_IN), 
        .ZN(n13431) );
  INV_X1 U16674 ( .A(n13420), .ZN(n13421) );
  NOR2_X1 U16675 ( .A1(n13422), .A2(n13421), .ZN(n13423) );
  NAND2_X1 U16676 ( .A1(n13424), .A2(n13423), .ZN(n20424) );
  INV_X1 U16677 ( .A(n13425), .ZN(n13426) );
  OAI22_X1 U16678 ( .A1(n9611), .A2(n15116), .B1(n13427), .B2(n20407), .ZN(
        n13428) );
  AOI21_X1 U16679 ( .B1(P1_EBX_REG_29__SCAN_IN), .B2(n20405), .A(n13428), .ZN(
        n13429) );
  OAI21_X1 U16680 ( .B1(P1_REIP_REG_29__SCAN_IN), .B2(n14667), .A(n13429), 
        .ZN(n13434) );
  NAND2_X1 U16681 ( .A1(n20410), .A2(n13430), .ZN(n14678) );
  NAND2_X1 U16682 ( .A1(n20420), .A2(n20410), .ZN(n14835) );
  OAI21_X1 U16683 ( .B1(n13431), .B2(n14678), .A(n14835), .ZN(n14589) );
  INV_X1 U16684 ( .A(n14589), .ZN(n13432) );
  NAND2_X1 U16685 ( .A1(n16850), .A2(n13630), .ZN(n13896) );
  INV_X1 U16686 ( .A(n20309), .ZN(n13628) );
  AND2_X1 U16687 ( .A1(n13436), .A2(n20272), .ZN(n13437) );
  AND2_X1 U16688 ( .A1(n14228), .A2(n13437), .ZN(n16865) );
  NOR2_X1 U16689 ( .A1(n14634), .A2(n19407), .ZN(n13497) );
  NOR2_X1 U16690 ( .A1(n13440), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13441) );
  OR2_X1 U16691 ( .A1(n13460), .A2(n13441), .ZN(n16304) );
  AND2_X1 U16692 ( .A1(n13455), .A2(n16328), .ZN(n13442) );
  OR2_X1 U16693 ( .A1(n13442), .A2(n13457), .ZN(n13576) );
  NOR2_X1 U16694 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n13452), .ZN(
        n13444) );
  NOR2_X1 U16695 ( .A1(n13443), .A2(n13444), .ZN(n16346) );
  AOI21_X1 U16696 ( .B1(n16368), .B2(n13450), .A(n13454), .ZN(n16370) );
  AOI21_X1 U16697 ( .B1(n13445), .B2(n16399), .A(n13451), .ZN(n16401) );
  AOI21_X1 U16698 ( .B1(n17199), .B2(n13447), .A(n13449), .ZN(n17191) );
  AOI21_X1 U16699 ( .B1(n16420), .B2(n13446), .A(n13448), .ZN(n15927) );
  OAI21_X1 U16700 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n13446), .ZN(n15941) );
  MUX2_X1 U16701 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n16773) );
  INV_X1 U16702 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13648) );
  MUX2_X1 U16703 ( .A(n13648), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n15954) );
  OAI21_X1 U16704 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n13448), .A(
        n13447), .ZN(n19581) );
  NOR2_X1 U16705 ( .A1(n17191), .A2(n15914), .ZN(n15898) );
  OAI21_X1 U16706 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n13449), .A(
        n13445), .ZN(n16409) );
  NAND2_X1 U16707 ( .A1(n15898), .A2(n16409), .ZN(n15887) );
  OAI21_X1 U16708 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n13451), .A(
        n13450), .ZN(n16387) );
  INV_X1 U16709 ( .A(n9685), .ZN(n15846) );
  INV_X1 U16710 ( .A(n13452), .ZN(n13453) );
  OAI21_X1 U16711 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n13454), .A(
        n13453), .ZN(n16359) );
  OAI21_X1 U16712 ( .B1(n13443), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n13455), .ZN(n16337) );
  INV_X1 U16713 ( .A(n13577), .ZN(n13456) );
  AND2_X1 U16714 ( .A1(n13576), .A2(n13456), .ZN(n15797) );
  NOR2_X1 U16715 ( .A1(n13457), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13458) );
  OR2_X1 U16716 ( .A1(n13440), .A2(n13458), .ZN(n16315) );
  NAND2_X1 U16717 ( .A1(n15797), .A2(n16315), .ZN(n19388) );
  INV_X1 U16718 ( .A(n19388), .ZN(n13459) );
  OAI21_X1 U16719 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n13460), .A(
        n9658), .ZN(n16293) );
  OAI21_X1 U16720 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n13462), .A(
        n13461), .ZN(n16285) );
  NOR2_X1 U16721 ( .A1(n15740), .A2(n15741), .ZN(n15723) );
  NAND2_X1 U16722 ( .A1(n15723), .A2(n15725), .ZN(n15722) );
  AOI21_X1 U16723 ( .B1(n16274), .B2(n13463), .A(n13464), .ZN(n16276) );
  NOR2_X1 U16724 ( .A1(n15722), .A2(n16276), .ZN(n15698) );
  OAI21_X1 U16725 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n13464), .A(
        n13466), .ZN(n16260) );
  NAND2_X1 U16726 ( .A1(n15698), .A2(n16260), .ZN(n13465) );
  INV_X1 U16727 ( .A(n13466), .ZN(n13468) );
  INV_X1 U16728 ( .A(n13467), .ZN(n13470) );
  OAI21_X1 U16729 ( .B1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n13468), .A(
        n13470), .ZN(n16245) );
  NAND2_X1 U16730 ( .A1(n15677), .A2(n16245), .ZN(n15668) );
  INV_X1 U16731 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n13471) );
  INV_X1 U16732 ( .A(n13469), .ZN(n13473) );
  AOI21_X1 U16733 ( .B1(n13471), .B2(n13470), .A(n13473), .ZN(n16239) );
  INV_X1 U16734 ( .A(n13472), .ZN(n13474) );
  OAI21_X1 U16735 ( .B1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n13473), .A(
        n13474), .ZN(n16228) );
  INV_X1 U16736 ( .A(n15637), .ZN(n13476) );
  AOI21_X1 U16737 ( .B1(n16218), .B2(n13474), .A(n13479), .ZN(n16220) );
  INV_X1 U16738 ( .A(n16220), .ZN(n13475) );
  NAND2_X1 U16739 ( .A1(n13476), .A2(n13475), .ZN(n13477) );
  INV_X1 U16740 ( .A(n13478), .ZN(n13482) );
  INV_X1 U16741 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15625) );
  INV_X1 U16742 ( .A(n13479), .ZN(n13480) );
  NAND2_X1 U16743 ( .A1(n15625), .A2(n13480), .ZN(n13481) );
  NAND2_X1 U16744 ( .A1(n13482), .A2(n13481), .ZN(n16210) );
  INV_X1 U16745 ( .A(n16761), .ZN(n19416) );
  OAI21_X1 U16746 ( .B1(n14603), .B2(n19416), .A(n14602), .ZN(n14604) );
  INV_X1 U16747 ( .A(n13483), .ZN(n13484) );
  NOR2_X1 U16748 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13777) );
  NOR2_X1 U16749 ( .A1(n13485), .A2(n13629), .ZN(n13486) );
  AND2_X1 U16750 ( .A1(n14228), .A2(n20272), .ZN(n13487) );
  NOR2_X1 U16751 ( .A1(n14059), .A2(n13487), .ZN(n13581) );
  NOR2_X1 U16752 ( .A1(n20306), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19741) );
  NAND2_X1 U16753 ( .A1(n13626), .A2(n19741), .ZN(n17233) );
  AND3_X1 U16754 ( .A1(n19417), .A2(n17200), .A3(n17233), .ZN(n13488) );
  AOI22_X1 U16755 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n13581), .B1(n19410), 
        .B2(P2_REIP_REG_31__SCAN_IN), .ZN(n13490) );
  NAND2_X1 U16756 ( .A1(n19404), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13489) );
  OAI211_X1 U16757 ( .C1(n14604), .C2(n19386), .A(n13490), .B(n13489), .ZN(
        n13495) );
  NAND2_X1 U16758 ( .A1(n20191), .A2(n20272), .ZN(n13491) );
  AND2_X1 U16759 ( .A1(n13633), .A2(n13491), .ZN(n13579) );
  AND2_X1 U16760 ( .A1(n15992), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n13492) );
  NOR2_X1 U16761 ( .A1(n13497), .A2(n13496), .ZN(n13500) );
  AND2_X1 U16762 ( .A1(n10884), .A2(n20191), .ZN(n13498) );
  NAND2_X1 U16763 ( .A1(n13500), .A2(n13499), .ZN(P2_U2824) );
  XNOR2_X1 U16764 ( .A(n13501), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15107) );
  AOI22_X1 U16765 ( .A1(n13502), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13088), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13509) );
  AOI22_X1 U16766 ( .A1(n13043), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13503), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13508) );
  AOI22_X1 U16767 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13504), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13507) );
  AOI22_X1 U16768 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12382), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13506) );
  NAND4_X1 U16769 ( .A1(n13509), .A2(n13508), .A3(n13507), .A4(n13506), .ZN(
        n13519) );
  AOI22_X1 U16770 ( .A1(n13510), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9623), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13517) );
  AOI22_X1 U16771 ( .A1(n13512), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n13511), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13516) );
  AOI22_X1 U16772 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9591), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13515) );
  NAND4_X1 U16773 ( .A1(n13517), .A2(n13516), .A3(n13515), .A4(n13514), .ZN(
        n13518) );
  NOR2_X1 U16774 ( .A1(n13519), .A2(n13518), .ZN(n13523) );
  NOR2_X1 U16775 ( .A1(n13521), .A2(n13520), .ZN(n13522) );
  XNOR2_X1 U16776 ( .A(n13523), .B(n13522), .ZN(n13529) );
  INV_X1 U16777 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n15016) );
  NAND2_X1 U16778 ( .A1(n21070), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13525) );
  OAI211_X1 U16779 ( .C1(n13526), .C2(n15016), .A(n13525), .B(n13524), .ZN(
        n13527) );
  AOI21_X1 U16780 ( .B1(n13529), .B2(n13528), .A(n13527), .ZN(n13530) );
  AOI22_X1 U16781 ( .A1(n12668), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n13532), .ZN(n13533) );
  INV_X1 U16782 ( .A(n13533), .ZN(n13534) );
  NAND2_X1 U16783 ( .A1(n13876), .A2(n12437), .ZN(n14646) );
  INV_X1 U16784 ( .A(n13535), .ZN(n13536) );
  NOR2_X1 U16785 ( .A1(n13536), .A2(n21142), .ZN(n14467) );
  NAND2_X1 U16786 ( .A1(n14467), .A2(n14544), .ZN(n13537) );
  NAND4_X1 U16787 ( .A1(n13538), .A2(n12319), .A3(n13950), .A4(n20626), .ZN(
        n13912) );
  NAND2_X1 U16788 ( .A1(n21221), .A2(n14650), .ZN(n14471) );
  OR2_X1 U16789 ( .A1(n13539), .A2(n14471), .ZN(n13877) );
  OAI21_X1 U16790 ( .B1(n13912), .B2(n14640), .A(n13877), .ZN(n13540) );
  INV_X1 U16791 ( .A(n13540), .ZN(n13541) );
  NAND2_X1 U16792 ( .A1(n14588), .A2(n13544), .ZN(n13560) );
  INV_X1 U16793 ( .A(n13871), .ZN(n14468) );
  NOR4_X1 U16794 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n13548) );
  NOR4_X1 U16795 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n13547) );
  NOR4_X1 U16796 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13546) );
  NOR4_X1 U16797 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n13545) );
  AND4_X1 U16798 ( .A1(n13548), .A2(n13547), .A3(n13546), .A4(n13545), .ZN(
        n13554) );
  NOR4_X1 U16799 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n13552) );
  NOR4_X1 U16800 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n13551) );
  NOR4_X1 U16801 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n13550) );
  INV_X1 U16802 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n13549) );
  AND4_X1 U16803 ( .A1(n13552), .A2(n13551), .A3(n13550), .A4(n13549), .ZN(
        n13553) );
  NAND2_X1 U16804 ( .A1(n13554), .A2(n13553), .ZN(n13555) );
  AOI22_X1 U16805 ( .A1(n15082), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n15076), .ZN(n13556) );
  INV_X1 U16806 ( .A(n13556), .ZN(n13558) );
  INV_X1 U16807 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n19643) );
  NOR2_X1 U16808 ( .A1(n15080), .A2(n19643), .ZN(n13557) );
  NOR2_X1 U16809 ( .A1(n13558), .A2(n13557), .ZN(n13559) );
  NAND2_X1 U16810 ( .A1(n13560), .A2(n13559), .ZN(P1_U2873) );
  NOR2_X1 U16811 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13562) );
  NOR4_X1 U16812 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13561) );
  NAND4_X1 U16813 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13562), .A4(n13561), .ZN(n13575) );
  INV_X1 U16814 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21213) );
  NOR3_X1 U16815 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n21213), .ZN(n13564) );
  NOR4_X1 U16816 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13563) );
  NAND4_X1 U16817 ( .A1(n20584), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13564), .A4(
        n13563), .ZN(U214) );
  NOR4_X1 U16818 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n13568) );
  NOR4_X1 U16819 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n13567) );
  NOR4_X1 U16820 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n13566) );
  NOR4_X1 U16821 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n13565) );
  AND4_X1 U16822 ( .A1(n13568), .A2(n13567), .A3(n13566), .A4(n13565), .ZN(
        n13573) );
  NOR4_X1 U16823 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n13571) );
  NOR4_X1 U16824 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n13570) );
  NOR4_X1 U16825 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n13569) );
  INV_X1 U16826 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20212) );
  AND4_X1 U16827 ( .A1(n13571), .A2(n13570), .A3(n13569), .A4(n20212), .ZN(
        n13572) );
  NAND2_X1 U16828 ( .A1(n13573), .A2(n13572), .ZN(n13574) );
  NOR2_X1 U16829 ( .A1(n19430), .A2(n13575), .ZN(n17268) );
  NAND2_X1 U16830 ( .A1(n17268), .A2(U214), .ZN(U212) );
  INV_X1 U16831 ( .A(n13576), .ZN(n16326) );
  AOI211_X1 U16832 ( .C1(n16326), .C2(n13577), .A(n15797), .B(n19386), .ZN(
        n13594) );
  INV_X1 U16833 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n13578) );
  AND2_X1 U16834 ( .A1(n13579), .A2(n13578), .ZN(n13580) );
  OAI22_X1 U16835 ( .A1(n19392), .A2(n11172), .B1(n16328), .B2(n19389), .ZN(
        n13593) );
  AOI22_X1 U16836 ( .A1(n13582), .A2(n15968), .B1(n19400), .B2(n16326), .ZN(
        n13583) );
  OAI211_X1 U16837 ( .C1(n20228), .C2(n15958), .A(n13583), .B(n17200), .ZN(
        n13592) );
  AOI21_X1 U16838 ( .B1(n13585), .B2(n15810), .A(n13584), .ZN(n16621) );
  INV_X1 U16839 ( .A(n16621), .ZN(n13590) );
  NAND2_X1 U16840 ( .A1(n14283), .A2(n13588), .ZN(n13589) );
  NAND2_X1 U16841 ( .A1(n13586), .A2(n13589), .ZN(n16616) );
  OAI22_X1 U16842 ( .A1(n13590), .A2(n15911), .B1(n16616), .B2(n19407), .ZN(
        n13591) );
  NAND2_X1 U16843 ( .A1(n14272), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17012) );
  NAND2_X1 U16844 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16991) );
  INV_X1 U16845 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n18421) );
  INV_X1 U16846 ( .A(n18352), .ZN(n18367) );
  NAND2_X1 U16847 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18373) );
  NAND2_X1 U16848 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16966) );
  NAND2_X1 U16849 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n18316) );
  NOR2_X1 U16850 ( .A1(n17709), .A2(n13596), .ZN(n13604) );
  AND2_X1 U16851 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n13604), .ZN(
        n13597) );
  NAND2_X1 U16852 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n18277) );
  NAND2_X1 U16853 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16949), .ZN(
        n16956) );
  OAI21_X1 U16854 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n13597), .A(
        n16956), .ZN(n13598) );
  INV_X1 U16855 ( .A(n13598), .ZN(n18276) );
  NAND2_X1 U16856 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n18251) );
  NAND2_X1 U16857 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n13600) );
  INV_X1 U16858 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n17412) );
  INV_X4 U16859 ( .A(n16881), .ZN(n17695) );
  NAND2_X1 U16860 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18301), .ZN(
        n13603) );
  INV_X1 U16861 ( .A(n13603), .ZN(n18273) );
  INV_X1 U16862 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n17728) );
  INV_X1 U16863 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n18303) );
  AOI21_X1 U16864 ( .B1(n18303), .B2(n13603), .A(n13604), .ZN(n18306) );
  INV_X1 U16865 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18291) );
  XNOR2_X1 U16866 ( .A(n18291), .B(n13604), .ZN(n18288) );
  NOR2_X1 U16867 ( .A1(n17485), .A2(n17695), .ZN(n13605) );
  NOR2_X1 U16868 ( .A1(n13605), .A2(n18276), .ZN(n17382) );
  INV_X1 U16869 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n21312) );
  NAND4_X1 U16870 ( .A1(n19349), .A2(n19338), .A3(n21312), .A4(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n17712) );
  AOI211_X1 U16871 ( .C1(n18276), .C2(n13605), .A(n17382), .B(n9767), .ZN(
        n13620) );
  INV_X1 U16872 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n18000) );
  NAND2_X1 U16873 ( .A1(n17708), .A2(n18000), .ZN(n17689) );
  NOR2_X2 U16874 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17689), .ZN(n17688) );
  NAND2_X1 U16875 ( .A1(n17688), .A2(n17992), .ZN(n17678) );
  NOR2_X2 U16876 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17678), .ZN(n17659) );
  NAND2_X1 U16877 ( .A1(n17659), .A2(n17653), .ZN(n17652) );
  NAND2_X1 U16878 ( .A1(n17631), .A2(n21250), .ZN(n17608) );
  NOR2_X2 U16879 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17608), .ZN(n17607) );
  NAND2_X1 U16880 ( .A1(n17607), .A2(n17604), .ZN(n17603) );
  INV_X1 U16881 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17582) );
  NAND2_X1 U16882 ( .A1(n17587), .A2(n17582), .ZN(n17581) );
  NOR2_X2 U16883 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17581), .ZN(n17561) );
  INV_X1 U16884 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n21278) );
  NAND2_X1 U16885 ( .A1(n17561), .A2(n21278), .ZN(n17557) );
  INV_X1 U16886 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17534) );
  NAND2_X1 U16887 ( .A1(n17542), .A2(n17534), .ZN(n17533) );
  NOR2_X2 U16888 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17533), .ZN(n17519) );
  INV_X1 U16889 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n17510) );
  NOR2_X2 U16890 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17509), .ZN(n17495) );
  INV_X1 U16891 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17927) );
  NAND2_X1 U16892 ( .A1(n17495), .A2(n17927), .ZN(n17487) );
  NOR2_X2 U16893 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17487), .ZN(n17481) );
  INV_X1 U16894 ( .A(n13606), .ZN(n13607) );
  NAND2_X1 U16895 ( .A1(n19335), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n13611) );
  AOI211_X4 U16896 ( .C1(n19222), .C2(n21312), .A(n13614), .B(n13611), .ZN(
        n17724) );
  AOI211_X1 U16897 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n17487), .A(n17481), .B(
        n17687), .ZN(n13619) );
  NAND2_X1 U16898 ( .A1(n19349), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19109) );
  INV_X1 U16899 ( .A(n19109), .ZN(n19225) );
  INV_X1 U16900 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n19223) );
  NAND3_X1 U16901 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19225), .A3(n19223), 
        .ZN(n19218) );
  NAND3_X1 U16902 ( .A1(n19218), .A2(n18739), .A3(n17712), .ZN(n13609) );
  AND2_X1 U16903 ( .A1(n19222), .A2(n21312), .ZN(n13610) );
  OAI21_X1 U16904 ( .B1(n19334), .B2(n19335), .A(n13610), .ZN(n19211) );
  NAND2_X1 U16905 ( .A1(n19211), .A2(n13611), .ZN(n13612) );
  AOI22_X1 U16906 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17700), .B1(
        n17725), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n13613) );
  INV_X1 U16907 ( .A(n13613), .ZN(n13618) );
  INV_X1 U16908 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n19285) );
  INV_X1 U16909 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n19286) );
  INV_X1 U16910 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n19283) );
  NOR3_X1 U16911 ( .A1(n19285), .A2(n19286), .A3(n19283), .ZN(n13615) );
  INV_X1 U16912 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n19279) );
  INV_X1 U16913 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n19277) );
  INV_X1 U16914 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n19269) );
  INV_X1 U16915 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n19257) );
  NAND2_X1 U16916 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n17716) );
  NOR2_X1 U16917 ( .A1(n21313), .A2(n17716), .ZN(n17686) );
  NAND2_X1 U16918 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n17686), .ZN(n17672) );
  NOR2_X1 U16919 ( .A1(n19257), .A2(n17672), .ZN(n17657) );
  AND3_X1 U16920 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .A3(n17657), .ZN(n17640) );
  NAND2_X1 U16921 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n17640), .ZN(n17630) );
  INV_X1 U16922 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n19267) );
  INV_X1 U16923 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n19265) );
  NAND3_X1 U16924 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(P3_REIP_REG_13__SCAN_IN), 
        .A3(n17572), .ZN(n17564) );
  NOR3_X1 U16925 ( .A1(n19279), .A2(n19277), .A3(n17564), .ZN(n17525) );
  NAND2_X1 U16926 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n17525), .ZN(n17379) );
  NOR2_X1 U16927 ( .A1(n17729), .A2(n17379), .ZN(n17517) );
  NAND2_X1 U16928 ( .A1(n13615), .A2(n17517), .ZN(n17492) );
  INV_X1 U16929 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n19289) );
  XOR2_X1 U16930 ( .A(P3_REIP_REG_22__SCAN_IN), .B(n19289), .Z(n13616) );
  INV_X1 U16931 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n19290) );
  INV_X1 U16932 ( .A(n13615), .ZN(n17378) );
  OR2_X1 U16933 ( .A1(n17379), .A2(n17721), .ZN(n17502) );
  NOR2_X1 U16934 ( .A1(n17658), .A2(n17721), .ZN(n17673) );
  OAI21_X1 U16935 ( .B1(n17378), .B2(n17502), .A(n17645), .ZN(n17501) );
  OAI22_X1 U16936 ( .A1(n17492), .A2(n13616), .B1(n19290), .B2(n17501), .ZN(
        n13617) );
  OR4_X1 U16937 ( .A1(n13620), .A2(n13619), .A3(n13618), .A4(n13617), .ZN(
        P3_U2649) );
  NOR3_X1 U16938 ( .A1(n20191), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n13438), 
        .ZN(n17234) );
  AND3_X1 U16939 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .A3(P2_STATE2_REG_2__SCAN_IN), .ZN(n17244) );
  NOR3_X1 U16940 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n13621) );
  NOR4_X1 U16941 ( .A1(n17234), .A2(n20319), .A3(n17244), .A4(n13621), .ZN(
        P2_U3178) );
  INV_X1 U16942 ( .A(n13896), .ZN(n13623) );
  NAND2_X1 U16943 ( .A1(n10895), .A2(n20191), .ZN(n13895) );
  INV_X1 U16944 ( .A(n14228), .ZN(n13622) );
  NAND3_X1 U16945 ( .A1(n13623), .A2(n13895), .A3(n13622), .ZN(n16856) );
  AND2_X1 U16946 ( .A1(n16856), .A2(n17236), .ZN(n20303) );
  OAI21_X1 U16947 ( .B1(n20303), .B2(n13625), .A(n13624), .ZN(P2_U2819) );
  INV_X1 U16948 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n21283) );
  INV_X1 U16949 ( .A(n20305), .ZN(n20268) );
  INV_X1 U16950 ( .A(n13626), .ZN(n13627) );
  OAI22_X1 U16951 ( .A1(n13628), .A2(n21283), .B1(n20268), .B2(n13627), .ZN(
        P2_U2816) );
  NOR2_X1 U16952 ( .A1(n10857), .A2(n13629), .ZN(n13708) );
  NAND2_X1 U16953 ( .A1(n13708), .A2(n13630), .ZN(n19412) );
  INV_X1 U16954 ( .A(P2_READREQUEST_REG_SCAN_IN), .ZN(n13631) );
  NAND2_X1 U16955 ( .A1(n19412), .A2(n13631), .ZN(n13634) );
  AND2_X1 U16956 ( .A1(n20305), .A2(n10955), .ZN(n13632) );
  OR2_X1 U16957 ( .A1(n13633), .A2(n13632), .ZN(n19356) );
  OAI22_X1 U16958 ( .A1(n13634), .A2(n19356), .B1(n20309), .B2(n10895), .ZN(
        n13635) );
  INV_X1 U16959 ( .A(n13635), .ZN(P2_U3612) );
  AND2_X1 U16960 ( .A1(n21383), .A2(n13636), .ZN(n14790) );
  AOI21_X1 U16961 ( .B1(n13637), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n14790), 
        .ZN(n13638) );
  NAND2_X1 U16962 ( .A1(n14372), .A2(n13638), .ZN(P1_U2801) );
  OAI21_X1 U16963 ( .B1(n13640), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n13639), .ZN(n16743) );
  INV_X1 U16964 ( .A(n13641), .ZN(n13643) );
  NAND2_X1 U16965 ( .A1(n13643), .A2(n13642), .ZN(n13644) );
  XNOR2_X1 U16966 ( .A(n13644), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16748) );
  AOI22_X1 U16967 ( .A1(n19586), .A2(n16748), .B1(n19584), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13646) );
  AND2_X1 U16968 ( .A1(n19571), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n16747) );
  INV_X1 U16969 ( .A(n16747), .ZN(n13645) );
  OAI211_X1 U16970 ( .C1(n16743), .C2(n19590), .A(n13646), .B(n13645), .ZN(
        n13647) );
  AOI21_X1 U16971 ( .B1(n17192), .B2(n13648), .A(n13647), .ZN(n13649) );
  OAI21_X1 U16972 ( .B1(n11572), .B2(n19573), .A(n13649), .ZN(P2_U3013) );
  AOI22_X1 U16973 ( .A1(n17975), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17974), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13653) );
  AOI22_X1 U16974 ( .A1(n17903), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17973), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13652) );
  NAND2_X1 U16975 ( .A1(n13685), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n13651) );
  NAND2_X1 U16976 ( .A1(n17818), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n13650) );
  NAND4_X1 U16977 ( .A1(n13653), .A2(n13652), .A3(n13651), .A4(n13650), .ZN(
        n13656) );
  INV_X1 U16978 ( .A(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13654) );
  OAI22_X1 U16979 ( .A1(n13654), .A2(n9568), .B1(n17981), .B2(n11954), .ZN(
        n13655) );
  OR2_X1 U16980 ( .A1(n13656), .A2(n13655), .ZN(n13664) );
  AOI22_X1 U16981 ( .A1(n17966), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17954), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13662) );
  AOI22_X1 U16982 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9581), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13661) );
  AOI22_X1 U16983 ( .A1(n14172), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13660) );
  AOI22_X1 U16984 ( .A1(n9576), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17967), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13659) );
  NAND4_X1 U16985 ( .A1(n13662), .A2(n13661), .A3(n13660), .A4(n13659), .ZN(
        n13663) );
  NOR2_X1 U16986 ( .A1(n13664), .A2(n13663), .ZN(n14237) );
  INV_X1 U16987 ( .A(n13665), .ZN(n13666) );
  NAND3_X1 U16988 ( .A1(n17863), .A2(n18770), .A3(n13666), .ZN(n13668) );
  NAND2_X1 U16989 ( .A1(n13667), .A2(n19180), .ZN(n13723) );
  NAND2_X1 U16990 ( .A1(n13668), .A2(n13723), .ZN(n13928) );
  AND3_X1 U16991 ( .A1(n18755), .A2(n19214), .A3(n19335), .ZN(n13669) );
  INV_X1 U16992 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n14193) );
  INV_X1 U16993 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n17705) );
  NAND2_X1 U16994 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17722) );
  NOR2_X1 U16995 ( .A1(n17705), .A2(n17722), .ZN(n17996) );
  NAND4_X2 U16996 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n18007), .A4(n17996), .ZN(n17995) );
  NAND4_X1 U16997 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(P3_EBX_REG_7__SCAN_IN), 
        .A3(P3_EBX_REG_6__SCAN_IN), .A4(P3_EBX_REG_5__SCAN_IN), .ZN(n13670) );
  NAND3_X1 U16998 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(P3_EBX_REG_8__SCAN_IN), 
        .A3(n13671), .ZN(n13675) );
  INV_X1 U16999 ( .A(n13675), .ZN(n13672) );
  INV_X1 U17000 ( .A(n18007), .ZN(n18015) );
  NOR2_X1 U17001 ( .A1(n18783), .A2(n18015), .ZN(n18011) );
  INV_X1 U17002 ( .A(n18011), .ZN(n18018) );
  OAI22_X1 U17003 ( .A1(n18016), .A2(n13672), .B1(P3_EBX_REG_13__SCAN_IN), 
        .B2(n18018), .ZN(n17986) );
  OAI21_X1 U17004 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n13672), .A(n17986), .ZN(
        n13673) );
  OAI21_X1 U17005 ( .B1(n14237), .B2(n18013), .A(n13673), .ZN(P3_U2690) );
  NAND3_X1 U17006 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_14__SCAN_IN), 
        .A3(P3_EBX_REG_13__SCAN_IN), .ZN(n14194) );
  NOR2_X1 U17007 ( .A1(n18016), .A2(n13835), .ZN(n14196) );
  NAND2_X1 U17008 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(P3_EBX_REG_13__SCAN_IN), 
        .ZN(n13674) );
  OAI21_X1 U17009 ( .B1(n13675), .B2(n13674), .A(n21278), .ZN(n13693) );
  AOI22_X1 U17010 ( .A1(n17966), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17954), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13680) );
  AOI22_X1 U17011 ( .A1(n9572), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9582), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13679) );
  AOI22_X1 U17012 ( .A1(n14172), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13678) );
  AOI22_X1 U17013 ( .A1(n9577), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17967), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13677) );
  NAND4_X1 U17014 ( .A1(n13680), .A2(n13679), .A3(n13678), .A4(n13677), .ZN(
        n13692) );
  INV_X1 U17015 ( .A(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13683) );
  AOI22_X1 U17016 ( .A1(n12119), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17973), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13682) );
  NAND2_X1 U17017 ( .A1(n11937), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n13681) );
  OAI211_X1 U17018 ( .C1(n13684), .C2(n13683), .A(n13682), .B(n13681), .ZN(
        n13691) );
  INV_X1 U17019 ( .A(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13687) );
  OAI22_X1 U17020 ( .A1(n13687), .A2(n17931), .B1(n12101), .B2(n13686), .ZN(
        n13690) );
  INV_X1 U17021 ( .A(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17795) );
  OAI22_X1 U17022 ( .A1(n13688), .A2(n17981), .B1(n17844), .B2(n17795), .ZN(
        n13689) );
  OR4_X1 U17023 ( .A1(n13692), .A2(n13691), .A3(n13690), .A4(n13689), .ZN(
        n18086) );
  AOI22_X1 U17024 ( .A1(n14196), .A2(n13693), .B1(n18016), .B2(n18086), .ZN(
        n13694) );
  INV_X1 U17025 ( .A(n13694), .ZN(P3_U2688) );
  INV_X1 U17026 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17991) );
  NOR4_X1 U17027 ( .A1(n17653), .A2(n17991), .A3(n17992), .A4(n17995), .ZN(
        n14511) );
  NAND2_X1 U17028 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n14511), .ZN(n13732) );
  OAI21_X1 U17029 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n14511), .A(n13732), .ZN(
        n13707) );
  AOI22_X1 U17030 ( .A1(n17966), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17954), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13698) );
  AOI22_X1 U17031 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9580), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13697) );
  AOI22_X1 U17032 ( .A1(n14172), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13696) );
  AOI22_X1 U17033 ( .A1(n9578), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17967), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13695) );
  NAND4_X1 U17034 ( .A1(n13698), .A2(n13697), .A3(n13696), .A4(n13695), .ZN(
        n13705) );
  AOI22_X1 U17035 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17818), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13701) );
  AOI22_X1 U17036 ( .A1(n17903), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17973), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13700) );
  AOI22_X1 U17037 ( .A1(n17975), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17974), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13699) );
  NAND3_X1 U17038 ( .A1(n13701), .A2(n13700), .A3(n13699), .ZN(n13704) );
  INV_X1 U17039 ( .A(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14169) );
  OAI22_X1 U17040 ( .A1(n17844), .A2(n14169), .B1(n17981), .B2(n13702), .ZN(
        n13703) );
  OR3_X1 U17041 ( .A1(n13705), .A2(n13704), .A3(n13703), .ZN(n18103) );
  NAND2_X1 U17042 ( .A1(n18016), .A2(n18103), .ZN(n13706) );
  OAI21_X1 U17043 ( .B1(n13707), .B2(n18016), .A(n13706), .ZN(P3_U2695) );
  INV_X1 U17044 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n13715) );
  INV_X1 U17045 ( .A(n13708), .ZN(n13709) );
  OAI21_X1 U17046 ( .B1(n13710), .B2(n13709), .A(n14059), .ZN(n13711) );
  INV_X1 U17047 ( .A(n13713), .ZN(n20312) );
  INV_X1 U17048 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n21346) );
  INV_X1 U17049 ( .A(P2_UWORD_REG_12__SCAN_IN), .ZN(n13714) );
  OAI222_X1 U17050 ( .A1(n13715), .A2(n19492), .B1(n13794), .B2(n21346), .C1(
        n20310), .C2(n13714), .ZN(P2_U2923) );
  INV_X1 U17051 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n13717) );
  INV_X1 U17052 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n14056) );
  INV_X1 U17053 ( .A(P2_UWORD_REG_11__SCAN_IN), .ZN(n13716) );
  OAI222_X1 U17054 ( .A1(n13717), .A2(n19492), .B1(n13794), .B2(n14056), .C1(
        n20310), .C2(n13716), .ZN(P2_U2924) );
  INV_X1 U17055 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n13719) );
  INV_X1 U17056 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n14050) );
  INV_X1 U17057 ( .A(P2_UWORD_REG_9__SCAN_IN), .ZN(n13718) );
  OAI222_X1 U17058 ( .A1(n13719), .A2(n19492), .B1(n13794), .B2(n14050), .C1(
        n20310), .C2(n13718), .ZN(P2_U2926) );
  INV_X1 U17059 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19438) );
  INV_X1 U17060 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n17330) );
  INV_X1 U17061 ( .A(P2_LWORD_REG_11__SCAN_IN), .ZN(n21298) );
  OAI222_X1 U17062 ( .A1(n19523), .A2(n19438), .B1(n19492), .B2(n17330), .C1(
        n20310), .C2(n21298), .ZN(P2_U2940) );
  INV_X1 U17063 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13720) );
  INV_X1 U17064 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n17336) );
  INV_X1 U17065 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n21331) );
  OAI222_X1 U17066 ( .A1(n13794), .A2(n13720), .B1(n19492), .B2(n17336), .C1(
        n20310), .C2(n21331), .ZN(P2_U2934) );
  NAND2_X1 U17067 ( .A1(n19185), .A2(n19222), .ZN(n13725) );
  NAND2_X1 U17068 ( .A1(n13722), .A2(n19334), .ZN(n18127) );
  OAI211_X1 U17069 ( .C1(n13725), .C2(n18127), .A(n13724), .B(n13723), .ZN(
        n13726) );
  NOR2_X1 U17070 ( .A1(n13929), .A2(n13726), .ZN(n19194) );
  INV_X1 U17071 ( .A(n19214), .ZN(n19220) );
  NAND2_X1 U17072 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n19341), .ZN(n19320) );
  INV_X1 U17073 ( .A(n19320), .ZN(n19229) );
  NAND2_X1 U17074 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n19229), .ZN(n13727) );
  NAND2_X1 U17075 ( .A1(n19338), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18753) );
  OAI211_X1 U17076 ( .C1(n19194), .C2(n19220), .A(n13727), .B(n18753), .ZN(
        n17103) );
  NOR2_X1 U17077 ( .A1(n18658), .A2(n13728), .ZN(n13787) );
  INV_X1 U17078 ( .A(n19350), .ZN(n13821) );
  NOR2_X1 U17079 ( .A1(n19171), .A2(n13821), .ZN(n13730) );
  INV_X1 U17080 ( .A(n19209), .ZN(n13814) );
  OAI22_X1 U17081 ( .A1(n13814), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n19223), .ZN(n13729) );
  OAI21_X1 U17082 ( .B1(n13730), .B2(n13729), .A(n17103), .ZN(n13731) );
  OAI21_X1 U17083 ( .B1(n17103), .B2(n14105), .A(n13731), .ZN(P3_U3290) );
  NOR2_X1 U17084 ( .A1(n21250), .A2(n13732), .ZN(n13839) );
  AOI21_X1 U17085 ( .B1(n21250), .B2(n13732), .A(n18016), .ZN(n13733) );
  INV_X1 U17086 ( .A(n13733), .ZN(n13748) );
  AOI22_X1 U17087 ( .A1(n17975), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17974), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13737) );
  AOI22_X1 U17088 ( .A1(n17903), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17973), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13736) );
  NAND2_X1 U17089 ( .A1(n17817), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n13735) );
  NAND2_X1 U17090 ( .A1(n17818), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n13734) );
  NAND4_X1 U17091 ( .A1(n13737), .A2(n13736), .A3(n13735), .A4(n13734), .ZN(
        n13740) );
  INV_X1 U17092 ( .A(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13738) );
  OAI22_X1 U17093 ( .A1(n17844), .A2(n13738), .B1(n17981), .B2(n18014), .ZN(
        n13739) );
  OR2_X1 U17094 ( .A1(n13740), .A2(n13739), .ZN(n13747) );
  AOI22_X1 U17095 ( .A1(n17966), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17954), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13745) );
  AOI22_X1 U17096 ( .A1(n9572), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9580), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13744) );
  AOI22_X1 U17097 ( .A1(n11960), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11944), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13743) );
  AOI22_X1 U17098 ( .A1(n9576), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17967), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13742) );
  NAND4_X1 U17099 ( .A1(n13745), .A2(n13744), .A3(n13743), .A4(n13742), .ZN(
        n13746) );
  NOR2_X1 U17100 ( .A1(n13747), .A2(n13746), .ZN(n14011) );
  OAI22_X1 U17101 ( .A1(n13839), .A2(n13748), .B1(n14011), .B2(n18013), .ZN(
        P3_U2694) );
  INV_X1 U17102 ( .A(n17103), .ZN(n13792) );
  NAND2_X1 U17103 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18658), .ZN(
        n13749) );
  NAND2_X1 U17104 ( .A1(n13754), .A2(n13749), .ZN(n13750) );
  NAND2_X1 U17105 ( .A1(n13750), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13757) );
  INV_X1 U17106 ( .A(n13784), .ZN(n13759) );
  AOI21_X1 U17107 ( .B1(n13753), .B2(n13752), .A(n13751), .ZN(n13816) );
  OAI21_X1 U17108 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n13754), .A(
        n13816), .ZN(n13755) );
  NAND2_X1 U17109 ( .A1(n13759), .A2(n13755), .ZN(n13756) );
  MUX2_X1 U17110 ( .A(n13757), .B(n13756), .S(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n13764) );
  NAND2_X1 U17111 ( .A1(n13759), .A2(n13758), .ZN(n13817) );
  NAND2_X1 U17112 ( .A1(n13760), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13819) );
  NAND2_X1 U17113 ( .A1(n13817), .A2(n13819), .ZN(n13766) );
  NOR3_X1 U17114 ( .A1(n13761), .A2(n13760), .A3(n17100), .ZN(n13762) );
  AOI21_X1 U17115 ( .B1(n19179), .B2(n13766), .A(n13762), .ZN(n13763) );
  NAND2_X1 U17116 ( .A1(n13764), .A2(n13763), .ZN(n19166) );
  NOR2_X1 U17117 ( .A1(n19223), .A2(n13980), .ZN(n13789) );
  OAI22_X1 U17118 ( .A1(n18710), .A2(n13765), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13790) );
  INV_X1 U17119 ( .A(n13790), .ZN(n13767) );
  INV_X1 U17120 ( .A(n13766), .ZN(n17704) );
  AOI222_X1 U17121 ( .A1(n19166), .A2(n19350), .B1(n13789), .B2(n13767), .C1(
        n17704), .C2(n19209), .ZN(n13769) );
  NAND2_X1 U17122 ( .A1(n13792), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13768) );
  OAI21_X1 U17123 ( .B1(n13792), .B2(n13769), .A(n13768), .ZN(P3_U3288) );
  NOR2_X1 U17124 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n13771) );
  OAI21_X1 U17125 ( .B1(n13772), .B2(n13771), .A(n13770), .ZN(n13773) );
  NOR2_X1 U17126 ( .A1(n13774), .A2(n20317), .ZN(n13775) );
  NOR2_X1 U17127 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20306), .ZN(
        n19658) );
  AOI211_X1 U17128 ( .C1(n19482), .C2(n20276), .A(n13775), .B(n19658), .ZN(
        n13783) );
  INV_X1 U17129 ( .A(n20319), .ZN(n13776) );
  OAI21_X1 U17130 ( .B1(n20307), .B2(n13777), .A(n13776), .ZN(n13778) );
  OAI21_X1 U17131 ( .B1(n20297), .B2(P2_FLUSH_REG_SCAN_IN), .A(n17244), .ZN(
        n13780) );
  INV_X1 U17132 ( .A(n13780), .ZN(n13781) );
  OR2_X1 U17133 ( .A1(n20133), .A2(n13781), .ZN(n20291) );
  INV_X1 U17134 ( .A(n20291), .ZN(n20294) );
  NAND2_X1 U17135 ( .A1(n20294), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n13782) );
  OAI21_X1 U17136 ( .B1(n13783), .B2(n20294), .A(n13782), .ZN(P2_U3605) );
  NAND2_X1 U17137 ( .A1(n18730), .A2(n14105), .ZN(n13813) );
  INV_X1 U17138 ( .A(n13813), .ZN(n13788) );
  NOR2_X1 U17139 ( .A1(n13785), .A2(n13784), .ZN(n17720) );
  INV_X1 U17140 ( .A(n17720), .ZN(n13786) );
  OAI22_X1 U17141 ( .A1(n13788), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n13787), .B2(n13786), .ZN(n19169) );
  AOI222_X1 U17142 ( .A1(n19169), .A2(n19350), .B1(n13790), .B2(n13789), .C1(
        n19209), .C2(n17720), .ZN(n13793) );
  NAND2_X1 U17143 ( .A1(n13792), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13791) );
  OAI21_X1 U17144 ( .B1(n13793), .B2(n13792), .A(n13791), .ZN(P3_U3289) );
  INV_X1 U17145 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n13796) );
  INV_X2 U17146 ( .A(n20310), .ZN(n19520) );
  AOI22_X1 U17147 ( .A1(n19489), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n19520), 
        .B2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13795) );
  OAI21_X1 U17148 ( .B1(n19492), .B2(n13796), .A(n13795), .ZN(P2_U2927) );
  INV_X1 U17149 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n13798) );
  AOI22_X1 U17150 ( .A1(n19489), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n19520), 
        .B2(P2_UWORD_REG_6__SCAN_IN), .ZN(n13797) );
  OAI21_X1 U17151 ( .B1(n19492), .B2(n13798), .A(n13797), .ZN(P2_U2929) );
  INV_X1 U17152 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n13800) );
  AOI22_X1 U17153 ( .A1(n19489), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n19520), 
        .B2(P2_UWORD_REG_2__SCAN_IN), .ZN(n13799) );
  OAI21_X1 U17154 ( .B1(n19492), .B2(n13800), .A(n13799), .ZN(P2_U2933) );
  INV_X1 U17155 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n13802) );
  AOI22_X1 U17156 ( .A1(n19489), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n19520), 
        .B2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13801) );
  OAI21_X1 U17157 ( .B1(n19492), .B2(n13802), .A(n13801), .ZN(P2_U2925) );
  INV_X1 U17158 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n13804) );
  AOI22_X1 U17159 ( .A1(n19489), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n19520), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n13803) );
  OAI21_X1 U17160 ( .B1(n19492), .B2(n13804), .A(n13803), .ZN(P2_U2935) );
  INV_X1 U17161 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n13806) );
  AOI22_X1 U17162 ( .A1(n19489), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n19520), 
        .B2(P2_UWORD_REG_7__SCAN_IN), .ZN(n13805) );
  OAI21_X1 U17163 ( .B1(n19492), .B2(n13806), .A(n13805), .ZN(P2_U2928) );
  INV_X1 U17164 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n13808) );
  AOI22_X1 U17165 ( .A1(n19489), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n19520), 
        .B2(P2_UWORD_REG_3__SCAN_IN), .ZN(n13807) );
  OAI21_X1 U17166 ( .B1(n19492), .B2(n13808), .A(n13807), .ZN(P2_U2932) );
  INV_X1 U17167 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n13810) );
  AOI22_X1 U17168 ( .A1(n19489), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n19520), 
        .B2(P2_UWORD_REG_5__SCAN_IN), .ZN(n13809) );
  OAI21_X1 U17169 ( .B1(n19492), .B2(n13810), .A(n13809), .ZN(P2_U2930) );
  INV_X1 U17170 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n13812) );
  AOI22_X1 U17171 ( .A1(n19489), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n19520), 
        .B2(P2_UWORD_REG_4__SCAN_IN), .ZN(n13811) );
  OAI21_X1 U17172 ( .B1(n19492), .B2(n13812), .A(n13811), .ZN(P2_U2931) );
  AOI22_X1 U17173 ( .A1(n13813), .A2(n13760), .B1(n19179), .B2(n13817), .ZN(
        n19195) );
  NAND2_X1 U17174 ( .A1(n19350), .A2(n19196), .ZN(n13815) );
  AOI21_X1 U17175 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13819), .A(
        n9578), .ZN(n14281) );
  OAI22_X1 U17176 ( .A1(n19195), .A2(n13815), .B1(n14281), .B2(n13814), .ZN(
        n13823) );
  OAI21_X1 U17177 ( .B1(n13760), .B2(n18730), .A(n13816), .ZN(n13820) );
  INV_X1 U17178 ( .A(n13817), .ZN(n13818) );
  AOI21_X1 U17179 ( .B1(n13820), .B2(n13819), .A(n13818), .ZN(n19193) );
  OAI21_X1 U17180 ( .B1(n19193), .B2(n13821), .A(n17103), .ZN(n13822) );
  AOI22_X1 U17181 ( .A1(n17103), .A2(n13823), .B1(n13822), .B2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13824) );
  INV_X1 U17182 ( .A(n13824), .ZN(P3_U3285) );
  AOI22_X1 U17183 ( .A1(n17948), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17947), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13828) );
  AOI22_X1 U17184 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17818), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13827) );
  AOI22_X1 U17185 ( .A1(n12119), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17973), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13826) );
  AOI22_X1 U17186 ( .A1(n17975), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17974), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13825) );
  NAND4_X1 U17187 ( .A1(n13828), .A2(n13827), .A3(n13826), .A4(n13825), .ZN(
        n13834) );
  AOI22_X1 U17188 ( .A1(n17966), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17954), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13832) );
  AOI22_X1 U17189 ( .A1(n9572), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9581), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13831) );
  AOI22_X1 U17190 ( .A1(n14172), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11944), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13830) );
  AOI22_X1 U17191 ( .A1(n9578), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17967), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13829) );
  NAND4_X1 U17192 ( .A1(n13832), .A2(n13831), .A3(n13830), .A4(n13829), .ZN(
        n13833) );
  OR2_X1 U17193 ( .A1(n13834), .A2(n13833), .ZN(n14207) );
  INV_X1 U17194 ( .A(n14207), .ZN(n13838) );
  NOR2_X1 U17195 ( .A1(n18016), .A2(n14043), .ZN(n17963) );
  OAI21_X1 U17196 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n13836), .A(n17963), .ZN(
        n13837) );
  OAI21_X1 U17197 ( .B1(n13838), .B2(n18013), .A(n13837), .ZN(P3_U2686) );
  NAND2_X1 U17198 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n13839), .ZN(n14073) );
  OAI21_X1 U17199 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n13839), .A(n14073), .ZN(
        n13854) );
  AOI22_X1 U17200 ( .A1(n17966), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17954), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13843) );
  AOI22_X1 U17201 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9583), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13842) );
  AOI22_X1 U17202 ( .A1(n14172), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13841) );
  AOI22_X1 U17203 ( .A1(n9578), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17967), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13840) );
  NAND4_X1 U17204 ( .A1(n13843), .A2(n13842), .A3(n13841), .A4(n13840), .ZN(
        n13852) );
  INV_X1 U17205 ( .A(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17766) );
  AOI22_X1 U17206 ( .A1(n17975), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17974), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13845) );
  NAND2_X1 U17207 ( .A1(n17973), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n13844) );
  OAI211_X1 U17208 ( .C1(n17766), .C2(n10404), .A(n13845), .B(n13844), .ZN(
        n13851) );
  INV_X1 U17209 ( .A(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13846) );
  OAI22_X1 U17210 ( .A1(n12101), .A2(n13847), .B1(n17931), .B2(n13846), .ZN(
        n13850) );
  INV_X1 U17211 ( .A(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13848) );
  OAI22_X1 U17212 ( .A1(n17844), .A2(n13848), .B1(n17981), .B2(n18009), .ZN(
        n13849) );
  OR4_X1 U17213 ( .A1(n13852), .A2(n13851), .A3(n13850), .A4(n13849), .ZN(
        n18097) );
  NAND2_X1 U17214 ( .A1(n18016), .A2(n18097), .ZN(n13853) );
  OAI21_X1 U17215 ( .B1(n13854), .B2(n18016), .A(n13853), .ZN(P3_U2693) );
  AND2_X1 U17216 ( .A1(n13305), .A2(n17135), .ZN(n15579) );
  NAND3_X1 U17217 ( .A1(n14640), .A2(n14550), .A3(n17153), .ZN(n13855) );
  AND2_X1 U17218 ( .A1(n13855), .A2(n21221), .ZN(n21215) );
  OAI21_X1 U17219 ( .B1(n15579), .B2(n13535), .A(n21215), .ZN(n13856) );
  AND2_X1 U17220 ( .A1(n13856), .A2(n14646), .ZN(n13874) );
  NAND2_X1 U17221 ( .A1(n12436), .A2(n12437), .ZN(n13867) );
  NAND2_X1 U17222 ( .A1(n13858), .A2(n20622), .ZN(n14475) );
  AND2_X1 U17223 ( .A1(n14475), .A2(n14486), .ZN(n13859) );
  NAND2_X1 U17224 ( .A1(n13857), .A2(n13859), .ZN(n13875) );
  AOI21_X1 U17225 ( .B1(n13861), .B2(n13860), .A(n14486), .ZN(n13863) );
  INV_X1 U17226 ( .A(n13271), .ZN(n13862) );
  OAI21_X1 U17227 ( .B1(n13863), .B2(n13862), .A(n17135), .ZN(n13866) );
  INV_X1 U17228 ( .A(n13864), .ZN(n13865) );
  NAND4_X1 U17229 ( .A1(n13867), .A2(n13875), .A3(n13866), .A4(n13865), .ZN(
        n14485) );
  INV_X1 U17230 ( .A(n13868), .ZN(n13869) );
  NAND3_X1 U17231 ( .A1(n13539), .A2(n13869), .A3(n12407), .ZN(n13870) );
  NOR2_X1 U17232 ( .A1(n13871), .A2(n12427), .ZN(n13872) );
  INV_X1 U17233 ( .A(n14648), .ZN(n13873) );
  MUX2_X1 U17234 ( .A(n13874), .B(n13873), .S(n17115), .Z(n13880) );
  OAI21_X1 U17235 ( .B1(n13876), .B2(n13305), .A(n13875), .ZN(n14476) );
  OAI21_X1 U17236 ( .B1(n14938), .B2(n12401), .A(n13877), .ZN(n13878) );
  NOR2_X1 U17237 ( .A1(n14476), .A2(n13878), .ZN(n13879) );
  INV_X1 U17238 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20339) );
  NAND2_X1 U17239 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n17185) );
  NAND2_X1 U17240 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n17141), .ZN(n17189) );
  OAI22_X1 U17241 ( .A1(n17117), .A2(n20330), .B1(n20339), .B2(n17189), .ZN(
        n13884) );
  NAND2_X1 U17242 ( .A1(n13884), .A2(n15586), .ZN(n14029) );
  INV_X1 U17243 ( .A(n20724), .ZN(n20961) );
  OR2_X1 U17244 ( .A1(n13881), .A2(n20961), .ZN(n13882) );
  XNOR2_X1 U17245 ( .A(n13882), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n20428) );
  INV_X1 U17246 ( .A(n13539), .ZN(n13883) );
  NAND2_X1 U17247 ( .A1(n20428), .A2(n13883), .ZN(n15559) );
  AOI21_X1 U17248 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n10368), .A(n13884), 
        .ZN(n15593) );
  INV_X1 U17249 ( .A(n15593), .ZN(n14026) );
  OAI22_X1 U17250 ( .A1(n14029), .A2(n15559), .B1(n12693), .B2(n14026), .ZN(
        P1_U3468) );
  XNOR2_X1 U17251 ( .A(n13885), .B(n14188), .ZN(n17025) );
  XOR2_X1 U17252 ( .A(n14187), .B(n13885), .Z(n17022) );
  OR3_X1 U17253 ( .A1(n18616), .A2(n18554), .A3(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18737) );
  AOI21_X1 U17254 ( .B1(n18729), .B2(n18737), .A(n18710), .ZN(n13886) );
  AOI21_X1 U17255 ( .B1(n17022), .B2(n18728), .A(n13886), .ZN(n13891) );
  INV_X1 U17256 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n19251) );
  NAND3_X1 U17257 ( .A1(n14119), .A2(n18710), .A3(n13887), .ZN(n13888) );
  OAI21_X1 U17258 ( .B1(n19251), .B2(n18739), .A(n13888), .ZN(n13889) );
  INV_X1 U17259 ( .A(n13889), .ZN(n13890) );
  OAI211_X1 U17260 ( .C1(n18734), .C2(n17025), .A(n13891), .B(n13890), .ZN(
        P3_U2861) );
  XNOR2_X1 U17261 ( .A(n13893), .B(n13894), .ZN(n16687) );
  NOR2_X1 U17262 ( .A1(n13896), .A2(n13895), .ZN(n13897) );
  AOI21_X1 U17263 ( .B1(n13898), .B2(n16847), .A(n13897), .ZN(n14226) );
  NAND2_X1 U17264 ( .A1(n13900), .A2(n13899), .ZN(n13901) );
  NAND2_X1 U17265 ( .A1(n14226), .A2(n13901), .ZN(n13902) );
  INV_X1 U17266 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19507) );
  INV_X1 U17267 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n13906) );
  OR2_X1 U17268 ( .A1(n19430), .A2(n13906), .ZN(n13908) );
  NAND2_X1 U17269 ( .A1(n19430), .A2(BUF2_REG_7__SCAN_IN), .ZN(n13907) );
  AND2_X1 U17270 ( .A1(n13908), .A2(n13907), .ZN(n19555) );
  OAI222_X1 U17271 ( .A1(n16687), .A2(n19441), .B1(n19445), .B2(n19507), .C1(
        n19485), .C2(n19555), .ZN(P2_U2912) );
  INV_X1 U17272 ( .A(n13909), .ZN(n13911) );
  OR2_X1 U17273 ( .A1(n14551), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13910) );
  AND2_X1 U17274 ( .A1(n13911), .A2(n13910), .ZN(n14972) );
  INV_X1 U17275 ( .A(n14972), .ZN(n20574) );
  NAND2_X1 U17276 ( .A1(n17115), .A2(n14648), .ZN(n13915) );
  INV_X1 U17277 ( .A(n13912), .ZN(n13913) );
  NAND2_X1 U17278 ( .A1(n13913), .A2(n14544), .ZN(n13914) );
  NAND2_X1 U17279 ( .A1(n13915), .A2(n13914), .ZN(n13916) );
  OAI21_X1 U17280 ( .B1(n13919), .B2(n13918), .A(n13917), .ZN(n14975) );
  OAI222_X1 U17281 ( .A1(n20574), .A2(n15013), .B1(n13313), .B2(n20447), .C1(
        n14975), .C2(n15011), .ZN(P1_U2872) );
  OAI21_X1 U17282 ( .B1(n20511), .B2(n13920), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13925) );
  OAI21_X1 U17283 ( .B1(n13922), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13921), .ZN(n20572) );
  INV_X1 U17284 ( .A(n20572), .ZN(n13923) );
  AOI22_X1 U17285 ( .A1(n20519), .A2(n13923), .B1(n20526), .B2(
        P1_REIP_REG_0__SCAN_IN), .ZN(n13924) );
  OAI211_X1 U17286 ( .C1(n14975), .C2(n20583), .A(n13925), .B(n13924), .ZN(
        P1_U2999) );
  INV_X1 U17287 ( .A(n13926), .ZN(n13927) );
  NAND2_X1 U17288 ( .A1(n18102), .A2(n13930), .ZN(n18126) );
  INV_X1 U17289 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n14210) );
  INV_X1 U17290 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n18209) );
  AOI21_X1 U17291 ( .B1(n17863), .B2(n18209), .A(n14009), .ZN(n13932) );
  INV_X1 U17292 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n18211) );
  OR2_X1 U17293 ( .A1(n14009), .A2(n18783), .ZN(n18020) );
  OR2_X1 U17294 ( .A1(n18209), .A2(n18020), .ZN(n13931) );
  OAI22_X1 U17295 ( .A1(n13932), .A2(n18211), .B1(P3_EAX_REG_1__SCAN_IN), .B2(
        n13931), .ZN(n13933) );
  AOI21_X1 U17296 ( .B1(n18104), .B2(n13934), .A(n13933), .ZN(n13935) );
  OAI21_X1 U17297 ( .B1(n18126), .B2(n14210), .A(n13935), .ZN(P3_U2734) );
  NAND2_X1 U17298 ( .A1(n14009), .A2(P3_EAX_REG_0__SCAN_IN), .ZN(n13936) );
  OAI21_X1 U17299 ( .B1(n18020), .B2(P3_EAX_REG_0__SCAN_IN), .A(n13936), .ZN(
        n13937) );
  AOI21_X1 U17300 ( .B1(n18104), .B2(n13938), .A(n13937), .ZN(n13939) );
  OAI21_X1 U17301 ( .B1(n18126), .B2(n18756), .A(n13939), .ZN(P3_U2735) );
  INV_X1 U17302 ( .A(n15857), .ZN(n13941) );
  AOI21_X1 U17303 ( .B1(n13943), .B2(n13942), .A(n13941), .ZN(n16678) );
  INV_X1 U17304 ( .A(n16678), .ZN(n13946) );
  INV_X1 U17305 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19505) );
  INV_X1 U17306 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n14463) );
  OR2_X1 U17307 ( .A1(n19430), .A2(n14463), .ZN(n13945) );
  NAND2_X1 U17308 ( .A1(n19430), .A2(BUF2_REG_8__SCAN_IN), .ZN(n13944) );
  AND2_X1 U17309 ( .A1(n13945), .A2(n13944), .ZN(n19557) );
  OAI222_X1 U17310 ( .A1(n13946), .A2(n19441), .B1(n19445), .B2(n19505), .C1(
        n19485), .C2(n19557), .ZN(P2_U2911) );
  OR2_X1 U17311 ( .A1(n13947), .A2(n14022), .ZN(n13956) );
  INV_X1 U17312 ( .A(n14646), .ZN(n13948) );
  OR2_X1 U17313 ( .A1(n14648), .A2(n13948), .ZN(n13972) );
  XNOR2_X1 U17314 ( .A(n13949), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13957) );
  NAND2_X1 U17315 ( .A1(n14022), .A2(n13950), .ZN(n13963) );
  INV_X1 U17316 ( .A(n13951), .ZN(n13952) );
  OAI211_X1 U17317 ( .C1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n15579), .B(n13952), .ZN(
        n13953) );
  OAI21_X1 U17318 ( .B1(n13963), .B2(n13957), .A(n13953), .ZN(n13954) );
  AOI21_X1 U17319 ( .B1(n13972), .B2(n13957), .A(n13954), .ZN(n13955) );
  NAND2_X1 U17320 ( .A1(n13956), .A2(n13955), .ZN(n15554) );
  INV_X1 U17321 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20555) );
  NOR2_X1 U17322 ( .A1(n13636), .A2(n20555), .ZN(n15589) );
  INV_X1 U17323 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14576) );
  INV_X1 U17324 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20569) );
  OAI22_X1 U17325 ( .A1(n14576), .A2(n20569), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15588) );
  INV_X1 U17326 ( .A(n15588), .ZN(n13959) );
  INV_X1 U17327 ( .A(n13957), .ZN(n13958) );
  AOI222_X1 U17328 ( .A1(n15554), .A2(n15586), .B1(n15589), .B2(n13959), .C1(
        n13958), .C2(n15591), .ZN(n13960) );
  MUX2_X1 U17329 ( .A(n13960), .B(n12649), .S(n15593), .Z(n13961) );
  INV_X1 U17330 ( .A(n13961), .ZN(P1_U3472) );
  INV_X1 U17331 ( .A(n20839), .ZN(n15576) );
  INV_X1 U17332 ( .A(n13963), .ZN(n13966) );
  AOI21_X1 U17333 ( .B1(n13949), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13964) );
  NOR2_X1 U17334 ( .A1(n13016), .A2(n13964), .ZN(n13975) );
  XNOR2_X1 U17335 ( .A(n13951), .B(n12681), .ZN(n13965) );
  AOI22_X1 U17336 ( .A1(n13966), .A2(n13975), .B1(n15579), .B2(n13965), .ZN(
        n13974) );
  INV_X1 U17337 ( .A(n13967), .ZN(n13971) );
  INV_X1 U17338 ( .A(n13968), .ZN(n13969) );
  MUX2_X1 U17339 ( .A(n13969), .B(n12681), .S(n13949), .Z(n13970) );
  NAND3_X1 U17340 ( .A1(n13972), .A2(n13971), .A3(n13970), .ZN(n13973) );
  OAI211_X1 U17341 ( .C1(n15576), .C2(n14022), .A(n13974), .B(n13973), .ZN(
        n15553) );
  AOI22_X1 U17342 ( .A1(n15553), .A2(n15586), .B1(n13975), .B2(n15591), .ZN(
        n13976) );
  MUX2_X1 U17343 ( .A(n13976), .B(n12681), .S(n15593), .Z(n13977) );
  INV_X1 U17344 ( .A(n13977), .ZN(P1_U3469) );
  AOI21_X1 U17345 ( .B1(n14156), .B2(n13979), .A(n13978), .ZN(n18457) );
  INV_X1 U17346 ( .A(n18457), .ZN(n13993) );
  NAND2_X1 U17347 ( .A1(n18658), .A2(n13980), .ZN(n18569) );
  INV_X1 U17348 ( .A(n18569), .ZN(n18715) );
  AOI21_X1 U17349 ( .B1(n19179), .B2(n13981), .A(n18715), .ZN(n13982) );
  OAI21_X1 U17350 ( .B1(n13983), .B2(n18713), .A(n13982), .ZN(n14154) );
  INV_X1 U17351 ( .A(n14154), .ZN(n13984) );
  OAI21_X1 U17352 ( .B1(n13984), .B2(n18616), .A(n18729), .ZN(n18695) );
  XNOR2_X1 U17353 ( .A(n13986), .B(n13985), .ZN(n18453) );
  INV_X1 U17354 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n13987) );
  OAI22_X1 U17355 ( .A1(n18734), .A2(n18453), .B1(n18739), .B2(n13987), .ZN(
        n13988) );
  AOI21_X1 U17356 ( .B1(n18695), .B2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n13988), .ZN(n13992) );
  OAI22_X1 U17357 ( .A1(n18718), .A2(n18712), .B1(n14118), .B2(n18709), .ZN(
        n18700) );
  NAND2_X1 U17358 ( .A1(n13989), .A2(n18700), .ZN(n18565) );
  NOR2_X1 U17359 ( .A1(n18616), .A2(n18565), .ZN(n13990) );
  NAND2_X1 U17360 ( .A1(n13990), .A2(n14156), .ZN(n13991) );
  OAI211_X1 U17361 ( .C1(n13993), .C2(n18629), .A(n13992), .B(n13991), .ZN(
        P3_U2856) );
  MUX2_X1 U17362 ( .A(n13994), .B(n11577), .S(n19429), .Z(n13995) );
  OAI21_X1 U17363 ( .B1(n16820), .B2(n16066), .A(n13995), .ZN(P2_U2887) );
  INV_X1 U17364 ( .A(n13997), .ZN(n14000) );
  INV_X1 U17365 ( .A(n13998), .ZN(n13999) );
  NAND2_X1 U17366 ( .A1(n14000), .A2(n13999), .ZN(n14001) );
  NOR2_X1 U17367 ( .A1(n11572), .A2(n16073), .ZN(n14002) );
  AOI21_X1 U17368 ( .B1(P2_EBX_REG_1__SCAN_IN), .B2(n16073), .A(n14002), .ZN(
        n14003) );
  OAI21_X1 U17369 ( .B1(n20275), .B2(n16066), .A(n14003), .ZN(P2_U2886) );
  MUX2_X1 U17370 ( .A(n15947), .B(n9613), .S(n19429), .Z(n14008) );
  OAI21_X1 U17371 ( .B1(n20288), .B2(n16066), .A(n14008), .ZN(P2_U2885) );
  INV_X1 U17372 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n21365) );
  INV_X1 U17373 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n18220) );
  NAND2_X1 U17374 ( .A1(n18101), .A2(n17863), .ZN(n18108) );
  NOR2_X1 U17375 ( .A1(n18220), .A2(n18108), .ZN(n14010) );
  AOI21_X1 U17376 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n18120), .A(n14010), .ZN(
        n14012) );
  NAND2_X1 U17377 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n14010), .ZN(n18099) );
  OAI222_X1 U17378 ( .A1(n21365), .A2(n18126), .B1(n14012), .B2(n14182), .C1(
        n18123), .C2(n14011), .ZN(P3_U2726) );
  AND2_X1 U17379 ( .A1(n12403), .A2(n12601), .ZN(n14015) );
  INV_X1 U17380 ( .A(n14015), .ZN(n14013) );
  AND2_X1 U17381 ( .A1(n14468), .A2(n14013), .ZN(n14014) );
  INV_X1 U17382 ( .A(DATAI_0_), .ZN(n14018) );
  NAND2_X1 U17383 ( .A1(n20584), .A2(BUF1_REG_0__SCAN_IN), .ZN(n14017) );
  OAI21_X1 U17384 ( .B1(n20584), .B2(n14018), .A(n14017), .ZN(n15077) );
  INV_X1 U17385 ( .A(n15077), .ZN(n20595) );
  INV_X1 U17386 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n21320) );
  OAI222_X1 U17387 ( .A1(n15101), .A2(n14975), .B1(n15100), .B2(n20595), .C1(
        n15098), .C2(n21320), .ZN(P1_U2904) );
  INV_X1 U17388 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18763) );
  AND2_X1 U17389 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n18121), .ZN(n14020) );
  AOI21_X1 U17390 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n18120), .A(n18121), .ZN(
        n14019) );
  OAI222_X1 U17391 ( .A1(n18123), .A2(n14021), .B1(n18126), .B2(n18763), .C1(
        n14020), .C2(n14019), .ZN(P3_U2733) );
  INV_X1 U17392 ( .A(n14022), .ZN(n15585) );
  MUX2_X1 U17393 ( .A(n15579), .B(n14024), .S(n14023), .Z(n14025) );
  AOI21_X1 U17394 ( .B1(n21386), .B2(n15585), .A(n14025), .ZN(n17119) );
  OAI22_X1 U17395 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n15566), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n13636), .ZN(n14027) );
  AOI22_X1 U17396 ( .A1(n15593), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n14027), .B2(n14026), .ZN(n14028) );
  OAI21_X1 U17397 ( .B1(n17119), .B2(n14029), .A(n14028), .ZN(P1_U3474) );
  INV_X1 U17398 ( .A(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14030) );
  OAI22_X1 U17399 ( .A1(n17997), .A2(n12101), .B1(n17931), .B2(n14030), .ZN(
        n14041) );
  AOI22_X1 U17400 ( .A1(n17966), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17954), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14034) );
  AOI22_X1 U17401 ( .A1(n9578), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17967), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14033) );
  AOI22_X1 U17402 ( .A1(n17932), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17953), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14032) );
  AOI22_X1 U17403 ( .A1(n9572), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9580), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14031) );
  NAND4_X1 U17404 ( .A1(n14034), .A2(n14033), .A3(n14032), .A4(n14031), .ZN(
        n14040) );
  INV_X1 U17405 ( .A(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14136) );
  AOI22_X1 U17406 ( .A1(n12119), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17973), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14036) );
  NAND2_X1 U17407 ( .A1(n17974), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n14035) );
  OAI211_X1 U17408 ( .C1(n14136), .C2(n14037), .A(n14036), .B(n14035), .ZN(
        n14039) );
  INV_X1 U17409 ( .A(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17824) );
  INV_X1 U17410 ( .A(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14133) );
  OAI22_X1 U17411 ( .A1(n17824), .A2(n9568), .B1(n17981), .B2(n14133), .ZN(
        n14038) );
  NOR4_X1 U17412 ( .A1(n14041), .A2(n14040), .A3(n14039), .A4(n14038), .ZN(
        n16873) );
  INV_X1 U17413 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n17961) );
  NOR2_X1 U17414 ( .A1(n17510), .A2(n17961), .ZN(n14045) );
  NOR2_X1 U17415 ( .A1(n18783), .A2(n14042), .ZN(n17962) );
  INV_X1 U17416 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n14044) );
  NAND3_X1 U17417 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(P3_EBX_REG_18__SCAN_IN), 
        .A3(n14043), .ZN(n17945) );
  NOR2_X1 U17418 ( .A1(n18016), .A2(n17862), .ZN(n17929) );
  OAI221_X1 U17419 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n14045), .C1(
        P3_EBX_REG_20__SCAN_IN), .C2(n17962), .A(n17929), .ZN(n14046) );
  OAI21_X1 U17420 ( .B1(n16873), .B2(n18013), .A(n14046), .ZN(P3_U2683) );
  NAND2_X1 U17421 ( .A1(n19567), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n14049) );
  INV_X1 U17422 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n17304) );
  OR2_X1 U17423 ( .A1(n19430), .A2(n17304), .ZN(n14048) );
  NAND2_X1 U17424 ( .A1(n19430), .A2(BUF2_REG_9__SCAN_IN), .ZN(n14047) );
  NAND2_X1 U17425 ( .A1(n14048), .A2(n14047), .ZN(n19439) );
  NAND2_X1 U17426 ( .A1(n19538), .A2(n19439), .ZN(n14057) );
  OAI211_X1 U17427 ( .C1(n14050), .C2(n14059), .A(n14049), .B(n14057), .ZN(
        P2_U2961) );
  NAND2_X1 U17428 ( .A1(n19567), .A2(P2_LWORD_REG_11__SCAN_IN), .ZN(n14053) );
  INV_X1 U17429 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n15026) );
  OR2_X1 U17430 ( .A1(n19430), .A2(n15026), .ZN(n14052) );
  NAND2_X1 U17431 ( .A1(n19430), .A2(BUF2_REG_11__SCAN_IN), .ZN(n14051) );
  NAND2_X1 U17432 ( .A1(n14052), .A2(n14051), .ZN(n19435) );
  NAND2_X1 U17433 ( .A1(n19538), .A2(n19435), .ZN(n14054) );
  OAI211_X1 U17434 ( .C1(n19438), .C2(n14059), .A(n14053), .B(n14054), .ZN(
        P2_U2978) );
  NAND2_X1 U17435 ( .A1(n19567), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n14055) );
  OAI211_X1 U17436 ( .C1(n14056), .C2(n14059), .A(n14055), .B(n14054), .ZN(
        P2_U2963) );
  INV_X1 U17437 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19503) );
  NAND2_X1 U17438 ( .A1(n19567), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n14058) );
  OAI211_X1 U17439 ( .C1(n19503), .C2(n14059), .A(n14058), .B(n14057), .ZN(
        P2_U2976) );
  AOI22_X1 U17440 ( .A1(n17975), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17974), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14064) );
  AOI22_X1 U17441 ( .A1(n12119), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17973), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14063) );
  NAND2_X1 U17442 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n14062) );
  NAND2_X1 U17443 ( .A1(n17818), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n14061) );
  NAND4_X1 U17444 ( .A1(n14064), .A2(n14063), .A3(n14062), .A4(n14061), .ZN(
        n14066) );
  INV_X1 U17445 ( .A(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17939) );
  OAI22_X1 U17446 ( .A1(n18002), .A2(n17981), .B1(n9568), .B2(n17939), .ZN(
        n14065) );
  OR2_X1 U17447 ( .A1(n14066), .A2(n14065), .ZN(n14072) );
  AOI22_X1 U17448 ( .A1(n17966), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17954), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14070) );
  AOI22_X1 U17449 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9582), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14069) );
  AOI22_X1 U17450 ( .A1(n14172), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11944), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14068) );
  AOI22_X1 U17451 ( .A1(n9577), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17967), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14067) );
  NAND4_X1 U17452 ( .A1(n14070), .A2(n14069), .A3(n14068), .A4(n14067), .ZN(
        n14071) );
  NOR2_X1 U17453 ( .A1(n14072), .A2(n14071), .ZN(n18093) );
  AOI21_X1 U17454 ( .B1(n17604), .B2(n14073), .A(n18016), .ZN(n14075) );
  NOR2_X1 U17455 ( .A1(n17604), .A2(n14073), .ZN(n14128) );
  INV_X1 U17456 ( .A(n14128), .ZN(n14074) );
  NAND2_X1 U17457 ( .A1(n14075), .A2(n14074), .ZN(n14076) );
  OAI21_X1 U17458 ( .B1(n18093), .B2(n18013), .A(n14076), .ZN(P3_U2692) );
  NAND2_X1 U17459 ( .A1(n15579), .A2(n14077), .ZN(n14078) );
  OAI22_X1 U17460 ( .A1(n14372), .A2(n17135), .B1(n17115), .B2(n14078), .ZN(
        n14079) );
  INV_X1 U17461 ( .A(n17153), .ZN(n14466) );
  NAND2_X1 U17462 ( .A1(n20453), .A2(n14486), .ZN(n14101) );
  NAND2_X1 U17463 ( .A1(n10368), .A2(n17141), .ZN(n20449) );
  INV_X2 U17464 ( .A(n20449), .ZN(n20473) );
  AOI22_X1 U17465 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20473), .B1(n20472), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n14080) );
  OAI21_X1 U17466 ( .B1(n15028), .B2(n14101), .A(n14080), .ZN(P1_U2909) );
  AOI22_X1 U17467 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20473), .B1(n20472), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n14081) );
  OAI21_X1 U17468 ( .B1(n15038), .B2(n14101), .A(n14081), .ZN(P1_U2911) );
  INV_X1 U17469 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n14083) );
  AOI22_X1 U17470 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20473), .B1(n20472), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n14082) );
  OAI21_X1 U17471 ( .B1(n14083), .B2(n14101), .A(n14082), .ZN(P1_U2912) );
  AOI22_X1 U17472 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20473), .B1(n20472), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n14084) );
  OAI21_X1 U17473 ( .B1(n15021), .B2(n14101), .A(n14084), .ZN(P1_U2907) );
  INV_X1 U17474 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n14086) );
  AOI22_X1 U17475 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20473), .B1(n20472), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n14085) );
  OAI21_X1 U17476 ( .B1(n14086), .B2(n14101), .A(n14085), .ZN(P1_U2908) );
  INV_X1 U17477 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n15065) );
  AOI22_X1 U17478 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20473), .B1(n20472), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n14087) );
  OAI21_X1 U17479 ( .B1(n15065), .B2(n14101), .A(n14087), .ZN(P1_U2918) );
  AOI22_X1 U17480 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20473), .B1(n20472), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n14088) );
  OAI21_X1 U17481 ( .B1(n15016), .B2(n14101), .A(n14088), .ZN(P1_U2906) );
  INV_X1 U17482 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n14090) );
  AOI22_X1 U17483 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20473), .B1(n20472), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n14089) );
  OAI21_X1 U17484 ( .B1(n14090), .B2(n14101), .A(n14089), .ZN(P1_U2917) );
  INV_X1 U17485 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n14092) );
  AOI22_X1 U17486 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20473), .B1(n20472), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n14091) );
  OAI21_X1 U17487 ( .B1(n14092), .B2(n14101), .A(n14091), .ZN(P1_U2920) );
  INV_X1 U17488 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n14094) );
  AOI22_X1 U17489 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20473), .B1(n20472), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n14093) );
  OAI21_X1 U17490 ( .B1(n14094), .B2(n14101), .A(n14093), .ZN(P1_U2915) );
  INV_X1 U17491 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n15069) );
  AOI22_X1 U17492 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20473), .B1(n20472), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n14095) );
  OAI21_X1 U17493 ( .B1(n15069), .B2(n14101), .A(n14095), .ZN(P1_U2919) );
  INV_X1 U17494 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14097) );
  AOI22_X1 U17495 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20473), .B1(n20472), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n14096) );
  OAI21_X1 U17496 ( .B1(n14097), .B2(n14101), .A(n14096), .ZN(P1_U2913) );
  INV_X1 U17497 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n21369) );
  AOI22_X1 U17498 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20473), .B1(n20472), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n14098) );
  OAI21_X1 U17499 ( .B1(n21369), .B2(n14101), .A(n14098), .ZN(P1_U2914) );
  INV_X1 U17500 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n15033) );
  AOI22_X1 U17501 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20473), .B1(n20472), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n14099) );
  OAI21_X1 U17502 ( .B1(n15033), .B2(n14101), .A(n14099), .ZN(P1_U2910) );
  AOI22_X1 U17503 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20473), .B1(n20472), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n14100) );
  OAI21_X1 U17504 ( .B1(n14102), .B2(n14101), .A(n14100), .ZN(P1_U2916) );
  INV_X1 U17505 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n14108) );
  AND2_X1 U17506 ( .A1(n19351), .A2(n14103), .ZN(n19353) );
  NOR3_X1 U17507 ( .A1(n17721), .A2(n19350), .A3(n17728), .ZN(n14104) );
  AOI21_X1 U17508 ( .B1(n19353), .B2(n14105), .A(n14104), .ZN(n14107) );
  OAI21_X1 U17509 ( .B1(n17725), .B2(n17724), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n14106) );
  OAI211_X1 U17510 ( .C1(n17673), .C2(n14108), .A(n14107), .B(n14106), .ZN(
        P3_U2671) );
  XNOR2_X2 U17511 ( .A(n14109), .B(n14110), .ZN(n16821) );
  NOR2_X1 U17512 ( .A1(n17207), .A2(n16073), .ZN(n14112) );
  AOI21_X1 U17513 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n16073), .A(n14112), .ZN(
        n14113) );
  OAI21_X1 U17514 ( .B1(n16821), .B2(n16066), .A(n14113), .ZN(P2_U2884) );
  XOR2_X1 U17515 ( .A(n14115), .B(n14114), .Z(n17014) );
  INV_X1 U17516 ( .A(n17014), .ZN(n14127) );
  AND3_X1 U17517 ( .A1(n18700), .A2(n18724), .A3(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14125) );
  OAI211_X1 U17518 ( .C1(n18712), .C2(n14116), .A(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n18569), .ZN(n14117) );
  AOI21_X1 U17519 ( .B1(n14118), .B2(n18576), .A(n14117), .ZN(n18708) );
  INV_X1 U17520 ( .A(n14119), .ZN(n14256) );
  OAI21_X1 U17521 ( .B1(n18708), .B2(n14256), .A(n18729), .ZN(n14124) );
  INV_X1 U17522 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n19255) );
  NOR2_X1 U17523 ( .A1(n14121), .A2(n14120), .ZN(n14122) );
  XOR2_X1 U17524 ( .A(n14122), .B(n18699), .Z(n17016) );
  OAI22_X1 U17525 ( .A1(n18739), .A2(n19255), .B1(n18629), .B2(n17016), .ZN(
        n14123) );
  AOI221_X1 U17526 ( .B1(n14125), .B2(n18699), .C1(n14124), .C2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n14123), .ZN(n14126) );
  OAI21_X1 U17527 ( .B1(n14127), .B2(n18734), .A(n14126), .ZN(P3_U2858) );
  NAND2_X1 U17528 ( .A1(n14128), .A2(n17863), .ZN(n14192) );
  NAND3_X1 U17529 ( .A1(n14192), .A2(P3_EBX_REG_12__SCAN_IN), .A3(n18013), 
        .ZN(n14144) );
  AOI22_X1 U17530 ( .A1(n17975), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17974), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14132) );
  AOI22_X1 U17531 ( .A1(n12119), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17973), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14131) );
  NAND2_X1 U17532 ( .A1(n17817), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n14130) );
  NAND2_X1 U17533 ( .A1(n17818), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n14129) );
  NAND4_X1 U17534 ( .A1(n14132), .A2(n14131), .A3(n14130), .A4(n14129), .ZN(
        n14135) );
  OAI22_X1 U17535 ( .A1(n17997), .A2(n17981), .B1(n9568), .B2(n14133), .ZN(
        n14134) );
  OR2_X1 U17536 ( .A1(n14135), .A2(n14134), .ZN(n14142) );
  AOI22_X1 U17537 ( .A1(n17966), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17954), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14140) );
  AOI22_X1 U17538 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9583), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14139) );
  AOI22_X1 U17539 ( .A1(n14172), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14138) );
  AOI22_X1 U17540 ( .A1(n9578), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17967), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14137) );
  NAND4_X1 U17541 ( .A1(n14140), .A2(n14139), .A3(n14138), .A4(n14137), .ZN(
        n14141) );
  NOR2_X1 U17542 ( .A1(n14142), .A2(n14141), .ZN(n14185) );
  OR2_X1 U17543 ( .A1(n18013), .A2(n14185), .ZN(n14143) );
  OAI211_X1 U17544 ( .C1(n14192), .C2(P3_EBX_REG_12__SCAN_IN), .A(n14144), .B(
        n14143), .ZN(P3_U2691) );
  OR2_X1 U17545 ( .A1(n14146), .A2(n14145), .ZN(n14147) );
  NAND2_X1 U17546 ( .A1(n14302), .A2(n14147), .ZN(n15312) );
  INV_X1 U17547 ( .A(DATAI_1_), .ZN(n14148) );
  INV_X1 U17548 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16182) );
  MUX2_X1 U17549 ( .A(n14148), .B(n16182), .S(n20584), .Z(n20604) );
  INV_X1 U17550 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20471) );
  OAI222_X1 U17551 ( .A1(n15101), .A2(n15312), .B1(n15100), .B2(n20604), .C1(
        n15098), .C2(n20471), .ZN(P1_U2903) );
  XNOR2_X1 U17552 ( .A(n14149), .B(n14550), .ZN(n20556) );
  INV_X1 U17553 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n14150) );
  OAI222_X1 U17554 ( .A1(n20556), .A2(n15013), .B1(n14150), .B2(n20447), .C1(
        n15312), .C2(n15011), .ZN(P1_U2871) );
  NAND2_X1 U17555 ( .A1(n14152), .A2(n14151), .ZN(n14153) );
  INV_X1 U17556 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n14155) );
  XOR2_X1 U17557 ( .A(n14153), .B(n14155), .Z(n17004) );
  INV_X1 U17558 ( .A(n17004), .ZN(n14162) );
  AOI221_X1 U17559 ( .B1(n14156), .B2(n14155), .C1(n18565), .C2(n14155), .A(
        n14257), .ZN(n14160) );
  XNOR2_X1 U17560 ( .A(n14157), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17009) );
  INV_X1 U17561 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n19260) );
  NOR2_X1 U17562 ( .A1(n18739), .A2(n19260), .ZN(n17005) );
  AOI21_X1 U17563 ( .B1(n18701), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n17005), .ZN(n14158) );
  OAI21_X1 U17564 ( .B1(n18734), .B2(n17009), .A(n14158), .ZN(n14159) );
  AOI21_X1 U17565 ( .B1(n14160), .B2(n18724), .A(n14159), .ZN(n14161) );
  OAI21_X1 U17566 ( .B1(n14162), .B2(n18629), .A(n14161), .ZN(P3_U2855) );
  INV_X1 U17567 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n18238) );
  INV_X1 U17568 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n21285) );
  INV_X1 U17569 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n18233) );
  NAND4_X1 U17570 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .A4(P3_EAX_REG_9__SCAN_IN), .ZN(n14163)
         );
  NOR4_X1 U17571 ( .A1(n21285), .A2(n18220), .A3(n18233), .A4(n14163), .ZN(
        n18084) );
  NAND2_X1 U17572 ( .A1(n18101), .A2(n18084), .ZN(n18085) );
  OAI211_X1 U17573 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n14164), .A(n18120), .B(
        n18019), .ZN(n14181) );
  NOR2_X2 U17574 ( .A1(n18775), .A2(n18120), .ZN(n18076) );
  AOI22_X1 U17575 ( .A1(n17975), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17974), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14168) );
  AOI22_X1 U17576 ( .A1(n12119), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17973), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14167) );
  NAND2_X1 U17577 ( .A1(n17817), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n14166) );
  NAND2_X1 U17578 ( .A1(n17818), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n14165) );
  NAND4_X1 U17579 ( .A1(n14168), .A2(n14167), .A3(n14166), .A4(n14165), .ZN(
        n14171) );
  INV_X1 U17580 ( .A(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n21347) );
  OAI22_X1 U17581 ( .A1(n17844), .A2(n21347), .B1(n17981), .B2(n14169), .ZN(
        n14170) );
  OR2_X1 U17582 ( .A1(n14171), .A2(n14170), .ZN(n14178) );
  AOI22_X1 U17583 ( .A1(n17966), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17954), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14176) );
  AOI22_X1 U17584 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9582), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14175) );
  AOI22_X1 U17585 ( .A1(n14172), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14174) );
  AOI22_X1 U17586 ( .A1(n9578), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17967), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14173) );
  NAND4_X1 U17587 ( .A1(n14176), .A2(n14175), .A3(n14174), .A4(n14173), .ZN(
        n14177) );
  NOR2_X1 U17588 ( .A1(n14178), .A2(n14177), .ZN(n14198) );
  NAND2_X1 U17589 ( .A1(n18779), .A2(n18102), .ZN(n18061) );
  INV_X1 U17590 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n16201) );
  OAI22_X1 U17591 ( .A1(n18123), .A2(n14198), .B1(n18061), .B2(n16201), .ZN(
        n14179) );
  AOI21_X1 U17592 ( .B1(n18076), .B2(BUF2_REG_0__SCAN_IN), .A(n14179), .ZN(
        n14180) );
  NAND2_X1 U17593 ( .A1(n14181), .A2(n14180), .ZN(P3_U2719) );
  INV_X1 U17594 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n18227) );
  INV_X1 U17595 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n18151) );
  NAND2_X1 U17596 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n14182), .ZN(n18096) );
  NOR2_X1 U17597 ( .A1(n18151), .A2(n18096), .ZN(n14183) );
  AOI21_X1 U17598 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n18120), .A(n14183), .ZN(
        n14184) );
  OAI222_X1 U17599 ( .A1(n18126), .A2(n18227), .B1(n18123), .B2(n14185), .C1(
        n14236), .C2(n14184), .ZN(P3_U2723) );
  NAND2_X1 U17600 ( .A1(n19178), .A2(n19180), .ZN(n14186) );
  NOR2_X2 U17601 ( .A1(n17362), .A2(n18178), .ZN(n18473) );
  INV_X1 U17602 ( .A(n18473), .ZN(n18488) );
  OR2_X1 U17603 ( .A1(n14188), .A2(n14187), .ZN(n18735) );
  AOI22_X1 U17604 ( .A1(n9600), .A2(n18735), .B1(n18693), .B2(
        P3_REIP_REG_0__SCAN_IN), .ZN(n14191) );
  NAND2_X1 U17605 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18741) );
  NAND2_X1 U17606 ( .A1(n19322), .A2(n18741), .ZN(n19340) );
  NAND2_X1 U17607 ( .A1(n19338), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18313) );
  NAND3_X1 U17608 ( .A1(n19223), .A2(n18495), .A3(n18313), .ZN(n14189) );
  NAND2_X1 U17609 ( .A1(n14189), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14190) );
  OAI211_X1 U17610 ( .C1(n18488), .C2(n18735), .A(n14191), .B(n14190), .ZN(
        P3_U2830) );
  NOR2_X1 U17611 ( .A1(n14193), .A2(n14192), .ZN(n17965) );
  NOR2_X1 U17612 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n14194), .ZN(n14195) );
  AOI22_X1 U17613 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n14196), .B1(n17965), 
        .B2(n14195), .ZN(n14197) );
  OAI21_X1 U17614 ( .B1(n14198), .B2(n18013), .A(n14197), .ZN(P3_U2687) );
  NAND2_X1 U17615 ( .A1(n15859), .A2(n14201), .ZN(n14202) );
  AND2_X1 U17616 ( .A1(n15828), .A2(n14202), .ZN(n16652) );
  INV_X1 U17617 ( .A(n16652), .ZN(n14205) );
  INV_X1 U17618 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n14373) );
  OR2_X1 U17619 ( .A1(n19430), .A2(n14373), .ZN(n14204) );
  NAND2_X1 U17620 ( .A1(n19430), .A2(BUF2_REG_10__SCAN_IN), .ZN(n14203) );
  AND2_X1 U17621 ( .A1(n14204), .A2(n14203), .ZN(n19559) );
  INV_X1 U17622 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n21366) );
  OAI222_X1 U17623 ( .A1(n14205), .A2(n19441), .B1(n19559), .B2(n19485), .C1(
        n21366), .C2(n19445), .ZN(P2_U2909) );
  INV_X1 U17624 ( .A(n18076), .ZN(n18060) );
  NOR2_X1 U17625 ( .A1(n18783), .A2(n18019), .ZN(n14206) );
  NAND2_X1 U17626 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n14206), .ZN(n18078) );
  OAI211_X1 U17627 ( .C1(n14206), .C2(P3_EAX_REG_17__SCAN_IN), .A(n18120), .B(
        n18078), .ZN(n14209) );
  AOI22_X1 U17628 ( .A1(n18104), .A2(n14207), .B1(BUF2_REG_17__SCAN_IN), .B2(
        n18075), .ZN(n14208) );
  OAI211_X1 U17629 ( .C1(n18060), .C2(n14210), .A(n14209), .B(n14208), .ZN(
        P3_U2718) );
  INV_X1 U17630 ( .A(n16821), .ZN(n20280) );
  OR2_X1 U17631 ( .A1(n17207), .A2(n16795), .ZN(n14223) );
  OR2_X1 U17632 ( .A1(n16847), .A2(n16848), .ZN(n16789) );
  NAND2_X1 U17633 ( .A1(n14211), .A2(n16834), .ZN(n16784) );
  AOI22_X1 U17634 ( .A1(n16789), .A2(n16784), .B1(n16785), .B2(n16787), .ZN(
        n14219) );
  INV_X1 U17635 ( .A(n16785), .ZN(n14213) );
  INV_X1 U17636 ( .A(n16784), .ZN(n14212) );
  AOI21_X1 U17637 ( .B1(n16787), .B2(n14213), .A(n14212), .ZN(n14217) );
  NAND2_X1 U17638 ( .A1(n14214), .A2(n9729), .ZN(n16792) );
  NAND2_X1 U17639 ( .A1(n16792), .A2(n9590), .ZN(n14216) );
  AND2_X1 U17640 ( .A1(n14217), .A2(n14216), .ZN(n14218) );
  MUX2_X1 U17641 ( .A(n14219), .B(n14218), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n14221) );
  AND2_X1 U17642 ( .A1(n14221), .A2(n14220), .ZN(n14222) );
  NAND2_X1 U17643 ( .A1(n14223), .A2(n14222), .ZN(n16835) );
  AOI22_X1 U17644 ( .A1(n20280), .A2(n17239), .B1(n20273), .B2(n16835), .ZN(
        n14235) );
  INV_X1 U17645 ( .A(n14224), .ZN(n14225) );
  AND2_X1 U17646 ( .A1(n14226), .A2(n14225), .ZN(n14232) );
  INV_X1 U17647 ( .A(n10857), .ZN(n14227) );
  NAND2_X1 U17648 ( .A1(n14228), .A2(n14227), .ZN(n14230) );
  MUX2_X1 U17649 ( .A(n14230), .B(n14229), .S(n16846), .Z(n14231) );
  INV_X1 U17650 ( .A(n17244), .ZN(n17243) );
  OAI22_X1 U17651 ( .A1(n17243), .A2(n13625), .B1(P2_STATE2_REG_0__SCAN_IN), 
        .B2(n20306), .ZN(n14233) );
  NAND2_X1 U17652 ( .A1(n16802), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14234) );
  OAI21_X1 U17653 ( .B1(n14235), .B2(n16802), .A(n14234), .ZN(P2_U3596) );
  INV_X1 U17654 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n18231) );
  AOI21_X1 U17655 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n18120), .A(n14236), .ZN(
        n14239) );
  NAND2_X1 U17656 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n14236), .ZN(n18092) );
  INV_X1 U17657 ( .A(n18092), .ZN(n14238) );
  OAI222_X1 U17658 ( .A1(n18231), .A2(n18126), .B1(n14239), .B2(n14238), .C1(
        n18123), .C2(n14237), .ZN(P3_U2722) );
  INV_X1 U17659 ( .A(n14240), .ZN(n14242) );
  NAND2_X1 U17660 ( .A1(n14241), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n14340) );
  XNOR2_X1 U17661 ( .A(n14383), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14249) );
  AOI21_X1 U17662 ( .B1(n14246), .B2(n14243), .A(n14245), .ZN(n17194) );
  INV_X1 U17663 ( .A(n17194), .ZN(n16720) );
  MUX2_X1 U17664 ( .A(n14247), .B(n16720), .S(n19429), .Z(n14248) );
  OAI21_X1 U17665 ( .B1(n14249), .B2(n16066), .A(n14248), .ZN(P2_U2882) );
  AOI21_X1 U17666 ( .B1(n14251), .B2(n18678), .A(n14250), .ZN(n14252) );
  INV_X1 U17667 ( .A(n14252), .ZN(n17002) );
  NAND2_X1 U17668 ( .A1(n14253), .A2(n18652), .ZN(n16997) );
  MUX2_X1 U17669 ( .A(n18652), .B(n16997), .S(n18365), .Z(n14254) );
  NAND2_X1 U17670 ( .A1(n14254), .A2(n18437), .ZN(n16999) );
  NAND2_X1 U17671 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n14255) );
  NOR3_X1 U17672 ( .A1(n18616), .A2(n14255), .A3(n18565), .ZN(n14260) );
  OAI21_X1 U17673 ( .B1(n14257), .B2(n14256), .A(n18729), .ZN(n14259) );
  INV_X1 U17674 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n19264) );
  NOR2_X1 U17675 ( .A1(n18739), .A2(n19264), .ZN(n14258) );
  AOI221_X1 U17676 ( .B1(n14260), .B2(n18678), .C1(n14259), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n14258), .ZN(n14261) );
  OAI21_X1 U17677 ( .B1(n18622), .B2(n16997), .A(n14261), .ZN(n14262) );
  AOI21_X1 U17678 ( .B1(n18672), .B2(n16999), .A(n14262), .ZN(n14263) );
  OAI21_X1 U17679 ( .B1(n17002), .B2(n18629), .A(n14263), .ZN(P3_U2854) );
  INV_X1 U17680 ( .A(n14264), .ZN(n14265) );
  NAND2_X1 U17681 ( .A1(n14383), .A2(n14265), .ZN(n14325) );
  NAND2_X1 U17682 ( .A1(n14325), .A2(n19426), .ZN(n14271) );
  AOI21_X1 U17683 ( .B1(n14383), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14270) );
  OAI21_X1 U17684 ( .B1(n14245), .B2(n14267), .A(n14266), .ZN(n16698) );
  MUX2_X1 U17685 ( .A(n16698), .B(n14268), .S(n16073), .Z(n14269) );
  OAI21_X1 U17686 ( .B1(n14271), .B2(n14270), .A(n14269), .ZN(P2_U2881) );
  INV_X1 U17687 ( .A(n19353), .ZN(n14280) );
  INV_X1 U17688 ( .A(n9767), .ZN(n19228) );
  NAND2_X1 U17689 ( .A1(n17728), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17691) );
  INV_X1 U17690 ( .A(n17691), .ZN(n17711) );
  AOI21_X1 U17691 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17711), .A(
        n17695), .ZN(n17710) );
  NOR2_X1 U17692 ( .A1(n17709), .A2(n18496), .ZN(n14273) );
  NAND2_X1 U17693 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n14272), .ZN(
        n17013) );
  OAI21_X1 U17694 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n14273), .A(
        n17013), .ZN(n18483) );
  XNOR2_X1 U17695 ( .A(n17710), .B(n18483), .ZN(n14277) );
  OAI21_X1 U17696 ( .B1(n17729), .B2(n17686), .A(n17644), .ZN(n14274) );
  INV_X1 U17697 ( .A(n14274), .ZN(n17703) );
  AOI221_X1 U17698 ( .B1(n17729), .B2(n21313), .C1(n17716), .C2(n21313), .A(
        n17703), .ZN(n14276) );
  OAI22_X1 U17699 ( .A1(n18477), .A2(n17726), .B1(n17706), .B2(n18000), .ZN(
        n14275) );
  AOI211_X1 U17700 ( .C1(n19228), .C2(n14277), .A(n14276), .B(n14275), .ZN(
        n14279) );
  OAI211_X1 U17701 ( .C1(n17708), .C2(n18000), .A(n17724), .B(n17689), .ZN(
        n14278) );
  OAI211_X1 U17702 ( .C1(n14281), .C2(n14280), .A(n14279), .B(n14278), .ZN(
        P3_U2668) );
  OAI21_X1 U17703 ( .B1(n15827), .B2(n14284), .A(n14283), .ZN(n16631) );
  INV_X1 U17704 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n14513) );
  OR2_X1 U17705 ( .A1(n19430), .A2(n14513), .ZN(n14286) );
  NAND2_X1 U17706 ( .A1(n19430), .A2(BUF2_REG_12__SCAN_IN), .ZN(n14285) );
  AND2_X1 U17707 ( .A1(n14286), .A2(n14285), .ZN(n19561) );
  INV_X1 U17708 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19500) );
  OAI222_X1 U17709 ( .A1(n16631), .A2(n19441), .B1(n19561), .B2(n19485), .C1(
        n19500), .C2(n19445), .ZN(P2_U2907) );
  INV_X1 U17710 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18785) );
  INV_X1 U17711 ( .A(n18108), .ZN(n18083) );
  INV_X1 U17712 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n18159) );
  INV_X1 U17713 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n18163) );
  NAND3_X1 U17714 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(P3_EAX_REG_2__SCAN_IN), 
        .A3(n18121), .ZN(n18116) );
  NOR2_X1 U17715 ( .A1(n18163), .A2(n18116), .ZN(n18119) );
  NAND2_X1 U17716 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n18119), .ZN(n18109) );
  NOR2_X1 U17717 ( .A1(n18159), .A2(n18109), .ZN(n18112) );
  AOI21_X1 U17718 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n18120), .A(n18112), .ZN(
        n14287) );
  OAI222_X1 U17719 ( .A1(n18123), .A2(n16880), .B1(n18126), .B2(n18785), .C1(
        n18083), .C2(n14287), .ZN(P3_U2728) );
  XOR2_X1 U17720 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B(n14325), .Z(n14293)
         );
  NAND2_X1 U17721 ( .A1(n14266), .A2(n14289), .ZN(n14290) );
  NAND2_X1 U17722 ( .A1(n14288), .A2(n14290), .ZN(n16691) );
  INV_X1 U17723 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n14291) );
  MUX2_X1 U17724 ( .A(n16691), .B(n14291), .S(n16073), .Z(n14292) );
  OAI21_X1 U17725 ( .B1(n14293), .B2(n16066), .A(n14292), .ZN(P2_U2880) );
  XNOR2_X1 U17726 ( .A(n14294), .B(n14295), .ZN(n14947) );
  NAND2_X1 U17727 ( .A1(n14296), .A2(n14297), .ZN(n14298) );
  AND2_X1 U17728 ( .A1(n20417), .A2(n14298), .ZN(n20534) );
  AOI22_X1 U17729 ( .A1(n20439), .A2(n20534), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n14996), .ZN(n14299) );
  OAI21_X1 U17730 ( .B1(n14947), .B2(n15011), .A(n14299), .ZN(P1_U2869) );
  INV_X1 U17731 ( .A(n14300), .ZN(n14301) );
  AOI21_X1 U17732 ( .B1(n14303), .B2(n14302), .A(n14301), .ZN(n14956) );
  INV_X1 U17733 ( .A(n14956), .ZN(n14320) );
  OAI21_X1 U17734 ( .B1(n14305), .B2(n14304), .A(n14296), .ZN(n14953) );
  INV_X1 U17735 ( .A(n14953), .ZN(n20541) );
  AOI22_X1 U17736 ( .A1(n20439), .A2(n20541), .B1(P1_EBX_REG_2__SCAN_IN), .B2(
        n14996), .ZN(n14306) );
  OAI21_X1 U17737 ( .B1(n14320), .B2(n15011), .A(n14306), .ZN(P1_U2870) );
  INV_X1 U17738 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n17298) );
  OR2_X1 U17739 ( .A1(n19430), .A2(n17298), .ZN(n14308) );
  NAND2_X1 U17740 ( .A1(n19430), .A2(BUF2_REG_13__SCAN_IN), .ZN(n14307) );
  NAND2_X1 U17741 ( .A1(n14308), .A2(n14307), .ZN(n19535) );
  AOI22_X1 U17742 ( .A1(n19434), .A2(n19535), .B1(P2_EAX_REG_13__SCAN_IN), 
        .B2(n19476), .ZN(n14309) );
  OAI21_X1 U17743 ( .B1(n16616), .B2(n19441), .A(n14309), .ZN(P2_U2906) );
  NAND2_X1 U17744 ( .A1(n20582), .A2(DATAI_3_), .ZN(n14311) );
  NAND2_X1 U17745 ( .A1(n20584), .A2(BUF1_REG_3__SCAN_IN), .ZN(n14310) );
  AND2_X1 U17746 ( .A1(n14311), .A2(n14310), .ZN(n20612) );
  INV_X1 U17747 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20467) );
  OAI222_X1 U17748 ( .A1(n15101), .A2(n14947), .B1(n15100), .B2(n20612), .C1(
        n15098), .C2(n20467), .ZN(P1_U2901) );
  OAI21_X1 U17749 ( .B1(n14314), .B2(n14313), .A(n14312), .ZN(n20542) );
  NAND2_X1 U17750 ( .A1(n14956), .A2(n20518), .ZN(n14317) );
  AND2_X1 U17751 ( .A1(n20577), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n20540) );
  NOR2_X1 U17752 ( .A1(n9869), .A2(n14951), .ZN(n14315) );
  AOI211_X1 U17753 ( .C1(n20511), .C2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n20540), .B(n14315), .ZN(n14316) );
  OAI211_X1 U17754 ( .C1(n20338), .C2(n20542), .A(n14317), .B(n14316), .ZN(
        P1_U2997) );
  NAND2_X1 U17755 ( .A1(n20582), .A2(DATAI_2_), .ZN(n14319) );
  NAND2_X1 U17756 ( .A1(n20584), .A2(BUF1_REG_2__SCAN_IN), .ZN(n14318) );
  AND2_X1 U17757 ( .A1(n14319), .A2(n14318), .ZN(n20608) );
  INV_X1 U17758 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20469) );
  OAI222_X1 U17759 ( .A1(n15101), .A2(n14320), .B1(n15100), .B2(n20608), .C1(
        n15098), .C2(n20469), .ZN(P1_U2902) );
  AND2_X1 U17760 ( .A1(n14288), .A2(n14321), .ZN(n14323) );
  OR2_X1 U17761 ( .A1(n14323), .A2(n14322), .ZN(n16681) );
  NOR2_X1 U17762 ( .A1(n14325), .A2(n14324), .ZN(n14327) );
  NAND2_X1 U17763 ( .A1(n14327), .A2(n14326), .ZN(n16056) );
  OAI211_X1 U17764 ( .C1(n14327), .C2(n14326), .A(n16056), .B(n19426), .ZN(
        n14329) );
  NAND2_X1 U17765 ( .A1(n16073), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n14328) );
  OAI211_X1 U17766 ( .C1(n16681), .C2(n16073), .A(n14329), .B(n14328), .ZN(
        P2_U2879) );
  XNOR2_X1 U17767 ( .A(n16056), .B(n16055), .ZN(n14334) );
  NOR2_X1 U17768 ( .A1(n14322), .A2(n14331), .ZN(n14332) );
  OR2_X1 U17769 ( .A1(n14330), .A2(n14332), .ZN(n16372) );
  MUX2_X1 U17770 ( .A(n16372), .B(n21360), .S(n16073), .Z(n14333) );
  OAI21_X1 U17771 ( .B1(n14334), .B2(n16066), .A(n14333), .ZN(P2_U2878) );
  AND2_X1 U17772 ( .A1(n14336), .A2(n14335), .ZN(n14337) );
  OR2_X1 U17773 ( .A1(n9594), .A2(n14337), .ZN(n20516) );
  INV_X1 U17774 ( .A(DATAI_4_), .ZN(n14339) );
  NAND2_X1 U17775 ( .A1(n20584), .A2(BUF1_REG_4__SCAN_IN), .ZN(n14338) );
  OAI21_X1 U17776 ( .B1(n20584), .B2(n14339), .A(n14338), .ZN(n15058) );
  INV_X1 U17777 ( .A(n15058), .ZN(n20616) );
  INV_X1 U17778 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20465) );
  OAI222_X1 U17779 ( .A1(n15101), .A2(n20516), .B1(n20616), .B2(n15100), .C1(
        n15098), .C2(n20465), .ZN(P1_U2900) );
  NAND2_X1 U17780 ( .A1(n14341), .A2(n14340), .ZN(n14343) );
  INV_X1 U17781 ( .A(n14383), .ZN(n14342) );
  OAI21_X1 U17782 ( .B1(n14344), .B2(n14343), .A(n14342), .ZN(n19411) );
  OR2_X1 U17783 ( .A1(n14346), .A2(n14345), .ZN(n14347) );
  NAND2_X1 U17784 ( .A1(n14348), .A2(n14347), .ZN(n19462) );
  INV_X1 U17785 ( .A(n19462), .ZN(n20286) );
  OR2_X1 U17786 ( .A1(n14350), .A2(n14349), .ZN(n14351) );
  NAND2_X1 U17787 ( .A1(n14352), .A2(n14351), .ZN(n19469) );
  INV_X1 U17788 ( .A(n19469), .ZN(n16759) );
  XNOR2_X1 U17789 ( .A(n19597), .B(n19469), .ZN(n19471) );
  OAI21_X1 U17790 ( .B1(n14355), .B2(n14354), .A(n14353), .ZN(n15966) );
  NOR2_X1 U17791 ( .A1(n16820), .A2(n15966), .ZN(n19478) );
  NOR2_X1 U17792 ( .A1(n19471), .A2(n19478), .ZN(n19470) );
  AOI21_X1 U17793 ( .B1(n16759), .B2(n20275), .A(n19470), .ZN(n19464) );
  XOR2_X1 U17794 ( .A(n19462), .B(n20288), .Z(n19465) );
  NOR2_X1 U17795 ( .A1(n19464), .A2(n19465), .ZN(n19463) );
  AOI21_X1 U17796 ( .B1(n20286), .B2(n20288), .A(n19463), .ZN(n19457) );
  NAND2_X1 U17797 ( .A1(n14358), .A2(n14357), .ZN(n14359) );
  NAND2_X1 U17798 ( .A1(n14356), .A2(n14359), .ZN(n17202) );
  XNOR2_X1 U17799 ( .A(n16821), .B(n17202), .ZN(n19458) );
  NOR2_X1 U17800 ( .A1(n19457), .A2(n19458), .ZN(n19456) );
  INV_X1 U17801 ( .A(n17202), .ZN(n20278) );
  NOR2_X1 U17802 ( .A1(n20280), .A2(n20278), .ZN(n14364) );
  AND2_X1 U17803 ( .A1(n14356), .A2(n14362), .ZN(n14363) );
  OR2_X1 U17804 ( .A1(n14361), .A2(n14363), .ZN(n19408) );
  OAI21_X1 U17805 ( .B1(n19456), .B2(n14364), .A(n19408), .ZN(n19453) );
  XOR2_X1 U17806 ( .A(n19411), .B(n19453), .Z(n14370) );
  INV_X1 U17807 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n14365) );
  OR2_X1 U17808 ( .A1(n19430), .A2(n14365), .ZN(n14367) );
  NAND2_X1 U17809 ( .A1(n19430), .A2(BUF2_REG_4__SCAN_IN), .ZN(n14366) );
  AND2_X1 U17810 ( .A1(n14367), .A2(n14366), .ZN(n19549) );
  INV_X1 U17811 ( .A(n19549), .ZN(n19626) );
  INV_X1 U17812 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19513) );
  OAI22_X1 U17813 ( .A1(n16191), .A2(n19408), .B1(n19445), .B2(n19513), .ZN(
        n14368) );
  AOI21_X1 U17814 ( .B1(n19626), .B2(n19434), .A(n14368), .ZN(n14369) );
  OAI21_X1 U17815 ( .B1(n14370), .B2(n19472), .A(n14369), .ZN(P2_U2915) );
  NOR2_X2 U17816 ( .A1(n20508), .A2(n20603), .ZN(n20493) );
  INV_X1 U17817 ( .A(DATAI_10_), .ZN(n14374) );
  MUX2_X1 U17818 ( .A(n14374), .B(n14373), .S(n20584), .Z(n15094) );
  INV_X1 U17819 ( .A(n15094), .ZN(n14375) );
  NAND2_X1 U17820 ( .A1(n20493), .A2(n14375), .ZN(n20499) );
  AND2_X2 U17821 ( .A1(n14379), .A2(n20603), .ZN(n20505) );
  AOI22_X1 U17822 ( .A1(n20505), .A2(P1_EAX_REG_26__SCAN_IN), .B1(n20508), 
        .B2(P1_UWORD_REG_10__SCAN_IN), .ZN(n14376) );
  NAND2_X1 U17823 ( .A1(n20499), .A2(n14376), .ZN(P1_U2947) );
  INV_X1 U17824 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n15085) );
  INV_X1 U17825 ( .A(n20493), .ZN(n14380) );
  INV_X1 U17826 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n14377) );
  NOR2_X1 U17827 ( .A1(n20582), .A2(n14377), .ZN(n14378) );
  AOI21_X1 U17828 ( .B1(DATAI_15_), .B2(n20582), .A(n14378), .ZN(n15084) );
  INV_X1 U17829 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20450) );
  OAI222_X1 U17830 ( .A1(n14381), .A2(n15085), .B1(n14380), .B2(n15084), .C1(
        n14379), .C2(n20450), .ZN(P1_U2967) );
  NAND2_X1 U17831 ( .A1(n14383), .A2(n14382), .ZN(n16057) );
  XNOR2_X1 U17832 ( .A(n16057), .B(n14424), .ZN(n14386) );
  NOR2_X1 U17833 ( .A1(n19429), .A2(n11172), .ZN(n14384) );
  AOI21_X1 U17834 ( .B1(n16621), .B2(n19429), .A(n14384), .ZN(n14385) );
  OAI21_X1 U17835 ( .B1(n14386), .B2(n16066), .A(n14385), .ZN(P2_U2874) );
  INV_X1 U17836 ( .A(DATAI_6_), .ZN(n14388) );
  NAND2_X1 U17837 ( .A1(n20584), .A2(BUF1_REG_6__SCAN_IN), .ZN(n14387) );
  OAI21_X1 U17838 ( .B1(n20584), .B2(n14388), .A(n14387), .ZN(n15049) );
  NAND2_X1 U17839 ( .A1(n20493), .A2(n15049), .ZN(n14396) );
  AOI22_X1 U17840 ( .A1(n20505), .A2(P1_EAX_REG_6__SCAN_IN), .B1(n20508), .B2(
        P1_LWORD_REG_6__SCAN_IN), .ZN(n14389) );
  NAND2_X1 U17841 ( .A1(n14396), .A2(n14389), .ZN(P1_U2958) );
  NAND2_X1 U17842 ( .A1(n20493), .A2(n15058), .ZN(n14419) );
  AOI22_X1 U17843 ( .A1(n20505), .A2(P1_EAX_REG_20__SCAN_IN), .B1(n20508), 
        .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n14390) );
  NAND2_X1 U17844 ( .A1(n14419), .A2(n14390), .ZN(P1_U2941) );
  INV_X1 U17845 ( .A(n20604), .ZN(n14391) );
  NAND2_X1 U17846 ( .A1(n20493), .A2(n14391), .ZN(n14402) );
  AOI22_X1 U17847 ( .A1(n20505), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n20508), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n14392) );
  NAND2_X1 U17848 ( .A1(n14402), .A2(n14392), .ZN(P1_U2938) );
  INV_X1 U17849 ( .A(n20612), .ZN(n14393) );
  NAND2_X1 U17850 ( .A1(n20493), .A2(n14393), .ZN(n14421) );
  AOI22_X1 U17851 ( .A1(n20505), .A2(P1_EAX_REG_19__SCAN_IN), .B1(n20508), 
        .B2(P1_UWORD_REG_3__SCAN_IN), .ZN(n14394) );
  NAND2_X1 U17852 ( .A1(n14421), .A2(n14394), .ZN(P1_U2940) );
  AOI22_X1 U17853 ( .A1(n20505), .A2(P1_EAX_REG_22__SCAN_IN), .B1(n20508), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n14395) );
  NAND2_X1 U17854 ( .A1(n14396), .A2(n14395), .ZN(P1_U2943) );
  NAND2_X1 U17855 ( .A1(n20582), .A2(DATAI_5_), .ZN(n14398) );
  NAND2_X1 U17856 ( .A1(n20584), .A2(BUF1_REG_5__SCAN_IN), .ZN(n14397) );
  INV_X1 U17857 ( .A(n20619), .ZN(n14399) );
  NAND2_X1 U17858 ( .A1(n20493), .A2(n14399), .ZN(n14415) );
  AOI22_X1 U17859 ( .A1(n20505), .A2(P1_EAX_REG_21__SCAN_IN), .B1(n20508), 
        .B2(P1_UWORD_REG_5__SCAN_IN), .ZN(n14400) );
  NAND2_X1 U17860 ( .A1(n14415), .A2(n14400), .ZN(P1_U2942) );
  AOI22_X1 U17861 ( .A1(n20505), .A2(P1_EAX_REG_1__SCAN_IN), .B1(n20508), .B2(
        P1_LWORD_REG_1__SCAN_IN), .ZN(n14401) );
  NAND2_X1 U17862 ( .A1(n14402), .A2(n14401), .ZN(P1_U2953) );
  NAND2_X1 U17863 ( .A1(n20582), .A2(DATAI_7_), .ZN(n14404) );
  NAND2_X1 U17864 ( .A1(n20584), .A2(BUF1_REG_7__SCAN_IN), .ZN(n14403) );
  INV_X1 U17865 ( .A(n20630), .ZN(n14405) );
  NAND2_X1 U17866 ( .A1(n20493), .A2(n14405), .ZN(n14411) );
  AOI22_X1 U17867 ( .A1(n20505), .A2(P1_EAX_REG_23__SCAN_IN), .B1(n20508), 
        .B2(P1_UWORD_REG_7__SCAN_IN), .ZN(n14406) );
  NAND2_X1 U17868 ( .A1(n14411), .A2(n14406), .ZN(P1_U2944) );
  NAND2_X1 U17869 ( .A1(n20493), .A2(n15077), .ZN(n14409) );
  AOI22_X1 U17870 ( .A1(n20505), .A2(P1_EAX_REG_0__SCAN_IN), .B1(n20508), .B2(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n14407) );
  NAND2_X1 U17871 ( .A1(n14409), .A2(n14407), .ZN(P1_U2952) );
  AOI22_X1 U17872 ( .A1(n20505), .A2(P1_EAX_REG_16__SCAN_IN), .B1(n20508), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n14408) );
  NAND2_X1 U17873 ( .A1(n14409), .A2(n14408), .ZN(P1_U2937) );
  AOI22_X1 U17874 ( .A1(n20505), .A2(P1_EAX_REG_7__SCAN_IN), .B1(n20508), .B2(
        P1_LWORD_REG_7__SCAN_IN), .ZN(n14410) );
  NAND2_X1 U17875 ( .A1(n14411), .A2(n14410), .ZN(P1_U2959) );
  INV_X1 U17876 ( .A(n20608), .ZN(n14412) );
  NAND2_X1 U17877 ( .A1(n20493), .A2(n14412), .ZN(n14417) );
  AOI22_X1 U17878 ( .A1(n20505), .A2(P1_EAX_REG_2__SCAN_IN), .B1(n20508), .B2(
        P1_LWORD_REG_2__SCAN_IN), .ZN(n14413) );
  NAND2_X1 U17879 ( .A1(n14417), .A2(n14413), .ZN(P1_U2954) );
  AOI22_X1 U17880 ( .A1(n20505), .A2(P1_EAX_REG_5__SCAN_IN), .B1(n20508), .B2(
        P1_LWORD_REG_5__SCAN_IN), .ZN(n14414) );
  NAND2_X1 U17881 ( .A1(n14415), .A2(n14414), .ZN(P1_U2957) );
  AOI22_X1 U17882 ( .A1(n20505), .A2(P1_EAX_REG_18__SCAN_IN), .B1(n20508), 
        .B2(P1_UWORD_REG_2__SCAN_IN), .ZN(n14416) );
  NAND2_X1 U17883 ( .A1(n14417), .A2(n14416), .ZN(P1_U2939) );
  AOI22_X1 U17884 ( .A1(n20505), .A2(P1_EAX_REG_4__SCAN_IN), .B1(n20508), .B2(
        P1_LWORD_REG_4__SCAN_IN), .ZN(n14418) );
  NAND2_X1 U17885 ( .A1(n14419), .A2(n14418), .ZN(P1_U2956) );
  AOI22_X1 U17886 ( .A1(n20505), .A2(P1_EAX_REG_3__SCAN_IN), .B1(n20508), .B2(
        P1_LWORD_REG_3__SCAN_IN), .ZN(n14420) );
  NAND2_X1 U17887 ( .A1(n14421), .A2(n14420), .ZN(P1_U2955) );
  OAI21_X1 U17888 ( .B1(n13584), .B2(n14423), .A(n16050), .ZN(n16608) );
  NOR2_X1 U17889 ( .A1(n16057), .A2(n14424), .ZN(n14426) );
  NAND2_X1 U17890 ( .A1(n14426), .A2(n14425), .ZN(n16048) );
  OAI211_X1 U17891 ( .C1(n14426), .C2(n14425), .A(n16048), .B(n19426), .ZN(
        n14428) );
  NAND2_X1 U17892 ( .A1(n16073), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n14427) );
  OAI211_X1 U17893 ( .C1(n16608), .C2(n16073), .A(n14428), .B(n14427), .ZN(
        P2_U2873) );
  XNOR2_X1 U17894 ( .A(n14429), .B(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14432) );
  INV_X1 U17895 ( .A(n14430), .ZN(n14431) );
  NOR2_X1 U17896 ( .A1(n14432), .A2(n14431), .ZN(n20512) );
  AOI21_X1 U17897 ( .B1(n14432), .B2(n14431), .A(n20512), .ZN(n20536) );
  NAND2_X1 U17898 ( .A1(n20536), .A2(n20519), .ZN(n14435) );
  AND2_X1 U17899 ( .A1(n20577), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n20533) );
  NOR2_X1 U17900 ( .A1(n9869), .A2(n14942), .ZN(n14433) );
  AOI211_X1 U17901 ( .C1(n20511), .C2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n20533), .B(n14433), .ZN(n14434) );
  OAI211_X1 U17902 ( .C1(n20583), .C2(n14947), .A(n14435), .B(n14434), .ZN(
        P1_U2996) );
  INV_X1 U17903 ( .A(n14436), .ZN(n14440) );
  INV_X1 U17904 ( .A(n9594), .ZN(n14439) );
  NAND2_X1 U17905 ( .A1(n9594), .A2(n14436), .ZN(n14447) );
  INV_X1 U17906 ( .A(n14447), .ZN(n14438) );
  AOI21_X1 U17907 ( .B1(n14440), .B2(n14439), .A(n14438), .ZN(n20412) );
  INV_X1 U17908 ( .A(n20412), .ZN(n14444) );
  INV_X1 U17909 ( .A(n14442), .ZN(n14452) );
  XNOR2_X1 U17910 ( .A(n14441), .B(n14452), .ZN(n17176) );
  OAI222_X1 U17911 ( .A1(n15011), .A2(n14444), .B1(n14443), .B2(n20447), .C1(
        n15013), .C2(n17176), .ZN(P1_U2867) );
  INV_X1 U17912 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n20463) );
  OAI222_X1 U17913 ( .A1(n15101), .A2(n14444), .B1(n20619), .B2(n15100), .C1(
        n15098), .C2(n20463), .ZN(P1_U2899) );
  INV_X1 U17914 ( .A(n14445), .ZN(n14446) );
  NAND2_X1 U17915 ( .A1(n14447), .A2(n14446), .ZN(n14448) );
  NAND2_X1 U17916 ( .A1(n15008), .A2(n14448), .ZN(n20394) );
  INV_X1 U17917 ( .A(n14450), .ZN(n14451) );
  AOI21_X1 U17918 ( .B1(n14441), .B2(n14452), .A(n14451), .ZN(n14453) );
  OR2_X1 U17919 ( .A1(n14449), .A2(n14453), .ZN(n17168) );
  OAI222_X1 U17920 ( .A1(n20394), .A2(n15011), .B1(n20391), .B2(n20447), .C1(
        n17168), .C2(n15013), .ZN(P1_U2866) );
  INV_X1 U17921 ( .A(n15049), .ZN(n20623) );
  INV_X1 U17922 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n20461) );
  OAI222_X1 U17923 ( .A1(n20394), .A2(n15101), .B1(n20623), .B2(n15100), .C1(
        n20461), .C2(n15098), .ZN(P1_U2898) );
  XNOR2_X1 U17924 ( .A(n14454), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14455) );
  XNOR2_X1 U17925 ( .A(n14456), .B(n14455), .ZN(n17173) );
  NAND2_X1 U17926 ( .A1(n17173), .A2(n20519), .ZN(n14459) );
  NOR2_X1 U17927 ( .A1(n15267), .A2(n21160), .ZN(n17169) );
  NOR2_X1 U17928 ( .A1(n9869), .A2(n20402), .ZN(n14457) );
  AOI211_X1 U17929 ( .C1(n20511), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n17169), .B(n14457), .ZN(n14458) );
  OAI211_X1 U17930 ( .C1(n20583), .C2(n20394), .A(n14459), .B(n14458), .ZN(
        P1_U2993) );
  INV_X1 U17931 ( .A(n14460), .ZN(n15007) );
  NOR2_X1 U17932 ( .A1(n15008), .A2(n15007), .ZN(n15010) );
  OAI21_X1 U17933 ( .B1(n15010), .B2(n14462), .A(n14461), .ZN(n15308) );
  INV_X1 U17934 ( .A(DATAI_8_), .ZN(n14464) );
  MUX2_X1 U17935 ( .A(n14464), .B(n14463), .S(n20584), .Z(n20476) );
  INV_X1 U17936 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n14465) );
  OAI222_X1 U17937 ( .A1(n15308), .A2(n15101), .B1(n20476), .B2(n15100), .C1(
        n14465), .C2(n15098), .ZN(P1_U2896) );
  OAI22_X1 U17938 ( .A1(n14467), .A2(n12427), .B1(n14466), .B2(n21216), .ZN(
        n14469) );
  AND2_X1 U17939 ( .A1(n14469), .A2(n14468), .ZN(n14470) );
  NAND2_X1 U17940 ( .A1(n17135), .A2(n17153), .ZN(n14473) );
  INV_X1 U17941 ( .A(n14471), .ZN(n14472) );
  NAND2_X1 U17942 ( .A1(n14473), .A2(n14472), .ZN(n14474) );
  INV_X1 U17943 ( .A(n14475), .ZN(n14477) );
  AOI21_X1 U17944 ( .B1(n17115), .B2(n14477), .A(n14476), .ZN(n14478) );
  OR2_X1 U17945 ( .A1(n14500), .A2(n20615), .ZN(n14481) );
  NAND4_X1 U17946 ( .A1(n14480), .A2(n14645), .A3(n14646), .A4(n14481), .ZN(
        n14482) );
  XNOR2_X1 U17947 ( .A(n14484), .B(n14483), .ZN(n17157) );
  INV_X1 U17948 ( .A(n14485), .ZN(n14490) );
  MUX2_X1 U17949 ( .A(n14487), .B(n20607), .S(n14486), .Z(n14488) );
  NAND3_X1 U17950 ( .A1(n14490), .A2(n14489), .A3(n14488), .ZN(n14491) );
  NAND2_X1 U17951 ( .A1(n14502), .A2(n15579), .ZN(n20579) );
  AND2_X2 U17952 ( .A1(n20545), .A2(n15515), .ZN(n20562) );
  INV_X1 U17953 ( .A(n20579), .ZN(n14492) );
  NOR2_X1 U17954 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n14492), .ZN(
        n20561) );
  NOR2_X1 U17955 ( .A1(n14494), .A2(n14493), .ZN(n20523) );
  NAND2_X1 U17956 ( .A1(n14495), .A2(n20523), .ZN(n17181) );
  INV_X1 U17957 ( .A(n17181), .ZN(n14499) );
  NOR2_X1 U17958 ( .A1(n20548), .A2(n20569), .ZN(n15513) );
  NAND2_X1 U17959 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n20523), .ZN(
        n14505) );
  INV_X1 U17960 ( .A(n14505), .ZN(n14557) );
  OAI21_X1 U17961 ( .B1(n20555), .B2(n20569), .A(n20548), .ZN(n15514) );
  NAND2_X1 U17962 ( .A1(n14557), .A2(n15514), .ZN(n15520) );
  NAND2_X1 U17963 ( .A1(n20571), .A2(n20555), .ZN(n14498) );
  INV_X1 U17964 ( .A(n14502), .ZN(n14496) );
  NAND2_X1 U17965 ( .A1(n14496), .A2(n15267), .ZN(n14497) );
  NAND2_X1 U17966 ( .A1(n14498), .A2(n14497), .ZN(n20554) );
  AOI21_X1 U17967 ( .B1(n20570), .B2(n15520), .A(n20554), .ZN(n15491) );
  OAI221_X1 U17968 ( .B1(n20545), .B2(n15513), .C1(n20545), .C2(n20523), .A(
        n15491), .ZN(n17178) );
  AOI21_X1 U17969 ( .B1(n20549), .B2(n14499), .A(n17178), .ZN(n17175) );
  OAI21_X1 U17970 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n20562), .A(
        n17175), .ZN(n15545) );
  OAI22_X1 U17971 ( .A1(n13298), .A2(n17135), .B1(n12406), .B2(n14500), .ZN(
        n14501) );
  OAI21_X1 U17972 ( .B1(n14449), .B2(n14504), .A(n15539), .ZN(n20379) );
  AOI22_X1 U17973 ( .A1(n20570), .A2(n15514), .B1(n20549), .B2(n15513), .ZN(
        n20539) );
  NOR2_X1 U17974 ( .A1(n20539), .A2(n14505), .ZN(n15541) );
  NAND3_X1 U17975 ( .A1(n15541), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        n14506), .ZN(n14507) );
  NAND2_X1 U17976 ( .A1(n20526), .A2(P1_REIP_REG_7__SCAN_IN), .ZN(n17159) );
  OAI211_X1 U17977 ( .C1(n20575), .C2(n20379), .A(n14507), .B(n17159), .ZN(
        n14508) );
  AOI21_X1 U17978 ( .B1(n15545), .B2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n14508), .ZN(n14509) );
  OAI21_X1 U17979 ( .B1(n20573), .B2(n17157), .A(n14509), .ZN(P1_U3024) );
  NOR3_X1 U17980 ( .A1(n18783), .A2(n17992), .A3(n17995), .ZN(n17989) );
  AOI21_X1 U17981 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17989), .A(
        P3_EBX_REG_7__SCAN_IN), .ZN(n14510) );
  NOR2_X1 U17982 ( .A1(n14511), .A2(n14510), .ZN(n14512) );
  MUX2_X1 U17983 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B(n14512), .S(n18013), 
        .Z(P3_U2696) );
  INV_X1 U17984 ( .A(DATAI_12_), .ZN(n14514) );
  MUX2_X1 U17985 ( .A(n14514), .B(n14513), .S(n20584), .Z(n20485) );
  OAI22_X1 U17986 ( .A1(n15070), .A2(n20485), .B1(n15098), .B2(n14086), .ZN(
        n14515) );
  AOI21_X1 U17987 ( .B1(BUF1_REG_28__SCAN_IN), .B2(n15072), .A(n14515), .ZN(
        n14517) );
  NAND2_X1 U17988 ( .A1(n15082), .A2(DATAI_28_), .ZN(n14516) );
  OAI211_X1 U17989 ( .C1(n14532), .C2(n15101), .A(n14517), .B(n14516), .ZN(
        P1_U2876) );
  INV_X1 U17990 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14521) );
  NAND2_X1 U17991 ( .A1(n14518), .A2(n14519), .ZN(n14520) );
  NAND2_X1 U17992 ( .A1(n9657), .A2(n14520), .ZN(n14522) );
  OAI222_X1 U17993 ( .A1(n15011), .A2(n14532), .B1(n14521), .B2(n20447), .C1(
        n14522), .C2(n15013), .ZN(P1_U2844) );
  INV_X1 U17994 ( .A(n14522), .ZN(n15338) );
  INV_X1 U17995 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n14529) );
  INV_X1 U17996 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n15123) );
  NOR3_X1 U17997 ( .A1(n14682), .A2(P1_REIP_REG_28__SCAN_IN), .A3(n15123), 
        .ZN(n14527) );
  INV_X1 U17998 ( .A(n14523), .ZN(n14525) );
  OAI22_X1 U17999 ( .A1(n14969), .A2(n14525), .B1(n14524), .B2(n20407), .ZN(
        n14526) );
  AOI211_X1 U18000 ( .C1(P1_EBX_REG_28__SCAN_IN), .C2(n20405), .A(n14527), .B(
        n14526), .ZN(n14528) );
  OAI21_X1 U18001 ( .B1(n14589), .B2(n14529), .A(n14528), .ZN(n14530) );
  AOI21_X1 U18002 ( .B1(n15338), .B2(n20404), .A(n14530), .ZN(n14531) );
  OAI21_X1 U18003 ( .B1(n14532), .B2(n20393), .A(n14531), .ZN(P1_U2812) );
  INV_X1 U18004 ( .A(n14537), .ZN(n14535) );
  INV_X1 U18005 ( .A(n14533), .ZN(n14534) );
  NAND2_X1 U18006 ( .A1(n14538), .A2(n9569), .ZN(n15139) );
  NAND2_X1 U18007 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15325) );
  NAND2_X1 U18008 ( .A1(n9569), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15113) );
  INV_X1 U18009 ( .A(n15113), .ZN(n14540) );
  NAND2_X1 U18010 ( .A1(n15102), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14542) );
  NOR2_X1 U18011 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15335) );
  INV_X1 U18012 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15328) );
  NAND2_X1 U18013 ( .A1(n10374), .A2(n15328), .ZN(n15114) );
  NOR2_X1 U18014 ( .A1(n15114), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14541) );
  INV_X1 U18015 ( .A(n14551), .ZN(n14545) );
  INV_X1 U18016 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14976) );
  INV_X1 U18017 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14543) );
  OAI22_X1 U18018 ( .A1(n14545), .A2(n14976), .B1(n14544), .B2(n14543), .ZN(
        n14660) );
  NAND2_X1 U18019 ( .A1(n14546), .A2(n14660), .ZN(n14548) );
  OAI21_X1 U18020 ( .B1(n9657), .B2(n14659), .A(n14658), .ZN(n14547) );
  OAI21_X1 U18021 ( .B1(n14548), .B2(n9657), .A(n14547), .ZN(n14549) );
  AOI22_X1 U18022 ( .A1(n14551), .A2(P1_EBX_REG_31__SCAN_IN), .B1(n14550), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14552) );
  INV_X1 U18023 ( .A(n20562), .ZN(n15519) );
  NOR2_X1 U18024 ( .A1(n15519), .A2(n20554), .ZN(n14566) );
  INV_X1 U18025 ( .A(n14566), .ZN(n14567) );
  NAND2_X1 U18026 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15506) );
  NAND2_X1 U18027 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15543) );
  INV_X1 U18028 ( .A(n15543), .ZN(n14555) );
  NAND2_X1 U18029 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n14555), .ZN(
        n15521) );
  NOR2_X1 U18030 ( .A1(n15506), .A2(n15521), .ZN(n15488) );
  AND2_X1 U18031 ( .A1(n15488), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15495) );
  NAND2_X1 U18032 ( .A1(n15495), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15470) );
  NOR2_X1 U18033 ( .A1(n15470), .A2(n15520), .ZN(n15403) );
  AND2_X1 U18034 ( .A1(n15435), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14570) );
  AND2_X1 U18035 ( .A1(n14556), .A2(n14570), .ZN(n14558) );
  AND2_X1 U18036 ( .A1(n15403), .A2(n14558), .ZN(n15406) );
  NAND2_X1 U18037 ( .A1(n20545), .A2(n15406), .ZN(n14559) );
  NAND2_X1 U18038 ( .A1(n15513), .A2(n14557), .ZN(n15490) );
  NOR2_X1 U18039 ( .A1(n15470), .A2(n15490), .ZN(n14568) );
  NAND2_X1 U18040 ( .A1(n14568), .A2(n14558), .ZN(n15404) );
  AOI21_X1 U18041 ( .B1(n14559), .B2(n15404), .A(n14571), .ZN(n14560) );
  OR2_X1 U18042 ( .A1(n14560), .A2(n20562), .ZN(n14561) );
  INV_X1 U18043 ( .A(n20554), .ZN(n20544) );
  NAND2_X1 U18044 ( .A1(n14561), .A2(n20544), .ZN(n15393) );
  AND2_X1 U18045 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14572) );
  NOR2_X1 U18046 ( .A1(n20562), .A2(n14572), .ZN(n14562) );
  OR2_X1 U18047 ( .A1(n15393), .A2(n14562), .ZN(n15378) );
  INV_X1 U18048 ( .A(n14563), .ZN(n14564) );
  NOR2_X1 U18049 ( .A1(n20562), .A2(n14564), .ZN(n15359) );
  NOR3_X1 U18050 ( .A1(n15378), .A2(n15359), .A3(n14565), .ZN(n15354) );
  NOR2_X1 U18051 ( .A1(n15354), .A2(n14566), .ZN(n15345) );
  AOI21_X1 U18052 ( .B1(n15325), .B2(n14567), .A(n15345), .ZN(n15329) );
  OAI211_X1 U18053 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n20562), .A(
        n15329), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15319) );
  NAND3_X1 U18054 ( .A1(n15319), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14567), .ZN(n14578) );
  NAND2_X1 U18055 ( .A1(n20526), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n14582) );
  AND2_X1 U18056 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15403), .ZN(
        n15427) );
  NAND2_X1 U18057 ( .A1(n20570), .A2(n15427), .ZN(n14569) );
  INV_X1 U18058 ( .A(n14568), .ZN(n15478) );
  NOR2_X1 U18059 ( .A1(n15482), .A2(n15478), .ZN(n15426) );
  INV_X1 U18060 ( .A(n14572), .ZN(n14573) );
  NAND2_X1 U18061 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14575) );
  NAND3_X1 U18062 ( .A1(n14578), .A2(n14582), .A3(n14577), .ZN(n14579) );
  AOI21_X1 U18063 ( .B1(n14587), .B2(n20560), .A(n14579), .ZN(n14580) );
  OAI21_X1 U18064 ( .B1(n14586), .B2(n20573), .A(n14580), .ZN(P1_U3000) );
  NAND2_X1 U18065 ( .A1(n20511), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14581) );
  OAI211_X1 U18066 ( .C1(n14583), .C2(n9869), .A(n14582), .B(n14581), .ZN(
        n14584) );
  OAI21_X1 U18067 ( .B1(n14586), .B2(n20338), .A(n14585), .ZN(P1_U2968) );
  INV_X1 U18068 ( .A(n14587), .ZN(n14598) );
  INV_X1 U18069 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14592) );
  OAI22_X1 U18070 ( .A1(n14598), .A2(n15013), .B1(n20447), .B2(n14592), .ZN(
        P1_U2841) );
  NAND2_X1 U18071 ( .A1(n14588), .A2(n20383), .ZN(n14597) );
  INV_X1 U18072 ( .A(n14835), .ZN(n14967) );
  NAND2_X1 U18073 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(P1_REIP_REG_29__SCAN_IN), 
        .ZN(n14593) );
  INV_X1 U18074 ( .A(n14593), .ZN(n14590) );
  OAI21_X1 U18075 ( .B1(n14967), .B2(n14590), .A(n14589), .ZN(n14672) );
  INV_X1 U18076 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14591) );
  OAI22_X1 U18077 ( .A1(n20424), .A2(n14592), .B1(n14591), .B2(n20407), .ZN(
        n14595) );
  NOR3_X1 U18078 ( .A1(n14667), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14593), 
        .ZN(n14594) );
  AOI211_X1 U18079 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n14672), .A(n14595), 
        .B(n14594), .ZN(n14596) );
  OAI211_X1 U18080 ( .C1(n14598), .C2(n20432), .A(n14597), .B(n14596), .ZN(
        P1_U2809) );
  NAND2_X1 U18081 ( .A1(n16073), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n14599) );
  OAI21_X1 U18082 ( .B1(n14600), .B2(n16073), .A(n14599), .ZN(P2_U2856) );
  INV_X1 U18083 ( .A(n14601), .ZN(n14611) );
  OAI21_X1 U18084 ( .B1(n14603), .B2(n14602), .A(n15942), .ZN(n14606) );
  INV_X1 U18085 ( .A(n14604), .ZN(n14605) );
  AOI22_X1 U18086 ( .A1(n19403), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19410), .ZN(n14608) );
  OAI21_X1 U18087 ( .B1(n10111), .B2(n19389), .A(n14608), .ZN(n14609) );
  INV_X1 U18088 ( .A(n14609), .ZN(n14610) );
  AOI21_X1 U18089 ( .B1(n16518), .B2(n16749), .A(n17216), .ZN(n14613) );
  OAI21_X1 U18090 ( .B1(n16515), .B2(n16749), .A(n14613), .ZN(n14624) );
  XOR2_X1 U18091 ( .A(n14615), .B(n14614), .Z(n14632) );
  AOI221_X1 U18092 ( .B1(n14616), .B2(n16562), .C1(n16749), .C2(n16515), .A(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14617) );
  INV_X1 U18093 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n20211) );
  NOR2_X1 U18094 ( .A1(n17200), .A2(n20211), .ZN(n14626) );
  AOI211_X1 U18095 ( .C1(n17209), .C2(n14632), .A(n14617), .B(n14626), .ZN(
        n14622) );
  INV_X1 U18096 ( .A(n14618), .ZN(n14627) );
  NAND2_X1 U18097 ( .A1(n14620), .A2(n14619), .ZN(n14628) );
  NAND3_X1 U18098 ( .A1(n17224), .A2(n14627), .A3(n14628), .ZN(n14621) );
  OAI211_X1 U18099 ( .C1(n20286), .C2(n17203), .A(n14622), .B(n14621), .ZN(
        n14623) );
  AOI21_X1 U18100 ( .B1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n14624), .A(
        n14623), .ZN(n14625) );
  OAI21_X1 U18101 ( .B1(n9613), .B2(n17227), .A(n14625), .ZN(P2_U3044) );
  AOI21_X1 U18102 ( .B1(n19584), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n14626), .ZN(n14630) );
  NAND3_X1 U18103 ( .A1(n14628), .A2(n19586), .A3(n14627), .ZN(n14629) );
  OAI211_X1 U18104 ( .C1(n19582), .C2(n15941), .A(n14630), .B(n14629), .ZN(
        n14631) );
  AOI21_X1 U18105 ( .B1(n14632), .B2(n19577), .A(n14631), .ZN(n14633) );
  OAI21_X1 U18106 ( .B1(n9613), .B2(n19573), .A(n14633), .ZN(P2_U3012) );
  AOI22_X1 U18107 ( .A1(n16193), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n19476), .ZN(n14639) );
  INV_X1 U18108 ( .A(n14635), .ZN(n14636) );
  INV_X1 U18109 ( .A(n16200), .ZN(n14637) );
  NAND2_X1 U18110 ( .A1(n14637), .A2(BUF2_REG_31__SCAN_IN), .ZN(n14638) );
  OAI211_X1 U18111 ( .C1(n14634), .C2(n16191), .A(n14639), .B(n14638), .ZN(
        P2_U2888) );
  OR2_X1 U18112 ( .A1(n14790), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n14643) );
  NAND2_X1 U18113 ( .A1(n14641), .A2(n14640), .ZN(n14642) );
  MUX2_X1 U18114 ( .A(n14643), .B(n14642), .S(n21219), .Z(P1_U3487) );
  NAND3_X1 U18115 ( .A1(n14646), .A2(n14645), .A3(n14644), .ZN(n14647) );
  MUX2_X1 U18116 ( .A(n14648), .B(n14647), .S(n17115), .Z(n14652) );
  INV_X1 U18117 ( .A(n13305), .ZN(n14649) );
  NOR2_X1 U18118 ( .A1(n14650), .A2(n14649), .ZN(n14651) );
  OR2_X1 U18119 ( .A1(n14652), .A2(n14651), .ZN(n14653) );
  NAND2_X1 U18120 ( .A1(n14653), .A2(n12408), .ZN(n17127) );
  INV_X1 U18121 ( .A(n17127), .ZN(n14657) );
  INV_X1 U18122 ( .A(n17115), .ZN(n14656) );
  INV_X1 U18123 ( .A(n13298), .ZN(n14655) );
  OAI22_X1 U18124 ( .A1(n14656), .A2(n12437), .B1(n14655), .B2(n14654), .ZN(
        n20331) );
  NOR2_X1 U18125 ( .A1(n20331), .A2(n21215), .ZN(n17131) );
  NOR2_X1 U18126 ( .A1(n17131), .A2(n20330), .ZN(n20340) );
  MUX2_X1 U18127 ( .A(P1_MORE_REG_SCAN_IN), .B(n14657), .S(n20340), .Z(
        P1_U3484) );
  INV_X1 U18128 ( .A(n9595), .ZN(n15111) );
  NAND2_X1 U18129 ( .A1(n15111), .A2(n20383), .ZN(n14674) );
  INV_X1 U18130 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n14666) );
  INV_X1 U18131 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14665) );
  OAI21_X1 U18132 ( .B1(n14667), .B2(n14666), .A(n14665), .ZN(n14671) );
  NOR2_X1 U18133 ( .A1(n20424), .A2(n14976), .ZN(n14670) );
  INV_X1 U18134 ( .A(n15107), .ZN(n14668) );
  OAI22_X1 U18135 ( .A1(n9611), .A2(n14668), .B1(n15109), .B2(n20407), .ZN(
        n14669) );
  AOI211_X1 U18136 ( .C1(n14672), .C2(n14671), .A(n14670), .B(n14669), .ZN(
        n14673) );
  OAI211_X1 U18137 ( .C1(n20432), .C2(n15323), .A(n14674), .B(n14673), .ZN(
        P1_U2810) );
  AOI21_X1 U18138 ( .B1(n14677), .B2(n14676), .A(n13126), .ZN(n15127) );
  INV_X1 U18139 ( .A(n15127), .ZN(n15032) );
  AND2_X1 U18140 ( .A1(n14835), .A2(n14678), .ZN(n14698) );
  OAI22_X1 U18141 ( .A1(n9611), .A2(n15125), .B1(n14679), .B2(n20407), .ZN(
        n14680) );
  AOI21_X1 U18142 ( .B1(n20405), .B2(P1_EBX_REG_27__SCAN_IN), .A(n14680), .ZN(
        n14681) );
  OAI21_X1 U18143 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(n14682), .A(n14681), 
        .ZN(n14687) );
  OR2_X1 U18144 ( .A1(n14683), .A2(n14684), .ZN(n14685) );
  NAND2_X1 U18145 ( .A1(n14518), .A2(n14685), .ZN(n15346) );
  NOR2_X1 U18146 ( .A1(n15346), .A2(n20432), .ZN(n14686) );
  AOI211_X1 U18147 ( .C1(P1_REIP_REG_27__SCAN_IN), .C2(n14698), .A(n14687), 
        .B(n14686), .ZN(n14688) );
  OAI21_X1 U18148 ( .B1(n15032), .B2(n20393), .A(n14688), .ZN(P1_U2813) );
  OAI21_X1 U18149 ( .B1(n14689), .B2(n14690), .A(n14676), .ZN(n15132) );
  INV_X1 U18150 ( .A(n14683), .ZN(n14693) );
  NAND2_X1 U18151 ( .A1(n14710), .A2(n14691), .ZN(n14692) );
  NAND2_X1 U18152 ( .A1(n14693), .A2(n14692), .ZN(n14980) );
  INV_X1 U18153 ( .A(n14980), .ZN(n15356) );
  OR2_X1 U18154 ( .A1(n14969), .A2(n15134), .ZN(n14702) );
  INV_X1 U18155 ( .A(n14694), .ZN(n14713) );
  NAND3_X1 U18156 ( .A1(n14713), .A2(P1_REIP_REG_25__SCAN_IN), .A3(n14695), 
        .ZN(n14696) );
  OAI22_X1 U18157 ( .A1(n20420), .A2(n14696), .B1(n20424), .B2(n14981), .ZN(
        n14697) );
  INV_X1 U18158 ( .A(n14697), .ZN(n14701) );
  NAND2_X1 U18159 ( .A1(n14698), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14700) );
  NAND2_X1 U18160 ( .A1(n20427), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14699) );
  NAND4_X1 U18161 ( .A1(n14702), .A2(n14701), .A3(n14700), .A4(n14699), .ZN(
        n14703) );
  AOI21_X1 U18162 ( .B1(n15356), .B2(n20404), .A(n14703), .ZN(n14704) );
  OAI21_X1 U18163 ( .B1(n15132), .B2(n20393), .A(n14704), .ZN(P1_U2814) );
  NAND2_X1 U18164 ( .A1(n14725), .A2(n14708), .ZN(n14709) );
  AND2_X1 U18165 ( .A1(n14710), .A2(n14709), .ZN(n15364) );
  INV_X1 U18166 ( .A(n14726), .ZN(n14711) );
  NAND2_X1 U18167 ( .A1(n20410), .A2(n14711), .ZN(n14712) );
  NAND2_X1 U18168 ( .A1(n14835), .A2(n14712), .ZN(n14739) );
  NOR2_X1 U18169 ( .A1(n14713), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14714) );
  AOI211_X1 U18170 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(P1_REIP_REG_24__SCAN_IN), .A(n14714), .B(n20420), .ZN(n14715) );
  AOI21_X1 U18171 ( .B1(P1_EBX_REG_25__SCAN_IN), .B2(n20405), .A(n14715), .ZN(
        n14717) );
  AOI22_X1 U18172 ( .A1(n10405), .A2(n15147), .B1(
        P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n20427), .ZN(n14716) );
  OAI211_X1 U18173 ( .C1(n14718), .C2(n14739), .A(n14717), .B(n14716), .ZN(
        n14719) );
  AOI21_X1 U18174 ( .B1(n15364), .B2(n20404), .A(n14719), .ZN(n14720) );
  OAI21_X1 U18175 ( .B1(n15145), .B2(n20393), .A(n14720), .ZN(P1_U2815) );
  INV_X1 U18176 ( .A(n14721), .ZN(n14722) );
  AOI21_X1 U18177 ( .B1(n14722), .B2(n9631), .A(n14706), .ZN(n15155) );
  INV_X1 U18178 ( .A(n15155), .ZN(n15045) );
  NAND2_X1 U18179 ( .A1(n14736), .A2(n14723), .ZN(n14724) );
  AND2_X1 U18180 ( .A1(n14725), .A2(n14724), .ZN(n15374) );
  NOR3_X1 U18181 ( .A1(n20420), .A2(P1_REIP_REG_24__SCAN_IN), .A3(n14726), 
        .ZN(n14729) );
  OAI22_X1 U18182 ( .A1(n9611), .A2(n15153), .B1(n14727), .B2(n20407), .ZN(
        n14728) );
  AOI211_X1 U18183 ( .C1(P1_EBX_REG_24__SCAN_IN), .C2(n20405), .A(n14729), .B(
        n14728), .ZN(n14730) );
  OAI21_X1 U18184 ( .B1(n14731), .B2(n14739), .A(n14730), .ZN(n14732) );
  AOI21_X1 U18185 ( .B1(n15374), .B2(n20404), .A(n14732), .ZN(n14733) );
  OAI21_X1 U18186 ( .B1(n15045), .B2(n20393), .A(n14733), .ZN(P1_U2816) );
  OR2_X1 U18187 ( .A1(n14746), .A2(n14734), .ZN(n14735) );
  NAND2_X1 U18188 ( .A1(n14736), .A2(n14735), .ZN(n14984) );
  INV_X1 U18189 ( .A(n14984), .ZN(n15383) );
  INV_X1 U18190 ( .A(n15163), .ZN(n14737) );
  INV_X1 U18191 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15159) );
  OAI22_X1 U18192 ( .A1(n14969), .A2(n14737), .B1(n15159), .B2(n20407), .ZN(
        n14743) );
  AOI21_X1 U18193 ( .B1(n20376), .B2(n14738), .A(P1_REIP_REG_23__SCAN_IN), 
        .ZN(n14740) );
  NOR2_X1 U18194 ( .A1(n14740), .A2(n14739), .ZN(n14742) );
  NOR2_X1 U18195 ( .A1(n20424), .A2(n14985), .ZN(n14741) );
  OR3_X1 U18196 ( .A1(n14743), .A2(n14742), .A3(n14741), .ZN(n14744) );
  AOI21_X1 U18197 ( .B1(n15383), .B2(n20404), .A(n14744), .ZN(n14745) );
  OAI21_X1 U18198 ( .B1(n15160), .B2(n20393), .A(n14745), .ZN(P1_U2817) );
  INV_X1 U18199 ( .A(n14746), .ZN(n14747) );
  OAI21_X1 U18200 ( .B1(n14748), .B2(n14761), .A(n14747), .ZN(n15388) );
  OR2_X1 U18201 ( .A1(n14749), .A2(n14760), .ZN(n14758) );
  AOI21_X1 U18202 ( .B1(n14750), .B2(n14758), .A(n9663), .ZN(n15171) );
  NAND2_X1 U18203 ( .A1(n15171), .A2(n20383), .ZN(n14757) );
  AOI21_X1 U18204 ( .B1(n14751), .B2(n20410), .A(n14967), .ZN(n14778) );
  INV_X1 U18205 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14986) );
  INV_X1 U18206 ( .A(n14751), .ZN(n14763) );
  OAI21_X1 U18207 ( .B1(n14763), .B2(P1_REIP_REG_22__SCAN_IN), .A(
        P1_REIP_REG_21__SCAN_IN), .ZN(n14752) );
  OAI211_X1 U18208 ( .C1(P1_REIP_REG_21__SCAN_IN), .C2(P1_REIP_REG_22__SCAN_IN), .A(n20376), .B(n14752), .ZN(n14753) );
  OAI21_X1 U18209 ( .B1(n14986), .B2(n20424), .A(n14753), .ZN(n14755) );
  OAI22_X1 U18210 ( .A1(n14969), .A2(n15169), .B1(n21302), .B2(n20407), .ZN(
        n14754) );
  AOI211_X1 U18211 ( .C1(P1_REIP_REG_22__SCAN_IN), .C2(n14778), .A(n14755), 
        .B(n14754), .ZN(n14756) );
  OAI211_X1 U18212 ( .C1(n15388), .C2(n20432), .A(n14757), .B(n14756), .ZN(
        P1_U2818) );
  INV_X1 U18213 ( .A(n14758), .ZN(n14759) );
  AOI21_X1 U18214 ( .B1(n14760), .B2(n14749), .A(n14759), .ZN(n15181) );
  INV_X1 U18215 ( .A(n15181), .ZN(n15057) );
  AOI21_X1 U18216 ( .B1(n14762), .B2(n14774), .A(n14761), .ZN(n15398) );
  INV_X1 U18217 ( .A(n14778), .ZN(n14767) );
  INV_X1 U18218 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n21183) );
  AOI22_X1 U18219 ( .A1(n10405), .A2(n15177), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n20427), .ZN(n14766) );
  NOR3_X1 U18220 ( .A1(n20420), .A2(P1_REIP_REG_21__SCAN_IN), .A3(n14763), 
        .ZN(n14764) );
  AOI21_X1 U18221 ( .B1(P1_EBX_REG_21__SCAN_IN), .B2(n20405), .A(n14764), .ZN(
        n14765) );
  OAI211_X1 U18222 ( .C1(n14767), .C2(n21183), .A(n14766), .B(n14765), .ZN(
        n14768) );
  AOI21_X1 U18223 ( .B1(n15398), .B2(n20404), .A(n14768), .ZN(n14769) );
  OAI21_X1 U18224 ( .B1(n15057), .B2(n20393), .A(n14769), .ZN(P1_U2819) );
  OAI21_X1 U18225 ( .B1(n14771), .B2(n14772), .A(n14749), .ZN(n15188) );
  INV_X1 U18226 ( .A(n14774), .ZN(n14775) );
  AOI21_X1 U18227 ( .B1(n14776), .B2(n14773), .A(n14775), .ZN(n15413) );
  NOR2_X1 U18228 ( .A1(n20420), .A2(n14777), .ZN(n14779) );
  OAI21_X1 U18229 ( .B1(P1_REIP_REG_20__SCAN_IN), .B2(n14779), .A(n14778), 
        .ZN(n14781) );
  AOI22_X1 U18230 ( .A1(n10405), .A2(n15191), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20427), .ZN(n14780) );
  OAI211_X1 U18231 ( .C1(n14782), .C2(n20424), .A(n14781), .B(n14780), .ZN(
        n14783) );
  AOI21_X1 U18232 ( .B1(n15413), .B2(n20404), .A(n14783), .ZN(n14784) );
  OAI21_X1 U18233 ( .B1(n15188), .B2(n20393), .A(n14784), .ZN(P1_U2820) );
  NOR2_X1 U18234 ( .A1(n14785), .A2(n14786), .ZN(n14787) );
  OR2_X1 U18235 ( .A1(n14771), .A2(n14787), .ZN(n15196) );
  OAI21_X1 U18236 ( .B1(n14788), .B2(n14789), .A(n14773), .ZN(n15417) );
  INV_X1 U18237 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n21176) );
  NOR4_X1 U18238 ( .A1(n20420), .A2(P1_REIP_REG_19__SCAN_IN), .A3(n14795), 
        .A4(n21176), .ZN(n14793) );
  NAND2_X1 U18239 ( .A1(n10405), .A2(n15199), .ZN(n14791) );
  NAND2_X1 U18240 ( .A1(n20410), .A2(n14790), .ZN(n20421) );
  OAI211_X1 U18241 ( .C1(n20407), .C2(n15195), .A(n14791), .B(n20421), .ZN(
        n14792) );
  AOI211_X1 U18242 ( .C1(P1_EBX_REG_19__SCAN_IN), .C2(n20405), .A(n14793), .B(
        n14792), .ZN(n14797) );
  INV_X1 U18243 ( .A(n14795), .ZN(n14794) );
  AOI21_X1 U18244 ( .B1(n14794), .B2(n20410), .A(n14967), .ZN(n14816) );
  NOR3_X1 U18245 ( .A1(n20420), .A2(P1_REIP_REG_18__SCAN_IN), .A3(n14795), 
        .ZN(n14803) );
  OAI21_X1 U18246 ( .B1(n14816), .B2(n14803), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n14796) );
  OAI211_X1 U18247 ( .C1(n15417), .C2(n20432), .A(n14797), .B(n14796), .ZN(
        n14798) );
  INV_X1 U18248 ( .A(n14798), .ZN(n14799) );
  OAI21_X1 U18249 ( .B1(n15196), .B2(n20393), .A(n14799), .ZN(P1_U2821) );
  INV_X1 U18250 ( .A(n14800), .ZN(n14802) );
  INV_X1 U18251 ( .A(n14785), .ZN(n14801) );
  AOI21_X1 U18252 ( .B1(n20405), .B2(P1_EBX_REG_18__SCAN_IN), .A(n14803), .ZN(
        n14805) );
  INV_X1 U18253 ( .A(n20421), .ZN(n20368) );
  AOI21_X1 U18254 ( .B1(n20427), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n20368), .ZN(n14804) );
  OAI211_X1 U18255 ( .C1(n15206), .C2(n14969), .A(n14805), .B(n14804), .ZN(
        n14810) );
  NOR2_X1 U18256 ( .A1(n14806), .A2(n14807), .ZN(n14808) );
  OR2_X1 U18257 ( .A1(n14788), .A2(n14808), .ZN(n15440) );
  NOR2_X1 U18258 ( .A1(n15440), .A2(n20432), .ZN(n14809) );
  AOI211_X1 U18259 ( .C1(n14816), .C2(P1_REIP_REG_18__SCAN_IN), .A(n14810), 
        .B(n14809), .ZN(n14811) );
  OAI21_X1 U18260 ( .B1(n15204), .B2(n20393), .A(n14811), .ZN(P1_U2822) );
  AOI21_X1 U18261 ( .B1(n14813), .B2(n9593), .A(n9635), .ZN(n15227) );
  INV_X1 U18262 ( .A(n15227), .ZN(n15075) );
  AND2_X1 U18263 ( .A1(n14830), .A2(n14814), .ZN(n14815) );
  NOR2_X1 U18264 ( .A1(n14806), .A2(n14815), .ZN(n15450) );
  INV_X1 U18265 ( .A(n14816), .ZN(n14823) );
  NAND2_X1 U18266 ( .A1(n20376), .A2(n14837), .ZN(n20356) );
  INV_X1 U18267 ( .A(n20356), .ZN(n14817) );
  AOI21_X1 U18268 ( .B1(n14818), .B2(n14817), .A(P1_REIP_REG_17__SCAN_IN), 
        .ZN(n14822) );
  AOI21_X1 U18269 ( .B1(n20427), .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n20368), .ZN(n14819) );
  OAI21_X1 U18270 ( .B1(n9611), .B2(n15225), .A(n14819), .ZN(n14820) );
  AOI21_X1 U18271 ( .B1(n20405), .B2(P1_EBX_REG_17__SCAN_IN), .A(n14820), .ZN(
        n14821) );
  OAI21_X1 U18272 ( .B1(n14823), .B2(n14822), .A(n14821), .ZN(n14824) );
  AOI21_X1 U18273 ( .B1(n15450), .B2(n20404), .A(n14824), .ZN(n14825) );
  OAI21_X1 U18274 ( .B1(n15075), .B2(n20393), .A(n14825), .ZN(P1_U2823) );
  OAI21_X1 U18275 ( .B1(n14826), .B2(n14827), .A(n9593), .ZN(n15240) );
  OAI21_X1 U18276 ( .B1(n14828), .B2(n14853), .A(n14829), .ZN(n14831) );
  NAND2_X1 U18277 ( .A1(n14831), .A2(n14830), .ZN(n15460) );
  INV_X1 U18278 ( .A(n15460), .ZN(n14847) );
  AND2_X1 U18279 ( .A1(n14835), .A2(n14832), .ZN(n14834) );
  OR2_X1 U18280 ( .A1(n20420), .A2(n14837), .ZN(n14833) );
  NAND2_X1 U18281 ( .A1(n14833), .A2(n20410), .ZN(n20371) );
  NOR2_X1 U18282 ( .A1(n14834), .A2(n20371), .ZN(n14885) );
  INV_X1 U18283 ( .A(n14885), .ZN(n14935) );
  AOI21_X1 U18284 ( .B1(n14855), .B2(n14835), .A(n14935), .ZN(n14868) );
  INV_X1 U18285 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n21174) );
  NAND2_X1 U18286 ( .A1(n20427), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14836) );
  OAI211_X1 U18287 ( .C1(n14969), .C2(n15236), .A(n20421), .B(n14836), .ZN(
        n14844) );
  NAND2_X1 U18288 ( .A1(n14837), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n14838) );
  OR2_X1 U18289 ( .A1(n20420), .A2(n14838), .ZN(n14931) );
  INV_X1 U18290 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n14839) );
  NOR2_X1 U18291 ( .A1(n14931), .A2(n14839), .ZN(n14913) );
  INV_X1 U18292 ( .A(n14913), .ZN(n14902) );
  INV_X1 U18293 ( .A(n14855), .ZN(n14840) );
  OAI211_X1 U18294 ( .C1(P1_REIP_REG_16__SCAN_IN), .C2(P1_REIP_REG_15__SCAN_IN), .A(n14841), .B(n14840), .ZN(n14842) );
  NOR2_X1 U18295 ( .A1(n14902), .A2(n14842), .ZN(n14843) );
  AOI211_X1 U18296 ( .C1(P1_EBX_REG_16__SCAN_IN), .C2(n20405), .A(n14844), .B(
        n14843), .ZN(n14845) );
  OAI21_X1 U18297 ( .B1(n14868), .B2(n21174), .A(n14845), .ZN(n14846) );
  AOI21_X1 U18298 ( .B1(n20404), .B2(n14847), .A(n14846), .ZN(n14848) );
  OAI21_X1 U18299 ( .B1(n15240), .B2(n20393), .A(n14848), .ZN(P1_U2824) );
  INV_X1 U18300 ( .A(n14918), .ZN(n14876) );
  OAI21_X1 U18301 ( .B1(n14876), .B2(n14849), .A(n14875), .ZN(n14850) );
  NAND2_X1 U18302 ( .A1(n14878), .A2(n14865), .ZN(n14864) );
  INV_X1 U18303 ( .A(n14851), .ZN(n14852) );
  AOI21_X1 U18304 ( .B1(n14864), .B2(n14852), .A(n14826), .ZN(n15247) );
  INV_X1 U18305 ( .A(n15247), .ZN(n15086) );
  XNOR2_X1 U18306 ( .A(n14828), .B(n14853), .ZN(n15463) );
  INV_X1 U18307 ( .A(n15463), .ZN(n14860) );
  INV_X1 U18308 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n21171) );
  NAND2_X1 U18309 ( .A1(n20427), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14854) );
  OAI211_X1 U18310 ( .C1(n9611), .C2(n15245), .A(n20421), .B(n14854), .ZN(
        n14857) );
  NOR3_X1 U18311 ( .A1(n14902), .A2(P1_REIP_REG_15__SCAN_IN), .A3(n14855), 
        .ZN(n14856) );
  AOI211_X1 U18312 ( .C1(P1_EBX_REG_15__SCAN_IN), .C2(n20405), .A(n14857), .B(
        n14856), .ZN(n14858) );
  OAI21_X1 U18313 ( .B1(n14868), .B2(n21171), .A(n14858), .ZN(n14859) );
  AOI21_X1 U18314 ( .B1(n20404), .B2(n14860), .A(n14859), .ZN(n14861) );
  OAI21_X1 U18315 ( .B1(n15086), .B2(n20393), .A(n14861), .ZN(P1_U2825) );
  OR2_X1 U18316 ( .A1(n14880), .A2(n14862), .ZN(n14863) );
  NAND2_X1 U18317 ( .A1(n14828), .A2(n14863), .ZN(n15476) );
  OAI21_X1 U18318 ( .B1(n14878), .B2(n14865), .A(n14864), .ZN(n15258) );
  INV_X1 U18319 ( .A(n15258), .ZN(n14866) );
  NAND2_X1 U18320 ( .A1(n14866), .A2(n20383), .ZN(n14873) );
  NAND2_X1 U18321 ( .A1(n20427), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14867) );
  OAI211_X1 U18322 ( .C1(n9611), .C2(n15254), .A(n20421), .B(n14867), .ZN(
        n14871) );
  INV_X1 U18323 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n15253) );
  NAND3_X1 U18324 ( .A1(n14913), .A2(P1_REIP_REG_11__SCAN_IN), .A3(
        P1_REIP_REG_12__SCAN_IN), .ZN(n14889) );
  INV_X1 U18325 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n21169) );
  OR2_X1 U18326 ( .A1(n14889), .A2(n21169), .ZN(n14869) );
  AOI21_X1 U18327 ( .B1(n15253), .B2(n14869), .A(n14868), .ZN(n14870) );
  AOI211_X1 U18328 ( .C1(P1_EBX_REG_14__SCAN_IN), .C2(n20405), .A(n14871), .B(
        n14870), .ZN(n14872) );
  OAI211_X1 U18329 ( .C1(n15476), .C2(n20432), .A(n14873), .B(n14872), .ZN(
        P1_U2826) );
  OAI21_X1 U18330 ( .B1(n14925), .B2(n14874), .A(n14875), .ZN(n14919) );
  OAI21_X1 U18331 ( .B1(n14919), .B2(n14876), .A(n14875), .ZN(n14894) );
  NAND2_X1 U18332 ( .A1(n14894), .A2(n14893), .ZN(n14892) );
  INV_X1 U18333 ( .A(n14877), .ZN(n14879) );
  AOI21_X1 U18334 ( .B1(n14892), .B2(n14879), .A(n14878), .ZN(n15271) );
  INV_X1 U18335 ( .A(n15271), .ZN(n15089) );
  AOI21_X1 U18336 ( .B1(n14881), .B2(n14897), .A(n14880), .ZN(n15485) );
  NAND2_X1 U18337 ( .A1(n20427), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14882) );
  OAI211_X1 U18338 ( .C1(n14969), .C2(n15269), .A(n20421), .B(n14882), .ZN(
        n14883) );
  AOI21_X1 U18339 ( .B1(n20405), .B2(P1_EBX_REG_13__SCAN_IN), .A(n14883), .ZN(
        n14888) );
  INV_X1 U18340 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n14884) );
  INV_X1 U18341 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n14912) );
  NOR2_X1 U18342 ( .A1(n14884), .A2(n14912), .ZN(n14886) );
  OAI21_X1 U18343 ( .B1(n14967), .B2(n14886), .A(n14885), .ZN(n14903) );
  NAND2_X1 U18344 ( .A1(n14903), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n14887) );
  OAI211_X1 U18345 ( .C1(P1_REIP_REG_13__SCAN_IN), .C2(n14889), .A(n14888), 
        .B(n14887), .ZN(n14890) );
  AOI21_X1 U18346 ( .B1(n20404), .B2(n15485), .A(n14890), .ZN(n14891) );
  OAI21_X1 U18347 ( .B1(n15089), .B2(n20393), .A(n14891), .ZN(P1_U2827) );
  OAI21_X1 U18348 ( .B1(n14894), .B2(n14893), .A(n14892), .ZN(n15280) );
  NAND2_X1 U18349 ( .A1(n20427), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14895) );
  OAI211_X1 U18350 ( .C1(n14969), .C2(n15276), .A(n20421), .B(n14895), .ZN(
        n14901) );
  AOI21_X1 U18351 ( .B1(n14898), .B2(n14896), .A(n10241), .ZN(n15499) );
  INV_X1 U18352 ( .A(n15499), .ZN(n14899) );
  NOR2_X1 U18353 ( .A1(n14899), .A2(n20432), .ZN(n14900) );
  AOI211_X1 U18354 ( .C1(P1_EBX_REG_12__SCAN_IN), .C2(n20405), .A(n14901), .B(
        n14900), .ZN(n14906) );
  NOR2_X1 U18355 ( .A1(n14902), .A2(n14912), .ZN(n14904) );
  OAI21_X1 U18356 ( .B1(n14904), .B2(P1_REIP_REG_12__SCAN_IN), .A(n14903), 
        .ZN(n14905) );
  OAI211_X1 U18357 ( .C1(n15280), .C2(n20393), .A(n14906), .B(n14905), .ZN(
        P1_U2828) );
  NAND2_X1 U18358 ( .A1(n20427), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n14907) );
  OAI211_X1 U18359 ( .C1(n14969), .C2(n15285), .A(n20421), .B(n14907), .ZN(
        n14908) );
  INV_X1 U18360 ( .A(n14908), .ZN(n14917) );
  OR2_X1 U18361 ( .A1(n14909), .A2(n14910), .ZN(n14911) );
  NAND2_X1 U18362 ( .A1(n14896), .A2(n14911), .ZN(n15505) );
  OR2_X1 U18363 ( .A1(n15505), .A2(n20432), .ZN(n14916) );
  NAND2_X1 U18364 ( .A1(n14913), .A2(n14912), .ZN(n14915) );
  OR2_X1 U18365 ( .A1(n20424), .A2(n14998), .ZN(n14914) );
  NAND4_X1 U18366 ( .A1(n14917), .A2(n14916), .A3(n14915), .A4(n14914), .ZN(
        n14921) );
  XNOR2_X1 U18367 ( .A(n14919), .B(n14918), .ZN(n15287) );
  INV_X1 U18368 ( .A(n15287), .ZN(n15092) );
  NOR2_X1 U18369 ( .A1(n15092), .A2(n20393), .ZN(n14920) );
  AOI211_X1 U18370 ( .C1(P1_REIP_REG_11__SCAN_IN), .C2(n14935), .A(n14921), 
        .B(n14920), .ZN(n14922) );
  INV_X1 U18371 ( .A(n14922), .ZN(P1_U2829) );
  AOI21_X1 U18372 ( .B1(n14926), .B2(n14924), .A(n14925), .ZN(n15299) );
  INV_X1 U18373 ( .A(n15299), .ZN(n15095) );
  NOR2_X1 U18374 ( .A1(n9746), .A2(n14927), .ZN(n14928) );
  OR2_X1 U18375 ( .A1(n14909), .A2(n14928), .ZN(n15526) );
  INV_X1 U18376 ( .A(n15526), .ZN(n14929) );
  AOI22_X1 U18377 ( .A1(n20404), .A2(n14929), .B1(n20405), .B2(
        P1_EBX_REG_10__SCAN_IN), .ZN(n14930) );
  OAI21_X1 U18378 ( .B1(P1_REIP_REG_10__SCAN_IN), .B2(n14931), .A(n14930), 
        .ZN(n14932) );
  AOI211_X1 U18379 ( .C1(n20427), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n14932), .B(n20368), .ZN(n14933) );
  OAI21_X1 U18380 ( .B1(n9611), .B2(n15297), .A(n14933), .ZN(n14934) );
  AOI21_X1 U18381 ( .B1(n14935), .B2(P1_REIP_REG_10__SCAN_IN), .A(n14934), 
        .ZN(n14936) );
  OAI21_X1 U18382 ( .B1(n15095), .B2(n20393), .A(n14936), .ZN(P1_U2830) );
  INV_X1 U18383 ( .A(n14939), .ZN(n14937) );
  NOR2_X1 U18384 ( .A1(n14939), .A2(n14938), .ZN(n20429) );
  NAND2_X1 U18385 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n14943) );
  NAND2_X1 U18386 ( .A1(n20376), .A2(n14943), .ZN(n14958) );
  NAND2_X1 U18387 ( .A1(n20410), .A2(n14958), .ZN(n14948) );
  AOI22_X1 U18388 ( .A1(n20427), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n14948), .ZN(n14941) );
  AOI22_X1 U18389 ( .A1(n20405), .A2(P1_EBX_REG_3__SCAN_IN), .B1(n20404), .B2(
        n20534), .ZN(n14940) );
  OAI211_X1 U18390 ( .C1(n14969), .C2(n14942), .A(n14941), .B(n14940), .ZN(
        n14945) );
  NOR3_X1 U18391 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n20420), .A3(n14943), .ZN(
        n14944) );
  AOI211_X1 U18392 ( .C1(n20429), .C2(n20839), .A(n14945), .B(n14944), .ZN(
        n14946) );
  OAI21_X1 U18393 ( .B1(n20433), .B2(n14947), .A(n14946), .ZN(P1_U2837) );
  INV_X1 U18394 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n21206) );
  INV_X1 U18395 ( .A(n20433), .ZN(n20411) );
  AOI22_X1 U18396 ( .A1(n20427), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n14948), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n14950) );
  INV_X1 U18397 ( .A(n13947), .ZN(n20593) );
  NAND2_X1 U18398 ( .A1(n20429), .A2(n20593), .ZN(n14949) );
  OAI211_X1 U18399 ( .C1(n9611), .C2(n14951), .A(n14950), .B(n14949), .ZN(
        n14955) );
  OAI22_X1 U18400 ( .A1(n20432), .A2(n14953), .B1(n14952), .B2(n20424), .ZN(
        n14954) );
  AOI211_X1 U18401 ( .C1(n14956), .C2(n20411), .A(n14955), .B(n14954), .ZN(
        n14957) );
  OAI21_X1 U18402 ( .B1(n14958), .B2(n21206), .A(n14957), .ZN(P1_U2838) );
  INV_X1 U18403 ( .A(n20429), .ZN(n14961) );
  OAI22_X1 U18404 ( .A1(n14961), .A2(n14960), .B1(n21206), .B2(n20410), .ZN(
        n14963) );
  OAI22_X1 U18405 ( .A1(n20432), .A2(n20556), .B1(P1_REIP_REG_1__SCAN_IN), 
        .B2(n20420), .ZN(n14962) );
  AOI211_X1 U18406 ( .C1(n20405), .C2(P1_EBX_REG_1__SCAN_IN), .A(n14963), .B(
        n14962), .ZN(n14965) );
  MUX2_X1 U18407 ( .A(n14969), .B(n20407), .S(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n14964) );
  OAI211_X1 U18408 ( .C1(n20433), .C2(n15312), .A(n14965), .B(n14964), .ZN(
        P1_U2839) );
  INV_X1 U18409 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n14966) );
  NOR2_X1 U18410 ( .A1(n14967), .A2(n14966), .ZN(n14971) );
  INV_X1 U18411 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14968) );
  AOI21_X1 U18412 ( .B1(n9611), .B2(n20407), .A(n14968), .ZN(n14970) );
  AOI211_X1 U18413 ( .C1(n20404), .C2(n14972), .A(n14971), .B(n14970), .ZN(
        n14974) );
  AOI22_X1 U18414 ( .A1(n20405), .A2(P1_EBX_REG_0__SCAN_IN), .B1(n21386), .B2(
        n20429), .ZN(n14973) );
  OAI211_X1 U18415 ( .C1(n20433), .C2(n14975), .A(n14974), .B(n14973), .ZN(
        P1_U2840) );
  INV_X1 U18416 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14978) );
  OAI222_X1 U18417 ( .A1(n15011), .A2(n15025), .B1(n14978), .B2(n20447), .C1(
        n15013), .C2(n14977), .ZN(P1_U2843) );
  OAI222_X1 U18418 ( .A1(n15011), .A2(n15032), .B1(n14979), .B2(n20447), .C1(
        n15346), .C2(n15013), .ZN(P1_U2845) );
  OAI222_X1 U18419 ( .A1(n15132), .A2(n15011), .B1(n14981), .B2(n20447), .C1(
        n14980), .C2(n15013), .ZN(P1_U2846) );
  AOI22_X1 U18420 ( .A1(n15364), .A2(n20439), .B1(P1_EBX_REG_25__SCAN_IN), 
        .B2(n14996), .ZN(n14982) );
  OAI21_X1 U18421 ( .B1(n15145), .B2(n15011), .A(n14982), .ZN(P1_U2847) );
  AOI22_X1 U18422 ( .A1(n15374), .A2(n20439), .B1(P1_EBX_REG_24__SCAN_IN), 
        .B2(n14996), .ZN(n14983) );
  OAI21_X1 U18423 ( .B1(n15045), .B2(n15011), .A(n14983), .ZN(P1_U2848) );
  OAI222_X1 U18424 ( .A1(n15160), .A2(n15011), .B1(n14985), .B2(n20447), .C1(
        n14984), .C2(n15013), .ZN(P1_U2849) );
  INV_X1 U18425 ( .A(n15171), .ZN(n15053) );
  OAI222_X1 U18426 ( .A1(n15053), .A2(n15011), .B1(n14986), .B2(n20447), .C1(
        n15388), .C2(n15013), .ZN(P1_U2850) );
  AOI22_X1 U18427 ( .A1(n15398), .A2(n20439), .B1(P1_EBX_REG_21__SCAN_IN), 
        .B2(n14996), .ZN(n14987) );
  OAI21_X1 U18428 ( .B1(n15057), .B2(n15011), .A(n14987), .ZN(P1_U2851) );
  AOI22_X1 U18429 ( .A1(n15413), .A2(n20439), .B1(P1_EBX_REG_20__SCAN_IN), 
        .B2(n14996), .ZN(n14988) );
  OAI21_X1 U18430 ( .B1(n15188), .B2(n15011), .A(n14988), .ZN(P1_U2852) );
  OAI222_X1 U18431 ( .A1(n15196), .A2(n15011), .B1(n14989), .B2(n20447), .C1(
        n15417), .C2(n15013), .ZN(P1_U2853) );
  INV_X1 U18432 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14990) );
  OAI222_X1 U18433 ( .A1(n15204), .A2(n15011), .B1(n14990), .B2(n20447), .C1(
        n15440), .C2(n15013), .ZN(P1_U2854) );
  AOI22_X1 U18434 ( .A1(n15450), .A2(n20439), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n14996), .ZN(n14991) );
  OAI21_X1 U18435 ( .B1(n15075), .B2(n15011), .A(n14991), .ZN(P1_U2855) );
  INV_X1 U18436 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14992) );
  OAI222_X1 U18437 ( .A1(n15240), .A2(n15011), .B1(n14992), .B2(n20447), .C1(
        n15460), .C2(n15013), .ZN(P1_U2856) );
  OAI222_X1 U18438 ( .A1(n15086), .A2(n15011), .B1(n14993), .B2(n20447), .C1(
        n15013), .C2(n15463), .ZN(P1_U2857) );
  INV_X1 U18439 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n14994) );
  OAI222_X1 U18440 ( .A1(n15258), .A2(n15011), .B1(n14994), .B2(n20447), .C1(
        n15476), .C2(n15013), .ZN(P1_U2858) );
  AOI22_X1 U18441 ( .A1(n15485), .A2(n20439), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n14996), .ZN(n14995) );
  OAI21_X1 U18442 ( .B1(n15089), .B2(n15011), .A(n14995), .ZN(P1_U2859) );
  AOI22_X1 U18443 ( .A1(n15499), .A2(n20439), .B1(P1_EBX_REG_12__SCAN_IN), 
        .B2(n14996), .ZN(n14997) );
  OAI21_X1 U18444 ( .B1(n15280), .B2(n15011), .A(n14997), .ZN(P1_U2860) );
  OAI22_X1 U18445 ( .A1(n15505), .A2(n15013), .B1(n14998), .B2(n20447), .ZN(
        n14999) );
  AOI21_X1 U18446 ( .B1(n15287), .B2(n20440), .A(n14999), .ZN(n15000) );
  INV_X1 U18447 ( .A(n15000), .ZN(P1_U2861) );
  INV_X1 U18448 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n15001) );
  OAI222_X1 U18449 ( .A1(n15095), .A2(n15011), .B1(n15001), .B2(n20447), .C1(
        n15526), .C2(n15013), .ZN(P1_U2862) );
  AOI21_X1 U18450 ( .B1(n15002), .B2(n14461), .A(n12740), .ZN(n20361) );
  INV_X1 U18451 ( .A(n20361), .ZN(n15097) );
  AND2_X1 U18452 ( .A1(n15003), .A2(n15004), .ZN(n15005) );
  OR2_X1 U18453 ( .A1(n15005), .A2(n9746), .ZN(n20357) );
  OAI222_X1 U18454 ( .A1(n15097), .A2(n15011), .B1(n15006), .B2(n20447), .C1(
        n20357), .C2(n15013), .ZN(P1_U2863) );
  AND2_X1 U18455 ( .A1(n15008), .A2(n15007), .ZN(n15009) );
  OAI222_X1 U18456 ( .A1(n20379), .A2(n15013), .B1(n15012), .B2(n20447), .C1(
        n20382), .C2(n15011), .ZN(P1_U2865) );
  INV_X1 U18457 ( .A(DATAI_14_), .ZN(n15015) );
  INV_X1 U18458 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n15014) );
  MUX2_X1 U18459 ( .A(n15015), .B(n15014), .S(n20584), .Z(n20491) );
  OAI22_X1 U18460 ( .A1(n15070), .A2(n20491), .B1(n15098), .B2(n15016), .ZN(
        n15017) );
  AOI21_X1 U18461 ( .B1(BUF1_REG_30__SCAN_IN), .B2(n15072), .A(n15017), .ZN(
        n15019) );
  NAND2_X1 U18462 ( .A1(n15082), .A2(DATAI_30_), .ZN(n15018) );
  OAI211_X1 U18463 ( .C1(n9596), .C2(n15101), .A(n15019), .B(n15018), .ZN(
        P1_U2874) );
  INV_X1 U18464 ( .A(DATAI_13_), .ZN(n15020) );
  MUX2_X1 U18465 ( .A(n15020), .B(n17298), .S(n20584), .Z(n20488) );
  OAI22_X1 U18466 ( .A1(n15070), .A2(n20488), .B1(n15098), .B2(n15021), .ZN(
        n15022) );
  AOI21_X1 U18467 ( .B1(BUF1_REG_29__SCAN_IN), .B2(n15072), .A(n15022), .ZN(
        n15024) );
  NAND2_X1 U18468 ( .A1(n15082), .A2(DATAI_29_), .ZN(n15023) );
  OAI211_X1 U18469 ( .C1(n15025), .C2(n15101), .A(n15024), .B(n15023), .ZN(
        P1_U2875) );
  INV_X1 U18470 ( .A(DATAI_11_), .ZN(n15027) );
  MUX2_X1 U18471 ( .A(n15027), .B(n15026), .S(n20584), .Z(n20482) );
  OAI22_X1 U18472 ( .A1(n15070), .A2(n20482), .B1(n15098), .B2(n15028), .ZN(
        n15029) );
  AOI21_X1 U18473 ( .B1(BUF1_REG_27__SCAN_IN), .B2(n15072), .A(n15029), .ZN(
        n15031) );
  NAND2_X1 U18474 ( .A1(n15082), .A2(DATAI_27_), .ZN(n15030) );
  OAI211_X1 U18475 ( .C1(n15032), .C2(n15101), .A(n15031), .B(n15030), .ZN(
        P1_U2877) );
  OAI22_X1 U18476 ( .A1(n15070), .A2(n15094), .B1(n15098), .B2(n15033), .ZN(
        n15034) );
  AOI21_X1 U18477 ( .B1(BUF1_REG_26__SCAN_IN), .B2(n15072), .A(n15034), .ZN(
        n15036) );
  NAND2_X1 U18478 ( .A1(n15082), .A2(DATAI_26_), .ZN(n15035) );
  OAI211_X1 U18479 ( .C1(n15132), .C2(n15101), .A(n15036), .B(n15035), .ZN(
        P1_U2878) );
  INV_X1 U18480 ( .A(DATAI_9_), .ZN(n15037) );
  MUX2_X1 U18481 ( .A(n15037), .B(n17304), .S(n20584), .Z(n20479) );
  OAI22_X1 U18482 ( .A1(n15070), .A2(n20479), .B1(n15098), .B2(n15038), .ZN(
        n15039) );
  AOI21_X1 U18483 ( .B1(n15072), .B2(BUF1_REG_25__SCAN_IN), .A(n15039), .ZN(
        n15041) );
  NAND2_X1 U18484 ( .A1(n15082), .A2(DATAI_25_), .ZN(n15040) );
  OAI211_X1 U18485 ( .C1(n15145), .C2(n15101), .A(n15041), .B(n15040), .ZN(
        P1_U2879) );
  OAI22_X1 U18486 ( .A1(n15070), .A2(n20476), .B1(n15098), .B2(n14083), .ZN(
        n15042) );
  AOI21_X1 U18487 ( .B1(n15072), .B2(BUF1_REG_24__SCAN_IN), .A(n15042), .ZN(
        n15044) );
  NAND2_X1 U18488 ( .A1(n15082), .A2(DATAI_24_), .ZN(n15043) );
  OAI211_X1 U18489 ( .C1(n15045), .C2(n15101), .A(n15044), .B(n15043), .ZN(
        P1_U2880) );
  OAI22_X1 U18490 ( .A1(n15070), .A2(n20630), .B1(n15098), .B2(n14097), .ZN(
        n15046) );
  AOI21_X1 U18491 ( .B1(n15072), .B2(BUF1_REG_23__SCAN_IN), .A(n15046), .ZN(
        n15048) );
  NAND2_X1 U18492 ( .A1(n15082), .A2(DATAI_23_), .ZN(n15047) );
  OAI211_X1 U18493 ( .C1(n15160), .C2(n15101), .A(n15048), .B(n15047), .ZN(
        P1_U2881) );
  INV_X1 U18494 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n19632) );
  INV_X1 U18495 ( .A(n15070), .ZN(n15078) );
  AOI22_X1 U18496 ( .A1(n15078), .A2(n15049), .B1(P1_EAX_REG_22__SCAN_IN), 
        .B2(n15076), .ZN(n15050) );
  OAI21_X1 U18497 ( .B1(n15080), .B2(n19632), .A(n15050), .ZN(n15051) );
  AOI21_X1 U18498 ( .B1(n15082), .B2(DATAI_22_), .A(n15051), .ZN(n15052) );
  OAI21_X1 U18499 ( .B1(n15053), .B2(n15101), .A(n15052), .ZN(P1_U2882) );
  OAI22_X1 U18500 ( .A1(n15070), .A2(n20619), .B1(n15098), .B2(n14094), .ZN(
        n15054) );
  AOI21_X1 U18501 ( .B1(n15072), .B2(BUF1_REG_21__SCAN_IN), .A(n15054), .ZN(
        n15056) );
  NAND2_X1 U18502 ( .A1(n15082), .A2(DATAI_21_), .ZN(n15055) );
  OAI211_X1 U18503 ( .C1(n15057), .C2(n15101), .A(n15056), .B(n15055), .ZN(
        P1_U2883) );
  INV_X1 U18504 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n17287) );
  AOI22_X1 U18505 ( .A1(n15078), .A2(n15058), .B1(P1_EAX_REG_20__SCAN_IN), 
        .B2(n15076), .ZN(n15059) );
  OAI21_X1 U18506 ( .B1(n15080), .B2(n17287), .A(n15059), .ZN(n15060) );
  AOI21_X1 U18507 ( .B1(n15082), .B2(DATAI_20_), .A(n15060), .ZN(n15061) );
  OAI21_X1 U18508 ( .B1(n15188), .B2(n15101), .A(n15061), .ZN(P1_U2884) );
  OAI22_X1 U18509 ( .A1(n15070), .A2(n20612), .B1(n15098), .B2(n14090), .ZN(
        n15062) );
  AOI21_X1 U18510 ( .B1(n15072), .B2(BUF1_REG_19__SCAN_IN), .A(n15062), .ZN(
        n15064) );
  NAND2_X1 U18511 ( .A1(n15082), .A2(DATAI_19_), .ZN(n15063) );
  OAI211_X1 U18512 ( .C1(n15196), .C2(n15101), .A(n15064), .B(n15063), .ZN(
        P1_U2885) );
  OAI22_X1 U18513 ( .A1(n15070), .A2(n20608), .B1(n15098), .B2(n15065), .ZN(
        n15066) );
  AOI21_X1 U18514 ( .B1(n15072), .B2(BUF1_REG_18__SCAN_IN), .A(n15066), .ZN(
        n15068) );
  NAND2_X1 U18515 ( .A1(n15082), .A2(DATAI_18_), .ZN(n15067) );
  OAI211_X1 U18516 ( .C1(n15204), .C2(n15101), .A(n15068), .B(n15067), .ZN(
        P1_U2886) );
  OAI22_X1 U18517 ( .A1(n15070), .A2(n20604), .B1(n15098), .B2(n15069), .ZN(
        n15071) );
  AOI21_X1 U18518 ( .B1(n15072), .B2(BUF1_REG_17__SCAN_IN), .A(n15071), .ZN(
        n15074) );
  NAND2_X1 U18519 ( .A1(n15082), .A2(DATAI_17_), .ZN(n15073) );
  OAI211_X1 U18520 ( .C1(n15075), .C2(n15101), .A(n15074), .B(n15073), .ZN(
        P1_U2887) );
  INV_X1 U18521 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n17294) );
  AOI22_X1 U18522 ( .A1(n15078), .A2(n15077), .B1(P1_EAX_REG_16__SCAN_IN), 
        .B2(n15076), .ZN(n15079) );
  OAI21_X1 U18523 ( .B1(n15080), .B2(n17294), .A(n15079), .ZN(n15081) );
  AOI21_X1 U18524 ( .B1(n15082), .B2(DATAI_16_), .A(n15081), .ZN(n15083) );
  OAI21_X1 U18525 ( .B1(n15240), .B2(n15101), .A(n15083), .ZN(P1_U2888) );
  OAI222_X1 U18526 ( .A1(n15086), .A2(n15101), .B1(n15098), .B2(n15085), .C1(
        n15100), .C2(n15084), .ZN(P1_U2889) );
  INV_X1 U18527 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n15087) );
  OAI222_X1 U18528 ( .A1(n15258), .A2(n15101), .B1(n20491), .B2(n15100), .C1(
        n15087), .C2(n15098), .ZN(P1_U2890) );
  INV_X1 U18529 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n15088) );
  OAI222_X1 U18530 ( .A1(n15089), .A2(n15101), .B1(n20488), .B2(n15100), .C1(
        n15088), .C2(n15098), .ZN(P1_U2891) );
  INV_X1 U18531 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n15090) );
  OAI222_X1 U18532 ( .A1(n15280), .A2(n15101), .B1(n20485), .B2(n15100), .C1(
        n15090), .C2(n15098), .ZN(P1_U2892) );
  INV_X1 U18533 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n15091) );
  OAI222_X1 U18534 ( .A1(n15092), .A2(n15101), .B1(n20482), .B2(n15100), .C1(
        n15091), .C2(n15098), .ZN(P1_U2893) );
  INV_X1 U18535 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n15093) );
  OAI222_X1 U18536 ( .A1(n15101), .A2(n15095), .B1(n15094), .B2(n15100), .C1(
        n15093), .C2(n15098), .ZN(P1_U2894) );
  INV_X1 U18537 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n15096) );
  OAI222_X1 U18538 ( .A1(n15097), .A2(n15101), .B1(n20479), .B2(n15100), .C1(
        n15096), .C2(n15098), .ZN(P1_U2895) );
  INV_X1 U18539 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n15099) );
  OAI222_X1 U18540 ( .A1(n20382), .A2(n15101), .B1(n20630), .B2(n15100), .C1(
        n15099), .C2(n15098), .ZN(P1_U2897) );
  INV_X1 U18541 ( .A(n15102), .ZN(n15105) );
  INV_X1 U18542 ( .A(n15114), .ZN(n15103) );
  NAND2_X1 U18543 ( .A1(n15107), .A2(n15200), .ZN(n15108) );
  NAND2_X1 U18544 ( .A1(n20526), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n15322) );
  OAI211_X1 U18545 ( .C1(n17161), .C2(n15109), .A(n15108), .B(n15322), .ZN(
        n15110) );
  OAI21_X1 U18546 ( .B1(n15324), .B2(n20338), .A(n15112), .ZN(P1_U2969) );
  NAND2_X1 U18547 ( .A1(n20526), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n15327) );
  NAND2_X1 U18548 ( .A1(n20511), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15115) );
  OAI211_X1 U18549 ( .C1(n15116), .C2(n9869), .A(n15327), .B(n15115), .ZN(
        n15117) );
  AOI21_X1 U18550 ( .B1(n15118), .B2(n20518), .A(n15117), .ZN(n15119) );
  OAI21_X1 U18551 ( .B1(n20338), .B2(n15333), .A(n15119), .ZN(P1_U2970) );
  INV_X1 U18552 ( .A(n15120), .ZN(n15121) );
  XNOR2_X1 U18553 ( .A(n15122), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15350) );
  NOR2_X1 U18554 ( .A1(n15267), .A2(n15123), .ZN(n15344) );
  AOI21_X1 U18555 ( .B1(n20511), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15344), .ZN(n15124) );
  OAI21_X1 U18556 ( .B1(n15125), .B2(n9869), .A(n15124), .ZN(n15126) );
  AOI21_X1 U18557 ( .B1(n15127), .B2(n20518), .A(n15126), .ZN(n15128) );
  OAI21_X1 U18558 ( .B1(n20338), .B2(n15350), .A(n15128), .ZN(P1_U2972) );
  OAI211_X1 U18559 ( .C1(n10374), .C2(n15158), .A(n15130), .B(n15129), .ZN(
        n15131) );
  XOR2_X1 U18560 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n15131), .Z(
        n15358) );
  INV_X1 U18561 ( .A(n15132), .ZN(n15136) );
  NAND2_X1 U18562 ( .A1(n20526), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n15352) );
  NAND2_X1 U18563 ( .A1(n20511), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15133) );
  OAI211_X1 U18564 ( .C1(n9869), .C2(n15134), .A(n15352), .B(n15133), .ZN(
        n15135) );
  AOI21_X1 U18565 ( .B1(n15136), .B2(n20518), .A(n15135), .ZN(n15137) );
  OAI21_X1 U18566 ( .B1(n20338), .B2(n15358), .A(n15137), .ZN(P1_U2973) );
  NAND2_X1 U18567 ( .A1(n14535), .A2(n15138), .ZN(n15141) );
  NAND2_X1 U18568 ( .A1(n15150), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15140) );
  MUX2_X1 U18569 ( .A(n15141), .B(n15140), .S(n9569), .Z(n15143) );
  XNOR2_X1 U18570 ( .A(n15143), .B(n15142), .ZN(n15366) );
  INV_X1 U18571 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15144) );
  NAND2_X1 U18572 ( .A1(n20577), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n15360) );
  OAI21_X1 U18573 ( .B1(n17161), .B2(n15144), .A(n15360), .ZN(n15146) );
  OAI21_X1 U18574 ( .B1(n20338), .B2(n15366), .A(n15148), .ZN(P1_U2974) );
  NOR2_X1 U18575 ( .A1(n15150), .A2(n15158), .ZN(n15149) );
  MUX2_X1 U18576 ( .A(n15150), .B(n15149), .S(n10374), .Z(n15151) );
  XNOR2_X1 U18577 ( .A(n15151), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15376) );
  NAND2_X1 U18578 ( .A1(n20526), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n15371) );
  NAND2_X1 U18579 ( .A1(n20511), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15152) );
  OAI211_X1 U18580 ( .C1(n9869), .C2(n15153), .A(n15371), .B(n15152), .ZN(
        n15154) );
  AOI21_X1 U18581 ( .B1(n15155), .B2(n20518), .A(n15154), .ZN(n15156) );
  OAI21_X1 U18582 ( .B1(n20338), .B2(n15376), .A(n15156), .ZN(P1_U2975) );
  XNOR2_X1 U18583 ( .A(n9569), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15157) );
  XNOR2_X1 U18584 ( .A(n15158), .B(n15157), .ZN(n15385) );
  NAND2_X1 U18585 ( .A1(n20526), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n15379) );
  OAI21_X1 U18586 ( .B1(n17161), .B2(n15159), .A(n15379), .ZN(n15162) );
  NOR2_X1 U18587 ( .A1(n15160), .A2(n20583), .ZN(n15161) );
  AOI211_X1 U18588 ( .C1(n15200), .C2(n15163), .A(n15162), .B(n15161), .ZN(
        n15164) );
  OAI21_X1 U18589 ( .B1(n15385), .B2(n20338), .A(n15164), .ZN(P1_U2976) );
  NAND2_X1 U18590 ( .A1(n15166), .A2(n15165), .ZN(n15167) );
  XOR2_X1 U18591 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n15167), .Z(
        n15392) );
  NAND2_X1 U18592 ( .A1(n20526), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n15386) );
  NAND2_X1 U18593 ( .A1(n20511), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15168) );
  OAI211_X1 U18594 ( .C1(n9869), .C2(n15169), .A(n15386), .B(n15168), .ZN(
        n15170) );
  AOI21_X1 U18595 ( .B1(n15171), .B2(n20518), .A(n15170), .ZN(n15172) );
  OAI21_X1 U18596 ( .B1(n20338), .B2(n15392), .A(n15172), .ZN(P1_U2977) );
  MUX2_X1 U18597 ( .A(n15174), .B(n15173), .S(n9569), .Z(n15176) );
  XNOR2_X1 U18598 ( .A(n15176), .B(n15175), .ZN(n15400) );
  NAND2_X1 U18599 ( .A1(n15200), .A2(n15177), .ZN(n15178) );
  NAND2_X1 U18600 ( .A1(n20526), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n15394) );
  OAI211_X1 U18601 ( .C1(n17161), .C2(n15179), .A(n15178), .B(n15394), .ZN(
        n15180) );
  AOI21_X1 U18602 ( .B1(n15181), .B2(n20518), .A(n15180), .ZN(n15182) );
  OAI21_X1 U18603 ( .B1(n20338), .B2(n15400), .A(n15182), .ZN(P1_U2978) );
  NAND2_X1 U18604 ( .A1(n13210), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15184) );
  MUX2_X1 U18605 ( .A(n15185), .B(n15184), .S(n9569), .Z(n15186) );
  XOR2_X1 U18606 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n15186), .Z(
        n15416) );
  NAND2_X1 U18607 ( .A1(n20526), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15408) );
  OAI21_X1 U18608 ( .B1(n17161), .B2(n15187), .A(n15408), .ZN(n15190) );
  NOR2_X1 U18609 ( .A1(n15188), .A2(n20583), .ZN(n15189) );
  AOI211_X1 U18610 ( .C1(n15200), .C2(n15191), .A(n15190), .B(n15189), .ZN(
        n15192) );
  OAI21_X1 U18611 ( .B1(n20338), .B2(n15416), .A(n15192), .ZN(P1_U2979) );
  NOR2_X1 U18612 ( .A1(n9569), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15193) );
  MUX2_X1 U18613 ( .A(n9569), .B(n15193), .S(n15183), .Z(n15194) );
  XNOR2_X1 U18614 ( .A(n15194), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15425) );
  NAND2_X1 U18615 ( .A1(n20526), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n15419) );
  OAI21_X1 U18616 ( .B1(n17161), .B2(n15195), .A(n15419), .ZN(n15198) );
  NOR2_X1 U18617 ( .A1(n15196), .A2(n20583), .ZN(n15197) );
  AOI211_X1 U18618 ( .C1(n15200), .C2(n15199), .A(n15198), .B(n15197), .ZN(
        n15201) );
  OAI21_X1 U18619 ( .B1(n20338), .B2(n15425), .A(n15201), .ZN(P1_U2980) );
  OAI21_X1 U18620 ( .B1(n15203), .B2(n15202), .A(n15183), .ZN(n15444) );
  INV_X1 U18621 ( .A(n15204), .ZN(n15208) );
  NAND2_X1 U18622 ( .A1(n20526), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n15436) );
  NAND2_X1 U18623 ( .A1(n20511), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15205) );
  OAI211_X1 U18624 ( .C1(n9869), .C2(n15206), .A(n15436), .B(n15205), .ZN(
        n15207) );
  AOI21_X1 U18625 ( .B1(n15208), .B2(n20518), .A(n15207), .ZN(n15209) );
  OAI21_X1 U18626 ( .B1(n20338), .B2(n15444), .A(n15209), .ZN(P1_U2981) );
  INV_X1 U18627 ( .A(n15212), .ZN(n15213) );
  INV_X1 U18628 ( .A(n15215), .ZN(n15216) );
  OR2_X1 U18629 ( .A1(n9569), .A2(n15216), .ZN(n15251) );
  AND2_X1 U18630 ( .A1(n10374), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15232) );
  NOR2_X1 U18631 ( .A1(n9569), .A2(n15217), .ZN(n15229) );
  NOR3_X1 U18632 ( .A1(n15249), .A2(n15232), .A3(n15229), .ZN(n15220) );
  INV_X1 U18633 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15219) );
  XNOR2_X1 U18634 ( .A(n9569), .B(n15219), .ZN(n15234) );
  NOR2_X1 U18635 ( .A1(n15222), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15221) );
  MUX2_X1 U18636 ( .A(n15222), .B(n15221), .S(n10374), .Z(n15223) );
  XNOR2_X1 U18637 ( .A(n15223), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15452) );
  NAND2_X1 U18638 ( .A1(n20526), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n15446) );
  NAND2_X1 U18639 ( .A1(n20511), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15224) );
  OAI211_X1 U18640 ( .C1(n9869), .C2(n15225), .A(n15446), .B(n15224), .ZN(
        n15226) );
  AOI21_X1 U18641 ( .B1(n15227), .B2(n20518), .A(n15226), .ZN(n15228) );
  OAI21_X1 U18642 ( .B1(n15452), .B2(n20338), .A(n15228), .ZN(P1_U2982) );
  INV_X1 U18643 ( .A(n15229), .ZN(n15230) );
  OAI211_X1 U18644 ( .C1(n15291), .C2(n15231), .A(n15251), .B(n15230), .ZN(
        n15243) );
  NOR2_X1 U18645 ( .A1(n15243), .A2(n15242), .ZN(n15241) );
  NOR2_X1 U18646 ( .A1(n15241), .A2(n15233), .ZN(n15235) );
  XNOR2_X1 U18647 ( .A(n15235), .B(n15234), .ZN(n15453) );
  NAND2_X1 U18648 ( .A1(n15453), .A2(n20519), .ZN(n15239) );
  AND2_X1 U18649 ( .A1(n20577), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n15457) );
  NOR2_X1 U18650 ( .A1(n9869), .A2(n15236), .ZN(n15237) );
  AOI211_X1 U18651 ( .C1(n20511), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n15457), .B(n15237), .ZN(n15238) );
  OAI211_X1 U18652 ( .C1(n20583), .C2(n15240), .A(n15239), .B(n15238), .ZN(
        P1_U2983) );
  AOI21_X1 U18653 ( .B1(n15243), .B2(n15242), .A(n15241), .ZN(n15468) );
  NAND2_X1 U18654 ( .A1(n20526), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n15461) );
  NAND2_X1 U18655 ( .A1(n20511), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15244) );
  OAI211_X1 U18656 ( .C1(n9869), .C2(n15245), .A(n15461), .B(n15244), .ZN(
        n15246) );
  AOI21_X1 U18657 ( .B1(n15247), .B2(n20518), .A(n15246), .ZN(n15248) );
  OAI21_X1 U18658 ( .B1(n15468), .B2(n20338), .A(n15248), .ZN(P1_U2984) );
  NAND2_X1 U18659 ( .A1(n15249), .A2(n15261), .ZN(n15250) );
  INV_X1 U18660 ( .A(n15264), .ZN(n15263) );
  INV_X1 U18661 ( .A(n15281), .ZN(n15290) );
  AOI21_X1 U18662 ( .B1(n15290), .B2(n15251), .A(n9569), .ZN(n15252) );
  NAND2_X1 U18663 ( .A1(n15469), .A2(n20519), .ZN(n15257) );
  NOR2_X1 U18664 ( .A1(n15267), .A2(n15253), .ZN(n15472) );
  NOR2_X1 U18665 ( .A1(n9869), .A2(n15254), .ZN(n15255) );
  AOI211_X1 U18666 ( .C1(n20511), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n15472), .B(n15255), .ZN(n15256) );
  OAI211_X1 U18667 ( .C1(n20583), .C2(n15258), .A(n15257), .B(n15256), .ZN(
        P1_U2985) );
  INV_X1 U18668 ( .A(n15291), .ZN(n15262) );
  INV_X1 U18669 ( .A(n15259), .ZN(n15260) );
  AOI22_X1 U18670 ( .A1(n15262), .A2(n15261), .B1(n10374), .B2(n15260), .ZN(
        n15275) );
  AOI21_X1 U18671 ( .B1(n10374), .B2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n15263), .ZN(n15274) );
  NAND2_X1 U18672 ( .A1(n15275), .A2(n15274), .ZN(n15273) );
  NAND2_X1 U18673 ( .A1(n15273), .A2(n15264), .ZN(n15266) );
  XNOR2_X1 U18674 ( .A(n9569), .B(n15482), .ZN(n15265) );
  XNOR2_X1 U18675 ( .A(n15266), .B(n15265), .ZN(n15487) );
  NOR2_X1 U18676 ( .A1(n15267), .A2(n21169), .ZN(n15479) );
  AOI21_X1 U18677 ( .B1(n20511), .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n15479), .ZN(n15268) );
  OAI21_X1 U18678 ( .B1(n15269), .B2(n9869), .A(n15268), .ZN(n15270) );
  AOI21_X1 U18679 ( .B1(n15271), .B2(n20518), .A(n15270), .ZN(n15272) );
  OAI21_X1 U18680 ( .B1(n15487), .B2(n20338), .A(n15272), .ZN(P1_U2986) );
  OAI21_X1 U18681 ( .B1(n15275), .B2(n15274), .A(n15273), .ZN(n15494) );
  NAND2_X1 U18682 ( .A1(n15494), .A2(n20519), .ZN(n15279) );
  AND2_X1 U18683 ( .A1(n20577), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n15498) );
  NOR2_X1 U18684 ( .A1(n9869), .A2(n15276), .ZN(n15277) );
  AOI211_X1 U18685 ( .C1(n20511), .C2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n15498), .B(n15277), .ZN(n15278) );
  OAI211_X1 U18686 ( .C1(n20583), .C2(n15280), .A(n15279), .B(n15278), .ZN(
        P1_U2987) );
  INV_X1 U18687 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15289) );
  NOR3_X1 U18688 ( .A1(n15291), .A2(n10374), .A3(n15289), .ZN(n15282) );
  NOR3_X1 U18689 ( .A1(n15281), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n9569), .ZN(n15294) );
  NOR2_X1 U18690 ( .A1(n15282), .A2(n15294), .ZN(n15283) );
  XNOR2_X1 U18691 ( .A(n15283), .B(n15493), .ZN(n15512) );
  NAND2_X1 U18692 ( .A1(n20526), .A2(P1_REIP_REG_11__SCAN_IN), .ZN(n15504) );
  NAND2_X1 U18693 ( .A1(n20511), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15284) );
  OAI211_X1 U18694 ( .C1(n9869), .C2(n15285), .A(n15504), .B(n15284), .ZN(
        n15286) );
  AOI21_X1 U18695 ( .B1(n15287), .B2(n20518), .A(n15286), .ZN(n15288) );
  OAI21_X1 U18696 ( .B1(n15512), .B2(n20338), .A(n15288), .ZN(P1_U2988) );
  NOR2_X1 U18697 ( .A1(n15290), .A2(n15289), .ZN(n15293) );
  XNOR2_X1 U18698 ( .A(n15291), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15292) );
  MUX2_X1 U18699 ( .A(n15293), .B(n15292), .S(n9569), .Z(n15295) );
  NOR2_X1 U18700 ( .A1(n15295), .A2(n15294), .ZN(n15529) );
  NAND2_X1 U18701 ( .A1(n20526), .A2(P1_REIP_REG_10__SCAN_IN), .ZN(n15524) );
  NAND2_X1 U18702 ( .A1(n20511), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15296) );
  OAI211_X1 U18703 ( .C1(n9869), .C2(n15297), .A(n15524), .B(n15296), .ZN(
        n15298) );
  AOI21_X1 U18704 ( .B1(n15299), .B2(n20518), .A(n15298), .ZN(n15300) );
  OAI21_X1 U18705 ( .B1(n15529), .B2(n20338), .A(n15300), .ZN(P1_U2989) );
  XNOR2_X1 U18706 ( .A(n9569), .B(n15530), .ZN(n15301) );
  XNOR2_X1 U18707 ( .A(n15302), .B(n15301), .ZN(n15537) );
  NAND2_X1 U18708 ( .A1(n20511), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15303) );
  NAND2_X1 U18709 ( .A1(n20526), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n15532) );
  OAI211_X1 U18710 ( .C1(n9869), .C2(n20359), .A(n15303), .B(n15532), .ZN(
        n15304) );
  AOI21_X1 U18711 ( .B1(n20361), .B2(n20518), .A(n15304), .ZN(n15305) );
  OAI21_X1 U18712 ( .B1(n15537), .B2(n20338), .A(n15305), .ZN(P1_U2990) );
  XOR2_X1 U18713 ( .A(n15307), .B(n15306), .Z(n15550) );
  INV_X1 U18714 ( .A(n15308), .ZN(n20441) );
  NAND2_X1 U18715 ( .A1(n20511), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15309) );
  NAND2_X1 U18716 ( .A1(n20526), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n15547) );
  OAI211_X1 U18717 ( .C1(n9869), .C2(n20369), .A(n15309), .B(n15547), .ZN(
        n15310) );
  AOI21_X1 U18718 ( .B1(n20441), .B2(n20518), .A(n15310), .ZN(n15311) );
  OAI21_X1 U18719 ( .B1(n15550), .B2(n20338), .A(n15311), .ZN(P1_U2991) );
  INV_X1 U18720 ( .A(n15312), .ZN(n15313) );
  NAND2_X1 U18721 ( .A1(n15313), .A2(n20518), .ZN(n15318) );
  OR2_X1 U18722 ( .A1(n15314), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20564) );
  NAND3_X1 U18723 ( .A1(n20564), .A2(n15315), .A3(n20519), .ZN(n15317) );
  MUX2_X1 U18724 ( .A(n9869), .B(n17161), .S(P1_PHYADDRPOINTER_REG_1__SCAN_IN), 
        .Z(n15316) );
  NAND2_X1 U18725 ( .A1(n20526), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20557) );
  NAND4_X1 U18726 ( .A1(n15318), .A2(n15317), .A3(n15316), .A4(n20557), .ZN(
        P1_U2998) );
  OAI21_X1 U18727 ( .B1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15320), .A(
        n15319), .ZN(n15321) );
  NAND3_X1 U18728 ( .A1(n10022), .A2(n10381), .A3(n15328), .ZN(n15326) );
  OAI211_X1 U18729 ( .C1(n15329), .C2(n15328), .A(n15327), .B(n15326), .ZN(
        n15330) );
  AOI21_X1 U18730 ( .B1(n15331), .B2(n20560), .A(n15330), .ZN(n15332) );
  OAI21_X1 U18731 ( .B1(n15333), .B2(n20573), .A(n15332), .ZN(P1_U3002) );
  INV_X1 U18732 ( .A(n15334), .ZN(n15337) );
  AOI211_X1 U18733 ( .C1(n15345), .C2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15337), .B(n15336), .ZN(n15340) );
  NAND2_X1 U18734 ( .A1(n15338), .A2(n20560), .ZN(n15339) );
  OAI211_X1 U18735 ( .C1(n15341), .C2(n20573), .A(n15340), .B(n15339), .ZN(
        P1_U3003) );
  NOR2_X1 U18736 ( .A1(n15342), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15343) );
  AOI211_X1 U18737 ( .C1(n15345), .C2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15344), .B(n15343), .ZN(n15349) );
  INV_X1 U18738 ( .A(n15346), .ZN(n15347) );
  NAND2_X1 U18739 ( .A1(n15347), .A2(n20560), .ZN(n15348) );
  OAI211_X1 U18740 ( .C1(n15350), .C2(n20573), .A(n15349), .B(n15348), .ZN(
        P1_U3004) );
  INV_X1 U18741 ( .A(n15362), .ZN(n15351) );
  AOI21_X1 U18742 ( .B1(n15351), .B2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15353) );
  OAI21_X1 U18743 ( .B1(n15354), .B2(n15353), .A(n15352), .ZN(n15355) );
  AOI21_X1 U18744 ( .B1(n15356), .B2(n20560), .A(n15355), .ZN(n15357) );
  OAI21_X1 U18745 ( .B1(n15358), .B2(n20573), .A(n15357), .ZN(P1_U3005) );
  OAI21_X1 U18746 ( .B1(n15378), .B2(n15359), .A(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15361) );
  OAI211_X1 U18747 ( .C1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n15362), .A(
        n15361), .B(n15360), .ZN(n15363) );
  AOI21_X1 U18748 ( .B1(n15364), .B2(n20560), .A(n15363), .ZN(n15365) );
  OAI21_X1 U18749 ( .B1(n15366), .B2(n20573), .A(n15365), .ZN(P1_U3006) );
  INV_X1 U18750 ( .A(n20549), .ZN(n15367) );
  AOI21_X1 U18751 ( .B1(n15515), .B2(n15367), .A(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15368) );
  OAI21_X1 U18752 ( .B1(n15378), .B2(n15368), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15372) );
  INV_X1 U18753 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15369) );
  NAND3_X1 U18754 ( .A1(n15377), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n15369), .ZN(n15370) );
  NAND3_X1 U18755 ( .A1(n15372), .A2(n15371), .A3(n15370), .ZN(n15373) );
  AOI21_X1 U18756 ( .B1(n15374), .B2(n20560), .A(n15373), .ZN(n15375) );
  OAI21_X1 U18757 ( .B1(n15376), .B2(n20573), .A(n15375), .ZN(P1_U3007) );
  INV_X1 U18758 ( .A(n15377), .ZN(n15381) );
  NAND2_X1 U18759 ( .A1(n15378), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15380) );
  OAI211_X1 U18760 ( .C1(n15381), .C2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15380), .B(n15379), .ZN(n15382) );
  AOI21_X1 U18761 ( .B1(n15383), .B2(n20560), .A(n15382), .ZN(n15384) );
  OAI21_X1 U18762 ( .B1(n15385), .B2(n20573), .A(n15384), .ZN(P1_U3008) );
  XNOR2_X1 U18763 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15387) );
  OAI21_X1 U18764 ( .B1(n15396), .B2(n15387), .A(n15386), .ZN(n15390) );
  NOR2_X1 U18765 ( .A1(n15388), .A2(n20575), .ZN(n15389) );
  AOI211_X1 U18766 ( .C1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n15393), .A(
        n15390), .B(n15389), .ZN(n15391) );
  OAI21_X1 U18767 ( .B1(n15392), .B2(n20573), .A(n15391), .ZN(P1_U3009) );
  NAND2_X1 U18768 ( .A1(n15393), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15395) );
  OAI211_X1 U18769 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n15396), .A(
        n15395), .B(n15394), .ZN(n15397) );
  AOI21_X1 U18770 ( .B1(n15398), .B2(n20560), .A(n15397), .ZN(n15399) );
  OAI21_X1 U18771 ( .B1(n15400), .B2(n20573), .A(n15399), .ZN(P1_U3010) );
  NOR3_X1 U18772 ( .A1(n20555), .A2(n15401), .A3(n15478), .ZN(n15402) );
  AOI21_X1 U18773 ( .B1(n20570), .B2(n15403), .A(n15402), .ZN(n15477) );
  INV_X1 U18774 ( .A(n20545), .ZN(n15518) );
  OAI21_X1 U18775 ( .B1(n15409), .B2(n15404), .A(n15518), .ZN(n15405) );
  OAI211_X1 U18776 ( .C1(n15406), .C2(n15515), .A(n20544), .B(n15405), .ZN(
        n15418) );
  INV_X1 U18777 ( .A(n15418), .ZN(n15407) );
  OAI21_X1 U18778 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n15477), .A(
        n15407), .ZN(n15412) );
  INV_X1 U18779 ( .A(n15408), .ZN(n15411) );
  NOR3_X1 U18780 ( .A1(n15421), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n15409), .ZN(n15410) );
  AOI211_X1 U18781 ( .C1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n15412), .A(
        n15411), .B(n15410), .ZN(n15415) );
  NAND2_X1 U18782 ( .A1(n15413), .A2(n20560), .ZN(n15414) );
  OAI211_X1 U18783 ( .C1(n15416), .C2(n20573), .A(n15415), .B(n15414), .ZN(
        P1_U3011) );
  INV_X1 U18784 ( .A(n15417), .ZN(n15423) );
  NAND2_X1 U18785 ( .A1(n15418), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15420) );
  OAI211_X1 U18786 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15421), .A(
        n15420), .B(n15419), .ZN(n15422) );
  AOI21_X1 U18787 ( .B1(n15423), .B2(n20560), .A(n15422), .ZN(n15424) );
  OAI21_X1 U18788 ( .B1(n15425), .B2(n20573), .A(n15424), .ZN(P1_U3012) );
  OR2_X1 U18789 ( .A1(n20562), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15432) );
  OR2_X1 U18790 ( .A1(n20545), .A2(n15426), .ZN(n15431) );
  INV_X1 U18791 ( .A(n15427), .ZN(n15428) );
  AND2_X1 U18792 ( .A1(n20570), .A2(n15428), .ZN(n15429) );
  NOR2_X1 U18793 ( .A1(n20554), .A2(n15429), .ZN(n15430) );
  NAND2_X1 U18794 ( .A1(n15432), .A2(n15483), .ZN(n15466) );
  NOR2_X1 U18795 ( .A1(n20562), .A2(n15435), .ZN(n15433) );
  NOR2_X1 U18796 ( .A1(n15466), .A2(n15433), .ZN(n15448) );
  INV_X1 U18797 ( .A(n15448), .ZN(n15439) );
  INV_X1 U18798 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15434) );
  NAND2_X1 U18799 ( .A1(n15435), .A2(n15434), .ZN(n15437) );
  OAI21_X1 U18800 ( .B1(n15462), .B2(n15437), .A(n15436), .ZN(n15438) );
  AOI21_X1 U18801 ( .B1(n15439), .B2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15438), .ZN(n15443) );
  INV_X1 U18802 ( .A(n15440), .ZN(n15441) );
  NAND2_X1 U18803 ( .A1(n15441), .A2(n20560), .ZN(n15442) );
  OAI211_X1 U18804 ( .C1(n15444), .C2(n20573), .A(n15443), .B(n15442), .ZN(
        P1_U3013) );
  INV_X1 U18805 ( .A(n15462), .ZN(n15445) );
  AOI21_X1 U18806 ( .B1(n15445), .B2(n15454), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15447) );
  OAI21_X1 U18807 ( .B1(n15448), .B2(n15447), .A(n15446), .ZN(n15449) );
  AOI21_X1 U18808 ( .B1(n15450), .B2(n20560), .A(n15449), .ZN(n15451) );
  OAI21_X1 U18809 ( .B1(n15452), .B2(n20573), .A(n15451), .ZN(P1_U3014) );
  NAND2_X1 U18810 ( .A1(n15453), .A2(n20563), .ZN(n15459) );
  NOR3_X1 U18811 ( .A1(n15462), .A2(n15455), .A3(n15454), .ZN(n15456) );
  AOI211_X1 U18812 ( .C1(n15466), .C2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n15457), .B(n15456), .ZN(n15458) );
  OAI211_X1 U18813 ( .C1(n20575), .C2(n15460), .A(n15459), .B(n15458), .ZN(
        P1_U3015) );
  OAI21_X1 U18814 ( .B1(n15462), .B2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15461), .ZN(n15465) );
  NOR2_X1 U18815 ( .A1(n15463), .A2(n20575), .ZN(n15464) );
  AOI211_X1 U18816 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n15466), .A(
        n15465), .B(n15464), .ZN(n15467) );
  OAI21_X1 U18817 ( .B1(n15468), .B2(n20573), .A(n15467), .ZN(P1_U3016) );
  INV_X1 U18818 ( .A(n15483), .ZN(n15473) );
  INV_X1 U18819 ( .A(n15541), .ZN(n17171) );
  NOR4_X1 U18820 ( .A1(n17171), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n15482), .A4(n15470), .ZN(n15471) );
  AOI211_X1 U18821 ( .C1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n15473), .A(
        n15472), .B(n15471), .ZN(n15474) );
  OAI211_X1 U18822 ( .C1(n20575), .C2(n15476), .A(n15475), .B(n15474), .ZN(
        P1_U3017) );
  OAI21_X1 U18823 ( .B1(n20579), .B2(n15478), .A(n15477), .ZN(n15480) );
  AOI21_X1 U18824 ( .B1(n15480), .B2(n15482), .A(n15479), .ZN(n15481) );
  OAI21_X1 U18825 ( .B1(n15483), .B2(n15482), .A(n15481), .ZN(n15484) );
  AOI21_X1 U18826 ( .B1(n15485), .B2(n20560), .A(n15484), .ZN(n15486) );
  OAI21_X1 U18827 ( .B1(n15487), .B2(n20573), .A(n15486), .ZN(P1_U3018) );
  INV_X1 U18828 ( .A(n15488), .ZN(n15489) );
  OAI21_X1 U18829 ( .B1(n15490), .B2(n15489), .A(n15518), .ZN(n15492) );
  OAI211_X1 U18830 ( .C1(n15495), .C2(n15515), .A(n15492), .B(n15491), .ZN(
        n15510) );
  AOI21_X1 U18831 ( .B1(n20549), .B2(n15493), .A(n15510), .ZN(n15503) );
  NAND2_X1 U18832 ( .A1(n15494), .A2(n20563), .ZN(n15501) );
  INV_X1 U18833 ( .A(n15495), .ZN(n15496) );
  NOR3_X1 U18834 ( .A1(n17171), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        n15496), .ZN(n15497) );
  AOI211_X1 U18835 ( .C1(n20560), .C2(n15499), .A(n15498), .B(n15497), .ZN(
        n15500) );
  OAI211_X1 U18836 ( .C1(n15503), .C2(n15502), .A(n15501), .B(n15500), .ZN(
        P1_U3019) );
  OAI21_X1 U18837 ( .B1(n15505), .B2(n20575), .A(n15504), .ZN(n15509) );
  NOR2_X1 U18838 ( .A1(n17171), .A2(n15521), .ZN(n15531) );
  INV_X1 U18839 ( .A(n15531), .ZN(n15507) );
  NOR3_X1 U18840 ( .A1(n15507), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        n15506), .ZN(n15508) );
  AOI211_X1 U18841 ( .C1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n15510), .A(
        n15509), .B(n15508), .ZN(n15511) );
  OAI21_X1 U18842 ( .B1(n15512), .B2(n20573), .A(n15511), .ZN(P1_U3020) );
  INV_X1 U18843 ( .A(n15513), .ZN(n15517) );
  OR2_X1 U18844 ( .A1(n15515), .A2(n15514), .ZN(n20551) );
  INV_X1 U18845 ( .A(n20551), .ZN(n15516) );
  AOI211_X1 U18846 ( .C1(n15518), .C2(n15517), .A(n20554), .B(n15516), .ZN(
        n20528) );
  OAI21_X1 U18847 ( .B1(n15521), .B2(n15520), .A(n15519), .ZN(n15522) );
  NAND2_X1 U18848 ( .A1(n20528), .A2(n15522), .ZN(n15535) );
  XNOR2_X1 U18849 ( .A(n15530), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15523) );
  NAND2_X1 U18850 ( .A1(n15531), .A2(n15523), .ZN(n15525) );
  OAI211_X1 U18851 ( .C1(n20575), .C2(n15526), .A(n15525), .B(n15524), .ZN(
        n15527) );
  AOI21_X1 U18852 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n15535), .A(
        n15527), .ZN(n15528) );
  OAI21_X1 U18853 ( .B1(n15529), .B2(n20573), .A(n15528), .ZN(P1_U3021) );
  NAND2_X1 U18854 ( .A1(n15531), .A2(n15530), .ZN(n15533) );
  OAI211_X1 U18855 ( .C1(n20575), .C2(n20357), .A(n15533), .B(n15532), .ZN(
        n15534) );
  AOI21_X1 U18856 ( .B1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15535), .A(
        n15534), .ZN(n15536) );
  OAI21_X1 U18857 ( .B1(n15537), .B2(n20573), .A(n15536), .ZN(P1_U3022) );
  INV_X1 U18858 ( .A(n15003), .ZN(n15538) );
  AOI21_X1 U18859 ( .B1(n15540), .B2(n15539), .A(n15538), .ZN(n20438) );
  OAI211_X1 U18860 ( .C1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n15541), .ZN(n15542) );
  INV_X1 U18861 ( .A(n15542), .ZN(n15544) );
  AOI22_X1 U18862 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n15545), .B1(
        n15544), .B2(n15543), .ZN(n15546) );
  NAND2_X1 U18863 ( .A1(n15547), .A2(n15546), .ZN(n15548) );
  AOI21_X1 U18864 ( .B1(n20438), .B2(n20560), .A(n15548), .ZN(n15549) );
  OAI21_X1 U18865 ( .B1(n15550), .B2(n20573), .A(n15549), .ZN(P1_U3023) );
  NAND2_X1 U18866 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20963), .ZN(n21385) );
  INV_X1 U18867 ( .A(n21385), .ZN(n15577) );
  NAND2_X1 U18868 ( .A1(n21383), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n15551) );
  OR2_X1 U18869 ( .A1(n20662), .A2(n15551), .ZN(n20869) );
  NAND3_X1 U18870 ( .A1(n20662), .A2(n21383), .A3(n21022), .ZN(n15552) );
  OAI211_X1 U18871 ( .C1(n14960), .C2(n15577), .A(n20869), .B(n15552), .ZN(
        n15568) );
  NOR2_X1 U18872 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n13636), .ZN(n15555) );
  MUX2_X1 U18873 ( .A(n15553), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n17117), .Z(n17126) );
  AOI22_X1 U18874 ( .A1(n15555), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n13636), .B2(n17126), .ZN(n15557) );
  MUX2_X1 U18875 ( .A(n15554), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n17117), .Z(n17120) );
  AOI22_X1 U18876 ( .A1(n17120), .A2(n13636), .B1(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n15555), .ZN(n15556) );
  INV_X1 U18877 ( .A(n17129), .ZN(n15558) );
  INV_X1 U18878 ( .A(n12276), .ZN(n15581) );
  NAND2_X1 U18879 ( .A1(n15558), .A2(n15581), .ZN(n17142) );
  AOI21_X1 U18880 ( .B1(n17117), .B2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n15560) );
  NAND2_X1 U18881 ( .A1(n15560), .A2(n15559), .ZN(n15562) );
  NAND2_X1 U18882 ( .A1(n12693), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n15561) );
  NOR2_X1 U18883 ( .A1(n17130), .A2(P1_FLUSH_REG_SCAN_IN), .ZN(n15563) );
  NAND2_X1 U18884 ( .A1(n17142), .A2(n15563), .ZN(n15565) );
  INV_X1 U18885 ( .A(n17189), .ZN(n15564) );
  NAND2_X1 U18886 ( .A1(n15565), .A2(n15564), .ZN(n15567) );
  MUX2_X1 U18887 ( .A(n15568), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        n21382), .Z(P1_U3477) );
  AND2_X1 U18888 ( .A1(n20662), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n15569) );
  NAND2_X1 U18889 ( .A1(n15569), .A2(n21383), .ZN(n20933) );
  INV_X1 U18890 ( .A(n15569), .ZN(n15573) );
  NAND2_X1 U18891 ( .A1(n15573), .A2(n21383), .ZN(n21074) );
  MUX2_X1 U18892 ( .A(n20933), .B(n21074), .S(n20585), .Z(n15570) );
  OAI21_X1 U18893 ( .B1(n15577), .B2(n13947), .A(n15570), .ZN(n15571) );
  MUX2_X1 U18894 ( .A(n15571), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        n21382), .Z(P1_U3476) );
  AOI21_X1 U18895 ( .B1(n20934), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20586), 
        .ZN(n15574) );
  NOR2_X1 U18896 ( .A1(n20807), .A2(n15573), .ZN(n20811) );
  NOR2_X1 U18897 ( .A1(n15574), .A2(n20811), .ZN(n15575) );
  OAI222_X1 U18898 ( .A1(n21017), .A2(n20869), .B1(n15577), .B2(n15576), .C1(
        n21075), .C2(n15575), .ZN(n15578) );
  MUX2_X1 U18899 ( .A(n15578), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        n21382), .Z(P1_U3475) );
  INV_X1 U18900 ( .A(n15579), .ZN(n15583) );
  INV_X1 U18901 ( .A(n13949), .ZN(n15580) );
  NAND2_X1 U18902 ( .A1(n15581), .A2(n15580), .ZN(n15587) );
  OAI22_X1 U18903 ( .A1(n15583), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n15587), .B2(n15582), .ZN(n15584) );
  AOI21_X1 U18904 ( .B1(n10366), .B2(n15585), .A(n15584), .ZN(n17116) );
  INV_X1 U18905 ( .A(n15586), .ZN(n20333) );
  INV_X1 U18906 ( .A(n15587), .ZN(n15590) );
  AOI22_X1 U18907 ( .A1(n15591), .A2(n15590), .B1(n15589), .B2(n15588), .ZN(
        n15592) );
  OAI21_X1 U18908 ( .B1(n17116), .B2(n20333), .A(n15592), .ZN(n15594) );
  MUX2_X1 U18909 ( .A(n15594), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n15593), .Z(P1_U3473) );
  NOR2_X1 U18910 ( .A1(n15596), .A2(n15595), .ZN(n15597) );
  INV_X1 U18911 ( .A(n15599), .ZN(n16432) );
  NAND2_X1 U18912 ( .A1(n16432), .A2(n19413), .ZN(n15608) );
  XNOR2_X1 U18913 ( .A(n15601), .B(n15600), .ZN(n15604) );
  AOI22_X1 U18914 ( .A1(n19403), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n19410), .ZN(n15603) );
  NAND2_X1 U18915 ( .A1(n19404), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15602) );
  OAI211_X1 U18916 ( .C1(n15604), .C2(n19417), .A(n15603), .B(n15602), .ZN(
        n15605) );
  AOI21_X1 U18917 ( .B1(n15606), .B2(n15968), .A(n15605), .ZN(n15607) );
  OAI211_X1 U18918 ( .C1(n19407), .C2(n16430), .A(n15608), .B(n15607), .ZN(
        P2_U2826) );
  AOI21_X1 U18919 ( .B1(n15612), .B2(n15942), .A(n19400), .ZN(n15616) );
  NAND2_X1 U18920 ( .A1(n15609), .A2(n15968), .ZN(n15614) );
  INV_X1 U18921 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n15610) );
  OAI22_X1 U18922 ( .A1(n19392), .A2(n15610), .B1(n20254), .B2(n15958), .ZN(
        n15613) );
  INV_X1 U18923 ( .A(n15615), .ZN(n15611) );
  NAND2_X1 U18924 ( .A1(n15617), .A2(n15618), .ZN(n15619) );
  NAND2_X1 U18925 ( .A1(n15620), .A2(n15619), .ZN(n16446) );
  AOI21_X1 U18926 ( .B1(n15622), .B2(n15621), .A(n11421), .ZN(n16437) );
  NAND2_X1 U18927 ( .A1(n16437), .A2(n19413), .ZN(n15631) );
  XOR2_X1 U18928 ( .A(n16210), .B(n15623), .Z(n15629) );
  AOI22_X1 U18929 ( .A1(n19403), .A2(P2_EBX_REG_27__SCAN_IN), .B1(
        P2_REIP_REG_27__SCAN_IN), .B2(n19410), .ZN(n15624) );
  OAI21_X1 U18930 ( .B1(n15625), .B2(n19389), .A(n15624), .ZN(n15628) );
  NOR2_X1 U18931 ( .A1(n15626), .A2(n19405), .ZN(n15627) );
  AOI211_X1 U18932 ( .C1(n15942), .C2(n15629), .A(n15628), .B(n15627), .ZN(
        n15630) );
  OAI211_X1 U18933 ( .C1(n19407), .C2(n16446), .A(n15631), .B(n15630), .ZN(
        P2_U2828) );
  OAI21_X1 U18934 ( .B1(n15632), .B2(n15633), .A(n15621), .ZN(n16460) );
  OR2_X1 U18935 ( .A1(n15634), .A2(n15635), .ZN(n15636) );
  AND2_X1 U18936 ( .A1(n15617), .A2(n15636), .ZN(n16458) );
  OAI21_X1 U18937 ( .B1(n15637), .B2(n19417), .A(n15957), .ZN(n15641) );
  NAND3_X1 U18938 ( .A1(n15637), .A2(n15967), .A3(n13475), .ZN(n15639) );
  AOI22_X1 U18939 ( .A1(n19403), .A2(P2_EBX_REG_26__SCAN_IN), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n19410), .ZN(n15638) );
  OAI211_X1 U18940 ( .C1(n19389), .C2(n16218), .A(n15639), .B(n15638), .ZN(
        n15640) );
  AOI21_X1 U18941 ( .B1(n16220), .B2(n15641), .A(n15640), .ZN(n15642) );
  OAI21_X1 U18942 ( .B1(n15643), .B2(n19405), .A(n15642), .ZN(n15644) );
  AOI21_X1 U18943 ( .B1(n16458), .B2(n19384), .A(n15644), .ZN(n15645) );
  OAI21_X1 U18944 ( .B1(n16460), .B2(n15911), .A(n15645), .ZN(P2_U2829) );
  INV_X1 U18945 ( .A(n15634), .ZN(n15647) );
  OAI21_X1 U18946 ( .B1(n15646), .B2(n15648), .A(n15647), .ZN(n16470) );
  INV_X1 U18947 ( .A(n15649), .ZN(n15650) );
  AOI21_X1 U18948 ( .B1(n15651), .B2(n15650), .A(n15632), .ZN(n16473) );
  NAND2_X1 U18949 ( .A1(n16473), .A2(n19413), .ZN(n15660) );
  XOR2_X1 U18950 ( .A(n16228), .B(n15652), .Z(n15658) );
  AOI22_X1 U18951 ( .A1(n19403), .A2(P2_EBX_REG_25__SCAN_IN), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n19410), .ZN(n15653) );
  OAI21_X1 U18952 ( .B1(n15654), .B2(n19389), .A(n15653), .ZN(n15657) );
  NOR2_X1 U18953 ( .A1(n15655), .A2(n19405), .ZN(n15656) );
  AOI211_X1 U18954 ( .C1(n15942), .C2(n15658), .A(n15657), .B(n15656), .ZN(
        n15659) );
  OAI211_X1 U18955 ( .C1(n19407), .C2(n16470), .A(n15660), .B(n15659), .ZN(
        P2_U2830) );
  NAND2_X1 U18956 ( .A1(n15676), .A2(n15661), .ZN(n15662) );
  NAND2_X1 U18957 ( .A1(n15650), .A2(n15662), .ZN(n16487) );
  AOI21_X1 U18958 ( .B1(n15664), .B2(n15663), .A(n15646), .ZN(n16479) );
  OAI22_X1 U18959 ( .A1(n19392), .A2(n16010), .B1(n20248), .B2(n15958), .ZN(
        n15667) );
  NOR3_X1 U18960 ( .A1(n15665), .A2(n16239), .A3(n19386), .ZN(n15666) );
  AOI211_X1 U18961 ( .C1(n19404), .C2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15667), .B(n15666), .ZN(n15671) );
  OAI21_X1 U18962 ( .B1(n15668), .B2(n19417), .A(n15957), .ZN(n15669) );
  NAND2_X1 U18963 ( .A1(n15669), .A2(n16239), .ZN(n15670) );
  OAI211_X1 U18964 ( .C1(n15672), .C2(n19405), .A(n15671), .B(n15670), .ZN(
        n15673) );
  AOI21_X1 U18965 ( .B1(n16479), .B2(n19384), .A(n15673), .ZN(n15674) );
  OAI21_X1 U18966 ( .B1(n16487), .B2(n15911), .A(n15674), .ZN(P2_U2831) );
  OAI21_X1 U18967 ( .B1(n9667), .B2(n11371), .A(n15676), .ZN(n16495) );
  XNOR2_X1 U18968 ( .A(n15677), .B(n16245), .ZN(n15680) );
  AOI22_X1 U18969 ( .A1(n19403), .A2(P2_EBX_REG_23__SCAN_IN), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n19410), .ZN(n15679) );
  NAND2_X1 U18970 ( .A1(n19404), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15678) );
  OAI211_X1 U18971 ( .C1(n15680), .C2(n19417), .A(n15679), .B(n15678), .ZN(
        n15681) );
  AOI21_X1 U18972 ( .B1(n15682), .B2(n15968), .A(n15681), .ZN(n15687) );
  INV_X1 U18973 ( .A(n15663), .ZN(n15684) );
  AOI21_X1 U18974 ( .B1(n15685), .B2(n15694), .A(n15684), .ZN(n16498) );
  NAND2_X1 U18975 ( .A1(n16498), .A2(n19384), .ZN(n15686) );
  OAI211_X1 U18976 ( .C1(n16495), .C2(n15911), .A(n15687), .B(n15686), .ZN(
        P2_U2832) );
  INV_X1 U18977 ( .A(n15688), .ZN(n15689) );
  AOI21_X1 U18978 ( .B1(n15689), .B2(n9634), .A(n9667), .ZN(n16511) );
  INV_X1 U18979 ( .A(n16511), .ZN(n16021) );
  OR2_X1 U18980 ( .A1(n15691), .A2(n15692), .ZN(n15693) );
  NAND2_X1 U18981 ( .A1(n15694), .A2(n15693), .ZN(n16509) );
  INV_X1 U18982 ( .A(n16509), .ZN(n16144) );
  NOR2_X1 U18983 ( .A1(n15695), .A2(n19405), .ZN(n15704) );
  AOI21_X1 U18984 ( .B1(n15698), .B2(n15942), .A(n19400), .ZN(n15702) );
  INV_X1 U18985 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n20245) );
  OAI22_X1 U18986 ( .A1(n19392), .A2(n15696), .B1(n20245), .B2(n15958), .ZN(
        n15700) );
  INV_X1 U18987 ( .A(n16260), .ZN(n15697) );
  NOR3_X1 U18988 ( .A1(n15698), .A2(n19386), .A3(n15697), .ZN(n15699) );
  AOI211_X1 U18989 ( .C1(n19404), .C2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15700), .B(n15699), .ZN(n15701) );
  OAI21_X1 U18990 ( .B1(n16260), .B2(n15702), .A(n15701), .ZN(n15703) );
  AOI211_X1 U18991 ( .C1(n16144), .C2(n19384), .A(n15704), .B(n15703), .ZN(
        n15705) );
  OAI21_X1 U18992 ( .B1(n16021), .B2(n15911), .A(n15705), .ZN(P2_U2833) );
  OAI21_X1 U18993 ( .B1(n11469), .B2(n15706), .A(n9634), .ZN(n16528) );
  INV_X1 U18994 ( .A(n15707), .ZN(n15709) );
  INV_X1 U18995 ( .A(n15708), .ZN(n15720) );
  AOI21_X1 U18996 ( .B1(n15709), .B2(n15720), .A(n15691), .ZN(n16526) );
  INV_X1 U18997 ( .A(n15710), .ZN(n15717) );
  OAI21_X1 U18998 ( .B1(n15722), .B2(n19417), .A(n15957), .ZN(n15715) );
  INV_X1 U18999 ( .A(n16276), .ZN(n15711) );
  NAND3_X1 U19000 ( .A1(n15722), .A2(n15967), .A3(n15711), .ZN(n15713) );
  AOI22_X1 U19001 ( .A1(n19403), .A2(P2_EBX_REG_21__SCAN_IN), .B1(
        P2_REIP_REG_21__SCAN_IN), .B2(n19410), .ZN(n15712) );
  OAI211_X1 U19002 ( .C1(n19389), .C2(n16274), .A(n15713), .B(n15712), .ZN(
        n15714) );
  AOI21_X1 U19003 ( .B1(n16276), .B2(n15715), .A(n15714), .ZN(n15716) );
  OAI21_X1 U19004 ( .B1(n15717), .B2(n19405), .A(n15716), .ZN(n15718) );
  AOI21_X1 U19005 ( .B1(n16526), .B2(n19384), .A(n15718), .ZN(n15719) );
  OAI21_X1 U19006 ( .B1(n16528), .B2(n15911), .A(n15719), .ZN(P2_U2834) );
  OAI21_X1 U19007 ( .B1(n9698), .B2(n15721), .A(n15720), .ZN(n16541) );
  NAND2_X1 U19008 ( .A1(n16533), .A2(n19413), .ZN(n15733) );
  OAI21_X1 U19009 ( .B1(n15723), .B2(n15725), .A(n15722), .ZN(n15724) );
  NOR2_X1 U19010 ( .A1(n15724), .A2(n19386), .ZN(n15730) );
  INV_X1 U19011 ( .A(n15725), .ZN(n15726) );
  AOI22_X1 U19012 ( .A1(n19410), .A2(P2_REIP_REG_20__SCAN_IN), .B1(n19400), 
        .B2(n15726), .ZN(n15728) );
  NAND2_X1 U19013 ( .A1(n19403), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n15727) );
  OAI211_X1 U19014 ( .C1(n19389), .C2(n10119), .A(n15728), .B(n15727), .ZN(
        n15729) );
  AOI211_X1 U19015 ( .C1(n15731), .C2(n15968), .A(n15730), .B(n15729), .ZN(
        n15732) );
  OAI211_X1 U19016 ( .C1(n19407), .C2(n16541), .A(n15733), .B(n15732), .ZN(
        P2_U2835) );
  INV_X1 U19017 ( .A(n15734), .ZN(n16172) );
  INV_X1 U19018 ( .A(n16032), .ZN(n15747) );
  OAI21_X1 U19019 ( .B1(n15741), .B2(n19417), .A(n15957), .ZN(n15739) );
  OAI21_X1 U19020 ( .B1(n15958), .B2(n20239), .A(n17200), .ZN(n15735) );
  AOI21_X1 U19021 ( .B1(n19403), .B2(P2_EBX_REG_19__SCAN_IN), .A(n15735), .ZN(
        n15736) );
  OAI21_X1 U19022 ( .B1(n15737), .B2(n19389), .A(n15736), .ZN(n15738) );
  AOI21_X1 U19023 ( .B1(n15740), .B2(n15739), .A(n15738), .ZN(n15744) );
  INV_X1 U19024 ( .A(n15740), .ZN(n15742) );
  NAND3_X1 U19025 ( .A1(n15742), .A2(n15967), .A3(n15741), .ZN(n15743) );
  OAI211_X1 U19026 ( .C1(n15745), .C2(n19405), .A(n15744), .B(n15743), .ZN(
        n15746) );
  AOI21_X1 U19027 ( .B1(n15747), .B2(n19413), .A(n15746), .ZN(n15748) );
  OAI21_X1 U19028 ( .B1(n16172), .B2(n19407), .A(n15748), .ZN(P2_U2836) );
  OAI21_X1 U19029 ( .B1(n11501), .B2(n15749), .A(n11543), .ZN(n16553) );
  NOR3_X1 U19030 ( .A1(n10192), .A2(n15750), .A3(n19386), .ZN(n15757) );
  OAI21_X1 U19031 ( .B1(n19417), .B2(n10193), .A(n15957), .ZN(n15751) );
  INV_X1 U19032 ( .A(n15751), .ZN(n15755) );
  INV_X1 U19033 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n20237) );
  OAI21_X1 U19034 ( .B1(n15958), .B2(n20237), .A(n17200), .ZN(n15752) );
  AOI21_X1 U19035 ( .B1(n19403), .B2(P2_EBX_REG_18__SCAN_IN), .A(n15752), .ZN(
        n15754) );
  NAND2_X1 U19036 ( .A1(n19404), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15753) );
  OAI211_X1 U19037 ( .C1(n16285), .C2(n15755), .A(n15754), .B(n15753), .ZN(
        n15756) );
  AOI211_X1 U19038 ( .C1(n15758), .C2(n15968), .A(n15757), .B(n15756), .ZN(
        n15763) );
  INV_X1 U19039 ( .A(n11542), .ZN(n15759) );
  AOI21_X1 U19040 ( .B1(n15761), .B2(n15760), .A(n15759), .ZN(n16551) );
  NAND2_X1 U19041 ( .A1(n16551), .A2(n19384), .ZN(n15762) );
  OAI211_X1 U19042 ( .C1(n16553), .C2(n15911), .A(n15763), .B(n15762), .ZN(
        P2_U2837) );
  INV_X1 U19043 ( .A(n15765), .ZN(n15764) );
  NOR3_X1 U19044 ( .A1(n15767), .A2(n19386), .A3(n15764), .ZN(n15772) );
  OAI21_X1 U19045 ( .B1(n15765), .B2(n19417), .A(n15957), .ZN(n15766) );
  NAND2_X1 U19046 ( .A1(n15767), .A2(n15766), .ZN(n15770) );
  INV_X1 U19047 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20235) );
  OAI21_X1 U19048 ( .B1(n20235), .B2(n15958), .A(n17200), .ZN(n15768) );
  AOI21_X1 U19049 ( .B1(n19403), .B2(P2_EBX_REG_17__SCAN_IN), .A(n15768), .ZN(
        n15769) );
  OAI211_X1 U19050 ( .C1(n11504), .C2(n19389), .A(n15770), .B(n15769), .ZN(
        n15771) );
  AOI211_X1 U19051 ( .C1(n15773), .C2(n15968), .A(n15772), .B(n15771), .ZN(
        n15777) );
  XOR2_X1 U19052 ( .A(n15775), .B(n15782), .Z(n16563) );
  NAND2_X1 U19053 ( .A1(n16563), .A2(n19384), .ZN(n15776) );
  OAI211_X1 U19054 ( .C1(n16566), .C2(n15911), .A(n15777), .B(n15776), .ZN(
        P2_U2838) );
  OR2_X1 U19055 ( .A1(n15779), .A2(n15780), .ZN(n15781) );
  NAND2_X1 U19056 ( .A1(n15782), .A2(n15781), .ZN(n16578) );
  AOI21_X1 U19057 ( .B1(n15783), .B2(n9731), .A(n11500), .ZN(n16582) );
  NAND2_X1 U19058 ( .A1(n16582), .A2(n19413), .ZN(n15794) );
  INV_X1 U19059 ( .A(n16293), .ZN(n15784) );
  NOR3_X1 U19060 ( .A1(n15784), .A2(n19387), .A3(n19386), .ZN(n15791) );
  NAND2_X1 U19061 ( .A1(n19387), .A2(n15942), .ZN(n15785) );
  AND2_X1 U19062 ( .A1(n15957), .A2(n15785), .ZN(n15789) );
  OAI21_X1 U19063 ( .B1(n15958), .B2(n20233), .A(n17200), .ZN(n15786) );
  AOI21_X1 U19064 ( .B1(n19403), .B2(P2_EBX_REG_16__SCAN_IN), .A(n15786), .ZN(
        n15788) );
  NAND2_X1 U19065 ( .A1(n19404), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15787) );
  OAI211_X1 U19066 ( .C1(n16293), .C2(n15789), .A(n15788), .B(n15787), .ZN(
        n15790) );
  AOI211_X1 U19067 ( .C1(n15792), .C2(n15968), .A(n15791), .B(n15790), .ZN(
        n15793) );
  OAI211_X1 U19068 ( .C1(n19407), .C2(n16578), .A(n15794), .B(n15793), .ZN(
        P2_U2839) );
  AND2_X1 U19069 ( .A1(n13586), .A2(n15795), .ZN(n15796) );
  NOR2_X1 U19070 ( .A1(n9665), .A2(n15796), .ZN(n16606) );
  AOI21_X1 U19071 ( .B1(n15942), .B2(n15797), .A(n19400), .ZN(n15800) );
  INV_X1 U19072 ( .A(n15797), .ZN(n15798) );
  NAND3_X1 U19073 ( .A1(n15967), .A2(n16315), .A3(n15798), .ZN(n15799) );
  OAI211_X1 U19074 ( .C1(n15800), .C2(n16315), .A(n17200), .B(n15799), .ZN(
        n15801) );
  AOI21_X1 U19075 ( .B1(n19410), .B2(P2_REIP_REG_14__SCAN_IN), .A(n15801), 
        .ZN(n15802) );
  OAI21_X1 U19076 ( .B1(n19392), .B2(n15803), .A(n15802), .ZN(n15804) );
  AOI21_X1 U19077 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19404), .A(
        n15804), .ZN(n15805) );
  OAI21_X1 U19078 ( .B1(n15806), .B2(n19405), .A(n15805), .ZN(n15807) );
  AOI21_X1 U19079 ( .B1(n16606), .B2(n19384), .A(n15807), .ZN(n15808) );
  OAI21_X1 U19080 ( .B1(n16608), .B2(n15911), .A(n15808), .ZN(P2_U2841) );
  INV_X1 U19081 ( .A(n15810), .ZN(n15811) );
  AOI21_X1 U19082 ( .B1(n15812), .B2(n15809), .A(n15811), .ZN(n16625) );
  INV_X1 U19083 ( .A(n16625), .ZN(n16062) );
  INV_X1 U19084 ( .A(n16631), .ZN(n15823) );
  AOI21_X1 U19085 ( .B1(n15942), .B2(n15813), .A(n19400), .ZN(n15816) );
  NAND3_X1 U19086 ( .A1(n15967), .A2(n16337), .A3(n15814), .ZN(n15815) );
  OAI211_X1 U19087 ( .C1(n15816), .C2(n16337), .A(n17200), .B(n15815), .ZN(
        n15818) );
  NOR2_X1 U19088 ( .A1(n15958), .A2(n20226), .ZN(n15817) );
  AOI211_X1 U19089 ( .C1(P2_EBX_REG_12__SCAN_IN), .C2(n19403), .A(n15818), .B(
        n15817), .ZN(n15820) );
  NAND2_X1 U19090 ( .A1(n19404), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15819) );
  OAI211_X1 U19091 ( .C1(n15821), .C2(n19405), .A(n15820), .B(n15819), .ZN(
        n15822) );
  AOI21_X1 U19092 ( .B1(n15823), .B2(n19384), .A(n15822), .ZN(n15824) );
  OAI21_X1 U19093 ( .B1(n16062), .B2(n15911), .A(n15824), .ZN(P2_U2843) );
  CLKBUF_X1 U19094 ( .A(n15825), .Z(n15844) );
  OAI21_X1 U19095 ( .B1(n10326), .B2(n11327), .A(n15809), .ZN(n16643) );
  AOI21_X1 U19096 ( .B1(n15829), .B2(n15828), .A(n15827), .ZN(n19436) );
  INV_X1 U19097 ( .A(n15836), .ZN(n15830) );
  NOR3_X1 U19098 ( .A1(n19386), .A2(n16346), .A3(n15830), .ZN(n15835) );
  INV_X1 U19099 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16344) );
  INV_X1 U19100 ( .A(n15831), .ZN(n15832) );
  AOI22_X1 U19101 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n19403), .B1(n15832), 
        .B2(n15968), .ZN(n15833) );
  OAI21_X1 U19102 ( .B1(n16344), .B2(n19389), .A(n15833), .ZN(n15834) );
  NOR3_X1 U19103 ( .A1(n15835), .A2(n19571), .A3(n15834), .ZN(n15839) );
  OAI21_X1 U19104 ( .B1(n15836), .B2(n19417), .A(n15957), .ZN(n15837) );
  NAND2_X1 U19105 ( .A1(n15837), .A2(n16346), .ZN(n15838) );
  OAI211_X1 U19106 ( .C1(n15958), .C2(n16343), .A(n15839), .B(n15838), .ZN(
        n15840) );
  AOI21_X1 U19107 ( .B1(n19436), .B2(n19384), .A(n15840), .ZN(n15841) );
  OAI21_X1 U19108 ( .B1(n16643), .B2(n15911), .A(n15841), .ZN(P2_U2844) );
  OR2_X1 U19109 ( .A1(n14330), .A2(n15842), .ZN(n15843) );
  NAND2_X1 U19110 ( .A1(n15844), .A2(n15843), .ZN(n16655) );
  NAND2_X1 U19111 ( .A1(n15845), .A2(n15968), .ZN(n15852) );
  AOI21_X1 U19112 ( .B1(n15942), .B2(n15846), .A(n19400), .ZN(n15848) );
  NAND3_X1 U19113 ( .A1(n15967), .A2(n16359), .A3(n9685), .ZN(n15847) );
  OAI211_X1 U19114 ( .C1(n15848), .C2(n16359), .A(n17200), .B(n15847), .ZN(
        n15850) );
  INV_X1 U19115 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n20223) );
  NOR2_X1 U19116 ( .A1(n15958), .A2(n20223), .ZN(n15849) );
  AOI211_X1 U19117 ( .C1(P2_EBX_REG_10__SCAN_IN), .C2(n19403), .A(n15850), .B(
        n15849), .ZN(n15851) );
  OAI211_X1 U19118 ( .C1(n19389), .C2(n15853), .A(n15852), .B(n15851), .ZN(
        n15854) );
  AOI21_X1 U19119 ( .B1(n16652), .B2(n19384), .A(n15854), .ZN(n15855) );
  OAI21_X1 U19120 ( .B1(n16655), .B2(n15911), .A(n15855), .ZN(P2_U2845) );
  NAND2_X1 U19121 ( .A1(n15857), .A2(n15856), .ZN(n15858) );
  NAND2_X1 U19122 ( .A1(n15859), .A2(n15858), .ZN(n19442) );
  INV_X1 U19123 ( .A(n16372), .ZN(n16663) );
  NAND2_X1 U19124 ( .A1(n16663), .A2(n19413), .ZN(n15871) );
  INV_X1 U19125 ( .A(n15861), .ZN(n15860) );
  OR2_X1 U19126 ( .A1(n16370), .A2(n15860), .ZN(n15868) );
  OAI21_X1 U19127 ( .B1(n15861), .B2(n19417), .A(n15957), .ZN(n15862) );
  NAND2_X1 U19128 ( .A1(n15862), .A2(n16370), .ZN(n15867) );
  AOI22_X1 U19129 ( .A1(P2_EBX_REG_9__SCAN_IN), .A2(n19403), .B1(n15863), .B2(
        n15968), .ZN(n15864) );
  OAI21_X1 U19130 ( .B1(n16368), .B2(n19389), .A(n15864), .ZN(n15865) );
  NOR2_X1 U19131 ( .A1(n19571), .A2(n15865), .ZN(n15866) );
  OAI211_X1 U19132 ( .C1(n19386), .C2(n15868), .A(n15867), .B(n15866), .ZN(
        n15869) );
  AOI21_X1 U19133 ( .B1(n19410), .B2(P2_REIP_REG_9__SCAN_IN), .A(n15869), .ZN(
        n15870) );
  OAI211_X1 U19134 ( .C1(n19407), .C2(n19442), .A(n15871), .B(n15870), .ZN(
        P2_U2846) );
  INV_X1 U19135 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n15881) );
  INV_X1 U19136 ( .A(n16387), .ZN(n15879) );
  OAI21_X1 U19137 ( .B1(n15872), .B2(n19417), .A(n15957), .ZN(n15878) );
  AOI22_X1 U19138 ( .A1(P2_EBX_REG_8__SCAN_IN), .A2(n19403), .B1(n15968), .B2(
        n15873), .ZN(n15874) );
  OAI211_X1 U19139 ( .C1(n20219), .C2(n15958), .A(n15874), .B(n17200), .ZN(
        n15877) );
  NOR3_X1 U19140 ( .A1(n15875), .A2(n19386), .A3(n15879), .ZN(n15876) );
  AOI211_X1 U19141 ( .C1(n15879), .C2(n15878), .A(n15877), .B(n15876), .ZN(
        n15880) );
  OAI21_X1 U19142 ( .B1(n19389), .B2(n15881), .A(n15880), .ZN(n15882) );
  AOI21_X1 U19143 ( .B1(n16678), .B2(n19384), .A(n15882), .ZN(n15883) );
  OAI21_X1 U19144 ( .B1(n16681), .B2(n15911), .A(n15883), .ZN(P2_U2847) );
  INV_X1 U19145 ( .A(n16691), .ZN(n15894) );
  OAI21_X1 U19146 ( .B1(n15887), .B2(n19417), .A(n15957), .ZN(n15891) );
  OAI22_X1 U19147 ( .A1(n15884), .A2(n19405), .B1(n16399), .B2(n19389), .ZN(
        n15885) );
  INV_X1 U19148 ( .A(n15885), .ZN(n15886) );
  OAI211_X1 U19149 ( .C1(n20217), .C2(n15958), .A(n15886), .B(n17200), .ZN(
        n15890) );
  INV_X1 U19150 ( .A(n15887), .ZN(n15888) );
  NOR3_X1 U19151 ( .A1(n19386), .A2(n16401), .A3(n15888), .ZN(n15889) );
  AOI211_X1 U19152 ( .C1(n16401), .C2(n15891), .A(n15890), .B(n15889), .ZN(
        n15892) );
  OAI21_X1 U19153 ( .B1(n19392), .B2(n14291), .A(n15892), .ZN(n15893) );
  AOI21_X1 U19154 ( .B1(n15894), .B2(n19413), .A(n15893), .ZN(n15895) );
  OAI21_X1 U19155 ( .B1(n19407), .B2(n16687), .A(n15895), .ZN(P2_U2848) );
  INV_X1 U19156 ( .A(n15896), .ZN(n16377) );
  NAND2_X1 U19157 ( .A1(n15942), .A2(n15898), .ZN(n15897) );
  AOI21_X1 U19158 ( .B1(n15957), .B2(n15897), .A(n16409), .ZN(n15902) );
  INV_X1 U19159 ( .A(n15898), .ZN(n15899) );
  NAND3_X1 U19160 ( .A1(n15967), .A2(n16409), .A3(n15899), .ZN(n15900) );
  NAND2_X1 U19161 ( .A1(n15900), .A2(n17200), .ZN(n15901) );
  AOI211_X1 U19162 ( .C1(n19410), .C2(P2_REIP_REG_6__SCAN_IN), .A(n15902), .B(
        n15901), .ZN(n15904) );
  NAND2_X1 U19163 ( .A1(n19403), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n15903) );
  OAI211_X1 U19164 ( .C1(n19389), .C2(n10112), .A(n15904), .B(n15903), .ZN(
        n15909) );
  OAI21_X1 U19165 ( .B1(n15907), .B2(n15906), .A(n15905), .ZN(n19446) );
  NOR2_X1 U19166 ( .A1(n19446), .A2(n19407), .ZN(n15908) );
  AOI211_X1 U19167 ( .C1(n15968), .C2(n16377), .A(n15909), .B(n15908), .ZN(
        n15910) );
  OAI21_X1 U19168 ( .B1(n15911), .B2(n16698), .A(n15910), .ZN(P2_U2849) );
  OAI21_X1 U19169 ( .B1(n14361), .B2(n15913), .A(n15912), .ZN(n19449) );
  NAND2_X1 U19170 ( .A1(n17194), .A2(n19413), .ZN(n15925) );
  NAND2_X1 U19171 ( .A1(n19403), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n15919) );
  OAI21_X1 U19172 ( .B1(n15914), .B2(n19417), .A(n15957), .ZN(n15917) );
  INV_X1 U19173 ( .A(n15914), .ZN(n15915) );
  NOR3_X1 U19174 ( .A1(n17191), .A2(n15915), .A3(n19386), .ZN(n15916) );
  AOI211_X1 U19175 ( .C1(n17191), .C2(n15917), .A(n19571), .B(n15916), .ZN(
        n15918) );
  OAI211_X1 U19176 ( .C1(n15958), .C2(n15920), .A(n15919), .B(n15918), .ZN(
        n15923) );
  NOR2_X1 U19177 ( .A1(n15921), .A2(n19405), .ZN(n15922) );
  AOI211_X1 U19178 ( .C1(n19404), .C2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n15923), .B(n15922), .ZN(n15924) );
  OAI211_X1 U19179 ( .C1(n19449), .C2(n19407), .A(n15925), .B(n15924), .ZN(
        P2_U2850) );
  NAND2_X1 U19180 ( .A1(n20278), .A2(n19384), .ZN(n15934) );
  OAI21_X1 U19181 ( .B1(n19417), .B2(n15928), .A(n15957), .ZN(n15926) );
  NAND2_X1 U19182 ( .A1(n15926), .A2(n15927), .ZN(n15930) );
  NAND3_X1 U19183 ( .A1(n15967), .A2(n10182), .A3(n15928), .ZN(n15929) );
  OAI211_X1 U19184 ( .C1(n15958), .C2(n17201), .A(n15930), .B(n15929), .ZN(
        n15932) );
  NOR2_X1 U19185 ( .A1(n19389), .A2(n16420), .ZN(n15931) );
  AOI211_X1 U19186 ( .C1(P2_EBX_REG_3__SCAN_IN), .C2(n19403), .A(n15932), .B(
        n15931), .ZN(n15933) );
  OAI211_X1 U19187 ( .C1(n19405), .C2(n15935), .A(n15934), .B(n15933), .ZN(
        n15936) );
  OAI21_X1 U19188 ( .B1(n16821), .B2(n19412), .A(n15937), .ZN(P2_U2852) );
  NOR2_X1 U19189 ( .A1(n19405), .A2(n15938), .ZN(n15949) );
  INV_X1 U19190 ( .A(n15939), .ZN(n15940) );
  AND2_X1 U19191 ( .A1(n16761), .A2(n15940), .ZN(n15956) );
  INV_X1 U19192 ( .A(n15941), .ZN(n15944) );
  OAI21_X1 U19193 ( .B1(n15956), .B2(n15944), .A(n15942), .ZN(n15943) );
  AOI21_X1 U19194 ( .B1(n15956), .B2(n15944), .A(n15943), .ZN(n15945) );
  AOI21_X1 U19195 ( .B1(n19410), .B2(P2_REIP_REG_2__SCAN_IN), .A(n15945), .ZN(
        n15946) );
  OAI21_X1 U19196 ( .B1(n19392), .B2(n15947), .A(n15946), .ZN(n15948) );
  AOI211_X1 U19197 ( .C1(n19404), .C2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n15949), .B(n15948), .ZN(n15950) );
  OAI21_X1 U19198 ( .B1(n20286), .B2(n19407), .A(n15950), .ZN(n15951) );
  AOI21_X1 U19199 ( .B1(n15952), .B2(n19413), .A(n15951), .ZN(n15953) );
  OAI21_X1 U19200 ( .B1(n20288), .B2(n19412), .A(n15953), .ZN(P2_U2853) );
  NAND2_X1 U19201 ( .A1(n16773), .A2(n15954), .ZN(n15955) );
  NAND2_X1 U19202 ( .A1(n15956), .A2(n15955), .ZN(n16775) );
  OAI22_X1 U19203 ( .A1(n16775), .A2(n19417), .B1(n15957), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15960) );
  NOR2_X1 U19204 ( .A1(n15958), .A2(n10958), .ZN(n15959) );
  AOI211_X1 U19205 ( .C1(n15968), .C2(n15961), .A(n15960), .B(n15959), .ZN(
        n15963) );
  AOI22_X1 U19206 ( .A1(n19403), .A2(P2_EBX_REG_1__SCAN_IN), .B1(n19404), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15962) );
  OAI211_X1 U19207 ( .C1(n16759), .C2(n19407), .A(n15963), .B(n15962), .ZN(
        n15964) );
  AOI21_X1 U19208 ( .B1(n16746), .B2(n19413), .A(n15964), .ZN(n15965) );
  OAI21_X1 U19209 ( .B1(n20275), .B2(n19412), .A(n15965), .ZN(P2_U2854) );
  INV_X1 U19210 ( .A(n15966), .ZN(n19481) );
  AOI22_X1 U19211 ( .A1(n19384), .A2(n19481), .B1(n19410), .B2(
        P2_REIP_REG_0__SCAN_IN), .ZN(n15972) );
  AOI22_X1 U19212 ( .A1(n15968), .A2(n17221), .B1(n15967), .B2(n16773), .ZN(
        n15971) );
  OAI21_X1 U19213 ( .B1(n19404), .B2(n19400), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15970) );
  NAND2_X1 U19214 ( .A1(n19403), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n15969) );
  NAND4_X1 U19215 ( .A1(n15972), .A2(n15971), .A3(n15970), .A4(n15969), .ZN(
        n15973) );
  AOI21_X1 U19216 ( .B1(n19593), .B2(n19413), .A(n15973), .ZN(n15974) );
  OAI21_X1 U19217 ( .B1(n16820), .B2(n19412), .A(n15974), .ZN(P2_U2855) );
  OR2_X1 U19218 ( .A1(n15976), .A2(n15975), .ZN(n16080) );
  NAND3_X1 U19219 ( .A1(n16080), .A2(n15977), .A3(n19426), .ZN(n15979) );
  NAND2_X1 U19220 ( .A1(n16073), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15978) );
  OAI211_X1 U19221 ( .C1(n16073), .C2(n15599), .A(n15979), .B(n15978), .ZN(
        P2_U2858) );
  NOR2_X1 U19222 ( .A1(n9666), .A2(n15980), .ZN(n15982) );
  XNOR2_X1 U19223 ( .A(n15982), .B(n15981), .ZN(n16091) );
  NAND2_X1 U19224 ( .A1(n16091), .A2(n19426), .ZN(n15984) );
  NAND2_X1 U19225 ( .A1(n16073), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n15983) );
  OAI211_X1 U19226 ( .C1(n11525), .C2(n16073), .A(n15984), .B(n15983), .ZN(
        P2_U2859) );
  OAI21_X1 U19227 ( .B1(n15987), .B2(n15986), .A(n15985), .ZN(n16106) );
  NAND2_X1 U19228 ( .A1(n16073), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n15989) );
  NAND2_X1 U19229 ( .A1(n16437), .A2(n19429), .ZN(n15988) );
  OAI211_X1 U19230 ( .C1(n16106), .C2(n16066), .A(n15989), .B(n15988), .ZN(
        P2_U2860) );
  NOR2_X1 U19231 ( .A1(n16001), .A2(n16000), .ZN(n15999) );
  NOR2_X1 U19232 ( .A1(n15999), .A2(n15990), .ZN(n15996) );
  NOR2_X1 U19233 ( .A1(n15992), .A2(n15991), .ZN(n15993) );
  XNOR2_X1 U19234 ( .A(n15994), .B(n15993), .ZN(n15995) );
  XNOR2_X1 U19235 ( .A(n15996), .B(n15995), .ZN(n16113) );
  NOR2_X1 U19236 ( .A1(n16460), .A2(n16073), .ZN(n15997) );
  AOI21_X1 U19237 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n16073), .A(n15997), .ZN(
        n15998) );
  OAI21_X1 U19238 ( .B1(n16113), .B2(n16066), .A(n15998), .ZN(P2_U2861) );
  INV_X1 U19239 ( .A(n16473), .ZN(n16004) );
  AOI21_X1 U19240 ( .B1(n16001), .B2(n16000), .A(n15999), .ZN(n16114) );
  NAND2_X1 U19241 ( .A1(n16114), .A2(n19426), .ZN(n16003) );
  NAND2_X1 U19242 ( .A1(n16073), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n16002) );
  OAI211_X1 U19243 ( .C1(n16004), .C2(n16073), .A(n16003), .B(n16002), .ZN(
        P2_U2862) );
  AOI21_X1 U19244 ( .B1(n16007), .B2(n16006), .A(n16005), .ZN(n16008) );
  XOR2_X1 U19245 ( .A(n16009), .B(n16008), .Z(n16128) );
  MUX2_X1 U19246 ( .A(n16487), .B(n16010), .S(n16073), .Z(n16011) );
  OAI21_X1 U19247 ( .B1(n16128), .B2(n16066), .A(n16011), .ZN(P2_U2863) );
  AOI21_X1 U19248 ( .B1(n16012), .B2(n16014), .A(n16013), .ZN(n16129) );
  NAND2_X1 U19249 ( .A1(n16129), .A2(n19426), .ZN(n16016) );
  NAND2_X1 U19250 ( .A1(n16073), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n16015) );
  OAI211_X1 U19251 ( .C1(n16495), .C2(n16073), .A(n16016), .B(n16015), .ZN(
        P2_U2864) );
  AOI21_X1 U19252 ( .B1(n16019), .B2(n16017), .A(n16018), .ZN(n16136) );
  AOI22_X1 U19253 ( .A1(n16136), .A2(n19426), .B1(P2_EBX_REG_22__SCAN_IN), 
        .B2(n16073), .ZN(n16020) );
  OAI21_X1 U19254 ( .B1(n16021), .B2(n16073), .A(n16020), .ZN(P2_U2865) );
  NAND2_X1 U19255 ( .A1(n16022), .A2(n16023), .ZN(n16024) );
  AND2_X1 U19256 ( .A1(n16017), .A2(n16024), .ZN(n16147) );
  AOI22_X1 U19257 ( .A1(n16147), .A2(n19426), .B1(P2_EBX_REG_21__SCAN_IN), 
        .B2(n16073), .ZN(n16025) );
  OAI21_X1 U19258 ( .B1(n16528), .B2(n16073), .A(n16025), .ZN(P2_U2866) );
  INV_X1 U19259 ( .A(n16533), .ZN(n16029) );
  OAI21_X1 U19260 ( .B1(n9730), .B2(n16026), .A(n16022), .ZN(n16162) );
  INV_X1 U19261 ( .A(n16162), .ZN(n16027) );
  AOI22_X1 U19262 ( .A1(n16027), .A2(n19426), .B1(P2_EBX_REG_20__SCAN_IN), 
        .B2(n16073), .ZN(n16028) );
  OAI21_X1 U19263 ( .B1(n16029), .B2(n16073), .A(n16028), .ZN(P2_U2867) );
  AOI21_X1 U19264 ( .B1(n10420), .B2(n16030), .A(n9730), .ZN(n16170) );
  AOI22_X1 U19265 ( .A1(n16170), .A2(n19426), .B1(P2_EBX_REG_19__SCAN_IN), 
        .B2(n16073), .ZN(n16031) );
  OAI21_X1 U19266 ( .B1(n16032), .B2(n16073), .A(n16031), .ZN(P2_U2868) );
  NOR2_X1 U19267 ( .A1(n16033), .A2(n16034), .ZN(n16035) );
  OR2_X1 U19268 ( .A1(n16036), .A2(n16035), .ZN(n16181) );
  OAI22_X1 U19269 ( .A1(n16181), .A2(n16066), .B1(n19429), .B2(n16037), .ZN(
        n16038) );
  INV_X1 U19270 ( .A(n16038), .ZN(n16039) );
  OAI21_X1 U19271 ( .B1(n16553), .B2(n16073), .A(n16039), .ZN(P2_U2869) );
  AOI21_X1 U19272 ( .B1(n16041), .B2(n16040), .A(n16033), .ZN(n16189) );
  AOI22_X1 U19273 ( .A1(n16189), .A2(n19426), .B1(P2_EBX_REG_17__SCAN_IN), 
        .B2(n16073), .ZN(n16042) );
  OAI21_X1 U19274 ( .B1(n16566), .B2(n16073), .A(n16042), .ZN(P2_U2870) );
  NOR2_X1 U19275 ( .A1(n16048), .A2(n16047), .ZN(n16044) );
  OAI21_X1 U19276 ( .B1(n16044), .B2(n16043), .A(n16040), .ZN(n16205) );
  NAND2_X1 U19277 ( .A1(n16582), .A2(n19429), .ZN(n16046) );
  NAND2_X1 U19278 ( .A1(n16073), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n16045) );
  OAI211_X1 U19279 ( .C1(n16205), .C2(n16066), .A(n16046), .B(n16045), .ZN(
        P2_U2871) );
  XNOR2_X1 U19280 ( .A(n16048), .B(n16047), .ZN(n16054) );
  NAND2_X1 U19281 ( .A1(n16050), .A2(n16049), .ZN(n16051) );
  NAND2_X1 U19282 ( .A1(n9731), .A2(n16051), .ZN(n19382) );
  NOR2_X1 U19283 ( .A1(n19382), .A2(n16073), .ZN(n16052) );
  AOI21_X1 U19284 ( .B1(P2_EBX_REG_15__SCAN_IN), .B2(n16073), .A(n16052), .ZN(
        n16053) );
  OAI21_X1 U19285 ( .B1(n16054), .B2(n16066), .A(n16053), .ZN(P2_U2872) );
  NOR2_X1 U19286 ( .A1(n16056), .A2(n16055), .ZN(n16070) );
  NAND2_X1 U19287 ( .A1(n16070), .A2(n16069), .ZN(n16068) );
  NOR2_X1 U19288 ( .A1(n16068), .A2(n16063), .ZN(n16059) );
  OAI211_X1 U19289 ( .C1(n16059), .C2(n16058), .A(n19426), .B(n16057), .ZN(
        n16061) );
  NAND2_X1 U19290 ( .A1(n16073), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n16060) );
  OAI211_X1 U19291 ( .C1(n16062), .C2(n16073), .A(n16061), .B(n16060), .ZN(
        P2_U2875) );
  XNOR2_X1 U19292 ( .A(n16068), .B(n16063), .ZN(n16067) );
  MUX2_X1 U19293 ( .A(n16064), .B(n16643), .S(n19429), .Z(n16065) );
  OAI21_X1 U19294 ( .B1(n16067), .B2(n16066), .A(n16065), .ZN(P2_U2876) );
  OAI211_X1 U19295 ( .C1(n16070), .C2(n16069), .A(n16068), .B(n19426), .ZN(
        n16072) );
  NAND2_X1 U19296 ( .A1(n16073), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n16071) );
  OAI211_X1 U19297 ( .C1(n16655), .C2(n16073), .A(n16072), .B(n16071), .ZN(
        P2_U2877) );
  INV_X1 U19298 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n16076) );
  NAND2_X1 U19299 ( .A1(n16193), .A2(BUF1_REG_30__SCAN_IN), .ZN(n16075) );
  MUX2_X1 U19300 ( .A(BUF1_REG_14__SCAN_IN), .B(BUF2_REG_14__SCAN_IN), .S(
        n19430), .Z(n19537) );
  AOI22_X1 U19301 ( .A1(n16197), .A2(n19537), .B1(n19476), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n16074) );
  OAI211_X1 U19302 ( .C1(n16076), .C2(n16200), .A(n16075), .B(n16074), .ZN(
        n16077) );
  AOI21_X1 U19303 ( .B1(n14612), .B2(n19477), .A(n16077), .ZN(n16078) );
  OAI21_X1 U19304 ( .B1(n16079), .B2(n19472), .A(n16078), .ZN(P2_U2889) );
  NAND3_X1 U19305 ( .A1(n16080), .A2(n15977), .A3(n19479), .ZN(n16090) );
  INV_X1 U19306 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n16082) );
  AOI22_X1 U19307 ( .A1(n16197), .A2(n19535), .B1(n19476), .B2(
        P2_EAX_REG_29__SCAN_IN), .ZN(n16081) );
  OAI21_X1 U19308 ( .B1(n16200), .B2(n16082), .A(n16081), .ZN(n16086) );
  INV_X1 U19309 ( .A(n16193), .ZN(n16084) );
  NOR2_X1 U19310 ( .A1(n16084), .A2(n16083), .ZN(n16085) );
  OR2_X1 U19311 ( .A1(n16086), .A2(n16085), .ZN(n16087) );
  NAND2_X1 U19312 ( .A1(n16090), .A2(n16089), .ZN(P2_U2890) );
  INV_X1 U19313 ( .A(n16091), .ZN(n16099) );
  INV_X1 U19314 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n16095) );
  NAND2_X1 U19315 ( .A1(n16193), .A2(BUF1_REG_28__SCAN_IN), .ZN(n16094) );
  INV_X1 U19316 ( .A(n19561), .ZN(n16092) );
  AOI22_X1 U19317 ( .A1(n16197), .A2(n16092), .B1(n19476), .B2(
        P2_EAX_REG_28__SCAN_IN), .ZN(n16093) );
  OAI211_X1 U19318 ( .C1(n16095), .C2(n16200), .A(n16094), .B(n16093), .ZN(
        n16096) );
  AOI21_X1 U19319 ( .B1(n16097), .B2(n19477), .A(n16096), .ZN(n16098) );
  OAI21_X1 U19320 ( .B1(n16099), .B2(n19472), .A(n16098), .ZN(P2_U2891) );
  INV_X1 U19321 ( .A(n16446), .ZN(n16104) );
  INV_X1 U19322 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n16102) );
  NAND2_X1 U19323 ( .A1(n16193), .A2(BUF1_REG_27__SCAN_IN), .ZN(n16101) );
  AOI22_X1 U19324 ( .A1(n16197), .A2(n19435), .B1(n19476), .B2(
        P2_EAX_REG_27__SCAN_IN), .ZN(n16100) );
  OAI211_X1 U19325 ( .C1(n16102), .C2(n16200), .A(n16101), .B(n16100), .ZN(
        n16103) );
  AOI21_X1 U19326 ( .B1(n16104), .B2(n19477), .A(n16103), .ZN(n16105) );
  OAI21_X1 U19327 ( .B1(n16106), .B2(n19472), .A(n16105), .ZN(P2_U2892) );
  INV_X1 U19328 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n16110) );
  NAND2_X1 U19329 ( .A1(n16193), .A2(BUF1_REG_26__SCAN_IN), .ZN(n16109) );
  INV_X1 U19330 ( .A(n19559), .ZN(n16107) );
  AOI22_X1 U19331 ( .A1(n16197), .A2(n16107), .B1(n19476), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n16108) );
  OAI211_X1 U19332 ( .C1(n16110), .C2(n16200), .A(n16109), .B(n16108), .ZN(
        n16111) );
  AOI21_X1 U19333 ( .B1(n16458), .B2(n19477), .A(n16111), .ZN(n16112) );
  OAI21_X1 U19334 ( .B1(n16113), .B2(n19472), .A(n16112), .ZN(P2_U2893) );
  INV_X1 U19335 ( .A(n16114), .ZN(n16121) );
  INV_X1 U19336 ( .A(n16470), .ZN(n16119) );
  INV_X1 U19337 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n16117) );
  NAND2_X1 U19338 ( .A1(n16193), .A2(BUF1_REG_25__SCAN_IN), .ZN(n16116) );
  AOI22_X1 U19339 ( .A1(n16197), .A2(n19439), .B1(n19476), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n16115) );
  OAI211_X1 U19340 ( .C1(n16117), .C2(n16200), .A(n16116), .B(n16115), .ZN(
        n16118) );
  AOI21_X1 U19341 ( .B1(n16119), .B2(n19477), .A(n16118), .ZN(n16120) );
  OAI21_X1 U19342 ( .B1(n16121), .B2(n19472), .A(n16120), .ZN(P2_U2894) );
  INV_X1 U19343 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n16125) );
  NAND2_X1 U19344 ( .A1(n16193), .A2(BUF1_REG_24__SCAN_IN), .ZN(n16124) );
  INV_X1 U19345 ( .A(n19557), .ZN(n16122) );
  AOI22_X1 U19346 ( .A1(n16197), .A2(n16122), .B1(n19476), .B2(
        P2_EAX_REG_24__SCAN_IN), .ZN(n16123) );
  OAI211_X1 U19347 ( .C1(n16125), .C2(n16200), .A(n16124), .B(n16123), .ZN(
        n16126) );
  AOI21_X1 U19348 ( .B1(n16479), .B2(n19477), .A(n16126), .ZN(n16127) );
  OAI21_X1 U19349 ( .B1(n16128), .B2(n19472), .A(n16127), .ZN(P2_U2895) );
  INV_X1 U19350 ( .A(n16129), .ZN(n16135) );
  INV_X1 U19351 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n16132) );
  NAND2_X1 U19352 ( .A1(n16193), .A2(BUF1_REG_23__SCAN_IN), .ZN(n16131) );
  INV_X1 U19353 ( .A(n19555), .ZN(n19646) );
  AOI22_X1 U19354 ( .A1(n16197), .A2(n19646), .B1(n19476), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n16130) );
  OAI211_X1 U19355 ( .C1(n16132), .C2(n16200), .A(n16131), .B(n16130), .ZN(
        n16133) );
  AOI21_X1 U19356 ( .B1(n16498), .B2(n19477), .A(n16133), .ZN(n16134) );
  OAI21_X1 U19357 ( .B1(n19472), .B2(n16135), .A(n16134), .ZN(P2_U2896) );
  INV_X1 U19358 ( .A(n16136), .ZN(n16146) );
  INV_X1 U19359 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n16142) );
  NAND2_X1 U19360 ( .A1(n16193), .A2(BUF1_REG_22__SCAN_IN), .ZN(n16141) );
  INV_X1 U19361 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16137) );
  OR2_X1 U19362 ( .A1(n19430), .A2(n16137), .ZN(n16139) );
  NAND2_X1 U19363 ( .A1(n19430), .A2(BUF2_REG_6__SCAN_IN), .ZN(n16138) );
  AND2_X1 U19364 ( .A1(n16139), .A2(n16138), .ZN(n19553) );
  INV_X1 U19365 ( .A(n19553), .ZN(n19635) );
  AOI22_X1 U19366 ( .A1(n16197), .A2(n19635), .B1(n19476), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n16140) );
  OAI211_X1 U19367 ( .C1(n16142), .C2(n16200), .A(n16141), .B(n16140), .ZN(
        n16143) );
  AOI21_X1 U19368 ( .B1(n16144), .B2(n19477), .A(n16143), .ZN(n16145) );
  OAI21_X1 U19369 ( .B1(n19472), .B2(n16146), .A(n16145), .ZN(P2_U2897) );
  INV_X1 U19370 ( .A(n16147), .ZN(n16156) );
  INV_X1 U19371 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n16153) );
  NAND2_X1 U19372 ( .A1(n16193), .A2(BUF1_REG_21__SCAN_IN), .ZN(n16152) );
  INV_X1 U19373 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16148) );
  OR2_X1 U19374 ( .A1(n19430), .A2(n16148), .ZN(n16150) );
  NAND2_X1 U19375 ( .A1(n19430), .A2(BUF2_REG_5__SCAN_IN), .ZN(n16149) );
  AND2_X1 U19376 ( .A1(n16150), .A2(n16149), .ZN(n19551) );
  INV_X1 U19377 ( .A(n19551), .ZN(n16828) );
  AOI22_X1 U19378 ( .A1(n16197), .A2(n16828), .B1(n19476), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n16151) );
  OAI211_X1 U19379 ( .C1(n16200), .C2(n16153), .A(n16152), .B(n16151), .ZN(
        n16154) );
  AOI21_X1 U19380 ( .B1(n16526), .B2(n19477), .A(n16154), .ZN(n16155) );
  OAI21_X1 U19381 ( .B1(n19472), .B2(n16156), .A(n16155), .ZN(P2_U2898) );
  INV_X1 U19382 ( .A(n16541), .ZN(n16160) );
  INV_X1 U19383 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n16872) );
  NAND2_X1 U19384 ( .A1(n16193), .A2(BUF1_REG_20__SCAN_IN), .ZN(n16158) );
  AOI22_X1 U19385 ( .A1(n16197), .A2(n19626), .B1(n19476), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n16157) );
  OAI211_X1 U19386 ( .C1(n16872), .C2(n16200), .A(n16158), .B(n16157), .ZN(
        n16159) );
  AOI21_X1 U19387 ( .B1(n16160), .B2(n19477), .A(n16159), .ZN(n16161) );
  OAI21_X1 U19388 ( .B1(n19472), .B2(n16162), .A(n16161), .ZN(P2_U2899) );
  INV_X1 U19389 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n16168) );
  NAND2_X1 U19390 ( .A1(n16193), .A2(BUF1_REG_19__SCAN_IN), .ZN(n16167) );
  INV_X1 U19391 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16163) );
  OR2_X1 U19392 ( .A1(n19430), .A2(n16163), .ZN(n16165) );
  NAND2_X1 U19393 ( .A1(n19430), .A2(BUF2_REG_3__SCAN_IN), .ZN(n16164) );
  AND2_X1 U19394 ( .A1(n16165), .A2(n16164), .ZN(n19547) );
  INV_X1 U19395 ( .A(n19547), .ZN(n19621) );
  AOI22_X1 U19396 ( .A1(n16197), .A2(n19621), .B1(n19476), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n16166) );
  OAI211_X1 U19397 ( .C1(n16168), .C2(n16200), .A(n16167), .B(n16166), .ZN(
        n16169) );
  AOI21_X1 U19398 ( .B1(n16170), .B2(n19479), .A(n16169), .ZN(n16171) );
  OAI21_X1 U19399 ( .B1(n16172), .B2(n16191), .A(n16171), .ZN(P2_U2900) );
  INV_X1 U19400 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n16178) );
  NAND2_X1 U19401 ( .A1(n16193), .A2(BUF1_REG_18__SCAN_IN), .ZN(n16177) );
  INV_X1 U19402 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16173) );
  OR2_X1 U19403 ( .A1(n19430), .A2(n16173), .ZN(n16175) );
  NAND2_X1 U19404 ( .A1(n19430), .A2(BUF2_REG_2__SCAN_IN), .ZN(n16174) );
  AND2_X1 U19405 ( .A1(n16175), .A2(n16174), .ZN(n19545) );
  INV_X1 U19406 ( .A(n19545), .ZN(n19616) );
  AOI22_X1 U19407 ( .A1(n16197), .A2(n19616), .B1(n19476), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n16176) );
  OAI211_X1 U19408 ( .C1(n16178), .C2(n16200), .A(n16177), .B(n16176), .ZN(
        n16179) );
  AOI21_X1 U19409 ( .B1(n16551), .B2(n19477), .A(n16179), .ZN(n16180) );
  OAI21_X1 U19410 ( .B1(n19472), .B2(n16181), .A(n16180), .ZN(P2_U2901) );
  INV_X1 U19411 ( .A(n16563), .ZN(n16192) );
  INV_X1 U19412 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n16187) );
  NAND2_X1 U19413 ( .A1(n16193), .A2(BUF1_REG_17__SCAN_IN), .ZN(n16186) );
  OR2_X1 U19414 ( .A1(n19430), .A2(n16182), .ZN(n16184) );
  NAND2_X1 U19415 ( .A1(n19430), .A2(BUF2_REG_1__SCAN_IN), .ZN(n16183) );
  AND2_X1 U19416 ( .A1(n16184), .A2(n16183), .ZN(n19543) );
  INV_X1 U19417 ( .A(n19543), .ZN(n19611) );
  AOI22_X1 U19418 ( .A1(n16197), .A2(n19611), .B1(n19476), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n16185) );
  OAI211_X1 U19419 ( .C1(n16187), .C2(n16200), .A(n16186), .B(n16185), .ZN(
        n16188) );
  AOI21_X1 U19420 ( .B1(n16189), .B2(n19479), .A(n16188), .ZN(n16190) );
  OAI21_X1 U19421 ( .B1(n16192), .B2(n16191), .A(n16190), .ZN(P2_U2902) );
  INV_X1 U19422 ( .A(n16578), .ZN(n16203) );
  NAND2_X1 U19423 ( .A1(n16193), .A2(BUF1_REG_16__SCAN_IN), .ZN(n16199) );
  INV_X1 U19424 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16194) );
  OR2_X1 U19425 ( .A1(n19430), .A2(n16194), .ZN(n16196) );
  NAND2_X1 U19426 ( .A1(n19430), .A2(BUF2_REG_0__SCAN_IN), .ZN(n16195) );
  AND2_X1 U19427 ( .A1(n16196), .A2(n16195), .ZN(n19541) );
  INV_X1 U19428 ( .A(n19541), .ZN(n16808) );
  AOI22_X1 U19429 ( .A1(n16197), .A2(n16808), .B1(n19476), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n16198) );
  OAI211_X1 U19430 ( .C1(n16201), .C2(n16200), .A(n16199), .B(n16198), .ZN(
        n16202) );
  AOI21_X1 U19431 ( .B1(n16203), .B2(n19477), .A(n16202), .ZN(n16204) );
  OAI21_X1 U19432 ( .B1(n16205), .B2(n19472), .A(n16204), .ZN(P2_U2903) );
  INV_X1 U19433 ( .A(n16606), .ZN(n16207) );
  AOI22_X1 U19434 ( .A1(n19434), .A2(n19537), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n19476), .ZN(n16206) );
  OAI21_X1 U19435 ( .B1(n16207), .B2(n19441), .A(n16206), .ZN(P2_U2905) );
  XNOR2_X1 U19436 ( .A(n16208), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16450) );
  NAND2_X1 U19437 ( .A1(n19571), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n16440) );
  NAND2_X1 U19438 ( .A1(n19584), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16209) );
  OAI211_X1 U19439 ( .C1(n19582), .C2(n16210), .A(n16440), .B(n16209), .ZN(
        n16211) );
  AOI21_X1 U19440 ( .B1(n16437), .B2(n19592), .A(n16211), .ZN(n16214) );
  AOI21_X1 U19441 ( .B1(n16438), .B2(n16212), .A(n11418), .ZN(n16448) );
  NAND2_X1 U19442 ( .A1(n16448), .A2(n19577), .ZN(n16213) );
  OAI211_X1 U19443 ( .C1(n16450), .C2(n19574), .A(n16214), .B(n16213), .ZN(
        P2_U2987) );
  OAI21_X1 U19444 ( .B1(n16230), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n16212), .ZN(n16464) );
  OAI21_X1 U19445 ( .B1(n16215), .B2(n16224), .A(n16225), .ZN(n16217) );
  XNOR2_X1 U19446 ( .A(n16217), .B(n16216), .ZN(n16462) );
  NAND2_X1 U19447 ( .A1(n19571), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n16455) );
  OAI21_X1 U19448 ( .B1(n17198), .B2(n16218), .A(n16455), .ZN(n16219) );
  AOI21_X1 U19449 ( .B1(n17192), .B2(n16220), .A(n16219), .ZN(n16221) );
  OAI21_X1 U19450 ( .B1(n16460), .B2(n19573), .A(n16221), .ZN(n16222) );
  AOI21_X1 U19451 ( .B1(n16462), .B2(n9627), .A(n16222), .ZN(n16223) );
  OAI21_X1 U19452 ( .B1(n19590), .B2(n16464), .A(n16223), .ZN(P2_U2988) );
  NAND2_X1 U19453 ( .A1(n9937), .A2(n16225), .ZN(n16226) );
  XNOR2_X1 U19454 ( .A(n16215), .B(n16226), .ZN(n16478) );
  NAND2_X1 U19455 ( .A1(n19571), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n16467) );
  NAND2_X1 U19456 ( .A1(n19584), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16227) );
  OAI211_X1 U19457 ( .C1(n19582), .C2(n16228), .A(n16467), .B(n16227), .ZN(
        n16229) );
  AOI21_X1 U19458 ( .B1(n16473), .B2(n19592), .A(n16229), .ZN(n16232) );
  INV_X1 U19459 ( .A(n16230), .ZN(n16475) );
  NAND2_X1 U19460 ( .A1(n16235), .A2(n16468), .ZN(n16474) );
  NAND3_X1 U19461 ( .A1(n16475), .A2(n19577), .A3(n16474), .ZN(n16231) );
  OAI211_X1 U19462 ( .C1(n16478), .C2(n19574), .A(n16232), .B(n16231), .ZN(
        P2_U2989) );
  INV_X1 U19463 ( .A(n16233), .ZN(n16234) );
  OAI21_X1 U19464 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n16234), .A(
        n16235), .ZN(n16491) );
  NAND2_X1 U19465 ( .A1(n9691), .A2(n16236), .ZN(n16237) );
  XNOR2_X1 U19466 ( .A(n16238), .B(n16237), .ZN(n16489) );
  NOR2_X1 U19467 ( .A1(n17200), .A2(n20248), .ZN(n16482) );
  AOI21_X1 U19468 ( .B1(n19584), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n16482), .ZN(n16241) );
  NAND2_X1 U19469 ( .A1(n17192), .A2(n16239), .ZN(n16240) );
  OAI211_X1 U19470 ( .C1(n16487), .C2(n19573), .A(n16241), .B(n16240), .ZN(
        n16242) );
  AOI21_X1 U19471 ( .B1(n16489), .B2(n9627), .A(n16242), .ZN(n16243) );
  OAI21_X1 U19472 ( .B1(n19590), .B2(n16491), .A(n16243), .ZN(P2_U2990) );
  INV_X1 U19473 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16257) );
  OAI21_X1 U19474 ( .B1(n16256), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16233), .ZN(n16502) );
  INV_X1 U19475 ( .A(n16495), .ZN(n16247) );
  NAND2_X1 U19476 ( .A1(n19571), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n16492) );
  NAND2_X1 U19477 ( .A1(n19584), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16244) );
  OAI211_X1 U19478 ( .C1(n19582), .C2(n16245), .A(n16492), .B(n16244), .ZN(
        n16246) );
  AOI21_X1 U19479 ( .B1(n16247), .B2(n19592), .A(n16246), .ZN(n16252) );
  OR2_X1 U19480 ( .A1(n16249), .A2(n16248), .ZN(n16499) );
  NAND3_X1 U19481 ( .A1(n16499), .A2(n16250), .A3(n9627), .ZN(n16251) );
  OAI211_X1 U19482 ( .C1(n16502), .C2(n19590), .A(n16252), .B(n16251), .ZN(
        P2_U2991) );
  NAND2_X1 U19483 ( .A1(n9736), .A2(n16253), .ZN(n16254) );
  XNOR2_X1 U19484 ( .A(n16255), .B(n16254), .ZN(n16514) );
  NAND2_X1 U19485 ( .A1(n16258), .A2(n16257), .ZN(n16503) );
  NAND3_X1 U19486 ( .A1(n10029), .A2(n19577), .A3(n16503), .ZN(n16263) );
  NAND2_X1 U19487 ( .A1(n19571), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n16504) );
  NAND2_X1 U19488 ( .A1(n19584), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16259) );
  OAI211_X1 U19489 ( .C1(n19582), .C2(n16260), .A(n16504), .B(n16259), .ZN(
        n16261) );
  AOI21_X1 U19490 ( .B1(n16511), .B2(n19592), .A(n16261), .ZN(n16262) );
  OAI211_X1 U19491 ( .C1(n16514), .C2(n19574), .A(n16263), .B(n16262), .ZN(
        P2_U2992) );
  INV_X1 U19492 ( .A(n16264), .ZN(n16267) );
  OAI21_X1 U19493 ( .B1(n16267), .B2(n16266), .A(n16265), .ZN(n16272) );
  INV_X1 U19494 ( .A(n16268), .ZN(n16269) );
  NOR2_X1 U19495 ( .A1(n16270), .A2(n16269), .ZN(n16271) );
  XNOR2_X1 U19496 ( .A(n16272), .B(n16271), .ZN(n16532) );
  INV_X1 U19497 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16523) );
  NAND2_X1 U19498 ( .A1(n19571), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n16521) );
  OAI21_X1 U19499 ( .B1(n17198), .B2(n16274), .A(n16521), .ZN(n16275) );
  AOI21_X1 U19500 ( .B1(n17192), .B2(n16276), .A(n16275), .ZN(n16277) );
  OAI21_X1 U19501 ( .B1(n16528), .B2(n19573), .A(n16277), .ZN(n16278) );
  AOI21_X1 U19502 ( .B1(n16530), .B2(n19577), .A(n16278), .ZN(n16279) );
  OAI21_X1 U19503 ( .B1(n16281), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n16280), .ZN(n16557) );
  NAND2_X1 U19504 ( .A1(n11536), .A2(n16282), .ZN(n16284) );
  XOR2_X1 U19505 ( .A(n16284), .B(n16283), .Z(n16555) );
  NOR2_X1 U19506 ( .A1(n17200), .A2(n20237), .ZN(n16545) );
  NOR2_X1 U19507 ( .A1(n16285), .A2(n19582), .ZN(n16286) );
  AOI211_X1 U19508 ( .C1(n19584), .C2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16545), .B(n16286), .ZN(n16287) );
  OAI21_X1 U19509 ( .B1(n16553), .B2(n19573), .A(n16287), .ZN(n16288) );
  AOI21_X1 U19510 ( .B1(n16555), .B2(n9627), .A(n16288), .ZN(n16289) );
  OAI21_X1 U19511 ( .B1(n19590), .B2(n16557), .A(n16289), .ZN(P2_U2996) );
  OAI21_X1 U19512 ( .B1(n16291), .B2(n16290), .A(n11495), .ZN(n16579) );
  NAND2_X1 U19513 ( .A1(n19571), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n16577) );
  NAND2_X1 U19514 ( .A1(n19584), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16292) );
  OAI211_X1 U19515 ( .C1(n16293), .C2(n19582), .A(n16577), .B(n16292), .ZN(
        n16294) );
  AOI21_X1 U19516 ( .B1(n16582), .B2(n19592), .A(n16294), .ZN(n16298) );
  INV_X1 U19517 ( .A(n16299), .ZN(n16570) );
  INV_X1 U19518 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16586) );
  OAI21_X1 U19519 ( .B1(n16570), .B2(n16590), .A(n16586), .ZN(n16296) );
  NAND3_X1 U19520 ( .A1(n16296), .A2(n19577), .A3(n16558), .ZN(n16297) );
  OAI211_X1 U19521 ( .C1(n16579), .C2(n19574), .A(n16298), .B(n16297), .ZN(
        P2_U2998) );
  XNOR2_X1 U19522 ( .A(n16299), .B(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16600) );
  NAND2_X1 U19523 ( .A1(n16301), .A2(n16300), .ZN(n16303) );
  XOR2_X1 U19524 ( .A(n16303), .B(n16302), .Z(n16598) );
  INV_X1 U19525 ( .A(n16304), .ZN(n19399) );
  INV_X1 U19526 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n19390) );
  NAND2_X1 U19527 ( .A1(n19571), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n16593) );
  OAI21_X1 U19528 ( .B1(n17198), .B2(n19390), .A(n16593), .ZN(n16305) );
  AOI21_X1 U19529 ( .B1(n17192), .B2(n19399), .A(n16305), .ZN(n16306) );
  OAI21_X1 U19530 ( .B1(n19382), .B2(n19573), .A(n16306), .ZN(n16307) );
  AOI21_X1 U19531 ( .B1(n16598), .B2(n9627), .A(n16307), .ZN(n16308) );
  OAI21_X1 U19532 ( .B1(n19590), .B2(n16600), .A(n16308), .ZN(P2_U2999) );
  INV_X1 U19533 ( .A(n16310), .ZN(n16602) );
  OAI21_X1 U19534 ( .B1(n16325), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n16570), .ZN(n16613) );
  NAND2_X1 U19535 ( .A1(n16312), .A2(n16311), .ZN(n16313) );
  XNOR2_X1 U19536 ( .A(n16314), .B(n16313), .ZN(n16611) );
  INV_X1 U19537 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n20230) );
  NOR2_X1 U19538 ( .A1(n17200), .A2(n20230), .ZN(n16605) );
  NOR2_X1 U19539 ( .A1(n19582), .A2(n16315), .ZN(n16316) );
  AOI211_X1 U19540 ( .C1(n19584), .C2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16605), .B(n16316), .ZN(n16317) );
  OAI21_X1 U19541 ( .B1(n16608), .B2(n19573), .A(n16317), .ZN(n16318) );
  AOI21_X1 U19542 ( .B1(n16611), .B2(n9627), .A(n16318), .ZN(n16319) );
  OAI21_X1 U19543 ( .B1(n16613), .B2(n19590), .A(n16319), .ZN(P2_U3000) );
  NAND2_X1 U19544 ( .A1(n16321), .A2(n16320), .ZN(n16322) );
  XNOR2_X1 U19545 ( .A(n16323), .B(n16322), .ZN(n16624) );
  INV_X1 U19546 ( .A(n16309), .ZN(n16324) );
  NAND2_X1 U19547 ( .A1(n17192), .A2(n16326), .ZN(n16327) );
  NAND2_X1 U19548 ( .A1(n19571), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n16615) );
  OAI211_X1 U19549 ( .C1(n17198), .C2(n16328), .A(n16327), .B(n16615), .ZN(
        n16329) );
  AOI21_X1 U19550 ( .B1(n16621), .B2(n19592), .A(n16329), .ZN(n16330) );
  XNOR2_X1 U19551 ( .A(n16309), .B(n16627), .ZN(n16636) );
  INV_X1 U19552 ( .A(n16331), .ZN(n16332) );
  NOR2_X1 U19553 ( .A1(n16333), .A2(n16332), .ZN(n16334) );
  XOR2_X1 U19554 ( .A(n16334), .B(n9716), .Z(n16633) );
  NAND2_X1 U19555 ( .A1(n16625), .A2(n19592), .ZN(n16336) );
  NOR2_X1 U19556 ( .A1(n17200), .A2(n20226), .ZN(n16626) );
  AOI21_X1 U19557 ( .B1(n19584), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16626), .ZN(n16335) );
  OAI211_X1 U19558 ( .C1(n19582), .C2(n16337), .A(n16336), .B(n16335), .ZN(
        n16338) );
  AOI21_X1 U19559 ( .B1(n16633), .B2(n9627), .A(n16338), .ZN(n16339) );
  OAI21_X1 U19560 ( .B1(n16636), .B2(n19590), .A(n16339), .ZN(P2_U3002) );
  OAI21_X1 U19561 ( .B1(n11474), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n16309), .ZN(n16647) );
  XNOR2_X1 U19562 ( .A(n16340), .B(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16341) );
  XNOR2_X1 U19563 ( .A(n16342), .B(n16341), .ZN(n16645) );
  NOR2_X1 U19564 ( .A1(n17200), .A2(n16343), .ZN(n16640) );
  NOR2_X1 U19565 ( .A1(n17198), .A2(n16344), .ZN(n16345) );
  AOI211_X1 U19566 ( .C1(n16346), .C2(n17192), .A(n16640), .B(n16345), .ZN(
        n16347) );
  OAI21_X1 U19567 ( .B1(n16643), .B2(n19573), .A(n16347), .ZN(n16348) );
  AOI21_X1 U19568 ( .B1(n16645), .B2(n9627), .A(n16348), .ZN(n16349) );
  OAI21_X1 U19569 ( .B1(n16647), .B2(n19590), .A(n16349), .ZN(P2_U3003) );
  NOR2_X1 U19570 ( .A1(n16350), .A2(n16665), .ZN(n16352) );
  OAI21_X1 U19571 ( .B1(n16352), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n16351), .ZN(n16659) );
  NAND2_X1 U19572 ( .A1(n16353), .A2(n16364), .ZN(n16358) );
  INV_X1 U19573 ( .A(n16354), .ZN(n16356) );
  NAND2_X1 U19574 ( .A1(n16356), .A2(n16355), .ZN(n16357) );
  XNOR2_X1 U19575 ( .A(n16358), .B(n16357), .ZN(n16657) );
  NOR2_X1 U19576 ( .A1(n17200), .A2(n20223), .ZN(n16651) );
  NOR2_X1 U19577 ( .A1(n19582), .A2(n16359), .ZN(n16360) );
  AOI211_X1 U19578 ( .C1(n19584), .C2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16651), .B(n16360), .ZN(n16361) );
  OAI21_X1 U19579 ( .B1(n16655), .B2(n19573), .A(n16361), .ZN(n16362) );
  AOI21_X1 U19580 ( .B1(n16657), .B2(n9627), .A(n16362), .ZN(n16363) );
  OAI21_X1 U19581 ( .B1(n16659), .B2(n19590), .A(n16363), .ZN(P2_U3004) );
  XNOR2_X1 U19582 ( .A(n11476), .B(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16670) );
  NAND2_X1 U19583 ( .A1(n16365), .A2(n16364), .ZN(n16366) );
  XNOR2_X1 U19584 ( .A(n16367), .B(n16366), .ZN(n16668) );
  NAND2_X1 U19585 ( .A1(n19571), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n16660) );
  OAI21_X1 U19586 ( .B1(n17198), .B2(n16368), .A(n16660), .ZN(n16369) );
  AOI21_X1 U19587 ( .B1(n17192), .B2(n16370), .A(n16369), .ZN(n16371) );
  OAI21_X1 U19588 ( .B1(n16372), .B2(n19573), .A(n16371), .ZN(n16373) );
  AOI21_X1 U19589 ( .B1(n16668), .B2(n9627), .A(n16373), .ZN(n16374) );
  OAI21_X1 U19590 ( .B1(n16670), .B2(n19590), .A(n16374), .ZN(P2_U3005) );
  XNOR2_X1 U19591 ( .A(n16375), .B(n16376), .ZN(n16685) );
  AOI21_X1 U19592 ( .B1(n16379), .B2(n16378), .A(n16377), .ZN(n16380) );
  XNOR2_X1 U19593 ( .A(n16380), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16407) );
  INV_X1 U19594 ( .A(n16380), .ZN(n16381) );
  AOI22_X1 U19595 ( .A1(n16407), .A2(n16408), .B1(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16381), .ZN(n16397) );
  INV_X1 U19596 ( .A(n16396), .ZN(n16382) );
  OAI21_X1 U19597 ( .B1(n16397), .B2(n16382), .A(n16395), .ZN(n16386) );
  NAND2_X1 U19598 ( .A1(n16384), .A2(n16383), .ZN(n16385) );
  XNOR2_X1 U19599 ( .A(n16386), .B(n16385), .ZN(n16683) );
  NOR2_X1 U19600 ( .A1(n17200), .A2(n20219), .ZN(n16677) );
  NOR2_X1 U19601 ( .A1(n19582), .A2(n16387), .ZN(n16388) );
  AOI211_X1 U19602 ( .C1(n19584), .C2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16677), .B(n16388), .ZN(n16389) );
  OAI21_X1 U19603 ( .B1(n16681), .B2(n19573), .A(n16389), .ZN(n16390) );
  AOI21_X1 U19604 ( .B1(n16683), .B2(n9627), .A(n16390), .ZN(n16391) );
  OAI21_X1 U19605 ( .B1(n16685), .B2(n19590), .A(n16391), .ZN(P2_U3006) );
  XNOR2_X1 U19606 ( .A(n16392), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16393) );
  XNOR2_X1 U19607 ( .A(n16394), .B(n16393), .ZN(n16696) );
  NAND2_X1 U19608 ( .A1(n16396), .A2(n16395), .ZN(n16398) );
  XOR2_X1 U19609 ( .A(n16398), .B(n16397), .Z(n16686) );
  NAND2_X1 U19610 ( .A1(n19571), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n16690) );
  OAI21_X1 U19611 ( .B1(n17198), .B2(n16399), .A(n16690), .ZN(n16400) );
  AOI21_X1 U19612 ( .B1(n17192), .B2(n16401), .A(n16400), .ZN(n16402) );
  OAI21_X1 U19613 ( .B1(n16691), .B2(n19573), .A(n16402), .ZN(n16403) );
  AOI21_X1 U19614 ( .B1(n16686), .B2(n9627), .A(n16403), .ZN(n16404) );
  OAI21_X1 U19615 ( .B1(n19590), .B2(n16696), .A(n16404), .ZN(P2_U3007) );
  OAI21_X1 U19616 ( .B1(n16405), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n16406), .ZN(n16708) );
  XOR2_X1 U19617 ( .A(n16408), .B(n16407), .Z(n16706) );
  INV_X1 U19618 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n20215) );
  OAI22_X1 U19619 ( .A1(n20215), .A2(n17200), .B1(n19582), .B2(n16409), .ZN(
        n16410) );
  AOI21_X1 U19620 ( .B1(n19584), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16410), .ZN(n16411) );
  OAI21_X1 U19621 ( .B1(n16698), .B2(n19573), .A(n16411), .ZN(n16412) );
  AOI21_X1 U19622 ( .B1(n16706), .B2(n9627), .A(n16412), .ZN(n16413) );
  OAI21_X1 U19623 ( .B1(n19590), .B2(n16708), .A(n16413), .ZN(P2_U3008) );
  XOR2_X1 U19624 ( .A(n16414), .B(n16415), .Z(n17210) );
  NAND2_X1 U19625 ( .A1(n17210), .A2(n19577), .ZN(n16424) );
  NOR2_X1 U19626 ( .A1(n16417), .A2(n16416), .ZN(n16418) );
  XNOR2_X1 U19627 ( .A(n16419), .B(n16418), .ZN(n17205) );
  NOR2_X1 U19628 ( .A1(n19582), .A2(n10182), .ZN(n16422) );
  OAI22_X1 U19629 ( .A1(n17198), .A2(n16420), .B1(n17201), .B2(n17200), .ZN(
        n16421) );
  AOI211_X1 U19630 ( .C1(n17205), .C2(n9627), .A(n16422), .B(n16421), .ZN(
        n16423) );
  OAI211_X1 U19631 ( .C1(n19573), .C2(n17207), .A(n16424), .B(n16423), .ZN(
        P2_U3011) );
  OAI21_X1 U19632 ( .B1(n16426), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n16425), .ZN(n16427) );
  AOI21_X1 U19633 ( .B1(n16428), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n16427), .ZN(n16429) );
  OAI21_X1 U19634 ( .B1(n16430), .B2(n17203), .A(n16429), .ZN(n16431) );
  AOI21_X1 U19635 ( .B1(n16432), .B2(n16745), .A(n16431), .ZN(n16435) );
  NAND2_X1 U19636 ( .A1(n16433), .A2(n17209), .ZN(n16434) );
  OAI211_X1 U19637 ( .C1(n16436), .C2(n16737), .A(n16435), .B(n16434), .ZN(
        P2_U3017) );
  NAND2_X1 U19638 ( .A1(n16437), .A2(n16745), .ZN(n16445) );
  NAND2_X1 U19639 ( .A1(n16439), .A2(n16438), .ZN(n16441) );
  NAND2_X1 U19640 ( .A1(n16441), .A2(n16440), .ZN(n16442) );
  AOI21_X1 U19641 ( .B1(n16443), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n16442), .ZN(n16444) );
  OAI211_X1 U19642 ( .C1(n17203), .C2(n16446), .A(n16445), .B(n16444), .ZN(
        n16447) );
  AOI21_X1 U19643 ( .B1(n17209), .B2(n16448), .A(n16447), .ZN(n16449) );
  OAI21_X1 U19644 ( .B1(n16450), .B2(n16737), .A(n16449), .ZN(P2_U3019) );
  INV_X1 U19645 ( .A(n16451), .ZN(n16453) );
  NAND2_X1 U19646 ( .A1(n16456), .A2(n16468), .ZN(n16452) );
  NAND3_X1 U19647 ( .A1(n16465), .A2(n16453), .A3(n16452), .ZN(n16454) );
  OAI211_X1 U19648 ( .C1(n16469), .C2(n16456), .A(n16455), .B(n16454), .ZN(
        n16457) );
  AOI21_X1 U19649 ( .B1(n16458), .B2(n17215), .A(n16457), .ZN(n16459) );
  OAI21_X1 U19650 ( .B1(n16460), .B2(n17227), .A(n16459), .ZN(n16461) );
  AOI21_X1 U19651 ( .B1(n16462), .B2(n17224), .A(n16461), .ZN(n16463) );
  OAI21_X1 U19652 ( .B1(n17226), .B2(n16464), .A(n16463), .ZN(P2_U3020) );
  NAND2_X1 U19653 ( .A1(n16465), .A2(n16468), .ZN(n16466) );
  OAI211_X1 U19654 ( .C1(n16469), .C2(n16468), .A(n16467), .B(n16466), .ZN(
        n16472) );
  NOR2_X1 U19655 ( .A1(n16470), .A2(n17203), .ZN(n16471) );
  AOI211_X1 U19656 ( .C1(n16473), .C2(n16745), .A(n16472), .B(n16471), .ZN(
        n16477) );
  NAND3_X1 U19657 ( .A1(n16475), .A2(n17209), .A3(n16474), .ZN(n16476) );
  OAI211_X1 U19658 ( .C1(n16478), .C2(n16737), .A(n16477), .B(n16476), .ZN(
        P2_U3021) );
  NAND2_X1 U19659 ( .A1(n16479), .A2(n17215), .ZN(n16486) );
  OAI21_X1 U19660 ( .B1(n16494), .B2(n16481), .A(n16480), .ZN(n16483) );
  AOI21_X1 U19661 ( .B1(n16484), .B2(n16483), .A(n16482), .ZN(n16485) );
  OAI211_X1 U19662 ( .C1(n16487), .C2(n17227), .A(n16486), .B(n16485), .ZN(
        n16488) );
  AOI21_X1 U19663 ( .B1(n16489), .B2(n17224), .A(n16488), .ZN(n16490) );
  OAI21_X1 U19664 ( .B1(n17226), .B2(n16491), .A(n16490), .ZN(P2_U3022) );
  NOR3_X1 U19665 ( .A1(n16649), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n16517), .ZN(n16506) );
  OAI21_X1 U19666 ( .B1(n16507), .B2(n16506), .A(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16493) );
  OAI211_X1 U19667 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n16494), .A(
        n16493), .B(n16492), .ZN(n16497) );
  NOR2_X1 U19668 ( .A1(n16495), .A2(n17227), .ZN(n16496) );
  AOI211_X1 U19669 ( .C1(n17215), .C2(n16498), .A(n16497), .B(n16496), .ZN(
        n16501) );
  NAND3_X1 U19670 ( .A1(n16499), .A2(n16250), .A3(n17224), .ZN(n16500) );
  OAI211_X1 U19671 ( .C1(n16502), .C2(n17226), .A(n16501), .B(n16500), .ZN(
        P2_U3023) );
  NAND3_X1 U19672 ( .A1(n10029), .A2(n17209), .A3(n16503), .ZN(n16513) );
  INV_X1 U19673 ( .A(n16504), .ZN(n16505) );
  AOI211_X1 U19674 ( .C1(n16507), .C2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n16506), .B(n16505), .ZN(n16508) );
  OAI21_X1 U19675 ( .B1(n16509), .B2(n17203), .A(n16508), .ZN(n16510) );
  AOI21_X1 U19676 ( .B1(n16511), .B2(n16745), .A(n16510), .ZN(n16512) );
  OAI211_X1 U19677 ( .C1(n16514), .C2(n16737), .A(n16513), .B(n16512), .ZN(
        P2_U3024) );
  OAI21_X1 U19678 ( .B1(n16519), .B2(n16515), .A(n16666), .ZN(n16516) );
  AOI21_X1 U19679 ( .B1(n16518), .B2(n16517), .A(n16516), .ZN(n16524) );
  INV_X1 U19680 ( .A(n16649), .ZN(n16520) );
  NAND3_X1 U19681 ( .A1(n16520), .A2(n16519), .A3(n16523), .ZN(n16522) );
  OAI211_X1 U19682 ( .C1(n16524), .C2(n16523), .A(n16522), .B(n16521), .ZN(
        n16525) );
  AOI21_X1 U19683 ( .B1(n16526), .B2(n17215), .A(n16525), .ZN(n16527) );
  OAI21_X1 U19684 ( .B1(n16528), .B2(n17227), .A(n16527), .ZN(n16529) );
  AOI21_X1 U19685 ( .B1(n16530), .B2(n17209), .A(n16529), .ZN(n16531) );
  OAI21_X1 U19686 ( .B1(n16532), .B2(n16737), .A(n16531), .ZN(P2_U3025) );
  NAND2_X1 U19687 ( .A1(n16533), .A2(n16745), .ZN(n16540) );
  XNOR2_X1 U19688 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16535) );
  NOR2_X1 U19689 ( .A1(n16535), .A2(n16534), .ZN(n16536) );
  AOI211_X1 U19690 ( .C1(n16538), .C2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n16537), .B(n16536), .ZN(n16539) );
  OAI211_X1 U19691 ( .C1(n17203), .C2(n16541), .A(n16540), .B(n16539), .ZN(
        n16542) );
  OAI21_X1 U19692 ( .B1(n17226), .B2(n16544), .A(n16543), .ZN(P2_U3026) );
  INV_X1 U19693 ( .A(n16545), .ZN(n16546) );
  OAI211_X1 U19694 ( .C1(n16549), .C2(n16548), .A(n16547), .B(n16546), .ZN(
        n16550) );
  AOI21_X1 U19695 ( .B1(n17215), .B2(n16551), .A(n16550), .ZN(n16552) );
  OAI21_X1 U19696 ( .B1(n17227), .B2(n16553), .A(n16552), .ZN(n16554) );
  AOI21_X1 U19697 ( .B1(n16555), .B2(n17224), .A(n16554), .ZN(n16556) );
  OAI21_X1 U19698 ( .B1(n17226), .B2(n16557), .A(n16556), .ZN(P2_U3028) );
  OAI21_X1 U19699 ( .B1(n17209), .B2(n16559), .A(n16558), .ZN(n16561) );
  INV_X1 U19700 ( .A(n16595), .ZN(n16560) );
  OAI211_X1 U19701 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n16562), .A(
        n16561), .B(n16560), .ZN(n16576) );
  AOI21_X1 U19702 ( .B1(n16586), .B2(n16750), .A(n16576), .ZN(n16575) );
  NAND2_X1 U19703 ( .A1(n16563), .A2(n17215), .ZN(n16564) );
  OAI211_X1 U19704 ( .C1(n16566), .C2(n17227), .A(n16565), .B(n16564), .ZN(
        n16567) );
  AOI21_X1 U19705 ( .B1(n16568), .B2(n17224), .A(n16567), .ZN(n16573) );
  INV_X1 U19706 ( .A(n16591), .ZN(n16569) );
  OAI21_X1 U19707 ( .B1(n16570), .B2(n17226), .A(n16569), .ZN(n16583) );
  NAND3_X1 U19708 ( .A1(n16583), .A2(n16571), .A3(n16574), .ZN(n16572) );
  OAI211_X1 U19709 ( .C1(n16575), .C2(n16574), .A(n16573), .B(n16572), .ZN(
        P2_U3029) );
  INV_X1 U19710 ( .A(n16576), .ZN(n16587) );
  OAI21_X1 U19711 ( .B1(n16578), .B2(n17203), .A(n16577), .ZN(n16581) );
  NOR2_X1 U19712 ( .A1(n16579), .A2(n16737), .ZN(n16580) );
  AOI211_X1 U19713 ( .C1(n16745), .C2(n16582), .A(n16581), .B(n16580), .ZN(
        n16585) );
  NAND3_X1 U19714 ( .A1(n16583), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        n16586), .ZN(n16584) );
  OAI211_X1 U19715 ( .C1(n16587), .C2(n16586), .A(n16585), .B(n16584), .ZN(
        P2_U3030) );
  INV_X1 U19716 ( .A(n15779), .ZN(n16588) );
  OAI21_X1 U19717 ( .B1(n9665), .B2(n16589), .A(n16588), .ZN(n19383) );
  NAND2_X1 U19718 ( .A1(n16591), .A2(n16590), .ZN(n16592) );
  OAI211_X1 U19719 ( .C1(n19383), .C2(n17203), .A(n16593), .B(n16592), .ZN(
        n16594) );
  AOI21_X1 U19720 ( .B1(n16595), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n16594), .ZN(n16596) );
  OAI21_X1 U19721 ( .B1(n17227), .B2(n19382), .A(n16596), .ZN(n16597) );
  AOI21_X1 U19722 ( .B1(n16598), .B2(n17224), .A(n16597), .ZN(n16599) );
  OAI21_X1 U19723 ( .B1(n17226), .B2(n16600), .A(n16599), .ZN(P2_U3031) );
  INV_X1 U19724 ( .A(n16603), .ZN(n16628) );
  AOI21_X1 U19725 ( .B1(n16628), .B2(n16602), .A(n16638), .ZN(n16618) );
  NOR2_X1 U19726 ( .A1(n16618), .A2(n16601), .ZN(n16610) );
  NOR3_X1 U19727 ( .A1(n16603), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n16602), .ZN(n16604) );
  AOI211_X1 U19728 ( .C1(n16606), .C2(n17215), .A(n16605), .B(n16604), .ZN(
        n16607) );
  OAI21_X1 U19729 ( .B1(n17227), .B2(n16608), .A(n16607), .ZN(n16609) );
  AOI211_X1 U19730 ( .C1(n16611), .C2(n17224), .A(n16610), .B(n16609), .ZN(
        n16612) );
  OAI21_X1 U19731 ( .B1(n16613), .B2(n17226), .A(n16612), .ZN(P2_U3032) );
  NAND2_X1 U19732 ( .A1(n16614), .A2(n17209), .ZN(n16623) );
  OAI21_X1 U19733 ( .B1(n16616), .B2(n17203), .A(n16615), .ZN(n16620) );
  AOI21_X1 U19734 ( .B1(n16628), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16617) );
  NOR2_X1 U19735 ( .A1(n16618), .A2(n16617), .ZN(n16619) );
  AOI211_X1 U19736 ( .C1(n16745), .C2(n16621), .A(n16620), .B(n16619), .ZN(
        n16622) );
  OAI211_X1 U19737 ( .C1(n16624), .C2(n16737), .A(n16623), .B(n16622), .ZN(
        P2_U3033) );
  NAND2_X1 U19738 ( .A1(n16625), .A2(n16745), .ZN(n16630) );
  AOI21_X1 U19739 ( .B1(n16628), .B2(n16627), .A(n16626), .ZN(n16629) );
  OAI211_X1 U19740 ( .C1(n17203), .C2(n16631), .A(n16630), .B(n16629), .ZN(
        n16632) );
  AOI21_X1 U19741 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16638), .A(
        n16632), .ZN(n16635) );
  NAND2_X1 U19742 ( .A1(n16633), .A2(n17224), .ZN(n16634) );
  OAI211_X1 U19743 ( .C1(n16636), .C2(n17226), .A(n16635), .B(n16634), .ZN(
        P2_U3034) );
  NOR2_X1 U19744 ( .A1(n16649), .A2(n16637), .ZN(n16639) );
  OAI21_X1 U19745 ( .B1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16639), .A(
        n16638), .ZN(n16642) );
  AOI21_X1 U19746 ( .B1(n19436), .B2(n17215), .A(n16640), .ZN(n16641) );
  OAI211_X1 U19747 ( .C1(n16643), .C2(n17227), .A(n16642), .B(n16641), .ZN(
        n16644) );
  AOI21_X1 U19748 ( .B1(n16645), .B2(n17224), .A(n16644), .ZN(n16646) );
  OAI21_X1 U19749 ( .B1(n16647), .B2(n17226), .A(n16646), .ZN(P2_U3035) );
  NAND2_X1 U19750 ( .A1(n16648), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16654) );
  NOR3_X1 U19751 ( .A1(n16649), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n16665), .ZN(n16650) );
  AOI211_X1 U19752 ( .C1(n17215), .C2(n16652), .A(n16651), .B(n16650), .ZN(
        n16653) );
  OAI211_X1 U19753 ( .C1(n16655), .C2(n17227), .A(n16654), .B(n16653), .ZN(
        n16656) );
  AOI21_X1 U19754 ( .B1(n16657), .B2(n17224), .A(n16656), .ZN(n16658) );
  OAI21_X1 U19755 ( .B1(n16659), .B2(n17226), .A(n16658), .ZN(P2_U3036) );
  OAI211_X1 U19756 ( .C1(n19442), .C2(n17203), .A(n16661), .B(n16660), .ZN(
        n16662) );
  AOI21_X1 U19757 ( .B1(n16663), .B2(n16745), .A(n16662), .ZN(n16664) );
  OAI21_X1 U19758 ( .B1(n16666), .B2(n16665), .A(n16664), .ZN(n16667) );
  AOI21_X1 U19759 ( .B1(n17224), .B2(n16668), .A(n16667), .ZN(n16669) );
  OAI21_X1 U19760 ( .B1(n16670), .B2(n17226), .A(n16669), .ZN(P2_U3037) );
  AND2_X1 U19761 ( .A1(n16672), .A2(n16671), .ZN(n16697) );
  NAND2_X1 U19762 ( .A1(n16697), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16680) );
  OAI211_X1 U19763 ( .C1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16674), .B(n16673), .ZN(n16675) );
  NOR2_X1 U19764 ( .A1(n17214), .A2(n16675), .ZN(n16676) );
  AOI211_X1 U19765 ( .C1(n16678), .C2(n17215), .A(n16677), .B(n16676), .ZN(
        n16679) );
  OAI211_X1 U19766 ( .C1(n16681), .C2(n17227), .A(n16680), .B(n16679), .ZN(
        n16682) );
  AOI21_X1 U19767 ( .B1(n16683), .B2(n17224), .A(n16682), .ZN(n16684) );
  OAI21_X1 U19768 ( .B1(n16685), .B2(n17226), .A(n16684), .ZN(P2_U3038) );
  NAND2_X1 U19769 ( .A1(n16686), .A2(n17224), .ZN(n16695) );
  NOR2_X1 U19770 ( .A1(n16687), .A2(n17203), .ZN(n16693) );
  NAND2_X1 U19771 ( .A1(n16688), .A2(n11074), .ZN(n16689) );
  OAI211_X1 U19772 ( .C1(n16691), .C2(n17227), .A(n16690), .B(n16689), .ZN(
        n16692) );
  AOI211_X1 U19773 ( .C1(n16697), .C2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n16693), .B(n16692), .ZN(n16694) );
  OAI211_X1 U19774 ( .C1(n16696), .C2(n17226), .A(n16695), .B(n16694), .ZN(
        P2_U3039) );
  INV_X1 U19775 ( .A(n16697), .ZN(n16704) );
  INV_X1 U19776 ( .A(n16698), .ZN(n16702) );
  OAI22_X1 U19777 ( .A1(n19446), .A2(n17203), .B1(n20215), .B2(n17200), .ZN(
        n16701) );
  NOR3_X1 U19778 ( .A1(n17214), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        n16699), .ZN(n16700) );
  AOI211_X1 U19779 ( .C1(n16702), .C2(n16745), .A(n16701), .B(n16700), .ZN(
        n16703) );
  OAI21_X1 U19780 ( .B1(n16704), .B2(n21322), .A(n16703), .ZN(n16705) );
  AOI21_X1 U19781 ( .B1(n16706), .B2(n17224), .A(n16705), .ZN(n16707) );
  OAI21_X1 U19782 ( .B1(n17226), .B2(n16708), .A(n16707), .ZN(P2_U3040) );
  NAND2_X1 U19783 ( .A1(n16711), .A2(n16710), .ZN(n16712) );
  XNOR2_X1 U19784 ( .A(n16709), .B(n16712), .ZN(n17195) );
  INV_X1 U19785 ( .A(n17195), .ZN(n16723) );
  AOI21_X1 U19786 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n17212), .A(
        n16713), .ZN(n16738) );
  XOR2_X1 U19787 ( .A(n16715), .B(n16714), .Z(n17193) );
  NOR2_X1 U19788 ( .A1(n17213), .A2(n17214), .ZN(n16739) );
  OAI221_X1 U19789 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C1(n16726), .C2(n11066), .A(
        n16739), .ZN(n16717) );
  NAND2_X1 U19790 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19571), .ZN(n16716) );
  OAI211_X1 U19791 ( .C1(n19449), .C2(n17203), .A(n16717), .B(n16716), .ZN(
        n16718) );
  AOI21_X1 U19792 ( .B1(n17224), .B2(n17193), .A(n16718), .ZN(n16719) );
  OAI21_X1 U19793 ( .B1(n16720), .B2(n17227), .A(n16719), .ZN(n16721) );
  AOI21_X1 U19794 ( .B1(n16738), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n16721), .ZN(n16722) );
  OAI21_X1 U19795 ( .B1(n16723), .B2(n17226), .A(n16722), .ZN(P2_U3041) );
  XNOR2_X1 U19796 ( .A(n16725), .B(n16726), .ZN(n16727) );
  XNOR2_X1 U19797 ( .A(n16724), .B(n16727), .ZN(n19578) );
  OAI21_X1 U19798 ( .B1(n16730), .B2(n16729), .A(n16728), .ZN(n19575) );
  NAND2_X1 U19799 ( .A1(n16732), .A2(n16731), .ZN(n16733) );
  NAND2_X1 U19800 ( .A1(n14243), .A2(n16733), .ZN(n19572) );
  INV_X1 U19801 ( .A(n19572), .ZN(n19425) );
  NOR2_X1 U19802 ( .A1(n11300), .A2(n17200), .ZN(n16735) );
  NOR2_X1 U19803 ( .A1(n19408), .A2(n17203), .ZN(n16734) );
  AOI211_X1 U19804 ( .C1(n19425), .C2(n16745), .A(n16735), .B(n16734), .ZN(
        n16736) );
  OAI21_X1 U19805 ( .B1(n19575), .B2(n16737), .A(n16736), .ZN(n16741) );
  MUX2_X1 U19806 ( .A(n16739), .B(n16738), .S(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(n16740) );
  AOI211_X1 U19807 ( .C1(n19578), .C2(n17209), .A(n16741), .B(n16740), .ZN(
        n16742) );
  INV_X1 U19808 ( .A(n16742), .ZN(P2_U3042) );
  OAI22_X1 U19809 ( .A1(n16759), .A2(n17203), .B1(n17226), .B2(n16743), .ZN(
        n16744) );
  AOI21_X1 U19810 ( .B1(n16746), .B2(n16745), .A(n16744), .ZN(n16754) );
  AOI21_X1 U19811 ( .B1(n17224), .B2(n16748), .A(n16747), .ZN(n16753) );
  NAND2_X1 U19812 ( .A1(n17216), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16752) );
  OAI211_X1 U19813 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n16750), .B(n16749), .ZN(n16751) );
  NAND4_X1 U19814 ( .A1(n16754), .A2(n16753), .A3(n16752), .A4(n16751), .ZN(
        P2_U3045) );
  INV_X1 U19815 ( .A(n16755), .ZN(n16756) );
  NAND2_X1 U19816 ( .A1(n20276), .A2(n16756), .ZN(n16757) );
  NAND2_X1 U19817 ( .A1(n20305), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20270) );
  MUX2_X1 U19818 ( .A(n16757), .B(n20270), .S(n20275), .Z(n16758) );
  OAI21_X1 U19819 ( .B1(n16759), .B2(n20306), .A(n16758), .ZN(n16760) );
  MUX2_X1 U19820 ( .A(n16760), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        n20294), .Z(P2_U3604) );
  INV_X1 U19821 ( .A(n16773), .ZN(n16762) );
  MUX2_X1 U19822 ( .A(n17217), .B(n16762), .S(n16761), .Z(n16769) );
  INV_X1 U19823 ( .A(n10953), .ZN(n16764) );
  NAND2_X1 U19824 ( .A1(n16764), .A2(n16763), .ZN(n16779) );
  INV_X1 U19825 ( .A(n16779), .ZN(n16766) );
  MUX2_X1 U19826 ( .A(n16766), .B(n16765), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n16767) );
  OAI21_X1 U19827 ( .B1(n11577), .B2(n16795), .A(n16767), .ZN(n16840) );
  AOI222_X1 U19828 ( .A1(n16769), .A2(P2_STATE2_REG_1__SCAN_IN), .B1(n16768), 
        .B2(n17239), .C1(n16840), .C2(n20273), .ZN(n16771) );
  NAND2_X1 U19829 ( .A1(n16802), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n16770) );
  OAI21_X1 U19830 ( .B1(n16771), .B2(n16802), .A(n16770), .ZN(P2_U3601) );
  NAND2_X1 U19831 ( .A1(n19416), .A2(n17217), .ZN(n16772) );
  OAI211_X1 U19832 ( .C1(n19416), .C2(n16773), .A(P2_STATE2_REG_1__SCAN_IN), 
        .B(n16772), .ZN(n16798) );
  NAND2_X1 U19833 ( .A1(n19416), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16774) );
  INV_X1 U19834 ( .A(n16797), .ZN(n16782) );
  INV_X1 U19835 ( .A(n20273), .ZN(n16801) );
  OR2_X1 U19836 ( .A1(n11572), .A2(n16795), .ZN(n16781) );
  INV_X1 U19837 ( .A(n10446), .ZN(n16777) );
  NAND2_X1 U19838 ( .A1(n16777), .A2(n16776), .ZN(n16778) );
  AOI22_X1 U19839 ( .A1(n16779), .A2(n16778), .B1(n16787), .B2(n10255), .ZN(
        n16780) );
  AND2_X1 U19840 ( .A1(n16781), .A2(n16780), .ZN(n16837) );
  INV_X1 U19841 ( .A(n17239), .ZN(n16799) );
  OAI222_X1 U19842 ( .A1(n16798), .A2(n16782), .B1(n16801), .B2(n16837), .C1(
        n16799), .C2(n20275), .ZN(n16783) );
  MUX2_X1 U19843 ( .A(n16783), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n16802), .Z(P2_U3600) );
  NAND2_X1 U19844 ( .A1(n9590), .A2(n16784), .ZN(n16790) );
  NOR2_X1 U19845 ( .A1(n16786), .A2(n16785), .ZN(n16788) );
  AOI22_X1 U19846 ( .A1(n16789), .A2(n16790), .B1(n16788), .B2(n16787), .ZN(
        n16794) );
  INV_X1 U19847 ( .A(n16790), .ZN(n16791) );
  NAND2_X1 U19848 ( .A1(n16792), .A2(n16791), .ZN(n16793) );
  OAI211_X1 U19849 ( .C1(n9613), .C2(n16795), .A(n16794), .B(n16793), .ZN(
        n16796) );
  INV_X1 U19850 ( .A(n16796), .ZN(n16833) );
  OAI222_X1 U19851 ( .A1(n20288), .A2(n16799), .B1(n16798), .B2(n16797), .C1(
        n16801), .C2(n16833), .ZN(n16800) );
  MUX2_X1 U19852 ( .A(n16800), .B(n10980), .S(n16802), .Z(P2_U3599) );
  NOR4_X1 U19853 ( .A1(n10857), .A2(n16852), .A3(n10884), .A4(n16801), .ZN(
        n16803) );
  MUX2_X1 U19854 ( .A(n16803), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n16802), .Z(P2_U3595) );
  INV_X1 U19855 ( .A(n20271), .ZN(n16804) );
  AOI21_X1 U19856 ( .B1(n19845), .B2(n16804), .A(n20268), .ZN(n16813) );
  INV_X1 U19857 ( .A(n16813), .ZN(n16807) );
  NOR2_X1 U19858 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19681) );
  NAND2_X1 U19859 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19681), .ZN(
        n16812) );
  INV_X1 U19860 ( .A(n19681), .ZN(n19683) );
  NOR2_X1 U19861 ( .A1(n19978), .A2(n19683), .ZN(n19732) );
  OAI21_X1 U19862 ( .B1(n16805), .B2(n19732), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n16806) );
  INV_X1 U19863 ( .A(n19734), .ZN(n16819) );
  INV_X2 U19864 ( .A(n19808), .ZN(n20133) );
  INV_X1 U19865 ( .A(n20127), .ZN(n16818) );
  AOI22_X1 U19866 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19639), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19638), .ZN(n20139) );
  INV_X1 U19867 ( .A(n20139), .ZN(n20047) );
  AOI22_X1 U19868 ( .A1(BUF2_REG_16__SCAN_IN), .A2(n19638), .B1(
        BUF1_REG_16__SCAN_IN), .B2(n19639), .ZN(n20084) );
  INV_X1 U19869 ( .A(n19732), .ZN(n19725) );
  NAND2_X1 U19870 ( .A1(n19644), .A2(n20311), .ZN(n20071) );
  OAI22_X1 U19871 ( .A1(n19718), .A2(n20084), .B1(n19725), .B2(n20071), .ZN(
        n16810) );
  AOI21_X1 U19872 ( .B1(n19733), .B2(n20047), .A(n16810), .ZN(n16817) );
  AOI21_X1 U19873 ( .B1(n16811), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n16815) );
  NAND2_X1 U19874 ( .A1(n16813), .A2(n16812), .ZN(n16814) );
  NAND2_X1 U19875 ( .A1(n19735), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n16816) );
  OAI211_X1 U19876 ( .C1(n16819), .C2(n16818), .A(n16817), .B(n16816), .ZN(
        P2_U3072) );
  OAI21_X1 U19877 ( .B1(n20065), .B2(n20031), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n16824) );
  INV_X1 U19878 ( .A(n19805), .ZN(n19739) );
  NAND3_X1 U19879 ( .A1(n19739), .A2(n19738), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n16825) );
  AND3_X1 U19880 ( .A1(n19911), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20040) );
  AND2_X1 U19881 ( .A1(n20040), .A2(n19682), .ZN(n20029) );
  OAI211_X1 U19882 ( .C1(n20029), .C2(n20306), .A(n16827), .B(n20133), .ZN(
        n16823) );
  INV_X1 U19883 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16832) );
  AOI22_X2 U19884 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19639), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19638), .ZN(n20171) );
  INV_X1 U19885 ( .A(n20171), .ZN(n20059) );
  AOI22_X1 U19886 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19639), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19638), .ZN(n20106) );
  INV_X1 U19887 ( .A(n20106), .ZN(n20166) );
  AOI22_X1 U19888 ( .A1(n20031), .A2(n20059), .B1(n20065), .B2(n20166), .ZN(
        n16831) );
  OAI21_X1 U19889 ( .B1(n16825), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20317), 
        .ZN(n16826) );
  AOI22_X1 U19890 ( .A1(n20030), .A2(n20165), .B1(n20029), .B2(n20164), .ZN(
        n16830) );
  OAI211_X1 U19891 ( .C1(n20035), .C2(n16832), .A(n16831), .B(n16830), .ZN(
        P2_U3149) );
  MUX2_X1 U19892 ( .A(n16834), .B(n16833), .S(n16836), .Z(n16863) );
  MUX2_X1 U19893 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n16835), .S(
        n16836), .Z(n16845) );
  INV_X1 U19894 ( .A(n16845), .ZN(n16862) );
  INV_X1 U19895 ( .A(n19978), .ZN(n19842) );
  AOI21_X1 U19896 ( .B1(n16837), .B2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        n19842), .ZN(n16841) );
  NAND2_X1 U19897 ( .A1(n16863), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n16839) );
  INV_X1 U19898 ( .A(n16836), .ZN(n16859) );
  AOI21_X1 U19899 ( .B1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n16837), .A(
        n16859), .ZN(n16838) );
  OAI211_X1 U19900 ( .C1(n16841), .C2(n16840), .A(n16839), .B(n16838), .ZN(
        n16842) );
  OAI21_X1 U19901 ( .B1(n19683), .B2(n16863), .A(n16842), .ZN(n16844) );
  AND2_X1 U19902 ( .A1(n16845), .A2(n16844), .ZN(n16843) );
  OAI221_X1 U19903 ( .B1(n16845), .B2(n16844), .C1(n20284), .C2(n16843), .A(
        n17156), .ZN(n16861) );
  NOR2_X1 U19904 ( .A1(P2_FLUSH_REG_SCAN_IN), .A2(P2_MORE_REG_SCAN_IN), .ZN(
        n16857) );
  MUX2_X1 U19905 ( .A(n16848), .B(n16847), .S(n16846), .Z(n16849) );
  AOI21_X1 U19906 ( .B1(n16851), .B2(n16850), .A(n16849), .ZN(n20301) );
  NOR3_X1 U19907 ( .A1(n10857), .A2(n16852), .A3(n10884), .ZN(n16853) );
  AOI21_X1 U19908 ( .B1(n16854), .B2(n20311), .A(n16853), .ZN(n16855) );
  OAI211_X1 U19909 ( .C1(n16857), .C2(n16856), .A(n20301), .B(n16855), .ZN(
        n16858) );
  AOI21_X1 U19910 ( .B1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n16859), .A(
        n16858), .ZN(n16860) );
  OAI211_X1 U19911 ( .C1(n16863), .C2(n16862), .A(n16861), .B(n16860), .ZN(
        n17237) );
  OAI21_X1 U19912 ( .B1(n17237), .B2(P2_STATE2_REG_1__SCAN_IN), .A(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n16867) );
  AOI211_X1 U19913 ( .C1(n16865), .C2(n16864), .A(n20307), .B(n20317), .ZN(
        n16866) );
  NAND2_X1 U19914 ( .A1(n16867), .A2(n16866), .ZN(n16869) );
  NAND2_X1 U19915 ( .A1(n16869), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n17245) );
  INV_X1 U19916 ( .A(n20191), .ZN(n20318) );
  NOR3_X1 U19917 ( .A1(n17245), .A2(P2_STATE2_REG_1__SCAN_IN), .A3(n20318), 
        .ZN(n16868) );
  AOI21_X1 U19918 ( .B1(n17236), .B2(n16869), .A(n16868), .ZN(n16871) );
  NOR2_X1 U19919 ( .A1(n16869), .A2(n20191), .ZN(n17238) );
  OAI21_X1 U19920 ( .B1(n17238), .B2(n17234), .A(P2_STATE2_REG_1__SCAN_IN), 
        .ZN(n16870) );
  OAI211_X1 U19921 ( .C1(n16871), .C2(n19741), .A(n19417), .B(n16870), .ZN(
        P2_U3177) );
  OAI22_X1 U19922 ( .A1(n18123), .A2(n16873), .B1(n18061), .B2(n16872), .ZN(
        n16875) );
  INV_X1 U19923 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n18188) );
  INV_X1 U19924 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n18184) );
  NAND2_X1 U19925 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n18077), .ZN(n18071) );
  AOI211_X1 U19926 ( .C1(n18188), .C2(n18071), .A(n18067), .B(n18102), .ZN(
        n16874) );
  AOI211_X1 U19927 ( .C1(BUF2_REG_4__SCAN_IN), .C2(n18076), .A(n16875), .B(
        n16874), .ZN(n16876) );
  INV_X1 U19928 ( .A(n16876), .ZN(P3_U2715) );
  NAND2_X1 U19929 ( .A1(n16877), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16879) );
  INV_X1 U19930 ( .A(n19232), .ZN(n19337) );
  NAND3_X1 U19931 ( .A1(n19322), .A2(n19349), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n19084) );
  NOR2_X2 U19932 ( .A1(n18856), .A2(n19084), .ZN(n16992) );
  OR2_X1 U19933 ( .A1(n16879), .A2(n18315), .ZN(n16896) );
  INV_X1 U19934 ( .A(n16990), .ZN(n18275) );
  NOR2_X1 U19935 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18275), .ZN(
        n17252) );
  NAND2_X1 U19936 ( .A1(n16992), .A2(n16879), .ZN(n17256) );
  OAI211_X1 U19937 ( .C1(n16910), .C2(n18313), .A(n18495), .B(n17256), .ZN(
        n17259) );
  NOR2_X1 U19938 ( .A1(n17252), .A2(n17259), .ZN(n16900) );
  INV_X1 U19939 ( .A(n16900), .ZN(n16888) );
  NOR2_X1 U19940 ( .A1(n19223), .A2(n21312), .ZN(n18368) );
  NAND2_X1 U19941 ( .A1(n18391), .A2(n17388), .ZN(n16885) );
  AOI21_X1 U19942 ( .B1(n9600), .B2(n16883), .A(n16882), .ZN(n16884) );
  OAI211_X1 U19943 ( .C1(n16886), .C2(n18380), .A(n16885), .B(n16884), .ZN(
        n16887) );
  AOI21_X1 U19944 ( .B1(n16888), .B2(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n16887), .ZN(n16889) );
  NOR2_X1 U19945 ( .A1(n16891), .A2(n16890), .ZN(n16892) );
  XOR2_X1 U19946 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n16892), .Z(
        n17037) );
  OR2_X1 U19947 ( .A1(n18407), .A2(n18381), .ZN(n16894) );
  INV_X1 U19948 ( .A(n18652), .ZN(n18360) );
  NAND2_X1 U19949 ( .A1(n18405), .A2(n18360), .ZN(n16893) );
  AND2_X2 U19950 ( .A1(n18438), .A2(n18568), .ZN(n18320) );
  NOR2_X1 U19951 ( .A1(n18350), .A2(n17027), .ZN(n16926) );
  NOR2_X1 U19952 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16895), .ZN(
        n17035) );
  NOR2_X1 U19953 ( .A1(n16896), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16902) );
  INV_X1 U19954 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n17401) );
  OAI22_X1 U19955 ( .A1(n18380), .A2(n17260), .B1(n17247), .B2(n18381), .ZN(
        n16897) );
  NOR2_X1 U19956 ( .A1(n18739), .A2(n19307), .ZN(n17034) );
  AOI21_X1 U19957 ( .B1(n16897), .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n17034), .ZN(n16899) );
  XNOR2_X1 U19958 ( .A(n17250), .B(n17401), .ZN(n17400) );
  NAND2_X1 U19959 ( .A1(n18391), .A2(n17400), .ZN(n16898) );
  OAI211_X1 U19960 ( .C1(n16900), .C2(n17401), .A(n16899), .B(n16898), .ZN(
        n16901) );
  AOI211_X1 U19961 ( .C1(n16926), .C2(n17035), .A(n16902), .B(n16901), .ZN(
        n16903) );
  OAI21_X1 U19962 ( .B1(n17037), .B2(n18451), .A(n16903), .ZN(P3_U2800) );
  NOR3_X1 U19963 ( .A1(n17027), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n17070), .ZN(n17057) );
  INV_X1 U19964 ( .A(n17057), .ZN(n16919) );
  INV_X1 U19965 ( .A(n17053), .ZN(n16904) );
  OAI21_X1 U19966 ( .B1(n9988), .B2(n17070), .A(n16904), .ZN(n16920) );
  OAI21_X1 U19967 ( .B1(n16920), .B2(n18357), .A(n16904), .ZN(n16906) );
  XNOR2_X1 U19968 ( .A(n18357), .B(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16905) );
  NAND2_X1 U19969 ( .A1(n16906), .A2(n16905), .ZN(n17051) );
  OAI211_X1 U19970 ( .C1(n16906), .C2(n16905), .A(n17051), .B(n18428), .ZN(
        n16918) );
  AOI21_X1 U19971 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18239), .A(
        n18313), .ZN(n16909) );
  AOI211_X1 U19972 ( .C1(n18368), .C2(n16907), .A(n18478), .B(n16909), .ZN(
        n18248) );
  OAI21_X1 U19973 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18275), .A(
        n18248), .ZN(n16924) );
  NOR2_X1 U19974 ( .A1(n17709), .A2(n16907), .ZN(n17384) );
  NAND2_X1 U19975 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17384), .ZN(
        n16921) );
  INV_X1 U19976 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16911) );
  AOI21_X1 U19977 ( .B1(n16921), .B2(n16911), .A(n16910), .ZN(n17424) );
  INV_X1 U19978 ( .A(n17424), .ZN(n16913) );
  NAND2_X1 U19979 ( .A1(n18693), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17060) );
  AOI22_X1 U19980 ( .A1(n18405), .A2(n17065), .B1(n9600), .B2(n17064), .ZN(
        n18241) );
  NAND2_X1 U19981 ( .A1(n18241), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16925) );
  NAND2_X1 U19982 ( .A1(n18380), .A2(n18381), .ZN(n18271) );
  NAND3_X1 U19983 ( .A1(n16925), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n18271), .ZN(n16912) );
  OAI211_X1 U19984 ( .C1(n18377), .C2(n16913), .A(n17060), .B(n16912), .ZN(
        n16916) );
  XNOR2_X1 U19985 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16914) );
  NOR3_X1 U19986 ( .A1(n18315), .A2(n16907), .A3(n16914), .ZN(n16915) );
  AOI211_X1 U19987 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n16924), .A(
        n16916), .B(n16915), .ZN(n16917) );
  OAI211_X1 U19988 ( .C1(n16919), .C2(n18350), .A(n16918), .B(n16917), .ZN(
        P3_U2802) );
  XNOR2_X1 U19989 ( .A(n16920), .B(n18365), .ZN(n17076) );
  INV_X1 U19990 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n19301) );
  OAI21_X1 U19991 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n17384), .A(
        n16921), .ZN(n17387) );
  OAI22_X1 U19992 ( .A1(n18739), .A2(n19301), .B1(n18377), .B2(n17387), .ZN(
        n16923) );
  NOR3_X1 U19993 ( .A1(n18315), .A2(n16907), .A3(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16922) );
  AOI211_X1 U19994 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n16924), .A(
        n16923), .B(n16922), .ZN(n16928) );
  OAI21_X1 U19995 ( .B1(n16926), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n16925), .ZN(n16927) );
  OAI211_X1 U19996 ( .C1(n17076), .C2(n18451), .A(n16928), .B(n16927), .ZN(
        P3_U2803) );
  INV_X1 U19997 ( .A(n16929), .ZN(n16930) );
  AOI21_X1 U19998 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n16930), .A(
        n18257), .ZN(n17093) );
  NOR2_X1 U19999 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n16931), .ZN(
        n17090) );
  INV_X1 U20000 ( .A(n16943), .ZN(n18249) );
  NOR2_X1 U20001 ( .A1(n16931), .A2(n18609), .ZN(n18255) );
  OAI22_X1 U20002 ( .A1(n18380), .A2(n18249), .B1(n18255), .B2(n18381), .ZN(
        n16954) );
  AOI22_X1 U20003 ( .A1(n18320), .A2(n17090), .B1(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n16954), .ZN(n16939) );
  NOR2_X1 U20004 ( .A1(n18315), .A2(n16932), .ZN(n18252) );
  INV_X1 U20005 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n16937) );
  AOI21_X1 U20006 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16949), .A(
        n18313), .ZN(n16933) );
  AOI211_X1 U20007 ( .C1(n16992), .C2(n16932), .A(n18478), .B(n16933), .ZN(
        n16951) );
  OAI21_X1 U20008 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18275), .A(
        n16951), .ZN(n18266) );
  NOR2_X1 U20009 ( .A1(n17709), .A2(n16932), .ZN(n16955) );
  INV_X1 U20010 ( .A(n16955), .ZN(n16934) );
  NOR3_X1 U20011 ( .A1(n17709), .A2(n16932), .A3(n16937), .ZN(n17383) );
  AOI21_X1 U20012 ( .B1(n16937), .B2(n16934), .A(n17383), .ZN(n17464) );
  AOI22_X1 U20013 ( .A1(n18693), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n18391), 
        .B2(n17464), .ZN(n16935) );
  INV_X1 U20014 ( .A(n16935), .ZN(n16936) );
  AOI221_X1 U20015 ( .B1(n18252), .B2(n16937), .C1(n18266), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n16936), .ZN(n16938) );
  OAI211_X1 U20016 ( .C1(n17093), .C2(n18451), .A(n16939), .B(n16938), .ZN(
        P3_U2806) );
  NAND2_X1 U20017 ( .A1(n18357), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16940) );
  OAI211_X1 U20018 ( .C1(n16941), .C2(n18269), .A(n18298), .B(n16940), .ZN(
        n16942) );
  XNOR2_X1 U20019 ( .A(n16942), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n18515) );
  INV_X1 U20020 ( .A(n18515), .ZN(n16960) );
  NAND3_X1 U20021 ( .A1(n18405), .A2(n18525), .A3(n16943), .ZN(n16948) );
  INV_X1 U20022 ( .A(n18609), .ZN(n16945) );
  INV_X1 U20023 ( .A(n18255), .ZN(n16944) );
  NAND3_X1 U20024 ( .A1(n9600), .A2(n16945), .A3(n16944), .ZN(n16947) );
  INV_X1 U20025 ( .A(n16946), .ZN(n18499) );
  AOI21_X1 U20026 ( .B1(n16948), .B2(n16947), .A(n18499), .ZN(n16953) );
  AOI21_X1 U20027 ( .B1(n16949), .B2(n16992), .A(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16950) );
  INV_X1 U20028 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n19293) );
  OAI22_X1 U20029 ( .A1(n16951), .A2(n16950), .B1(n18739), .B2(n19293), .ZN(
        n16952) );
  AOI211_X1 U20030 ( .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n16954), .A(
        n16953), .B(n16952), .ZN(n16959) );
  INV_X1 U20031 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16957) );
  AOI21_X1 U20032 ( .B1(n16957), .B2(n16956), .A(n16955), .ZN(n17474) );
  OAI21_X1 U20033 ( .B1(n18391), .B2(n16990), .A(n17474), .ZN(n16958) );
  OAI211_X1 U20034 ( .C1(n16960), .C2(n18451), .A(n16959), .B(n16958), .ZN(
        P3_U2807) );
  NAND2_X1 U20035 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16961), .ZN(
        n18369) );
  NOR2_X1 U20036 ( .A1(n16965), .A2(n18369), .ZN(n17562) );
  AOI21_X1 U20037 ( .B1(n18368), .B2(n16962), .A(n18478), .ZN(n18353) );
  OAI21_X1 U20038 ( .B1(n17562), .B2(n18313), .A(n18353), .ZN(n16976) );
  INV_X1 U20039 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16963) );
  INV_X1 U20040 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17560) );
  INV_X1 U20041 ( .A(n17562), .ZN(n17548) );
  NOR2_X1 U20042 ( .A1(n17560), .A2(n17548), .ZN(n17503) );
  INV_X1 U20043 ( .A(n17503), .ZN(n16974) );
  AND2_X1 U20044 ( .A1(n18338), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17527) );
  AOI21_X1 U20045 ( .B1(n16963), .B2(n16974), .A(n17527), .ZN(n17541) );
  AOI22_X1 U20046 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n16976), .B1(
        n18391), .B2(n17541), .ZN(n16968) );
  INV_X1 U20047 ( .A(n16961), .ZN(n16964) );
  NOR2_X1 U20048 ( .A1(n16964), .A2(n18315), .ZN(n18388) );
  INV_X1 U20049 ( .A(n18388), .ZN(n18375) );
  NOR2_X1 U20050 ( .A1(n16965), .A2(n18375), .ZN(n16977) );
  OAI211_X1 U20051 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n16977), .B(n16966), .ZN(n16967) );
  OAI211_X1 U20052 ( .C1(n19279), .C2(n18739), .A(n16968), .B(n16967), .ZN(
        n16969) );
  INV_X1 U20053 ( .A(n16969), .ZN(n16973) );
  AOI21_X1 U20054 ( .B1(n18365), .B2(n18343), .A(n16970), .ZN(n16971) );
  XOR2_X1 U20055 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n16971), .Z(
        n18595) );
  AND2_X1 U20056 ( .A1(n18405), .A2(n18343), .ZN(n16983) );
  AND2_X1 U20057 ( .A1(n9600), .A2(n18609), .ZN(n16985) );
  AOI22_X1 U20058 ( .A1(n18595), .A2(n18428), .B1(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18272), .ZN(n16972) );
  OAI211_X1 U20059 ( .C1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n18350), .A(
        n16973), .B(n16972), .ZN(P3_U2814) );
  OAI21_X1 U20060 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17562), .A(
        n16974), .ZN(n17550) );
  OAI22_X1 U20061 ( .A1(n18739), .A2(n19277), .B1(n18377), .B2(n17550), .ZN(
        n16975) );
  AOI221_X1 U20062 ( .B1(n16977), .B2(n17560), .C1(n16976), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n16975), .ZN(n16988) );
  NAND2_X1 U20063 ( .A1(n18361), .A2(n16978), .ZN(n18602) );
  AND2_X1 U20064 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16984) );
  NAND3_X1 U20065 ( .A1(n18360), .A2(n16984), .A3(n18664), .ZN(n16981) );
  OAI21_X1 U20066 ( .B1(n18619), .B2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n16979), .ZN(n16980) );
  AOI21_X1 U20067 ( .B1(n18358), .B2(n16981), .A(n16980), .ZN(n16982) );
  XOR2_X1 U20068 ( .A(n16982), .B(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .Z(
        n18607) );
  AOI22_X1 U20069 ( .A1(n16983), .A2(n18602), .B1(n18428), .B2(n18607), .ZN(
        n16987) );
  NAND2_X1 U20070 ( .A1(n16984), .A2(n9659), .ZN(n18351) );
  NAND2_X1 U20071 ( .A1(n16978), .A2(n18351), .ZN(n18608) );
  NAND2_X1 U20072 ( .A1(n18608), .A2(n16985), .ZN(n16986) );
  NAND3_X1 U20073 ( .A1(n16988), .A2(n16987), .A3(n16986), .ZN(P3_U2815) );
  INV_X1 U20074 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17637) );
  INV_X1 U20075 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17656) );
  NOR3_X1 U20076 ( .A1(n17709), .A2(n17632), .A3(n17656), .ZN(n17003) );
  INV_X1 U20077 ( .A(n17003), .ZN(n16989) );
  NAND2_X1 U20078 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18456), .ZN(
        n17674) );
  INV_X1 U20079 ( .A(n17674), .ZN(n17661) );
  NAND2_X1 U20080 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17661), .ZN(
        n17660) );
  NOR2_X1 U20081 ( .A1(n16991), .A2(n17660), .ZN(n17619) );
  AOI21_X1 U20082 ( .B1(n17637), .B2(n16989), .A(n17619), .ZN(n17634) );
  INV_X1 U20083 ( .A(n17632), .ZN(n16994) );
  NAND2_X1 U20084 ( .A1(n16994), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16993) );
  INV_X1 U20085 ( .A(n16991), .ZN(n18401) );
  AOI211_X1 U20086 ( .C1(n17637), .C2(n16993), .A(n18401), .B(n18857), .ZN(
        n16996) );
  INV_X1 U20087 ( .A(n18368), .ZN(n17098) );
  OAI21_X1 U20088 ( .B1(n17098), .B2(n16994), .A(n18495), .ZN(n17006) );
  INV_X1 U20089 ( .A(n17006), .ZN(n18372) );
  OAI22_X1 U20090 ( .A1(n18372), .A2(n17637), .B1(n18739), .B2(n19264), .ZN(
        n16995) );
  AOI211_X1 U20091 ( .C1(n17634), .C2(n18426), .A(n16996), .B(n16995), .ZN(
        n17001) );
  INV_X1 U20092 ( .A(n16997), .ZN(n16998) );
  AOI22_X1 U20093 ( .A1(n18428), .A2(n16999), .B1(n18405), .B2(n16998), .ZN(
        n17000) );
  OAI211_X1 U20094 ( .C1(n18381), .C2(n17002), .A(n17001), .B(n17000), .ZN(
        P3_U2822) );
  AOI21_X1 U20095 ( .B1(n17656), .B2(n17660), .A(n17003), .ZN(n17648) );
  NAND2_X1 U20096 ( .A1(n17004), .A2(n9600), .ZN(n17008) );
  NOR2_X1 U20097 ( .A1(n17632), .A2(n18857), .ZN(n18400) );
  AOI221_X1 U20098 ( .B1(n18400), .B2(n17656), .C1(n17006), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n17005), .ZN(n17007) );
  OAI211_X1 U20099 ( .C1(n17009), .C2(n18488), .A(n17008), .B(n17007), .ZN(
        n17010) );
  AOI21_X1 U20100 ( .B1(n18426), .B2(n17648), .A(n17010), .ZN(n17011) );
  INV_X1 U20101 ( .A(n17011), .ZN(P3_U2823) );
  OAI21_X1 U20102 ( .B1(n14272), .B2(n17098), .A(n18495), .ZN(n18480) );
  INV_X1 U20103 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17015) );
  NOR2_X1 U20104 ( .A1(n17709), .A2(n17012), .ZN(n17675) );
  AOI21_X1 U20105 ( .B1(n17015), .B2(n17013), .A(n17675), .ZN(n17694) );
  AOI22_X1 U20106 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18480), .B1(
        n17694), .B2(n18426), .ZN(n17020) );
  AOI22_X1 U20107 ( .A1(n18473), .A2(n17014), .B1(n18693), .B2(
        P3_REIP_REG_4__SCAN_IN), .ZN(n17019) );
  NAND2_X1 U20108 ( .A1(n14272), .A2(n17015), .ZN(n17690) );
  OAI22_X1 U20109 ( .A1(n18381), .A2(n17016), .B1(n18857), .B2(n17690), .ZN(
        n17017) );
  INV_X1 U20110 ( .A(n17017), .ZN(n17018) );
  NAND3_X1 U20111 ( .A1(n17020), .A2(n17019), .A3(n17018), .ZN(P3_U2826) );
  OAI22_X1 U20112 ( .A1(n17709), .A2(n18455), .B1(n18490), .B2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17021) );
  INV_X1 U20113 ( .A(n17021), .ZN(n17024) );
  AOI22_X1 U20114 ( .A1(n9600), .A2(n17022), .B1(n18693), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17023) );
  OAI211_X1 U20115 ( .C1(n18488), .C2(n17025), .A(n17024), .B(n17023), .ZN(
        P3_U2829) );
  INV_X1 U20116 ( .A(n17026), .ZN(n18500) );
  NOR3_X1 U20117 ( .A1(n18500), .A2(n17027), .A3(n18616), .ZN(n17028) );
  AOI21_X1 U20118 ( .B1(n17044), .B2(n18728), .A(n17028), .ZN(n17029) );
  OAI21_X1 U20119 ( .B1(n18622), .B2(n17065), .A(n17029), .ZN(n17111) );
  OAI22_X1 U20120 ( .A1(n17247), .A2(n18629), .B1(n17260), .B2(n18622), .ZN(
        n17030) );
  NOR2_X1 U20121 ( .A1(n18701), .A2(n17030), .ZN(n17107) );
  AOI21_X1 U20122 ( .B1(n17107), .B2(n17032), .A(n17031), .ZN(n17033) );
  AOI211_X1 U20123 ( .C1(n17035), .C2(n17111), .A(n17034), .B(n17033), .ZN(
        n17036) );
  OAI21_X1 U20124 ( .B1(n17037), .B2(n18689), .A(n17036), .ZN(P3_U2832) );
  INV_X1 U20125 ( .A(n17112), .ZN(n17038) );
  NOR2_X1 U20126 ( .A1(n17065), .A2(n17038), .ZN(n17262) );
  INV_X1 U20127 ( .A(n19183), .ZN(n17043) );
  NAND3_X1 U20128 ( .A1(n17040), .A2(n17039), .A3(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17041) );
  NAND4_X1 U20129 ( .A1(n17051), .A2(n17043), .A3(n17042), .A4(n17041), .ZN(
        n17048) );
  NAND2_X1 U20130 ( .A1(n17044), .A2(n17112), .ZN(n17249) );
  NAND2_X1 U20131 ( .A1(n18712), .A2(n18730), .ZN(n18669) );
  AOI21_X1 U20132 ( .B1(n17070), .B2(n18669), .A(n17045), .ZN(n17109) );
  INV_X1 U20133 ( .A(n17109), .ZN(n17046) );
  AOI211_X1 U20134 ( .C1(n19178), .C2(n17249), .A(n18616), .B(n17046), .ZN(
        n17047) );
  OAI211_X1 U20135 ( .C1(n17262), .C2(n18524), .A(n17048), .B(n17047), .ZN(
        n17049) );
  NAND3_X1 U20136 ( .A1(n17049), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n18739), .ZN(n17062) );
  NOR2_X1 U20137 ( .A1(n17050), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n17052) );
  OAI211_X1 U20138 ( .C1(n17053), .C2(n17052), .A(n17051), .B(n18672), .ZN(
        n17061) );
  INV_X1 U20139 ( .A(n19178), .ZN(n18655) );
  OR2_X1 U20140 ( .A1(n18407), .A2(n18655), .ZN(n17055) );
  NAND2_X1 U20141 ( .A1(n18653), .A2(n18360), .ZN(n17054) );
  NAND2_X1 U20142 ( .A1(n17055), .A2(n17054), .ZN(n18567) );
  NAND2_X1 U20143 ( .A1(n18567), .A2(n18568), .ZN(n17056) );
  INV_X1 U20144 ( .A(n18532), .ZN(n17058) );
  NAND3_X1 U20145 ( .A1(n17058), .A2(n18724), .A3(n17057), .ZN(n17059) );
  NAND4_X1 U20146 ( .A1(n17062), .A2(n17061), .A3(n17060), .A4(n17059), .ZN(
        P3_U2834) );
  NOR2_X1 U20147 ( .A1(n18532), .A2(n18499), .ZN(n18514) );
  AOI22_X1 U20148 ( .A1(n18658), .A2(n17063), .B1(n18680), .B2(n18509), .ZN(
        n17069) );
  AOI22_X1 U20149 ( .A1(n17065), .A2(n18653), .B1(n19178), .B2(n17064), .ZN(
        n17068) );
  OR2_X1 U20150 ( .A1(n18715), .A2(n17066), .ZN(n17085) );
  OAI21_X1 U20151 ( .B1(n18501), .B2(n17085), .A(n18576), .ZN(n18502) );
  NAND4_X1 U20152 ( .A1(n17069), .A2(n17068), .A3(n17067), .A4(n18502), .ZN(
        n17080) );
  AOI211_X1 U20153 ( .C1(n18680), .C2(n12028), .A(n17070), .B(n17080), .ZN(
        n17071) );
  OAI22_X1 U20154 ( .A1(n17071), .A2(n18616), .B1(n17070), .B2(n18729), .ZN(
        n17072) );
  OAI221_X1 U20155 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17073), 
        .C1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n18514), .A(n17072), .ZN(
        n17075) );
  NAND2_X1 U20156 ( .A1(n18693), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17074) );
  OAI211_X1 U20157 ( .C1(n17076), .C2(n18689), .A(n17075), .B(n17074), .ZN(
        P3_U2835) );
  INV_X1 U20158 ( .A(n17077), .ZN(n17078) );
  AOI21_X1 U20159 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17079), .A(
        n17078), .ZN(n18242) );
  AND2_X1 U20160 ( .A1(n17080), .A2(n18739), .ZN(n17081) );
  OAI21_X1 U20161 ( .B1(n17081), .B2(n18701), .A(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17083) );
  NOR4_X1 U20162 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18501), .A3(
        n18499), .A4(n18509), .ZN(n18244) );
  AOI22_X1 U20163 ( .A1(n18244), .A2(n18560), .B1(n18693), .B2(
        P3_REIP_REG_26__SCAN_IN), .ZN(n17082) );
  OAI211_X1 U20164 ( .C1(n18242), .C2(n18689), .A(n17083), .B(n17082), .ZN(
        P3_U2836) );
  OAI22_X1 U20165 ( .A1(n18249), .A2(n18524), .B1(n18255), .B2(n18655), .ZN(
        n17084) );
  AOI211_X1 U20166 ( .C1(n18576), .C2(n17085), .A(n18701), .B(n17084), .ZN(
        n17087) );
  OAI21_X1 U20167 ( .B1(n18499), .B2(n18571), .A(n19179), .ZN(n18503) );
  NAND3_X1 U20168 ( .A1(n18503), .A2(n17087), .A3(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17086) );
  NAND2_X1 U20169 ( .A1(n17086), .A2(n18739), .ZN(n18517) );
  AOI211_X1 U20170 ( .C1(n17088), .C2(n17087), .A(n12022), .B(n18517), .ZN(
        n17089) );
  AOI21_X1 U20171 ( .B1(n17090), .B2(n18560), .A(n17089), .ZN(n17092) );
  NAND2_X1 U20172 ( .A1(n18693), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n17091) );
  OAI211_X1 U20173 ( .C1(n17093), .C2(n18689), .A(n17092), .B(n17091), .ZN(
        P3_U2838) );
  INV_X1 U20174 ( .A(n19084), .ZN(n18748) );
  NOR2_X1 U20175 ( .A1(n19322), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18791) );
  INV_X1 U20176 ( .A(n18791), .ZN(n17097) );
  NOR2_X1 U20177 ( .A1(n17094), .A2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n18740) );
  INV_X1 U20178 ( .A(n18740), .ZN(n17095) );
  NOR3_X1 U20179 ( .A1(n17095), .A2(n17972), .A3(P3_FLUSH_REG_SCAN_IN), .ZN(
        n17096) );
  OAI21_X1 U20180 ( .B1(n17096), .B2(n19320), .A(n18856), .ZN(n18752) );
  NAND2_X1 U20181 ( .A1(n17097), .A2(n18752), .ZN(n18744) );
  NOR2_X1 U20182 ( .A1(n18748), .A2(n18744), .ZN(n17099) );
  AOI21_X1 U20183 ( .B1(n18741), .B2(n17098), .A(P3_STATE2_REG_3__SCAN_IN), 
        .ZN(n18746) );
  INV_X1 U20184 ( .A(n18746), .ZN(n18745) );
  NAND2_X1 U20185 ( .A1(n12171), .A2(n18745), .ZN(n18925) );
  OAI22_X1 U20186 ( .A1(n12171), .A2(n17099), .B1(n18925), .B2(n18744), .ZN(
        P3_U2864) );
  INV_X1 U20187 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17102) );
  NOR2_X1 U20188 ( .A1(n18740), .A2(n17100), .ZN(n19187) );
  NAND3_X1 U20189 ( .A1(n17103), .A2(n19350), .A3(n19187), .ZN(n17101) );
  OAI21_X1 U20190 ( .B1(n17103), .B2(n17102), .A(n17101), .ZN(P3_U3284) );
  XNOR2_X1 U20191 ( .A(n17105), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17265) );
  NAND2_X1 U20192 ( .A1(n17106), .A2(n18593), .ZN(n17108) );
  OAI221_X1 U20193 ( .B1(n18616), .B2(n17109), .C1(n18616), .C2(n17108), .A(
        n17107), .ZN(n17110) );
  AOI22_X1 U20194 ( .A1(n18693), .A2(P3_REIP_REG_29__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n17110), .ZN(n17114) );
  NAND3_X1 U20195 ( .A1(n17112), .A2(n17248), .A3(n17111), .ZN(n17113) );
  OAI211_X1 U20196 ( .C1(n17265), .C2(n18689), .A(n17114), .B(n17113), .ZN(
        P3_U2833) );
  NOR2_X1 U20197 ( .A1(n17115), .A2(n17143), .ZN(n17150) );
  INV_X1 U20198 ( .A(n17120), .ZN(n17124) );
  AOI211_X1 U20199 ( .C1(n17118), .C2(n17119), .A(n17117), .B(n17116), .ZN(
        n17122) );
  OAI21_X1 U20200 ( .B1(n17119), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n20958), .ZN(n17121) );
  OAI22_X1 U20201 ( .A1(n17122), .A2(n17121), .B1(n17120), .B2(n20840), .ZN(
        n17123) );
  OAI21_X1 U20202 ( .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n17124), .A(
        n17123), .ZN(n17125) );
  AOI222_X1 U20203 ( .A1(n20589), .A2(n17126), .B1(n20589), .B2(n17125), .C1(
        n17126), .C2(n17125), .ZN(n17134) );
  AND3_X1 U20204 ( .A1(n17129), .A2(n17128), .A3(n17127), .ZN(n17133) );
  AOI221_X1 U20205 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(n17131), .C1(
        P1_MORE_REG_SCAN_IN), .C2(n17131), .A(n17130), .ZN(n17132) );
  OAI211_X1 U20206 ( .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n17134), .A(
        n17133), .B(n17132), .ZN(n17145) );
  NOR3_X1 U20207 ( .A1(n13298), .A2(n17135), .A3(n17153), .ZN(n17138) );
  NAND3_X1 U20208 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21142), .A3(n10368), 
        .ZN(n17136) );
  AOI22_X1 U20209 ( .A1(n17138), .A2(n17137), .B1(n21134), .B2(n17136), .ZN(
        n17184) );
  INV_X1 U20210 ( .A(n17184), .ZN(n17139) );
  AOI221_X1 U20211 ( .B1(n13636), .B2(n10368), .C1(n13636), .C2(n17145), .A(
        n17139), .ZN(n17140) );
  INV_X1 U20212 ( .A(n17140), .ZN(n17190) );
  NAND2_X1 U20213 ( .A1(n17190), .A2(n10368), .ZN(n17149) );
  OAI211_X1 U20214 ( .C1(n12693), .C2(P1_FLUSH_REG_SCAN_IN), .A(n17142), .B(
        n17141), .ZN(n21387) );
  OAI211_X1 U20215 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n21221), .A(n21387), 
        .B(n17143), .ZN(n17144) );
  AOI21_X1 U20216 ( .B1(n17146), .B2(n17145), .A(n17144), .ZN(n17147) );
  AND2_X1 U20217 ( .A1(n17190), .A2(n17147), .ZN(n17148) );
  OAI22_X1 U20218 ( .A1(n17150), .A2(n17149), .B1(n17148), .B2(n10368), .ZN(
        P1_U3161) );
  INV_X1 U20219 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n21150) );
  INV_X1 U20220 ( .A(HOLD), .ZN(n20199) );
  INV_X1 U20221 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n21151) );
  NAND2_X1 U20222 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n17151) );
  OAI21_X1 U20223 ( .B1(n20199), .B2(n21150), .A(n17151), .ZN(n17152) );
  OAI21_X1 U20224 ( .B1(n20199), .B2(n21151), .A(n17152), .ZN(n17154) );
  OAI211_X1 U20225 ( .C1(n21221), .C2(n21150), .A(n17154), .B(n17153), .ZN(
        P1_U3195) );
  INV_X1 U20226 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n21268) );
  NOR2_X1 U20227 ( .A1(n21268), .A2(n17155), .ZN(P1_U2905) );
  NOR2_X1 U20228 ( .A1(n17156), .A2(n20291), .ZN(P2_U3047) );
  OAI222_X1 U20229 ( .A1(n9869), .A2(n20387), .B1(n17157), .B2(n20338), .C1(
        n20583), .C2(n20382), .ZN(n17158) );
  INV_X1 U20230 ( .A(n17158), .ZN(n17160) );
  OAI211_X1 U20231 ( .C1(n12605), .C2(n17161), .A(n17160), .B(n17159), .ZN(
        P1_U2992) );
  AOI22_X1 U20232 ( .A1(n20511), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n20577), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n17167) );
  OR2_X1 U20233 ( .A1(n17163), .A2(n17162), .ZN(n17164) );
  AND2_X1 U20234 ( .A1(n17165), .A2(n17164), .ZN(n17177) );
  AOI22_X1 U20235 ( .A1(n20412), .A2(n20518), .B1(n20519), .B2(n17177), .ZN(
        n17166) );
  OAI211_X1 U20236 ( .C1(n9869), .C2(n20415), .A(n17167), .B(n17166), .ZN(
        P1_U2994) );
  INV_X1 U20237 ( .A(n17168), .ZN(n20389) );
  AOI21_X1 U20238 ( .B1(n20560), .B2(n20389), .A(n17169), .ZN(n17170) );
  OAI21_X1 U20239 ( .B1(n17171), .B2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n17170), .ZN(n17172) );
  AOI21_X1 U20240 ( .B1(n17173), .B2(n20563), .A(n17172), .ZN(n17174) );
  OAI21_X1 U20241 ( .B1(n17175), .B2(n13178), .A(n17174), .ZN(P1_U3025) );
  INV_X1 U20242 ( .A(n17176), .ZN(n20403) );
  AOI22_X1 U20243 ( .A1(n20560), .A2(n20403), .B1(n20526), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n17180) );
  AOI22_X1 U20244 ( .A1(n17178), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B1(
        n20563), .B2(n17177), .ZN(n17179) );
  OAI211_X1 U20245 ( .C1(n20539), .C2(n17181), .A(n17180), .B(n17179), .ZN(
        P1_U3026) );
  NAND2_X1 U20246 ( .A1(n20963), .A2(n21221), .ZN(n17188) );
  NAND4_X1 U20247 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_0__SCAN_IN), .A3(n21070), .A4(n21221), .ZN(n17182) );
  AND2_X1 U20248 ( .A1(n17183), .A2(n17182), .ZN(n21135) );
  AOI21_X1 U20249 ( .B1(n21135), .B2(n17185), .A(n17184), .ZN(n17187) );
  AOI21_X1 U20250 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n17190), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n17186) );
  AOI211_X1 U20251 ( .C1(n21218), .C2(n17188), .A(n17187), .B(n17186), .ZN(
        P1_U3162) );
  OAI221_X1 U20252 ( .B1(n20963), .B2(P1_STATE2_REG_0__SCAN_IN), .C1(n20963), 
        .C2(n17190), .A(n17189), .ZN(P1_U3466) );
  AOI22_X1 U20253 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19571), .B1(n17192), 
        .B2(n17191), .ZN(n17197) );
  AOI222_X1 U20254 ( .A1(n17195), .A2(n19577), .B1(n19592), .B2(n17194), .C1(
        n17193), .C2(n9627), .ZN(n17196) );
  OAI211_X1 U20255 ( .C1(n17199), .C2(n17198), .A(n17197), .B(n17196), .ZN(
        P2_U3009) );
  OAI22_X1 U20256 ( .A1(n17203), .A2(n17202), .B1(n17201), .B2(n17200), .ZN(
        n17204) );
  AOI21_X1 U20257 ( .B1(n17205), .B2(n17224), .A(n17204), .ZN(n17206) );
  OAI21_X1 U20258 ( .B1(n17207), .B2(n17227), .A(n17206), .ZN(n17208) );
  AOI21_X1 U20259 ( .B1(n17210), .B2(n17209), .A(n17208), .ZN(n17211) );
  OAI221_X1 U20260 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n17214), .C1(
        n17213), .C2(n17212), .A(n17211), .ZN(P2_U3043) );
  AOI22_X1 U20261 ( .A1(n17216), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n17215), .B2(n19481), .ZN(n17231) );
  AND2_X1 U20262 ( .A1(n17218), .A2(n17217), .ZN(n17220) );
  OR2_X1 U20263 ( .A1(n17220), .A2(n17219), .ZN(n19589) );
  NOR2_X1 U20264 ( .A1(n17221), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17222) );
  NOR2_X1 U20265 ( .A1(n17223), .A2(n17222), .ZN(n19585) );
  NAND2_X1 U20266 ( .A1(n17224), .A2(n19585), .ZN(n17225) );
  OAI21_X1 U20267 ( .B1(n19589), .B2(n17226), .A(n17225), .ZN(n17229) );
  INV_X1 U20268 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n19375) );
  NAND2_X1 U20269 ( .A1(n19571), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n19587) );
  OAI21_X1 U20270 ( .B1(n17227), .B2(n11577), .A(n19587), .ZN(n17228) );
  NOR2_X1 U20271 ( .A1(n17229), .A2(n17228), .ZN(n17230) );
  OAI211_X1 U20272 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n17232), .A(
        n17231), .B(n17230), .ZN(P2_U3046) );
  INV_X1 U20273 ( .A(n17233), .ZN(n17235) );
  AOI211_X1 U20274 ( .C1(n17237), .C2(n17236), .A(n17235), .B(n17234), .ZN(
        n17242) );
  AOI21_X1 U20275 ( .B1(n17239), .B2(n20319), .A(n17238), .ZN(n17240) );
  OAI21_X1 U20276 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n17240), .A(n17245), 
        .ZN(n17241) );
  OAI211_X1 U20277 ( .C1(n20297), .C2(n17243), .A(n17242), .B(n17241), .ZN(
        P2_U3176) );
  AOI21_X1 U20278 ( .B1(n17245), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n17244), 
        .ZN(n17246) );
  INV_X1 U20279 ( .A(n17246), .ZN(P2_U3593) );
  AOI211_X1 U20280 ( .C1(n17249), .C2(n17248), .A(n17247), .B(n18381), .ZN(
        n17258) );
  NAND2_X1 U20281 ( .A1(n18693), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n17254) );
  AOI21_X1 U20282 ( .B1(n17251), .B2(n17412), .A(n17250), .ZN(n17410) );
  OAI21_X1 U20283 ( .B1(n17252), .B2(n18391), .A(n17410), .ZN(n17253) );
  OAI211_X1 U20284 ( .C1(n17256), .C2(n17255), .A(n17254), .B(n17253), .ZN(
        n17257) );
  AOI211_X1 U20285 ( .C1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n17259), .A(
        n17258), .B(n17257), .ZN(n17264) );
  INV_X1 U20286 ( .A(n17260), .ZN(n17261) );
  OAI211_X1 U20287 ( .C1(n17262), .C2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n18405), .B(n17261), .ZN(n17263) );
  OAI211_X1 U20288 ( .C1(n17265), .C2(n18451), .A(n17264), .B(n17263), .ZN(
        P3_U2801) );
  NOR3_X1 U20289 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n17267) );
  NOR4_X1 U20290 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n17266) );
  NAND4_X1 U20291 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n17267), .A3(n17266), .A4(
        U215), .ZN(U213) );
  INV_X1 U20292 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19486) );
  INV_X2 U20293 ( .A(U214), .ZN(n17314) );
  NOR2_X2 U20294 ( .A1(n17314), .A2(n17268), .ZN(n17317) );
  OAI222_X1 U20295 ( .A1(U212), .A2(n19486), .B1(n17316), .B2(n19643), .C1(
        U214), .C2(n21268), .ZN(U216) );
  AOI222_X1 U20296 ( .A1(n17313), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n17317), 
        .B2(BUF1_REG_30__SCAN_IN), .C1(n17314), .C2(P1_DATAO_REG_30__SCAN_IN), 
        .ZN(n17269) );
  INV_X1 U20297 ( .A(n17269), .ZN(U217) );
  AOI222_X1 U20298 ( .A1(n17313), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(n17317), 
        .B2(BUF1_REG_29__SCAN_IN), .C1(n17314), .C2(P1_DATAO_REG_29__SCAN_IN), 
        .ZN(n17270) );
  INV_X1 U20299 ( .A(n17270), .ZN(U218) );
  INV_X1 U20300 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n17272) );
  AOI22_X1 U20301 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n17314), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n17313), .ZN(n17271) );
  OAI21_X1 U20302 ( .B1(n17272), .B2(n17316), .A(n17271), .ZN(U219) );
  INV_X1 U20303 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n17274) );
  AOI22_X1 U20304 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n17314), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n17313), .ZN(n17273) );
  OAI21_X1 U20305 ( .B1(n17274), .B2(n17316), .A(n17273), .ZN(U220) );
  INV_X1 U20306 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n17276) );
  AOI22_X1 U20307 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n17314), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n17313), .ZN(n17275) );
  OAI21_X1 U20308 ( .B1(n17276), .B2(n17316), .A(n17275), .ZN(U221) );
  INV_X1 U20309 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n17278) );
  AOI22_X1 U20310 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n17314), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n17313), .ZN(n17277) );
  OAI21_X1 U20311 ( .B1(n17278), .B2(n17316), .A(n17277), .ZN(U222) );
  INV_X1 U20312 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n17280) );
  AOI22_X1 U20313 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n17314), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n17313), .ZN(n17279) );
  OAI21_X1 U20314 ( .B1(n17280), .B2(n17316), .A(n17279), .ZN(U223) );
  INV_X1 U20315 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n17282) );
  AOI22_X1 U20316 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n17314), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n17313), .ZN(n17281) );
  OAI21_X1 U20317 ( .B1(n17282), .B2(n17316), .A(n17281), .ZN(U224) );
  AOI22_X1 U20318 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n17314), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n17313), .ZN(n17283) );
  OAI21_X1 U20319 ( .B1(n19632), .B2(n17316), .A(n17283), .ZN(U225) );
  INV_X1 U20320 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n17285) );
  AOI22_X1 U20321 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n17314), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n17313), .ZN(n17284) );
  OAI21_X1 U20322 ( .B1(n17285), .B2(n17316), .A(n17284), .ZN(U226) );
  AOI22_X1 U20323 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n17314), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n17313), .ZN(n17286) );
  OAI21_X1 U20324 ( .B1(n17287), .B2(n17316), .A(n17286), .ZN(U227) );
  INV_X1 U20325 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n17289) );
  AOI22_X1 U20326 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n17314), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n17313), .ZN(n17288) );
  OAI21_X1 U20327 ( .B1(n17289), .B2(n17316), .A(n17288), .ZN(U228) );
  INV_X1 U20328 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n17291) );
  AOI22_X1 U20329 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n17314), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n17313), .ZN(n17290) );
  OAI21_X1 U20330 ( .B1(n17291), .B2(n17316), .A(n17290), .ZN(U229) );
  AOI222_X1 U20331 ( .A1(n17313), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n17317), 
        .B2(BUF1_REG_17__SCAN_IN), .C1(n17314), .C2(P1_DATAO_REG_17__SCAN_IN), 
        .ZN(n17292) );
  INV_X1 U20332 ( .A(n17292), .ZN(U230) );
  AOI22_X1 U20333 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n17314), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n17313), .ZN(n17293) );
  OAI21_X1 U20334 ( .B1(n17294), .B2(n17316), .A(n17293), .ZN(U231) );
  AOI22_X1 U20335 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n17314), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n17313), .ZN(n17295) );
  OAI21_X1 U20336 ( .B1(n14377), .B2(n17316), .A(n17295), .ZN(U232) );
  AOI22_X1 U20337 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n17314), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n17313), .ZN(n17296) );
  OAI21_X1 U20338 ( .B1(n15014), .B2(n17316), .A(n17296), .ZN(U233) );
  AOI22_X1 U20339 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n17314), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n17313), .ZN(n17297) );
  OAI21_X1 U20340 ( .B1(n17298), .B2(n17316), .A(n17297), .ZN(U234) );
  INV_X1 U20341 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n21295) );
  AOI22_X1 U20342 ( .A1(BUF1_REG_12__SCAN_IN), .A2(n17317), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n17313), .ZN(n17299) );
  OAI21_X1 U20343 ( .B1(n21295), .B2(U214), .A(n17299), .ZN(U235) );
  AOI222_X1 U20344 ( .A1(n17313), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n17317), 
        .B2(BUF1_REG_11__SCAN_IN), .C1(n17314), .C2(P1_DATAO_REG_11__SCAN_IN), 
        .ZN(n17300) );
  INV_X1 U20345 ( .A(n17300), .ZN(U236) );
  INV_X1 U20346 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n17302) );
  AOI22_X1 U20347 ( .A1(BUF1_REG_10__SCAN_IN), .A2(n17317), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n17314), .ZN(n17301) );
  OAI21_X1 U20348 ( .B1(n17302), .B2(U212), .A(n17301), .ZN(U237) );
  AOI22_X1 U20349 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n17314), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n17313), .ZN(n17303) );
  OAI21_X1 U20350 ( .B1(n17304), .B2(n17316), .A(n17303), .ZN(U238) );
  INV_X1 U20351 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n17306) );
  AOI22_X1 U20352 ( .A1(BUF1_REG_8__SCAN_IN), .A2(n17317), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n17314), .ZN(n17305) );
  OAI21_X1 U20353 ( .B1(n17306), .B2(U212), .A(n17305), .ZN(U239) );
  AOI22_X1 U20354 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n17314), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n17313), .ZN(n17307) );
  OAI21_X1 U20355 ( .B1(n13906), .B2(n17316), .A(n17307), .ZN(U240) );
  INV_X1 U20356 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n17325) );
  AOI22_X1 U20357 ( .A1(BUF1_REG_6__SCAN_IN), .A2(n17317), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n17314), .ZN(n17308) );
  OAI21_X1 U20358 ( .B1(n17325), .B2(U212), .A(n17308), .ZN(U241) );
  INV_X1 U20359 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n17324) );
  AOI22_X1 U20360 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n17317), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n17314), .ZN(n17309) );
  OAI21_X1 U20361 ( .B1(n17324), .B2(U212), .A(n17309), .ZN(U242) );
  INV_X1 U20362 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n17323) );
  AOI22_X1 U20363 ( .A1(BUF1_REG_4__SCAN_IN), .A2(n17317), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n17314), .ZN(n17310) );
  OAI21_X1 U20364 ( .B1(n17323), .B2(U212), .A(n17310), .ZN(U243) );
  INV_X1 U20365 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n17322) );
  AOI22_X1 U20366 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n17317), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n17314), .ZN(n17311) );
  OAI21_X1 U20367 ( .B1(n17322), .B2(U212), .A(n17311), .ZN(U244) );
  INV_X1 U20368 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n17321) );
  AOI22_X1 U20369 ( .A1(BUF1_REG_2__SCAN_IN), .A2(n17317), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n17314), .ZN(n17312) );
  OAI21_X1 U20370 ( .B1(n17321), .B2(U212), .A(n17312), .ZN(U245) );
  AOI22_X1 U20371 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n17314), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n17313), .ZN(n17315) );
  OAI21_X1 U20372 ( .B1(n16182), .B2(n17316), .A(n17315), .ZN(U246) );
  INV_X1 U20373 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n17319) );
  AOI22_X1 U20374 ( .A1(BUF1_REG_0__SCAN_IN), .A2(n17317), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n17314), .ZN(n17318) );
  OAI21_X1 U20375 ( .B1(n17319), .B2(U212), .A(n17318), .ZN(U247) );
  INV_X1 U20376 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18756) );
  AOI22_X1 U20377 ( .A1(n17348), .A2(n17319), .B1(n18756), .B2(U215), .ZN(U251) );
  OAI22_X1 U20378 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n17348), .ZN(n17320) );
  INV_X1 U20379 ( .A(n17320), .ZN(U252) );
  AOI22_X1 U20380 ( .A1(n17348), .A2(n17321), .B1(n18763), .B2(U215), .ZN(U253) );
  INV_X1 U20381 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18767) );
  AOI22_X1 U20382 ( .A1(n17348), .A2(n17322), .B1(n18767), .B2(U215), .ZN(U254) );
  INV_X1 U20383 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18772) );
  AOI22_X1 U20384 ( .A1(n17348), .A2(n17323), .B1(n18772), .B2(U215), .ZN(U255) );
  INV_X1 U20385 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18776) );
  AOI22_X1 U20386 ( .A1(n17348), .A2(n17324), .B1(n18776), .B2(U215), .ZN(U256) );
  INV_X1 U20387 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18780) );
  AOI22_X1 U20388 ( .A1(n17348), .A2(n17325), .B1(n18780), .B2(U215), .ZN(U257) );
  OAI22_X1 U20389 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n17348), .ZN(n17326) );
  INV_X1 U20390 ( .A(n17326), .ZN(U258) );
  OAI22_X1 U20391 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n17348), .ZN(n17327) );
  INV_X1 U20392 ( .A(n17327), .ZN(U259) );
  OAI22_X1 U20393 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n17348), .ZN(n17328) );
  INV_X1 U20394 ( .A(n17328), .ZN(U260) );
  OAI22_X1 U20395 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n17348), .ZN(n17329) );
  INV_X1 U20396 ( .A(n17329), .ZN(U261) );
  INV_X1 U20397 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n18225) );
  AOI22_X1 U20398 ( .A1(n17349), .A2(n17330), .B1(n18225), .B2(U215), .ZN(U262) );
  OAI22_X1 U20399 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n17348), .ZN(n17331) );
  INV_X1 U20400 ( .A(n17331), .ZN(U263) );
  OAI22_X1 U20401 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n17348), .ZN(n17332) );
  INV_X1 U20402 ( .A(n17332), .ZN(U264) );
  OAI22_X1 U20403 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n17348), .ZN(n17333) );
  INV_X1 U20404 ( .A(n17333), .ZN(U265) );
  OAI22_X1 U20405 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n17348), .ZN(n17334) );
  INV_X1 U20406 ( .A(n17334), .ZN(U266) );
  OAI22_X1 U20407 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17349), .ZN(n17335) );
  INV_X1 U20408 ( .A(n17335), .ZN(U267) );
  AOI22_X1 U20409 ( .A1(n17348), .A2(n17336), .B1(n16187), .B2(U215), .ZN(U268) );
  OAI22_X1 U20410 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17349), .ZN(n17337) );
  INV_X1 U20411 ( .A(n17337), .ZN(U269) );
  OAI22_X1 U20412 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17349), .ZN(n17338) );
  INV_X1 U20413 ( .A(n17338), .ZN(U270) );
  OAI22_X1 U20414 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17349), .ZN(n17339) );
  INV_X1 U20415 ( .A(n17339), .ZN(U271) );
  OAI22_X1 U20416 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n17349), .ZN(n17340) );
  INV_X1 U20417 ( .A(n17340), .ZN(U272) );
  OAI22_X1 U20418 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n17348), .ZN(n17341) );
  INV_X1 U20419 ( .A(n17341), .ZN(U273) );
  OAI22_X1 U20420 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17349), .ZN(n17342) );
  INV_X1 U20421 ( .A(n17342), .ZN(U274) );
  OAI22_X1 U20422 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17349), .ZN(n17343) );
  INV_X1 U20423 ( .A(n17343), .ZN(U275) );
  OAI22_X1 U20424 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17348), .ZN(n17344) );
  INV_X1 U20425 ( .A(n17344), .ZN(U276) );
  OAI22_X1 U20426 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17348), .ZN(n17345) );
  INV_X1 U20427 ( .A(n17345), .ZN(U277) );
  OAI22_X1 U20428 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17348), .ZN(n17346) );
  INV_X1 U20429 ( .A(n17346), .ZN(U278) );
  OAI22_X1 U20430 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n17348), .ZN(n17347) );
  INV_X1 U20431 ( .A(n17347), .ZN(U279) );
  INV_X1 U20432 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n19491) );
  AOI22_X1 U20433 ( .A1(n17348), .A2(n19491), .B1(n16082), .B2(U215), .ZN(U280) );
  INV_X1 U20434 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n19488) );
  AOI22_X1 U20435 ( .A1(n17349), .A2(n19488), .B1(n16076), .B2(U215), .ZN(U281) );
  INV_X1 U20436 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19641) );
  AOI22_X1 U20437 ( .A1(n17349), .A2(n19486), .B1(n19641), .B2(U215), .ZN(U282) );
  INV_X1 U20438 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n18128) );
  AOI222_X1 U20439 ( .A1(n18128), .A2(P3_DATAO_REG_30__SCAN_IN), .B1(n19486), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n21268), .C2(
        P1_DATAO_REG_30__SCAN_IN), .ZN(n17350) );
  INV_X2 U20440 ( .A(n17352), .ZN(n17351) );
  INV_X1 U20441 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19268) );
  INV_X1 U20442 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20224) );
  AOI22_X1 U20443 ( .A1(n17351), .A2(n19268), .B1(n20224), .B2(n17352), .ZN(
        U347) );
  INV_X1 U20444 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19266) );
  INV_X1 U20445 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20222) );
  AOI22_X1 U20446 ( .A1(n17351), .A2(n19266), .B1(n20222), .B2(n17352), .ZN(
        U348) );
  INV_X1 U20447 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19263) );
  INV_X1 U20448 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20220) );
  AOI22_X1 U20449 ( .A1(n17351), .A2(n19263), .B1(n20220), .B2(n17352), .ZN(
        U349) );
  INV_X1 U20450 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19262) );
  INV_X1 U20451 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20218) );
  AOI22_X1 U20452 ( .A1(n17351), .A2(n19262), .B1(n20218), .B2(n17352), .ZN(
        U350) );
  INV_X1 U20453 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19259) );
  INV_X1 U20454 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20216) );
  AOI22_X1 U20455 ( .A1(n17351), .A2(n19259), .B1(n20216), .B2(n17352), .ZN(
        U351) );
  INV_X1 U20456 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19258) );
  INV_X1 U20457 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20214) );
  AOI22_X1 U20458 ( .A1(n17351), .A2(n19258), .B1(n20214), .B2(n17352), .ZN(
        U352) );
  INV_X1 U20459 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19256) );
  INV_X1 U20460 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20213) );
  AOI22_X1 U20461 ( .A1(n17351), .A2(n19256), .B1(n20213), .B2(n17352), .ZN(
        U353) );
  INV_X1 U20462 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19254) );
  AOI22_X1 U20463 ( .A1(n17351), .A2(n19254), .B1(n20212), .B2(n17352), .ZN(
        U354) );
  INV_X1 U20464 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19309) );
  INV_X1 U20465 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20261) );
  AOI22_X1 U20466 ( .A1(n17351), .A2(n19309), .B1(n20261), .B2(n17352), .ZN(
        U355) );
  INV_X1 U20467 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19305) );
  INV_X1 U20468 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20257) );
  AOI22_X1 U20469 ( .A1(n17351), .A2(n19305), .B1(n20257), .B2(n17352), .ZN(
        U356) );
  INV_X1 U20470 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19303) );
  INV_X1 U20471 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20255) );
  AOI22_X1 U20472 ( .A1(n17351), .A2(n19303), .B1(n20255), .B2(n17352), .ZN(
        U357) );
  INV_X1 U20473 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19300) );
  INV_X1 U20474 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20253) );
  AOI22_X1 U20475 ( .A1(n17351), .A2(n19300), .B1(n20253), .B2(n17352), .ZN(
        U358) );
  INV_X1 U20476 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19299) );
  INV_X1 U20477 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20252) );
  AOI22_X1 U20478 ( .A1(n17351), .A2(n19299), .B1(n20252), .B2(n17352), .ZN(
        U359) );
  INV_X1 U20479 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19297) );
  INV_X1 U20480 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20250) );
  AOI22_X1 U20481 ( .A1(n17351), .A2(n19297), .B1(n20250), .B2(n17352), .ZN(
        U360) );
  INV_X1 U20482 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19295) );
  INV_X1 U20483 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20249) );
  AOI22_X1 U20484 ( .A1(n17351), .A2(n19295), .B1(n20249), .B2(n17352), .ZN(
        U361) );
  INV_X1 U20485 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19292) );
  INV_X1 U20486 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20247) );
  AOI22_X1 U20487 ( .A1(n17351), .A2(n19292), .B1(n20247), .B2(n17352), .ZN(
        U362) );
  INV_X1 U20488 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19291) );
  INV_X1 U20489 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20246) );
  AOI22_X1 U20490 ( .A1(n17351), .A2(n19291), .B1(n20246), .B2(n17352), .ZN(
        U363) );
  INV_X1 U20491 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19288) );
  INV_X1 U20492 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20244) );
  AOI22_X1 U20493 ( .A1(n17351), .A2(n19288), .B1(n20244), .B2(n17352), .ZN(
        U364) );
  INV_X1 U20494 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n19253) );
  INV_X1 U20495 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20210) );
  AOI22_X1 U20496 ( .A1(n17351), .A2(n19253), .B1(n20210), .B2(n17352), .ZN(
        U365) );
  INV_X1 U20497 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19287) );
  INV_X1 U20498 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20242) );
  AOI22_X1 U20499 ( .A1(n17351), .A2(n19287), .B1(n20242), .B2(n17352), .ZN(
        U366) );
  INV_X1 U20500 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n21368) );
  INV_X1 U20501 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20240) );
  AOI22_X1 U20502 ( .A1(n17351), .A2(n21368), .B1(n20240), .B2(n17352), .ZN(
        U367) );
  INV_X1 U20503 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19284) );
  INV_X1 U20504 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20238) );
  AOI22_X1 U20505 ( .A1(n17351), .A2(n19284), .B1(n20238), .B2(n17352), .ZN(
        U368) );
  INV_X1 U20506 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19281) );
  INV_X1 U20507 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20236) );
  AOI22_X1 U20508 ( .A1(n17351), .A2(n19281), .B1(n20236), .B2(n17352), .ZN(
        U369) );
  INV_X1 U20509 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19280) );
  INV_X1 U20510 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20234) );
  AOI22_X1 U20511 ( .A1(n17351), .A2(n19280), .B1(n20234), .B2(n17352), .ZN(
        U370) );
  INV_X1 U20512 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19278) );
  INV_X1 U20513 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20232) );
  AOI22_X1 U20514 ( .A1(n17351), .A2(n19278), .B1(n20232), .B2(n17352), .ZN(
        U371) );
  INV_X1 U20515 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19276) );
  INV_X1 U20516 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20231) );
  AOI22_X1 U20517 ( .A1(n17351), .A2(n19276), .B1(n20231), .B2(n17352), .ZN(
        U372) );
  INV_X1 U20518 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19274) );
  INV_X1 U20519 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20229) );
  AOI22_X1 U20520 ( .A1(n17351), .A2(n19274), .B1(n20229), .B2(n17352), .ZN(
        U373) );
  INV_X1 U20521 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19272) );
  INV_X1 U20522 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20227) );
  AOI22_X1 U20523 ( .A1(n17351), .A2(n19272), .B1(n20227), .B2(n17352), .ZN(
        U374) );
  INV_X1 U20524 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19270) );
  INV_X1 U20525 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20225) );
  AOI22_X1 U20526 ( .A1(n17351), .A2(n19270), .B1(n20225), .B2(n17352), .ZN(
        U375) );
  INV_X1 U20527 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n19250) );
  INV_X1 U20528 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20209) );
  AOI22_X1 U20529 ( .A1(n17351), .A2(n19250), .B1(n20209), .B2(n17352), .ZN(
        U376) );
  NAND2_X1 U20530 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n21319), .ZN(n19240) );
  NAND2_X1 U20531 ( .A1(n19235), .A2(n17353), .ZN(n19236) );
  OAI21_X1 U20532 ( .B1(n19240), .B2(n17353), .A(n19236), .ZN(n19319) );
  AOI21_X1 U20533 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n19319), .ZN(n17354) );
  INV_X1 U20534 ( .A(n17354), .ZN(P3_U2633) );
  NAND2_X1 U20535 ( .A1(n19350), .A2(n19349), .ZN(n17357) );
  OAI21_X1 U20536 ( .B1(n17355), .B2(n18173), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n17356) );
  OAI21_X1 U20537 ( .B1(n17357), .B2(n19338), .A(n17356), .ZN(P3_U2634) );
  INV_X1 U20538 ( .A(n19234), .ZN(n17359) );
  AOI22_X1 U20539 ( .A1(P3_D_C_N_REG_SCAN_IN), .A2(n19347), .B1(n17359), .B2(
        n19235), .ZN(n17358) );
  OAI21_X1 U20540 ( .B1(P3_CODEFETCH_REG_SCAN_IN), .B2(n19347), .A(n17358), 
        .ZN(P3_U2635) );
  OAI21_X1 U20541 ( .B1(n17359), .B2(BS16), .A(n19319), .ZN(n19317) );
  OAI21_X1 U20542 ( .B1(n19319), .B2(n21312), .A(n19317), .ZN(P3_U2636) );
  NAND3_X1 U20543 ( .A1(n17361), .A2(n19185), .A3(n17360), .ZN(n19204) );
  AND2_X1 U20544 ( .A1(n19214), .A2(n19204), .ZN(n19331) );
  INV_X1 U20545 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n21335) );
  OAI21_X1 U20546 ( .B1(n19331), .B2(n21335), .A(n17362), .ZN(P3_U2637) );
  NOR4_X1 U20547 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n17366) );
  NOR4_X1 U20548 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n17365) );
  NOR4_X1 U20549 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n17364) );
  NOR4_X1 U20550 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n17363) );
  NAND4_X1 U20551 ( .A1(n17366), .A2(n17365), .A3(n17364), .A4(n17363), .ZN(
        n17372) );
  NOR4_X1 U20552 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n17370) );
  AOI211_X1 U20553 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_13__SCAN_IN), .B(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n17369) );
  NOR4_X1 U20554 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n17368) );
  NOR4_X1 U20555 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n17367) );
  NAND4_X1 U20556 ( .A1(n17370), .A2(n17369), .A3(n17368), .A4(n17367), .ZN(
        n17371) );
  NOR2_X1 U20557 ( .A1(n17372), .A2(n17371), .ZN(n19329) );
  INV_X1 U20558 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n17374) );
  NOR3_X1 U20559 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n17375) );
  OAI21_X1 U20560 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n17375), .A(n19329), .ZN(
        n17373) );
  OAI21_X1 U20561 ( .B1(n19329), .B2(n17374), .A(n17373), .ZN(P3_U2638) );
  INV_X1 U20562 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19318) );
  AOI21_X1 U20563 ( .B1(n19251), .B2(n19318), .A(n17375), .ZN(n17377) );
  INV_X1 U20564 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n17376) );
  INV_X1 U20565 ( .A(n19329), .ZN(n19326) );
  AOI22_X1 U20566 ( .A1(n19329), .A2(n17377), .B1(n17376), .B2(n19326), .ZN(
        P3_U2639) );
  INV_X1 U20567 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n17397) );
  INV_X1 U20568 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n19307) );
  INV_X1 U20569 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n19294) );
  NOR4_X1 U20570 ( .A1(n19289), .A2(n19290), .A3(n17379), .A4(n17378), .ZN(
        n17475) );
  NAND2_X1 U20571 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n17475), .ZN(n17470) );
  NOR2_X1 U20572 ( .A1(n19294), .A2(n17470), .ZN(n17390) );
  NAND2_X1 U20573 ( .A1(n17658), .A2(n17390), .ZN(n17455) );
  NAND2_X1 U20574 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .ZN(n17380) );
  NAND4_X1 U20575 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n17420), .ZN(n17389) );
  NOR3_X1 U20576 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n19307), .A3(n17389), 
        .ZN(n17381) );
  AOI21_X1 U20577 ( .B1(n17725), .B2(P3_EBX_REG_31__SCAN_IN), .A(n17381), .ZN(
        n17396) );
  INV_X1 U20578 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n17864) );
  NAND2_X1 U20579 ( .A1(n17481), .A2(n17864), .ZN(n17480) );
  INV_X1 U20580 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n17865) );
  NAND2_X1 U20581 ( .A1(n17462), .A2(n17865), .ZN(n17458) );
  NOR2_X2 U20582 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17458), .ZN(n17443) );
  INV_X1 U20583 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17439) );
  NAND2_X1 U20584 ( .A1(n17443), .A2(n17439), .ZN(n17438) );
  INV_X1 U20585 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17737) );
  NAND2_X1 U20586 ( .A1(n17421), .A2(n17737), .ZN(n17398) );
  NOR2_X1 U20587 ( .A1(n17687), .A2(n17398), .ZN(n17404) );
  INV_X1 U20588 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17742) );
  NOR2_X1 U20589 ( .A1(n17463), .A2(n17695), .ZN(n17453) );
  NAND2_X1 U20590 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18239), .ZN(
        n17385) );
  OAI21_X1 U20591 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n17383), .A(
        n17385), .ZN(n18254) );
  INV_X1 U20592 ( .A(n18254), .ZN(n17454) );
  NOR2_X1 U20593 ( .A1(n17453), .A2(n17454), .ZN(n17452) );
  NOR2_X1 U20594 ( .A1(n17452), .A2(n17695), .ZN(n17444) );
  INV_X1 U20595 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17386) );
  AOI21_X1 U20596 ( .B1(n17386), .B2(n17385), .A(n17384), .ZN(n18240) );
  NOR2_X1 U20597 ( .A1(n17444), .A2(n18240), .ZN(n17445) );
  NOR2_X1 U20598 ( .A1(n17445), .A2(n17695), .ZN(n17432) );
  INV_X1 U20599 ( .A(n17387), .ZN(n17433) );
  INV_X1 U20600 ( .A(n17695), .ZN(n17388) );
  NOR2_X1 U20601 ( .A1(n17423), .A2(n17424), .ZN(n17422) );
  NOR2_X1 U20602 ( .A1(n17422), .A2(n17695), .ZN(n17409) );
  NAND2_X1 U20603 ( .A1(n17388), .A2(n19228), .ZN(n17727) );
  NOR3_X1 U20604 ( .A1(n17400), .A2(n17399), .A3(n17727), .ZN(n17394) );
  NOR2_X1 U20605 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n17389), .ZN(n17403) );
  INV_X1 U20606 ( .A(n17403), .ZN(n17392) );
  NAND3_X1 U20607 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n17391) );
  NAND4_X1 U20608 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(P3_REIP_REG_26__SCAN_IN), 
        .A3(n17390), .A4(n17644), .ZN(n17419) );
  OAI21_X1 U20609 ( .B1(n17391), .B2(n17419), .A(n17645), .ZN(n17411) );
  AOI21_X1 U20610 ( .B1(n17392), .B2(n17411), .A(n19310), .ZN(n17393) );
  OAI211_X1 U20611 ( .C1(n17397), .C2(n17726), .A(n17396), .B(n17395), .ZN(
        P3_U2640) );
  NAND2_X1 U20612 ( .A1(n17724), .A2(n17398), .ZN(n17417) );
  OAI22_X1 U20613 ( .A1(n17401), .A2(n17726), .B1(n19307), .B2(n17411), .ZN(
        n17402) );
  OAI21_X1 U20614 ( .B1(n17725), .B2(n17404), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n17405) );
  OAI211_X1 U20615 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n17417), .A(n17406), .B(
        n17405), .ZN(P3_U2641) );
  NOR2_X1 U20616 ( .A1(n17421), .A2(n17737), .ZN(n17418) );
  INV_X1 U20617 ( .A(n17407), .ZN(n17408) );
  AOI211_X1 U20618 ( .C1(n17410), .C2(n17409), .A(n17408), .B(n9767), .ZN(
        n17414) );
  INV_X1 U20619 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n19304) );
  OAI22_X1 U20620 ( .A1(n17412), .A2(n17726), .B1(n19304), .B2(n17411), .ZN(
        n17413) );
  AOI211_X1 U20621 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n17725), .A(n17414), .B(
        n17413), .ZN(n17416) );
  NAND4_X1 U20622 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n17420), .A4(n19304), .ZN(n17415) );
  OAI211_X1 U20623 ( .C1(n17418), .C2(n17417), .A(n17416), .B(n17415), .ZN(
        P3_U2642) );
  NAND2_X1 U20624 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n17420), .ZN(n17430) );
  AOI22_X1 U20625 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17700), .B1(
        n17725), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n17429) );
  NAND2_X1 U20626 ( .A1(n17645), .A2(n17419), .ZN(n17450) );
  NAND2_X1 U20627 ( .A1(n17420), .A2(n19301), .ZN(n17434) );
  NAND2_X1 U20628 ( .A1(n17450), .A2(n17434), .ZN(n17427) );
  AOI211_X1 U20629 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n17438), .A(n17421), .B(
        n17687), .ZN(n17426) );
  AOI211_X1 U20630 ( .C1(n17424), .C2(n17423), .A(n17422), .B(n9767), .ZN(
        n17425) );
  AOI211_X1 U20631 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n17427), .A(n17426), 
        .B(n17425), .ZN(n17428) );
  OAI211_X1 U20632 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n17430), .A(n17429), 
        .B(n17428), .ZN(P3_U2643) );
  AOI211_X1 U20633 ( .C1(n17433), .C2(n17432), .A(n17431), .B(n9767), .ZN(
        n17437) );
  INV_X1 U20634 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17435) );
  OAI21_X1 U20635 ( .B1(n17726), .B2(n17435), .A(n17434), .ZN(n17436) );
  AOI211_X1 U20636 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n17725), .A(n17437), .B(
        n17436), .ZN(n17441) );
  OAI211_X1 U20637 ( .C1(n17443), .C2(n17439), .A(n17724), .B(n17438), .ZN(
        n17440) );
  OAI211_X1 U20638 ( .C1(n17450), .C2(n19301), .A(n17441), .B(n17440), .ZN(
        P3_U2644) );
  INV_X1 U20639 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n19296) );
  INV_X1 U20640 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n19298) );
  OAI21_X1 U20641 ( .B1(n19296), .B2(n17455), .A(n19298), .ZN(n17442) );
  INV_X1 U20642 ( .A(n17442), .ZN(n17451) );
  AOI22_X1 U20643 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17700), .B1(
        n17725), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n17449) );
  AOI211_X1 U20644 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n17458), .A(n17443), .B(
        n17687), .ZN(n17447) );
  AOI211_X1 U20645 ( .C1(n18240), .C2(n17444), .A(n17445), .B(n9767), .ZN(
        n17446) );
  NOR2_X1 U20646 ( .A1(n17447), .A2(n17446), .ZN(n17448) );
  OAI211_X1 U20647 ( .C1(n17451), .C2(n17450), .A(n17449), .B(n17448), .ZN(
        P3_U2645) );
  NAND2_X1 U20648 ( .A1(n17658), .A2(n17470), .ZN(n17476) );
  NAND2_X1 U20649 ( .A1(n17644), .A2(n17476), .ZN(n17471) );
  AOI21_X1 U20650 ( .B1(n17658), .B2(n19294), .A(n17471), .ZN(n17461) );
  AOI211_X1 U20651 ( .C1(n17454), .C2(n17453), .A(n17452), .B(n9767), .ZN(
        n17457) );
  OAI22_X1 U20652 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n17455), .B1(n17865), 
        .B2(n17706), .ZN(n17456) );
  AOI211_X1 U20653 ( .C1(n17700), .C2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n17457), .B(n17456), .ZN(n17460) );
  OAI211_X1 U20654 ( .C1(n17462), .C2(n17865), .A(n17724), .B(n17458), .ZN(
        n17459) );
  OAI211_X1 U20655 ( .C1(n17461), .C2(n19296), .A(n17460), .B(n17459), .ZN(
        P3_U2646) );
  NAND2_X1 U20656 ( .A1(n17658), .A2(n19294), .ZN(n17469) );
  AOI22_X1 U20657 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n17700), .B1(
        n17725), .B2(P3_EBX_REG_24__SCAN_IN), .ZN(n17468) );
  AOI211_X1 U20658 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n17480), .A(n17462), .B(
        n17687), .ZN(n17466) );
  AOI211_X1 U20659 ( .C1(n17464), .C2(n9747), .A(n17463), .B(n9767), .ZN(
        n17465) );
  AOI211_X1 U20660 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n17471), .A(n17466), 
        .B(n17465), .ZN(n17467) );
  OAI211_X1 U20661 ( .C1(n17470), .C2(n17469), .A(n17468), .B(n17467), .ZN(
        P3_U2647) );
  INV_X1 U20662 ( .A(n17471), .ZN(n17484) );
  AOI211_X1 U20663 ( .C1(n17474), .C2(n17473), .A(n17472), .B(n9767), .ZN(
        n17479) );
  INV_X1 U20664 ( .A(n17475), .ZN(n17477) );
  OAI22_X1 U20665 ( .A1(n17706), .A2(n17864), .B1(n17477), .B2(n17476), .ZN(
        n17478) );
  AOI211_X1 U20666 ( .C1(n17700), .C2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n17479), .B(n17478), .ZN(n17483) );
  OAI211_X1 U20667 ( .C1(n17481), .C2(n17864), .A(n17724), .B(n17480), .ZN(
        n17482) );
  OAI211_X1 U20668 ( .C1(n17484), .C2(n19293), .A(n17483), .B(n17482), .ZN(
        P3_U2648) );
  AOI211_X1 U20669 ( .C1(n18288), .C2(n17486), .A(n17485), .B(n9767), .ZN(
        n17490) );
  OAI211_X1 U20670 ( .C1(n17495), .C2(n17927), .A(n17724), .B(n17487), .ZN(
        n17488) );
  OAI21_X1 U20671 ( .B1(n17927), .B2(n17706), .A(n17488), .ZN(n17489) );
  AOI211_X1 U20672 ( .C1(n17700), .C2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n17490), .B(n17489), .ZN(n17491) );
  OAI221_X1 U20673 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(n17492), .C1(n19289), 
        .C2(n17501), .A(n17491), .ZN(P3_U2650) );
  AOI22_X1 U20674 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n17700), .B1(
        n17725), .B2(P3_EBX_REG_20__SCAN_IN), .ZN(n17500) );
  NAND2_X1 U20675 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n17511) );
  NOR2_X1 U20676 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n17511), .ZN(n17498) );
  AOI211_X1 U20677 ( .C1(n18306), .C2(n17494), .A(n17493), .B(n9767), .ZN(
        n17497) );
  AOI211_X1 U20678 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17509), .A(n17495), .B(
        n17687), .ZN(n17496) );
  AOI211_X1 U20679 ( .C1(n17498), .C2(n17517), .A(n17497), .B(n17496), .ZN(
        n17499) );
  OAI211_X1 U20680 ( .C1(n19286), .C2(n17501), .A(n17500), .B(n17499), .ZN(
        P3_U2651) );
  NAND2_X1 U20681 ( .A1(n17645), .A2(n17502), .ZN(n17530) );
  INV_X1 U20682 ( .A(n17530), .ZN(n17521) );
  NOR2_X1 U20683 ( .A1(n17709), .A2(n9751), .ZN(n18314) );
  NAND2_X1 U20684 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18314), .ZN(
        n17515) );
  AOI21_X1 U20685 ( .B1(n17503), .B2(n17728), .A(n17695), .ZN(n17540) );
  AOI21_X1 U20686 ( .B1(n17388), .B2(n17515), .A(n17540), .ZN(n17506) );
  INV_X1 U20687 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n21269) );
  AOI21_X1 U20688 ( .B1(n21269), .B2(n17515), .A(n18273), .ZN(n17504) );
  INV_X1 U20689 ( .A(n17504), .ZN(n18318) );
  OAI21_X1 U20690 ( .B1(n17506), .B2(n18318), .A(n19228), .ZN(n17505) );
  AOI21_X1 U20691 ( .B1(n17506), .B2(n18318), .A(n17505), .ZN(n17508) );
  OAI22_X1 U20692 ( .A1(n21269), .A2(n17726), .B1(n17706), .B2(n17510), .ZN(
        n17507) );
  AOI211_X1 U20693 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(n17521), .A(n17508), 
        .B(n17507), .ZN(n17514) );
  OAI211_X1 U20694 ( .C1(n17519), .C2(n17510), .A(n17724), .B(n17509), .ZN(
        n17513) );
  OAI211_X1 U20695 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(P3_REIP_REG_18__SCAN_IN), .A(n17517), .B(n17511), .ZN(n17512) );
  NAND4_X1 U20696 ( .A1(n17514), .A2(n18739), .A3(n17513), .A4(n17512), .ZN(
        P3_U2652) );
  AOI22_X1 U20697 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17700), .B1(
        n17725), .B2(P3_EBX_REG_18__SCAN_IN), .ZN(n17524) );
  AOI21_X1 U20698 ( .B1(n18314), .B2(n17728), .A(n17695), .ZN(n17516) );
  OAI21_X1 U20699 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n18314), .A(
        n17515), .ZN(n18324) );
  XNOR2_X1 U20700 ( .A(n17516), .B(n18324), .ZN(n17518) );
  AOI22_X1 U20701 ( .A1(n19228), .A2(n17518), .B1(n17517), .B2(n19283), .ZN(
        n17523) );
  AOI211_X1 U20702 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n17533), .A(n17519), .B(
        n17687), .ZN(n17520) );
  AOI211_X1 U20703 ( .C1(P3_REIP_REG_18__SCAN_IN), .C2(n17521), .A(n18693), 
        .B(n17520), .ZN(n17522) );
  NAND3_X1 U20704 ( .A1(n17524), .A2(n17523), .A3(n17522), .ZN(P3_U2653) );
  INV_X1 U20705 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17537) );
  AOI21_X1 U20706 ( .B1(n17658), .B2(n17525), .A(P3_REIP_REG_17__SCAN_IN), 
        .ZN(n17531) );
  INV_X1 U20707 ( .A(n18314), .ZN(n17526) );
  OAI21_X1 U20708 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n17527), .A(
        n17526), .ZN(n18339) );
  OAI21_X1 U20709 ( .B1(n17541), .B2(n17540), .A(n17388), .ZN(n17528) );
  XNOR2_X1 U20710 ( .A(n18339), .B(n17528), .ZN(n17529) );
  OAI22_X1 U20711 ( .A1(n17531), .A2(n17530), .B1(n9767), .B2(n17529), .ZN(
        n17532) );
  AOI211_X1 U20712 ( .C1(n17725), .C2(P3_EBX_REG_17__SCAN_IN), .A(n18693), .B(
        n17532), .ZN(n17536) );
  OAI211_X1 U20713 ( .C1(n17542), .C2(n17534), .A(n17724), .B(n17533), .ZN(
        n17535) );
  OAI211_X1 U20714 ( .C1(n17726), .C2(n17537), .A(n17536), .B(n17535), .ZN(
        P3_U2654) );
  AOI221_X1 U20715 ( .B1(n19277), .B2(n17658), .C1(n17564), .C2(n17658), .A(
        n17721), .ZN(n17547) );
  NOR4_X1 U20716 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n17729), .A3(n19277), 
        .A4(n17564), .ZN(n17538) );
  AOI211_X1 U20717 ( .C1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n17700), .A(
        n18693), .B(n17538), .ZN(n17546) );
  NOR2_X1 U20718 ( .A1(n17541), .A2(n17540), .ZN(n17539) );
  AOI211_X1 U20719 ( .C1(n17541), .C2(n17540), .A(n17539), .B(n9767), .ZN(
        n17544) );
  AOI211_X1 U20720 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17557), .A(n17542), .B(
        n17687), .ZN(n17543) );
  AOI211_X1 U20721 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17725), .A(n17544), .B(
        n17543), .ZN(n17545) );
  OAI211_X1 U20722 ( .C1(n17547), .C2(n19279), .A(n17546), .B(n17545), .ZN(
        P3_U2655) );
  AOI21_X1 U20723 ( .B1(n17564), .B2(n17658), .A(n17721), .ZN(n17571) );
  INV_X1 U20724 ( .A(n17571), .ZN(n17556) );
  OAI21_X1 U20725 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17548), .A(
        n17388), .ZN(n17551) );
  OAI21_X1 U20726 ( .B1(n17551), .B2(n17550), .A(n19228), .ZN(n17549) );
  AOI21_X1 U20727 ( .B1(n17551), .B2(n17550), .A(n17549), .ZN(n17555) );
  NOR2_X1 U20728 ( .A1(n17729), .A2(n17564), .ZN(n17552) );
  NAND2_X1 U20729 ( .A1(n17552), .A2(n19277), .ZN(n17553) );
  OAI211_X1 U20730 ( .C1(n17706), .C2(n21278), .A(n18739), .B(n17553), .ZN(
        n17554) );
  AOI211_X1 U20731 ( .C1(n17556), .C2(P3_REIP_REG_15__SCAN_IN), .A(n17555), 
        .B(n17554), .ZN(n17559) );
  OAI211_X1 U20732 ( .C1(n17561), .C2(n21278), .A(n17724), .B(n17557), .ZN(
        n17558) );
  OAI211_X1 U20733 ( .C1(n17726), .C2(n17560), .A(n17559), .B(n17558), .ZN(
        P3_U2656) );
  INV_X1 U20734 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n19275) );
  AOI21_X1 U20735 ( .B1(n17725), .B2(P3_EBX_REG_14__SCAN_IN), .A(n18693), .ZN(
        n17570) );
  AOI211_X1 U20736 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17581), .A(n17561), .B(
        n17687), .ZN(n17568) );
  OR2_X1 U20737 ( .A1(n18373), .A2(n18369), .ZN(n17573) );
  AOI21_X1 U20738 ( .B1(n18354), .B2(n17573), .A(n17562), .ZN(n18356) );
  OAI21_X1 U20739 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17573), .A(
        n17388), .ZN(n17563) );
  XOR2_X1 U20740 ( .A(n18356), .B(n17563), .Z(n17566) );
  INV_X1 U20741 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n19273) );
  NAND3_X1 U20742 ( .A1(n17564), .A2(n17658), .A3(n17572), .ZN(n17565) );
  OAI22_X1 U20743 ( .A1(n9767), .A2(n17566), .B1(n19273), .B2(n17565), .ZN(
        n17567) );
  AOI211_X1 U20744 ( .C1(n17700), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n17568), .B(n17567), .ZN(n17569) );
  OAI211_X1 U20745 ( .C1(n19275), .C2(n17571), .A(n17570), .B(n17569), .ZN(
        P3_U2657) );
  INV_X1 U20746 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17585) );
  NAND2_X1 U20747 ( .A1(n17658), .A2(n17572), .ZN(n17579) );
  INV_X1 U20748 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n19271) );
  OAI21_X1 U20749 ( .B1(n17591), .B2(n17729), .A(n17644), .ZN(n17586) );
  AOI21_X1 U20750 ( .B1(n17658), .B2(n19271), .A(n17586), .ZN(n17578) );
  INV_X1 U20751 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n18387) );
  NOR2_X1 U20752 ( .A1(n18387), .A2(n18369), .ZN(n17588) );
  OAI21_X1 U20753 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17588), .A(
        n17573), .ZN(n18376) );
  INV_X1 U20754 ( .A(n17588), .ZN(n17574) );
  OAI21_X1 U20755 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17574), .A(
        n17388), .ZN(n17576) );
  AOI21_X1 U20756 ( .B1(n18376), .B2(n17576), .A(n9767), .ZN(n17575) );
  OAI21_X1 U20757 ( .B1(n18376), .B2(n17576), .A(n17575), .ZN(n17577) );
  OAI221_X1 U20758 ( .B1(P3_REIP_REG_13__SCAN_IN), .B2(n17579), .C1(n19273), 
        .C2(n17578), .A(n17577), .ZN(n17580) );
  AOI211_X1 U20759 ( .C1(n17725), .C2(P3_EBX_REG_13__SCAN_IN), .A(n18693), .B(
        n17580), .ZN(n17584) );
  OAI211_X1 U20760 ( .C1(n17587), .C2(n17582), .A(n17724), .B(n17581), .ZN(
        n17583) );
  OAI211_X1 U20761 ( .C1(n17726), .C2(n17585), .A(n17584), .B(n17583), .ZN(
        P3_U2658) );
  INV_X1 U20762 ( .A(n17586), .ZN(n17600) );
  AOI211_X1 U20763 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17603), .A(n17587), .B(
        n17687), .ZN(n17595) );
  AOI21_X1 U20764 ( .B1(n18387), .B2(n18369), .A(n17588), .ZN(n18390) );
  AOI21_X1 U20765 ( .B1(n16961), .B2(n17711), .A(n17695), .ZN(n17589) );
  XOR2_X1 U20766 ( .A(n18390), .B(n17589), .Z(n17592) );
  NOR2_X1 U20767 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17729), .ZN(n17590) );
  AOI22_X1 U20768 ( .A1(n19228), .A2(n17592), .B1(n17591), .B2(n17590), .ZN(
        n17593) );
  OAI211_X1 U20769 ( .C1(n18387), .C2(n17726), .A(n17593), .B(n18739), .ZN(
        n17594) );
  AOI211_X1 U20770 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17725), .A(n17595), .B(
        n17594), .ZN(n17596) );
  OAI21_X1 U20771 ( .B1(n19271), .B2(n17600), .A(n17596), .ZN(P3_U2659) );
  NAND2_X1 U20772 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_9__SCAN_IN), 
        .ZN(n17612) );
  INV_X1 U20773 ( .A(n17612), .ZN(n17597) );
  NOR2_X1 U20774 ( .A1(n17729), .A2(n17630), .ZN(n17626) );
  AOI21_X1 U20775 ( .B1(n17597), .B2(n17626), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n17601) );
  NAND2_X1 U20776 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17619), .ZN(
        n17618) );
  NOR2_X1 U20777 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17618), .ZN(
        n17610) );
  AOI21_X1 U20778 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17610), .A(
        n17695), .ZN(n17598) );
  NOR2_X1 U20779 ( .A1(n18421), .A2(n17618), .ZN(n17609) );
  OAI21_X1 U20780 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17609), .A(
        n18369), .ZN(n18419) );
  XOR2_X1 U20781 ( .A(n17598), .B(n18419), .Z(n17599) );
  OAI22_X1 U20782 ( .A1(n17601), .A2(n17600), .B1(n9767), .B2(n17599), .ZN(
        n17602) );
  AOI211_X1 U20783 ( .C1(n17725), .C2(P3_EBX_REG_11__SCAN_IN), .A(n18693), .B(
        n17602), .ZN(n17606) );
  OAI211_X1 U20784 ( .C1(n17607), .C2(n17604), .A(n17724), .B(n17603), .ZN(
        n17605) );
  OAI211_X1 U20785 ( .C1(n17726), .C2(n18402), .A(n17606), .B(n17605), .ZN(
        P3_U2660) );
  AOI211_X1 U20786 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17608), .A(n17607), .B(
        n17687), .ZN(n17616) );
  AOI21_X1 U20787 ( .B1(n17658), .B2(n17630), .A(n17721), .ZN(n17643) );
  AOI21_X1 U20788 ( .B1(n18421), .B2(n17618), .A(n17609), .ZN(n18427) );
  NOR2_X1 U20789 ( .A1(n17610), .A2(n17695), .ZN(n17620) );
  AOI21_X1 U20790 ( .B1(n18427), .B2(n17620), .A(n9767), .ZN(n17611) );
  OAI21_X1 U20791 ( .B1(n18427), .B2(n17620), .A(n17611), .ZN(n17614) );
  OAI211_X1 U20792 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(P3_REIP_REG_9__SCAN_IN), 
        .A(n17626), .B(n17612), .ZN(n17613) );
  OAI211_X1 U20793 ( .C1(n17643), .C2(n19267), .A(n17614), .B(n17613), .ZN(
        n17615) );
  AOI211_X1 U20794 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17725), .A(n17616), .B(
        n17615), .ZN(n17617) );
  OAI211_X1 U20795 ( .C1(n18421), .C2(n17726), .A(n17617), .B(n18739), .ZN(
        P3_U2661) );
  AOI21_X1 U20796 ( .B1(n17724), .B2(n17631), .A(n17725), .ZN(n17629) );
  OAI21_X1 U20797 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17619), .A(
        n17618), .ZN(n18444) );
  INV_X1 U20798 ( .A(n17620), .ZN(n17622) );
  AOI211_X1 U20799 ( .C1(n18440), .C2(n17728), .A(n17695), .B(n18444), .ZN(
        n17621) );
  AOI211_X1 U20800 ( .C1(n18444), .C2(n17622), .A(n17621), .B(n9767), .ZN(
        n17623) );
  AOI211_X1 U20801 ( .C1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n17700), .A(
        n18693), .B(n17623), .ZN(n17628) );
  INV_X1 U20802 ( .A(n17643), .ZN(n17625) );
  NOR3_X1 U20803 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n17631), .A3(n17687), .ZN(
        n17624) );
  AOI221_X1 U20804 ( .B1(n17626), .B2(n19265), .C1(n17625), .C2(
        P3_REIP_REG_9__SCAN_IN), .A(n17624), .ZN(n17627) );
  OAI211_X1 U20805 ( .C1(n17629), .C2(n21250), .A(n17628), .B(n17627), .ZN(
        P3_U2662) );
  AND2_X1 U20806 ( .A1(n17630), .A2(n17658), .ZN(n17641) );
  AOI211_X1 U20807 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17652), .A(n17631), .B(
        n17687), .ZN(n17639) );
  NOR2_X1 U20808 ( .A1(n17632), .A2(n17691), .ZN(n17662) );
  AOI21_X1 U20809 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n17662), .A(
        n17695), .ZN(n17633) );
  XOR2_X1 U20810 ( .A(n17634), .B(n17633), .Z(n17635) );
  AOI22_X1 U20811 ( .A1(n17725), .A2(P3_EBX_REG_8__SCAN_IN), .B1(n19228), .B2(
        n17635), .ZN(n17636) );
  OAI211_X1 U20812 ( .C1(n17637), .C2(n17726), .A(n17636), .B(n18739), .ZN(
        n17638) );
  AOI211_X1 U20813 ( .C1(n17641), .C2(n17640), .A(n17639), .B(n17638), .ZN(
        n17642) );
  OAI21_X1 U20814 ( .B1(n17643), .B2(n19264), .A(n17642), .ZN(P3_U2663) );
  NAND3_X1 U20815 ( .A1(n17658), .A2(P3_REIP_REG_6__SCAN_IN), .A3(n17657), 
        .ZN(n17650) );
  NAND2_X1 U20816 ( .A1(n17657), .A2(n17644), .ZN(n17683) );
  OAI21_X1 U20817 ( .B1(n13987), .B2(n17683), .A(n17645), .ZN(n17670) );
  NOR2_X1 U20818 ( .A1(n17662), .A2(n17695), .ZN(n17647) );
  AOI21_X1 U20819 ( .B1(n17648), .B2(n17647), .A(n9767), .ZN(n17646) );
  OAI21_X1 U20820 ( .B1(n17648), .B2(n17647), .A(n17646), .ZN(n17649) );
  OAI221_X1 U20821 ( .B1(P3_REIP_REG_7__SCAN_IN), .B2(n17650), .C1(n19260), 
        .C2(n17670), .A(n17649), .ZN(n17651) );
  AOI211_X1 U20822 ( .C1(n17725), .C2(P3_EBX_REG_7__SCAN_IN), .A(n18693), .B(
        n17651), .ZN(n17655) );
  OAI211_X1 U20823 ( .C1(n17659), .C2(n17653), .A(n17724), .B(n17652), .ZN(
        n17654) );
  OAI211_X1 U20824 ( .C1(n17726), .C2(n17656), .A(n17655), .B(n17654), .ZN(
        P3_U2664) );
  AOI21_X1 U20825 ( .B1(n17658), .B2(n17657), .A(P3_REIP_REG_6__SCAN_IN), .ZN(
        n17671) );
  AOI22_X1 U20826 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17700), .B1(
        n17725), .B2(P3_EBX_REG_6__SCAN_IN), .ZN(n17669) );
  AOI211_X1 U20827 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17678), .A(n17659), .B(
        n17687), .ZN(n17667) );
  OAI21_X1 U20828 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17661), .A(
        n17660), .ZN(n18460) );
  INV_X1 U20829 ( .A(n18460), .ZN(n17663) );
  NOR3_X1 U20830 ( .A1(n17663), .A2(n17662), .A3(n17727), .ZN(n17666) );
  NAND2_X1 U20831 ( .A1(n17388), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17664) );
  NAND2_X1 U20832 ( .A1(n19228), .A2(n17664), .ZN(n17730) );
  AOI211_X1 U20833 ( .C1(n17388), .C2(n17674), .A(n18460), .B(n17730), .ZN(
        n17665) );
  NOR4_X1 U20834 ( .A1(n18693), .A2(n17667), .A3(n17666), .A4(n17665), .ZN(
        n17668) );
  OAI211_X1 U20835 ( .C1(n17671), .C2(n17670), .A(n17669), .B(n17668), .ZN(
        P3_U2665) );
  OAI22_X1 U20836 ( .A1(n17673), .A2(n19257), .B1(n17729), .B2(n17672), .ZN(
        n17682) );
  OAI21_X1 U20837 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n17675), .A(
        n17674), .ZN(n18469) );
  AOI21_X1 U20838 ( .B1(n17728), .B2(n17675), .A(n17695), .ZN(n17676) );
  INV_X1 U20839 ( .A(n17676), .ZN(n17692) );
  AOI21_X1 U20840 ( .B1(n18469), .B2(n17692), .A(n9767), .ZN(n17677) );
  OAI21_X1 U20841 ( .B1(n18469), .B2(n17692), .A(n17677), .ZN(n17680) );
  OAI211_X1 U20842 ( .C1(n17688), .C2(n17992), .A(n17724), .B(n17678), .ZN(
        n17679) );
  OAI211_X1 U20843 ( .C1(n17992), .C2(n17706), .A(n17680), .B(n17679), .ZN(
        n17681) );
  AOI21_X1 U20844 ( .B1(n17683), .B2(n17682), .A(n17681), .ZN(n17684) );
  OAI211_X1 U20845 ( .C1(n18464), .C2(n17726), .A(n17684), .B(n18739), .ZN(
        P3_U2666) );
  NOR2_X1 U20846 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n17729), .ZN(n17685) );
  AOI22_X1 U20847 ( .A1(n17725), .A2(P3_EBX_REG_4__SCAN_IN), .B1(n17686), .B2(
        n17685), .ZN(n17702) );
  AOI211_X1 U20848 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17689), .A(n17688), .B(
        n17687), .ZN(n17699) );
  OAI22_X1 U20849 ( .A1(n17694), .A2(n17692), .B1(n17691), .B2(n17690), .ZN(
        n17693) );
  AOI21_X1 U20850 ( .B1(n17695), .B2(n17694), .A(n17693), .ZN(n17697) );
  OAI21_X1 U20851 ( .B1(n17948), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n19353), .ZN(n17696) );
  OAI211_X1 U20852 ( .C1(n17697), .C2(n9767), .A(n18739), .B(n17696), .ZN(
        n17698) );
  AOI211_X1 U20853 ( .C1(n17700), .C2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n17699), .B(n17698), .ZN(n17701) );
  OAI211_X1 U20854 ( .C1(n19255), .C2(n17703), .A(n17702), .B(n17701), .ZN(
        P3_U2667) );
  AOI22_X1 U20855 ( .A1(n17721), .A2(P3_REIP_REG_2__SCAN_IN), .B1(n19353), 
        .B2(n17704), .ZN(n17719) );
  INV_X1 U20856 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n19252) );
  AOI21_X1 U20857 ( .B1(n19251), .B2(n19252), .A(n17729), .ZN(n17717) );
  NOR2_X1 U20858 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17723) );
  OAI21_X1 U20859 ( .B1(n17723), .B2(n17705), .A(n17724), .ZN(n17707) );
  OAI22_X1 U20860 ( .A1(n17708), .A2(n17707), .B1(n17706), .B2(n17705), .ZN(
        n17715) );
  AOI22_X1 U20861 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18496), .B1(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17709), .ZN(n18489) );
  OAI21_X1 U20862 ( .B1(n17711), .B2(n18489), .A(n17710), .ZN(n17713) );
  AOI221_X1 U20863 ( .B1(n17388), .B2(n17713), .C1(n18489), .C2(n17713), .A(
        n9767), .ZN(n17714) );
  AOI211_X1 U20864 ( .C1(n17717), .C2(n17716), .A(n17715), .B(n17714), .ZN(
        n17718) );
  OAI211_X1 U20865 ( .C1(n18496), .C2(n17726), .A(n17719), .B(n17718), .ZN(
        P3_U2669) );
  AOI22_X1 U20866 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17721), .B1(n19353), 
        .B2(n17720), .ZN(n17735) );
  INV_X1 U20867 ( .A(n17722), .ZN(n18006) );
  NOR2_X1 U20868 ( .A1(n17723), .A2(n18006), .ZN(n18010) );
  AOI22_X1 U20869 ( .A1(n17725), .A2(P3_EBX_REG_1__SCAN_IN), .B1(n17724), .B2(
        n18010), .ZN(n17734) );
  OAI21_X1 U20870 ( .B1(n17728), .B2(n17727), .A(n17726), .ZN(n17732) );
  OAI22_X1 U20871 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17730), .B1(
        P3_REIP_REG_1__SCAN_IN), .B2(n17729), .ZN(n17731) );
  AOI21_X1 U20872 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17732), .A(
        n17731), .ZN(n17733) );
  NAND3_X1 U20873 ( .A1(n17735), .A2(n17734), .A3(n17733), .ZN(P3_U2670) );
  INV_X1 U20874 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n21262) );
  NAND4_X1 U20875 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(P3_EBX_REG_23__SCAN_IN), .A4(P3_EBX_REG_22__SCAN_IN), .ZN(n17736)
         );
  NOR4_X1 U20876 ( .A1(n17737), .A2(n21262), .A3(n17927), .A4(n17736), .ZN(
        n17738) );
  NAND4_X1 U20877 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .A3(n17862), .A4(n17738), .ZN(n17741) );
  NOR2_X1 U20878 ( .A1(n17742), .A2(n17741), .ZN(n17861) );
  NAND2_X1 U20879 ( .A1(n18013), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17740) );
  NAND2_X1 U20880 ( .A1(n17861), .A2(n17863), .ZN(n17739) );
  OAI22_X1 U20881 ( .A1(n17861), .A2(n17740), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17739), .ZN(P3_U2672) );
  NAND2_X1 U20882 ( .A1(n17742), .A2(n17741), .ZN(n17743) );
  NAND2_X1 U20883 ( .A1(n17743), .A2(n18013), .ZN(n17860) );
  AOI22_X1 U20884 ( .A1(n17948), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17947), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17747) );
  AOI22_X1 U20885 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17818), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17746) );
  AOI22_X1 U20886 ( .A1(n12119), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17973), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17745) );
  AOI22_X1 U20887 ( .A1(n17975), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17974), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17744) );
  NAND4_X1 U20888 ( .A1(n17747), .A2(n17746), .A3(n17745), .A4(n17744), .ZN(
        n17753) );
  AOI22_X1 U20889 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17954), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17751) );
  AOI22_X1 U20890 ( .A1(n9577), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9581), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17750) );
  AOI22_X1 U20891 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17749) );
  AOI22_X1 U20892 ( .A1(n11960), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17834), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17748) );
  NAND4_X1 U20893 ( .A1(n17751), .A2(n17750), .A3(n17749), .A4(n17748), .ZN(
        n17752) );
  NOR2_X1 U20894 ( .A1(n17753), .A2(n17752), .ZN(n17867) );
  INV_X1 U20895 ( .A(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17940) );
  INV_X1 U20896 ( .A(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17754) );
  OAI22_X1 U20897 ( .A1(n17940), .A2(n17981), .B1(n17844), .B2(n17754), .ZN(
        n17755) );
  INV_X1 U20898 ( .A(n17755), .ZN(n17759) );
  AOI22_X1 U20899 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17818), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17758) );
  AOI22_X1 U20900 ( .A1(n12119), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17973), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17757) );
  AOI22_X1 U20901 ( .A1(n17975), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17974), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17756) );
  NAND4_X1 U20902 ( .A1(n17759), .A2(n17758), .A3(n17757), .A4(n17756), .ZN(
        n17765) );
  AOI22_X1 U20903 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17954), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17763) );
  AOI22_X1 U20904 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9580), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17762) );
  AOI22_X1 U20905 ( .A1(n14172), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17761) );
  AOI22_X1 U20906 ( .A1(n9576), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17834), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17760) );
  NAND4_X1 U20907 ( .A1(n17763), .A2(n17762), .A3(n17761), .A4(n17760), .ZN(
        n17764) );
  OR2_X1 U20908 ( .A1(n17765), .A2(n17764), .ZN(n17882) );
  AOI22_X1 U20909 ( .A1(n17948), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17947), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17771) );
  AOI22_X1 U20910 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17818), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17770) );
  AOI22_X1 U20911 ( .A1(n17903), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17973), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17769) );
  AOI22_X1 U20912 ( .A1(n17975), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17767), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17768) );
  NAND4_X1 U20913 ( .A1(n17771), .A2(n17770), .A3(n17769), .A4(n17768), .ZN(
        n17777) );
  AOI22_X1 U20914 ( .A1(n9578), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9573), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17775) );
  AOI22_X1 U20915 ( .A1(n17954), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9583), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17774) );
  AOI22_X1 U20916 ( .A1(n17953), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17773) );
  AOI22_X1 U20917 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17834), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17772) );
  NAND4_X1 U20918 ( .A1(n17775), .A2(n17774), .A3(n17773), .A4(n17772), .ZN(
        n17776) );
  NOR2_X1 U20919 ( .A1(n17777), .A2(n17776), .ZN(n17887) );
  AOI22_X1 U20920 ( .A1(n17975), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17974), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17781) );
  AOI22_X1 U20921 ( .A1(n12119), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17973), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17780) );
  NAND2_X1 U20922 ( .A1(n17817), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n17779) );
  NAND2_X1 U20923 ( .A1(n17818), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n17778) );
  NAND4_X1 U20924 ( .A1(n17781), .A2(n17780), .A3(n17779), .A4(n17778), .ZN(
        n17784) );
  INV_X1 U20925 ( .A(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17782) );
  OAI22_X1 U20926 ( .A1(n17844), .A2(n17782), .B1(n17981), .B2(n21347), .ZN(
        n17783) );
  OR2_X1 U20927 ( .A1(n17784), .A2(n17783), .ZN(n17790) );
  AOI22_X1 U20928 ( .A1(n9578), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17954), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17788) );
  AOI22_X1 U20929 ( .A1(n9574), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17953), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17787) );
  AOI22_X1 U20930 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17786) );
  AOI22_X1 U20931 ( .A1(n9581), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17834), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17785) );
  NAND4_X1 U20932 ( .A1(n17788), .A2(n17787), .A3(n17786), .A4(n17785), .ZN(
        n17789) );
  NOR2_X1 U20933 ( .A1(n17790), .A2(n17789), .ZN(n17897) );
  AOI22_X1 U20934 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n17975), .B1(
        n17974), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17794) );
  AOI22_X1 U20935 ( .A1(n12119), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17973), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17793) );
  NAND2_X1 U20936 ( .A1(n17818), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n17792) );
  NAND2_X1 U20937 ( .A1(n17817), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n17791) );
  NAND4_X1 U20938 ( .A1(n17794), .A2(n17793), .A3(n17792), .A4(n17791), .ZN(
        n17797) );
  INV_X1 U20939 ( .A(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n21247) );
  OAI22_X1 U20940 ( .A1(n21247), .A2(n17844), .B1(n17981), .B2(n17795), .ZN(
        n17796) );
  OR2_X1 U20941 ( .A1(n17797), .A2(n17796), .ZN(n17803) );
  AOI22_X1 U20942 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n17954), .B1(
        n9580), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17801) );
  AOI22_X1 U20943 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17953), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17800) );
  AOI22_X1 U20944 ( .A1(n9576), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17799) );
  AOI22_X1 U20945 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17834), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17798) );
  NAND4_X1 U20946 ( .A1(n17801), .A2(n17800), .A3(n17799), .A4(n17798), .ZN(
        n17802) );
  NOR2_X1 U20947 ( .A1(n17803), .A2(n17802), .ZN(n17898) );
  NOR2_X1 U20948 ( .A1(n17897), .A2(n17898), .ZN(n17896) );
  INV_X1 U20949 ( .A(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17805) );
  INV_X1 U20950 ( .A(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17804) );
  OAI22_X1 U20951 ( .A1(n17844), .A2(n17805), .B1(n17981), .B2(n17804), .ZN(
        n17806) );
  INV_X1 U20952 ( .A(n17806), .ZN(n17810) );
  AOI22_X1 U20953 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17818), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17809) );
  AOI22_X1 U20954 ( .A1(n12119), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17973), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17808) );
  AOI22_X1 U20955 ( .A1(n17975), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17974), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17807) );
  NAND4_X1 U20956 ( .A1(n17810), .A2(n17809), .A3(n17808), .A4(n17807), .ZN(
        n17816) );
  AOI22_X1 U20957 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17954), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17814) );
  AOI22_X1 U20958 ( .A1(n9572), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9582), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17813) );
  AOI22_X1 U20959 ( .A1(n14172), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17812) );
  AOI22_X1 U20960 ( .A1(n9577), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17834), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17811) );
  NAND4_X1 U20961 ( .A1(n17814), .A2(n17813), .A3(n17812), .A4(n17811), .ZN(
        n17815) );
  OR2_X1 U20962 ( .A1(n17816), .A2(n17815), .ZN(n17892) );
  NAND2_X1 U20963 ( .A1(n17896), .A2(n17892), .ZN(n17891) );
  NOR2_X1 U20964 ( .A1(n17887), .A2(n17891), .ZN(n17886) );
  NAND2_X1 U20965 ( .A1(n17882), .A2(n17886), .ZN(n17881) );
  AOI22_X1 U20966 ( .A1(n17975), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17974), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17822) );
  AOI22_X1 U20967 ( .A1(n12119), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17973), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17821) );
  NAND2_X1 U20968 ( .A1(n17817), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n17820) );
  NAND2_X1 U20969 ( .A1(n17818), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n17819) );
  NAND4_X1 U20970 ( .A1(n17822), .A2(n17821), .A3(n17820), .A4(n17819), .ZN(
        n17826) );
  INV_X1 U20971 ( .A(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17823) );
  OAI22_X1 U20972 ( .A1(n17824), .A2(n17981), .B1(n17844), .B2(n17823), .ZN(
        n17825) );
  OR2_X1 U20973 ( .A1(n17826), .A2(n17825), .ZN(n17832) );
  AOI22_X1 U20974 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17954), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17830) );
  AOI22_X1 U20975 ( .A1(n9572), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9581), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17829) );
  AOI22_X1 U20976 ( .A1(n14172), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17828) );
  AOI22_X1 U20977 ( .A1(n9578), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17834), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17827) );
  NAND4_X1 U20978 ( .A1(n17830), .A2(n17829), .A3(n17828), .A4(n17827), .ZN(
        n17831) );
  NOR2_X1 U20979 ( .A1(n17832), .A2(n17831), .ZN(n17875) );
  NOR2_X1 U20980 ( .A1(n17881), .A2(n17875), .ZN(n17877) );
  AOI22_X1 U20981 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17954), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17838) );
  AOI22_X1 U20982 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9582), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17837) );
  AOI22_X1 U20983 ( .A1(n17953), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17836) );
  AOI22_X1 U20984 ( .A1(n9577), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17834), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17835) );
  NAND4_X1 U20985 ( .A1(n17838), .A2(n17837), .A3(n17836), .A4(n17835), .ZN(
        n17847) );
  AOI22_X1 U20986 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17818), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17841) );
  AOI22_X1 U20987 ( .A1(n12119), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17973), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17840) );
  AOI22_X1 U20988 ( .A1(n17975), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17974), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17839) );
  NAND3_X1 U20989 ( .A1(n17841), .A2(n17840), .A3(n17839), .ZN(n17846) );
  INV_X1 U20990 ( .A(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17843) );
  INV_X1 U20991 ( .A(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17842) );
  OAI22_X1 U20992 ( .A1(n17844), .A2(n17843), .B1(n17981), .B2(n17842), .ZN(
        n17845) );
  OR3_X1 U20993 ( .A1(n17847), .A2(n17846), .A3(n17845), .ZN(n17872) );
  NAND2_X1 U20994 ( .A1(n17877), .A2(n17872), .ZN(n17871) );
  NOR2_X1 U20995 ( .A1(n17867), .A2(n17871), .ZN(n17866) );
  AOI22_X1 U20996 ( .A1(n17966), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17954), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17851) );
  AOI22_X1 U20997 ( .A1(n14172), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17850) );
  AOI22_X1 U20998 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n9574), .B1(
        n9583), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17849) );
  AOI22_X1 U20999 ( .A1(n9576), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17967), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17848) );
  NAND4_X1 U21000 ( .A1(n17851), .A2(n17850), .A3(n17849), .A4(n17848), .ZN(
        n17858) );
  AOI22_X1 U21001 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n17972), .B1(
        n17818), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17854) );
  AOI22_X1 U21002 ( .A1(n17903), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17973), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17853) );
  AOI22_X1 U21003 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n17975), .B1(
        n17974), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17852) );
  NAND3_X1 U21004 ( .A1(n17854), .A2(n17853), .A3(n17852), .ZN(n17857) );
  INV_X1 U21005 ( .A(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17855) );
  OAI22_X1 U21006 ( .A1(n21247), .A2(n17981), .B1(n17844), .B2(n17855), .ZN(
        n17856) );
  OR3_X1 U21007 ( .A1(n17858), .A2(n17857), .A3(n17856), .ZN(n17859) );
  XNOR2_X1 U21008 ( .A(n17866), .B(n17859), .ZN(n18024) );
  OAI22_X1 U21009 ( .A1(n17861), .A2(n17860), .B1(n18024), .B2(n18013), .ZN(
        P3_U2673) );
  NAND2_X1 U21010 ( .A1(n17863), .A2(n17862), .ZN(n17926) );
  NAND2_X1 U21011 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17902), .ZN(n17895) );
  NAND2_X1 U21012 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17901), .ZN(n17885) );
  NAND2_X1 U21013 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n17884), .ZN(n17874) );
  INV_X1 U21014 ( .A(n17874), .ZN(n17880) );
  NAND2_X1 U21015 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17880), .ZN(n17870) );
  AOI21_X1 U21016 ( .B1(n17867), .B2(n17871), .A(n17866), .ZN(n18028) );
  INV_X1 U21017 ( .A(n18028), .ZN(n17869) );
  NAND3_X1 U21018 ( .A1(n17870), .A2(P3_EBX_REG_29__SCAN_IN), .A3(n18013), 
        .ZN(n17868) );
  OAI221_X1 U21019 ( .B1(n17870), .B2(P3_EBX_REG_29__SCAN_IN), .C1(n18013), 
        .C2(n17869), .A(n17868), .ZN(P3_U2674) );
  OAI21_X1 U21020 ( .B1(n17877), .B2(n17872), .A(n17871), .ZN(n18035) );
  NAND3_X1 U21021 ( .A1(n17874), .A2(P3_EBX_REG_28__SCAN_IN), .A3(n18013), 
        .ZN(n17873) );
  OAI221_X1 U21022 ( .B1(n17874), .B2(P3_EBX_REG_28__SCAN_IN), .C1(n18013), 
        .C2(n18035), .A(n17873), .ZN(P3_U2675) );
  AOI21_X1 U21023 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n18013), .A(n17884), .ZN(
        n17879) );
  AND2_X1 U21024 ( .A1(n17881), .A2(n17875), .ZN(n17876) );
  NOR2_X1 U21025 ( .A1(n17877), .A2(n17876), .ZN(n18036) );
  INV_X1 U21026 ( .A(n18036), .ZN(n17878) );
  OAI22_X1 U21027 ( .A1(n17880), .A2(n17879), .B1(n18013), .B2(n17878), .ZN(
        P3_U2676) );
  AOI21_X1 U21028 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n18013), .A(n17890), .ZN(
        n17883) );
  OAI21_X1 U21029 ( .B1(n17886), .B2(n17882), .A(n17881), .ZN(n18044) );
  OAI22_X1 U21030 ( .A1(n17884), .A2(n17883), .B1(n18013), .B2(n18044), .ZN(
        P3_U2677) );
  INV_X1 U21031 ( .A(n17885), .ZN(n17894) );
  AOI21_X1 U21032 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n18013), .A(n17894), .ZN(
        n17889) );
  AOI21_X1 U21033 ( .B1(n17887), .B2(n17891), .A(n17886), .ZN(n18045) );
  INV_X1 U21034 ( .A(n18045), .ZN(n17888) );
  OAI22_X1 U21035 ( .A1(n17890), .A2(n17889), .B1(n18013), .B2(n17888), .ZN(
        P3_U2678) );
  AOI21_X1 U21036 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n18013), .A(n17901), .ZN(
        n17893) );
  OAI21_X1 U21037 ( .B1(n17896), .B2(n17892), .A(n17891), .ZN(n18054) );
  OAI22_X1 U21038 ( .A1(n17894), .A2(n17893), .B1(n18013), .B2(n18054), .ZN(
        P3_U2679) );
  INV_X1 U21039 ( .A(n17895), .ZN(n17915) );
  AOI21_X1 U21040 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n18013), .A(n17915), .ZN(
        n17900) );
  AOI21_X1 U21041 ( .B1(n17898), .B2(n17897), .A(n17896), .ZN(n18055) );
  INV_X1 U21042 ( .A(n18055), .ZN(n17899) );
  OAI22_X1 U21043 ( .A1(n17901), .A2(n17900), .B1(n18013), .B2(n17899), .ZN(
        P3_U2680) );
  AOI21_X1 U21044 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n18013), .A(n17902), .ZN(
        n17914) );
  AOI22_X1 U21045 ( .A1(n17948), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17947), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17907) );
  AOI22_X1 U21046 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17818), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17906) );
  AOI22_X1 U21047 ( .A1(n12119), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17973), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17905) );
  AOI22_X1 U21048 ( .A1(n17975), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17974), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17904) );
  NAND4_X1 U21049 ( .A1(n17907), .A2(n17906), .A3(n17905), .A4(n17904), .ZN(
        n17913) );
  AOI22_X1 U21050 ( .A1(n17966), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17954), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17911) );
  AOI22_X1 U21051 ( .A1(n9577), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9573), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17910) );
  AOI22_X1 U21052 ( .A1(n9583), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17953), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17909) );
  AOI22_X1 U21053 ( .A1(n17932), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17967), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17908) );
  NAND4_X1 U21054 ( .A1(n17911), .A2(n17910), .A3(n17909), .A4(n17908), .ZN(
        n17912) );
  NOR2_X1 U21055 ( .A1(n17913), .A2(n17912), .ZN(n18062) );
  OAI22_X1 U21056 ( .A1(n17915), .A2(n17914), .B1(n18062), .B2(n18013), .ZN(
        P3_U2681) );
  AOI22_X1 U21057 ( .A1(n17948), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17947), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17919) );
  AOI22_X1 U21058 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17818), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17918) );
  AOI22_X1 U21059 ( .A1(n12119), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17973), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17917) );
  AOI22_X1 U21060 ( .A1(n17975), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17974), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17916) );
  NAND4_X1 U21061 ( .A1(n17919), .A2(n17918), .A3(n17917), .A4(n17916), .ZN(
        n17925) );
  AOI22_X1 U21062 ( .A1(n9576), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9574), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17923) );
  AOI22_X1 U21063 ( .A1(n17954), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9582), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17922) );
  AOI22_X1 U21064 ( .A1(n17966), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11944), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17921) );
  AOI22_X1 U21065 ( .A1(n11960), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17967), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17920) );
  NAND4_X1 U21066 ( .A1(n17923), .A2(n17922), .A3(n17921), .A4(n17920), .ZN(
        n17924) );
  NOR2_X1 U21067 ( .A1(n17925), .A2(n17924), .ZN(n18070) );
  INV_X1 U21068 ( .A(n17926), .ZN(n17928) );
  AOI22_X1 U21069 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17929), .B1(n17928), 
        .B2(n17927), .ZN(n17930) );
  OAI21_X1 U21070 ( .B1(n18070), .B2(n18013), .A(n17930), .ZN(P3_U2682) );
  INV_X1 U21071 ( .A(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n21279) );
  OAI22_X1 U21072 ( .A1(n18002), .A2(n12101), .B1(n17931), .B2(n21279), .ZN(
        n17944) );
  AOI22_X1 U21073 ( .A1(n17966), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9574), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17936) );
  AOI22_X1 U21074 ( .A1(n17954), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9580), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17935) );
  AOI22_X1 U21075 ( .A1(n9576), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17953), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17934) );
  AOI22_X1 U21076 ( .A1(n17932), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17967), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17933) );
  NAND4_X1 U21077 ( .A1(n17936), .A2(n17935), .A3(n17934), .A4(n17933), .ZN(
        n17943) );
  AOI22_X1 U21078 ( .A1(n17975), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17974), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17938) );
  AOI22_X1 U21079 ( .A1(n12119), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17973), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17937) );
  NAND2_X1 U21080 ( .A1(n17938), .A2(n17937), .ZN(n17942) );
  OAI22_X1 U21081 ( .A1(n17940), .A2(n9568), .B1(n17981), .B2(n17939), .ZN(
        n17941) );
  NOR4_X1 U21082 ( .A1(n17944), .A2(n17943), .A3(n17942), .A4(n17941), .ZN(
        n18074) );
  OAI221_X1 U21083 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(P3_EBX_REG_18__SCAN_IN), 
        .C1(P3_EBX_REG_19__SCAN_IN), .C2(n17962), .A(n17945), .ZN(n17946) );
  AOI22_X1 U21084 ( .A1(n18016), .A2(n18074), .B1(n17946), .B2(n18013), .ZN(
        P3_U2684) );
  AOI22_X1 U21085 ( .A1(n17948), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17947), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17952) );
  AOI22_X1 U21086 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17818), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17951) );
  AOI22_X1 U21087 ( .A1(n17975), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17973), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17950) );
  AOI22_X1 U21088 ( .A1(n17974), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12119), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17949) );
  NAND4_X1 U21089 ( .A1(n17952), .A2(n17951), .A3(n17950), .A4(n17949), .ZN(
        n17960) );
  AOI22_X1 U21090 ( .A1(n17966), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9572), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17958) );
  AOI22_X1 U21091 ( .A1(n9577), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17953), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17957) );
  AOI22_X1 U21092 ( .A1(n9583), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11944), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17956) );
  AOI22_X1 U21093 ( .A1(n17954), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17967), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17955) );
  NAND4_X1 U21094 ( .A1(n17958), .A2(n17957), .A3(n17956), .A4(n17955), .ZN(
        n17959) );
  NOR2_X1 U21095 ( .A1(n17960), .A2(n17959), .ZN(n18082) );
  AOI22_X1 U21096 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17963), .B1(n17962), 
        .B2(n17961), .ZN(n17964) );
  OAI21_X1 U21097 ( .B1(n18082), .B2(n18013), .A(n17964), .ZN(P3_U2685) );
  NAND2_X1 U21098 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17965), .ZN(n17988) );
  AOI22_X1 U21099 ( .A1(n17966), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17954), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17971) );
  AOI22_X1 U21100 ( .A1(n9572), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9581), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17970) );
  AOI22_X1 U21101 ( .A1(n11960), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17932), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17969) );
  AOI22_X1 U21102 ( .A1(n9576), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17967), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17968) );
  NAND4_X1 U21103 ( .A1(n17971), .A2(n17970), .A3(n17969), .A4(n17968), .ZN(
        n17985) );
  AOI22_X1 U21104 ( .A1(n17972), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17818), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17978) );
  AOI22_X1 U21105 ( .A1(n12119), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17973), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17977) );
  AOI22_X1 U21106 ( .A1(n17975), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17974), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17976) );
  NAND3_X1 U21107 ( .A1(n17978), .A2(n17977), .A3(n17976), .ZN(n17984) );
  INV_X1 U21108 ( .A(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17979) );
  OAI22_X1 U21109 ( .A1(n17982), .A2(n17981), .B1(n9568), .B2(n17979), .ZN(
        n17983) );
  OR3_X1 U21110 ( .A1(n17985), .A2(n17984), .A3(n17983), .ZN(n18089) );
  AOI22_X1 U21111 ( .A1(n17986), .A2(P3_EBX_REG_14__SCAN_IN), .B1(n18016), 
        .B2(n18089), .ZN(n17987) );
  OAI21_X1 U21112 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17988), .A(n17987), .ZN(
        P3_U2689) );
  OAI21_X1 U21113 ( .B1(n17992), .B2(n17995), .A(n18013), .ZN(n17993) );
  AOI22_X1 U21114 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18016), .B1(
        n17989), .B2(n17991), .ZN(n17990) );
  OAI21_X1 U21115 ( .B1(n17991), .B2(n17993), .A(n17990), .ZN(P3_U2697) );
  AND2_X1 U21116 ( .A1(n17992), .A2(n17995), .ZN(n17994) );
  OAI22_X1 U21117 ( .A1(n17994), .A2(n17993), .B1(n11954), .B2(n18013), .ZN(
        P3_U2698) );
  INV_X1 U21118 ( .A(n17995), .ZN(n17999) );
  NAND2_X1 U21119 ( .A1(n17996), .A2(n18011), .ZN(n18005) );
  NOR2_X1 U21120 ( .A1(n18000), .A2(n18005), .ZN(n18004) );
  AOI21_X1 U21121 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n18013), .A(n18004), .ZN(
        n17998) );
  OAI22_X1 U21122 ( .A1(n17999), .A2(n17998), .B1(n17997), .B2(n18013), .ZN(
        P3_U2699) );
  OAI21_X1 U21123 ( .B1(n18000), .B2(n18016), .A(n18005), .ZN(n18001) );
  INV_X1 U21124 ( .A(n18001), .ZN(n18003) );
  OAI22_X1 U21125 ( .A1(n18004), .A2(n18003), .B1(n18002), .B2(n18013), .ZN(
        P3_U2700) );
  OAI221_X1 U21126 ( .B1(P3_EBX_REG_2__SCAN_IN), .B2(n18007), .C1(
        P3_EBX_REG_2__SCAN_IN), .C2(n18006), .A(n18005), .ZN(n18008) );
  AOI22_X1 U21127 ( .A1(n18016), .A2(n18009), .B1(n18008), .B2(n18013), .ZN(
        P3_U2701) );
  AOI22_X1 U21128 ( .A1(P3_EBX_REG_1__SCAN_IN), .A2(n18015), .B1(n18011), .B2(
        n18010), .ZN(n18012) );
  OAI21_X1 U21129 ( .B1(n18014), .B2(n18013), .A(n18012), .ZN(P3_U2702) );
  AOI22_X1 U21130 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18016), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n18015), .ZN(n18017) );
  OAI21_X1 U21131 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n18018), .A(n18017), .ZN(
        P3_U2703) );
  INV_X1 U21132 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n18201) );
  INV_X1 U21133 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n18197) );
  INV_X1 U21134 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n18192) );
  INV_X1 U21135 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n18190) );
  INV_X1 U21136 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n18207) );
  OR2_X1 U21137 ( .A1(n9661), .A2(n18207), .ZN(n18023) );
  NAND2_X1 U21138 ( .A1(n18120), .A2(n9661), .ZN(n18027) );
  OAI21_X1 U21139 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n18020), .A(n18027), .ZN(
        n18021) );
  AOI22_X1 U21140 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n18075), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n18021), .ZN(n18022) );
  OAI21_X1 U21141 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n18023), .A(n18022), .ZN(
        P3_U2704) );
  OAI22_X1 U21142 ( .A1(n18024), .A2(n18123), .B1(n16076), .B2(n18061), .ZN(
        n18025) );
  AOI21_X1 U21143 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n18076), .A(n18025), .ZN(
        n18026) );
  OAI221_X1 U21144 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n9661), .C1(n18207), 
        .C2(n18027), .A(n18026), .ZN(P3_U2705) );
  AOI22_X1 U21145 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18076), .B1(n18104), .B2(
        n18028), .ZN(n18031) );
  OAI211_X1 U21146 ( .C1(n18029), .C2(P3_EAX_REG_29__SCAN_IN), .A(n18120), .B(
        n9661), .ZN(n18030) );
  OAI211_X1 U21147 ( .C1(n18061), .C2(n16082), .A(n18031), .B(n18030), .ZN(
        P3_U2706) );
  AOI22_X1 U21148 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n18076), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n18075), .ZN(n18034) );
  OAI211_X1 U21149 ( .C1(n18037), .C2(P3_EAX_REG_28__SCAN_IN), .A(n18120), .B(
        n18032), .ZN(n18033) );
  OAI211_X1 U21150 ( .C1(n18035), .C2(n18123), .A(n18034), .B(n18033), .ZN(
        P3_U2707) );
  AOI22_X1 U21151 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18076), .B1(n18104), .B2(
        n18036), .ZN(n18040) );
  AOI211_X1 U21152 ( .C1(n18201), .C2(n18041), .A(n18037), .B(n18102), .ZN(
        n18038) );
  INV_X1 U21153 ( .A(n18038), .ZN(n18039) );
  OAI211_X1 U21154 ( .C1(n18061), .C2(n16102), .A(n18040), .B(n18039), .ZN(
        P3_U2708) );
  AOI22_X1 U21155 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18076), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n18075), .ZN(n18043) );
  OAI211_X1 U21156 ( .C1(n18046), .C2(P3_EAX_REG_26__SCAN_IN), .A(n18120), .B(
        n18041), .ZN(n18042) );
  OAI211_X1 U21157 ( .C1(n18044), .C2(n18123), .A(n18043), .B(n18042), .ZN(
        P3_U2709) );
  AOI22_X1 U21158 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18075), .B1(n18104), .B2(
        n18045), .ZN(n18049) );
  AOI211_X1 U21159 ( .C1(n18197), .C2(n18050), .A(n18046), .B(n18102), .ZN(
        n18047) );
  INV_X1 U21160 ( .A(n18047), .ZN(n18048) );
  OAI211_X1 U21161 ( .C1(n18060), .C2(n21365), .A(n18049), .B(n18048), .ZN(
        P3_U2710) );
  AOI22_X1 U21162 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18076), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n18075), .ZN(n18053) );
  OAI211_X1 U21163 ( .C1(n18051), .C2(P3_EAX_REG_24__SCAN_IN), .A(n18120), .B(
        n18050), .ZN(n18052) );
  OAI211_X1 U21164 ( .C1(n18054), .C2(n18123), .A(n18053), .B(n18052), .ZN(
        P3_U2711) );
  AOI22_X1 U21165 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18075), .B1(n18104), .B2(
        n18055), .ZN(n18059) );
  OAI211_X1 U21166 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n18057), .A(n18056), .B(
        n18120), .ZN(n18058) );
  OAI211_X1 U21167 ( .C1(n18060), .C2(n18785), .A(n18059), .B(n18058), .ZN(
        P3_U2712) );
  NAND2_X1 U21168 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n18067), .ZN(n18066) );
  NAND3_X1 U21169 ( .A1(n18120), .A2(P3_EAX_REG_22__SCAN_IN), .A3(n18066), 
        .ZN(n18065) );
  OAI22_X1 U21170 ( .A1(n18062), .A2(n18123), .B1(n16142), .B2(n18061), .ZN(
        n18063) );
  AOI21_X1 U21171 ( .B1(BUF2_REG_6__SCAN_IN), .B2(n18076), .A(n18063), .ZN(
        n18064) );
  OAI211_X1 U21172 ( .C1(P3_EAX_REG_22__SCAN_IN), .C2(n18066), .A(n18065), .B(
        n18064), .ZN(P3_U2713) );
  AOI22_X1 U21173 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n18076), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n18075), .ZN(n18069) );
  OAI211_X1 U21174 ( .C1(n18067), .C2(P3_EAX_REG_21__SCAN_IN), .A(n18120), .B(
        n18066), .ZN(n18068) );
  OAI211_X1 U21175 ( .C1(n18070), .C2(n18123), .A(n18069), .B(n18068), .ZN(
        P3_U2714) );
  AOI22_X1 U21176 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18076), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n18075), .ZN(n18073) );
  OAI211_X1 U21177 ( .C1(n18077), .C2(P3_EAX_REG_19__SCAN_IN), .A(n18120), .B(
        n18071), .ZN(n18072) );
  OAI211_X1 U21178 ( .C1(n18074), .C2(n18123), .A(n18073), .B(n18072), .ZN(
        P3_U2716) );
  AOI22_X1 U21179 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n18076), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n18075), .ZN(n18081) );
  AOI211_X1 U21180 ( .C1(n18184), .C2(n18078), .A(n18077), .B(n18102), .ZN(
        n18079) );
  INV_X1 U21181 ( .A(n18079), .ZN(n18080) );
  OAI211_X1 U21182 ( .C1(n18082), .C2(n18123), .A(n18081), .B(n18080), .ZN(
        P3_U2717) );
  NAND2_X1 U21183 ( .A1(n18084), .A2(n18083), .ZN(n18088) );
  NAND2_X1 U21184 ( .A1(n18120), .A2(n18085), .ZN(n18091) );
  INV_X1 U21185 ( .A(n18126), .ZN(n18105) );
  AOI22_X1 U21186 ( .A1(n18105), .A2(BUF2_REG_15__SCAN_IN), .B1(n18104), .B2(
        n18086), .ZN(n18087) );
  OAI221_X1 U21187 ( .B1(P3_EAX_REG_15__SCAN_IN), .B2(n18088), .C1(n18238), 
        .C2(n18091), .A(n18087), .ZN(P3_U2720) );
  AOI22_X1 U21188 ( .A1(n18105), .A2(BUF2_REG_14__SCAN_IN), .B1(n18104), .B2(
        n18089), .ZN(n18090) );
  OAI221_X1 U21189 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n18092), .C1(n18233), 
        .C2(n18091), .A(n18090), .ZN(P3_U2721) );
  NAND2_X1 U21190 ( .A1(n18120), .A2(n18096), .ZN(n18100) );
  OAI22_X1 U21191 ( .A1(n18126), .A2(n18225), .B1(n18093), .B2(n18123), .ZN(
        n18094) );
  INV_X1 U21192 ( .A(n18094), .ZN(n18095) );
  OAI221_X1 U21193 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n18096), .C1(n18151), 
        .C2(n18100), .A(n18095), .ZN(P3_U2724) );
  INV_X1 U21194 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n18223) );
  AOI22_X1 U21195 ( .A1(n18105), .A2(BUF2_REG_10__SCAN_IN), .B1(n18104), .B2(
        n18097), .ZN(n18098) );
  OAI221_X1 U21196 ( .B1(n18100), .B2(n18223), .C1(n18100), .C2(n18099), .A(
        n18098), .ZN(P3_U2725) );
  OR2_X1 U21197 ( .A1(n18102), .A2(n18101), .ZN(n18107) );
  AOI22_X1 U21198 ( .A1(n18105), .A2(BUF2_REG_8__SCAN_IN), .B1(n18104), .B2(
        n18103), .ZN(n18106) );
  OAI221_X1 U21199 ( .B1(P3_EAX_REG_8__SCAN_IN), .B2(n18108), .C1(n18220), 
        .C2(n18107), .A(n18106), .ZN(P3_U2727) );
  INV_X1 U21200 ( .A(n18109), .ZN(n18115) );
  AOI21_X1 U21201 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n18120), .A(n18115), .ZN(
        n18111) );
  OAI222_X1 U21202 ( .A1(n18780), .A2(n18126), .B1(n18112), .B2(n18111), .C1(
        n18123), .C2(n18110), .ZN(P3_U2729) );
  AOI21_X1 U21203 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n18120), .A(n18119), .ZN(
        n18114) );
  OAI222_X1 U21204 ( .A1(n18776), .A2(n18126), .B1(n18115), .B2(n18114), .C1(
        n18123), .C2(n18113), .ZN(P3_U2730) );
  INV_X1 U21205 ( .A(n18116), .ZN(n18125) );
  AOI21_X1 U21206 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n18120), .A(n18125), .ZN(
        n18118) );
  OAI222_X1 U21207 ( .A1(n18772), .A2(n18126), .B1(n18119), .B2(n18118), .C1(
        n18123), .C2(n18117), .ZN(P3_U2731) );
  AOI22_X1 U21208 ( .A1(n18121), .A2(P3_EAX_REG_2__SCAN_IN), .B1(
        P3_EAX_REG_3__SCAN_IN), .B2(n18120), .ZN(n18124) );
  OAI222_X1 U21209 ( .A1(n18767), .A2(n18126), .B1(n18125), .B2(n18124), .C1(
        n18123), .C2(n18122), .ZN(P3_U2732) );
  INV_X1 U21210 ( .A(n18313), .ZN(n18370) );
  NAND2_X1 U21211 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18370), .ZN(n19342) );
  NOR2_X1 U21212 ( .A1(n18166), .A2(n18128), .ZN(P3_U2736) );
  NAND2_X1 U21213 ( .A1(n18164), .A2(n18755), .ZN(n18144) );
  INV_X2 U21214 ( .A(n19342), .ZN(n18170) );
  AOI22_X1 U21215 ( .A1(n18170), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n18169), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18129) );
  OAI21_X1 U21216 ( .B1(n18207), .B2(n18144), .A(n18129), .ZN(P3_U2737) );
  INV_X1 U21217 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n18205) );
  AOI22_X1 U21218 ( .A1(n18170), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18169), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18130) );
  OAI21_X1 U21219 ( .B1(n18205), .B2(n18144), .A(n18130), .ZN(P3_U2738) );
  INV_X1 U21220 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n18203) );
  AOI22_X1 U21221 ( .A1(n18170), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18169), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18131) );
  OAI21_X1 U21222 ( .B1(n18203), .B2(n18144), .A(n18131), .ZN(P3_U2739) );
  AOI22_X1 U21223 ( .A1(P3_DATAO_REG_27__SCAN_IN), .A2(n18169), .B1(n18170), 
        .B2(P3_UWORD_REG_11__SCAN_IN), .ZN(n18132) );
  OAI21_X1 U21224 ( .B1(n18201), .B2(n18144), .A(n18132), .ZN(P3_U2740) );
  INV_X1 U21225 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n18199) );
  AOI22_X1 U21226 ( .A1(n18170), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n18169), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18133) );
  OAI21_X1 U21227 ( .B1(n18199), .B2(n18144), .A(n18133), .ZN(P3_U2741) );
  AOI22_X1 U21228 ( .A1(n18170), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18169), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18134) );
  OAI21_X1 U21229 ( .B1(n18197), .B2(n18144), .A(n18134), .ZN(P3_U2742) );
  INV_X1 U21230 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n18195) );
  AOI22_X1 U21231 ( .A1(n18170), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n18169), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18135) );
  OAI21_X1 U21232 ( .B1(n18195), .B2(n18144), .A(n18135), .ZN(P3_U2743) );
  INV_X1 U21233 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n21299) );
  AOI22_X1 U21234 ( .A1(n18170), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n18169), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18136) );
  OAI21_X1 U21235 ( .B1(n21299), .B2(n18144), .A(n18136), .ZN(P3_U2744) );
  AOI22_X1 U21236 ( .A1(n18170), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18169), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18137) );
  OAI21_X1 U21237 ( .B1(n18192), .B2(n18144), .A(n18137), .ZN(P3_U2745) );
  AOI22_X1 U21238 ( .A1(n18170), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n18169), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18138) );
  OAI21_X1 U21239 ( .B1(n18190), .B2(n18144), .A(n18138), .ZN(P3_U2746) );
  AOI22_X1 U21240 ( .A1(n18170), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18169), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18139) );
  OAI21_X1 U21241 ( .B1(n18188), .B2(n18144), .A(n18139), .ZN(P3_U2747) );
  INV_X1 U21242 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n18186) );
  AOI22_X1 U21243 ( .A1(n18170), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n18169), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18140) );
  OAI21_X1 U21244 ( .B1(n18186), .B2(n18144), .A(n18140), .ZN(P3_U2748) );
  AOI22_X1 U21245 ( .A1(n18170), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n18169), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18141) );
  OAI21_X1 U21246 ( .B1(n18184), .B2(n18144), .A(n18141), .ZN(P3_U2749) );
  INV_X1 U21247 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n18182) );
  AOI22_X1 U21248 ( .A1(n18170), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n18169), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18142) );
  OAI21_X1 U21249 ( .B1(n18182), .B2(n18144), .A(n18142), .ZN(P3_U2750) );
  INV_X1 U21250 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n18180) );
  AOI22_X1 U21251 ( .A1(n18170), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n18169), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18143) );
  OAI21_X1 U21252 ( .B1(n18180), .B2(n18144), .A(n18143), .ZN(P3_U2751) );
  INV_X1 U21253 ( .A(P3_DATAO_REG_15__SCAN_IN), .ZN(n21314) );
  AOI22_X1 U21254 ( .A1(P3_EAX_REG_15__SCAN_IN), .A2(n18164), .B1(n18170), 
        .B2(P3_LWORD_REG_15__SCAN_IN), .ZN(n18145) );
  OAI21_X1 U21255 ( .B1(n21314), .B2(n18166), .A(n18145), .ZN(P3_U2752) );
  AOI22_X1 U21256 ( .A1(n18170), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n18169), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18146) );
  OAI21_X1 U21257 ( .B1(n18233), .B2(n18172), .A(n18146), .ZN(P3_U2753) );
  INV_X1 U21258 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n18148) );
  AOI22_X1 U21259 ( .A1(n18170), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n18169), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18147) );
  OAI21_X1 U21260 ( .B1(n18148), .B2(n18172), .A(n18147), .ZN(P3_U2754) );
  AOI22_X1 U21261 ( .A1(n18170), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n18169), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18149) );
  OAI21_X1 U21262 ( .B1(n21285), .B2(n18172), .A(n18149), .ZN(P3_U2755) );
  AOI22_X1 U21263 ( .A1(n18170), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18169), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18150) );
  OAI21_X1 U21264 ( .B1(n18151), .B2(n18172), .A(n18150), .ZN(P3_U2756) );
  AOI22_X1 U21265 ( .A1(n18170), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18169), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18152) );
  OAI21_X1 U21266 ( .B1(n18223), .B2(n18172), .A(n18152), .ZN(P3_U2757) );
  INV_X1 U21267 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n18154) );
  AOI22_X1 U21268 ( .A1(n18170), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n18169), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18153) );
  OAI21_X1 U21269 ( .B1(n18154), .B2(n18172), .A(n18153), .ZN(P3_U2758) );
  AOI22_X1 U21270 ( .A1(n18170), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18169), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18155) );
  OAI21_X1 U21271 ( .B1(n18220), .B2(n18172), .A(n18155), .ZN(P3_U2759) );
  INV_X1 U21272 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n18157) );
  AOI22_X1 U21273 ( .A1(n18170), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n18169), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18156) );
  OAI21_X1 U21274 ( .B1(n18157), .B2(n18172), .A(n18156), .ZN(P3_U2760) );
  AOI22_X1 U21275 ( .A1(n18170), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n18169), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18158) );
  OAI21_X1 U21276 ( .B1(n18159), .B2(n18172), .A(n18158), .ZN(P3_U2761) );
  INV_X1 U21277 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n18161) );
  AOI22_X1 U21278 ( .A1(n18170), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18169), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18160) );
  OAI21_X1 U21279 ( .B1(n18161), .B2(n18172), .A(n18160), .ZN(P3_U2762) );
  AOI22_X1 U21280 ( .A1(n18170), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18169), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18162) );
  OAI21_X1 U21281 ( .B1(n18163), .B2(n18172), .A(n18162), .ZN(P3_U2763) );
  INV_X1 U21282 ( .A(P3_DATAO_REG_3__SCAN_IN), .ZN(n21328) );
  AOI22_X1 U21283 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n18164), .B1(n18170), .B2(
        P3_LWORD_REG_3__SCAN_IN), .ZN(n18165) );
  OAI21_X1 U21284 ( .B1(n21328), .B2(n18166), .A(n18165), .ZN(P3_U2764) );
  INV_X1 U21285 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n18213) );
  AOI22_X1 U21286 ( .A1(n18170), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n18169), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18167) );
  OAI21_X1 U21287 ( .B1(n18213), .B2(n18172), .A(n18167), .ZN(P3_U2765) );
  AOI22_X1 U21288 ( .A1(n18170), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n18169), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18168) );
  OAI21_X1 U21289 ( .B1(n18211), .B2(n18172), .A(n18168), .ZN(P3_U2766) );
  AOI22_X1 U21290 ( .A1(n18170), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n18169), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18171) );
  OAI21_X1 U21291 ( .B1(n18209), .B2(n18172), .A(n18171), .ZN(P3_U2767) );
  OR2_X1 U21292 ( .A1(n18175), .A2(n19335), .ZN(n19212) );
  INV_X1 U21293 ( .A(n18173), .ZN(n18177) );
  INV_X1 U21294 ( .A(n19222), .ZN(n19343) );
  AND2_X1 U21295 ( .A1(n19335), .A2(n19343), .ZN(n18174) );
  NOR2_X1 U21296 ( .A1(n18175), .A2(n18174), .ZN(n18176) );
  AOI22_X1 U21297 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n18235), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n18234), .ZN(n18179) );
  OAI21_X1 U21298 ( .B1(n18180), .B2(n18237), .A(n18179), .ZN(P3_U2768) );
  AOI22_X1 U21299 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18235), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n18234), .ZN(n18181) );
  OAI21_X1 U21300 ( .B1(n18182), .B2(n18237), .A(n18181), .ZN(P3_U2769) );
  AOI22_X1 U21301 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n18235), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n18234), .ZN(n18183) );
  OAI21_X1 U21302 ( .B1(n18184), .B2(n18237), .A(n18183), .ZN(P3_U2770) );
  AOI22_X1 U21303 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18235), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n18234), .ZN(n18185) );
  OAI21_X1 U21304 ( .B1(n18186), .B2(n18237), .A(n18185), .ZN(P3_U2771) );
  AOI22_X1 U21305 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n18235), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n18234), .ZN(n18187) );
  OAI21_X1 U21306 ( .B1(n18188), .B2(n18237), .A(n18187), .ZN(P3_U2772) );
  AOI22_X1 U21307 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n18235), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n18234), .ZN(n18189) );
  OAI21_X1 U21308 ( .B1(n18190), .B2(n18237), .A(n18189), .ZN(P3_U2773) );
  AOI22_X1 U21309 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n18235), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n18234), .ZN(n18191) );
  OAI21_X1 U21310 ( .B1(n18192), .B2(n18237), .A(n18191), .ZN(P3_U2774) );
  AOI22_X1 U21311 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18235), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n18234), .ZN(n18193) );
  OAI21_X1 U21312 ( .B1(n21299), .B2(n18237), .A(n18193), .ZN(P3_U2775) );
  AOI22_X1 U21313 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18235), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n18234), .ZN(n18194) );
  OAI21_X1 U21314 ( .B1(n18195), .B2(n18237), .A(n18194), .ZN(P3_U2776) );
  AOI22_X1 U21315 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18235), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n18234), .ZN(n18196) );
  OAI21_X1 U21316 ( .B1(n18197), .B2(n18237), .A(n18196), .ZN(P3_U2777) );
  AOI22_X1 U21317 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18235), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n18234), .ZN(n18198) );
  OAI21_X1 U21318 ( .B1(n18199), .B2(n18237), .A(n18198), .ZN(P3_U2778) );
  AOI22_X1 U21319 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18235), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n18234), .ZN(n18200) );
  OAI21_X1 U21320 ( .B1(n18201), .B2(n18237), .A(n18200), .ZN(P3_U2779) );
  AOI22_X1 U21321 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n18235), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n18234), .ZN(n18202) );
  OAI21_X1 U21322 ( .B1(n18203), .B2(n18237), .A(n18202), .ZN(P3_U2780) );
  AOI22_X1 U21323 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18235), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n18234), .ZN(n18204) );
  OAI21_X1 U21324 ( .B1(n18205), .B2(n18237), .A(n18204), .ZN(P3_U2781) );
  AOI22_X1 U21325 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18235), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n18234), .ZN(n18206) );
  OAI21_X1 U21326 ( .B1(n18207), .B2(n18237), .A(n18206), .ZN(P3_U2782) );
  AOI22_X1 U21327 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n18235), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n18234), .ZN(n18208) );
  OAI21_X1 U21328 ( .B1(n18209), .B2(n18237), .A(n18208), .ZN(P3_U2783) );
  AOI22_X1 U21329 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18235), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n18234), .ZN(n18210) );
  OAI21_X1 U21330 ( .B1(n18211), .B2(n18237), .A(n18210), .ZN(P3_U2784) );
  AOI22_X1 U21331 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n18235), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n18234), .ZN(n18212) );
  OAI21_X1 U21332 ( .B1(n18213), .B2(n18237), .A(n18212), .ZN(P3_U2785) );
  AOI22_X1 U21333 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n18228), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n18234), .ZN(n18214) );
  OAI21_X1 U21334 ( .B1(n18767), .B2(n18230), .A(n18214), .ZN(P3_U2786) );
  AOI22_X1 U21335 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n18228), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n18234), .ZN(n18215) );
  OAI21_X1 U21336 ( .B1(n18772), .B2(n18230), .A(n18215), .ZN(P3_U2787) );
  AOI22_X1 U21337 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n18228), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n18234), .ZN(n18216) );
  OAI21_X1 U21338 ( .B1(n18776), .B2(n18230), .A(n18216), .ZN(P3_U2788) );
  AOI22_X1 U21339 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n18228), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n18234), .ZN(n18217) );
  OAI21_X1 U21340 ( .B1(n18780), .B2(n18230), .A(n18217), .ZN(P3_U2789) );
  AOI22_X1 U21341 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n18228), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n18234), .ZN(n18218) );
  OAI21_X1 U21342 ( .B1(n18785), .B2(n18230), .A(n18218), .ZN(P3_U2790) );
  AOI22_X1 U21343 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18235), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n18234), .ZN(n18219) );
  OAI21_X1 U21344 ( .B1(n18220), .B2(n18237), .A(n18219), .ZN(P3_U2791) );
  AOI22_X1 U21345 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n18228), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n18234), .ZN(n18221) );
  OAI21_X1 U21346 ( .B1(n21365), .B2(n18230), .A(n18221), .ZN(P3_U2792) );
  AOI22_X1 U21347 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18235), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n18234), .ZN(n18222) );
  OAI21_X1 U21348 ( .B1(n18223), .B2(n18237), .A(n18222), .ZN(P3_U2793) );
  AOI22_X1 U21349 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n18228), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n18234), .ZN(n18224) );
  OAI21_X1 U21350 ( .B1(n18225), .B2(n18230), .A(n18224), .ZN(P3_U2794) );
  AOI22_X1 U21351 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n18228), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n18234), .ZN(n18226) );
  OAI21_X1 U21352 ( .B1(n18227), .B2(n18230), .A(n18226), .ZN(P3_U2795) );
  AOI22_X1 U21353 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n18228), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n18234), .ZN(n18229) );
  OAI21_X1 U21354 ( .B1(n18231), .B2(n18230), .A(n18229), .ZN(P3_U2796) );
  AOI22_X1 U21355 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18235), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n18234), .ZN(n18232) );
  OAI21_X1 U21356 ( .B1(n18233), .B2(n18237), .A(n18232), .ZN(P3_U2797) );
  AOI22_X1 U21357 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n18235), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n18234), .ZN(n18236) );
  OAI21_X1 U21358 ( .B1(n18238), .B2(n18237), .A(n18236), .ZN(P3_U2798) );
  AOI21_X1 U21359 ( .B1(n18239), .B2(n16992), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n18247) );
  AOI22_X1 U21360 ( .A1(n18693), .A2(P3_REIP_REG_26__SCAN_IN), .B1(n18240), 
        .B2(n18426), .ZN(n18246) );
  OAI22_X1 U21361 ( .A1(n18242), .A2(n18451), .B1(n18241), .B2(n12028), .ZN(
        n18243) );
  AOI21_X1 U21362 ( .B1(n18320), .B2(n18244), .A(n18243), .ZN(n18245) );
  OAI211_X1 U21363 ( .C1(n18248), .C2(n18247), .A(n18246), .B(n18245), .ZN(
        P3_U2804) );
  NAND2_X1 U21364 ( .A1(n18249), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n18250) );
  XOR2_X1 U21365 ( .A(n18250), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n18513) );
  OAI211_X1 U21366 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n18252), .B(n18251), .ZN(n18253) );
  NAND2_X1 U21367 ( .A1(n18693), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n18508) );
  OAI211_X1 U21368 ( .C1(n18377), .C2(n18254), .A(n18253), .B(n18508), .ZN(
        n18265) );
  NAND2_X1 U21369 ( .A1(n18255), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n18256) );
  XOR2_X1 U21370 ( .A(n18256), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n18497) );
  XNOR2_X1 U21371 ( .A(n18257), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n18260) );
  NOR2_X1 U21372 ( .A1(n18258), .A2(n18509), .ZN(n18259) );
  MUX2_X1 U21373 ( .A(n18260), .B(n18259), .S(n18365), .Z(n18261) );
  INV_X1 U21374 ( .A(n18261), .ZN(n18262) );
  OAI21_X1 U21375 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n18263), .A(
        n18262), .ZN(n18498) );
  OAI22_X1 U21376 ( .A1(n18381), .A2(n18497), .B1(n18451), .B2(n18498), .ZN(
        n18264) );
  AOI211_X1 U21377 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n18266), .A(
        n18265), .B(n18264), .ZN(n18267) );
  OAI21_X1 U21378 ( .B1(n18380), .B2(n18513), .A(n18267), .ZN(P3_U2805) );
  INV_X1 U21379 ( .A(n18522), .ZN(n18530) );
  NOR2_X1 U21380 ( .A1(n18343), .A2(n18530), .ZN(n18268) );
  OAI21_X1 U21381 ( .B1(n18269), .B2(n18268), .A(n18298), .ZN(n18270) );
  INV_X1 U21382 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18531) );
  XNOR2_X1 U21383 ( .A(n18270), .B(n18531), .ZN(n18536) );
  INV_X1 U21384 ( .A(n18271), .ZN(n18307) );
  OAI21_X1 U21385 ( .B1(n18307), .B2(n18522), .A(n18329), .ZN(n18294) );
  OAI21_X1 U21386 ( .B1(n18273), .B2(n18313), .A(n18495), .ZN(n18274) );
  AOI21_X1 U21387 ( .B1(n18368), .B2(n13596), .A(n18274), .ZN(n18302) );
  OAI21_X1 U21388 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18275), .A(
        n18302), .ZN(n18290) );
  AOI22_X1 U21389 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n18290), .B1(
        n18391), .B2(n18276), .ZN(n18279) );
  NOR2_X1 U21390 ( .A1(n18315), .A2(n13596), .ZN(n18292) );
  OAI211_X1 U21391 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n18292), .B(n18277), .ZN(n18278) );
  OAI211_X1 U21392 ( .C1(n19290), .C2(n18739), .A(n18279), .B(n18278), .ZN(
        n18280) );
  AOI21_X1 U21393 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n18294), .A(
        n18280), .ZN(n18282) );
  NAND3_X1 U21394 ( .A1(n18320), .A2(n18522), .A3(n18531), .ZN(n18281) );
  OAI211_X1 U21395 ( .C1(n18451), .C2(n18536), .A(n18282), .B(n18281), .ZN(
        P3_U2808) );
  INV_X1 U21396 ( .A(n18331), .ZN(n18285) );
  INV_X1 U21397 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18577) );
  INV_X1 U21398 ( .A(n18573), .ZN(n18283) );
  NOR4_X1 U21399 ( .A1(n18343), .A2(n18577), .A3(n18357), .A4(n18283), .ZN(
        n18311) );
  AOI22_X1 U21400 ( .A1(n18285), .A2(n18284), .B1(n18311), .B2(n18542), .ZN(
        n18287) );
  XNOR2_X1 U21401 ( .A(n18287), .B(n18286), .ZN(n18546) );
  OAI22_X1 U21402 ( .A1(n18739), .A2(n19289), .B1(n18377), .B2(n10203), .ZN(
        n18289) );
  AOI221_X1 U21403 ( .B1(n18292), .B2(n18291), .C1(n18290), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n18289), .ZN(n18296) );
  NOR3_X1 U21404 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18519), .A3(
        n18293), .ZN(n18537) );
  AOI22_X1 U21405 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18294), .B1(
        n18320), .B2(n18537), .ZN(n18295) );
  OAI211_X1 U21406 ( .C1(n18546), .C2(n18451), .A(n18296), .B(n18295), .ZN(
        P3_U2809) );
  INV_X1 U21407 ( .A(n18330), .ZN(n18310) );
  NAND2_X1 U21408 ( .A1(n18310), .A2(n18299), .ZN(n18297) );
  OAI211_X1 U21409 ( .C1(n18311), .C2(n18299), .A(n18298), .B(n18297), .ZN(
        n18300) );
  XOR2_X1 U21410 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n18300), .Z(
        n18558) );
  INV_X1 U21411 ( .A(n18301), .ZN(n18304) );
  AOI221_X1 U21412 ( .B1(n18304), .B2(n18303), .C1(n18857), .C2(n18303), .A(
        n18302), .ZN(n18305) );
  NOR2_X1 U21413 ( .A1(n18739), .A2(n19286), .ZN(n18547) );
  AOI211_X1 U21414 ( .C1(n18306), .C2(n18426), .A(n18305), .B(n18547), .ZN(
        n18309) );
  NAND2_X1 U21415 ( .A1(n18538), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n18551) );
  INV_X1 U21416 ( .A(n18551), .ZN(n18521) );
  OAI21_X1 U21417 ( .B1(n18307), .B2(n18521), .A(n18329), .ZN(n18321) );
  NOR2_X1 U21418 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18551), .ZN(
        n18548) );
  AOI22_X1 U21419 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18321), .B1(
        n18320), .B2(n18548), .ZN(n18308) );
  OAI211_X1 U21420 ( .C1(n18451), .C2(n18558), .A(n18309), .B(n18308), .ZN(
        P3_U2810) );
  NOR2_X1 U21421 ( .A1(n18331), .A2(n18310), .ZN(n18334) );
  NOR2_X1 U21422 ( .A1(n18334), .A2(n18311), .ZN(n18312) );
  XOR2_X1 U21423 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B(n18312), .Z(
        n18564) );
  AOI21_X1 U21424 ( .B1(n18368), .B2(n9751), .A(n18478), .ZN(n18340) );
  OAI21_X1 U21425 ( .B1(n18314), .B2(n18313), .A(n18340), .ZN(n18326) );
  NOR2_X1 U21426 ( .A1(n18315), .A2(n9751), .ZN(n18328) );
  OAI211_X1 U21427 ( .C1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n18328), .B(n18316), .ZN(n18317) );
  NAND2_X1 U21428 ( .A1(n18693), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18562) );
  OAI211_X1 U21429 ( .C1(n18377), .C2(n18318), .A(n18317), .B(n18562), .ZN(
        n18319) );
  AOI21_X1 U21430 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n18326), .A(
        n18319), .ZN(n18323) );
  NOR2_X1 U21431 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18519), .ZN(
        n18559) );
  AOI22_X1 U21432 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18321), .B1(
        n18320), .B2(n18559), .ZN(n18322) );
  OAI211_X1 U21433 ( .C1(n18564), .C2(n18451), .A(n18323), .B(n18322), .ZN(
        P3_U2811) );
  NAND2_X1 U21434 ( .A1(n18573), .A2(n18577), .ZN(n18582) );
  INV_X1 U21435 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n18327) );
  OAI22_X1 U21436 ( .A1(n18739), .A2(n19283), .B1(n18377), .B2(n18324), .ZN(
        n18325) );
  AOI221_X1 U21437 ( .B1(n18328), .B2(n18327), .C1(n18326), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n18325), .ZN(n18337) );
  NOR2_X1 U21438 ( .A1(n18357), .A2(n18577), .ZN(n18333) );
  NOR2_X1 U21439 ( .A1(n18333), .A2(n18330), .ZN(n18332) );
  MUX2_X1 U21440 ( .A(n18333), .B(n18332), .S(n18331), .Z(n18335) );
  OR2_X1 U21441 ( .A1(n18335), .A2(n18334), .ZN(n18578) );
  AOI22_X1 U21442 ( .A1(n18347), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B1(
        n18428), .B2(n18578), .ZN(n18336) );
  OAI211_X1 U21443 ( .C1(n18350), .C2(n18582), .A(n18337), .B(n18336), .ZN(
        P3_U2812) );
  NAND2_X1 U21444 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18583), .ZN(
        n18589) );
  AOI21_X1 U21445 ( .B1(n18338), .B2(n16992), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18341) );
  OAI22_X1 U21446 ( .A1(n18341), .A2(n18340), .B1(n18490), .B2(n18339), .ZN(
        n18342) );
  AOI21_X1 U21447 ( .B1(n18693), .B2(P3_REIP_REG_17__SCAN_IN), .A(n18342), 
        .ZN(n18349) );
  AOI22_X1 U21448 ( .A1(n18344), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B1(
        n18573), .B2(n18343), .ZN(n18346) );
  NAND2_X1 U21449 ( .A1(n18346), .A2(n18345), .ZN(n18586) );
  AOI22_X1 U21450 ( .A1(n18347), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B1(
        n18428), .B2(n18586), .ZN(n18348) );
  OAI211_X1 U21451 ( .C1(n18350), .C2(n18589), .A(n18349), .B(n18348), .ZN(
        P3_U2813) );
  OAI221_X1 U21452 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n9659), .A(n18351), .ZN(
        n18628) );
  NAND2_X1 U21453 ( .A1(n18352), .A2(n18400), .ZN(n18404) );
  AOI221_X1 U21454 ( .B1(n18373), .B2(n18354), .C1(n18404), .C2(n18354), .A(
        n18353), .ZN(n18355) );
  NOR2_X1 U21455 ( .A1(n18739), .A2(n19275), .ZN(n18621) );
  AOI211_X1 U21456 ( .C1(n18356), .C2(n18426), .A(n18355), .B(n18621), .ZN(
        n18364) );
  INV_X1 U21457 ( .A(n18600), .ZN(n18615) );
  OR2_X1 U21458 ( .A1(n18652), .A2(n18357), .ZN(n18434) );
  OAI22_X1 U21459 ( .A1(n18358), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n18615), .B2(n18434), .ZN(n18359) );
  XNOR2_X1 U21460 ( .A(n18359), .B(n18619), .ZN(n18625) );
  AOI21_X1 U21461 ( .B1(n18360), .B2(n18600), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18362) );
  NOR2_X1 U21462 ( .A1(n18362), .A2(n9586), .ZN(n18623) );
  AOI22_X1 U21463 ( .A1(n18428), .A2(n18625), .B1(n18405), .B2(n18623), .ZN(
        n18363) );
  OAI211_X1 U21464 ( .C1(n18381), .C2(n18628), .A(n18364), .B(n18363), .ZN(
        P3_U2816) );
  INV_X1 U21465 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18644) );
  NOR2_X1 U21466 ( .A1(n18652), .A2(n18630), .ZN(n18632) );
  AOI22_X1 U21467 ( .A1(n18392), .A2(n18644), .B1(n18365), .B2(n18632), .ZN(
        n18366) );
  XNOR2_X1 U21468 ( .A(n18366), .B(n18384), .ZN(n18639) );
  AOI22_X1 U21469 ( .A1(n18370), .A2(n18369), .B1(n18368), .B2(n18367), .ZN(
        n18371) );
  NAND2_X1 U21470 ( .A1(n18372), .A2(n18371), .ZN(n18389) );
  NOR2_X1 U21471 ( .A1(n18739), .A2(n19273), .ZN(n18379) );
  OAI21_X1 U21472 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n18373), .ZN(n18374) );
  OAI22_X1 U21473 ( .A1(n18377), .A2(n18376), .B1(n18375), .B2(n18374), .ZN(
        n18378) );
  AOI211_X1 U21474 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n18389), .A(
        n18379), .B(n18378), .ZN(n18386) );
  OAI22_X1 U21475 ( .A1(n9659), .A2(n18381), .B1(n18632), .B2(n18380), .ZN(
        n18395) );
  INV_X1 U21476 ( .A(n18438), .ZN(n18382) );
  OAI21_X1 U21477 ( .B1(n18382), .B2(n18630), .A(n18384), .ZN(n18383) );
  OAI21_X1 U21478 ( .B1(n18395), .B2(n18384), .A(n18383), .ZN(n18385) );
  OAI211_X1 U21479 ( .C1(n18451), .C2(n18639), .A(n18386), .B(n18385), .ZN(
        P3_U2817) );
  AOI22_X1 U21480 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18389), .B1(
        n18388), .B2(n18387), .ZN(n18399) );
  AOI22_X1 U21481 ( .A1(n18693), .A2(P3_REIP_REG_12__SCAN_IN), .B1(n18391), 
        .B2(n18390), .ZN(n18398) );
  NOR2_X1 U21482 ( .A1(n18434), .A2(n18676), .ZN(n18433) );
  NOR2_X1 U21483 ( .A1(n18409), .A2(n18415), .ZN(n18393) );
  AOI21_X1 U21484 ( .B1(n18433), .B2(n18393), .A(n18392), .ZN(n18394) );
  XNOR2_X1 U21485 ( .A(n18394), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n18640) );
  AOI22_X1 U21486 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18395), .B1(
        n18428), .B2(n18640), .ZN(n18397) );
  NAND3_X1 U21487 ( .A1(n18438), .A2(n18664), .A3(n18644), .ZN(n18396) );
  NAND4_X1 U21488 ( .A1(n18399), .A2(n18398), .A3(n18397), .A4(n18396), .ZN(
        P3_U2818) );
  NAND2_X1 U21489 ( .A1(n18401), .A2(n18400), .ZN(n18439) );
  NOR2_X1 U21490 ( .A1(n18440), .A2(n18439), .ZN(n18420) );
  NAND2_X1 U21491 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n18420), .ZN(
        n18423) );
  OAI21_X1 U21492 ( .B1(n18455), .B2(n18402), .A(n18423), .ZN(n18403) );
  AOI22_X1 U21493 ( .A1(n18693), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18404), 
        .B2(n18403), .ZN(n18418) );
  NAND2_X1 U21494 ( .A1(n18438), .A2(n18649), .ZN(n18408) );
  AND2_X1 U21495 ( .A1(n18405), .A2(n18652), .ZN(n18406) );
  AOI21_X1 U21496 ( .B1(n18407), .B2(n9600), .A(n18406), .ZN(n18448) );
  AND2_X1 U21497 ( .A1(n18408), .A2(n18448), .ZN(n18432) );
  NOR2_X1 U21498 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18649), .ZN(
        n18648) );
  NAND2_X1 U21499 ( .A1(n18433), .A2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n18411) );
  NOR2_X1 U21500 ( .A1(n18437), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n18424) );
  NAND2_X1 U21501 ( .A1(n18424), .A2(n18409), .ZN(n18410) );
  NAND2_X1 U21502 ( .A1(n18411), .A2(n18410), .ZN(n18412) );
  XNOR2_X1 U21503 ( .A(n18412), .B(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18668) );
  INV_X1 U21504 ( .A(n18668), .ZN(n18413) );
  AOI22_X1 U21505 ( .A1(n18438), .A2(n18648), .B1(n18428), .B2(n18413), .ZN(
        n18414) );
  OAI21_X1 U21506 ( .B1(n18432), .B2(n18415), .A(n18414), .ZN(n18416) );
  INV_X1 U21507 ( .A(n18416), .ZN(n18417) );
  OAI211_X1 U21508 ( .C1(n18490), .C2(n18419), .A(n18418), .B(n18417), .ZN(
        P3_U2819) );
  AOI21_X1 U21509 ( .B1(n18438), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18431) );
  INV_X1 U21510 ( .A(n18420), .ZN(n18442) );
  OAI21_X1 U21511 ( .B1(n18455), .B2(n18421), .A(n18442), .ZN(n18422) );
  AOI22_X1 U21512 ( .A1(n18693), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n18423), 
        .B2(n18422), .ZN(n18430) );
  NOR2_X1 U21513 ( .A1(n18433), .A2(n18424), .ZN(n18425) );
  XNOR2_X1 U21514 ( .A(n18425), .B(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n18671) );
  AOI22_X1 U21515 ( .A1(n18428), .A2(n18671), .B1(n18427), .B2(n18426), .ZN(
        n18429) );
  OAI211_X1 U21516 ( .C1(n18432), .C2(n18431), .A(n18430), .B(n18429), .ZN(
        P3_U2820) );
  INV_X1 U21517 ( .A(n18433), .ZN(n18436) );
  NAND3_X1 U21518 ( .A1(n18437), .A2(n18434), .A3(n18676), .ZN(n18435) );
  OAI211_X1 U21519 ( .C1(n18676), .C2(n18437), .A(n18436), .B(n18435), .ZN(
        n18690) );
  NAND2_X1 U21520 ( .A1(n18438), .A2(n18676), .ZN(n18447) );
  OAI21_X1 U21521 ( .B1(n18455), .B2(n18440), .A(n18439), .ZN(n18441) );
  AOI22_X1 U21522 ( .A1(n18693), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n18442), 
        .B2(n18441), .ZN(n18443) );
  OAI21_X1 U21523 ( .B1(n18490), .B2(n18444), .A(n18443), .ZN(n18445) );
  INV_X1 U21524 ( .A(n18445), .ZN(n18446) );
  OAI211_X1 U21525 ( .C1(n18448), .C2(n18676), .A(n18447), .B(n18446), .ZN(
        n18449) );
  INV_X1 U21526 ( .A(n18449), .ZN(n18450) );
  OAI21_X1 U21527 ( .B1(n18690), .B2(n18451), .A(n18450), .ZN(P3_U2821) );
  NAND2_X1 U21528 ( .A1(n18456), .A2(n16992), .ZN(n18452) );
  OAI22_X1 U21529 ( .A1(n18488), .A2(n18453), .B1(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18452), .ZN(n18454) );
  AOI21_X1 U21530 ( .B1(n18693), .B2(P3_REIP_REG_6__SCAN_IN), .A(n18454), .ZN(
        n18459) );
  AOI21_X1 U21531 ( .B1(n16992), .B2(n18456), .A(n18455), .ZN(n18466) );
  AOI22_X1 U21532 ( .A1(n9600), .A2(n18457), .B1(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18466), .ZN(n18458) );
  OAI211_X1 U21533 ( .C1(n18490), .C2(n18460), .A(n18459), .B(n18458), .ZN(
        P3_U2824) );
  XOR2_X1 U21534 ( .A(n18461), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(
        n18694) );
  AOI22_X1 U21535 ( .A1(n18473), .A2(n18694), .B1(n18693), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n18468) );
  AOI21_X1 U21536 ( .B1(n9760), .B2(n18463), .A(n18462), .ZN(n18692) );
  OAI21_X1 U21537 ( .B1(n18478), .B2(n17012), .A(n18464), .ZN(n18465) );
  AOI22_X1 U21538 ( .A1(n9600), .A2(n18692), .B1(n18466), .B2(n18465), .ZN(
        n18467) );
  OAI211_X1 U21539 ( .C1(n18490), .C2(n18469), .A(n18468), .B(n18467), .ZN(
        P3_U2825) );
  NAND2_X1 U21540 ( .A1(n18471), .A2(n18470), .ZN(n18472) );
  XNOR2_X1 U21541 ( .A(n18472), .B(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n18703) );
  AOI22_X1 U21542 ( .A1(n18693), .A2(P3_REIP_REG_3__SCAN_IN), .B1(n18473), 
        .B2(n18703), .ZN(n18482) );
  AOI21_X1 U21543 ( .B1(n18476), .B2(n18475), .A(n18474), .ZN(n18702) );
  OAI21_X1 U21544 ( .B1(n18478), .B2(n18496), .A(n18477), .ZN(n18479) );
  AOI22_X1 U21545 ( .A1(n9600), .A2(n18702), .B1(n18480), .B2(n18479), .ZN(
        n18481) );
  OAI211_X1 U21546 ( .C1(n18490), .C2(n18483), .A(n18482), .B(n18481), .ZN(
        P3_U2827) );
  XNOR2_X1 U21547 ( .A(n18485), .B(n18484), .ZN(n18722) );
  NAND2_X1 U21548 ( .A1(n18693), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18725) );
  INV_X1 U21549 ( .A(n18725), .ZN(n18492) );
  XNOR2_X1 U21550 ( .A(n18487), .B(n18486), .ZN(n18721) );
  OAI22_X1 U21551 ( .A1(n18490), .A2(n18489), .B1(n18721), .B2(n18488), .ZN(
        n18491) );
  AOI211_X1 U21552 ( .C1(n9600), .C2(n18722), .A(n18492), .B(n18491), .ZN(
        n18494) );
  OAI221_X1 U21553 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18857), .C1(
        n18496), .C2(n18495), .A(n18494), .ZN(P3_U2828) );
  OAI22_X1 U21554 ( .A1(n18689), .A2(n18498), .B1(n18629), .B2(n18497), .ZN(
        n18511) );
  NOR3_X1 U21555 ( .A1(n18500), .A2(n18501), .A3(n18499), .ZN(n18506) );
  INV_X1 U21556 ( .A(n18501), .ZN(n18504) );
  OAI211_X1 U21557 ( .C1(n18504), .C2(n18712), .A(n18503), .B(n18502), .ZN(
        n18505) );
  OAI221_X1 U21558 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n18506), 
        .C1(n18509), .C2(n18505), .A(n18724), .ZN(n18507) );
  OAI211_X1 U21559 ( .C1(n18729), .C2(n18509), .A(n18508), .B(n18507), .ZN(
        n18510) );
  NOR2_X1 U21560 ( .A1(n18511), .A2(n18510), .ZN(n18512) );
  OAI21_X1 U21561 ( .B1(n18513), .B2(n18622), .A(n18512), .ZN(P3_U2837) );
  AOI21_X1 U21562 ( .B1(n18514), .B2(n18729), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18518) );
  AOI22_X1 U21563 ( .A1(n18693), .A2(P3_REIP_REG_23__SCAN_IN), .B1(n18672), 
        .B2(n18515), .ZN(n18516) );
  OAI21_X1 U21564 ( .B1(n18518), .B2(n18517), .A(n18516), .ZN(P3_U2839) );
  INV_X1 U21565 ( .A(n18669), .ZN(n18663) );
  OAI21_X1 U21566 ( .B1(n18519), .B2(n18571), .A(n19179), .ZN(n18520) );
  OAI221_X1 U21567 ( .B1(n18730), .B2(n18570), .C1(n18730), .C2(n18521), .A(
        n18520), .ZN(n18549) );
  NAND2_X1 U21568 ( .A1(n18524), .A2(n18655), .ZN(n18550) );
  INV_X1 U21569 ( .A(n18550), .ZN(n18661) );
  OAI22_X1 U21570 ( .A1(n18730), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n18522), .B2(n18661), .ZN(n18523) );
  NOR2_X1 U21571 ( .A1(n18549), .A2(n18523), .ZN(n18541) );
  NOR2_X1 U21572 ( .A1(n18525), .A2(n18524), .ZN(n18603) );
  AOI21_X1 U21573 ( .B1(n18609), .B2(n19178), .A(n18603), .ZN(n18539) );
  OAI211_X1 U21574 ( .C1(n18526), .C2(n18663), .A(n18541), .B(n18539), .ZN(
        n18527) );
  AOI211_X1 U21575 ( .C1(n18528), .C2(n18658), .A(n18527), .B(n18531), .ZN(
        n18529) );
  AOI221_X1 U21576 ( .B1(n18532), .B2(n18531), .C1(n18530), .C2(n18531), .A(
        n18529), .ZN(n18533) );
  AOI22_X1 U21577 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18701), .B1(
        n18724), .B2(n18533), .ZN(n18535) );
  NAND2_X1 U21578 ( .A1(n18693), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n18534) );
  OAI211_X1 U21579 ( .C1(n18536), .C2(n18689), .A(n18535), .B(n18534), .ZN(
        P3_U2840) );
  AOI22_X1 U21580 ( .A1(n18693), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n18560), 
        .B2(n18537), .ZN(n18545) );
  AOI21_X1 U21581 ( .B1(n18538), .B2(n18592), .A(n18683), .ZN(n18540) );
  NAND2_X1 U21582 ( .A1(n18539), .A2(n18724), .ZN(n18594) );
  NOR2_X1 U21583 ( .A1(n18540), .A2(n18594), .ZN(n18553) );
  OAI211_X1 U21584 ( .C1(n18554), .C2(n18542), .A(n18541), .B(n18553), .ZN(
        n18543) );
  NAND3_X1 U21585 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18739), .A3(
        n18543), .ZN(n18544) );
  OAI211_X1 U21586 ( .C1(n18546), .C2(n18689), .A(n18545), .B(n18544), .ZN(
        P3_U2841) );
  AOI21_X1 U21587 ( .B1(n18548), .B2(n18560), .A(n18547), .ZN(n18557) );
  AOI21_X1 U21588 ( .B1(n18551), .B2(n18550), .A(n18549), .ZN(n18552) );
  AOI21_X1 U21589 ( .B1(n18553), .B2(n18552), .A(n18693), .ZN(n18561) );
  NOR3_X1 U21590 ( .A1(n18554), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n19349), .ZN(n18555) );
  OAI21_X1 U21591 ( .B1(n18561), .B2(n18555), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18556) );
  OAI211_X1 U21592 ( .C1(n18558), .C2(n18689), .A(n18557), .B(n18556), .ZN(
        P3_U2842) );
  AOI22_X1 U21593 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18561), .B1(
        n18560), .B2(n18559), .ZN(n18563) );
  OAI211_X1 U21594 ( .C1(n18564), .C2(n18689), .A(n18563), .B(n18562), .ZN(
        P3_U2843) );
  NOR2_X1 U21595 ( .A1(n18566), .A2(n18565), .ZN(n18601) );
  NAND2_X1 U21596 ( .A1(n18568), .A2(n18677), .ZN(n18599) );
  NAND3_X1 U21597 ( .A1(n18570), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n18569), .ZN(n18575) );
  NAND2_X1 U21598 ( .A1(n19179), .A2(n18571), .ZN(n18572) );
  AOI22_X1 U21599 ( .A1(n18573), .A2(n18572), .B1(n18661), .B2(n18712), .ZN(
        n18574) );
  AOI211_X1 U21600 ( .C1(n18576), .C2(n18575), .A(n18574), .B(n18594), .ZN(
        n18584) );
  AOI221_X1 U21601 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18584), 
        .C1(n18713), .C2(n18584), .A(n18577), .ZN(n18579) );
  AOI22_X1 U21602 ( .A1(n18579), .A2(n18739), .B1(n18672), .B2(n18578), .ZN(
        n18581) );
  NAND2_X1 U21603 ( .A1(n18693), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18580) );
  OAI211_X1 U21604 ( .C1(n18582), .C2(n18599), .A(n18581), .B(n18580), .ZN(
        P3_U2844) );
  NOR3_X1 U21605 ( .A1(n18584), .A2(n18693), .A3(n18583), .ZN(n18585) );
  AOI21_X1 U21606 ( .B1(n18672), .B2(n18586), .A(n18585), .ZN(n18588) );
  NAND2_X1 U21607 ( .A1(n18693), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n18587) );
  OAI211_X1 U21608 ( .C1(n18589), .C2(n18599), .A(n18588), .B(n18587), .ZN(
        P3_U2845) );
  INV_X1 U21609 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18598) );
  OAI21_X1 U21610 ( .B1(n18678), .B2(n18679), .A(n18680), .ZN(n18660) );
  OAI21_X1 U21611 ( .B1(n18650), .B2(n18712), .A(n18660), .ZN(n18613) );
  AOI21_X1 U21612 ( .B1(n18590), .B2(n18669), .A(n18613), .ZN(n18591) );
  OAI211_X1 U21613 ( .C1(n18592), .C2(n18683), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n18591), .ZN(n18604) );
  OAI221_X1 U21614 ( .B1(n18594), .B2(n18593), .C1(n18594), .C2(n18604), .A(
        n18739), .ZN(n18597) );
  AOI22_X1 U21615 ( .A1(n18693), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n18672), 
        .B2(n18595), .ZN(n18596) );
  OAI221_X1 U21616 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18599), 
        .C1(n18598), .C2(n18597), .A(n18596), .ZN(P3_U2846) );
  NAND2_X1 U21617 ( .A1(n18601), .A2(n18600), .ZN(n18618) );
  OAI21_X1 U21618 ( .B1(n18619), .B2(n18618), .A(n16978), .ZN(n18605) );
  AOI22_X1 U21619 ( .A1(n18605), .A2(n18604), .B1(n18603), .B2(n18602), .ZN(
        n18612) );
  OAI22_X1 U21620 ( .A1(n18739), .A2(n19277), .B1(n16978), .B2(n18729), .ZN(
        n18606) );
  AOI21_X1 U21621 ( .B1(n18672), .B2(n18607), .A(n18606), .ZN(n18611) );
  NAND3_X1 U21622 ( .A1(n18728), .A2(n18609), .A3(n18608), .ZN(n18610) );
  OAI211_X1 U21623 ( .C1(n18612), .C2(n18616), .A(n18611), .B(n18610), .ZN(
        P3_U2847) );
  AOI221_X1 U21624 ( .B1(n18630), .B2(n18658), .C1(n18657), .C2(n18658), .A(
        n18613), .ZN(n18635) );
  OAI211_X1 U21625 ( .C1(n18683), .C2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n18635), .ZN(n18614) );
  AOI21_X1 U21626 ( .B1(n18669), .B2(n18615), .A(n18614), .ZN(n18617) );
  AOI211_X1 U21627 ( .C1(n18619), .C2(n18618), .A(n18617), .B(n18616), .ZN(
        n18620) );
  AOI211_X1 U21628 ( .C1(n18701), .C2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n18621), .B(n18620), .ZN(n18627) );
  INV_X1 U21629 ( .A(n18622), .ZN(n18624) );
  AOI22_X1 U21630 ( .A1(n18625), .A2(n18672), .B1(n18624), .B2(n18623), .ZN(
        n18626) );
  OAI211_X1 U21631 ( .C1(n18629), .C2(n18628), .A(n18627), .B(n18626), .ZN(
        P3_U2848) );
  NOR2_X1 U21632 ( .A1(n18630), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18631) );
  AOI22_X1 U21633 ( .A1(n18693), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18677), 
        .B2(n18631), .ZN(n18638) );
  INV_X1 U21634 ( .A(n18632), .ZN(n18633) );
  INV_X1 U21635 ( .A(n18664), .ZN(n18641) );
  AOI22_X1 U21636 ( .A1(n18653), .A2(n18633), .B1(n18641), .B2(n18669), .ZN(
        n18634) );
  OAI211_X1 U21637 ( .C1(n9659), .C2(n18655), .A(n18635), .B(n18634), .ZN(
        n18643) );
  OAI21_X1 U21638 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18663), .A(
        n18724), .ZN(n18636) );
  OAI211_X1 U21639 ( .C1(n18643), .C2(n18636), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18739), .ZN(n18637) );
  OAI211_X1 U21640 ( .C1(n18639), .C2(n18689), .A(n18638), .B(n18637), .ZN(
        P3_U2849) );
  AOI22_X1 U21641 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18701), .B1(
        n18672), .B2(n18640), .ZN(n18647) );
  NOR2_X1 U21642 ( .A1(n18642), .A2(n18641), .ZN(n18645) );
  OAI221_X1 U21643 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18645), 
        .C1(n18644), .C2(n18643), .A(n18724), .ZN(n18646) );
  OAI211_X1 U21644 ( .C1(n19271), .C2(n18739), .A(n18647), .B(n18646), .ZN(
        P3_U2850) );
  AOI22_X1 U21645 ( .A1(n18693), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18677), 
        .B2(n18648), .ZN(n18667) );
  INV_X1 U21646 ( .A(n18649), .ZN(n18662) );
  OAI21_X1 U21647 ( .B1(n18650), .B2(n18712), .A(n18724), .ZN(n18651) );
  AOI21_X1 U21648 ( .B1(n18653), .B2(n18652), .A(n18651), .ZN(n18654) );
  OAI21_X1 U21649 ( .B1(n18656), .B2(n18655), .A(n18654), .ZN(n18686) );
  AOI221_X1 U21650 ( .B1(n18676), .B2(n18658), .C1(n18657), .C2(n18658), .A(
        n18686), .ZN(n18659) );
  OAI211_X1 U21651 ( .C1(n18662), .C2(n18661), .A(n18660), .B(n18659), .ZN(
        n18670) );
  OAI22_X1 U21652 ( .A1(n18683), .A2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n18664), .B2(n18663), .ZN(n18665) );
  OAI211_X1 U21653 ( .C1(n18670), .C2(n18665), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18739), .ZN(n18666) );
  OAI211_X1 U21654 ( .C1(n18668), .C2(n18689), .A(n18667), .B(n18666), .ZN(
        P3_U2851) );
  OAI221_X1 U21655 ( .B1(n18670), .B2(n18676), .C1(n18670), .C2(n18669), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18675) );
  AOI22_X1 U21656 ( .A1(n18693), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n18672), 
        .B2(n18671), .ZN(n18674) );
  NAND3_X1 U21657 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18677), .A3(
        n18409), .ZN(n18673) );
  OAI211_X1 U21658 ( .C1(n18693), .C2(n18675), .A(n18674), .B(n18673), .ZN(
        P3_U2852) );
  AOI22_X1 U21659 ( .A1(n18693), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n18677), 
        .B2(n18676), .ZN(n18688) );
  NAND2_X1 U21660 ( .A1(n18680), .A2(n18678), .ZN(n18682) );
  NAND2_X1 U21661 ( .A1(n18680), .A2(n18679), .ZN(n18681) );
  OAI211_X1 U21662 ( .C1(n18684), .C2(n18683), .A(n18682), .B(n18681), .ZN(
        n18685) );
  OAI211_X1 U21663 ( .C1(n18686), .C2(n18685), .A(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B(n18739), .ZN(n18687) );
  OAI211_X1 U21664 ( .C1(n18690), .C2(n18689), .A(n18688), .B(n18687), .ZN(
        P3_U2853) );
  NAND4_X1 U21665 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18724), .A3(
        n18691), .A4(n18700), .ZN(n18698) );
  AOI22_X1 U21666 ( .A1(n18693), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n18728), 
        .B2(n18692), .ZN(n18697) );
  INV_X1 U21667 ( .A(n18734), .ZN(n18704) );
  AOI22_X1 U21668 ( .A1(n18695), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B1(
        n18704), .B2(n18694), .ZN(n18696) );
  OAI211_X1 U21669 ( .C1(n18699), .C2(n18698), .A(n18697), .B(n18696), .ZN(
        P3_U2857) );
  OAI21_X1 U21670 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n18700), .A(
        n18724), .ZN(n18707) );
  AOI22_X1 U21671 ( .A1(n18693), .A2(P3_REIP_REG_3__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n18701), .ZN(n18706) );
  AOI22_X1 U21672 ( .A1(n18704), .A2(n18703), .B1(n18728), .B2(n18702), .ZN(
        n18705) );
  OAI211_X1 U21673 ( .C1(n18708), .C2(n18707), .A(n18706), .B(n18705), .ZN(
        P3_U2859) );
  OR2_X1 U21674 ( .A1(n18710), .A2(n18709), .ZN(n18717) );
  NAND2_X1 U21675 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18711) );
  OAI22_X1 U21676 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18713), .B1(
        n18712), .B2(n18711), .ZN(n18714) );
  NOR2_X1 U21677 ( .A1(n18715), .A2(n18714), .ZN(n18716) );
  MUX2_X1 U21678 ( .A(n18717), .B(n18716), .S(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n18720) );
  NAND2_X1 U21679 ( .A1(n19179), .A2(n18718), .ZN(n18719) );
  OAI211_X1 U21680 ( .C1(n18721), .C2(n19183), .A(n18720), .B(n18719), .ZN(
        n18723) );
  AOI22_X1 U21681 ( .A1(n18724), .A2(n18723), .B1(n18728), .B2(n18722), .ZN(
        n18726) );
  OAI211_X1 U21682 ( .C1(n18729), .C2(n18727), .A(n18726), .B(n18725), .ZN(
        P3_U2860) );
  NAND2_X1 U21683 ( .A1(n18728), .A2(n18735), .ZN(n18733) );
  OAI21_X1 U21684 ( .B1(n18693), .B2(n18730), .A(n18729), .ZN(n18731) );
  NAND2_X1 U21685 ( .A1(n18731), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18732) );
  OAI211_X1 U21686 ( .C1(n18735), .C2(n18734), .A(n18733), .B(n18732), .ZN(
        n18736) );
  INV_X1 U21687 ( .A(n18736), .ZN(n18738) );
  OAI211_X1 U21688 ( .C1(n14108), .C2(n18739), .A(n18738), .B(n18737), .ZN(
        P3_U2862) );
  NAND2_X1 U21689 ( .A1(n12101), .A2(n18740), .ZN(n18742) );
  AOI21_X1 U21690 ( .B1(n18742), .B2(n21335), .A(n18741), .ZN(n19215) );
  OAI21_X1 U21691 ( .B1(n19215), .B2(n18791), .A(n18752), .ZN(n18743) );
  OAI221_X1 U21692 ( .B1(n21323), .B2(n19340), .C1(n21323), .C2(n18752), .A(
        n18743), .ZN(P3_U2863) );
  NAND2_X1 U21693 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18901) );
  AOI21_X1 U21694 ( .B1(n18901), .B2(n18745), .A(n18744), .ZN(n18751) );
  NOR3_X1 U21695 ( .A1(n12171), .A2(n18791), .A3(n18746), .ZN(n18747) );
  OAI21_X1 U21696 ( .B1(n18748), .B2(n18747), .A(n18752), .ZN(n18749) );
  AOI22_X1 U21697 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18751), .B1(
        n18749), .B2(n12172), .ZN(P3_U2865) );
  NAND2_X1 U21698 ( .A1(n19189), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18880) );
  INV_X1 U21699 ( .A(n18880), .ZN(n18927) );
  NOR2_X1 U21700 ( .A1(n19016), .A2(n18927), .ZN(n18750) );
  OAI22_X1 U21701 ( .A1(n18751), .A2(n19189), .B1(n18750), .B2(n18749), .ZN(
        P3_U2866) );
  NOR2_X1 U21702 ( .A1(n19188), .A2(n18752), .ZN(P3_U2867) );
  NOR2_X1 U21703 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19174) );
  NAND2_X1 U21704 ( .A1(n12172), .A2(n19189), .ZN(n18834) );
  INV_X1 U21705 ( .A(n18834), .ZN(n18792) );
  NAND2_X1 U21706 ( .A1(n19174), .A2(n18792), .ZN(n18790) );
  NOR2_X1 U21707 ( .A1(n18754), .A2(n18753), .ZN(n18784) );
  NAND2_X1 U21708 ( .A1(n18784), .A2(n18755), .ZN(n19118) );
  NOR2_X1 U21709 ( .A1(n19189), .A2(n18901), .ZN(n19113) );
  NAND2_X1 U21710 ( .A1(n21323), .A2(n19113), .ZN(n19108) );
  AND2_X1 U21711 ( .A1(n16992), .A2(BUF2_REG_16__SCAN_IN), .ZN(n19111) );
  NOR2_X2 U21712 ( .A1(n18856), .A2(n18756), .ZN(n19110) );
  NAND2_X1 U21713 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19113), .ZN(
        n19165) );
  AOI21_X1 U21714 ( .B1(n18790), .B2(n19165), .A(n19225), .ZN(n18786) );
  AOI22_X1 U21715 ( .A1(n19088), .A2(n19111), .B1(n19110), .B2(n18786), .ZN(
        n18759) );
  NOR2_X1 U21716 ( .A1(n12172), .A2(n19189), .ZN(n19062) );
  NOR2_X1 U21717 ( .A1(n21323), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18970) );
  NAND2_X1 U21718 ( .A1(n19062), .A2(n18970), .ZN(n19082) );
  INV_X1 U21719 ( .A(n19082), .ZN(n19160) );
  NOR2_X1 U21720 ( .A1(n19160), .A2(n19088), .ZN(n19083) );
  AOI221_X1 U21721 ( .B1(n19083), .B2(n19165), .C1(n19084), .C2(n19165), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18757) );
  OAI21_X1 U21722 ( .B1(n18851), .B2(n18757), .A(n19087), .ZN(n18787) );
  NOR2_X2 U21723 ( .A1(n16125), .A2(n18857), .ZN(n19115) );
  AOI22_X1 U21724 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18787), .B1(
        n19160), .B2(n19115), .ZN(n18758) );
  OAI211_X1 U21725 ( .C1(n18790), .C2(n19118), .A(n18759), .B(n18758), .ZN(
        P3_U2868) );
  NAND2_X1 U21726 ( .A1(n18784), .A2(n19335), .ZN(n19124) );
  AND2_X1 U21727 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n16992), .ZN(n19120) );
  AND2_X1 U21728 ( .A1(n19087), .A2(BUF2_REG_1__SCAN_IN), .ZN(n19119) );
  AOI22_X1 U21729 ( .A1(n19160), .A2(n19120), .B1(n18786), .B2(n19119), .ZN(
        n18761) );
  NOR2_X2 U21730 ( .A1(n18857), .A2(n16187), .ZN(n19121) );
  AOI22_X1 U21731 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18787), .B1(
        n19088), .B2(n19121), .ZN(n18760) );
  OAI211_X1 U21732 ( .C1(n18790), .C2(n19124), .A(n18761), .B(n18760), .ZN(
        P3_U2869) );
  NAND2_X1 U21733 ( .A1(n18762), .A2(n18784), .ZN(n19130) );
  AND2_X1 U21734 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n16992), .ZN(n19127) );
  NOR2_X2 U21735 ( .A1(n18856), .A2(n18763), .ZN(n19125) );
  AOI22_X1 U21736 ( .A1(n19160), .A2(n19127), .B1(n18786), .B2(n19125), .ZN(
        n18765) );
  NOR2_X2 U21737 ( .A1(n18857), .A2(n16178), .ZN(n19126) );
  AOI22_X1 U21738 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18787), .B1(
        n19088), .B2(n19126), .ZN(n18764) );
  OAI211_X1 U21739 ( .C1(n18790), .C2(n19130), .A(n18765), .B(n18764), .ZN(
        P3_U2870) );
  NAND2_X1 U21740 ( .A1(n18784), .A2(n18766), .ZN(n19136) );
  NOR2_X2 U21741 ( .A1(n16102), .A2(n18857), .ZN(n19133) );
  NOR2_X2 U21742 ( .A1(n18856), .A2(n18767), .ZN(n19131) );
  AOI22_X1 U21743 ( .A1(n19160), .A2(n19133), .B1(n18786), .B2(n19131), .ZN(
        n18769) );
  AND2_X1 U21744 ( .A1(n16992), .A2(BUF2_REG_19__SCAN_IN), .ZN(n19132) );
  AOI22_X1 U21745 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18787), .B1(
        n19088), .B2(n19132), .ZN(n18768) );
  OAI211_X1 U21746 ( .C1(n18790), .C2(n19136), .A(n18769), .B(n18768), .ZN(
        P3_U2871) );
  INV_X1 U21747 ( .A(n18770), .ZN(n18771) );
  NAND2_X1 U21748 ( .A1(n18771), .A2(n18784), .ZN(n19142) );
  NOR2_X2 U21749 ( .A1(n18857), .A2(n16872), .ZN(n19139) );
  NOR2_X2 U21750 ( .A1(n18856), .A2(n18772), .ZN(n19137) );
  AOI22_X1 U21751 ( .A1(n19088), .A2(n19139), .B1(n18786), .B2(n19137), .ZN(
        n18774) );
  AND2_X1 U21752 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n16992), .ZN(n19138) );
  AOI22_X1 U21753 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18787), .B1(
        n19160), .B2(n19138), .ZN(n18773) );
  OAI211_X1 U21754 ( .C1(n18790), .C2(n19142), .A(n18774), .B(n18773), .ZN(
        P3_U2872) );
  NAND2_X1 U21755 ( .A1(n18784), .A2(n18775), .ZN(n19148) );
  NOR2_X2 U21756 ( .A1(n16082), .A2(n18857), .ZN(n19145) );
  NOR2_X2 U21757 ( .A1(n18856), .A2(n18776), .ZN(n19143) );
  AOI22_X1 U21758 ( .A1(n19160), .A2(n19145), .B1(n18786), .B2(n19143), .ZN(
        n18778) );
  AOI22_X1 U21759 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18787), .B1(
        n19088), .B2(n19144), .ZN(n18777) );
  OAI211_X1 U21760 ( .C1(n18790), .C2(n19148), .A(n18778), .B(n18777), .ZN(
        P3_U2873) );
  NAND2_X1 U21761 ( .A1(n18784), .A2(n18779), .ZN(n19154) );
  NOR2_X2 U21762 ( .A1(n16142), .A2(n18857), .ZN(n19150) );
  NOR2_X2 U21763 ( .A1(n18780), .A2(n18856), .ZN(n19149) );
  AOI22_X1 U21764 ( .A1(n19088), .A2(n19150), .B1(n18786), .B2(n19149), .ZN(
        n18782) );
  NOR2_X2 U21765 ( .A1(n16076), .A2(n18857), .ZN(n19151) );
  AOI22_X1 U21766 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18787), .B1(
        n19160), .B2(n19151), .ZN(n18781) );
  OAI211_X1 U21767 ( .C1(n18790), .C2(n19154), .A(n18782), .B(n18781), .ZN(
        P3_U2874) );
  NAND2_X1 U21768 ( .A1(n18784), .A2(n18783), .ZN(n19164) );
  NOR2_X2 U21769 ( .A1(n16132), .A2(n18857), .ZN(n19159) );
  NOR2_X2 U21770 ( .A1(n18785), .A2(n18856), .ZN(n19156) );
  AOI22_X1 U21771 ( .A1(n19088), .A2(n19159), .B1(n18786), .B2(n19156), .ZN(
        n18789) );
  NOR2_X2 U21772 ( .A1(n18857), .A2(n19641), .ZN(n19158) );
  AOI22_X1 U21773 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18787), .B1(
        n19160), .B2(n19158), .ZN(n18788) );
  OAI211_X1 U21774 ( .C1(n18790), .C2(n19164), .A(n18789), .B(n18788), .ZN(
        P3_U2875) );
  NAND2_X1 U21775 ( .A1(n18970), .A2(n18792), .ZN(n18811) );
  NAND2_X1 U21776 ( .A1(n12171), .A2(n19109), .ZN(n19059) );
  NOR2_X1 U21777 ( .A1(n18834), .A2(n19059), .ZN(n18807) );
  AOI22_X1 U21778 ( .A1(n19115), .A2(n19088), .B1(n19110), .B2(n18807), .ZN(
        n18794) );
  NOR2_X1 U21779 ( .A1(n18856), .A2(n18791), .ZN(n19112) );
  AND2_X1 U21780 ( .A1(n12171), .A2(n19112), .ZN(n19061) );
  AOI22_X1 U21781 ( .A1(n16992), .A2(n19113), .B1(n18792), .B2(n19061), .ZN(
        n18808) );
  AOI22_X1 U21782 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18808), .B1(
        n18829), .B2(n19111), .ZN(n18793) );
  OAI211_X1 U21783 ( .C1(n19118), .C2(n18811), .A(n18794), .B(n18793), .ZN(
        P3_U2876) );
  AOI22_X1 U21784 ( .A1(n19088), .A2(n19120), .B1(n19119), .B2(n18807), .ZN(
        n18796) );
  AOI22_X1 U21785 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18808), .B1(
        n18829), .B2(n19121), .ZN(n18795) );
  OAI211_X1 U21786 ( .C1(n19124), .C2(n18811), .A(n18796), .B(n18795), .ZN(
        P3_U2877) );
  AOI22_X1 U21787 ( .A1(n18829), .A2(n19126), .B1(n19125), .B2(n18807), .ZN(
        n18798) );
  AOI22_X1 U21788 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18808), .B1(
        n19088), .B2(n19127), .ZN(n18797) );
  OAI211_X1 U21789 ( .C1(n19130), .C2(n18811), .A(n18798), .B(n18797), .ZN(
        P3_U2878) );
  AOI22_X1 U21790 ( .A1(n19088), .A2(n19133), .B1(n19131), .B2(n18807), .ZN(
        n18800) );
  AOI22_X1 U21791 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18808), .B1(
        n18829), .B2(n19132), .ZN(n18799) );
  OAI211_X1 U21792 ( .C1(n19136), .C2(n18811), .A(n18800), .B(n18799), .ZN(
        P3_U2879) );
  AOI22_X1 U21793 ( .A1(n19088), .A2(n19138), .B1(n19137), .B2(n18807), .ZN(
        n18802) );
  AOI22_X1 U21794 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18808), .B1(
        n18829), .B2(n19139), .ZN(n18801) );
  OAI211_X1 U21795 ( .C1(n19142), .C2(n18811), .A(n18802), .B(n18801), .ZN(
        P3_U2880) );
  AOI22_X1 U21796 ( .A1(n19088), .A2(n19145), .B1(n19143), .B2(n18807), .ZN(
        n18804) );
  AOI22_X1 U21797 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18808), .B1(
        n18829), .B2(n19144), .ZN(n18803) );
  OAI211_X1 U21798 ( .C1(n19148), .C2(n18811), .A(n18804), .B(n18803), .ZN(
        P3_U2881) );
  AOI22_X1 U21799 ( .A1(n19088), .A2(n19151), .B1(n19149), .B2(n18807), .ZN(
        n18806) );
  AOI22_X1 U21800 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18808), .B1(
        n18829), .B2(n19150), .ZN(n18805) );
  OAI211_X1 U21801 ( .C1(n19154), .C2(n18811), .A(n18806), .B(n18805), .ZN(
        P3_U2882) );
  AOI22_X1 U21802 ( .A1(n18829), .A2(n19159), .B1(n19156), .B2(n18807), .ZN(
        n18810) );
  AOI22_X1 U21803 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18808), .B1(
        n19088), .B2(n19158), .ZN(n18809) );
  OAI211_X1 U21804 ( .C1(n19164), .C2(n18811), .A(n18810), .B(n18809), .ZN(
        P3_U2883) );
  NOR2_X1 U21805 ( .A1(n12171), .A2(n18834), .ZN(n18881) );
  NAND2_X1 U21806 ( .A1(n18881), .A2(n21323), .ZN(n18833) );
  NOR2_X1 U21807 ( .A1(n18875), .A2(n18897), .ZN(n18858) );
  NOR2_X1 U21808 ( .A1(n19225), .A2(n18858), .ZN(n18828) );
  AOI22_X1 U21809 ( .A1(n19115), .A2(n18829), .B1(n19110), .B2(n18828), .ZN(
        n18815) );
  NOR2_X1 U21810 ( .A1(n18851), .A2(n18829), .ZN(n18812) );
  OAI21_X1 U21811 ( .B1(n18812), .B2(n19084), .A(n18858), .ZN(n18813) );
  OAI211_X1 U21812 ( .C1(n18897), .C2(n19322), .A(n19087), .B(n18813), .ZN(
        n18830) );
  AOI22_X1 U21813 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18830), .B1(
        n18851), .B2(n19111), .ZN(n18814) );
  OAI211_X1 U21814 ( .C1(n19118), .C2(n18833), .A(n18815), .B(n18814), .ZN(
        P3_U2884) );
  AOI22_X1 U21815 ( .A1(n18829), .A2(n19120), .B1(n19119), .B2(n18828), .ZN(
        n18817) );
  AOI22_X1 U21816 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18830), .B1(
        n18851), .B2(n19121), .ZN(n18816) );
  OAI211_X1 U21817 ( .C1(n19124), .C2(n18833), .A(n18817), .B(n18816), .ZN(
        P3_U2885) );
  AOI22_X1 U21818 ( .A1(n18851), .A2(n19126), .B1(n19125), .B2(n18828), .ZN(
        n18819) );
  AOI22_X1 U21819 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18830), .B1(
        n18829), .B2(n19127), .ZN(n18818) );
  OAI211_X1 U21820 ( .C1(n19130), .C2(n18833), .A(n18819), .B(n18818), .ZN(
        P3_U2886) );
  AOI22_X1 U21821 ( .A1(n18829), .A2(n19133), .B1(n19131), .B2(n18828), .ZN(
        n18821) );
  AOI22_X1 U21822 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18830), .B1(
        n18851), .B2(n19132), .ZN(n18820) );
  OAI211_X1 U21823 ( .C1(n19136), .C2(n18833), .A(n18821), .B(n18820), .ZN(
        P3_U2887) );
  AOI22_X1 U21824 ( .A1(n18851), .A2(n19139), .B1(n19137), .B2(n18828), .ZN(
        n18823) );
  AOI22_X1 U21825 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18830), .B1(
        n18829), .B2(n19138), .ZN(n18822) );
  OAI211_X1 U21826 ( .C1(n19142), .C2(n18833), .A(n18823), .B(n18822), .ZN(
        P3_U2888) );
  AOI22_X1 U21827 ( .A1(n18829), .A2(n19145), .B1(n19143), .B2(n18828), .ZN(
        n18825) );
  AOI22_X1 U21828 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18830), .B1(
        n18851), .B2(n19144), .ZN(n18824) );
  OAI211_X1 U21829 ( .C1(n19148), .C2(n18833), .A(n18825), .B(n18824), .ZN(
        P3_U2889) );
  AOI22_X1 U21830 ( .A1(n18829), .A2(n19151), .B1(n19149), .B2(n18828), .ZN(
        n18827) );
  AOI22_X1 U21831 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18830), .B1(
        n18851), .B2(n19150), .ZN(n18826) );
  OAI211_X1 U21832 ( .C1(n19154), .C2(n18833), .A(n18827), .B(n18826), .ZN(
        P3_U2890) );
  AOI22_X1 U21833 ( .A1(n18851), .A2(n19159), .B1(n19156), .B2(n18828), .ZN(
        n18832) );
  AOI22_X1 U21834 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18830), .B1(
        n18829), .B2(n19158), .ZN(n18831) );
  OAI211_X1 U21835 ( .C1(n19164), .C2(n18833), .A(n18832), .B(n18831), .ZN(
        P3_U2891) );
  NAND2_X1 U21836 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18881), .ZN(
        n18855) );
  AND2_X1 U21837 ( .A1(n19109), .A2(n18881), .ZN(n18850) );
  AOI22_X1 U21838 ( .A1(n19115), .A2(n18851), .B1(n19110), .B2(n18850), .ZN(
        n18837) );
  OAI21_X1 U21839 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18834), .A(n18855), 
        .ZN(n18835) );
  NAND3_X1 U21840 ( .A1(n19087), .A2(n18925), .A3(n18835), .ZN(n18852) );
  AOI22_X1 U21841 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18852), .B1(
        n19111), .B2(n18875), .ZN(n18836) );
  OAI211_X1 U21842 ( .C1(n19118), .C2(n18855), .A(n18837), .B(n18836), .ZN(
        P3_U2892) );
  AOI22_X1 U21843 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18852), .B1(
        n19119), .B2(n18850), .ZN(n18839) );
  AOI22_X1 U21844 ( .A1(n18851), .A2(n19120), .B1(n19121), .B2(n18875), .ZN(
        n18838) );
  OAI211_X1 U21845 ( .C1(n19124), .C2(n18855), .A(n18839), .B(n18838), .ZN(
        P3_U2893) );
  AOI22_X1 U21846 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18852), .B1(
        n19125), .B2(n18850), .ZN(n18841) );
  AOI22_X1 U21847 ( .A1(n18851), .A2(n19127), .B1(n19126), .B2(n18875), .ZN(
        n18840) );
  OAI211_X1 U21848 ( .C1(n19130), .C2(n18855), .A(n18841), .B(n18840), .ZN(
        P3_U2894) );
  AOI22_X1 U21849 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18852), .B1(
        n19131), .B2(n18850), .ZN(n18843) );
  AOI22_X1 U21850 ( .A1(n18851), .A2(n19133), .B1(n19132), .B2(n18875), .ZN(
        n18842) );
  OAI211_X1 U21851 ( .C1(n19136), .C2(n18855), .A(n18843), .B(n18842), .ZN(
        P3_U2895) );
  AOI22_X1 U21852 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18852), .B1(
        n19137), .B2(n18850), .ZN(n18845) );
  AOI22_X1 U21853 ( .A1(n18851), .A2(n19138), .B1(n19139), .B2(n18875), .ZN(
        n18844) );
  OAI211_X1 U21854 ( .C1(n19142), .C2(n18855), .A(n18845), .B(n18844), .ZN(
        P3_U2896) );
  AOI22_X1 U21855 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18852), .B1(
        n19143), .B2(n18850), .ZN(n18847) );
  AOI22_X1 U21856 ( .A1(n18851), .A2(n19145), .B1(n19144), .B2(n18875), .ZN(
        n18846) );
  OAI211_X1 U21857 ( .C1(n19148), .C2(n18855), .A(n18847), .B(n18846), .ZN(
        P3_U2897) );
  AOI22_X1 U21858 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18852), .B1(
        n19149), .B2(n18850), .ZN(n18849) );
  AOI22_X1 U21859 ( .A1(n18851), .A2(n19151), .B1(n19150), .B2(n18875), .ZN(
        n18848) );
  OAI211_X1 U21860 ( .C1(n19154), .C2(n18855), .A(n18849), .B(n18848), .ZN(
        P3_U2898) );
  AOI22_X1 U21861 ( .A1(n18851), .A2(n19158), .B1(n19156), .B2(n18850), .ZN(
        n18854) );
  AOI22_X1 U21862 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18852), .B1(
        n19159), .B2(n18875), .ZN(n18853) );
  OAI211_X1 U21863 ( .C1(n19164), .C2(n18855), .A(n18854), .B(n18853), .ZN(
        P3_U2899) );
  NAND2_X1 U21864 ( .A1(n19174), .A2(n18927), .ZN(n18879) );
  INV_X1 U21865 ( .A(n18855), .ZN(n18920) );
  NOR2_X1 U21866 ( .A1(n18920), .A2(n18944), .ZN(n18903) );
  NOR2_X1 U21867 ( .A1(n19225), .A2(n18903), .ZN(n18874) );
  AOI22_X1 U21868 ( .A1(n19110), .A2(n18874), .B1(n19111), .B2(n18897), .ZN(
        n18861) );
  OAI22_X1 U21869 ( .A1(n18858), .A2(n18857), .B1(n18903), .B2(n18856), .ZN(
        n18859) );
  OAI21_X1 U21870 ( .B1(n18944), .B2(n19322), .A(n18859), .ZN(n18876) );
  AOI22_X1 U21871 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18876), .B1(
        n19115), .B2(n18875), .ZN(n18860) );
  OAI211_X1 U21872 ( .C1(n19118), .C2(n18879), .A(n18861), .B(n18860), .ZN(
        P3_U2900) );
  AOI22_X1 U21873 ( .A1(n19120), .A2(n18875), .B1(n19119), .B2(n18874), .ZN(
        n18863) );
  AOI22_X1 U21874 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18876), .B1(
        n19121), .B2(n18897), .ZN(n18862) );
  OAI211_X1 U21875 ( .C1(n19124), .C2(n18879), .A(n18863), .B(n18862), .ZN(
        P3_U2901) );
  AOI22_X1 U21876 ( .A1(n19127), .A2(n18875), .B1(n19125), .B2(n18874), .ZN(
        n18865) );
  AOI22_X1 U21877 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18876), .B1(
        n19126), .B2(n18897), .ZN(n18864) );
  OAI211_X1 U21878 ( .C1(n19130), .C2(n18879), .A(n18865), .B(n18864), .ZN(
        P3_U2902) );
  AOI22_X1 U21879 ( .A1(n19133), .A2(n18875), .B1(n19131), .B2(n18874), .ZN(
        n18867) );
  AOI22_X1 U21880 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18876), .B1(
        n19132), .B2(n18897), .ZN(n18866) );
  OAI211_X1 U21881 ( .C1(n19136), .C2(n18879), .A(n18867), .B(n18866), .ZN(
        P3_U2903) );
  AOI22_X1 U21882 ( .A1(n19137), .A2(n18874), .B1(n19139), .B2(n18897), .ZN(
        n18869) );
  AOI22_X1 U21883 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18876), .B1(
        n19138), .B2(n18875), .ZN(n18868) );
  OAI211_X1 U21884 ( .C1(n19142), .C2(n18879), .A(n18869), .B(n18868), .ZN(
        P3_U2904) );
  AOI22_X1 U21885 ( .A1(n19143), .A2(n18874), .B1(n19145), .B2(n18875), .ZN(
        n18871) );
  AOI22_X1 U21886 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18876), .B1(
        n19144), .B2(n18897), .ZN(n18870) );
  OAI211_X1 U21887 ( .C1(n19148), .C2(n18879), .A(n18871), .B(n18870), .ZN(
        P3_U2905) );
  AOI22_X1 U21888 ( .A1(n19150), .A2(n18897), .B1(n19149), .B2(n18874), .ZN(
        n18873) );
  AOI22_X1 U21889 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18876), .B1(
        n19151), .B2(n18875), .ZN(n18872) );
  OAI211_X1 U21890 ( .C1(n19154), .C2(n18879), .A(n18873), .B(n18872), .ZN(
        P3_U2906) );
  AOI22_X1 U21891 ( .A1(n19159), .A2(n18897), .B1(n19156), .B2(n18874), .ZN(
        n18878) );
  AOI22_X1 U21892 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18876), .B1(
        n19158), .B2(n18875), .ZN(n18877) );
  OAI211_X1 U21893 ( .C1(n19164), .C2(n18879), .A(n18878), .B(n18877), .ZN(
        P3_U2907) );
  NAND2_X1 U21894 ( .A1(n18970), .A2(n18927), .ZN(n18902) );
  NOR2_X1 U21895 ( .A1(n18880), .A2(n19059), .ZN(n18896) );
  AOI22_X1 U21896 ( .A1(n19115), .A2(n18897), .B1(n19110), .B2(n18896), .ZN(
        n18883) );
  AOI22_X1 U21897 ( .A1(n16992), .A2(n18881), .B1(n18927), .B2(n19061), .ZN(
        n18898) );
  AOI22_X1 U21898 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18898), .B1(
        n19111), .B2(n18920), .ZN(n18882) );
  OAI211_X1 U21899 ( .C1(n19118), .C2(n18902), .A(n18883), .B(n18882), .ZN(
        P3_U2908) );
  AOI22_X1 U21900 ( .A1(n19120), .A2(n18897), .B1(n19119), .B2(n18896), .ZN(
        n18885) );
  AOI22_X1 U21901 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18898), .B1(
        n19121), .B2(n18920), .ZN(n18884) );
  OAI211_X1 U21902 ( .C1(n19124), .C2(n18902), .A(n18885), .B(n18884), .ZN(
        P3_U2909) );
  AOI22_X1 U21903 ( .A1(n19127), .A2(n18897), .B1(n19125), .B2(n18896), .ZN(
        n18887) );
  AOI22_X1 U21904 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18898), .B1(
        n19126), .B2(n18920), .ZN(n18886) );
  OAI211_X1 U21905 ( .C1(n19130), .C2(n18902), .A(n18887), .B(n18886), .ZN(
        P3_U2910) );
  AOI22_X1 U21906 ( .A1(n19133), .A2(n18897), .B1(n19131), .B2(n18896), .ZN(
        n18889) );
  AOI22_X1 U21907 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18898), .B1(
        n19132), .B2(n18920), .ZN(n18888) );
  OAI211_X1 U21908 ( .C1(n19136), .C2(n18902), .A(n18889), .B(n18888), .ZN(
        P3_U2911) );
  AOI22_X1 U21909 ( .A1(n19138), .A2(n18897), .B1(n19137), .B2(n18896), .ZN(
        n18891) );
  AOI22_X1 U21910 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18898), .B1(
        n19139), .B2(n18920), .ZN(n18890) );
  OAI211_X1 U21911 ( .C1(n19142), .C2(n18902), .A(n18891), .B(n18890), .ZN(
        P3_U2912) );
  AOI22_X1 U21912 ( .A1(n19144), .A2(n18920), .B1(n19143), .B2(n18896), .ZN(
        n18893) );
  AOI22_X1 U21913 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18898), .B1(
        n19145), .B2(n18897), .ZN(n18892) );
  OAI211_X1 U21914 ( .C1(n19148), .C2(n18902), .A(n18893), .B(n18892), .ZN(
        P3_U2913) );
  AOI22_X1 U21915 ( .A1(n19150), .A2(n18920), .B1(n19149), .B2(n18896), .ZN(
        n18895) );
  AOI22_X1 U21916 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18898), .B1(
        n19151), .B2(n18897), .ZN(n18894) );
  OAI211_X1 U21917 ( .C1(n19154), .C2(n18902), .A(n18895), .B(n18894), .ZN(
        P3_U2914) );
  AOI22_X1 U21918 ( .A1(n19158), .A2(n18897), .B1(n19156), .B2(n18896), .ZN(
        n18900) );
  AOI22_X1 U21919 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18898), .B1(
        n19159), .B2(n18920), .ZN(n18899) );
  OAI211_X1 U21920 ( .C1(n19164), .C2(n18902), .A(n18900), .B(n18899), .ZN(
        P3_U2915) );
  NOR2_X1 U21921 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18901), .ZN(
        n18972) );
  NAND2_X1 U21922 ( .A1(n18972), .A2(n21323), .ZN(n18924) );
  INV_X1 U21923 ( .A(n18924), .ZN(n18988) );
  NOR2_X1 U21924 ( .A1(n18965), .A2(n18988), .ZN(n18948) );
  NOR2_X1 U21925 ( .A1(n19225), .A2(n18948), .ZN(n18919) );
  AOI22_X1 U21926 ( .A1(n19110), .A2(n18919), .B1(n19111), .B2(n18944), .ZN(
        n18906) );
  OAI21_X1 U21927 ( .B1(n18903), .B2(n19084), .A(n18948), .ZN(n18904) );
  OAI211_X1 U21928 ( .C1(n18988), .C2(n19322), .A(n19087), .B(n18904), .ZN(
        n18921) );
  AOI22_X1 U21929 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18921), .B1(
        n19115), .B2(n18920), .ZN(n18905) );
  OAI211_X1 U21930 ( .C1(n19118), .C2(n18924), .A(n18906), .B(n18905), .ZN(
        P3_U2916) );
  AOI22_X1 U21931 ( .A1(n19120), .A2(n18920), .B1(n19119), .B2(n18919), .ZN(
        n18908) );
  AOI22_X1 U21932 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18921), .B1(
        n19121), .B2(n18944), .ZN(n18907) );
  OAI211_X1 U21933 ( .C1(n19124), .C2(n18924), .A(n18908), .B(n18907), .ZN(
        P3_U2917) );
  AOI22_X1 U21934 ( .A1(n19126), .A2(n18944), .B1(n19125), .B2(n18919), .ZN(
        n18910) );
  AOI22_X1 U21935 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18921), .B1(
        n19127), .B2(n18920), .ZN(n18909) );
  OAI211_X1 U21936 ( .C1(n19130), .C2(n18924), .A(n18910), .B(n18909), .ZN(
        P3_U2918) );
  AOI22_X1 U21937 ( .A1(n19133), .A2(n18920), .B1(n19131), .B2(n18919), .ZN(
        n18912) );
  AOI22_X1 U21938 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18921), .B1(
        n19132), .B2(n18944), .ZN(n18911) );
  OAI211_X1 U21939 ( .C1(n19136), .C2(n18924), .A(n18912), .B(n18911), .ZN(
        P3_U2919) );
  AOI22_X1 U21940 ( .A1(n19138), .A2(n18920), .B1(n19137), .B2(n18919), .ZN(
        n18914) );
  AOI22_X1 U21941 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18921), .B1(
        n19139), .B2(n18944), .ZN(n18913) );
  OAI211_X1 U21942 ( .C1(n19142), .C2(n18924), .A(n18914), .B(n18913), .ZN(
        P3_U2920) );
  AOI22_X1 U21943 ( .A1(n19143), .A2(n18919), .B1(n19145), .B2(n18920), .ZN(
        n18916) );
  AOI22_X1 U21944 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18921), .B1(
        n19144), .B2(n18944), .ZN(n18915) );
  OAI211_X1 U21945 ( .C1(n19148), .C2(n18924), .A(n18916), .B(n18915), .ZN(
        P3_U2921) );
  AOI22_X1 U21946 ( .A1(n19151), .A2(n18920), .B1(n19149), .B2(n18919), .ZN(
        n18918) );
  AOI22_X1 U21947 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18921), .B1(
        n19150), .B2(n18944), .ZN(n18917) );
  OAI211_X1 U21948 ( .C1(n19154), .C2(n18924), .A(n18918), .B(n18917), .ZN(
        P3_U2922) );
  AOI22_X1 U21949 ( .A1(n19159), .A2(n18944), .B1(n19156), .B2(n18919), .ZN(
        n18923) );
  AOI22_X1 U21950 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18921), .B1(
        n19158), .B2(n18920), .ZN(n18922) );
  OAI211_X1 U21951 ( .C1(n19164), .C2(n18924), .A(n18923), .B(n18922), .ZN(
        P3_U2923) );
  NAND2_X1 U21952 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18972), .ZN(
        n18947) );
  AND2_X1 U21953 ( .A1(n19109), .A2(n18972), .ZN(n18942) );
  AOI22_X1 U21954 ( .A1(n19110), .A2(n18942), .B1(n19111), .B2(n18965), .ZN(
        n18929) );
  INV_X1 U21955 ( .A(n18947), .ZN(n19010) );
  AND2_X1 U21956 ( .A1(n19087), .A2(n18925), .ZN(n18926) );
  OAI211_X1 U21957 ( .C1(n19010), .C2(n19322), .A(n18927), .B(n18926), .ZN(
        n18943) );
  AOI22_X1 U21958 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18943), .B1(
        n19115), .B2(n18944), .ZN(n18928) );
  OAI211_X1 U21959 ( .C1(n19118), .C2(n18947), .A(n18929), .B(n18928), .ZN(
        P3_U2924) );
  AOI22_X1 U21960 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18943), .B1(
        n19119), .B2(n18942), .ZN(n18931) );
  AOI22_X1 U21961 ( .A1(n19121), .A2(n18965), .B1(n19120), .B2(n18944), .ZN(
        n18930) );
  OAI211_X1 U21962 ( .C1(n19124), .C2(n18947), .A(n18931), .B(n18930), .ZN(
        P3_U2925) );
  AOI22_X1 U21963 ( .A1(n19127), .A2(n18944), .B1(n19125), .B2(n18942), .ZN(
        n18933) );
  AOI22_X1 U21964 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18943), .B1(
        n19126), .B2(n18965), .ZN(n18932) );
  OAI211_X1 U21965 ( .C1(n19130), .C2(n18947), .A(n18933), .B(n18932), .ZN(
        P3_U2926) );
  AOI22_X1 U21966 ( .A1(n19133), .A2(n18944), .B1(n19131), .B2(n18942), .ZN(
        n18935) );
  AOI22_X1 U21967 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18943), .B1(
        n19132), .B2(n18965), .ZN(n18934) );
  OAI211_X1 U21968 ( .C1(n19136), .C2(n18947), .A(n18935), .B(n18934), .ZN(
        P3_U2927) );
  AOI22_X1 U21969 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18943), .B1(
        n19137), .B2(n18942), .ZN(n18937) );
  AOI22_X1 U21970 ( .A1(n19138), .A2(n18944), .B1(n19139), .B2(n18965), .ZN(
        n18936) );
  OAI211_X1 U21971 ( .C1(n19142), .C2(n18947), .A(n18937), .B(n18936), .ZN(
        P3_U2928) );
  AOI22_X1 U21972 ( .A1(n19144), .A2(n18965), .B1(n19143), .B2(n18942), .ZN(
        n18939) );
  AOI22_X1 U21973 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18943), .B1(
        n19145), .B2(n18944), .ZN(n18938) );
  OAI211_X1 U21974 ( .C1(n19148), .C2(n18947), .A(n18939), .B(n18938), .ZN(
        P3_U2929) );
  AOI22_X1 U21975 ( .A1(n19151), .A2(n18944), .B1(n19149), .B2(n18942), .ZN(
        n18941) );
  AOI22_X1 U21976 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18943), .B1(
        n19150), .B2(n18965), .ZN(n18940) );
  OAI211_X1 U21977 ( .C1(n19154), .C2(n18947), .A(n18941), .B(n18940), .ZN(
        P3_U2930) );
  AOI22_X1 U21978 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18943), .B1(
        n19156), .B2(n18942), .ZN(n18946) );
  AOI22_X1 U21979 ( .A1(n19158), .A2(n18944), .B1(n19159), .B2(n18965), .ZN(
        n18945) );
  OAI211_X1 U21980 ( .C1(n19164), .C2(n18947), .A(n18946), .B(n18945), .ZN(
        P3_U2931) );
  NAND2_X1 U21981 ( .A1(n19174), .A2(n19016), .ZN(n18969) );
  NOR2_X1 U21982 ( .A1(n19010), .A2(n19032), .ZN(n18993) );
  NOR2_X1 U21983 ( .A1(n19225), .A2(n18993), .ZN(n18964) );
  AOI22_X1 U21984 ( .A1(n19110), .A2(n18964), .B1(n19111), .B2(n18988), .ZN(
        n18951) );
  OAI21_X1 U21985 ( .B1(n18948), .B2(n19084), .A(n18993), .ZN(n18949) );
  OAI211_X1 U21986 ( .C1(n19032), .C2(n19322), .A(n19087), .B(n18949), .ZN(
        n18966) );
  AOI22_X1 U21987 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18966), .B1(
        n19115), .B2(n18965), .ZN(n18950) );
  OAI211_X1 U21988 ( .C1(n19118), .C2(n18969), .A(n18951), .B(n18950), .ZN(
        P3_U2932) );
  AOI22_X1 U21989 ( .A1(n19120), .A2(n18965), .B1(n19119), .B2(n18964), .ZN(
        n18953) );
  AOI22_X1 U21990 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18966), .B1(
        n19121), .B2(n18988), .ZN(n18952) );
  OAI211_X1 U21991 ( .C1(n19124), .C2(n18969), .A(n18953), .B(n18952), .ZN(
        P3_U2933) );
  AOI22_X1 U21992 ( .A1(n19127), .A2(n18965), .B1(n19125), .B2(n18964), .ZN(
        n18955) );
  AOI22_X1 U21993 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18966), .B1(
        n19126), .B2(n18988), .ZN(n18954) );
  OAI211_X1 U21994 ( .C1(n19130), .C2(n18969), .A(n18955), .B(n18954), .ZN(
        P3_U2934) );
  AOI22_X1 U21995 ( .A1(n19132), .A2(n18988), .B1(n19131), .B2(n18964), .ZN(
        n18957) );
  AOI22_X1 U21996 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18966), .B1(
        n19133), .B2(n18965), .ZN(n18956) );
  OAI211_X1 U21997 ( .C1(n19136), .C2(n18969), .A(n18957), .B(n18956), .ZN(
        P3_U2935) );
  AOI22_X1 U21998 ( .A1(n19137), .A2(n18964), .B1(n19139), .B2(n18988), .ZN(
        n18959) );
  AOI22_X1 U21999 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18966), .B1(
        n19138), .B2(n18965), .ZN(n18958) );
  OAI211_X1 U22000 ( .C1(n19142), .C2(n18969), .A(n18959), .B(n18958), .ZN(
        P3_U2936) );
  AOI22_X1 U22001 ( .A1(n19143), .A2(n18964), .B1(n19145), .B2(n18965), .ZN(
        n18961) );
  AOI22_X1 U22002 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18966), .B1(
        n19144), .B2(n18988), .ZN(n18960) );
  OAI211_X1 U22003 ( .C1(n19148), .C2(n18969), .A(n18961), .B(n18960), .ZN(
        P3_U2937) );
  AOI22_X1 U22004 ( .A1(n19150), .A2(n18988), .B1(n19149), .B2(n18964), .ZN(
        n18963) );
  AOI22_X1 U22005 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18966), .B1(
        n19151), .B2(n18965), .ZN(n18962) );
  OAI211_X1 U22006 ( .C1(n19154), .C2(n18969), .A(n18963), .B(n18962), .ZN(
        P3_U2938) );
  AOI22_X1 U22007 ( .A1(n19159), .A2(n18988), .B1(n19156), .B2(n18964), .ZN(
        n18968) );
  AOI22_X1 U22008 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18966), .B1(
        n19158), .B2(n18965), .ZN(n18967) );
  OAI211_X1 U22009 ( .C1(n19164), .C2(n18969), .A(n18968), .B(n18967), .ZN(
        P3_U2939) );
  NAND2_X1 U22010 ( .A1(n18970), .A2(n19016), .ZN(n18992) );
  INV_X1 U22011 ( .A(n19016), .ZN(n18971) );
  NOR2_X1 U22012 ( .A1(n18971), .A2(n19059), .ZN(n18987) );
  AOI22_X1 U22013 ( .A1(n19110), .A2(n18987), .B1(n19111), .B2(n19010), .ZN(
        n18974) );
  AOI22_X1 U22014 ( .A1(n16992), .A2(n18972), .B1(n19016), .B2(n19061), .ZN(
        n18989) );
  AOI22_X1 U22015 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18989), .B1(
        n19115), .B2(n18988), .ZN(n18973) );
  OAI211_X1 U22016 ( .C1(n19118), .C2(n18992), .A(n18974), .B(n18973), .ZN(
        P3_U2940) );
  AOI22_X1 U22017 ( .A1(n19121), .A2(n19010), .B1(n19119), .B2(n18987), .ZN(
        n18976) );
  AOI22_X1 U22018 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18989), .B1(
        n19120), .B2(n18988), .ZN(n18975) );
  OAI211_X1 U22019 ( .C1(n19124), .C2(n18992), .A(n18976), .B(n18975), .ZN(
        P3_U2941) );
  AOI22_X1 U22020 ( .A1(n19126), .A2(n19010), .B1(n19125), .B2(n18987), .ZN(
        n18978) );
  AOI22_X1 U22021 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18989), .B1(
        n19127), .B2(n18988), .ZN(n18977) );
  OAI211_X1 U22022 ( .C1(n19130), .C2(n18992), .A(n18978), .B(n18977), .ZN(
        P3_U2942) );
  AOI22_X1 U22023 ( .A1(n19132), .A2(n19010), .B1(n19131), .B2(n18987), .ZN(
        n18980) );
  AOI22_X1 U22024 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18989), .B1(
        n19133), .B2(n18988), .ZN(n18979) );
  OAI211_X1 U22025 ( .C1(n19136), .C2(n18992), .A(n18980), .B(n18979), .ZN(
        P3_U2943) );
  AOI22_X1 U22026 ( .A1(n19137), .A2(n18987), .B1(n19139), .B2(n19010), .ZN(
        n18982) );
  AOI22_X1 U22027 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18989), .B1(
        n19138), .B2(n18988), .ZN(n18981) );
  OAI211_X1 U22028 ( .C1(n19142), .C2(n18992), .A(n18982), .B(n18981), .ZN(
        P3_U2944) );
  AOI22_X1 U22029 ( .A1(n19144), .A2(n19010), .B1(n19143), .B2(n18987), .ZN(
        n18984) );
  AOI22_X1 U22030 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18989), .B1(
        n19145), .B2(n18988), .ZN(n18983) );
  OAI211_X1 U22031 ( .C1(n19148), .C2(n18992), .A(n18984), .B(n18983), .ZN(
        P3_U2945) );
  AOI22_X1 U22032 ( .A1(n19150), .A2(n19010), .B1(n19149), .B2(n18987), .ZN(
        n18986) );
  AOI22_X1 U22033 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18989), .B1(
        n19151), .B2(n18988), .ZN(n18985) );
  OAI211_X1 U22034 ( .C1(n19154), .C2(n18992), .A(n18986), .B(n18985), .ZN(
        P3_U2946) );
  AOI22_X1 U22035 ( .A1(n19159), .A2(n19010), .B1(n19156), .B2(n18987), .ZN(
        n18991) );
  AOI22_X1 U22036 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18989), .B1(
        n19158), .B2(n18988), .ZN(n18990) );
  OAI211_X1 U22037 ( .C1(n19164), .C2(n18992), .A(n18991), .B(n18990), .ZN(
        P3_U2947) );
  NAND2_X1 U22038 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19016), .ZN(
        n19015) );
  INV_X1 U22039 ( .A(n19015), .ZN(n19063) );
  NAND2_X1 U22040 ( .A1(n21323), .A2(n19063), .ZN(n19014) );
  NOR2_X1 U22041 ( .A1(n19078), .A2(n19054), .ZN(n19037) );
  NOR2_X1 U22042 ( .A1(n19225), .A2(n19037), .ZN(n19009) );
  AOI22_X1 U22043 ( .A1(n19110), .A2(n19009), .B1(n19111), .B2(n19032), .ZN(
        n18996) );
  OAI21_X1 U22044 ( .B1(n18993), .B2(n19084), .A(n19037), .ZN(n18994) );
  OAI211_X1 U22045 ( .C1(n19078), .C2(n19322), .A(n19087), .B(n18994), .ZN(
        n19011) );
  AOI22_X1 U22046 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19011), .B1(
        n19115), .B2(n19010), .ZN(n18995) );
  OAI211_X1 U22047 ( .C1(n19118), .C2(n19014), .A(n18996), .B(n18995), .ZN(
        P3_U2948) );
  AOI22_X1 U22048 ( .A1(n19120), .A2(n19010), .B1(n19119), .B2(n19009), .ZN(
        n18998) );
  AOI22_X1 U22049 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19011), .B1(
        n19121), .B2(n19032), .ZN(n18997) );
  OAI211_X1 U22050 ( .C1(n19124), .C2(n19014), .A(n18998), .B(n18997), .ZN(
        P3_U2949) );
  AOI22_X1 U22051 ( .A1(n19126), .A2(n19032), .B1(n19125), .B2(n19009), .ZN(
        n19000) );
  AOI22_X1 U22052 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19011), .B1(
        n19127), .B2(n19010), .ZN(n18999) );
  OAI211_X1 U22053 ( .C1(n19130), .C2(n19014), .A(n19000), .B(n18999), .ZN(
        P3_U2950) );
  AOI22_X1 U22054 ( .A1(n19133), .A2(n19010), .B1(n19131), .B2(n19009), .ZN(
        n19002) );
  AOI22_X1 U22055 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19011), .B1(
        n19132), .B2(n19032), .ZN(n19001) );
  OAI211_X1 U22056 ( .C1(n19136), .C2(n19014), .A(n19002), .B(n19001), .ZN(
        P3_U2951) );
  AOI22_X1 U22057 ( .A1(n19138), .A2(n19010), .B1(n19137), .B2(n19009), .ZN(
        n19004) );
  AOI22_X1 U22058 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19011), .B1(
        n19139), .B2(n19032), .ZN(n19003) );
  OAI211_X1 U22059 ( .C1(n19142), .C2(n19014), .A(n19004), .B(n19003), .ZN(
        P3_U2952) );
  AOI22_X1 U22060 ( .A1(n19143), .A2(n19009), .B1(n19145), .B2(n19010), .ZN(
        n19006) );
  AOI22_X1 U22061 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19011), .B1(
        n19144), .B2(n19032), .ZN(n19005) );
  OAI211_X1 U22062 ( .C1(n19148), .C2(n19014), .A(n19006), .B(n19005), .ZN(
        P3_U2953) );
  AOI22_X1 U22063 ( .A1(n19151), .A2(n19010), .B1(n19149), .B2(n19009), .ZN(
        n19008) );
  AOI22_X1 U22064 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19011), .B1(
        n19150), .B2(n19032), .ZN(n19007) );
  OAI211_X1 U22065 ( .C1(n19154), .C2(n19014), .A(n19008), .B(n19007), .ZN(
        P3_U2954) );
  AOI22_X1 U22066 ( .A1(n19159), .A2(n19032), .B1(n19156), .B2(n19009), .ZN(
        n19013) );
  AOI22_X1 U22067 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19011), .B1(
        n19158), .B2(n19010), .ZN(n19012) );
  OAI211_X1 U22068 ( .C1(n19164), .C2(n19014), .A(n19013), .B(n19012), .ZN(
        P3_U2955) );
  NOR2_X2 U22069 ( .A1(n21323), .A2(n19015), .ZN(n19104) );
  NOR2_X1 U22070 ( .A1(n19225), .A2(n19015), .ZN(n19031) );
  AOI22_X1 U22071 ( .A1(n19110), .A2(n19031), .B1(n19111), .B2(n19054), .ZN(
        n19018) );
  AOI22_X1 U22072 ( .A1(n16992), .A2(n19016), .B1(n19063), .B2(n19112), .ZN(
        n19033) );
  AOI22_X1 U22073 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19033), .B1(
        n19115), .B2(n19032), .ZN(n19017) );
  OAI211_X1 U22074 ( .C1(n19118), .C2(n19036), .A(n19018), .B(n19017), .ZN(
        P3_U2956) );
  AOI22_X1 U22075 ( .A1(n19121), .A2(n19054), .B1(n19119), .B2(n19031), .ZN(
        n19020) );
  AOI22_X1 U22076 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19033), .B1(
        n19120), .B2(n19032), .ZN(n19019) );
  OAI211_X1 U22077 ( .C1(n19124), .C2(n19036), .A(n19020), .B(n19019), .ZN(
        P3_U2957) );
  AOI22_X1 U22078 ( .A1(n19126), .A2(n19054), .B1(n19125), .B2(n19031), .ZN(
        n19022) );
  AOI22_X1 U22079 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19033), .B1(
        n19127), .B2(n19032), .ZN(n19021) );
  OAI211_X1 U22080 ( .C1(n19130), .C2(n19036), .A(n19022), .B(n19021), .ZN(
        P3_U2958) );
  AOI22_X1 U22081 ( .A1(n19133), .A2(n19032), .B1(n19131), .B2(n19031), .ZN(
        n19024) );
  AOI22_X1 U22082 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19033), .B1(
        n19132), .B2(n19054), .ZN(n19023) );
  OAI211_X1 U22083 ( .C1(n19136), .C2(n19036), .A(n19024), .B(n19023), .ZN(
        P3_U2959) );
  AOI22_X1 U22084 ( .A1(n19137), .A2(n19031), .B1(n19139), .B2(n19054), .ZN(
        n19026) );
  AOI22_X1 U22085 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19033), .B1(
        n19138), .B2(n19032), .ZN(n19025) );
  OAI211_X1 U22086 ( .C1(n19142), .C2(n19036), .A(n19026), .B(n19025), .ZN(
        P3_U2960) );
  AOI22_X1 U22087 ( .A1(n19143), .A2(n19031), .B1(n19145), .B2(n19032), .ZN(
        n19028) );
  AOI22_X1 U22088 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19033), .B1(
        n19144), .B2(n19054), .ZN(n19027) );
  OAI211_X1 U22089 ( .C1(n19148), .C2(n19036), .A(n19028), .B(n19027), .ZN(
        P3_U2961) );
  AOI22_X1 U22090 ( .A1(n19151), .A2(n19032), .B1(n19149), .B2(n19031), .ZN(
        n19030) );
  AOI22_X1 U22091 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19033), .B1(
        n19150), .B2(n19054), .ZN(n19029) );
  OAI211_X1 U22092 ( .C1(n19154), .C2(n19036), .A(n19030), .B(n19029), .ZN(
        P3_U2962) );
  AOI22_X1 U22093 ( .A1(n19159), .A2(n19054), .B1(n19156), .B2(n19031), .ZN(
        n19035) );
  AOI22_X1 U22094 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19033), .B1(
        n19158), .B2(n19032), .ZN(n19034) );
  OAI211_X1 U22095 ( .C1(n19164), .C2(n19036), .A(n19035), .B(n19034), .ZN(
        P3_U2963) );
  NAND2_X1 U22096 ( .A1(n19174), .A2(n19062), .ZN(n19058) );
  AOI21_X1 U22097 ( .B1(n19058), .B2(n19036), .A(n19225), .ZN(n19053) );
  AOI22_X1 U22098 ( .A1(n19110), .A2(n19053), .B1(n19111), .B2(n19078), .ZN(
        n19040) );
  INV_X1 U22099 ( .A(n19058), .ZN(n19157) );
  AOI221_X1 U22100 ( .B1(n19037), .B2(n19036), .C1(n19084), .C2(n19036), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n19038) );
  OAI21_X1 U22101 ( .B1(n19157), .B2(n19038), .A(n19087), .ZN(n19055) );
  AOI22_X1 U22102 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19055), .B1(
        n19115), .B2(n19054), .ZN(n19039) );
  OAI211_X1 U22103 ( .C1(n19118), .C2(n19058), .A(n19040), .B(n19039), .ZN(
        P3_U2964) );
  AOI22_X1 U22104 ( .A1(n19120), .A2(n19054), .B1(n19119), .B2(n19053), .ZN(
        n19042) );
  AOI22_X1 U22105 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19055), .B1(
        n19121), .B2(n19078), .ZN(n19041) );
  OAI211_X1 U22106 ( .C1(n19124), .C2(n19058), .A(n19042), .B(n19041), .ZN(
        P3_U2965) );
  AOI22_X1 U22107 ( .A1(n19127), .A2(n19054), .B1(n19125), .B2(n19053), .ZN(
        n19044) );
  AOI22_X1 U22108 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19055), .B1(
        n19126), .B2(n19078), .ZN(n19043) );
  OAI211_X1 U22109 ( .C1(n19130), .C2(n19058), .A(n19044), .B(n19043), .ZN(
        P3_U2966) );
  AOI22_X1 U22110 ( .A1(n19133), .A2(n19054), .B1(n19131), .B2(n19053), .ZN(
        n19046) );
  AOI22_X1 U22111 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19055), .B1(
        n19132), .B2(n19078), .ZN(n19045) );
  OAI211_X1 U22112 ( .C1(n19136), .C2(n19058), .A(n19046), .B(n19045), .ZN(
        P3_U2967) );
  AOI22_X1 U22113 ( .A1(n19138), .A2(n19054), .B1(n19137), .B2(n19053), .ZN(
        n19048) );
  AOI22_X1 U22114 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19055), .B1(
        n19139), .B2(n19078), .ZN(n19047) );
  OAI211_X1 U22115 ( .C1(n19142), .C2(n19058), .A(n19048), .B(n19047), .ZN(
        P3_U2968) );
  AOI22_X1 U22116 ( .A1(n19143), .A2(n19053), .B1(n19145), .B2(n19054), .ZN(
        n19050) );
  AOI22_X1 U22117 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19055), .B1(
        n19144), .B2(n19078), .ZN(n19049) );
  OAI211_X1 U22118 ( .C1(n19148), .C2(n19058), .A(n19050), .B(n19049), .ZN(
        P3_U2969) );
  AOI22_X1 U22119 ( .A1(n19151), .A2(n19054), .B1(n19149), .B2(n19053), .ZN(
        n19052) );
  AOI22_X1 U22120 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19055), .B1(
        n19150), .B2(n19078), .ZN(n19051) );
  OAI211_X1 U22121 ( .C1(n19154), .C2(n19058), .A(n19052), .B(n19051), .ZN(
        P3_U2970) );
  AOI22_X1 U22122 ( .A1(n19158), .A2(n19054), .B1(n19156), .B2(n19053), .ZN(
        n19057) );
  AOI22_X1 U22123 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19055), .B1(
        n19159), .B2(n19078), .ZN(n19056) );
  OAI211_X1 U22124 ( .C1(n19164), .C2(n19058), .A(n19057), .B(n19056), .ZN(
        P3_U2971) );
  INV_X1 U22125 ( .A(n19062), .ZN(n19060) );
  NOR2_X1 U22126 ( .A1(n19060), .A2(n19059), .ZN(n19114) );
  AOI22_X1 U22127 ( .A1(n19110), .A2(n19114), .B1(n19111), .B2(n19104), .ZN(
        n19065) );
  AOI22_X1 U22128 ( .A1(n16992), .A2(n19063), .B1(n19062), .B2(n19061), .ZN(
        n19079) );
  AOI22_X1 U22129 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19079), .B1(
        n19115), .B2(n19078), .ZN(n19064) );
  OAI211_X1 U22130 ( .C1(n19082), .C2(n19118), .A(n19065), .B(n19064), .ZN(
        P3_U2972) );
  AOI22_X1 U22131 ( .A1(n19120), .A2(n19078), .B1(n19119), .B2(n19114), .ZN(
        n19067) );
  AOI22_X1 U22132 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19079), .B1(
        n19121), .B2(n19104), .ZN(n19066) );
  OAI211_X1 U22133 ( .C1(n19082), .C2(n19124), .A(n19067), .B(n19066), .ZN(
        P3_U2973) );
  AOI22_X1 U22134 ( .A1(n19127), .A2(n19078), .B1(n19125), .B2(n19114), .ZN(
        n19069) );
  AOI22_X1 U22135 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19079), .B1(
        n19126), .B2(n19104), .ZN(n19068) );
  OAI211_X1 U22136 ( .C1(n19082), .C2(n19130), .A(n19069), .B(n19068), .ZN(
        P3_U2974) );
  AOI22_X1 U22137 ( .A1(n19132), .A2(n19104), .B1(n19131), .B2(n19114), .ZN(
        n19071) );
  AOI22_X1 U22138 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19079), .B1(
        n19133), .B2(n19078), .ZN(n19070) );
  OAI211_X1 U22139 ( .C1(n19082), .C2(n19136), .A(n19071), .B(n19070), .ZN(
        P3_U2975) );
  AOI22_X1 U22140 ( .A1(n19137), .A2(n19114), .B1(n19139), .B2(n19104), .ZN(
        n19073) );
  AOI22_X1 U22141 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19079), .B1(
        n19138), .B2(n19078), .ZN(n19072) );
  OAI211_X1 U22142 ( .C1(n19082), .C2(n19142), .A(n19073), .B(n19072), .ZN(
        P3_U2976) );
  AOI22_X1 U22143 ( .A1(n19144), .A2(n19104), .B1(n19143), .B2(n19114), .ZN(
        n19075) );
  AOI22_X1 U22144 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19079), .B1(
        n19145), .B2(n19078), .ZN(n19074) );
  OAI211_X1 U22145 ( .C1(n19082), .C2(n19148), .A(n19075), .B(n19074), .ZN(
        P3_U2977) );
  AOI22_X1 U22146 ( .A1(n19151), .A2(n19078), .B1(n19149), .B2(n19114), .ZN(
        n19077) );
  AOI22_X1 U22147 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19079), .B1(
        n19150), .B2(n19104), .ZN(n19076) );
  OAI211_X1 U22148 ( .C1(n19082), .C2(n19154), .A(n19077), .B(n19076), .ZN(
        P3_U2978) );
  AOI22_X1 U22149 ( .A1(n19159), .A2(n19104), .B1(n19156), .B2(n19114), .ZN(
        n19081) );
  AOI22_X1 U22150 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19079), .B1(
        n19158), .B2(n19078), .ZN(n19080) );
  OAI211_X1 U22151 ( .C1(n19082), .C2(n19164), .A(n19081), .B(n19080), .ZN(
        P3_U2979) );
  NOR2_X1 U22152 ( .A1(n19225), .A2(n19083), .ZN(n19103) );
  AOI22_X1 U22153 ( .A1(n19110), .A2(n19103), .B1(n19111), .B2(n19157), .ZN(
        n19090) );
  NOR2_X1 U22154 ( .A1(n19157), .A2(n19104), .ZN(n19085) );
  OAI21_X1 U22155 ( .B1(n19085), .B2(n19084), .A(n19083), .ZN(n19086) );
  OAI211_X1 U22156 ( .C1(n19088), .C2(n19322), .A(n19087), .B(n19086), .ZN(
        n19105) );
  AOI22_X1 U22157 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19105), .B1(
        n19115), .B2(n19104), .ZN(n19089) );
  OAI211_X1 U22158 ( .C1(n19108), .C2(n19118), .A(n19090), .B(n19089), .ZN(
        P3_U2980) );
  AOI22_X1 U22159 ( .A1(n19121), .A2(n19157), .B1(n19119), .B2(n19103), .ZN(
        n19092) );
  AOI22_X1 U22160 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19105), .B1(
        n19120), .B2(n19104), .ZN(n19091) );
  OAI211_X1 U22161 ( .C1(n19108), .C2(n19124), .A(n19092), .B(n19091), .ZN(
        P3_U2981) );
  AOI22_X1 U22162 ( .A1(n19127), .A2(n19104), .B1(n19125), .B2(n19103), .ZN(
        n19094) );
  AOI22_X1 U22163 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19105), .B1(
        n19126), .B2(n19157), .ZN(n19093) );
  OAI211_X1 U22164 ( .C1(n19108), .C2(n19130), .A(n19094), .B(n19093), .ZN(
        P3_U2982) );
  AOI22_X1 U22165 ( .A1(n19132), .A2(n19157), .B1(n19131), .B2(n19103), .ZN(
        n19096) );
  AOI22_X1 U22166 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19105), .B1(
        n19133), .B2(n19104), .ZN(n19095) );
  OAI211_X1 U22167 ( .C1(n19108), .C2(n19136), .A(n19096), .B(n19095), .ZN(
        P3_U2983) );
  AOI22_X1 U22168 ( .A1(n19138), .A2(n19104), .B1(n19137), .B2(n19103), .ZN(
        n19098) );
  AOI22_X1 U22169 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19105), .B1(
        n19139), .B2(n19157), .ZN(n19097) );
  OAI211_X1 U22170 ( .C1(n19108), .C2(n19142), .A(n19098), .B(n19097), .ZN(
        P3_U2984) );
  AOI22_X1 U22171 ( .A1(n19144), .A2(n19157), .B1(n19143), .B2(n19103), .ZN(
        n19100) );
  AOI22_X1 U22172 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19105), .B1(
        n19145), .B2(n19104), .ZN(n19099) );
  OAI211_X1 U22173 ( .C1(n19108), .C2(n19148), .A(n19100), .B(n19099), .ZN(
        P3_U2985) );
  AOI22_X1 U22174 ( .A1(n19150), .A2(n19157), .B1(n19149), .B2(n19103), .ZN(
        n19102) );
  AOI22_X1 U22175 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19105), .B1(
        n19151), .B2(n19104), .ZN(n19101) );
  OAI211_X1 U22176 ( .C1(n19108), .C2(n19154), .A(n19102), .B(n19101), .ZN(
        P3_U2986) );
  AOI22_X1 U22177 ( .A1(n19158), .A2(n19104), .B1(n19156), .B2(n19103), .ZN(
        n19107) );
  AOI22_X1 U22178 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19105), .B1(
        n19159), .B2(n19157), .ZN(n19106) );
  OAI211_X1 U22179 ( .C1(n19108), .C2(n19164), .A(n19107), .B(n19106), .ZN(
        P3_U2987) );
  AND2_X1 U22180 ( .A1(n19109), .A2(n19113), .ZN(n19155) );
  AOI22_X1 U22181 ( .A1(n19160), .A2(n19111), .B1(n19110), .B2(n19155), .ZN(
        n19117) );
  AOI22_X1 U22182 ( .A1(n16992), .A2(n19114), .B1(n19113), .B2(n19112), .ZN(
        n19161) );
  AOI22_X1 U22183 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19161), .B1(
        n19115), .B2(n19157), .ZN(n19116) );
  OAI211_X1 U22184 ( .C1(n19165), .C2(n19118), .A(n19117), .B(n19116), .ZN(
        P3_U2988) );
  AOI22_X1 U22185 ( .A1(n19120), .A2(n19157), .B1(n19119), .B2(n19155), .ZN(
        n19123) );
  AOI22_X1 U22186 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19161), .B1(
        n19160), .B2(n19121), .ZN(n19122) );
  OAI211_X1 U22187 ( .C1(n19165), .C2(n19124), .A(n19123), .B(n19122), .ZN(
        P3_U2989) );
  AOI22_X1 U22188 ( .A1(n19160), .A2(n19126), .B1(n19125), .B2(n19155), .ZN(
        n19129) );
  AOI22_X1 U22189 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19161), .B1(
        n19127), .B2(n19157), .ZN(n19128) );
  OAI211_X1 U22190 ( .C1(n19165), .C2(n19130), .A(n19129), .B(n19128), .ZN(
        P3_U2990) );
  AOI22_X1 U22191 ( .A1(n19160), .A2(n19132), .B1(n19131), .B2(n19155), .ZN(
        n19135) );
  AOI22_X1 U22192 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19161), .B1(
        n19133), .B2(n19157), .ZN(n19134) );
  OAI211_X1 U22193 ( .C1(n19165), .C2(n19136), .A(n19135), .B(n19134), .ZN(
        P3_U2991) );
  AOI22_X1 U22194 ( .A1(n19138), .A2(n19157), .B1(n19137), .B2(n19155), .ZN(
        n19141) );
  AOI22_X1 U22195 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19161), .B1(
        n19160), .B2(n19139), .ZN(n19140) );
  OAI211_X1 U22196 ( .C1(n19165), .C2(n19142), .A(n19141), .B(n19140), .ZN(
        P3_U2992) );
  AOI22_X1 U22197 ( .A1(n19160), .A2(n19144), .B1(n19143), .B2(n19155), .ZN(
        n19147) );
  AOI22_X1 U22198 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19161), .B1(
        n19145), .B2(n19157), .ZN(n19146) );
  OAI211_X1 U22199 ( .C1(n19165), .C2(n19148), .A(n19147), .B(n19146), .ZN(
        P3_U2993) );
  AOI22_X1 U22200 ( .A1(n19160), .A2(n19150), .B1(n19149), .B2(n19155), .ZN(
        n19153) );
  AOI22_X1 U22201 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19161), .B1(
        n19151), .B2(n19157), .ZN(n19152) );
  OAI211_X1 U22202 ( .C1(n19165), .C2(n19154), .A(n19153), .B(n19152), .ZN(
        P3_U2994) );
  AOI22_X1 U22203 ( .A1(n19158), .A2(n19157), .B1(n19156), .B2(n19155), .ZN(
        n19163) );
  AOI22_X1 U22204 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19161), .B1(
        n19160), .B2(n19159), .ZN(n19162) );
  OAI211_X1 U22205 ( .C1(n19165), .C2(n19164), .A(n19163), .B(n19162), .ZN(
        P3_U2995) );
  NOR2_X1 U22206 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19208) );
  NAND2_X1 U22207 ( .A1(n19194), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n19168) );
  INV_X1 U22208 ( .A(n19194), .ZN(n19192) );
  NAND2_X1 U22209 ( .A1(n19166), .A2(n19192), .ZN(n19167) );
  INV_X1 U22210 ( .A(n19169), .ZN(n19173) );
  INV_X1 U22211 ( .A(n19171), .ZN(n19170) );
  NOR3_X1 U22212 ( .A1(n19170), .A2(n21323), .A3(n12171), .ZN(n19172) );
  OAI22_X1 U22213 ( .A1(n19173), .A2(n19172), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n19171), .ZN(n19175) );
  AOI222_X1 U22214 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19191), 
        .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n19176), .C1(n19191), 
        .C2(n19176), .ZN(n19207) );
  INV_X1 U22215 ( .A(n19177), .ZN(n19182) );
  NOR2_X1 U22216 ( .A1(n19179), .A2(n19178), .ZN(n19181) );
  OAI222_X1 U22217 ( .A1(n19185), .A2(n19184), .B1(n19183), .B2(n19182), .C1(
        n19181), .C2(n19180), .ZN(n19332) );
  NOR2_X1 U22218 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(P3_MORE_REG_SCAN_IN), .ZN(
        n19205) );
  AOI211_X1 U22219 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n19194), .A(
        n19187), .B(n19186), .ZN(n19203) );
  OAI21_X1 U22220 ( .B1(n19189), .B2(n19207), .A(n19188), .ZN(n19190) );
  INV_X1 U22221 ( .A(n19190), .ZN(n19201) );
  INV_X1 U22222 ( .A(n19191), .ZN(n19200) );
  NAND2_X1 U22223 ( .A1(n19193), .A2(n19192), .ZN(n19198) );
  NOR2_X1 U22224 ( .A1(n19195), .A2(n19194), .ZN(n19197) );
  MUX2_X1 U22225 ( .A(n19198), .B(n19197), .S(n19196), .Z(n19199) );
  OAI21_X1 U22226 ( .B1(n19201), .B2(n19200), .A(n19199), .ZN(n19202) );
  OAI211_X1 U22227 ( .C1(n19205), .C2(n19204), .A(n19203), .B(n19202), .ZN(
        n19206) );
  AOI211_X1 U22228 ( .C1(n19208), .C2(n19207), .A(n19332), .B(n19206), .ZN(
        n19221) );
  AOI22_X1 U22229 ( .A1(n19343), .A2(n18170), .B1(n19209), .B2(n19232), .ZN(
        n19210) );
  INV_X1 U22230 ( .A(n19210), .ZN(n19217) );
  OR2_X1 U22231 ( .A1(n19212), .A2(n19211), .ZN(n19213) );
  NAND3_X1 U22232 ( .A1(n19221), .A2(n19214), .A3(n19213), .ZN(n19321) );
  OAI21_X1 U22233 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n19222), .A(n19321), 
        .ZN(n19224) );
  NOR2_X1 U22234 ( .A1(n19215), .A2(n19224), .ZN(n19216) );
  MUX2_X1 U22235 ( .A(n19217), .B(n19216), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n19219) );
  OAI211_X1 U22236 ( .C1(n19221), .C2(n19220), .A(n19219), .B(n19218), .ZN(
        P3_U2996) );
  NOR2_X1 U22237 ( .A1(n19222), .A2(n19342), .ZN(n19227) );
  NOR4_X1 U22238 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n19338), .A3(n19223), 
        .A4(n19222), .ZN(n19230) );
  NOR4_X1 U22239 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n19225), .A3(n19338), 
        .A4(n19224), .ZN(n19226) );
  OR4_X1 U22240 ( .A1(n19228), .A2(n19227), .A3(n19230), .A4(n19226), .ZN(
        P3_U2997) );
  NOR3_X1 U22241 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .ZN(n19231) );
  NOR4_X1 U22242 ( .A1(n19232), .A2(n19231), .A3(n19230), .A4(n19229), .ZN(
        P3_U2998) );
  AND2_X1 U22243 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n19233), .ZN(
        P3_U2999) );
  AND2_X1 U22244 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n19233), .ZN(
        P3_U3000) );
  AND2_X1 U22245 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n19233), .ZN(
        P3_U3001) );
  AND2_X1 U22246 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n19233), .ZN(
        P3_U3002) );
  AND2_X1 U22247 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n19233), .ZN(
        P3_U3003) );
  AND2_X1 U22248 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n19233), .ZN(
        P3_U3004) );
  AND2_X1 U22249 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n19233), .ZN(
        P3_U3005) );
  AND2_X1 U22250 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n19233), .ZN(
        P3_U3006) );
  AND2_X1 U22251 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n19233), .ZN(
        P3_U3007) );
  AND2_X1 U22252 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n19233), .ZN(
        P3_U3008) );
  AND2_X1 U22253 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n19233), .ZN(
        P3_U3009) );
  AND2_X1 U22254 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n19233), .ZN(
        P3_U3010) );
  AND2_X1 U22255 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n19233), .ZN(
        P3_U3011) );
  AND2_X1 U22256 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n19233), .ZN(
        P3_U3012) );
  AND2_X1 U22257 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n19233), .ZN(
        P3_U3013) );
  AND2_X1 U22258 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n19233), .ZN(
        P3_U3014) );
  AND2_X1 U22259 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n19233), .ZN(
        P3_U3015) );
  AND2_X1 U22260 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n19233), .ZN(
        P3_U3016) );
  INV_X1 U22261 ( .A(P3_DATAWIDTH_REG_13__SCAN_IN), .ZN(n21334) );
  NOR2_X1 U22262 ( .A1(n21334), .A2(n19319), .ZN(P3_U3017) );
  AND2_X1 U22263 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n19233), .ZN(
        P3_U3018) );
  AND2_X1 U22264 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n19233), .ZN(
        P3_U3019) );
  AND2_X1 U22265 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n19233), .ZN(
        P3_U3020) );
  AND2_X1 U22266 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n19233), .ZN(P3_U3021) );
  AND2_X1 U22267 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n19233), .ZN(P3_U3022) );
  AND2_X1 U22268 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n19233), .ZN(P3_U3023) );
  AND2_X1 U22269 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n19233), .ZN(P3_U3024) );
  AND2_X1 U22270 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n19233), .ZN(P3_U3025) );
  AND2_X1 U22271 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n19233), .ZN(P3_U3026) );
  AND2_X1 U22272 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n19233), .ZN(P3_U3027) );
  AND2_X1 U22273 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n19233), .ZN(P3_U3028) );
  INV_X1 U22274 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19241) );
  AOI21_X1 U22275 ( .B1(HOLD), .B2(n19234), .A(n19241), .ZN(n19238) );
  AOI21_X1 U22276 ( .B1(n19343), .B2(P3_STATE_REG_1__SCAN_IN), .A(n19235), 
        .ZN(n19249) );
  INV_X1 U22277 ( .A(NA), .ZN(n21141) );
  OAI21_X1 U22278 ( .B1(n21141), .B2(n19236), .A(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n19248) );
  INV_X1 U22279 ( .A(n19248), .ZN(n19237) );
  OAI22_X1 U22280 ( .A1(n19261), .A2(n19238), .B1(n19249), .B2(n19237), .ZN(
        P3_U3029) );
  NAND3_X1 U22281 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(HOLD), .A3(n21319), .ZN(
        n19239) );
  OAI221_X1 U22282 ( .B1(n19241), .B2(HOLD), .C1(n19241), .C2(n19240), .A(
        n19239), .ZN(n19242) );
  AOI22_X1 U22283 ( .A1(n19343), .A2(P3_STATE_REG_1__SCAN_IN), .B1(
        P3_STATE_REG_0__SCAN_IN), .B2(n19242), .ZN(n19244) );
  NAND2_X1 U22284 ( .A1(n19244), .A2(n19243), .ZN(P3_U3030) );
  NAND2_X1 U22285 ( .A1(n19343), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19245) );
  OAI222_X1 U22286 ( .A1(n20199), .A2(n21319), .B1(P3_STATE_REG_1__SCAN_IN), 
        .B2(P3_REQUESTPENDING_REG_SCAN_IN), .C1(n19245), .C2(NA), .ZN(n19246)
         );
  OAI211_X1 U22287 ( .C1(P3_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P3_STATE_REG_0__SCAN_IN), .B(n19246), .ZN(n19247) );
  OAI21_X1 U22288 ( .B1(n19249), .B2(n19248), .A(n19247), .ZN(P3_U3031) );
  OAI222_X1 U22289 ( .A1(n19251), .A2(n19306), .B1(n19250), .B2(n19261), .C1(
        n19252), .C2(n19311), .ZN(P3_U3032) );
  OAI222_X1 U22290 ( .A1(n19311), .A2(n21313), .B1(n19253), .B2(n19308), .C1(
        n19252), .C2(n19306), .ZN(P3_U3033) );
  OAI222_X1 U22291 ( .A1(n19311), .A2(n19255), .B1(n19254), .B2(n19261), .C1(
        n21313), .C2(n19306), .ZN(P3_U3034) );
  OAI222_X1 U22292 ( .A1(n19311), .A2(n19257), .B1(n19256), .B2(n19261), .C1(
        n19255), .C2(n19306), .ZN(P3_U3035) );
  OAI222_X1 U22293 ( .A1(n19311), .A2(n13987), .B1(n19258), .B2(n19261), .C1(
        n19257), .C2(n19306), .ZN(P3_U3036) );
  OAI222_X1 U22294 ( .A1(n19311), .A2(n19260), .B1(n19259), .B2(n19261), .C1(
        n13987), .C2(n19306), .ZN(P3_U3037) );
  OAI222_X1 U22295 ( .A1(n19311), .A2(n19264), .B1(n19262), .B2(n19261), .C1(
        n19260), .C2(n19306), .ZN(P3_U3038) );
  OAI222_X1 U22296 ( .A1(n19264), .A2(n19306), .B1(n19263), .B2(n19261), .C1(
        n19265), .C2(n19311), .ZN(P3_U3039) );
  OAI222_X1 U22297 ( .A1(n19311), .A2(n19267), .B1(n19266), .B2(n19261), .C1(
        n19265), .C2(n19306), .ZN(P3_U3040) );
  OAI222_X1 U22298 ( .A1(n19311), .A2(n19269), .B1(n19268), .B2(n19261), .C1(
        n19267), .C2(n19306), .ZN(P3_U3041) );
  OAI222_X1 U22299 ( .A1(n19311), .A2(n19271), .B1(n19270), .B2(n19261), .C1(
        n19269), .C2(n19306), .ZN(P3_U3042) );
  OAI222_X1 U22300 ( .A1(n19311), .A2(n19273), .B1(n19272), .B2(n19261), .C1(
        n19271), .C2(n19306), .ZN(P3_U3043) );
  OAI222_X1 U22301 ( .A1(n19311), .A2(n19275), .B1(n19274), .B2(n19261), .C1(
        n19273), .C2(n19306), .ZN(P3_U3044) );
  OAI222_X1 U22302 ( .A1(n19311), .A2(n19277), .B1(n19276), .B2(n19261), .C1(
        n19275), .C2(n19306), .ZN(P3_U3045) );
  OAI222_X1 U22303 ( .A1(n19311), .A2(n19279), .B1(n19278), .B2(n19261), .C1(
        n19277), .C2(n19306), .ZN(P3_U3046) );
  INV_X1 U22304 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n19282) );
  OAI222_X1 U22305 ( .A1(n19311), .A2(n19282), .B1(n19280), .B2(n19308), .C1(
        n19279), .C2(n19306), .ZN(P3_U3047) );
  OAI222_X1 U22306 ( .A1(n19282), .A2(n19306), .B1(n19281), .B2(n19308), .C1(
        n19283), .C2(n19311), .ZN(P3_U3048) );
  OAI222_X1 U22307 ( .A1(n19311), .A2(n19285), .B1(n19284), .B2(n19308), .C1(
        n19283), .C2(n19306), .ZN(P3_U3049) );
  OAI222_X1 U22308 ( .A1(n19285), .A2(n19306), .B1(n21368), .B2(n19308), .C1(
        n19286), .C2(n19311), .ZN(P3_U3050) );
  OAI222_X1 U22309 ( .A1(n19311), .A2(n19289), .B1(n19287), .B2(n19308), .C1(
        n19286), .C2(n19306), .ZN(P3_U3051) );
  OAI222_X1 U22310 ( .A1(n19289), .A2(n19306), .B1(n19288), .B2(n19308), .C1(
        n19290), .C2(n19311), .ZN(P3_U3052) );
  OAI222_X1 U22311 ( .A1(n19311), .A2(n19293), .B1(n19291), .B2(n19308), .C1(
        n19290), .C2(n19306), .ZN(P3_U3053) );
  OAI222_X1 U22312 ( .A1(n19293), .A2(n19306), .B1(n19292), .B2(n19308), .C1(
        n19294), .C2(n19311), .ZN(P3_U3054) );
  OAI222_X1 U22313 ( .A1(n19311), .A2(n19296), .B1(n19295), .B2(n19308), .C1(
        n19294), .C2(n19306), .ZN(P3_U3055) );
  OAI222_X1 U22314 ( .A1(n19311), .A2(n19298), .B1(n19297), .B2(n19308), .C1(
        n19296), .C2(n19306), .ZN(P3_U3056) );
  OAI222_X1 U22315 ( .A1(n19311), .A2(n19301), .B1(n19299), .B2(n19308), .C1(
        n19298), .C2(n19306), .ZN(P3_U3057) );
  INV_X1 U22316 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n19302) );
  OAI222_X1 U22317 ( .A1(n19306), .A2(n19301), .B1(n19300), .B2(n19308), .C1(
        n19302), .C2(n19311), .ZN(P3_U3058) );
  OAI222_X1 U22318 ( .A1(n19311), .A2(n19304), .B1(n19303), .B2(n19308), .C1(
        n19302), .C2(n19306), .ZN(P3_U3059) );
  OAI222_X1 U22319 ( .A1(n19311), .A2(n19307), .B1(n19305), .B2(n19308), .C1(
        n19304), .C2(n19306), .ZN(P3_U3060) );
  OAI222_X1 U22320 ( .A1(n19311), .A2(n19310), .B1(n19309), .B2(n19308), .C1(
        n19307), .C2(n19306), .ZN(P3_U3061) );
  OAI22_X1 U22321 ( .A1(n19347), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n19261), .ZN(n19312) );
  INV_X1 U22322 ( .A(n19312), .ZN(P3_U3274) );
  OAI22_X1 U22323 ( .A1(n19347), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n19261), .ZN(n19313) );
  INV_X1 U22324 ( .A(n19313), .ZN(P3_U3275) );
  OAI22_X1 U22325 ( .A1(n19347), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n19261), .ZN(n19314) );
  INV_X1 U22326 ( .A(n19314), .ZN(P3_U3276) );
  OAI22_X1 U22327 ( .A1(n19347), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n19261), .ZN(n19315) );
  INV_X1 U22328 ( .A(n19315), .ZN(P3_U3277) );
  OAI21_X1 U22329 ( .B1(n19319), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n19317), 
        .ZN(n19316) );
  INV_X1 U22330 ( .A(n19316), .ZN(P3_U3280) );
  OAI21_X1 U22331 ( .B1(n19319), .B2(n19318), .A(n19317), .ZN(P3_U3281) );
  OAI221_X1 U22332 ( .B1(n19322), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n19322), 
        .C2(n19321), .A(n19320), .ZN(P3_U3282) );
  AOI211_X1 U22333 ( .C1(P3_REIP_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_REIP_REG_1__SCAN_IN), .B(
        P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19323) );
  AOI21_X1 U22334 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n19323), .ZN(n19325) );
  INV_X1 U22335 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19324) );
  AOI22_X1 U22336 ( .A1(n19329), .A2(n19325), .B1(n19324), .B2(n19326), .ZN(
        P3_U3292) );
  NOR2_X1 U22337 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .ZN(n19328) );
  INV_X1 U22338 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19327) );
  AOI22_X1 U22339 ( .A1(n19329), .A2(n19328), .B1(n19327), .B2(n19326), .ZN(
        P3_U3293) );
  INV_X1 U22340 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n19352) );
  OAI22_X1 U22341 ( .A1(n19347), .A2(n19352), .B1(P3_W_R_N_REG_SCAN_IN), .B2(
        n19261), .ZN(n19330) );
  INV_X1 U22342 ( .A(n19330), .ZN(P3_U3294) );
  MUX2_X1 U22343 ( .A(P3_MORE_REG_SCAN_IN), .B(n19332), .S(n19331), .Z(
        P3_U3295) );
  OAI21_X1 U22344 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n19335), .A(n19334), 
        .ZN(n19336) );
  AOI211_X1 U22345 ( .C1(n9771), .C2(n19336), .A(n19343), .B(n19349), .ZN(
        n19339) );
  OAI21_X1 U22346 ( .B1(n19339), .B2(n19338), .A(n19337), .ZN(n19346) );
  OAI22_X1 U22347 ( .A1(n19343), .A2(n19342), .B1(n19341), .B2(n19340), .ZN(
        n19344) );
  NOR2_X1 U22348 ( .A1(n19351), .A2(n19344), .ZN(n19345) );
  MUX2_X1 U22349 ( .A(n19346), .B(P3_REQUESTPENDING_REG_SCAN_IN), .S(n19345), 
        .Z(P3_U3296) );
  OAI22_X1 U22350 ( .A1(n19347), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n19261), .ZN(n19348) );
  INV_X1 U22351 ( .A(n19348), .ZN(P3_U3297) );
  AOI21_X1 U22352 ( .B1(n19350), .B2(n19349), .A(n19351), .ZN(n19355) );
  AOI22_X1 U22353 ( .A1(n19355), .A2(n19352), .B1(n19351), .B2(n9771), .ZN(
        P3_U3298) );
  INV_X1 U22354 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n19354) );
  AOI21_X1 U22355 ( .B1(n19355), .B2(n19354), .A(n19353), .ZN(P3_U3299) );
  AOI21_X1 U22356 ( .B1(n19412), .B2(P2_MEMORYFETCH_REG_SCAN_IN), .A(n19356), 
        .ZN(n19357) );
  INV_X1 U22357 ( .A(n19357), .ZN(P2_U2814) );
  NAND2_X1 U22358 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20208), .ZN(n20200) );
  NAND2_X1 U22359 ( .A1(n20195), .A2(n20190), .ZN(n20196) );
  OAI21_X1 U22360 ( .B1(n20195), .B2(n20200), .A(n20196), .ZN(n20267) );
  AOI21_X1 U22361 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n20267), .ZN(n19358) );
  INV_X1 U22362 ( .A(n19358), .ZN(P2_U2815) );
  INV_X1 U22363 ( .A(n20202), .ZN(n19360) );
  AOI22_X1 U22364 ( .A1(P2_D_C_N_REG_SCAN_IN), .A2(n20326), .B1(n19360), .B2(
        n20195), .ZN(n19359) );
  OAI21_X1 U22365 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(n20326), .A(n19359), 
        .ZN(P2_U2817) );
  OAI21_X1 U22366 ( .B1(n19360), .B2(BS16), .A(n20267), .ZN(n20265) );
  OAI21_X1 U22367 ( .B1(n20267), .B2(n20272), .A(n20265), .ZN(P2_U2818) );
  NOR4_X1 U22368 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19370) );
  NOR4_X1 U22369 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19369) );
  INV_X1 U22370 ( .A(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n21292) );
  INV_X1 U22371 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20266) );
  NOR4_X1 U22372 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19361) );
  OAI21_X1 U22373 ( .B1(n21292), .B2(n20266), .A(n19361), .ZN(n19367) );
  NOR4_X1 U22374 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19365) );
  NOR4_X1 U22375 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19364) );
  NOR4_X1 U22376 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19363) );
  NOR4_X1 U22377 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19362) );
  NAND4_X1 U22378 ( .A1(n19365), .A2(n19364), .A3(n19363), .A4(n19362), .ZN(
        n19366) );
  NOR4_X1 U22379 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_3__SCAN_IN), .A3(n19367), .A4(n19366), .ZN(n19368) );
  NAND3_X1 U22380 ( .A1(n19370), .A2(n19369), .A3(n19368), .ZN(n19372) );
  NOR2_X1 U22381 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19372), .ZN(n19374) );
  INV_X1 U22382 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19371) );
  AOI22_X1 U22383 ( .A1(n19374), .A2(n19375), .B1(n19372), .B2(n19371), .ZN(
        P2_U2820) );
  INV_X1 U22384 ( .A(n19372), .ZN(n19381) );
  NOR2_X1 U22385 ( .A1(n19381), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19373)
         );
  NAND4_X1 U22386 ( .A1(n19381), .A2(n19375), .A3(n21292), .A4(n20266), .ZN(
        n19379) );
  OAI21_X1 U22387 ( .B1(n19374), .B2(n19373), .A(n19379), .ZN(P2_U2821) );
  NAND2_X1 U22388 ( .A1(n19374), .A2(n20266), .ZN(n19378) );
  OAI21_X1 U22389 ( .B1(n19375), .B2(n10958), .A(n19381), .ZN(n19376) );
  OAI21_X1 U22390 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19381), .A(n19376), 
        .ZN(n19377) );
  OAI221_X1 U22391 ( .B1(n19378), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19378), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19377), .ZN(P2_U2822) );
  INV_X1 U22392 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19380) );
  OAI211_X1 U22393 ( .C1(n19381), .C2(n19380), .A(n19379), .B(n19378), .ZN(
        P2_U2823) );
  INV_X1 U22394 ( .A(n19382), .ZN(n19385) );
  INV_X1 U22395 ( .A(n19383), .ZN(n19432) );
  AOI22_X1 U22396 ( .A1(n19385), .A2(n19413), .B1(n19432), .B2(n19384), .ZN(
        n19402) );
  AOI211_X1 U22397 ( .C1(n19399), .C2(n19388), .A(n19387), .B(n19386), .ZN(
        n19398) );
  OAI22_X1 U22398 ( .A1(n19392), .A2(n19391), .B1(n19390), .B2(n19389), .ZN(
        n19393) );
  NOR2_X1 U22399 ( .A1(n19571), .A2(n19393), .ZN(n19395) );
  NAND2_X1 U22400 ( .A1(n19410), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n19394) );
  OAI211_X1 U22401 ( .C1(n19396), .C2(n19405), .A(n19395), .B(n19394), .ZN(
        n19397) );
  AOI211_X1 U22402 ( .C1(n19400), .C2(n19399), .A(n19398), .B(n19397), .ZN(
        n19401) );
  NAND2_X1 U22403 ( .A1(n19402), .A2(n19401), .ZN(P2_U2840) );
  AOI22_X1 U22404 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19404), .B1(
        P2_EBX_REG_4__SCAN_IN), .B2(n19403), .ZN(n19424) );
  OAI22_X1 U22405 ( .A1(n19408), .A2(n19407), .B1(n19406), .B2(n19405), .ZN(
        n19409) );
  AOI211_X1 U22406 ( .C1(P2_REIP_REG_4__SCAN_IN), .C2(n19410), .A(n19571), .B(
        n19409), .ZN(n19423) );
  INV_X1 U22407 ( .A(n19411), .ZN(n19452) );
  INV_X1 U22408 ( .A(n19412), .ZN(n19414) );
  AOI22_X1 U22409 ( .A1(n19452), .A2(n19414), .B1(n19413), .B2(n19425), .ZN(
        n19422) );
  INV_X1 U22410 ( .A(n19581), .ZN(n19420) );
  NOR2_X1 U22411 ( .A1(n19416), .A2(n19415), .ZN(n19419) );
  AOI21_X1 U22412 ( .B1(n19419), .B2(n19420), .A(n19417), .ZN(n19418) );
  OAI21_X1 U22413 ( .B1(n19420), .B2(n19419), .A(n19418), .ZN(n19421) );
  NAND4_X1 U22414 ( .A1(n19424), .A2(n19423), .A3(n19422), .A4(n19421), .ZN(
        P2_U2851) );
  AOI22_X1 U22415 ( .A1(n19452), .A2(n19426), .B1(n19429), .B2(n19425), .ZN(
        n19427) );
  OAI21_X1 U22416 ( .B1(n19429), .B2(n19428), .A(n19427), .ZN(P2_U2883) );
  AOI22_X1 U22417 ( .A1(n19431), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n19430), .ZN(n19570) );
  AOI22_X1 U22418 ( .A1(n19432), .A2(n19451), .B1(P2_EAX_REG_15__SCAN_IN), 
        .B2(n19476), .ZN(n19433) );
  OAI21_X1 U22419 ( .B1(n19485), .B2(n19570), .A(n19433), .ZN(P2_U2904) );
  AOI22_X1 U22420 ( .A1(n19436), .A2(n19451), .B1(n19435), .B2(n19434), .ZN(
        n19437) );
  OAI21_X1 U22421 ( .B1(n19445), .B2(n19438), .A(n19437), .ZN(P2_U2908) );
  INV_X1 U22422 ( .A(n19439), .ZN(n19440) );
  OAI22_X1 U22423 ( .A1(n19442), .A2(n19441), .B1(n19440), .B2(n19485), .ZN(
        n19443) );
  INV_X1 U22424 ( .A(n19443), .ZN(n19444) );
  OAI21_X1 U22425 ( .B1(n19445), .B2(n19503), .A(n19444), .ZN(P2_U2910) );
  INV_X1 U22426 ( .A(n19446), .ZN(n19447) );
  AOI22_X1 U22427 ( .A1(n19447), .A2(n19451), .B1(P2_EAX_REG_6__SCAN_IN), .B2(
        n19476), .ZN(n19448) );
  OAI21_X1 U22428 ( .B1(n19553), .B2(n19485), .A(n19448), .ZN(P2_U2913) );
  INV_X1 U22429 ( .A(n19449), .ZN(n19450) );
  AOI22_X1 U22430 ( .A1(n19451), .A2(n19450), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n19476), .ZN(n19455) );
  NAND3_X1 U22431 ( .A1(n19453), .A2(n19452), .A3(n19479), .ZN(n19454) );
  OAI211_X1 U22432 ( .C1(n19551), .C2(n19485), .A(n19455), .B(n19454), .ZN(
        P2_U2914) );
  AOI22_X1 U22433 ( .A1(n19477), .A2(n20278), .B1(n19476), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n19461) );
  AOI21_X1 U22434 ( .B1(n19458), .B2(n19457), .A(n19456), .ZN(n19459) );
  OR2_X1 U22435 ( .A1(n19459), .A2(n19472), .ZN(n19460) );
  OAI211_X1 U22436 ( .C1(n19547), .C2(n19485), .A(n19461), .B(n19460), .ZN(
        P2_U2916) );
  AOI22_X1 U22437 ( .A1(n19477), .A2(n19462), .B1(n19476), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n19468) );
  AOI21_X1 U22438 ( .B1(n19465), .B2(n19464), .A(n19463), .ZN(n19466) );
  OR2_X1 U22439 ( .A1(n19466), .A2(n19472), .ZN(n19467) );
  OAI211_X1 U22440 ( .C1(n19545), .C2(n19485), .A(n19468), .B(n19467), .ZN(
        P2_U2917) );
  AOI22_X1 U22441 ( .A1(n19477), .A2(n19469), .B1(n19476), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n19475) );
  AOI21_X1 U22442 ( .B1(n19478), .B2(n19471), .A(n19470), .ZN(n19473) );
  OR2_X1 U22443 ( .A1(n19473), .A2(n19472), .ZN(n19474) );
  OAI211_X1 U22444 ( .C1(n19543), .C2(n19485), .A(n19475), .B(n19474), .ZN(
        P2_U2918) );
  AOI22_X1 U22445 ( .A1(n19477), .A2(n19481), .B1(n19476), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n19484) );
  INV_X1 U22446 ( .A(n19478), .ZN(n19480) );
  OAI211_X1 U22447 ( .C1(n19482), .C2(n19481), .A(n19480), .B(n19479), .ZN(
        n19483) );
  OAI211_X1 U22448 ( .C1(n19541), .C2(n19485), .A(n19484), .B(n19483), .ZN(
        P2_U2919) );
  NOR2_X1 U22449 ( .A1(n19492), .A2(n19486), .ZN(P2_U2920) );
  AOI22_X1 U22450 ( .A1(n19489), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n19520), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n19487) );
  OAI21_X1 U22451 ( .B1(n19492), .B2(n19488), .A(n19487), .ZN(P2_U2921) );
  AOI22_X1 U22452 ( .A1(n19489), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n19520), 
        .B2(P2_UWORD_REG_13__SCAN_IN), .ZN(n19490) );
  OAI21_X1 U22453 ( .B1(n19492), .B2(n19491), .A(n19490), .ZN(P2_U2922) );
  INV_X1 U22454 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19494) );
  AOI22_X1 U22455 ( .A1(n19521), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n19520), 
        .B2(P2_LWORD_REG_15__SCAN_IN), .ZN(n19493) );
  OAI21_X1 U22456 ( .B1(n19494), .B2(n19523), .A(n19493), .ZN(P2_U2936) );
  INV_X1 U22457 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19496) );
  AOI22_X1 U22458 ( .A1(n19521), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n19520), 
        .B2(P2_LWORD_REG_14__SCAN_IN), .ZN(n19495) );
  OAI21_X1 U22459 ( .B1(n19496), .B2(n19523), .A(n19495), .ZN(P2_U2937) );
  INV_X1 U22460 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19498) );
  AOI22_X1 U22461 ( .A1(n19521), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n19520), 
        .B2(P2_LWORD_REG_13__SCAN_IN), .ZN(n19497) );
  OAI21_X1 U22462 ( .B1(n19498), .B2(n19523), .A(n19497), .ZN(P2_U2938) );
  AOI22_X1 U22463 ( .A1(n19521), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n19520), 
        .B2(P2_LWORD_REG_12__SCAN_IN), .ZN(n19499) );
  OAI21_X1 U22464 ( .B1(n19500), .B2(n19523), .A(n19499), .ZN(P2_U2939) );
  AOI22_X1 U22465 ( .A1(n19521), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n19520), 
        .B2(P2_LWORD_REG_10__SCAN_IN), .ZN(n19501) );
  OAI21_X1 U22466 ( .B1(n21366), .B2(n19523), .A(n19501), .ZN(P2_U2941) );
  AOI22_X1 U22467 ( .A1(n19521), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n19520), 
        .B2(P2_LWORD_REG_9__SCAN_IN), .ZN(n19502) );
  OAI21_X1 U22468 ( .B1(n19503), .B2(n19523), .A(n19502), .ZN(P2_U2942) );
  AOI22_X1 U22469 ( .A1(n19521), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n19520), 
        .B2(P2_LWORD_REG_8__SCAN_IN), .ZN(n19504) );
  OAI21_X1 U22470 ( .B1(n19505), .B2(n19523), .A(n19504), .ZN(P2_U2943) );
  AOI22_X1 U22471 ( .A1(n19521), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n19520), 
        .B2(P2_LWORD_REG_7__SCAN_IN), .ZN(n19506) );
  OAI21_X1 U22472 ( .B1(n19507), .B2(n19523), .A(n19506), .ZN(P2_U2944) );
  INV_X1 U22473 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19509) );
  AOI22_X1 U22474 ( .A1(n19521), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n19520), 
        .B2(P2_LWORD_REG_6__SCAN_IN), .ZN(n19508) );
  OAI21_X1 U22475 ( .B1(n19509), .B2(n19523), .A(n19508), .ZN(P2_U2945) );
  INV_X1 U22476 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19511) );
  AOI22_X1 U22477 ( .A1(n19521), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n19520), 
        .B2(P2_LWORD_REG_5__SCAN_IN), .ZN(n19510) );
  OAI21_X1 U22478 ( .B1(n19511), .B2(n19523), .A(n19510), .ZN(P2_U2946) );
  AOI22_X1 U22479 ( .A1(n19521), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n19520), 
        .B2(P2_LWORD_REG_4__SCAN_IN), .ZN(n19512) );
  OAI21_X1 U22480 ( .B1(n19513), .B2(n19523), .A(n19512), .ZN(P2_U2947) );
  AOI22_X1 U22481 ( .A1(n19521), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n19520), 
        .B2(P2_LWORD_REG_3__SCAN_IN), .ZN(n19514) );
  OAI21_X1 U22482 ( .B1(n19515), .B2(n19523), .A(n19514), .ZN(P2_U2948) );
  INV_X1 U22483 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19517) );
  AOI22_X1 U22484 ( .A1(n19521), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n19520), 
        .B2(P2_LWORD_REG_2__SCAN_IN), .ZN(n19516) );
  OAI21_X1 U22485 ( .B1(n19517), .B2(n19523), .A(n19516), .ZN(P2_U2949) );
  INV_X1 U22486 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19519) );
  AOI22_X1 U22487 ( .A1(n19521), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(n19520), 
        .B2(P2_LWORD_REG_1__SCAN_IN), .ZN(n19518) );
  OAI21_X1 U22488 ( .B1(n19519), .B2(n19523), .A(n19518), .ZN(P2_U2950) );
  AOI22_X1 U22489 ( .A1(n19521), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(n19520), 
        .B2(P2_LWORD_REG_0__SCAN_IN), .ZN(n19522) );
  OAI21_X1 U22490 ( .B1(n10475), .B2(n19523), .A(n19522), .ZN(P2_U2951) );
  AOI22_X1 U22491 ( .A1(n19567), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_16__SCAN_IN), .B2(n19566), .ZN(n19524) );
  OAI21_X1 U22492 ( .B1(n19541), .B2(n19569), .A(n19524), .ZN(P2_U2952) );
  AOI22_X1 U22493 ( .A1(n19567), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(
        P2_EAX_REG_17__SCAN_IN), .B2(n19566), .ZN(n19525) );
  OAI21_X1 U22494 ( .B1(n19543), .B2(n19569), .A(n19525), .ZN(P2_U2953) );
  AOI22_X1 U22495 ( .A1(n10400), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_18__SCAN_IN), .B2(n19566), .ZN(n19526) );
  OAI21_X1 U22496 ( .B1(n19545), .B2(n19569), .A(n19526), .ZN(P2_U2954) );
  AOI22_X1 U22497 ( .A1(n10400), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_19__SCAN_IN), .B2(n19566), .ZN(n19527) );
  OAI21_X1 U22498 ( .B1(n19547), .B2(n19569), .A(n19527), .ZN(P2_U2955) );
  AOI22_X1 U22499 ( .A1(n10400), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n19566), .ZN(n19528) );
  OAI21_X1 U22500 ( .B1(n19549), .B2(n19569), .A(n19528), .ZN(P2_U2956) );
  AOI22_X1 U22501 ( .A1(n10400), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_21__SCAN_IN), .B2(n19566), .ZN(n19529) );
  OAI21_X1 U22502 ( .B1(n19551), .B2(n19569), .A(n19529), .ZN(P2_U2957) );
  AOI22_X1 U22503 ( .A1(n10400), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n19566), .ZN(n19530) );
  OAI21_X1 U22504 ( .B1(n19553), .B2(n19569), .A(n19530), .ZN(P2_U2958) );
  AOI22_X1 U22505 ( .A1(n10400), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(
        P2_EAX_REG_23__SCAN_IN), .B2(n19566), .ZN(n19531) );
  OAI21_X1 U22506 ( .B1(n19555), .B2(n19569), .A(n19531), .ZN(P2_U2959) );
  AOI22_X1 U22507 ( .A1(n10400), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_24__SCAN_IN), .B2(n19566), .ZN(n19532) );
  OAI21_X1 U22508 ( .B1(n19557), .B2(n19569), .A(n19532), .ZN(P2_U2960) );
  AOI22_X1 U22509 ( .A1(n10400), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(
        P2_EAX_REG_26__SCAN_IN), .B2(n19566), .ZN(n19533) );
  OAI21_X1 U22510 ( .B1(n19559), .B2(n19569), .A(n19533), .ZN(P2_U2962) );
  AOI22_X1 U22511 ( .A1(n10400), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_28__SCAN_IN), .B2(n19566), .ZN(n19534) );
  OAI21_X1 U22512 ( .B1(n19561), .B2(n19569), .A(n19534), .ZN(P2_U2964) );
  AOI22_X1 U22513 ( .A1(n19567), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n19566), .ZN(n19536) );
  NAND2_X1 U22514 ( .A1(n19538), .A2(n19535), .ZN(n19562) );
  NAND2_X1 U22515 ( .A1(n19536), .A2(n19562), .ZN(P2_U2965) );
  AOI22_X1 U22516 ( .A1(n10400), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_30__SCAN_IN), .B2(n19566), .ZN(n19539) );
  NAND2_X1 U22517 ( .A1(n19538), .A2(n19537), .ZN(n19564) );
  NAND2_X1 U22518 ( .A1(n19539), .A2(n19564), .ZN(P2_U2966) );
  AOI22_X1 U22519 ( .A1(n10400), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_0__SCAN_IN), .B2(n19566), .ZN(n19540) );
  OAI21_X1 U22520 ( .B1(n19541), .B2(n19569), .A(n19540), .ZN(P2_U2967) );
  AOI22_X1 U22521 ( .A1(n10400), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(
        P2_EAX_REG_1__SCAN_IN), .B2(n19566), .ZN(n19542) );
  OAI21_X1 U22522 ( .B1(n19543), .B2(n19569), .A(n19542), .ZN(P2_U2968) );
  AOI22_X1 U22523 ( .A1(n10400), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_2__SCAN_IN), .B2(n19566), .ZN(n19544) );
  OAI21_X1 U22524 ( .B1(n19545), .B2(n19569), .A(n19544), .ZN(P2_U2969) );
  AOI22_X1 U22525 ( .A1(n10400), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_3__SCAN_IN), .B2(n19566), .ZN(n19546) );
  OAI21_X1 U22526 ( .B1(n19547), .B2(n19569), .A(n19546), .ZN(P2_U2970) );
  AOI22_X1 U22527 ( .A1(n19567), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_4__SCAN_IN), .B2(n19566), .ZN(n19548) );
  OAI21_X1 U22528 ( .B1(n19549), .B2(n19569), .A(n19548), .ZN(P2_U2971) );
  AOI22_X1 U22529 ( .A1(n19567), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_5__SCAN_IN), .B2(n19566), .ZN(n19550) );
  OAI21_X1 U22530 ( .B1(n19551), .B2(n19569), .A(n19550), .ZN(P2_U2972) );
  AOI22_X1 U22531 ( .A1(n19567), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_6__SCAN_IN), .B2(n19566), .ZN(n19552) );
  OAI21_X1 U22532 ( .B1(n19553), .B2(n19569), .A(n19552), .ZN(P2_U2973) );
  AOI22_X1 U22533 ( .A1(n19567), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(
        P2_EAX_REG_7__SCAN_IN), .B2(n19566), .ZN(n19554) );
  OAI21_X1 U22534 ( .B1(n19555), .B2(n19569), .A(n19554), .ZN(P2_U2974) );
  AOI22_X1 U22535 ( .A1(n19567), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_8__SCAN_IN), .B2(n19566), .ZN(n19556) );
  OAI21_X1 U22536 ( .B1(n19557), .B2(n19569), .A(n19556), .ZN(P2_U2975) );
  AOI22_X1 U22537 ( .A1(n19567), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(
        P2_EAX_REG_10__SCAN_IN), .B2(n19566), .ZN(n19558) );
  OAI21_X1 U22538 ( .B1(n19559), .B2(n19569), .A(n19558), .ZN(P2_U2977) );
  AOI22_X1 U22539 ( .A1(n19567), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_12__SCAN_IN), .B2(n19566), .ZN(n19560) );
  OAI21_X1 U22540 ( .B1(n19561), .B2(n19569), .A(n19560), .ZN(P2_U2979) );
  AOI22_X1 U22541 ( .A1(n19567), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_13__SCAN_IN), .B2(n19566), .ZN(n19563) );
  NAND2_X1 U22542 ( .A1(n19563), .A2(n19562), .ZN(P2_U2980) );
  AOI22_X1 U22543 ( .A1(n19567), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_14__SCAN_IN), .B2(n19566), .ZN(n19565) );
  NAND2_X1 U22544 ( .A1(n19565), .A2(n19564), .ZN(P2_U2981) );
  AOI22_X1 U22545 ( .A1(n19567), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(
        P2_EAX_REG_15__SCAN_IN), .B2(n19566), .ZN(n19568) );
  OAI21_X1 U22546 ( .B1(n19570), .B2(n19569), .A(n19568), .ZN(P2_U2982) );
  AOI22_X1 U22547 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19584), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19571), .ZN(n19580) );
  OAI22_X1 U22548 ( .A1(n19575), .A2(n19574), .B1(n19573), .B2(n19572), .ZN(
        n19576) );
  AOI21_X1 U22549 ( .B1(n19578), .B2(n19577), .A(n19576), .ZN(n19579) );
  OAI211_X1 U22550 ( .C1(n19582), .C2(n19581), .A(n19580), .B(n19579), .ZN(
        P2_U3010) );
  NOR2_X1 U22551 ( .A1(n19584), .A2(n19583), .ZN(n19596) );
  INV_X1 U22552 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19595) );
  NAND2_X1 U22553 ( .A1(n19586), .A2(n19585), .ZN(n19588) );
  OAI211_X1 U22554 ( .C1(n19590), .C2(n19589), .A(n19588), .B(n19587), .ZN(
        n19591) );
  AOI21_X1 U22555 ( .B1(n19593), .B2(n19592), .A(n19591), .ZN(n19594) );
  OAI21_X1 U22556 ( .B1(n19596), .B2(n19595), .A(n19594), .ZN(P2_U3014) );
  NOR2_X1 U22557 ( .A1(n19871), .A2(n19683), .ZN(n19645) );
  INV_X1 U22558 ( .A(n19645), .ZN(n19633) );
  OAI22_X1 U22559 ( .A1(n20187), .A2(n20139), .B1(n19633), .B2(n20071), .ZN(
        n19599) );
  INV_X1 U22560 ( .A(n19599), .ZN(n19609) );
  AOI21_X1 U22561 ( .B1(n20187), .B2(n19680), .A(n20272), .ZN(n19600) );
  NOR2_X1 U22562 ( .A1(n19600), .A2(n20268), .ZN(n19604) );
  AOI21_X1 U22563 ( .B1(n19605), .B2(n20306), .A(n20305), .ZN(n19601) );
  AOI21_X1 U22564 ( .B1(n19604), .B2(n19603), .A(n19601), .ZN(n19602) );
  OAI21_X2 U22565 ( .B1(n19602), .B2(n19645), .A(n20133), .ZN(n19648) );
  INV_X1 U22566 ( .A(n19603), .ZN(n20179) );
  OAI21_X1 U22567 ( .B1(n20179), .B2(n19645), .A(n19604), .ZN(n19607) );
  OAI21_X1 U22568 ( .B1(n19605), .B2(n19645), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19606) );
  AOI22_X1 U22569 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19648), .B1(
        n20127), .B2(n19647), .ZN(n19608) );
  OAI211_X1 U22570 ( .C1(n20084), .C2(n19680), .A(n19609), .B(n19608), .ZN(
        P2_U3048) );
  AOI22_X1 U22571 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19639), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19638), .ZN(n20089) );
  AOI22_X2 U22572 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19639), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19638), .ZN(n20145) );
  NAND2_X1 U22573 ( .A1(n19644), .A2(n10884), .ZN(n20085) );
  OAI22_X1 U22574 ( .A1(n20187), .A2(n20145), .B1(n19633), .B2(n20085), .ZN(
        n19610) );
  INV_X1 U22575 ( .A(n19610), .ZN(n19613) );
  AOI22_X1 U22576 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19648), .B1(
        n20141), .B2(n19647), .ZN(n19612) );
  OAI211_X1 U22577 ( .C1(n20089), .C2(n19680), .A(n19613), .B(n19612), .ZN(
        P2_U3049) );
  AOI22_X2 U22578 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n19638), .B1(
        BUF1_REG_18__SCAN_IN), .B2(n19639), .ZN(n20151) );
  AOI22_X1 U22579 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19639), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19638), .ZN(n20094) );
  NAND2_X1 U22580 ( .A1(n19644), .A2(n19614), .ZN(n20090) );
  OAI22_X1 U22581 ( .A1(n20187), .A2(n20094), .B1(n19633), .B2(n20090), .ZN(
        n19615) );
  INV_X1 U22582 ( .A(n19615), .ZN(n19618) );
  AOI22_X1 U22583 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19648), .B1(
        n20147), .B2(n19647), .ZN(n19617) );
  OAI211_X1 U22584 ( .C1(n20151), .C2(n19680), .A(n19618), .B(n19617), .ZN(
        P2_U3050) );
  AOI22_X2 U22585 ( .A1(BUF2_REG_19__SCAN_IN), .A2(n19638), .B1(
        BUF1_REG_19__SCAN_IN), .B2(n19639), .ZN(n20157) );
  AOI22_X1 U22586 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19638), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n19639), .ZN(n20096) );
  NAND2_X1 U22587 ( .A1(n19644), .A2(n19619), .ZN(n20095) );
  OAI22_X1 U22588 ( .A1(n20187), .A2(n20096), .B1(n19633), .B2(n20095), .ZN(
        n19620) );
  INV_X1 U22589 ( .A(n19620), .ZN(n19623) );
  AOI22_X1 U22590 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19648), .B1(
        n20153), .B2(n19647), .ZN(n19622) );
  OAI211_X1 U22591 ( .C1(n20157), .C2(n19680), .A(n19623), .B(n19622), .ZN(
        P2_U3051) );
  AOI22_X1 U22592 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n19638), .B1(
        BUF1_REG_20__SCAN_IN), .B2(n19639), .ZN(n20163) );
  AOI22_X1 U22593 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19639), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19638), .ZN(n20104) );
  NAND2_X1 U22594 ( .A1(n19644), .A2(n19624), .ZN(n20100) );
  OAI22_X1 U22595 ( .A1(n20187), .A2(n20104), .B1(n19633), .B2(n20100), .ZN(
        n19625) );
  INV_X1 U22596 ( .A(n19625), .ZN(n19628) );
  AOI22_X1 U22597 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19648), .B1(
        n20159), .B2(n19647), .ZN(n19627) );
  OAI211_X1 U22598 ( .C1(n20163), .C2(n19680), .A(n19628), .B(n19627), .ZN(
        P2_U3052) );
  INV_X1 U22599 ( .A(n20164), .ZN(n20105) );
  OAI22_X1 U22600 ( .A1(n20187), .A2(n20171), .B1(n20105), .B2(n19633), .ZN(
        n19629) );
  INV_X1 U22601 ( .A(n19629), .ZN(n19631) );
  AOI22_X1 U22602 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19648), .B1(
        n20165), .B2(n19647), .ZN(n19630) );
  OAI211_X1 U22603 ( .C1(n20106), .C2(n19680), .A(n19631), .B(n19630), .ZN(
        P2_U3053) );
  INV_X1 U22604 ( .A(n19638), .ZN(n19640) );
  INV_X1 U22605 ( .A(n19639), .ZN(n19642) );
  AOI22_X1 U22606 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19638), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n19639), .ZN(n20111) );
  AND2_X1 U22607 ( .A1(n19644), .A2(n10889), .ZN(n20172) );
  INV_X1 U22608 ( .A(n20172), .ZN(n20110) );
  OAI22_X1 U22609 ( .A1(n20187), .A2(n20111), .B1(n19633), .B2(n20110), .ZN(
        n19634) );
  INV_X1 U22610 ( .A(n19634), .ZN(n19637) );
  AOI22_X1 U22611 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19648), .B1(
        n20173), .B2(n19647), .ZN(n19636) );
  OAI211_X1 U22612 ( .C1(n20177), .C2(n19680), .A(n19637), .B(n19636), .ZN(
        P2_U3054) );
  AOI22_X2 U22613 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19639), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19638), .ZN(n20188) );
  INV_X1 U22614 ( .A(n20187), .ZN(n20167) );
  AOI22_X1 U22615 ( .A1(n20182), .A2(n20167), .B1(n19645), .B2(n20178), .ZN(
        n19650) );
  AOI22_X1 U22616 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19648), .B1(
        n20180), .B2(n19647), .ZN(n19649) );
  OAI211_X1 U22617 ( .C1(n20188), .C2(n19680), .A(n19650), .B(n19649), .ZN(
        P2_U3055) );
  NAND2_X1 U22618 ( .A1(n19911), .A2(n19681), .ZN(n19657) );
  INV_X1 U22619 ( .A(n19651), .ZN(n19653) );
  INV_X1 U22620 ( .A(n19657), .ZN(n19652) );
  NAND2_X1 U22621 ( .A1(n19652), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19655) );
  NAND3_X1 U22622 ( .A1(n19653), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19655), 
        .ZN(n19659) );
  INV_X1 U22623 ( .A(n19659), .ZN(n19654) );
  AOI211_X2 U22624 ( .C1(n20317), .C2(n19657), .A(n19741), .B(n19654), .ZN(
        n19676) );
  INV_X1 U22625 ( .A(n19655), .ZN(n19675) );
  AOI22_X1 U22626 ( .A1(n19676), .A2(n20127), .B1(n20126), .B2(n19675), .ZN(
        n19662) );
  NAND3_X1 U22627 ( .A1(n19845), .A2(n19870), .A3(n20306), .ZN(n19656) );
  OAI21_X1 U22628 ( .B1(n19658), .B2(n19657), .A(n19656), .ZN(n19660) );
  NAND3_X1 U22629 ( .A1(n19660), .A2(n20133), .A3(n19659), .ZN(n19677) );
  INV_X1 U22630 ( .A(n20084), .ZN(n20136) );
  AOI22_X1 U22631 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19677), .B1(
        n19708), .B2(n20136), .ZN(n19661) );
  OAI211_X1 U22632 ( .C1(n20139), .C2(n19680), .A(n19662), .B(n19661), .ZN(
        P2_U3056) );
  AOI22_X1 U22633 ( .A1(n19676), .A2(n20141), .B1(n20140), .B2(n19675), .ZN(
        n19664) );
  INV_X1 U22634 ( .A(n20089), .ZN(n20142) );
  AOI22_X1 U22635 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19677), .B1(
        n19708), .B2(n20142), .ZN(n19663) );
  OAI211_X1 U22636 ( .C1(n20145), .C2(n19680), .A(n19664), .B(n19663), .ZN(
        P2_U3057) );
  AOI22_X1 U22637 ( .A1(n19676), .A2(n20147), .B1(n20146), .B2(n19675), .ZN(
        n19666) );
  INV_X1 U22638 ( .A(n20151), .ZN(n20013) );
  AOI22_X1 U22639 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19677), .B1(
        n19708), .B2(n20013), .ZN(n19665) );
  OAI211_X1 U22640 ( .C1(n20094), .C2(n19680), .A(n19666), .B(n19665), .ZN(
        P2_U3058) );
  AOI22_X1 U22641 ( .A1(n19676), .A2(n20153), .B1(n20152), .B2(n19675), .ZN(
        n19668) );
  INV_X1 U22642 ( .A(n20157), .ZN(n20017) );
  AOI22_X1 U22643 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19677), .B1(
        n19708), .B2(n20017), .ZN(n19667) );
  OAI211_X1 U22644 ( .C1(n20096), .C2(n19680), .A(n19668), .B(n19667), .ZN(
        P2_U3059) );
  AOI22_X1 U22645 ( .A1(n19676), .A2(n20159), .B1(n20158), .B2(n19675), .ZN(
        n19670) );
  INV_X1 U22646 ( .A(n20163), .ZN(n20021) );
  AOI22_X1 U22647 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19677), .B1(
        n19708), .B2(n20021), .ZN(n19669) );
  OAI211_X1 U22648 ( .C1(n20104), .C2(n19680), .A(n19670), .B(n19669), .ZN(
        P2_U3060) );
  AOI22_X1 U22649 ( .A1(n19676), .A2(n20165), .B1(n20164), .B2(n19675), .ZN(
        n19672) );
  AOI22_X1 U22650 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19677), .B1(
        n19708), .B2(n20166), .ZN(n19671) );
  OAI211_X1 U22651 ( .C1(n20171), .C2(n19680), .A(n19672), .B(n19671), .ZN(
        P2_U3061) );
  AOI22_X1 U22652 ( .A1(n19676), .A2(n20173), .B1(n20172), .B2(n19675), .ZN(
        n19674) );
  AOI22_X1 U22653 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19677), .B1(
        n19708), .B2(n20025), .ZN(n19673) );
  OAI211_X1 U22654 ( .C1(n20111), .C2(n19680), .A(n19674), .B(n19673), .ZN(
        P2_U3062) );
  AOI22_X1 U22655 ( .A1(n19676), .A2(n20180), .B1(n20178), .B2(n19675), .ZN(
        n19679) );
  INV_X1 U22656 ( .A(n20188), .ZN(n20032) );
  AOI22_X1 U22657 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19677), .B1(
        n19708), .B2(n20032), .ZN(n19678) );
  OAI211_X1 U22658 ( .C1(n20123), .C2(n19680), .A(n19679), .B(n19678), .ZN(
        P2_U3063) );
  NAND2_X1 U22659 ( .A1(n19805), .A2(n19681), .ZN(n19686) );
  NAND2_X1 U22660 ( .A1(n19682), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19949) );
  OR2_X1 U22661 ( .A1(n19949), .A2(n19683), .ZN(n19688) );
  INV_X1 U22662 ( .A(n19688), .ZN(n19706) );
  OAI21_X1 U22663 ( .B1(n19687), .B2(n19706), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19684) );
  OAI21_X1 U22664 ( .B1(n19686), .B2(n20268), .A(n19684), .ZN(n19707) );
  AOI22_X1 U22665 ( .A1(n19707), .A2(n20127), .B1(n20126), .B2(n19706), .ZN(
        n19693) );
  OAI21_X1 U22666 ( .B1(n19733), .B2(n19708), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19685) );
  NAND2_X1 U22667 ( .A1(n19686), .A2(n19685), .ZN(n19691) );
  INV_X1 U22668 ( .A(n19687), .ZN(n19689) );
  OAI211_X1 U22669 ( .C1(n19689), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19688), 
        .B(n20268), .ZN(n19690) );
  NAND3_X1 U22670 ( .A1(n19691), .A2(n20133), .A3(n19690), .ZN(n19709) );
  AOI22_X1 U22671 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19709), .B1(
        n19708), .B2(n20047), .ZN(n19692) );
  OAI211_X1 U22672 ( .C1(n20084), .C2(n19726), .A(n19693), .B(n19692), .ZN(
        P2_U3064) );
  AOI22_X1 U22673 ( .A1(n19707), .A2(n20141), .B1(n19706), .B2(n20140), .ZN(
        n19695) );
  INV_X1 U22674 ( .A(n20145), .ZN(n20050) );
  AOI22_X1 U22675 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19709), .B1(
        n19708), .B2(n20050), .ZN(n19694) );
  OAI211_X1 U22676 ( .C1(n20089), .C2(n19726), .A(n19695), .B(n19694), .ZN(
        P2_U3065) );
  AOI22_X1 U22677 ( .A1(n19707), .A2(n20147), .B1(n19706), .B2(n20146), .ZN(
        n19697) );
  INV_X1 U22678 ( .A(n20094), .ZN(n20148) );
  AOI22_X1 U22679 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19709), .B1(
        n19708), .B2(n20148), .ZN(n19696) );
  OAI211_X1 U22680 ( .C1(n20151), .C2(n19726), .A(n19697), .B(n19696), .ZN(
        P2_U3066) );
  AOI22_X1 U22681 ( .A1(n19707), .A2(n20153), .B1(n19706), .B2(n20152), .ZN(
        n19699) );
  INV_X1 U22682 ( .A(n20096), .ZN(n20154) );
  AOI22_X1 U22683 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19709), .B1(
        n19708), .B2(n20154), .ZN(n19698) );
  OAI211_X1 U22684 ( .C1(n20157), .C2(n19726), .A(n19699), .B(n19698), .ZN(
        P2_U3067) );
  AOI22_X1 U22685 ( .A1(n19707), .A2(n20159), .B1(n19706), .B2(n20158), .ZN(
        n19701) );
  INV_X1 U22686 ( .A(n20104), .ZN(n20160) );
  AOI22_X1 U22687 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19709), .B1(
        n19708), .B2(n20160), .ZN(n19700) );
  OAI211_X1 U22688 ( .C1(n20163), .C2(n19726), .A(n19701), .B(n19700), .ZN(
        P2_U3068) );
  AOI22_X1 U22689 ( .A1(n19707), .A2(n20165), .B1(n20164), .B2(n19706), .ZN(
        n19703) );
  AOI22_X1 U22690 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19709), .B1(
        n19708), .B2(n20059), .ZN(n19702) );
  OAI211_X1 U22691 ( .C1(n20106), .C2(n19726), .A(n19703), .B(n19702), .ZN(
        P2_U3069) );
  AOI22_X1 U22692 ( .A1(n19707), .A2(n20173), .B1(n19706), .B2(n20172), .ZN(
        n19705) );
  INV_X1 U22693 ( .A(n20111), .ZN(n20174) );
  AOI22_X1 U22694 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19709), .B1(
        n19708), .B2(n20174), .ZN(n19704) );
  OAI211_X1 U22695 ( .C1(n20177), .C2(n19726), .A(n19705), .B(n19704), .ZN(
        P2_U3070) );
  AOI22_X1 U22696 ( .A1(n19707), .A2(n20180), .B1(n19706), .B2(n20178), .ZN(
        n19711) );
  AOI22_X1 U22697 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19709), .B1(
        n19708), .B2(n20182), .ZN(n19710) );
  OAI211_X1 U22698 ( .C1(n20188), .C2(n19726), .A(n19711), .B(n19710), .ZN(
        P2_U3071) );
  OAI22_X1 U22699 ( .A1(n19718), .A2(n20089), .B1(n19725), .B2(n20085), .ZN(
        n19712) );
  INV_X1 U22700 ( .A(n19712), .ZN(n19714) );
  AOI22_X1 U22701 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19735), .B1(
        n20141), .B2(n19734), .ZN(n19713) );
  OAI211_X1 U22702 ( .C1(n20145), .C2(n19726), .A(n19714), .B(n19713), .ZN(
        P2_U3073) );
  OAI22_X1 U22703 ( .A1(n19718), .A2(n20151), .B1(n19725), .B2(n20090), .ZN(
        n19715) );
  INV_X1 U22704 ( .A(n19715), .ZN(n19717) );
  AOI22_X1 U22705 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19735), .B1(
        n20147), .B2(n19734), .ZN(n19716) );
  OAI211_X1 U22706 ( .C1(n20094), .C2(n19726), .A(n19717), .B(n19716), .ZN(
        P2_U3074) );
  OAI22_X1 U22707 ( .A1(n19726), .A2(n20096), .B1(n19725), .B2(n20095), .ZN(
        n19719) );
  INV_X1 U22708 ( .A(n19719), .ZN(n19721) );
  AOI22_X1 U22709 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19735), .B1(
        n20153), .B2(n19734), .ZN(n19720) );
  OAI211_X1 U22710 ( .C1(n20157), .C2(n19718), .A(n19721), .B(n19720), .ZN(
        P2_U3075) );
  OAI22_X1 U22711 ( .A1(n19726), .A2(n20104), .B1(n19725), .B2(n20100), .ZN(
        n19722) );
  INV_X1 U22712 ( .A(n19722), .ZN(n19724) );
  AOI22_X1 U22713 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19735), .B1(
        n20159), .B2(n19734), .ZN(n19723) );
  OAI211_X1 U22714 ( .C1(n20163), .C2(n19718), .A(n19724), .B(n19723), .ZN(
        P2_U3076) );
  OAI22_X1 U22715 ( .A1(n19726), .A2(n20171), .B1(n20105), .B2(n19725), .ZN(
        n19727) );
  INV_X1 U22716 ( .A(n19727), .ZN(n19729) );
  AOI22_X1 U22717 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19735), .B1(
        n20165), .B2(n19734), .ZN(n19728) );
  OAI211_X1 U22718 ( .C1(n20106), .C2(n19718), .A(n19729), .B(n19728), .ZN(
        P2_U3077) );
  AOI22_X1 U22719 ( .A1(n20025), .A2(n19763), .B1(n19732), .B2(n20172), .ZN(
        n19731) );
  AOI22_X1 U22720 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19735), .B1(
        n20173), .B2(n19734), .ZN(n19730) );
  OAI211_X1 U22721 ( .C1(n20111), .C2(n19726), .A(n19731), .B(n19730), .ZN(
        P2_U3078) );
  AOI22_X1 U22722 ( .A1(n20182), .A2(n19733), .B1(n19732), .B2(n20178), .ZN(
        n19737) );
  AOI22_X1 U22723 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19735), .B1(
        n20180), .B2(n19734), .ZN(n19736) );
  OAI211_X1 U22724 ( .C1(n20188), .C2(n19718), .A(n19737), .B(n19736), .ZN(
        P2_U3079) );
  NAND3_X1 U22725 ( .A1(n19739), .A2(n19738), .A3(n20284), .ZN(n19743) );
  NAND2_X1 U22726 ( .A1(n20284), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19816) );
  NOR2_X1 U22727 ( .A1(n19871), .A2(n19816), .ZN(n19761) );
  NOR3_X1 U22728 ( .A1(n19740), .A2(n19761), .A3(n20317), .ZN(n19742) );
  AOI211_X2 U22729 ( .C1(n20317), .C2(n19743), .A(n19741), .B(n19742), .ZN(
        n19762) );
  AOI22_X1 U22730 ( .A1(n19762), .A2(n20127), .B1(n20126), .B2(n19761), .ZN(
        n19747) );
  OAI21_X1 U22731 ( .B1(n19763), .B2(n19756), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19744) );
  AOI211_X1 U22732 ( .C1(n19744), .C2(n19743), .A(n19808), .B(n19742), .ZN(
        n19745) );
  AOI22_X1 U22733 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19764), .B1(
        n19763), .B2(n20047), .ZN(n19746) );
  OAI211_X1 U22734 ( .C1(n20084), .C2(n19794), .A(n19747), .B(n19746), .ZN(
        P2_U3080) );
  AOI22_X1 U22735 ( .A1(n19762), .A2(n20141), .B1(n20140), .B2(n19761), .ZN(
        n19749) );
  AOI22_X1 U22736 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19764), .B1(
        n19756), .B2(n20142), .ZN(n19748) );
  OAI211_X1 U22737 ( .C1(n20145), .C2(n19718), .A(n19749), .B(n19748), .ZN(
        P2_U3081) );
  AOI22_X1 U22738 ( .A1(n19762), .A2(n20147), .B1(n20146), .B2(n19761), .ZN(
        n19751) );
  AOI22_X1 U22739 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19764), .B1(
        n19756), .B2(n20013), .ZN(n19750) );
  OAI211_X1 U22740 ( .C1(n20094), .C2(n19718), .A(n19751), .B(n19750), .ZN(
        P2_U3082) );
  AOI22_X1 U22741 ( .A1(n19762), .A2(n20153), .B1(n20152), .B2(n19761), .ZN(
        n19753) );
  AOI22_X1 U22742 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19764), .B1(
        n19763), .B2(n20154), .ZN(n19752) );
  OAI211_X1 U22743 ( .C1(n20157), .C2(n19794), .A(n19753), .B(n19752), .ZN(
        P2_U3083) );
  AOI22_X1 U22744 ( .A1(n19762), .A2(n20159), .B1(n20158), .B2(n19761), .ZN(
        n19755) );
  AOI22_X1 U22745 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19764), .B1(
        n19756), .B2(n20021), .ZN(n19754) );
  OAI211_X1 U22746 ( .C1(n20104), .C2(n19718), .A(n19755), .B(n19754), .ZN(
        P2_U3084) );
  AOI22_X1 U22747 ( .A1(n19762), .A2(n20165), .B1(n20164), .B2(n19761), .ZN(
        n19758) );
  AOI22_X1 U22748 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19764), .B1(
        n19756), .B2(n20166), .ZN(n19757) );
  OAI211_X1 U22749 ( .C1(n20171), .C2(n19718), .A(n19758), .B(n19757), .ZN(
        P2_U3085) );
  AOI22_X1 U22750 ( .A1(n19762), .A2(n20173), .B1(n20172), .B2(n19761), .ZN(
        n19760) );
  AOI22_X1 U22751 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19764), .B1(
        n19763), .B2(n20174), .ZN(n19759) );
  OAI211_X1 U22752 ( .C1(n20177), .C2(n19794), .A(n19760), .B(n19759), .ZN(
        P2_U3086) );
  AOI22_X1 U22753 ( .A1(n19762), .A2(n20180), .B1(n20178), .B2(n19761), .ZN(
        n19766) );
  AOI22_X1 U22754 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19764), .B1(
        n19763), .B2(n20182), .ZN(n19765) );
  OAI211_X1 U22755 ( .C1(n20188), .C2(n19794), .A(n19766), .B(n19765), .ZN(
        P2_U3087) );
  NOR2_X1 U22756 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19816), .ZN(
        n19771) );
  NAND2_X1 U22757 ( .A1(n19771), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19798) );
  OAI22_X1 U22758 ( .A1(n19839), .A2(n20084), .B1(n19798), .B2(n20071), .ZN(
        n19767) );
  INV_X1 U22759 ( .A(n19767), .ZN(n19778) );
  INV_X1 U22760 ( .A(n19845), .ZN(n19768) );
  OAI21_X1 U22761 ( .B1(n19768), .B2(n20043), .A(n20305), .ZN(n19776) );
  OAI21_X1 U22762 ( .B1(n19773), .B2(n20317), .A(n20306), .ZN(n19769) );
  AOI21_X1 U22763 ( .B1(n19769), .B2(n19798), .A(n19808), .ZN(n19770) );
  INV_X1 U22764 ( .A(n19771), .ZN(n19775) );
  INV_X1 U22765 ( .A(n19798), .ZN(n19772) );
  OAI21_X1 U22766 ( .B1(n19773), .B2(n19772), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19774) );
  AOI22_X1 U22767 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19801), .B1(
        n20127), .B2(n19800), .ZN(n19777) );
  OAI211_X1 U22768 ( .C1(n20139), .C2(n19794), .A(n19778), .B(n19777), .ZN(
        P2_U3088) );
  OAI22_X1 U22769 ( .A1(n19839), .A2(n20089), .B1(n19798), .B2(n20085), .ZN(
        n19779) );
  INV_X1 U22770 ( .A(n19779), .ZN(n19781) );
  AOI22_X1 U22771 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19801), .B1(
        n20141), .B2(n19800), .ZN(n19780) );
  OAI211_X1 U22772 ( .C1(n20145), .C2(n19794), .A(n19781), .B(n19780), .ZN(
        P2_U3089) );
  OAI22_X1 U22773 ( .A1(n19794), .A2(n20094), .B1(n19798), .B2(n20090), .ZN(
        n19782) );
  INV_X1 U22774 ( .A(n19782), .ZN(n19784) );
  AOI22_X1 U22775 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19801), .B1(
        n20147), .B2(n19800), .ZN(n19783) );
  OAI211_X1 U22776 ( .C1(n20151), .C2(n19839), .A(n19784), .B(n19783), .ZN(
        P2_U3090) );
  OAI22_X1 U22777 ( .A1(n19839), .A2(n20157), .B1(n19798), .B2(n20095), .ZN(
        n19785) );
  INV_X1 U22778 ( .A(n19785), .ZN(n19787) );
  AOI22_X1 U22779 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19801), .B1(
        n20153), .B2(n19800), .ZN(n19786) );
  OAI211_X1 U22780 ( .C1(n20096), .C2(n19794), .A(n19787), .B(n19786), .ZN(
        P2_U3091) );
  OAI22_X1 U22781 ( .A1(n19794), .A2(n20104), .B1(n19798), .B2(n20100), .ZN(
        n19788) );
  INV_X1 U22782 ( .A(n19788), .ZN(n19790) );
  AOI22_X1 U22783 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19801), .B1(
        n20159), .B2(n19800), .ZN(n19789) );
  OAI211_X1 U22784 ( .C1(n20163), .C2(n19839), .A(n19790), .B(n19789), .ZN(
        P2_U3092) );
  OAI22_X1 U22785 ( .A1(n19839), .A2(n20106), .B1(n20105), .B2(n19798), .ZN(
        n19791) );
  INV_X1 U22786 ( .A(n19791), .ZN(n19793) );
  AOI22_X1 U22787 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19801), .B1(
        n20165), .B2(n19800), .ZN(n19792) );
  OAI211_X1 U22788 ( .C1(n20171), .C2(n19794), .A(n19793), .B(n19792), .ZN(
        P2_U3093) );
  OAI22_X1 U22789 ( .A1(n19794), .A2(n20111), .B1(n19798), .B2(n20110), .ZN(
        n19795) );
  INV_X1 U22790 ( .A(n19795), .ZN(n19797) );
  AOI22_X1 U22791 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19801), .B1(
        n20173), .B2(n19800), .ZN(n19796) );
  OAI211_X1 U22792 ( .C1(n20177), .C2(n19839), .A(n19797), .B(n19796), .ZN(
        P2_U3094) );
  INV_X1 U22793 ( .A(n20178), .ZN(n20116) );
  OAI22_X1 U22794 ( .A1(n19839), .A2(n20188), .B1(n19798), .B2(n20116), .ZN(
        n19799) );
  INV_X1 U22795 ( .A(n19799), .ZN(n19803) );
  AOI22_X1 U22796 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19801), .B1(
        n20180), .B2(n19800), .ZN(n19802) );
  OAI211_X1 U22797 ( .C1(n20123), .C2(n19794), .A(n19803), .B(n19802), .ZN(
        P2_U3095) );
  INV_X1 U22798 ( .A(n19839), .ZN(n19817) );
  OAI21_X1 U22799 ( .B1(n19817), .B2(n19866), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19807) );
  INV_X1 U22800 ( .A(n19816), .ZN(n19841) );
  NAND2_X1 U22801 ( .A1(n19805), .A2(n19841), .ZN(n19806) );
  NAND2_X1 U22802 ( .A1(n19807), .A2(n19806), .ZN(n19812) );
  NAND2_X1 U22803 ( .A1(n19814), .A2(n20306), .ZN(n19810) );
  NOR3_X2 U22804 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n20130), .ZN(n19834) );
  NOR2_X1 U22805 ( .A1(n20305), .A2(n19834), .ZN(n19809) );
  AOI21_X1 U22806 ( .B1(n19810), .B2(n19809), .A(n19808), .ZN(n19811) );
  INV_X1 U22807 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n19820) );
  INV_X1 U22808 ( .A(n19813), .ZN(n19951) );
  OAI21_X1 U22809 ( .B1(n19814), .B2(n19834), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19815) );
  OAI21_X1 U22810 ( .B1(n19816), .B2(n19951), .A(n19815), .ZN(n19835) );
  AOI22_X1 U22811 ( .A1(n19835), .A2(n20127), .B1(n20126), .B2(n19834), .ZN(
        n19819) );
  AOI22_X1 U22812 ( .A1(n19817), .A2(n20047), .B1(n19866), .B2(n20136), .ZN(
        n19818) );
  OAI211_X1 U22813 ( .C1(n19821), .C2(n19820), .A(n19819), .B(n19818), .ZN(
        P2_U3096) );
  AOI22_X1 U22814 ( .A1(n19835), .A2(n20141), .B1(n20140), .B2(n19834), .ZN(
        n19823) );
  AOI22_X1 U22815 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19836), .B1(
        n19866), .B2(n20142), .ZN(n19822) );
  OAI211_X1 U22816 ( .C1(n20145), .C2(n19839), .A(n19823), .B(n19822), .ZN(
        P2_U3097) );
  AOI22_X1 U22817 ( .A1(n19835), .A2(n20147), .B1(n20146), .B2(n19834), .ZN(
        n19825) );
  AOI22_X1 U22818 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19836), .B1(
        n19866), .B2(n20013), .ZN(n19824) );
  OAI211_X1 U22819 ( .C1(n20094), .C2(n19839), .A(n19825), .B(n19824), .ZN(
        P2_U3098) );
  AOI22_X1 U22820 ( .A1(n19835), .A2(n20153), .B1(n20152), .B2(n19834), .ZN(
        n19827) );
  AOI22_X1 U22821 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19836), .B1(
        n19866), .B2(n20017), .ZN(n19826) );
  OAI211_X1 U22822 ( .C1(n20096), .C2(n19839), .A(n19827), .B(n19826), .ZN(
        P2_U3099) );
  AOI22_X1 U22823 ( .A1(n19835), .A2(n20159), .B1(n20158), .B2(n19834), .ZN(
        n19829) );
  AOI22_X1 U22824 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19836), .B1(
        n19866), .B2(n20021), .ZN(n19828) );
  OAI211_X1 U22825 ( .C1(n20104), .C2(n19839), .A(n19829), .B(n19828), .ZN(
        P2_U3100) );
  AOI22_X1 U22826 ( .A1(n19835), .A2(n20165), .B1(n20164), .B2(n19834), .ZN(
        n19831) );
  AOI22_X1 U22827 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19836), .B1(
        n19866), .B2(n20166), .ZN(n19830) );
  OAI211_X1 U22828 ( .C1(n20171), .C2(n19839), .A(n19831), .B(n19830), .ZN(
        P2_U3101) );
  AOI22_X1 U22829 ( .A1(n19835), .A2(n20173), .B1(n20172), .B2(n19834), .ZN(
        n19833) );
  AOI22_X1 U22830 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19836), .B1(
        n19866), .B2(n20025), .ZN(n19832) );
  OAI211_X1 U22831 ( .C1(n20111), .C2(n19839), .A(n19833), .B(n19832), .ZN(
        P2_U3102) );
  AOI22_X1 U22832 ( .A1(n19835), .A2(n20180), .B1(n20178), .B2(n19834), .ZN(
        n19838) );
  AOI22_X1 U22833 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19836), .B1(
        n19866), .B2(n20032), .ZN(n19837) );
  OAI211_X1 U22834 ( .C1(n20123), .C2(n19839), .A(n19838), .B(n19837), .ZN(
        P2_U3103) );
  NOR2_X1 U22835 ( .A1(n20130), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19849) );
  INV_X1 U22836 ( .A(n19849), .ZN(n19844) );
  NAND2_X1 U22837 ( .A1(n19842), .A2(n19841), .ZN(n19875) );
  INV_X1 U22838 ( .A(n19875), .ZN(n19878) );
  OAI21_X1 U22839 ( .B1(n19846), .B2(n19878), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19843) );
  OAI21_X1 U22840 ( .B1(n19844), .B2(n20268), .A(n19843), .ZN(n19865) );
  AOI22_X1 U22841 ( .A1(n19865), .A2(n20127), .B1(n20126), .B2(n19878), .ZN(
        n19852) );
  NAND2_X1 U22842 ( .A1(n19845), .A2(n20069), .ZN(n20269) );
  INV_X1 U22843 ( .A(n20269), .ZN(n19850) );
  INV_X1 U22844 ( .A(n19846), .ZN(n19847) );
  OAI211_X1 U22845 ( .C1(n19847), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19875), 
        .B(n20268), .ZN(n19848) );
  OAI211_X1 U22846 ( .C1(n19850), .C2(n19849), .A(n20133), .B(n19848), .ZN(
        n19867) );
  AOI22_X1 U22847 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19867), .B1(
        n19866), .B2(n20047), .ZN(n19851) );
  OAI211_X1 U22848 ( .C1(n20084), .C2(n19909), .A(n19852), .B(n19851), .ZN(
        P2_U3104) );
  AOI22_X1 U22849 ( .A1(n19865), .A2(n20141), .B1(n19878), .B2(n20140), .ZN(
        n19854) );
  AOI22_X1 U22850 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19867), .B1(
        n19866), .B2(n20050), .ZN(n19853) );
  OAI211_X1 U22851 ( .C1(n20089), .C2(n19909), .A(n19854), .B(n19853), .ZN(
        P2_U3105) );
  AOI22_X1 U22852 ( .A1(n19865), .A2(n20147), .B1(n19878), .B2(n20146), .ZN(
        n19856) );
  AOI22_X1 U22853 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19867), .B1(
        n19866), .B2(n20148), .ZN(n19855) );
  OAI211_X1 U22854 ( .C1(n20151), .C2(n19909), .A(n19856), .B(n19855), .ZN(
        P2_U3106) );
  AOI22_X1 U22855 ( .A1(n19865), .A2(n20153), .B1(n19878), .B2(n20152), .ZN(
        n19858) );
  AOI22_X1 U22856 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19867), .B1(
        n19866), .B2(n20154), .ZN(n19857) );
  OAI211_X1 U22857 ( .C1(n20157), .C2(n19909), .A(n19858), .B(n19857), .ZN(
        P2_U3107) );
  AOI22_X1 U22858 ( .A1(n19865), .A2(n20159), .B1(n19878), .B2(n20158), .ZN(
        n19860) );
  AOI22_X1 U22859 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19867), .B1(
        n19866), .B2(n20160), .ZN(n19859) );
  OAI211_X1 U22860 ( .C1(n20163), .C2(n19909), .A(n19860), .B(n19859), .ZN(
        P2_U3108) );
  AOI22_X1 U22861 ( .A1(n19865), .A2(n20165), .B1(n20164), .B2(n19878), .ZN(
        n19862) );
  AOI22_X1 U22862 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19867), .B1(
        n19866), .B2(n20059), .ZN(n19861) );
  OAI211_X1 U22863 ( .C1(n20106), .C2(n19909), .A(n19862), .B(n19861), .ZN(
        P2_U3109) );
  AOI22_X1 U22864 ( .A1(n19865), .A2(n20173), .B1(n19878), .B2(n20172), .ZN(
        n19864) );
  AOI22_X1 U22865 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19867), .B1(
        n19866), .B2(n20174), .ZN(n19863) );
  OAI211_X1 U22866 ( .C1(n20177), .C2(n19909), .A(n19864), .B(n19863), .ZN(
        P2_U3110) );
  AOI22_X1 U22867 ( .A1(n19865), .A2(n20180), .B1(n19878), .B2(n20178), .ZN(
        n19869) );
  AOI22_X1 U22868 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19867), .B1(
        n19866), .B2(n20182), .ZN(n19868) );
  OAI211_X1 U22869 ( .C1(n20188), .C2(n19909), .A(n19869), .B(n19868), .ZN(
        P2_U3111) );
  NOR2_X1 U22870 ( .A1(n20284), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19981) );
  INV_X1 U22871 ( .A(n19981), .ZN(n19979) );
  NOR2_X1 U22872 ( .A1(n19979), .A2(n19871), .ZN(n19879) );
  INV_X1 U22873 ( .A(n19879), .ZN(n19903) );
  OAI22_X1 U22874 ( .A1(n19909), .A2(n20139), .B1(n19903), .B2(n20071), .ZN(
        n19872) );
  INV_X1 U22875 ( .A(n19872), .ZN(n19884) );
  NAND2_X1 U22876 ( .A1(n19947), .A2(n19909), .ZN(n19873) );
  AOI21_X1 U22877 ( .B1(n19873), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n20268), 
        .ZN(n19877) );
  OAI21_X1 U22878 ( .B1(n19880), .B2(n20317), .A(n20306), .ZN(n19874) );
  AOI21_X1 U22879 ( .B1(n19877), .B2(n19875), .A(n19874), .ZN(n19876) );
  OAI21_X2 U22880 ( .B1(n19879), .B2(n19876), .A(n20133), .ZN(n19906) );
  OAI21_X1 U22881 ( .B1(n19878), .B2(n19879), .A(n19877), .ZN(n19882) );
  OAI21_X1 U22882 ( .B1(n19880), .B2(n19879), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19881) );
  AOI22_X1 U22883 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19906), .B1(
        n20127), .B2(n19905), .ZN(n19883) );
  OAI211_X1 U22884 ( .C1(n20084), .C2(n19947), .A(n19884), .B(n19883), .ZN(
        P2_U3112) );
  OAI22_X1 U22885 ( .A1(n19947), .A2(n20089), .B1(n19903), .B2(n20085), .ZN(
        n19885) );
  INV_X1 U22886 ( .A(n19885), .ZN(n19887) );
  AOI22_X1 U22887 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19906), .B1(
        n19905), .B2(n20141), .ZN(n19886) );
  OAI211_X1 U22888 ( .C1(n20145), .C2(n19909), .A(n19887), .B(n19886), .ZN(
        P2_U3113) );
  OAI22_X1 U22889 ( .A1(n19947), .A2(n20151), .B1(n19903), .B2(n20090), .ZN(
        n19888) );
  INV_X1 U22890 ( .A(n19888), .ZN(n19890) );
  AOI22_X1 U22891 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19906), .B1(
        n19905), .B2(n20147), .ZN(n19889) );
  OAI211_X1 U22892 ( .C1(n20094), .C2(n19909), .A(n19890), .B(n19889), .ZN(
        P2_U3114) );
  OAI22_X1 U22893 ( .A1(n19909), .A2(n20096), .B1(n19903), .B2(n20095), .ZN(
        n19891) );
  INV_X1 U22894 ( .A(n19891), .ZN(n19893) );
  AOI22_X1 U22895 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19906), .B1(
        n19905), .B2(n20153), .ZN(n19892) );
  OAI211_X1 U22896 ( .C1(n20157), .C2(n19947), .A(n19893), .B(n19892), .ZN(
        P2_U3115) );
  OAI22_X1 U22897 ( .A1(n19947), .A2(n20163), .B1(n19903), .B2(n20100), .ZN(
        n19894) );
  INV_X1 U22898 ( .A(n19894), .ZN(n19896) );
  AOI22_X1 U22899 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19906), .B1(
        n19905), .B2(n20159), .ZN(n19895) );
  OAI211_X1 U22900 ( .C1(n20104), .C2(n19909), .A(n19896), .B(n19895), .ZN(
        P2_U3116) );
  OAI22_X1 U22901 ( .A1(n19909), .A2(n20171), .B1(n20105), .B2(n19903), .ZN(
        n19897) );
  INV_X1 U22902 ( .A(n19897), .ZN(n19899) );
  AOI22_X1 U22903 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19906), .B1(
        n19905), .B2(n20165), .ZN(n19898) );
  OAI211_X1 U22904 ( .C1(n20106), .C2(n19947), .A(n19899), .B(n19898), .ZN(
        P2_U3117) );
  OAI22_X1 U22905 ( .A1(n19909), .A2(n20111), .B1(n19903), .B2(n20110), .ZN(
        n19900) );
  INV_X1 U22906 ( .A(n19900), .ZN(n19902) );
  AOI22_X1 U22907 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19906), .B1(
        n19905), .B2(n20173), .ZN(n19901) );
  OAI211_X1 U22908 ( .C1(n20177), .C2(n19947), .A(n19902), .B(n19901), .ZN(
        P2_U3118) );
  OAI22_X1 U22909 ( .A1(n19947), .A2(n20188), .B1(n19903), .B2(n20116), .ZN(
        n19904) );
  INV_X1 U22910 ( .A(n19904), .ZN(n19908) );
  AOI22_X1 U22911 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19906), .B1(
        n19905), .B2(n20180), .ZN(n19907) );
  OAI211_X1 U22912 ( .C1(n20123), .C2(n19909), .A(n19908), .B(n19907), .ZN(
        P2_U3119) );
  NAND2_X1 U22913 ( .A1(n19911), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19912) );
  NOR2_X1 U22914 ( .A1(n19979), .A2(n19912), .ZN(n19953) );
  INV_X1 U22915 ( .A(n19953), .ZN(n19936) );
  NOR2_X1 U22916 ( .A1(n20071), .A2(n19936), .ZN(n19913) );
  AOI21_X1 U22917 ( .B1(n19974), .B2(n20136), .A(n19913), .ZN(n19923) );
  NAND2_X1 U22918 ( .A1(n20280), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20132) );
  OAI21_X1 U22919 ( .B1(n20132), .B2(n19914), .A(n20305), .ZN(n19921) );
  NOR2_X1 U22920 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19979), .ZN(
        n19917) );
  INV_X1 U22921 ( .A(n19918), .ZN(n19915) );
  OAI211_X1 U22922 ( .C1(n19915), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19936), 
        .B(n20268), .ZN(n19916) );
  INV_X1 U22923 ( .A(n19917), .ZN(n19920) );
  OAI21_X1 U22924 ( .B1(n19918), .B2(n19953), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19919) );
  AOI22_X1 U22925 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19944), .B1(
        n20127), .B2(n19943), .ZN(n19922) );
  OAI211_X1 U22926 ( .C1(n20139), .C2(n19947), .A(n19923), .B(n19922), .ZN(
        P2_U3120) );
  NOR2_X1 U22927 ( .A1(n20085), .A2(n19936), .ZN(n19924) );
  AOI21_X1 U22928 ( .B1(n19974), .B2(n20142), .A(n19924), .ZN(n19926) );
  AOI22_X1 U22929 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19944), .B1(
        n20141), .B2(n19943), .ZN(n19925) );
  OAI211_X1 U22930 ( .C1(n20145), .C2(n19947), .A(n19926), .B(n19925), .ZN(
        P2_U3121) );
  INV_X1 U22931 ( .A(n19974), .ZN(n19940) );
  OAI22_X1 U22932 ( .A1(n19947), .A2(n20094), .B1(n19936), .B2(n20090), .ZN(
        n19927) );
  INV_X1 U22933 ( .A(n19927), .ZN(n19929) );
  AOI22_X1 U22934 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19944), .B1(
        n20147), .B2(n19943), .ZN(n19928) );
  OAI211_X1 U22935 ( .C1(n20151), .C2(n19940), .A(n19929), .B(n19928), .ZN(
        P2_U3122) );
  OAI22_X1 U22936 ( .A1(n19947), .A2(n20096), .B1(n19936), .B2(n20095), .ZN(
        n19930) );
  INV_X1 U22937 ( .A(n19930), .ZN(n19932) );
  AOI22_X1 U22938 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19944), .B1(
        n20153), .B2(n19943), .ZN(n19931) );
  OAI211_X1 U22939 ( .C1(n20157), .C2(n19940), .A(n19932), .B(n19931), .ZN(
        P2_U3123) );
  NOR2_X1 U22940 ( .A1(n20100), .A2(n19936), .ZN(n19933) );
  AOI21_X1 U22941 ( .B1(n19974), .B2(n20021), .A(n19933), .ZN(n19935) );
  AOI22_X1 U22942 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19944), .B1(
        n20159), .B2(n19943), .ZN(n19934) );
  OAI211_X1 U22943 ( .C1(n20104), .C2(n19947), .A(n19935), .B(n19934), .ZN(
        P2_U3124) );
  OAI22_X1 U22944 ( .A1(n19947), .A2(n20171), .B1(n20105), .B2(n19936), .ZN(
        n19937) );
  INV_X1 U22945 ( .A(n19937), .ZN(n19939) );
  AOI22_X1 U22946 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19944), .B1(
        n20165), .B2(n19943), .ZN(n19938) );
  OAI211_X1 U22947 ( .C1(n20106), .C2(n19940), .A(n19939), .B(n19938), .ZN(
        P2_U3125) );
  AOI22_X1 U22948 ( .A1(n20025), .A2(n19974), .B1(n19953), .B2(n20172), .ZN(
        n19942) );
  AOI22_X1 U22949 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19944), .B1(
        n20173), .B2(n19943), .ZN(n19941) );
  OAI211_X1 U22950 ( .C1(n20111), .C2(n19947), .A(n19942), .B(n19941), .ZN(
        P2_U3126) );
  AOI22_X1 U22951 ( .A1(n19974), .A2(n20032), .B1(n19953), .B2(n20178), .ZN(
        n19946) );
  AOI22_X1 U22952 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19944), .B1(
        n20180), .B2(n19943), .ZN(n19945) );
  OAI211_X1 U22953 ( .C1(n20123), .C2(n19947), .A(n19946), .B(n19945), .ZN(
        P2_U3127) );
  NOR2_X1 U22954 ( .A1(n19979), .A2(n19949), .ZN(n19972) );
  OAI21_X1 U22955 ( .B1(n11052), .B2(n19972), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19950) );
  OAI21_X1 U22956 ( .B1(n19979), .B2(n19951), .A(n19950), .ZN(n19973) );
  AOI22_X1 U22957 ( .A1(n19973), .A2(n20127), .B1(n19972), .B2(n20126), .ZN(
        n19959) );
  INV_X1 U22958 ( .A(n11052), .ZN(n19956) );
  OR2_X1 U22959 ( .A1(n19974), .A2(n19952), .ZN(n19954) );
  AOI21_X1 U22960 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n19954), .A(n19953), 
        .ZN(n19955) );
  AOI211_X1 U22961 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19956), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19955), .ZN(n19957) );
  AOI22_X1 U22962 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19975), .B1(
        n19974), .B2(n20047), .ZN(n19958) );
  OAI211_X1 U22963 ( .C1(n20084), .C2(n20006), .A(n19959), .B(n19958), .ZN(
        P2_U3128) );
  AOI22_X1 U22964 ( .A1(n19973), .A2(n20141), .B1(n19972), .B2(n20140), .ZN(
        n19961) );
  AOI22_X1 U22965 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19975), .B1(
        n19974), .B2(n20050), .ZN(n19960) );
  OAI211_X1 U22966 ( .C1(n20089), .C2(n20006), .A(n19961), .B(n19960), .ZN(
        P2_U3129) );
  AOI22_X1 U22967 ( .A1(n19973), .A2(n20147), .B1(n19972), .B2(n20146), .ZN(
        n19963) );
  AOI22_X1 U22968 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19975), .B1(
        n19974), .B2(n20148), .ZN(n19962) );
  OAI211_X1 U22969 ( .C1(n20151), .C2(n20006), .A(n19963), .B(n19962), .ZN(
        P2_U3130) );
  AOI22_X1 U22970 ( .A1(n19973), .A2(n20153), .B1(n19972), .B2(n20152), .ZN(
        n19965) );
  AOI22_X1 U22971 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19975), .B1(
        n19974), .B2(n20154), .ZN(n19964) );
  OAI211_X1 U22972 ( .C1(n20157), .C2(n20006), .A(n19965), .B(n19964), .ZN(
        P2_U3131) );
  AOI22_X1 U22973 ( .A1(n19973), .A2(n20159), .B1(n19972), .B2(n20158), .ZN(
        n19967) );
  AOI22_X1 U22974 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19975), .B1(
        n19974), .B2(n20160), .ZN(n19966) );
  OAI211_X1 U22975 ( .C1(n20163), .C2(n20006), .A(n19967), .B(n19966), .ZN(
        P2_U3132) );
  AOI22_X1 U22976 ( .A1(n19973), .A2(n20165), .B1(n20164), .B2(n19972), .ZN(
        n19969) );
  AOI22_X1 U22977 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19975), .B1(
        n19974), .B2(n20059), .ZN(n19968) );
  OAI211_X1 U22978 ( .C1(n20106), .C2(n20006), .A(n19969), .B(n19968), .ZN(
        P2_U3133) );
  AOI22_X1 U22979 ( .A1(n19973), .A2(n20173), .B1(n19972), .B2(n20172), .ZN(
        n19971) );
  AOI22_X1 U22980 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19975), .B1(
        n19974), .B2(n20174), .ZN(n19970) );
  OAI211_X1 U22981 ( .C1(n20177), .C2(n20006), .A(n19971), .B(n19970), .ZN(
        P2_U3134) );
  AOI22_X1 U22982 ( .A1(n19973), .A2(n20180), .B1(n19972), .B2(n20178), .ZN(
        n19977) );
  AOI22_X1 U22983 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19975), .B1(
        n19974), .B2(n20182), .ZN(n19976) );
  OAI211_X1 U22984 ( .C1(n20188), .C2(n20006), .A(n19977), .B(n19976), .ZN(
        P2_U3135) );
  NOR2_X1 U22985 ( .A1(n19979), .A2(n19978), .ZN(n20001) );
  NAND2_X1 U22986 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19981), .ZN(
        n19983) );
  OAI21_X1 U22987 ( .B1(n19983), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20317), 
        .ZN(n19982) );
  AOI22_X1 U22988 ( .A1(n20002), .A2(n20127), .B1(n20126), .B2(n20001), .ZN(
        n19988) );
  OAI21_X1 U22989 ( .B1(n20132), .B2(n20271), .A(n19983), .ZN(n19985) );
  AND2_X1 U22990 ( .A1(n19985), .A2(n19984), .ZN(n19986) );
  OAI211_X1 U22991 ( .C1(n20001), .C2(n20306), .A(n19986), .B(n20133), .ZN(
        n20003) );
  AOI22_X1 U22992 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20003), .B1(
        n20031), .B2(n20136), .ZN(n19987) );
  OAI211_X1 U22993 ( .C1(n20139), .C2(n20006), .A(n19988), .B(n19987), .ZN(
        P2_U3136) );
  AOI22_X1 U22994 ( .A1(n20002), .A2(n20141), .B1(n20140), .B2(n20001), .ZN(
        n19990) );
  AOI22_X1 U22995 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20003), .B1(
        n20031), .B2(n20142), .ZN(n19989) );
  OAI211_X1 U22996 ( .C1(n20145), .C2(n20006), .A(n19990), .B(n19989), .ZN(
        P2_U3137) );
  AOI22_X1 U22997 ( .A1(n20002), .A2(n20147), .B1(n20146), .B2(n20001), .ZN(
        n19992) );
  AOI22_X1 U22998 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20003), .B1(
        n20031), .B2(n20013), .ZN(n19991) );
  OAI211_X1 U22999 ( .C1(n20094), .C2(n20006), .A(n19992), .B(n19991), .ZN(
        P2_U3138) );
  AOI22_X1 U23000 ( .A1(n20002), .A2(n20153), .B1(n20152), .B2(n20001), .ZN(
        n19994) );
  AOI22_X1 U23001 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20003), .B1(
        n20031), .B2(n20017), .ZN(n19993) );
  OAI211_X1 U23002 ( .C1(n20096), .C2(n20006), .A(n19994), .B(n19993), .ZN(
        P2_U3139) );
  AOI22_X1 U23003 ( .A1(n20002), .A2(n20159), .B1(n20158), .B2(n20001), .ZN(
        n19996) );
  AOI22_X1 U23004 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20003), .B1(
        n20031), .B2(n20021), .ZN(n19995) );
  OAI211_X1 U23005 ( .C1(n20104), .C2(n20006), .A(n19996), .B(n19995), .ZN(
        P2_U3140) );
  AOI22_X1 U23006 ( .A1(n20002), .A2(n20165), .B1(n20164), .B2(n20001), .ZN(
        n19998) );
  AOI22_X1 U23007 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20003), .B1(
        n20031), .B2(n20166), .ZN(n19997) );
  OAI211_X1 U23008 ( .C1(n20171), .C2(n20006), .A(n19998), .B(n19997), .ZN(
        P2_U3141) );
  AOI22_X1 U23009 ( .A1(n20002), .A2(n20173), .B1(n20172), .B2(n20001), .ZN(
        n20000) );
  AOI22_X1 U23010 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20003), .B1(
        n20031), .B2(n20025), .ZN(n19999) );
  OAI211_X1 U23011 ( .C1(n20111), .C2(n20006), .A(n20000), .B(n19999), .ZN(
        P2_U3142) );
  AOI22_X1 U23012 ( .A1(n20002), .A2(n20180), .B1(n20178), .B2(n20001), .ZN(
        n20005) );
  AOI22_X1 U23013 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20003), .B1(
        n20031), .B2(n20032), .ZN(n20004) );
  OAI211_X1 U23014 ( .C1(n20123), .C2(n20006), .A(n20005), .B(n20004), .ZN(
        P2_U3143) );
  INV_X1 U23015 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n20009) );
  AOI22_X1 U23016 ( .A1(n20030), .A2(n20127), .B1(n20029), .B2(n20126), .ZN(
        n20008) );
  AOI22_X1 U23017 ( .A1(n20031), .A2(n20047), .B1(n20065), .B2(n20136), .ZN(
        n20007) );
  OAI211_X1 U23018 ( .C1(n20035), .C2(n20009), .A(n20008), .B(n20007), .ZN(
        P2_U3144) );
  INV_X1 U23019 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n20012) );
  AOI22_X1 U23020 ( .A1(n20030), .A2(n20141), .B1(n20029), .B2(n20140), .ZN(
        n20011) );
  AOI22_X1 U23021 ( .A1(n20065), .A2(n20142), .B1(n20031), .B2(n20050), .ZN(
        n20010) );
  OAI211_X1 U23022 ( .C1(n20035), .C2(n20012), .A(n20011), .B(n20010), .ZN(
        P2_U3145) );
  INV_X1 U23023 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n20016) );
  AOI22_X1 U23024 ( .A1(n20030), .A2(n20147), .B1(n20029), .B2(n20146), .ZN(
        n20015) );
  AOI22_X1 U23025 ( .A1(n20065), .A2(n20013), .B1(n20031), .B2(n20148), .ZN(
        n20014) );
  OAI211_X1 U23026 ( .C1(n20035), .C2(n20016), .A(n20015), .B(n20014), .ZN(
        P2_U3146) );
  INV_X1 U23027 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n20020) );
  AOI22_X1 U23028 ( .A1(n20030), .A2(n20153), .B1(n20029), .B2(n20152), .ZN(
        n20019) );
  AOI22_X1 U23029 ( .A1(n20031), .A2(n20154), .B1(n20065), .B2(n20017), .ZN(
        n20018) );
  OAI211_X1 U23030 ( .C1(n20035), .C2(n20020), .A(n20019), .B(n20018), .ZN(
        P2_U3147) );
  INV_X1 U23031 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n20024) );
  AOI22_X1 U23032 ( .A1(n20030), .A2(n20159), .B1(n20029), .B2(n20158), .ZN(
        n20023) );
  AOI22_X1 U23033 ( .A1(n20065), .A2(n20021), .B1(n20031), .B2(n20160), .ZN(
        n20022) );
  OAI211_X1 U23034 ( .C1(n20035), .C2(n20024), .A(n20023), .B(n20022), .ZN(
        P2_U3148) );
  INV_X1 U23035 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n20028) );
  AOI22_X1 U23036 ( .A1(n20030), .A2(n20173), .B1(n20029), .B2(n20172), .ZN(
        n20027) );
  AOI22_X1 U23037 ( .A1(n20031), .A2(n20174), .B1(n20065), .B2(n20025), .ZN(
        n20026) );
  OAI211_X1 U23038 ( .C1(n20035), .C2(n20028), .A(n20027), .B(n20026), .ZN(
        P2_U3150) );
  AOI22_X1 U23039 ( .A1(n20030), .A2(n20180), .B1(n20029), .B2(n20178), .ZN(
        n20034) );
  AOI22_X1 U23040 ( .A1(n20065), .A2(n20032), .B1(n20031), .B2(n20182), .ZN(
        n20033) );
  OAI211_X1 U23041 ( .C1(n20035), .C2(n10591), .A(n20034), .B(n20033), .ZN(
        P2_U3151) );
  INV_X1 U23042 ( .A(n20043), .ZN(n20036) );
  NAND2_X1 U23043 ( .A1(n20040), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20075) );
  AND2_X1 U23044 ( .A1(n20075), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20038) );
  NAND2_X1 U23045 ( .A1(n20039), .A2(n20038), .ZN(n20045) );
  INV_X1 U23046 ( .A(n20040), .ZN(n20042) );
  OAI21_X1 U23047 ( .B1(n20042), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20317), 
        .ZN(n20041) );
  INV_X1 U23048 ( .A(n20075), .ZN(n20078) );
  AOI22_X1 U23049 ( .A1(n20064), .A2(n20127), .B1(n20078), .B2(n20126), .ZN(
        n20049) );
  OAI21_X1 U23050 ( .B1(n20132), .B2(n20043), .A(n20042), .ZN(n20046) );
  NAND2_X1 U23051 ( .A1(n20075), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20044) );
  NAND4_X1 U23052 ( .A1(n20046), .A2(n20133), .A3(n20045), .A4(n20044), .ZN(
        n20066) );
  AOI22_X1 U23053 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20066), .B1(
        n20065), .B2(n20047), .ZN(n20048) );
  OAI211_X1 U23054 ( .C1(n20084), .C2(n20122), .A(n20049), .B(n20048), .ZN(
        P2_U3152) );
  AOI22_X1 U23055 ( .A1(n20064), .A2(n20141), .B1(n20078), .B2(n20140), .ZN(
        n20052) );
  AOI22_X1 U23056 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20066), .B1(
        n20065), .B2(n20050), .ZN(n20051) );
  OAI211_X1 U23057 ( .C1(n20089), .C2(n20122), .A(n20052), .B(n20051), .ZN(
        P2_U3153) );
  AOI22_X1 U23058 ( .A1(n20064), .A2(n20147), .B1(n20078), .B2(n20146), .ZN(
        n20054) );
  AOI22_X1 U23059 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20066), .B1(
        n20065), .B2(n20148), .ZN(n20053) );
  OAI211_X1 U23060 ( .C1(n20151), .C2(n20122), .A(n20054), .B(n20053), .ZN(
        P2_U3154) );
  AOI22_X1 U23061 ( .A1(n20064), .A2(n20153), .B1(n20078), .B2(n20152), .ZN(
        n20056) );
  AOI22_X1 U23062 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20066), .B1(
        n20065), .B2(n20154), .ZN(n20055) );
  OAI211_X1 U23063 ( .C1(n20157), .C2(n20122), .A(n20056), .B(n20055), .ZN(
        P2_U3155) );
  AOI22_X1 U23064 ( .A1(n20064), .A2(n20159), .B1(n20078), .B2(n20158), .ZN(
        n20058) );
  AOI22_X1 U23065 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20066), .B1(
        n20065), .B2(n20160), .ZN(n20057) );
  OAI211_X1 U23066 ( .C1(n20163), .C2(n20122), .A(n20058), .B(n20057), .ZN(
        P2_U3156) );
  AOI22_X1 U23067 ( .A1(n20064), .A2(n20165), .B1(n20164), .B2(n20078), .ZN(
        n20061) );
  AOI22_X1 U23068 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20066), .B1(
        n20065), .B2(n20059), .ZN(n20060) );
  OAI211_X1 U23069 ( .C1(n20106), .C2(n20122), .A(n20061), .B(n20060), .ZN(
        P2_U3157) );
  AOI22_X1 U23070 ( .A1(n20064), .A2(n20173), .B1(n20078), .B2(n20172), .ZN(
        n20063) );
  AOI22_X1 U23071 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20066), .B1(
        n20065), .B2(n20174), .ZN(n20062) );
  OAI211_X1 U23072 ( .C1(n20177), .C2(n20122), .A(n20063), .B(n20062), .ZN(
        P2_U3158) );
  AOI22_X1 U23073 ( .A1(n20064), .A2(n20180), .B1(n20078), .B2(n20178), .ZN(
        n20068) );
  AOI22_X1 U23074 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20066), .B1(
        n20065), .B2(n20182), .ZN(n20067) );
  OAI211_X1 U23075 ( .C1(n20188), .C2(n20122), .A(n20068), .B(n20067), .ZN(
        P2_U3159) );
  NOR3_X1 U23076 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20284), .A3(
        n20130), .ZN(n20079) );
  INV_X1 U23077 ( .A(n20079), .ZN(n20115) );
  OAI22_X1 U23078 ( .A1(n20122), .A2(n20139), .B1(n20071), .B2(n20115), .ZN(
        n20072) );
  INV_X1 U23079 ( .A(n20072), .ZN(n20083) );
  AOI21_X1 U23080 ( .B1(n20170), .B2(n20122), .A(n20272), .ZN(n20073) );
  NOR2_X1 U23081 ( .A1(n20073), .A2(n20268), .ZN(n20077) );
  OAI21_X1 U23082 ( .B1(n11057), .B2(n20317), .A(n20306), .ZN(n20074) );
  AOI21_X1 U23083 ( .B1(n20077), .B2(n20075), .A(n20074), .ZN(n20076) );
  OAI21_X2 U23084 ( .B1(n20076), .B2(n20079), .A(n20133), .ZN(n20119) );
  OAI21_X1 U23085 ( .B1(n20079), .B2(n20078), .A(n20077), .ZN(n20081) );
  OAI21_X1 U23086 ( .B1(n11057), .B2(n20079), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20080) );
  AOI22_X1 U23087 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20119), .B1(
        n20127), .B2(n20118), .ZN(n20082) );
  OAI211_X1 U23088 ( .C1(n20084), .C2(n20170), .A(n20083), .B(n20082), .ZN(
        P2_U3160) );
  OAI22_X1 U23089 ( .A1(n20122), .A2(n20145), .B1(n20085), .B2(n20115), .ZN(
        n20086) );
  INV_X1 U23090 ( .A(n20086), .ZN(n20088) );
  AOI22_X1 U23091 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20119), .B1(
        n20141), .B2(n20118), .ZN(n20087) );
  OAI211_X1 U23092 ( .C1(n20089), .C2(n20170), .A(n20088), .B(n20087), .ZN(
        P2_U3161) );
  OAI22_X1 U23093 ( .A1(n20170), .A2(n20151), .B1(n20090), .B2(n20115), .ZN(
        n20091) );
  INV_X1 U23094 ( .A(n20091), .ZN(n20093) );
  AOI22_X1 U23095 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20119), .B1(
        n20147), .B2(n20118), .ZN(n20092) );
  OAI211_X1 U23096 ( .C1(n20094), .C2(n20122), .A(n20093), .B(n20092), .ZN(
        P2_U3162) );
  OAI22_X1 U23097 ( .A1(n20122), .A2(n20096), .B1(n20095), .B2(n20115), .ZN(
        n20097) );
  INV_X1 U23098 ( .A(n20097), .ZN(n20099) );
  AOI22_X1 U23099 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20119), .B1(
        n20153), .B2(n20118), .ZN(n20098) );
  OAI211_X1 U23100 ( .C1(n20157), .C2(n20170), .A(n20099), .B(n20098), .ZN(
        P2_U3163) );
  OAI22_X1 U23101 ( .A1(n20170), .A2(n20163), .B1(n20100), .B2(n20115), .ZN(
        n20101) );
  INV_X1 U23102 ( .A(n20101), .ZN(n20103) );
  AOI22_X1 U23103 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20119), .B1(
        n20159), .B2(n20118), .ZN(n20102) );
  OAI211_X1 U23104 ( .C1(n20104), .C2(n20122), .A(n20103), .B(n20102), .ZN(
        P2_U3164) );
  OAI22_X1 U23105 ( .A1(n20170), .A2(n20106), .B1(n20105), .B2(n20115), .ZN(
        n20107) );
  INV_X1 U23106 ( .A(n20107), .ZN(n20109) );
  AOI22_X1 U23107 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20119), .B1(
        n20165), .B2(n20118), .ZN(n20108) );
  OAI211_X1 U23108 ( .C1(n20171), .C2(n20122), .A(n20109), .B(n20108), .ZN(
        P2_U3165) );
  OAI22_X1 U23109 ( .A1(n20122), .A2(n20111), .B1(n20115), .B2(n20110), .ZN(
        n20112) );
  INV_X1 U23110 ( .A(n20112), .ZN(n20114) );
  AOI22_X1 U23111 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20119), .B1(
        n20173), .B2(n20118), .ZN(n20113) );
  OAI211_X1 U23112 ( .C1(n20177), .C2(n20170), .A(n20114), .B(n20113), .ZN(
        P2_U3166) );
  OAI22_X1 U23113 ( .A1(n20170), .A2(n20188), .B1(n20116), .B2(n20115), .ZN(
        n20117) );
  INV_X1 U23114 ( .A(n20117), .ZN(n20121) );
  AOI22_X1 U23115 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20119), .B1(
        n20180), .B2(n20118), .ZN(n20120) );
  OAI211_X1 U23116 ( .C1(n20123), .C2(n20122), .A(n20121), .B(n20120), .ZN(
        P2_U3167) );
  OR2_X1 U23117 ( .A1(n20284), .A2(n20130), .ZN(n20125) );
  OAI21_X1 U23118 ( .B1(n20128), .B2(n20179), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20124) );
  OAI21_X1 U23119 ( .B1(n20125), .B2(n20268), .A(n20124), .ZN(n20181) );
  AOI22_X1 U23120 ( .A1(n20181), .A2(n20127), .B1(n20179), .B2(n20126), .ZN(
        n20138) );
  INV_X1 U23121 ( .A(n20128), .ZN(n20129) );
  AOI21_X1 U23122 ( .B1(n20129), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20135) );
  OAI22_X1 U23123 ( .A1(n20132), .A2(n20131), .B1(n20130), .B2(n20284), .ZN(
        n20134) );
  OAI211_X1 U23124 ( .C1(n20179), .C2(n20135), .A(n20134), .B(n20133), .ZN(
        n20184) );
  AOI22_X1 U23125 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20184), .B1(
        n20167), .B2(n20136), .ZN(n20137) );
  OAI211_X1 U23126 ( .C1(n20139), .C2(n20170), .A(n20138), .B(n20137), .ZN(
        P2_U3168) );
  AOI22_X1 U23127 ( .A1(n20181), .A2(n20141), .B1(n20179), .B2(n20140), .ZN(
        n20144) );
  AOI22_X1 U23128 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20184), .B1(
        n20167), .B2(n20142), .ZN(n20143) );
  OAI211_X1 U23129 ( .C1(n20145), .C2(n20170), .A(n20144), .B(n20143), .ZN(
        P2_U3169) );
  AOI22_X1 U23130 ( .A1(n20181), .A2(n20147), .B1(n20179), .B2(n20146), .ZN(
        n20150) );
  INV_X1 U23131 ( .A(n20170), .ZN(n20183) );
  AOI22_X1 U23132 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20184), .B1(
        n20183), .B2(n20148), .ZN(n20149) );
  OAI211_X1 U23133 ( .C1(n20151), .C2(n20187), .A(n20150), .B(n20149), .ZN(
        P2_U3170) );
  AOI22_X1 U23134 ( .A1(n20181), .A2(n20153), .B1(n20179), .B2(n20152), .ZN(
        n20156) );
  AOI22_X1 U23135 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20184), .B1(
        n20183), .B2(n20154), .ZN(n20155) );
  OAI211_X1 U23136 ( .C1(n20157), .C2(n20187), .A(n20156), .B(n20155), .ZN(
        P2_U3171) );
  AOI22_X1 U23137 ( .A1(n20181), .A2(n20159), .B1(n20179), .B2(n20158), .ZN(
        n20162) );
  AOI22_X1 U23138 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20184), .B1(
        n20183), .B2(n20160), .ZN(n20161) );
  OAI211_X1 U23139 ( .C1(n20163), .C2(n20187), .A(n20162), .B(n20161), .ZN(
        P2_U3172) );
  AOI22_X1 U23140 ( .A1(n20181), .A2(n20165), .B1(n20179), .B2(n20164), .ZN(
        n20169) );
  AOI22_X1 U23141 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20184), .B1(
        n20167), .B2(n20166), .ZN(n20168) );
  OAI211_X1 U23142 ( .C1(n20171), .C2(n20170), .A(n20169), .B(n20168), .ZN(
        P2_U3173) );
  AOI22_X1 U23143 ( .A1(n20181), .A2(n20173), .B1(n20179), .B2(n20172), .ZN(
        n20176) );
  AOI22_X1 U23144 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20184), .B1(
        n20183), .B2(n20174), .ZN(n20175) );
  OAI211_X1 U23145 ( .C1(n20177), .C2(n20187), .A(n20176), .B(n20175), .ZN(
        P2_U3174) );
  AOI22_X1 U23146 ( .A1(n20181), .A2(n20180), .B1(n20179), .B2(n20178), .ZN(
        n20186) );
  AOI22_X1 U23147 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20184), .B1(
        n20183), .B2(n20182), .ZN(n20185) );
  OAI211_X1 U23148 ( .C1(n20188), .C2(n20187), .A(n20186), .B(n20185), .ZN(
        P2_U3175) );
  AND2_X1 U23149 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n20189), .ZN(
        P2_U3179) );
  AND2_X1 U23150 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n20189), .ZN(
        P2_U3180) );
  AND2_X1 U23151 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n20189), .ZN(
        P2_U3181) );
  AND2_X1 U23152 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n20189), .ZN(
        P2_U3182) );
  AND2_X1 U23153 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n20189), .ZN(
        P2_U3183) );
  AND2_X1 U23154 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20189), .ZN(
        P2_U3184) );
  AND2_X1 U23155 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n20189), .ZN(
        P2_U3185) );
  AND2_X1 U23156 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n20189), .ZN(
        P2_U3186) );
  AND2_X1 U23157 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20189), .ZN(
        P2_U3187) );
  AND2_X1 U23158 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n20189), .ZN(
        P2_U3188) );
  AND2_X1 U23159 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20189), .ZN(
        P2_U3189) );
  AND2_X1 U23160 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20189), .ZN(
        P2_U3190) );
  AND2_X1 U23161 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20189), .ZN(
        P2_U3191) );
  AND2_X1 U23162 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n20189), .ZN(
        P2_U3192) );
  AND2_X1 U23163 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n20189), .ZN(
        P2_U3193) );
  AND2_X1 U23164 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n20189), .ZN(
        P2_U3194) );
  AND2_X1 U23165 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n20189), .ZN(
        P2_U3195) );
  AND2_X1 U23166 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n20189), .ZN(
        P2_U3196) );
  AND2_X1 U23167 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n20189), .ZN(
        P2_U3197) );
  AND2_X1 U23168 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n20189), .ZN(
        P2_U3198) );
  AND2_X1 U23169 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n20189), .ZN(
        P2_U3199) );
  AND2_X1 U23170 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n20189), .ZN(
        P2_U3200) );
  AND2_X1 U23171 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n20189), .ZN(P2_U3201) );
  AND2_X1 U23172 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n20189), .ZN(P2_U3202) );
  AND2_X1 U23173 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n20189), .ZN(P2_U3203) );
  AND2_X1 U23174 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20189), .ZN(P2_U3204) );
  AND2_X1 U23175 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n20189), .ZN(P2_U3205) );
  AND2_X1 U23176 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n20189), .ZN(P2_U3206) );
  AND2_X1 U23177 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n20189), .ZN(P2_U3207) );
  AND2_X1 U23178 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n20189), .ZN(P2_U3208) );
  OAI21_X1 U23179 ( .B1(n21141), .B2(n20196), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n20207) );
  INV_X1 U23180 ( .A(n20207), .ZN(n20194) );
  NOR2_X1 U23181 ( .A1(n20191), .A2(n20190), .ZN(n20201) );
  INV_X1 U23182 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20324) );
  NOR3_X1 U23183 ( .A1(n20201), .A2(n20324), .A3(n20195), .ZN(n20193) );
  OAI211_X1 U23184 ( .C1(HOLD), .C2(n20324), .A(n20326), .B(n20202), .ZN(
        n20192) );
  OAI21_X1 U23185 ( .B1(n20194), .B2(n20193), .A(n20192), .ZN(P2_U3209) );
  NOR2_X1 U23186 ( .A1(n20313), .A2(n20201), .ZN(n20198) );
  NOR2_X1 U23187 ( .A1(HOLD), .A2(n20195), .ZN(n20206) );
  OAI211_X1 U23188 ( .C1(n20206), .C2(n20208), .A(
        P2_REQUESTPENDING_REG_SCAN_IN), .B(n20196), .ZN(n20197) );
  OAI211_X1 U23189 ( .C1(n20200), .C2(n20199), .A(n20198), .B(n20197), .ZN(
        P2_U3210) );
  INV_X1 U23190 ( .A(n20201), .ZN(n20205) );
  OAI22_X1 U23191 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n20202), .B1(NA), 
        .B2(n20205), .ZN(n20203) );
  OAI211_X1 U23192 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n20203), .ZN(n20204) );
  OAI221_X1 U23193 ( .B1(n20207), .B2(n20206), .C1(n20207), .C2(n20205), .A(
        n20204), .ZN(P2_U3211) );
  OAI222_X1 U23194 ( .A1(n20258), .A2(n20211), .B1(n20209), .B2(n20260), .C1(
        n10958), .C2(n20259), .ZN(P2_U3212) );
  OAI222_X1 U23195 ( .A1(n20259), .A2(n20211), .B1(n20210), .B2(n20260), .C1(
        n17201), .C2(n20258), .ZN(P2_U3213) );
  OAI222_X1 U23196 ( .A1(n20259), .A2(n17201), .B1(n20212), .B2(n20260), .C1(
        n11300), .C2(n20258), .ZN(P2_U3214) );
  OAI222_X1 U23197 ( .A1(n20258), .A2(n15920), .B1(n20213), .B2(n20260), .C1(
        n11300), .C2(n20259), .ZN(P2_U3215) );
  OAI222_X1 U23198 ( .A1(n20258), .A2(n20215), .B1(n20214), .B2(n20260), .C1(
        n15920), .C2(n20259), .ZN(P2_U3216) );
  OAI222_X1 U23199 ( .A1(n20258), .A2(n20217), .B1(n20216), .B2(n20260), .C1(
        n20215), .C2(n20259), .ZN(P2_U3217) );
  INV_X2 U23200 ( .A(n20326), .ZN(n20260) );
  OAI222_X1 U23201 ( .A1(n20258), .A2(n20219), .B1(n20218), .B2(n20260), .C1(
        n20217), .C2(n20259), .ZN(P2_U3218) );
  INV_X1 U23202 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n20221) );
  OAI222_X1 U23203 ( .A1(n20258), .A2(n20221), .B1(n20220), .B2(n20260), .C1(
        n20219), .C2(n20259), .ZN(P2_U3219) );
  OAI222_X1 U23204 ( .A1(n20258), .A2(n20223), .B1(n20222), .B2(n20260), .C1(
        n20221), .C2(n20259), .ZN(P2_U3220) );
  OAI222_X1 U23205 ( .A1(n20258), .A2(n16343), .B1(n20224), .B2(n20260), .C1(
        n20223), .C2(n20259), .ZN(P2_U3221) );
  OAI222_X1 U23206 ( .A1(n20258), .A2(n20226), .B1(n20225), .B2(n20260), .C1(
        n16343), .C2(n20259), .ZN(P2_U3222) );
  OAI222_X1 U23207 ( .A1(n20258), .A2(n20228), .B1(n20227), .B2(n20260), .C1(
        n20226), .C2(n20259), .ZN(P2_U3223) );
  OAI222_X1 U23208 ( .A1(n20258), .A2(n20230), .B1(n20229), .B2(n20260), .C1(
        n20228), .C2(n20259), .ZN(P2_U3224) );
  OAI222_X1 U23209 ( .A1(n20258), .A2(n11340), .B1(n20231), .B2(n20260), .C1(
        n20230), .C2(n20259), .ZN(P2_U3225) );
  OAI222_X1 U23210 ( .A1(n20258), .A2(n20233), .B1(n20232), .B2(n20260), .C1(
        n11340), .C2(n20259), .ZN(P2_U3226) );
  OAI222_X1 U23211 ( .A1(n20258), .A2(n20235), .B1(n20234), .B2(n20260), .C1(
        n20233), .C2(n20259), .ZN(P2_U3227) );
  OAI222_X1 U23212 ( .A1(n20258), .A2(n20237), .B1(n20236), .B2(n20260), .C1(
        n20235), .C2(n20259), .ZN(P2_U3228) );
  OAI222_X1 U23213 ( .A1(n20258), .A2(n20239), .B1(n20238), .B2(n20260), .C1(
        n20237), .C2(n20259), .ZN(P2_U3229) );
  OAI222_X1 U23214 ( .A1(n20258), .A2(n20241), .B1(n20240), .B2(n20260), .C1(
        n20239), .C2(n20259), .ZN(P2_U3230) );
  INV_X1 U23215 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20243) );
  OAI222_X1 U23216 ( .A1(n20258), .A2(n20243), .B1(n20242), .B2(n20260), .C1(
        n20241), .C2(n20259), .ZN(P2_U3231) );
  OAI222_X1 U23217 ( .A1(n20258), .A2(n20245), .B1(n20244), .B2(n20260), .C1(
        n20243), .C2(n20259), .ZN(P2_U3232) );
  OAI222_X1 U23218 ( .A1(n20258), .A2(n11369), .B1(n20246), .B2(n20260), .C1(
        n20245), .C2(n20259), .ZN(P2_U3233) );
  OAI222_X1 U23219 ( .A1(n20258), .A2(n20248), .B1(n20247), .B2(n20260), .C1(
        n11369), .C2(n20259), .ZN(P2_U3234) );
  OAI222_X1 U23220 ( .A1(n20258), .A2(n11377), .B1(n20249), .B2(n20260), .C1(
        n20248), .C2(n20259), .ZN(P2_U3235) );
  INV_X1 U23221 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20251) );
  OAI222_X1 U23222 ( .A1(n20258), .A2(n20251), .B1(n20250), .B2(n20260), .C1(
        n11377), .C2(n20259), .ZN(P2_U3236) );
  OAI222_X1 U23223 ( .A1(n20258), .A2(n11386), .B1(n20252), .B2(n20260), .C1(
        n20251), .C2(n20259), .ZN(P2_U3237) );
  OAI222_X1 U23224 ( .A1(n20259), .A2(n11386), .B1(n20253), .B2(n20260), .C1(
        n20254), .C2(n20258), .ZN(P2_U3238) );
  INV_X1 U23225 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20256) );
  OAI222_X1 U23226 ( .A1(n20258), .A2(n20256), .B1(n20255), .B2(n20260), .C1(
        n20254), .C2(n20259), .ZN(P2_U3239) );
  OAI222_X1 U23227 ( .A1(n20258), .A2(n11480), .B1(n20257), .B2(n20260), .C1(
        n20256), .C2(n20259), .ZN(P2_U3240) );
  OAI222_X1 U23228 ( .A1(n20258), .A2(n11403), .B1(n20261), .B2(n20260), .C1(
        n11480), .C2(n20259), .ZN(P2_U3241) );
  OAI22_X1 U23229 ( .A1(n20326), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n20260), .ZN(n20262) );
  INV_X1 U23230 ( .A(n20262), .ZN(P2_U3585) );
  MUX2_X1 U23231 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n20326), .Z(P2_U3586) );
  MUX2_X1 U23232 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .B(P2_BE_N_REG_1__SCAN_IN), .S(n20326), .Z(P2_U3587) );
  OAI22_X1 U23233 ( .A1(n20326), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n20260), .ZN(n20263) );
  INV_X1 U23234 ( .A(n20263), .ZN(P2_U3588) );
  OAI21_X1 U23235 ( .B1(n20267), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20265), 
        .ZN(n20264) );
  INV_X1 U23236 ( .A(n20264), .ZN(P2_U3591) );
  OAI21_X1 U23237 ( .B1(n20267), .B2(n20266), .A(n20265), .ZN(P2_U3592) );
  OR2_X1 U23238 ( .A1(n20269), .A2(n20268), .ZN(n20282) );
  OR2_X1 U23239 ( .A1(n20271), .A2(n20270), .ZN(n20285) );
  OR2_X1 U23240 ( .A1(n20273), .A2(n20272), .ZN(n20274) );
  OR2_X1 U23241 ( .A1(n20275), .A2(n20274), .ZN(n20277) );
  NAND2_X1 U23242 ( .A1(n20277), .A2(n20276), .ZN(n20287) );
  NAND2_X1 U23243 ( .A1(n20285), .A2(n20287), .ZN(n20279) );
  AOI22_X1 U23244 ( .A1(n20280), .A2(n20279), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20278), .ZN(n20281) );
  AND2_X1 U23245 ( .A1(n20282), .A2(n20281), .ZN(n20283) );
  AOI22_X1 U23246 ( .A1(n20294), .A2(n20284), .B1(n20283), .B2(n20291), .ZN(
        P2_U3602) );
  INV_X1 U23247 ( .A(n20285), .ZN(n20290) );
  OAI22_X1 U23248 ( .A1(n20288), .A2(n20287), .B1(n20286), .B2(n20306), .ZN(
        n20289) );
  NOR2_X1 U23249 ( .A1(n20290), .A2(n20289), .ZN(n20292) );
  AOI22_X1 U23250 ( .A1(n20294), .A2(n20293), .B1(n20292), .B2(n20291), .ZN(
        P2_U3603) );
  INV_X1 U23251 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20295) );
  AOI22_X1 U23252 ( .A1(n20260), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20295), 
        .B2(n20326), .ZN(P2_U3608) );
  INV_X1 U23253 ( .A(n20296), .ZN(n20300) );
  AOI22_X1 U23254 ( .A1(n20300), .A2(n20299), .B1(n20298), .B2(n20297), .ZN(
        n20302) );
  NAND2_X1 U23255 ( .A1(n20302), .A2(n20301), .ZN(n20304) );
  MUX2_X1 U23256 ( .A(P2_MORE_REG_SCAN_IN), .B(n20304), .S(n20303), .Z(
        P2_U3609) );
  AOI21_X1 U23257 ( .B1(n20307), .B2(n20306), .A(n20305), .ZN(n20308) );
  OAI211_X1 U23258 ( .C1(n20318), .C2(n20310), .A(n20309), .B(n20308), .ZN(
        n20325) );
  NOR3_X1 U23259 ( .A1(n20313), .A2(n20311), .A3(n13438), .ZN(n20316) );
  AOI21_X1 U23260 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n20313), .A(n20312), 
        .ZN(n20315) );
  MUX2_X1 U23261 ( .A(n20316), .B(n20315), .S(n20314), .Z(n20322) );
  OAI22_X1 U23262 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20319), .B1(n20318), 
        .B2(n20317), .ZN(n20320) );
  INV_X1 U23263 ( .A(n20320), .ZN(n20321) );
  OAI21_X1 U23264 ( .B1(n20322), .B2(n20321), .A(n20325), .ZN(n20323) );
  OAI21_X1 U23265 ( .B1(n20325), .B2(n20324), .A(n20323), .ZN(P2_U3610) );
  OAI22_X1 U23266 ( .A1(n20326), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n20260), .ZN(n20327) );
  INV_X1 U23267 ( .A(n20327), .ZN(P2_U3611) );
  NOR2_X1 U23268 ( .A1(n21150), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20336) );
  NOR2_X1 U23269 ( .A1(n20336), .A2(n21137), .ZN(n20329) );
  INV_X1 U23270 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n20328) );
  NAND2_X2 U23271 ( .A1(n21137), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n21198) );
  AOI21_X1 U23272 ( .B1(n20329), .B2(n20328), .A(n21214), .ZN(P1_U2802) );
  NAND2_X1 U23273 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21070), .ZN(n20334) );
  OAI21_X1 U23274 ( .B1(n20331), .B2(n20330), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20332) );
  OAI21_X1 U23275 ( .B1(n20334), .B2(n20333), .A(n20332), .ZN(P1_U2803) );
  NOR2_X1 U23276 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20337) );
  OAI21_X1 U23277 ( .B1(n20337), .B2(P1_D_C_N_REG_SCAN_IN), .A(n21198), .ZN(
        n20335) );
  OAI21_X1 U23278 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n21198), .A(n20335), 
        .ZN(P1_U2804) );
  OAI21_X2 U23279 ( .B1(n21137), .B2(n20336), .A(n21198), .ZN(n21136) );
  OAI21_X1 U23280 ( .B1(BS16), .B2(n20337), .A(n21204), .ZN(n21202) );
  OAI21_X1 U23281 ( .B1(n21204), .B2(n21022), .A(n21202), .ZN(P1_U2805) );
  OAI21_X1 U23282 ( .B1(n20340), .B2(n20339), .A(n20338), .ZN(P1_U2806) );
  NOR4_X1 U23283 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20344) );
  NOR4_X1 U23284 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_15__SCAN_IN), .A3(P1_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20343) );
  NOR4_X1 U23285 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .A3(P1_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n20342) );
  NOR4_X1 U23286 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20341) );
  NAND4_X1 U23287 ( .A1(n20344), .A2(n20343), .A3(n20342), .A4(n20341), .ZN(
        n20350) );
  NOR4_X1 U23288 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_2__SCAN_IN), .A3(P1_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_5__SCAN_IN), .ZN(n20348) );
  AOI211_X1 U23289 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_12__SCAN_IN), .B(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n20347) );
  NOR4_X1 U23290 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_11__SCAN_IN), .A3(P1_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n20346) );
  NOR4_X1 U23291 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_7__SCAN_IN), .A3(P1_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_9__SCAN_IN), .ZN(n20345) );
  NAND4_X1 U23292 ( .A1(n20348), .A2(n20347), .A3(n20346), .A4(n20345), .ZN(
        n20349) );
  NOR2_X1 U23293 ( .A1(n20350), .A2(n20349), .ZN(n21212) );
  INV_X1 U23294 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20352) );
  NOR3_X1 U23295 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20353) );
  OAI21_X1 U23296 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20353), .A(n21212), .ZN(
        n20351) );
  OAI21_X1 U23297 ( .B1(n21212), .B2(n20352), .A(n20351), .ZN(P1_U2807) );
  INV_X1 U23298 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21203) );
  AOI21_X1 U23299 ( .B1(n21206), .B2(n21203), .A(n20353), .ZN(n20355) );
  INV_X1 U23300 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20354) );
  INV_X1 U23301 ( .A(n21212), .ZN(n21209) );
  AOI22_X1 U23302 ( .A1(n21212), .A2(n20355), .B1(n20354), .B2(n21209), .ZN(
        P1_U2808) );
  OAI22_X1 U23303 ( .A1(n20432), .A2(n20357), .B1(n20356), .B2(
        P1_REIP_REG_9__SCAN_IN), .ZN(n20358) );
  INV_X1 U23304 ( .A(n20358), .ZN(n20365) );
  AOI22_X1 U23305 ( .A1(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n20427), .B1(
        P1_REIP_REG_9__SCAN_IN), .B2(n20371), .ZN(n20364) );
  AOI21_X1 U23306 ( .B1(n20405), .B2(P1_EBX_REG_9__SCAN_IN), .A(n20368), .ZN(
        n20363) );
  INV_X1 U23307 ( .A(n20359), .ZN(n20360) );
  AOI22_X1 U23308 ( .A1(n20361), .A2(n20383), .B1(n10405), .B2(n20360), .ZN(
        n20362) );
  NAND4_X1 U23309 ( .A1(n20365), .A2(n20364), .A3(n20363), .A4(n20362), .ZN(
        P1_U2831) );
  AOI22_X1 U23310 ( .A1(n20438), .A2(n20404), .B1(n20405), .B2(
        P1_EBX_REG_8__SCAN_IN), .ZN(n20375) );
  NOR3_X1 U23311 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n20420), .A3(n20366), .ZN(
        n20367) );
  AOI211_X1 U23312 ( .C1(n20427), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n20368), .B(n20367), .ZN(n20374) );
  INV_X1 U23313 ( .A(n20369), .ZN(n20370) );
  AOI22_X1 U23314 ( .A1(n20441), .A2(n20383), .B1(n10405), .B2(n20370), .ZN(
        n20373) );
  NAND2_X1 U23315 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n20371), .ZN(n20372) );
  NAND4_X1 U23316 ( .A1(n20375), .A2(n20374), .A3(n20373), .A4(n20372), .ZN(
        P1_U2832) );
  NAND2_X1 U23317 ( .A1(n20376), .A2(n20396), .ZN(n20377) );
  OR2_X1 U23318 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20377), .ZN(n20378) );
  OAI211_X1 U23319 ( .C1(n20407), .C2(n12605), .A(n20421), .B(n20378), .ZN(
        n20381) );
  NOR2_X1 U23320 ( .A1(n20432), .A2(n20379), .ZN(n20380) );
  AOI211_X1 U23321 ( .C1(P1_EBX_REG_7__SCAN_IN), .C2(n20405), .A(n20381), .B(
        n20380), .ZN(n20386) );
  INV_X1 U23322 ( .A(n20382), .ZN(n20384) );
  OAI21_X1 U23323 ( .B1(n20420), .B2(n20396), .A(n20410), .ZN(n20388) );
  AOI22_X1 U23324 ( .A1(n20384), .A2(n20383), .B1(P1_REIP_REG_7__SCAN_IN), 
        .B2(n20388), .ZN(n20385) );
  OAI211_X1 U23325 ( .C1(n20387), .C2(n14969), .A(n20386), .B(n20385), .ZN(
        P1_U2833) );
  AOI22_X1 U23326 ( .A1(n20404), .A2(n20389), .B1(P1_REIP_REG_6__SCAN_IN), 
        .B2(n20388), .ZN(n20400) );
  NAND2_X1 U23327 ( .A1(n20427), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n20390) );
  OAI211_X1 U23328 ( .C1(n20424), .C2(n20391), .A(n20390), .B(n20421), .ZN(
        n20392) );
  INV_X1 U23329 ( .A(n20392), .ZN(n20399) );
  OR2_X1 U23330 ( .A1(n20394), .A2(n20393), .ZN(n20398) );
  OR3_X1 U23331 ( .A1(n20420), .A2(n20396), .A3(n20395), .ZN(n20397) );
  AND4_X1 U23332 ( .A1(n20400), .A2(n20399), .A3(n20398), .A4(n20397), .ZN(
        n20401) );
  OAI21_X1 U23333 ( .B1(n20402), .B2(n14969), .A(n20401), .ZN(P1_U2834) );
  NOR2_X1 U23334 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n20420), .ZN(n20409) );
  AOI22_X1 U23335 ( .A1(n20405), .A2(P1_EBX_REG_5__SCAN_IN), .B1(n20404), .B2(
        n20403), .ZN(n20406) );
  OAI211_X1 U23336 ( .C1(n20407), .C2(n12612), .A(n20406), .B(n20421), .ZN(
        n20408) );
  AOI21_X1 U23337 ( .B1(n20409), .B2(n20419), .A(n20408), .ZN(n20414) );
  OAI21_X1 U23338 ( .B1(n20420), .B2(n20419), .A(n20410), .ZN(n20436) );
  AOI22_X1 U23339 ( .A1(n20412), .A2(n20411), .B1(P1_REIP_REG_5__SCAN_IN), 
        .B2(n20436), .ZN(n20413) );
  OAI211_X1 U23340 ( .C1(n20415), .C2(n9611), .A(n20414), .B(n20413), .ZN(
        P1_U2835) );
  AND2_X1 U23341 ( .A1(n20417), .A2(n20416), .ZN(n20418) );
  OR2_X1 U23342 ( .A1(n20418), .A2(n14441), .ZN(n20525) );
  OR2_X1 U23343 ( .A1(n20420), .A2(n20419), .ZN(n20423) );
  OAI21_X1 U23344 ( .B1(n20423), .B2(n20422), .A(n20421), .ZN(n20426) );
  NOR2_X1 U23345 ( .A1(n20424), .A2(n20446), .ZN(n20425) );
  AOI211_X1 U23346 ( .C1(n20427), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20426), .B(n20425), .ZN(n20431) );
  NAND2_X1 U23347 ( .A1(n20429), .A2(n20428), .ZN(n20430) );
  OAI211_X1 U23348 ( .C1(n20525), .C2(n20432), .A(n20431), .B(n20430), .ZN(
        n20435) );
  NOR2_X1 U23349 ( .A1(n20516), .A2(n20433), .ZN(n20434) );
  OAI21_X1 U23350 ( .B1(n20522), .B2(n9611), .A(n20437), .ZN(P1_U2836) );
  AOI22_X1 U23351 ( .A1(n20441), .A2(n20440), .B1(n20439), .B2(n20438), .ZN(
        n20442) );
  OAI21_X1 U23352 ( .B1(n20447), .B2(n20443), .A(n20442), .ZN(P1_U2864) );
  OAI22_X1 U23353 ( .A1(n20516), .A2(n15011), .B1(n15013), .B2(n20525), .ZN(
        n20444) );
  INV_X1 U23354 ( .A(n20444), .ZN(n20445) );
  OAI21_X1 U23355 ( .B1(n20447), .B2(n20446), .A(n20445), .ZN(P1_U2868) );
  AOI22_X1 U23356 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n20453), .B1(n20472), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20448) );
  OAI21_X1 U23357 ( .B1(n20450), .B2(n20449), .A(n20448), .ZN(P1_U2921) );
  AOI22_X1 U23358 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20473), .B1(n20472), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20451) );
  OAI21_X1 U23359 ( .B1(n15087), .B2(n20475), .A(n20451), .ZN(P1_U2922) );
  AOI22_X1 U23360 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20473), .B1(n20472), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20452) );
  OAI21_X1 U23361 ( .B1(n15088), .B2(n20475), .A(n20452), .ZN(P1_U2923) );
  AOI222_X1 U23362 ( .A1(n20473), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n20453), 
        .B2(P1_EAX_REG_12__SCAN_IN), .C1(P1_DATAO_REG_12__SCAN_IN), .C2(n20472), .ZN(n20454) );
  INV_X1 U23363 ( .A(n20454), .ZN(P1_U2924) );
  AOI22_X1 U23364 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20473), .B1(n20472), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20455) );
  OAI21_X1 U23365 ( .B1(n15091), .B2(n20475), .A(n20455), .ZN(P1_U2925) );
  AOI22_X1 U23366 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20473), .B1(n20472), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20456) );
  OAI21_X1 U23367 ( .B1(n15093), .B2(n20475), .A(n20456), .ZN(P1_U2926) );
  AOI22_X1 U23368 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20473), .B1(n20472), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20457) );
  OAI21_X1 U23369 ( .B1(n15096), .B2(n20475), .A(n20457), .ZN(P1_U2927) );
  AOI22_X1 U23370 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20473), .B1(n20472), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20458) );
  OAI21_X1 U23371 ( .B1(n14465), .B2(n20475), .A(n20458), .ZN(P1_U2928) );
  AOI22_X1 U23372 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20473), .B1(n20472), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20459) );
  OAI21_X1 U23373 ( .B1(n15099), .B2(n20475), .A(n20459), .ZN(P1_U2929) );
  AOI22_X1 U23374 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20473), .B1(n20472), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20460) );
  OAI21_X1 U23375 ( .B1(n20461), .B2(n20475), .A(n20460), .ZN(P1_U2930) );
  AOI22_X1 U23376 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20473), .B1(n20472), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20462) );
  OAI21_X1 U23377 ( .B1(n20463), .B2(n20475), .A(n20462), .ZN(P1_U2931) );
  AOI22_X1 U23378 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20473), .B1(n20472), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20464) );
  OAI21_X1 U23379 ( .B1(n20465), .B2(n20475), .A(n20464), .ZN(P1_U2932) );
  AOI22_X1 U23380 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20473), .B1(n20472), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20466) );
  OAI21_X1 U23381 ( .B1(n20467), .B2(n20475), .A(n20466), .ZN(P1_U2933) );
  AOI22_X1 U23382 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20473), .B1(n20472), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20468) );
  OAI21_X1 U23383 ( .B1(n20469), .B2(n20475), .A(n20468), .ZN(P1_U2934) );
  AOI22_X1 U23384 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20473), .B1(n20472), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20470) );
  OAI21_X1 U23385 ( .B1(n20471), .B2(n20475), .A(n20470), .ZN(P1_U2935) );
  AOI22_X1 U23386 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20473), .B1(n20472), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20474) );
  OAI21_X1 U23387 ( .B1(n21320), .B2(n20475), .A(n20474), .ZN(P1_U2936) );
  AOI22_X1 U23388 ( .A1(n20505), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20508), .ZN(n20478) );
  INV_X1 U23389 ( .A(n20476), .ZN(n20477) );
  NAND2_X1 U23390 ( .A1(n20493), .A2(n20477), .ZN(n20495) );
  NAND2_X1 U23391 ( .A1(n20478), .A2(n20495), .ZN(P1_U2945) );
  AOI22_X1 U23392 ( .A1(n20505), .A2(P1_EAX_REG_25__SCAN_IN), .B1(n20508), 
        .B2(P1_UWORD_REG_9__SCAN_IN), .ZN(n20481) );
  INV_X1 U23393 ( .A(n20479), .ZN(n20480) );
  NAND2_X1 U23394 ( .A1(n20493), .A2(n20480), .ZN(n20497) );
  NAND2_X1 U23395 ( .A1(n20481), .A2(n20497), .ZN(P1_U2946) );
  AOI22_X1 U23396 ( .A1(n20505), .A2(P1_EAX_REG_27__SCAN_IN), .B1(n20508), 
        .B2(P1_UWORD_REG_11__SCAN_IN), .ZN(n20484) );
  INV_X1 U23397 ( .A(n20482), .ZN(n20483) );
  NAND2_X1 U23398 ( .A1(n20493), .A2(n20483), .ZN(n20501) );
  NAND2_X1 U23399 ( .A1(n20484), .A2(n20501), .ZN(P1_U2948) );
  AOI22_X1 U23400 ( .A1(n20505), .A2(P1_EAX_REG_28__SCAN_IN), .B1(n20508), 
        .B2(P1_UWORD_REG_12__SCAN_IN), .ZN(n20487) );
  INV_X1 U23401 ( .A(n20485), .ZN(n20486) );
  NAND2_X1 U23402 ( .A1(n20493), .A2(n20486), .ZN(n20503) );
  NAND2_X1 U23403 ( .A1(n20487), .A2(n20503), .ZN(P1_U2949) );
  AOI22_X1 U23404 ( .A1(n20505), .A2(P1_EAX_REG_29__SCAN_IN), .B1(n20508), 
        .B2(P1_UWORD_REG_13__SCAN_IN), .ZN(n20490) );
  INV_X1 U23405 ( .A(n20488), .ZN(n20489) );
  NAND2_X1 U23406 ( .A1(n20493), .A2(n20489), .ZN(n20506) );
  NAND2_X1 U23407 ( .A1(n20490), .A2(n20506), .ZN(P1_U2950) );
  AOI22_X1 U23408 ( .A1(n20505), .A2(P1_EAX_REG_30__SCAN_IN), .B1(n20508), 
        .B2(P1_UWORD_REG_14__SCAN_IN), .ZN(n20494) );
  INV_X1 U23409 ( .A(n20491), .ZN(n20492) );
  NAND2_X1 U23410 ( .A1(n20493), .A2(n20492), .ZN(n20509) );
  NAND2_X1 U23411 ( .A1(n20494), .A2(n20509), .ZN(P1_U2951) );
  AOI22_X1 U23412 ( .A1(n20505), .A2(P1_EAX_REG_8__SCAN_IN), .B1(n20508), .B2(
        P1_LWORD_REG_8__SCAN_IN), .ZN(n20496) );
  NAND2_X1 U23413 ( .A1(n20496), .A2(n20495), .ZN(P1_U2960) );
  AOI22_X1 U23414 ( .A1(n20505), .A2(P1_EAX_REG_9__SCAN_IN), .B1(n20508), .B2(
        P1_LWORD_REG_9__SCAN_IN), .ZN(n20498) );
  NAND2_X1 U23415 ( .A1(n20498), .A2(n20497), .ZN(P1_U2961) );
  AOI22_X1 U23416 ( .A1(n20505), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n20508), 
        .B2(P1_LWORD_REG_10__SCAN_IN), .ZN(n20500) );
  NAND2_X1 U23417 ( .A1(n20500), .A2(n20499), .ZN(P1_U2962) );
  AOI22_X1 U23418 ( .A1(n20505), .A2(P1_EAX_REG_11__SCAN_IN), .B1(n20508), 
        .B2(P1_LWORD_REG_11__SCAN_IN), .ZN(n20502) );
  NAND2_X1 U23419 ( .A1(n20502), .A2(n20501), .ZN(P1_U2963) );
  AOI22_X1 U23420 ( .A1(n20505), .A2(P1_EAX_REG_12__SCAN_IN), .B1(n20508), 
        .B2(P1_LWORD_REG_12__SCAN_IN), .ZN(n20504) );
  NAND2_X1 U23421 ( .A1(n20504), .A2(n20503), .ZN(P1_U2964) );
  AOI22_X1 U23422 ( .A1(n20505), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n20508), 
        .B2(P1_LWORD_REG_13__SCAN_IN), .ZN(n20507) );
  NAND2_X1 U23423 ( .A1(n20507), .A2(n20506), .ZN(P1_U2965) );
  AOI22_X1 U23424 ( .A1(n20505), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n20508), 
        .B2(P1_LWORD_REG_14__SCAN_IN), .ZN(n20510) );
  NAND2_X1 U23425 ( .A1(n20510), .A2(n20509), .ZN(P1_U2966) );
  AOI22_X1 U23426 ( .A1(n20511), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20577), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20521) );
  AOI21_X1 U23427 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n14429), .A(
        n20512), .ZN(n20515) );
  XNOR2_X1 U23428 ( .A(n20513), .B(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n20514) );
  XNOR2_X1 U23429 ( .A(n20515), .B(n20514), .ZN(n20529) );
  INV_X1 U23430 ( .A(n20516), .ZN(n20517) );
  AOI22_X1 U23431 ( .A1(n20529), .A2(n20519), .B1(n20518), .B2(n20517), .ZN(
        n20520) );
  OAI211_X1 U23432 ( .C1(n9869), .C2(n20522), .A(n20521), .B(n20520), .ZN(
        P1_U2995) );
  INV_X1 U23433 ( .A(n20523), .ZN(n20524) );
  OAI21_X1 U23434 ( .B1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n20524), .ZN(n20532) );
  INV_X1 U23435 ( .A(n20525), .ZN(n20527) );
  AOI22_X1 U23436 ( .A1(n20560), .A2(n20527), .B1(n20526), .B2(
        P1_REIP_REG_4__SCAN_IN), .ZN(n20531) );
  INV_X1 U23437 ( .A(n20528), .ZN(n20535) );
  AOI22_X1 U23438 ( .A1(n20529), .A2(n20563), .B1(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n20535), .ZN(n20530) );
  OAI211_X1 U23439 ( .C1(n20539), .C2(n20532), .A(n20531), .B(n20530), .ZN(
        P1_U3027) );
  AOI21_X1 U23440 ( .B1(n20560), .B2(n20534), .A(n20533), .ZN(n20538) );
  AOI22_X1 U23441 ( .A1(n20536), .A2(n20563), .B1(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n20535), .ZN(n20537) );
  OAI211_X1 U23442 ( .C1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n20539), .A(
        n20538), .B(n20537), .ZN(P1_U3028) );
  AOI21_X1 U23443 ( .B1(n20560), .B2(n20541), .A(n20540), .ZN(n20553) );
  INV_X1 U23444 ( .A(n20542), .ZN(n20547) );
  NAND3_X1 U23445 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n20570), .ZN(n20543) );
  OAI211_X1 U23446 ( .C1(n20545), .C2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n20544), .B(n20543), .ZN(n20546) );
  AOI22_X1 U23447 ( .A1(n20547), .A2(n20563), .B1(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20546), .ZN(n20552) );
  NAND3_X1 U23448 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20549), .A3(
        n20548), .ZN(n20550) );
  NAND4_X1 U23449 ( .A1(n20553), .A2(n20552), .A3(n20551), .A4(n20550), .ZN(
        P1_U3029) );
  AOI21_X1 U23450 ( .B1(n20570), .B2(n20555), .A(n20554), .ZN(n20580) );
  INV_X1 U23451 ( .A(n20556), .ZN(n20559) );
  INV_X1 U23452 ( .A(n20557), .ZN(n20558) );
  AOI21_X1 U23453 ( .B1(n20560), .B2(n20559), .A(n20558), .ZN(n20568) );
  OR3_X1 U23454 ( .A1(n20562), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n20561), .ZN(n20566) );
  NAND3_X1 U23455 ( .A1(n20564), .A2(n15315), .A3(n20563), .ZN(n20565) );
  AND2_X1 U23456 ( .A1(n20566), .A2(n20565), .ZN(n20567) );
  OAI211_X1 U23457 ( .C1(n20580), .C2(n20569), .A(n20568), .B(n20567), .ZN(
        P1_U3030) );
  NOR3_X1 U23458 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n20571), .A3(
        n20570), .ZN(n20581) );
  OAI22_X1 U23459 ( .A1(n20575), .A2(n20574), .B1(n20573), .B2(n20572), .ZN(
        n20576) );
  AOI21_X1 U23460 ( .B1(n20577), .B2(P1_REIP_REG_0__SCAN_IN), .A(n20576), .ZN(
        n20578) );
  OAI221_X1 U23461 ( .B1(n20581), .B2(n20580), .C1(n20581), .C2(n20579), .A(
        n20578), .ZN(P1_U3031) );
  AND2_X1 U23462 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n21382), .ZN(
        P1_U3032) );
  AOI22_X1 U23463 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20629), .B1(DATAI_16_), 
        .B2(n20628), .ZN(n21032) );
  NOR2_X2 U23464 ( .A1(n20627), .A2(n12427), .ZN(n21072) );
  NAND2_X1 U23465 ( .A1(n20589), .A2(n20840), .ZN(n20693) );
  AOI22_X1 U23466 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20629), .B1(DATAI_24_), 
        .B2(n20628), .ZN(n21085) );
  INV_X1 U23467 ( .A(n21085), .ZN(n21029) );
  AOI22_X1 U23468 ( .A1(n21072), .A2(n10413), .B1(n21127), .B2(n21029), .ZN(
        n20602) );
  OR2_X1 U23469 ( .A1(n20597), .A2(n21070), .ZN(n21019) );
  INV_X1 U23470 ( .A(n21019), .ZN(n20590) );
  NAND2_X1 U23471 ( .A1(n20660), .A2(n20591), .ZN(n20592) );
  AOI21_X1 U23472 ( .B1(n20592), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n21075), 
        .ZN(n20596) );
  OR2_X1 U23473 ( .A1(n20839), .A2(n20593), .ZN(n20665) );
  OR2_X1 U23474 ( .A1(n20665), .A2(n10366), .ZN(n20599) );
  OR2_X1 U23475 ( .A1(n20841), .A2(n20897), .ZN(n20726) );
  AOI22_X1 U23476 ( .A1(n20596), .A2(n20599), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20726), .ZN(n20594) );
  NOR2_X2 U23477 ( .A1(n20729), .A2(n20595), .ZN(n21073) );
  INV_X1 U23478 ( .A(n20596), .ZN(n20600) );
  INV_X1 U23479 ( .A(n20597), .ZN(n20598) );
  NOR2_X1 U23480 ( .A1(n20598), .A2(n21070), .ZN(n20730) );
  INV_X1 U23481 ( .A(n20730), .ZN(n20902) );
  AOI22_X1 U23482 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20632), .B1(
        n21073), .B2(n20631), .ZN(n20601) );
  OAI211_X1 U23483 ( .C1(n21032), .C2(n20660), .A(n20602), .B(n20601), .ZN(
        P1_U3033) );
  AOI22_X1 U23484 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n20629), .B1(DATAI_17_), 
        .B2(n20628), .ZN(n21036) );
  NOR2_X2 U23485 ( .A1(n20627), .A2(n20603), .ZN(n21086) );
  AOI22_X1 U23486 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20629), .B1(DATAI_25_), 
        .B2(n20628), .ZN(n21091) );
  INV_X1 U23487 ( .A(n21091), .ZN(n21033) );
  AOI22_X1 U23488 ( .A1(n21086), .A2(n10413), .B1(n21127), .B2(n21033), .ZN(
        n20606) );
  NOR2_X2 U23489 ( .A1(n20729), .A2(n20604), .ZN(n21087) );
  AOI22_X1 U23490 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20632), .B1(
        n21087), .B2(n20631), .ZN(n20605) );
  OAI211_X1 U23491 ( .C1(n21036), .C2(n20660), .A(n20606), .B(n20605), .ZN(
        P1_U3034) );
  AOI22_X1 U23492 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20629), .B1(DATAI_18_), 
        .B2(n20628), .ZN(n21040) );
  NOR2_X2 U23493 ( .A1(n20627), .A2(n20607), .ZN(n21092) );
  AOI22_X1 U23494 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20629), .B1(DATAI_26_), 
        .B2(n20628), .ZN(n21097) );
  INV_X1 U23495 ( .A(n21097), .ZN(n21037) );
  AOI22_X1 U23496 ( .A1(n21092), .A2(n10413), .B1(n21127), .B2(n21037), .ZN(
        n20610) );
  NOR2_X2 U23497 ( .A1(n20729), .A2(n20608), .ZN(n21093) );
  AOI22_X1 U23498 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20632), .B1(
        n21093), .B2(n20631), .ZN(n20609) );
  OAI211_X1 U23499 ( .C1(n21040), .C2(n20660), .A(n20610), .B(n20609), .ZN(
        P1_U3035) );
  AOI22_X1 U23500 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20629), .B1(DATAI_19_), 
        .B2(n20628), .ZN(n21044) );
  NOR2_X2 U23501 ( .A1(n20627), .A2(n20611), .ZN(n21098) );
  AOI22_X1 U23502 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20629), .B1(DATAI_27_), 
        .B2(n20628), .ZN(n21103) );
  INV_X1 U23503 ( .A(n21103), .ZN(n21041) );
  AOI22_X1 U23504 ( .A1(n21098), .A2(n10413), .B1(n21127), .B2(n21041), .ZN(
        n20614) );
  NOR2_X2 U23505 ( .A1(n20729), .A2(n20612), .ZN(n21099) );
  AOI22_X1 U23506 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20632), .B1(
        n21099), .B2(n20631), .ZN(n20613) );
  OAI211_X1 U23507 ( .C1(n21044), .C2(n20660), .A(n20614), .B(n20613), .ZN(
        P1_U3036) );
  AOI22_X1 U23508 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20629), .B1(DATAI_20_), 
        .B2(n20628), .ZN(n21048) );
  NOR2_X2 U23509 ( .A1(n20627), .A2(n20615), .ZN(n21104) );
  AOI22_X1 U23510 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20629), .B1(DATAI_28_), 
        .B2(n20628), .ZN(n21109) );
  INV_X1 U23511 ( .A(n21109), .ZN(n21045) );
  AOI22_X1 U23512 ( .A1(n21104), .A2(n10413), .B1(n21127), .B2(n21045), .ZN(
        n20618) );
  NOR2_X2 U23513 ( .A1(n20729), .A2(n20616), .ZN(n21105) );
  AOI22_X1 U23514 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20632), .B1(
        n21105), .B2(n20631), .ZN(n20617) );
  OAI211_X1 U23515 ( .C1(n21048), .C2(n20660), .A(n20618), .B(n20617), .ZN(
        P1_U3037) );
  AOI22_X1 U23516 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n20629), .B1(DATAI_21_), 
        .B2(n20628), .ZN(n21052) );
  AOI22_X1 U23517 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20629), .B1(DATAI_29_), 
        .B2(n20628), .ZN(n21115) );
  AOI22_X1 U23518 ( .A1(n9565), .A2(n10413), .B1(n21127), .B2(n21049), .ZN(
        n20621) );
  NOR2_X2 U23519 ( .A1(n20729), .A2(n20619), .ZN(n21111) );
  AOI22_X1 U23520 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20632), .B1(
        n21111), .B2(n20631), .ZN(n20620) );
  OAI211_X1 U23521 ( .C1(n21052), .C2(n20660), .A(n20621), .B(n20620), .ZN(
        P1_U3038) );
  AOI22_X1 U23522 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20629), .B1(DATAI_22_), 
        .B2(n20628), .ZN(n21056) );
  NOR2_X2 U23523 ( .A1(n20627), .A2(n20622), .ZN(n21116) );
  INV_X1 U23524 ( .A(n21121), .ZN(n21053) );
  AOI22_X1 U23525 ( .A1(n21116), .A2(n10413), .B1(n21127), .B2(n21053), .ZN(
        n20625) );
  NOR2_X2 U23526 ( .A1(n20729), .A2(n20623), .ZN(n21117) );
  AOI22_X1 U23527 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20632), .B1(
        n21117), .B2(n20631), .ZN(n20624) );
  OAI211_X1 U23528 ( .C1(n21056), .C2(n20660), .A(n20625), .B(n20624), .ZN(
        P1_U3039) );
  AOI22_X1 U23529 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20629), .B1(DATAI_23_), 
        .B2(n20628), .ZN(n21064) );
  INV_X1 U23530 ( .A(n21132), .ZN(n21059) );
  AOI22_X1 U23531 ( .A1(n9567), .A2(n10413), .B1(n21127), .B2(n21059), .ZN(
        n20634) );
  NOR2_X2 U23532 ( .A1(n20729), .A2(n20630), .ZN(n21125) );
  AOI22_X1 U23533 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20632), .B1(
        n21125), .B2(n20631), .ZN(n20633) );
  OAI211_X1 U23534 ( .C1(n21064), .C2(n20660), .A(n20634), .B(n20633), .ZN(
        P1_U3040) );
  OR2_X1 U23535 ( .A1(n20635), .A2(n21075), .ZN(n20868) );
  NOR2_X1 U23536 ( .A1(n20693), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20638) );
  INV_X1 U23537 ( .A(n20638), .ZN(n20637) );
  NOR2_X1 U23538 ( .A1(n20988), .A2(n20637), .ZN(n20655) );
  INV_X1 U23539 ( .A(n20655), .ZN(n20636) );
  OAI222_X1 U23540 ( .A1(n20868), .A2(n20665), .B1(n21070), .B2(n20637), .C1(
        n21075), .C2(n20636), .ZN(n20656) );
  AOI22_X1 U23541 ( .A1(n21073), .A2(n20656), .B1(n21072), .B2(n20655), .ZN(
        n20641) );
  NOR2_X1 U23542 ( .A1(n20697), .A2(n20869), .ZN(n20639) );
  INV_X1 U23543 ( .A(n21032), .ZN(n21082) );
  AOI22_X1 U23544 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20657), .B1(
        n20682), .B2(n21082), .ZN(n20640) );
  OAI211_X1 U23545 ( .C1(n21085), .C2(n20660), .A(n20641), .B(n20640), .ZN(
        P1_U3041) );
  AOI22_X1 U23546 ( .A1(n21087), .A2(n20656), .B1(n21086), .B2(n20655), .ZN(
        n20643) );
  INV_X1 U23547 ( .A(n20660), .ZN(n20650) );
  AOI22_X1 U23548 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20657), .B1(
        n20650), .B2(n21033), .ZN(n20642) );
  OAI211_X1 U23549 ( .C1(n21036), .C2(n20692), .A(n20643), .B(n20642), .ZN(
        P1_U3042) );
  AOI22_X1 U23550 ( .A1(n21093), .A2(n20656), .B1(n21092), .B2(n20655), .ZN(
        n20645) );
  INV_X1 U23551 ( .A(n21040), .ZN(n21094) );
  AOI22_X1 U23552 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20657), .B1(
        n20682), .B2(n21094), .ZN(n20644) );
  OAI211_X1 U23553 ( .C1(n21097), .C2(n20660), .A(n20645), .B(n20644), .ZN(
        P1_U3043) );
  AOI22_X1 U23554 ( .A1(n21099), .A2(n20656), .B1(n21098), .B2(n20655), .ZN(
        n20647) );
  AOI22_X1 U23555 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20657), .B1(
        n20650), .B2(n21041), .ZN(n20646) );
  OAI211_X1 U23556 ( .C1(n21044), .C2(n20692), .A(n20647), .B(n20646), .ZN(
        P1_U3044) );
  AOI22_X1 U23557 ( .A1(n21105), .A2(n20656), .B1(n21104), .B2(n20655), .ZN(
        n20649) );
  INV_X1 U23558 ( .A(n21048), .ZN(n21106) );
  AOI22_X1 U23559 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20657), .B1(
        n20682), .B2(n21106), .ZN(n20648) );
  OAI211_X1 U23560 ( .C1(n21109), .C2(n20660), .A(n20649), .B(n20648), .ZN(
        P1_U3045) );
  AOI22_X1 U23561 ( .A1(n21111), .A2(n20656), .B1(n9565), .B2(n20655), .ZN(
        n20652) );
  AOI22_X1 U23562 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20657), .B1(
        n20650), .B2(n21049), .ZN(n20651) );
  OAI211_X1 U23563 ( .C1(n21052), .C2(n20692), .A(n20652), .B(n20651), .ZN(
        P1_U3046) );
  AOI22_X1 U23564 ( .A1(n21117), .A2(n20656), .B1(n21116), .B2(n20655), .ZN(
        n20654) );
  INV_X1 U23565 ( .A(n21056), .ZN(n21118) );
  AOI22_X1 U23566 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20657), .B1(
        n20682), .B2(n21118), .ZN(n20653) );
  OAI211_X1 U23567 ( .C1(n21121), .C2(n20660), .A(n20654), .B(n20653), .ZN(
        P1_U3047) );
  AOI22_X1 U23568 ( .A1(n21125), .A2(n20656), .B1(n9567), .B2(n20655), .ZN(
        n20659) );
  INV_X1 U23569 ( .A(n21064), .ZN(n21126) );
  AOI22_X1 U23570 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20657), .B1(
        n20682), .B2(n21126), .ZN(n20658) );
  OAI211_X1 U23571 ( .C1(n21132), .C2(n20660), .A(n20659), .B(n20658), .ZN(
        P1_U3048) );
  INV_X1 U23572 ( .A(n20693), .ZN(n20663) );
  NAND2_X1 U23573 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20663), .ZN(
        n20700) );
  NOR2_X1 U23574 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20700), .ZN(
        n20687) );
  AOI22_X1 U23575 ( .A1(n21072), .A2(n20687), .B1(n20682), .B2(n21029), .ZN(
        n20673) );
  NAND2_X1 U23576 ( .A1(n20723), .A2(n20692), .ZN(n20664) );
  AOI21_X1 U23577 ( .B1(n20664), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n21075), 
        .ZN(n20668) );
  INV_X1 U23578 ( .A(n20665), .ZN(n20695) );
  NAND2_X1 U23579 ( .A1(n20695), .A2(n10366), .ZN(n20670) );
  INV_X1 U23580 ( .A(n20897), .ZN(n20842) );
  NOR2_X1 U23581 ( .A1(n20842), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20669) );
  NOR2_X1 U23582 ( .A1(n20669), .A2(n21070), .ZN(n20780) );
  INV_X1 U23583 ( .A(n20898), .ZN(n20666) );
  AOI211_X1 U23584 ( .C1(n20668), .C2(n20670), .A(n20780), .B(n20666), .ZN(
        n20667) );
  INV_X1 U23585 ( .A(n20668), .ZN(n20671) );
  INV_X1 U23586 ( .A(n20669), .ZN(n20783) );
  AOI22_X1 U23587 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20689), .B1(
        n21073), .B2(n20688), .ZN(n20672) );
  OAI211_X1 U23588 ( .C1(n21032), .C2(n20723), .A(n20673), .B(n20672), .ZN(
        P1_U3049) );
  AOI22_X1 U23589 ( .A1(n21086), .A2(n20687), .B1(n20682), .B2(n21033), .ZN(
        n20675) );
  AOI22_X1 U23590 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20689), .B1(
        n21087), .B2(n20688), .ZN(n20674) );
  OAI211_X1 U23591 ( .C1(n21036), .C2(n20723), .A(n20675), .B(n20674), .ZN(
        P1_U3050) );
  AOI22_X1 U23592 ( .A1(n21092), .A2(n20687), .B1(n20713), .B2(n21094), .ZN(
        n20677) );
  AOI22_X1 U23593 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20689), .B1(
        n21093), .B2(n20688), .ZN(n20676) );
  OAI211_X1 U23594 ( .C1(n21097), .C2(n20692), .A(n20677), .B(n20676), .ZN(
        P1_U3051) );
  INV_X1 U23595 ( .A(n21044), .ZN(n21100) );
  AOI22_X1 U23596 ( .A1(n21098), .A2(n20687), .B1(n20713), .B2(n21100), .ZN(
        n20679) );
  AOI22_X1 U23597 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20689), .B1(
        n21099), .B2(n20688), .ZN(n20678) );
  OAI211_X1 U23598 ( .C1(n21103), .C2(n20692), .A(n20679), .B(n20678), .ZN(
        P1_U3052) );
  AOI22_X1 U23599 ( .A1(n21104), .A2(n20687), .B1(n20713), .B2(n21106), .ZN(
        n20681) );
  AOI22_X1 U23600 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20689), .B1(
        n21105), .B2(n20688), .ZN(n20680) );
  OAI211_X1 U23601 ( .C1(n21109), .C2(n20692), .A(n20681), .B(n20680), .ZN(
        P1_U3053) );
  AOI22_X1 U23602 ( .A1(n9565), .A2(n20687), .B1(n20682), .B2(n21049), .ZN(
        n20684) );
  AOI22_X1 U23603 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20689), .B1(
        n21111), .B2(n20688), .ZN(n20683) );
  OAI211_X1 U23604 ( .C1(n21052), .C2(n20723), .A(n20684), .B(n20683), .ZN(
        P1_U3054) );
  AOI22_X1 U23605 ( .A1(n21116), .A2(n20687), .B1(n20713), .B2(n21118), .ZN(
        n20686) );
  AOI22_X1 U23606 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20689), .B1(
        n21117), .B2(n20688), .ZN(n20685) );
  OAI211_X1 U23607 ( .C1(n21121), .C2(n20692), .A(n20686), .B(n20685), .ZN(
        P1_U3055) );
  AOI22_X1 U23608 ( .A1(n9567), .A2(n20687), .B1(n20713), .B2(n21126), .ZN(
        n20691) );
  AOI22_X1 U23609 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20689), .B1(
        n21125), .B2(n20688), .ZN(n20690) );
  OAI211_X1 U23610 ( .C1(n21132), .C2(n20692), .A(n20691), .B(n20690), .ZN(
        P1_U3056) );
  NOR2_X1 U23611 ( .A1(n21065), .A2(n20693), .ZN(n20718) );
  AOI22_X1 U23612 ( .A1(n21072), .A2(n20718), .B1(n20742), .B2(n21082), .ZN(
        n20704) );
  AND2_X1 U23613 ( .A1(n20694), .A2(n21386), .ZN(n21066) );
  AOI21_X1 U23614 ( .B1(n20695), .B2(n21066), .A(n20718), .ZN(n20702) );
  INV_X1 U23615 ( .A(n21074), .ZN(n20696) );
  AOI21_X1 U23616 ( .B1(n20697), .B2(n21383), .A(n20696), .ZN(n20701) );
  INV_X1 U23617 ( .A(n20701), .ZN(n20698) );
  AOI22_X1 U23618 ( .A1(n20702), .A2(n20698), .B1(n21075), .B2(n20700), .ZN(
        n20699) );
  NAND2_X1 U23619 ( .A1(n21080), .A2(n20699), .ZN(n20720) );
  AOI22_X1 U23620 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20720), .B1(
        n21073), .B2(n20719), .ZN(n20703) );
  OAI211_X1 U23621 ( .C1(n21085), .C2(n20723), .A(n20704), .B(n20703), .ZN(
        P1_U3057) );
  INV_X1 U23622 ( .A(n21036), .ZN(n21088) );
  AOI22_X1 U23623 ( .A1(n21086), .A2(n20718), .B1(n20742), .B2(n21088), .ZN(
        n20706) );
  AOI22_X1 U23624 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20720), .B1(
        n21087), .B2(n20719), .ZN(n20705) );
  OAI211_X1 U23625 ( .C1(n21091), .C2(n20723), .A(n20706), .B(n20705), .ZN(
        P1_U3058) );
  AOI22_X1 U23626 ( .A1(n21092), .A2(n20718), .B1(n20713), .B2(n21037), .ZN(
        n20708) );
  AOI22_X1 U23627 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20720), .B1(
        n21093), .B2(n20719), .ZN(n20707) );
  OAI211_X1 U23628 ( .C1(n21040), .C2(n20751), .A(n20708), .B(n20707), .ZN(
        P1_U3059) );
  AOI22_X1 U23629 ( .A1(n21098), .A2(n20718), .B1(n20742), .B2(n21100), .ZN(
        n20710) );
  AOI22_X1 U23630 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20720), .B1(
        n21099), .B2(n20719), .ZN(n20709) );
  OAI211_X1 U23631 ( .C1(n21103), .C2(n20723), .A(n20710), .B(n20709), .ZN(
        P1_U3060) );
  AOI22_X1 U23632 ( .A1(n21104), .A2(n20718), .B1(n20713), .B2(n21045), .ZN(
        n20712) );
  AOI22_X1 U23633 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20720), .B1(
        n21105), .B2(n20719), .ZN(n20711) );
  OAI211_X1 U23634 ( .C1(n21048), .C2(n20751), .A(n20712), .B(n20711), .ZN(
        P1_U3061) );
  AOI22_X1 U23635 ( .A1(n9565), .A2(n20718), .B1(n20713), .B2(n21049), .ZN(
        n20715) );
  AOI22_X1 U23636 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20720), .B1(
        n21111), .B2(n20719), .ZN(n20714) );
  OAI211_X1 U23637 ( .C1(n21052), .C2(n20751), .A(n20715), .B(n20714), .ZN(
        P1_U3062) );
  AOI22_X1 U23638 ( .A1(n21116), .A2(n20718), .B1(n20742), .B2(n21118), .ZN(
        n20717) );
  AOI22_X1 U23639 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20720), .B1(
        n21117), .B2(n20719), .ZN(n20716) );
  OAI211_X1 U23640 ( .C1(n21121), .C2(n20723), .A(n20717), .B(n20716), .ZN(
        P1_U3063) );
  AOI22_X1 U23641 ( .A1(n9567), .A2(n20718), .B1(n20742), .B2(n21126), .ZN(
        n20722) );
  AOI22_X1 U23642 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20720), .B1(
        n21125), .B2(n20719), .ZN(n20721) );
  OAI211_X1 U23643 ( .C1(n21132), .C2(n20723), .A(n20722), .B(n20721), .ZN(
        P1_U3064) );
  NOR2_X1 U23644 ( .A1(n13947), .A2(n20724), .ZN(n20809) );
  NAND3_X1 U23645 ( .A1(n20809), .A2(n21383), .A3(n14960), .ZN(n20725) );
  OAI21_X1 U23646 ( .B1(n20726), .B2(n21019), .A(n20725), .ZN(n20747) );
  AOI22_X1 U23647 ( .A1(n21073), .A2(n20747), .B1(n21072), .B2(n10419), .ZN(
        n20733) );
  AOI21_X1 U23648 ( .B1(n20751), .B2(n20777), .A(n21022), .ZN(n20727) );
  AOI21_X1 U23649 ( .B1(n20809), .B2(n14960), .A(n20727), .ZN(n20728) );
  NOR2_X1 U23650 ( .A1(n20728), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20731) );
  AOI22_X1 U23651 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20748), .B1(
        n20742), .B2(n21029), .ZN(n20732) );
  OAI211_X1 U23652 ( .C1(n21032), .C2(n20777), .A(n20733), .B(n20732), .ZN(
        P1_U3065) );
  AOI22_X1 U23653 ( .A1(n21087), .A2(n20747), .B1(n21086), .B2(n10419), .ZN(
        n20735) );
  AOI22_X1 U23654 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20748), .B1(
        n20742), .B2(n21033), .ZN(n20734) );
  OAI211_X1 U23655 ( .C1(n21036), .C2(n20777), .A(n20735), .B(n20734), .ZN(
        P1_U3066) );
  AOI22_X1 U23656 ( .A1(n21093), .A2(n20747), .B1(n21092), .B2(n10419), .ZN(
        n20737) );
  AOI22_X1 U23657 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20748), .B1(
        n20767), .B2(n21094), .ZN(n20736) );
  OAI211_X1 U23658 ( .C1(n21097), .C2(n20751), .A(n20737), .B(n20736), .ZN(
        P1_U3067) );
  AOI22_X1 U23659 ( .A1(n21099), .A2(n20747), .B1(n21098), .B2(n10419), .ZN(
        n20739) );
  AOI22_X1 U23660 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20748), .B1(
        n20767), .B2(n21100), .ZN(n20738) );
  OAI211_X1 U23661 ( .C1(n21103), .C2(n20751), .A(n20739), .B(n20738), .ZN(
        P1_U3068) );
  AOI22_X1 U23662 ( .A1(n21105), .A2(n20747), .B1(n21104), .B2(n10419), .ZN(
        n20741) );
  AOI22_X1 U23663 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20748), .B1(
        n20767), .B2(n21106), .ZN(n20740) );
  OAI211_X1 U23664 ( .C1(n21109), .C2(n20751), .A(n20741), .B(n20740), .ZN(
        P1_U3069) );
  AOI22_X1 U23665 ( .A1(n21111), .A2(n20747), .B1(n9565), .B2(n10419), .ZN(
        n20744) );
  AOI22_X1 U23666 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20748), .B1(
        n20742), .B2(n21049), .ZN(n20743) );
  OAI211_X1 U23667 ( .C1(n21052), .C2(n20777), .A(n20744), .B(n20743), .ZN(
        P1_U3070) );
  AOI22_X1 U23668 ( .A1(n21117), .A2(n20747), .B1(n21116), .B2(n10419), .ZN(
        n20746) );
  AOI22_X1 U23669 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20748), .B1(
        n20767), .B2(n21118), .ZN(n20745) );
  OAI211_X1 U23670 ( .C1(n21121), .C2(n20751), .A(n20746), .B(n20745), .ZN(
        P1_U3071) );
  AOI22_X1 U23671 ( .A1(n21125), .A2(n20747), .B1(n9567), .B2(n10419), .ZN(
        n20750) );
  AOI22_X1 U23672 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20748), .B1(
        n20767), .B2(n21126), .ZN(n20749) );
  OAI211_X1 U23673 ( .C1(n21132), .C2(n20751), .A(n20750), .B(n20749), .ZN(
        P1_U3072) );
  INV_X1 U23674 ( .A(n20809), .ZN(n20754) );
  NOR2_X1 U23675 ( .A1(n20778), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20755) );
  INV_X1 U23676 ( .A(n20755), .ZN(n20753) );
  NOR2_X1 U23677 ( .A1(n20988), .A2(n20753), .ZN(n20772) );
  INV_X1 U23678 ( .A(n20772), .ZN(n20752) );
  OAI222_X1 U23679 ( .A1(n20868), .A2(n20754), .B1(n21070), .B2(n20753), .C1(
        n21075), .C2(n20752), .ZN(n20773) );
  AOI22_X1 U23680 ( .A1(n21073), .A2(n20773), .B1(n21072), .B2(n20772), .ZN(
        n20758) );
  NOR2_X1 U23681 ( .A1(n20807), .A2(n20869), .ZN(n20756) );
  AOI22_X1 U23682 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20774), .B1(
        n20801), .B2(n21082), .ZN(n20757) );
  OAI211_X1 U23683 ( .C1(n21085), .C2(n20777), .A(n20758), .B(n20757), .ZN(
        P1_U3073) );
  AOI22_X1 U23684 ( .A1(n21087), .A2(n20773), .B1(n21086), .B2(n20772), .ZN(
        n20760) );
  AOI22_X1 U23685 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20774), .B1(
        n20767), .B2(n21033), .ZN(n20759) );
  OAI211_X1 U23686 ( .C1(n21036), .C2(n20798), .A(n20760), .B(n20759), .ZN(
        P1_U3074) );
  AOI22_X1 U23687 ( .A1(n21093), .A2(n20773), .B1(n21092), .B2(n20772), .ZN(
        n20762) );
  AOI22_X1 U23688 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20774), .B1(
        n20767), .B2(n21037), .ZN(n20761) );
  OAI211_X1 U23689 ( .C1(n21040), .C2(n20798), .A(n20762), .B(n20761), .ZN(
        P1_U3075) );
  AOI22_X1 U23690 ( .A1(n21099), .A2(n20773), .B1(n21098), .B2(n20772), .ZN(
        n20764) );
  AOI22_X1 U23691 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20774), .B1(
        n20801), .B2(n21100), .ZN(n20763) );
  OAI211_X1 U23692 ( .C1(n21103), .C2(n20777), .A(n20764), .B(n20763), .ZN(
        P1_U3076) );
  AOI22_X1 U23693 ( .A1(n21105), .A2(n20773), .B1(n21104), .B2(n20772), .ZN(
        n20766) );
  AOI22_X1 U23694 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20774), .B1(
        n20767), .B2(n21045), .ZN(n20765) );
  OAI211_X1 U23695 ( .C1(n21048), .C2(n20798), .A(n20766), .B(n20765), .ZN(
        P1_U3077) );
  AOI22_X1 U23696 ( .A1(n21111), .A2(n20773), .B1(n9565), .B2(n20772), .ZN(
        n20769) );
  AOI22_X1 U23697 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20774), .B1(
        n20767), .B2(n21049), .ZN(n20768) );
  OAI211_X1 U23698 ( .C1(n21052), .C2(n20798), .A(n20769), .B(n20768), .ZN(
        P1_U3078) );
  AOI22_X1 U23699 ( .A1(n21117), .A2(n20773), .B1(n21116), .B2(n20772), .ZN(
        n20771) );
  AOI22_X1 U23700 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20774), .B1(
        n20801), .B2(n21118), .ZN(n20770) );
  OAI211_X1 U23701 ( .C1(n21121), .C2(n20777), .A(n20771), .B(n20770), .ZN(
        P1_U3079) );
  AOI22_X1 U23702 ( .A1(n21125), .A2(n20773), .B1(n9567), .B2(n20772), .ZN(
        n20776) );
  AOI22_X1 U23703 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20774), .B1(
        n20801), .B2(n21126), .ZN(n20775) );
  OAI211_X1 U23704 ( .C1(n21132), .C2(n20777), .A(n20776), .B(n20775), .ZN(
        P1_U3080) );
  NOR2_X1 U23705 ( .A1(n21069), .A2(n20778), .ZN(n20815) );
  INV_X1 U23706 ( .A(n20815), .ZN(n20810) );
  NOR2_X1 U23707 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20810), .ZN(
        n20802) );
  AOI22_X1 U23708 ( .A1(n21072), .A2(n20802), .B1(n20801), .B2(n21029), .ZN(
        n20787) );
  NAND2_X1 U23709 ( .A1(n20837), .A2(n20798), .ZN(n20779) );
  AOI21_X1 U23710 ( .B1(n20779), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n21075), 
        .ZN(n20782) );
  NAND2_X1 U23711 ( .A1(n20809), .A2(n10366), .ZN(n20784) );
  AOI21_X1 U23712 ( .B1(n20782), .B2(n20784), .A(n20780), .ZN(n20781) );
  INV_X1 U23713 ( .A(n20782), .ZN(n20785) );
  AOI22_X1 U23714 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20804), .B1(
        n21073), .B2(n20803), .ZN(n20786) );
  OAI211_X1 U23715 ( .C1(n21032), .C2(n20837), .A(n20787), .B(n20786), .ZN(
        P1_U3081) );
  AOI22_X1 U23716 ( .A1(n21086), .A2(n20802), .B1(n20828), .B2(n21088), .ZN(
        n20789) );
  AOI22_X1 U23717 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20804), .B1(
        n21087), .B2(n20803), .ZN(n20788) );
  OAI211_X1 U23718 ( .C1(n21091), .C2(n20798), .A(n20789), .B(n20788), .ZN(
        P1_U3082) );
  AOI22_X1 U23719 ( .A1(n21092), .A2(n20802), .B1(n20828), .B2(n21094), .ZN(
        n20791) );
  AOI22_X1 U23720 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20804), .B1(
        n21093), .B2(n20803), .ZN(n20790) );
  OAI211_X1 U23721 ( .C1(n21097), .C2(n20798), .A(n20791), .B(n20790), .ZN(
        P1_U3083) );
  AOI22_X1 U23722 ( .A1(n21098), .A2(n20802), .B1(n20801), .B2(n21041), .ZN(
        n20793) );
  AOI22_X1 U23723 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20804), .B1(
        n21099), .B2(n20803), .ZN(n20792) );
  OAI211_X1 U23724 ( .C1(n21044), .C2(n20837), .A(n20793), .B(n20792), .ZN(
        P1_U3084) );
  AOI22_X1 U23725 ( .A1(n21104), .A2(n20802), .B1(n20828), .B2(n21106), .ZN(
        n20795) );
  AOI22_X1 U23726 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20804), .B1(
        n21105), .B2(n20803), .ZN(n20794) );
  OAI211_X1 U23727 ( .C1(n21109), .C2(n20798), .A(n20795), .B(n20794), .ZN(
        P1_U3085) );
  INV_X1 U23728 ( .A(n21052), .ZN(n21112) );
  AOI22_X1 U23729 ( .A1(n9565), .A2(n20802), .B1(n20828), .B2(n21112), .ZN(
        n20797) );
  AOI22_X1 U23730 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20804), .B1(
        n21111), .B2(n20803), .ZN(n20796) );
  OAI211_X1 U23731 ( .C1(n21115), .C2(n20798), .A(n20797), .B(n20796), .ZN(
        P1_U3086) );
  AOI22_X1 U23732 ( .A1(n21116), .A2(n20802), .B1(n20801), .B2(n21053), .ZN(
        n20800) );
  AOI22_X1 U23733 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20804), .B1(
        n21117), .B2(n20803), .ZN(n20799) );
  OAI211_X1 U23734 ( .C1(n21056), .C2(n20837), .A(n20800), .B(n20799), .ZN(
        P1_U3087) );
  AOI22_X1 U23735 ( .A1(n9567), .A2(n20802), .B1(n20801), .B2(n21059), .ZN(
        n20806) );
  AOI22_X1 U23736 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20804), .B1(
        n21125), .B2(n20803), .ZN(n20805) );
  OAI211_X1 U23737 ( .C1(n21064), .C2(n20837), .A(n20806), .B(n20805), .ZN(
        P1_U3088) );
  INV_X1 U23738 ( .A(n20808), .ZN(n20832) );
  AOI21_X1 U23739 ( .B1(n20809), .B2(n21066), .A(n20832), .ZN(n20812) );
  OAI22_X1 U23740 ( .A1(n20812), .A2(n21075), .B1(n20810), .B2(n21070), .ZN(
        n20833) );
  AOI22_X1 U23741 ( .A1(n21073), .A2(n20833), .B1(n21072), .B2(n20832), .ZN(
        n20817) );
  INV_X1 U23742 ( .A(n20811), .ZN(n20813) );
  NAND2_X1 U23743 ( .A1(n20813), .A2(n20812), .ZN(n20814) );
  AOI22_X1 U23744 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20834), .B1(
        n20828), .B2(n21029), .ZN(n20816) );
  OAI211_X1 U23745 ( .C1(n21032), .C2(n20831), .A(n20817), .B(n20816), .ZN(
        P1_U3089) );
  AOI22_X1 U23746 ( .A1(n21087), .A2(n20833), .B1(n21086), .B2(n20832), .ZN(
        n20819) );
  AOI22_X1 U23747 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20834), .B1(
        n20828), .B2(n21033), .ZN(n20818) );
  OAI211_X1 U23748 ( .C1(n21036), .C2(n20831), .A(n20819), .B(n20818), .ZN(
        P1_U3090) );
  AOI22_X1 U23749 ( .A1(n21093), .A2(n20833), .B1(n21092), .B2(n20832), .ZN(
        n20821) );
  AOI22_X1 U23750 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20834), .B1(
        n20862), .B2(n21094), .ZN(n20820) );
  OAI211_X1 U23751 ( .C1(n21097), .C2(n20837), .A(n20821), .B(n20820), .ZN(
        P1_U3091) );
  AOI22_X1 U23752 ( .A1(n21099), .A2(n20833), .B1(n21098), .B2(n20832), .ZN(
        n20823) );
  AOI22_X1 U23753 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20834), .B1(
        n20828), .B2(n21041), .ZN(n20822) );
  OAI211_X1 U23754 ( .C1(n21044), .C2(n20831), .A(n20823), .B(n20822), .ZN(
        P1_U3092) );
  AOI22_X1 U23755 ( .A1(n21105), .A2(n20833), .B1(n21104), .B2(n20832), .ZN(
        n20825) );
  AOI22_X1 U23756 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20834), .B1(
        n20828), .B2(n21045), .ZN(n20824) );
  OAI211_X1 U23757 ( .C1(n21048), .C2(n20831), .A(n20825), .B(n20824), .ZN(
        P1_U3093) );
  AOI22_X1 U23758 ( .A1(n21111), .A2(n20833), .B1(n9565), .B2(n20832), .ZN(
        n20827) );
  AOI22_X1 U23759 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20834), .B1(
        n20862), .B2(n21112), .ZN(n20826) );
  OAI211_X1 U23760 ( .C1(n21115), .C2(n20837), .A(n20827), .B(n20826), .ZN(
        P1_U3094) );
  AOI22_X1 U23761 ( .A1(n21117), .A2(n20833), .B1(n21116), .B2(n20832), .ZN(
        n20830) );
  AOI22_X1 U23762 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20834), .B1(
        n20828), .B2(n21053), .ZN(n20829) );
  OAI211_X1 U23763 ( .C1(n21056), .C2(n20831), .A(n20830), .B(n20829), .ZN(
        P1_U3095) );
  AOI22_X1 U23764 ( .A1(n21125), .A2(n20833), .B1(n9567), .B2(n20832), .ZN(
        n20836) );
  AOI22_X1 U23765 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20834), .B1(
        n20862), .B2(n21126), .ZN(n20835) );
  OAI211_X1 U23766 ( .C1(n21132), .C2(n20837), .A(n20836), .B(n20835), .ZN(
        P1_U3096) );
  INV_X1 U23767 ( .A(n20959), .ZN(n20838) );
  NAND2_X1 U23768 ( .A1(n20839), .A2(n13947), .ZN(n20896) );
  INV_X1 U23769 ( .A(n20896), .ZN(n20930) );
  NAND2_X1 U23770 ( .A1(n20840), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20929) );
  AOI21_X1 U23771 ( .B1(n20930), .B2(n14960), .A(n10412), .ZN(n20844) );
  NAND2_X1 U23772 ( .A1(n20842), .A2(n20841), .ZN(n20965) );
  OAI22_X1 U23773 ( .A1(n20844), .A2(n21075), .B1(n20902), .B2(n20965), .ZN(
        n20861) );
  AOI22_X1 U23774 ( .A1(n21073), .A2(n20861), .B1(n21072), .B2(n10412), .ZN(
        n20848) );
  INV_X1 U23775 ( .A(n20892), .ZN(n20843) );
  OAI21_X1 U23776 ( .B1(n20843), .B2(n20862), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20845) );
  NAND2_X1 U23777 ( .A1(n20845), .A2(n20844), .ZN(n20846) );
  AOI22_X1 U23778 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20863), .B1(
        n20862), .B2(n21029), .ZN(n20847) );
  OAI211_X1 U23779 ( .C1(n21032), .C2(n20892), .A(n20848), .B(n20847), .ZN(
        P1_U3097) );
  AOI22_X1 U23780 ( .A1(n21087), .A2(n20861), .B1(n21086), .B2(n10412), .ZN(
        n20850) );
  AOI22_X1 U23781 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20863), .B1(
        n20862), .B2(n21033), .ZN(n20849) );
  OAI211_X1 U23782 ( .C1(n21036), .C2(n20892), .A(n20850), .B(n20849), .ZN(
        P1_U3098) );
  AOI22_X1 U23783 ( .A1(n21093), .A2(n20861), .B1(n21092), .B2(n10412), .ZN(
        n20852) );
  AOI22_X1 U23784 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20863), .B1(
        n20862), .B2(n21037), .ZN(n20851) );
  OAI211_X1 U23785 ( .C1(n21040), .C2(n20892), .A(n20852), .B(n20851), .ZN(
        P1_U3099) );
  AOI22_X1 U23786 ( .A1(n21099), .A2(n20861), .B1(n21098), .B2(n10412), .ZN(
        n20854) );
  AOI22_X1 U23787 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20863), .B1(
        n20862), .B2(n21041), .ZN(n20853) );
  OAI211_X1 U23788 ( .C1(n21044), .C2(n20892), .A(n20854), .B(n20853), .ZN(
        P1_U3100) );
  AOI22_X1 U23789 ( .A1(n21105), .A2(n20861), .B1(n21104), .B2(n10412), .ZN(
        n20856) );
  AOI22_X1 U23790 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20863), .B1(
        n20862), .B2(n21045), .ZN(n20855) );
  OAI211_X1 U23791 ( .C1(n21048), .C2(n20892), .A(n20856), .B(n20855), .ZN(
        P1_U3101) );
  AOI22_X1 U23792 ( .A1(n21111), .A2(n20861), .B1(n9565), .B2(n10412), .ZN(
        n20858) );
  AOI22_X1 U23793 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20863), .B1(
        n20862), .B2(n21049), .ZN(n20857) );
  OAI211_X1 U23794 ( .C1(n21052), .C2(n20892), .A(n20858), .B(n20857), .ZN(
        P1_U3102) );
  AOI22_X1 U23795 ( .A1(n21117), .A2(n20861), .B1(n21116), .B2(n10412), .ZN(
        n20860) );
  AOI22_X1 U23796 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20863), .B1(
        n20862), .B2(n21053), .ZN(n20859) );
  OAI211_X1 U23797 ( .C1(n21056), .C2(n20892), .A(n20860), .B(n20859), .ZN(
        P1_U3103) );
  AOI22_X1 U23798 ( .A1(n21125), .A2(n20861), .B1(n9567), .B2(n10412), .ZN(
        n20865) );
  AOI22_X1 U23799 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20863), .B1(
        n20862), .B2(n21059), .ZN(n20864) );
  OAI211_X1 U23800 ( .C1(n21064), .C2(n20892), .A(n20865), .B(n20864), .ZN(
        P1_U3104) );
  NOR2_X1 U23801 ( .A1(n20929), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20870) );
  INV_X1 U23802 ( .A(n20870), .ZN(n20867) );
  NOR2_X1 U23803 ( .A1(n20988), .A2(n20867), .ZN(n20887) );
  INV_X1 U23804 ( .A(n20887), .ZN(n20866) );
  OAI222_X1 U23805 ( .A1(n20868), .A2(n20896), .B1(n21070), .B2(n20867), .C1(
        n21075), .C2(n20866), .ZN(n20888) );
  AOI22_X1 U23806 ( .A1(n21073), .A2(n20888), .B1(n21072), .B2(n20887), .ZN(
        n20874) );
  NOR2_X1 U23807 ( .A1(n20934), .A2(n20869), .ZN(n20871) );
  NAND2_X1 U23808 ( .A1(n20928), .A2(n20872), .ZN(n20919) );
  AOI22_X1 U23809 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20889), .B1(
        n20921), .B2(n21082), .ZN(n20873) );
  OAI211_X1 U23810 ( .C1(n21085), .C2(n20892), .A(n20874), .B(n20873), .ZN(
        P1_U3105) );
  AOI22_X1 U23811 ( .A1(n21087), .A2(n20888), .B1(n21086), .B2(n20887), .ZN(
        n20876) );
  AOI22_X1 U23812 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20889), .B1(
        n20921), .B2(n21088), .ZN(n20875) );
  OAI211_X1 U23813 ( .C1(n21091), .C2(n20892), .A(n20876), .B(n20875), .ZN(
        P1_U3106) );
  AOI22_X1 U23814 ( .A1(n21093), .A2(n20888), .B1(n21092), .B2(n20887), .ZN(
        n20878) );
  AOI22_X1 U23815 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20889), .B1(
        n20921), .B2(n21094), .ZN(n20877) );
  OAI211_X1 U23816 ( .C1(n21097), .C2(n20892), .A(n20878), .B(n20877), .ZN(
        P1_U3107) );
  AOI22_X1 U23817 ( .A1(n21099), .A2(n20888), .B1(n21098), .B2(n20887), .ZN(
        n20880) );
  AOI22_X1 U23818 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20889), .B1(
        n20921), .B2(n21100), .ZN(n20879) );
  OAI211_X1 U23819 ( .C1(n21103), .C2(n20892), .A(n20880), .B(n20879), .ZN(
        P1_U3108) );
  AOI22_X1 U23820 ( .A1(n21105), .A2(n20888), .B1(n21104), .B2(n20887), .ZN(
        n20882) );
  AOI22_X1 U23821 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20889), .B1(
        n20921), .B2(n21106), .ZN(n20881) );
  OAI211_X1 U23822 ( .C1(n21109), .C2(n20892), .A(n20882), .B(n20881), .ZN(
        P1_U3109) );
  AOI22_X1 U23823 ( .A1(n21111), .A2(n20888), .B1(n9565), .B2(n20887), .ZN(
        n20884) );
  AOI22_X1 U23824 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20889), .B1(
        n20921), .B2(n21112), .ZN(n20883) );
  OAI211_X1 U23825 ( .C1(n21115), .C2(n20892), .A(n20884), .B(n20883), .ZN(
        P1_U3110) );
  AOI22_X1 U23826 ( .A1(n21117), .A2(n20888), .B1(n21116), .B2(n20887), .ZN(
        n20886) );
  AOI22_X1 U23827 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20889), .B1(
        n20921), .B2(n21118), .ZN(n20885) );
  OAI211_X1 U23828 ( .C1(n21121), .C2(n20892), .A(n20886), .B(n20885), .ZN(
        P1_U3111) );
  AOI22_X1 U23829 ( .A1(n21125), .A2(n20888), .B1(n9567), .B2(n20887), .ZN(
        n20891) );
  AOI22_X1 U23830 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20889), .B1(
        n20921), .B2(n21126), .ZN(n20890) );
  OAI211_X1 U23831 ( .C1(n21132), .C2(n20892), .A(n20891), .B(n20890), .ZN(
        P1_U3112) );
  INV_X1 U23832 ( .A(n20929), .ZN(n20894) );
  NAND2_X1 U23833 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20894), .ZN(
        n20932) );
  NOR2_X1 U23834 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20932), .ZN(
        n20920) );
  AOI22_X1 U23835 ( .A1(n20921), .A2(n21029), .B1(n21072), .B2(n20920), .ZN(
        n20906) );
  AOI21_X1 U23836 ( .B1(n20957), .B2(n20919), .A(n21022), .ZN(n20895) );
  NOR2_X1 U23837 ( .A1(n20895), .A2(n21075), .ZN(n20901) );
  OR2_X1 U23838 ( .A1(n20896), .A2(n14960), .ZN(n20903) );
  NAND2_X1 U23839 ( .A1(n20897), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21018) );
  NAND2_X1 U23840 ( .A1(n21018), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21026) );
  OAI211_X1 U23841 ( .C1(n20963), .C2(n20920), .A(n21026), .B(n20898), .ZN(
        n20899) );
  AOI21_X1 U23842 ( .B1(n20901), .B2(n20903), .A(n20899), .ZN(n20900) );
  INV_X1 U23843 ( .A(n20901), .ZN(n20904) );
  AOI22_X1 U23844 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20923), .B1(
        n21073), .B2(n20922), .ZN(n20905) );
  OAI211_X1 U23845 ( .C1(n21032), .C2(n20957), .A(n20906), .B(n20905), .ZN(
        P1_U3113) );
  AOI22_X1 U23846 ( .A1(n20946), .A2(n21088), .B1(n21086), .B2(n20920), .ZN(
        n20908) );
  AOI22_X1 U23847 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20923), .B1(
        n21087), .B2(n20922), .ZN(n20907) );
  OAI211_X1 U23848 ( .C1(n21091), .C2(n20919), .A(n20908), .B(n20907), .ZN(
        P1_U3114) );
  AOI22_X1 U23849 ( .A1(n20921), .A2(n21037), .B1(n21092), .B2(n20920), .ZN(
        n20910) );
  AOI22_X1 U23850 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20923), .B1(
        n21093), .B2(n20922), .ZN(n20909) );
  OAI211_X1 U23851 ( .C1(n21040), .C2(n20957), .A(n20910), .B(n20909), .ZN(
        P1_U3115) );
  AOI22_X1 U23852 ( .A1(n20921), .A2(n21041), .B1(n21098), .B2(n20920), .ZN(
        n20912) );
  AOI22_X1 U23853 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20923), .B1(
        n21099), .B2(n20922), .ZN(n20911) );
  OAI211_X1 U23854 ( .C1(n21044), .C2(n20957), .A(n20912), .B(n20911), .ZN(
        P1_U3116) );
  AOI22_X1 U23855 ( .A1(n20946), .A2(n21106), .B1(n21104), .B2(n20920), .ZN(
        n20914) );
  AOI22_X1 U23856 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20923), .B1(
        n21105), .B2(n20922), .ZN(n20913) );
  OAI211_X1 U23857 ( .C1(n21109), .C2(n20919), .A(n20914), .B(n20913), .ZN(
        P1_U3117) );
  AOI22_X1 U23858 ( .A1(n20921), .A2(n21049), .B1(n9565), .B2(n20920), .ZN(
        n20916) );
  AOI22_X1 U23859 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20923), .B1(
        n21111), .B2(n20922), .ZN(n20915) );
  OAI211_X1 U23860 ( .C1(n21052), .C2(n20957), .A(n20916), .B(n20915), .ZN(
        P1_U3118) );
  AOI22_X1 U23861 ( .A1(n20946), .A2(n21118), .B1(n21116), .B2(n20920), .ZN(
        n20918) );
  AOI22_X1 U23862 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20923), .B1(
        n21117), .B2(n20922), .ZN(n20917) );
  OAI211_X1 U23863 ( .C1(n21121), .C2(n20919), .A(n20918), .B(n20917), .ZN(
        P1_U3119) );
  AOI22_X1 U23864 ( .A1(n20921), .A2(n21059), .B1(n9567), .B2(n20920), .ZN(
        n20925) );
  AOI22_X1 U23865 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20923), .B1(
        n21125), .B2(n20922), .ZN(n20924) );
  OAI211_X1 U23866 ( .C1(n21064), .C2(n20957), .A(n20925), .B(n20924), .ZN(
        P1_U3120) );
  INV_X1 U23867 ( .A(n20926), .ZN(n20927) );
  NOR2_X1 U23868 ( .A1(n21065), .A2(n20929), .ZN(n20951) );
  AOI21_X1 U23869 ( .B1(n20930), .B2(n21066), .A(n20951), .ZN(n20931) );
  OAI22_X1 U23870 ( .A1(n20931), .A2(n21075), .B1(n20932), .B2(n21070), .ZN(
        n20952) );
  AOI22_X1 U23871 ( .A1(n21073), .A2(n20952), .B1(n21072), .B2(n20951), .ZN(
        n20937) );
  OAI21_X1 U23872 ( .B1(n20934), .B2(n20933), .A(n20932), .ZN(n20935) );
  NAND2_X1 U23873 ( .A1(n20935), .A2(n21080), .ZN(n20954) );
  AOI22_X1 U23874 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20954), .B1(
        n20946), .B2(n21029), .ZN(n20936) );
  OAI211_X1 U23875 ( .C1(n21032), .C2(n20987), .A(n20937), .B(n20936), .ZN(
        P1_U3121) );
  AOI22_X1 U23876 ( .A1(n21087), .A2(n20952), .B1(n21086), .B2(n20951), .ZN(
        n20939) );
  INV_X1 U23877 ( .A(n20987), .ZN(n20953) );
  AOI22_X1 U23878 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20954), .B1(
        n20953), .B2(n21088), .ZN(n20938) );
  OAI211_X1 U23879 ( .C1(n21091), .C2(n20957), .A(n20939), .B(n20938), .ZN(
        P1_U3122) );
  AOI22_X1 U23880 ( .A1(n21093), .A2(n20952), .B1(n21092), .B2(n20951), .ZN(
        n20941) );
  AOI22_X1 U23881 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20954), .B1(
        n20946), .B2(n21037), .ZN(n20940) );
  OAI211_X1 U23882 ( .C1(n21040), .C2(n20987), .A(n20941), .B(n20940), .ZN(
        P1_U3123) );
  AOI22_X1 U23883 ( .A1(n21099), .A2(n20952), .B1(n21098), .B2(n20951), .ZN(
        n20943) );
  AOI22_X1 U23884 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20954), .B1(
        n20953), .B2(n21100), .ZN(n20942) );
  OAI211_X1 U23885 ( .C1(n21103), .C2(n20957), .A(n20943), .B(n20942), .ZN(
        P1_U3124) );
  AOI22_X1 U23886 ( .A1(n21105), .A2(n20952), .B1(n21104), .B2(n20951), .ZN(
        n20945) );
  AOI22_X1 U23887 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20954), .B1(
        n20953), .B2(n21106), .ZN(n20944) );
  OAI211_X1 U23888 ( .C1(n21109), .C2(n20957), .A(n20945), .B(n20944), .ZN(
        P1_U3125) );
  AOI22_X1 U23889 ( .A1(n21111), .A2(n20952), .B1(n9565), .B2(n20951), .ZN(
        n20948) );
  AOI22_X1 U23890 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20954), .B1(
        n20946), .B2(n21049), .ZN(n20947) );
  OAI211_X1 U23891 ( .C1(n21052), .C2(n20987), .A(n20948), .B(n20947), .ZN(
        P1_U3126) );
  AOI22_X1 U23892 ( .A1(n21117), .A2(n20952), .B1(n21116), .B2(n20951), .ZN(
        n20950) );
  AOI22_X1 U23893 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20954), .B1(
        n20953), .B2(n21118), .ZN(n20949) );
  OAI211_X1 U23894 ( .C1(n21121), .C2(n20957), .A(n20950), .B(n20949), .ZN(
        P1_U3127) );
  AOI22_X1 U23895 ( .A1(n21125), .A2(n20952), .B1(n9567), .B2(n20951), .ZN(
        n20956) );
  AOI22_X1 U23896 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20954), .B1(
        n20953), .B2(n21126), .ZN(n20955) );
  OAI211_X1 U23897 ( .C1(n21132), .C2(n20957), .A(n20956), .B(n20955), .ZN(
        P1_U3128) );
  NAND2_X1 U23898 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21068) );
  AOI22_X1 U23899 ( .A1(n21072), .A2(n10418), .B1(n20982), .B2(n21082), .ZN(
        n20969) );
  NAND2_X1 U23900 ( .A1(n20987), .A2(n21015), .ZN(n20960) );
  AOI21_X1 U23901 ( .B1(n20960), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n21075), 
        .ZN(n20964) );
  OR2_X1 U23902 ( .A1(n13947), .A2(n20961), .ZN(n21021) );
  OR2_X1 U23903 ( .A1(n21021), .A2(n10366), .ZN(n20966) );
  AOI22_X1 U23904 ( .A1(n20964), .A2(n20966), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20965), .ZN(n20962) );
  INV_X1 U23905 ( .A(n20964), .ZN(n20967) );
  AOI22_X1 U23906 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20984), .B1(
        n21073), .B2(n20983), .ZN(n20968) );
  OAI211_X1 U23907 ( .C1(n21085), .C2(n20987), .A(n20969), .B(n20968), .ZN(
        P1_U3129) );
  AOI22_X1 U23908 ( .A1(n21086), .A2(n10418), .B1(n20982), .B2(n21088), .ZN(
        n20971) );
  AOI22_X1 U23909 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20984), .B1(
        n21087), .B2(n20983), .ZN(n20970) );
  OAI211_X1 U23910 ( .C1(n21091), .C2(n20987), .A(n20971), .B(n20970), .ZN(
        P1_U3130) );
  AOI22_X1 U23911 ( .A1(n21092), .A2(n10418), .B1(n20982), .B2(n21094), .ZN(
        n20973) );
  AOI22_X1 U23912 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20984), .B1(
        n21093), .B2(n20983), .ZN(n20972) );
  OAI211_X1 U23913 ( .C1(n21097), .C2(n20987), .A(n20973), .B(n20972), .ZN(
        P1_U3131) );
  AOI22_X1 U23914 ( .A1(n21098), .A2(n10418), .B1(n20982), .B2(n21100), .ZN(
        n20975) );
  AOI22_X1 U23915 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20984), .B1(
        n21099), .B2(n20983), .ZN(n20974) );
  OAI211_X1 U23916 ( .C1(n21103), .C2(n20987), .A(n20975), .B(n20974), .ZN(
        P1_U3132) );
  AOI22_X1 U23917 ( .A1(n21104), .A2(n10418), .B1(n20982), .B2(n21106), .ZN(
        n20977) );
  AOI22_X1 U23918 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20984), .B1(
        n21105), .B2(n20983), .ZN(n20976) );
  OAI211_X1 U23919 ( .C1(n21109), .C2(n20987), .A(n20977), .B(n20976), .ZN(
        P1_U3133) );
  AOI22_X1 U23920 ( .A1(n9565), .A2(n10418), .B1(n20982), .B2(n21112), .ZN(
        n20979) );
  AOI22_X1 U23921 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20984), .B1(
        n21111), .B2(n20983), .ZN(n20978) );
  OAI211_X1 U23922 ( .C1(n21115), .C2(n20987), .A(n20979), .B(n20978), .ZN(
        P1_U3134) );
  AOI22_X1 U23923 ( .A1(n21116), .A2(n10418), .B1(n20982), .B2(n21118), .ZN(
        n20981) );
  AOI22_X1 U23924 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20984), .B1(
        n21117), .B2(n20983), .ZN(n20980) );
  OAI211_X1 U23925 ( .C1(n21121), .C2(n20987), .A(n20981), .B(n20980), .ZN(
        P1_U3135) );
  AOI22_X1 U23926 ( .A1(n9567), .A2(n10418), .B1(n20982), .B2(n21126), .ZN(
        n20986) );
  AOI22_X1 U23927 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20984), .B1(
        n21125), .B2(n20983), .ZN(n20985) );
  OAI211_X1 U23928 ( .C1(n21132), .C2(n20987), .A(n20986), .B(n20985), .ZN(
        P1_U3136) );
  INV_X1 U23929 ( .A(n21021), .ZN(n21067) );
  INV_X1 U23930 ( .A(n20635), .ZN(n20989) );
  NOR3_X2 U23931 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20988), .A3(
        n21068), .ZN(n21010) );
  AOI21_X1 U23932 ( .B1(n21067), .B2(n20989), .A(n21010), .ZN(n20991) );
  NOR2_X1 U23933 ( .A1(n21068), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20994) );
  INV_X1 U23934 ( .A(n20994), .ZN(n20990) );
  OAI22_X1 U23935 ( .A1(n20991), .A2(n21075), .B1(n20990), .B2(n21070), .ZN(
        n21011) );
  AOI22_X1 U23936 ( .A1(n21073), .A2(n21011), .B1(n21072), .B2(n21010), .ZN(
        n20997) );
  INV_X1 U23937 ( .A(n21017), .ZN(n21076) );
  NAND2_X1 U23938 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n21076), .ZN(n20992) );
  NAND2_X1 U23939 ( .A1(n20992), .A2(n20991), .ZN(n20993) );
  AOI22_X1 U23940 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n21012), .B1(
        n21060), .B2(n21082), .ZN(n20996) );
  OAI211_X1 U23941 ( .C1(n21085), .C2(n21015), .A(n20997), .B(n20996), .ZN(
        P1_U3137) );
  AOI22_X1 U23942 ( .A1(n21087), .A2(n21011), .B1(n21086), .B2(n21010), .ZN(
        n20999) );
  AOI22_X1 U23943 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n21012), .B1(
        n21060), .B2(n21088), .ZN(n20998) );
  OAI211_X1 U23944 ( .C1(n21091), .C2(n21015), .A(n20999), .B(n20998), .ZN(
        P1_U3138) );
  AOI22_X1 U23945 ( .A1(n21093), .A2(n21011), .B1(n21092), .B2(n21010), .ZN(
        n21001) );
  AOI22_X1 U23946 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n21012), .B1(
        n21060), .B2(n21094), .ZN(n21000) );
  OAI211_X1 U23947 ( .C1(n21097), .C2(n21015), .A(n21001), .B(n21000), .ZN(
        P1_U3139) );
  AOI22_X1 U23948 ( .A1(n21099), .A2(n21011), .B1(n21098), .B2(n21010), .ZN(
        n21003) );
  AOI22_X1 U23949 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n21012), .B1(
        n21060), .B2(n21100), .ZN(n21002) );
  OAI211_X1 U23950 ( .C1(n21103), .C2(n21015), .A(n21003), .B(n21002), .ZN(
        P1_U3140) );
  AOI22_X1 U23951 ( .A1(n21105), .A2(n21011), .B1(n21104), .B2(n21010), .ZN(
        n21005) );
  AOI22_X1 U23952 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n21012), .B1(
        n21060), .B2(n21106), .ZN(n21004) );
  OAI211_X1 U23953 ( .C1(n21109), .C2(n21015), .A(n21005), .B(n21004), .ZN(
        P1_U3141) );
  AOI22_X1 U23954 ( .A1(n21111), .A2(n21011), .B1(n9565), .B2(n21010), .ZN(
        n21007) );
  AOI22_X1 U23955 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n21012), .B1(
        n21060), .B2(n21112), .ZN(n21006) );
  OAI211_X1 U23956 ( .C1(n21115), .C2(n21015), .A(n21007), .B(n21006), .ZN(
        P1_U3142) );
  AOI22_X1 U23957 ( .A1(n21117), .A2(n21011), .B1(n21116), .B2(n21010), .ZN(
        n21009) );
  AOI22_X1 U23958 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n21012), .B1(
        n21060), .B2(n21118), .ZN(n21008) );
  OAI211_X1 U23959 ( .C1(n21121), .C2(n21015), .A(n21009), .B(n21008), .ZN(
        P1_U3143) );
  AOI22_X1 U23960 ( .A1(n21125), .A2(n21011), .B1(n9567), .B2(n21010), .ZN(
        n21014) );
  AOI22_X1 U23961 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n21012), .B1(
        n21060), .B2(n21126), .ZN(n21013) );
  OAI211_X1 U23962 ( .C1(n21132), .C2(n21015), .A(n21014), .B(n21013), .ZN(
        P1_U3144) );
  NAND2_X1 U23963 ( .A1(n10366), .A2(n21383), .ZN(n21020) );
  OAI22_X1 U23964 ( .A1(n21021), .A2(n21020), .B1(n21019), .B2(n21018), .ZN(
        n21058) );
  NOR3_X2 U23965 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21069), .A3(
        n21068), .ZN(n21057) );
  AOI22_X1 U23966 ( .A1(n21073), .A2(n21058), .B1(n21072), .B2(n21057), .ZN(
        n21031) );
  INV_X1 U23967 ( .A(n21060), .ZN(n21023) );
  AOI21_X1 U23968 ( .B1(n21023), .B2(n21131), .A(n21022), .ZN(n21024) );
  AOI21_X1 U23969 ( .B1(n21067), .B2(n10366), .A(n21024), .ZN(n21025) );
  NOR2_X1 U23970 ( .A1(n21025), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21028) );
  AOI22_X1 U23971 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n21061), .B1(
        n21060), .B2(n21029), .ZN(n21030) );
  OAI211_X1 U23972 ( .C1(n21032), .C2(n21131), .A(n21031), .B(n21030), .ZN(
        P1_U3145) );
  AOI22_X1 U23973 ( .A1(n21087), .A2(n21058), .B1(n21086), .B2(n21057), .ZN(
        n21035) );
  AOI22_X1 U23974 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n21061), .B1(
        n21060), .B2(n21033), .ZN(n21034) );
  OAI211_X1 U23975 ( .C1(n21036), .C2(n21131), .A(n21035), .B(n21034), .ZN(
        P1_U3146) );
  AOI22_X1 U23976 ( .A1(n21093), .A2(n21058), .B1(n21092), .B2(n21057), .ZN(
        n21039) );
  AOI22_X1 U23977 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n21061), .B1(
        n21060), .B2(n21037), .ZN(n21038) );
  OAI211_X1 U23978 ( .C1(n21040), .C2(n21131), .A(n21039), .B(n21038), .ZN(
        P1_U3147) );
  AOI22_X1 U23979 ( .A1(n21099), .A2(n21058), .B1(n21098), .B2(n21057), .ZN(
        n21043) );
  AOI22_X1 U23980 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n21061), .B1(
        n21060), .B2(n21041), .ZN(n21042) );
  OAI211_X1 U23981 ( .C1(n21044), .C2(n21131), .A(n21043), .B(n21042), .ZN(
        P1_U3148) );
  AOI22_X1 U23982 ( .A1(n21105), .A2(n21058), .B1(n21104), .B2(n21057), .ZN(
        n21047) );
  AOI22_X1 U23983 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n21061), .B1(
        n21060), .B2(n21045), .ZN(n21046) );
  OAI211_X1 U23984 ( .C1(n21048), .C2(n21131), .A(n21047), .B(n21046), .ZN(
        P1_U3149) );
  AOI22_X1 U23985 ( .A1(n21111), .A2(n21058), .B1(n9565), .B2(n21057), .ZN(
        n21051) );
  AOI22_X1 U23986 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n21061), .B1(
        n21060), .B2(n21049), .ZN(n21050) );
  OAI211_X1 U23987 ( .C1(n21052), .C2(n21131), .A(n21051), .B(n21050), .ZN(
        P1_U3150) );
  AOI22_X1 U23988 ( .A1(n21117), .A2(n21058), .B1(n21116), .B2(n21057), .ZN(
        n21055) );
  AOI22_X1 U23989 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n21061), .B1(
        n21060), .B2(n21053), .ZN(n21054) );
  OAI211_X1 U23990 ( .C1(n21056), .C2(n21131), .A(n21055), .B(n21054), .ZN(
        P1_U3151) );
  AOI22_X1 U23991 ( .A1(n21125), .A2(n21058), .B1(n9567), .B2(n21057), .ZN(
        n21063) );
  AOI22_X1 U23992 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n21061), .B1(
        n21060), .B2(n21059), .ZN(n21062) );
  OAI211_X1 U23993 ( .C1(n21064), .C2(n21131), .A(n21063), .B(n21062), .ZN(
        P1_U3152) );
  NOR2_X1 U23994 ( .A1(n21065), .A2(n21068), .ZN(n21122) );
  AOI21_X1 U23995 ( .B1(n21067), .B2(n21066), .A(n21122), .ZN(n21077) );
  NOR2_X1 U23996 ( .A1(n21069), .A2(n21068), .ZN(n21081) );
  INV_X1 U23997 ( .A(n21081), .ZN(n21071) );
  OAI22_X1 U23998 ( .A1(n21077), .A2(n21075), .B1(n21071), .B2(n21070), .ZN(
        n21124) );
  AOI22_X1 U23999 ( .A1(n21073), .A2(n21124), .B1(n21072), .B2(n21122), .ZN(
        n21084) );
  OAI21_X1 U24000 ( .B1(n21076), .B2(n21075), .A(n21074), .ZN(n21078) );
  NAND2_X1 U24001 ( .A1(n21078), .A2(n21077), .ZN(n21079) );
  AOI22_X1 U24002 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n21128), .B1(
        n21127), .B2(n21082), .ZN(n21083) );
  OAI211_X1 U24003 ( .C1(n21085), .C2(n21131), .A(n21084), .B(n21083), .ZN(
        P1_U3153) );
  AOI22_X1 U24004 ( .A1(n21087), .A2(n21124), .B1(n21086), .B2(n21122), .ZN(
        n21090) );
  AOI22_X1 U24005 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n21128), .B1(
        n21127), .B2(n21088), .ZN(n21089) );
  OAI211_X1 U24006 ( .C1(n21091), .C2(n21131), .A(n21090), .B(n21089), .ZN(
        P1_U3154) );
  AOI22_X1 U24007 ( .A1(n21093), .A2(n21124), .B1(n21092), .B2(n21122), .ZN(
        n21096) );
  AOI22_X1 U24008 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n21128), .B1(
        n21127), .B2(n21094), .ZN(n21095) );
  OAI211_X1 U24009 ( .C1(n21097), .C2(n21131), .A(n21096), .B(n21095), .ZN(
        P1_U3155) );
  AOI22_X1 U24010 ( .A1(n21099), .A2(n21124), .B1(n21098), .B2(n21122), .ZN(
        n21102) );
  AOI22_X1 U24011 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n21128), .B1(
        n21127), .B2(n21100), .ZN(n21101) );
  OAI211_X1 U24012 ( .C1(n21103), .C2(n21131), .A(n21102), .B(n21101), .ZN(
        P1_U3156) );
  AOI22_X1 U24013 ( .A1(n21105), .A2(n21124), .B1(n21104), .B2(n21122), .ZN(
        n21108) );
  AOI22_X1 U24014 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n21128), .B1(
        n21127), .B2(n21106), .ZN(n21107) );
  OAI211_X1 U24015 ( .C1(n21109), .C2(n21131), .A(n21108), .B(n21107), .ZN(
        P1_U3157) );
  AOI22_X1 U24016 ( .A1(n21111), .A2(n21124), .B1(n9565), .B2(n21122), .ZN(
        n21114) );
  AOI22_X1 U24017 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n21128), .B1(
        n21127), .B2(n21112), .ZN(n21113) );
  OAI211_X1 U24018 ( .C1(n21115), .C2(n21131), .A(n21114), .B(n21113), .ZN(
        P1_U3158) );
  AOI22_X1 U24019 ( .A1(n21117), .A2(n21124), .B1(n21116), .B2(n21122), .ZN(
        n21120) );
  AOI22_X1 U24020 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n21128), .B1(
        n21127), .B2(n21118), .ZN(n21119) );
  OAI211_X1 U24021 ( .C1(n21121), .C2(n21131), .A(n21120), .B(n21119), .ZN(
        P1_U3159) );
  AOI22_X1 U24022 ( .A1(n21125), .A2(n21124), .B1(n9567), .B2(n21122), .ZN(
        n21130) );
  AOI22_X1 U24023 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n21128), .B1(
        n21127), .B2(n21126), .ZN(n21129) );
  OAI211_X1 U24024 ( .C1(n21132), .C2(n21131), .A(n21130), .B(n21129), .ZN(
        P1_U3160) );
  NAND3_X1 U24025 ( .A1(n21135), .A2(n21134), .A3(n21133), .ZN(P1_U3163) );
  AND2_X1 U24026 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n21136), .ZN(
        P1_U3164) );
  AND2_X1 U24027 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n21136), .ZN(
        P1_U3165) );
  AND2_X1 U24028 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n21136), .ZN(
        P1_U3166) );
  AND2_X1 U24029 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n21136), .ZN(
        P1_U3167) );
  AND2_X1 U24030 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n21136), .ZN(
        P1_U3168) );
  AND2_X1 U24031 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n21136), .ZN(
        P1_U3169) );
  AND2_X1 U24032 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n21136), .ZN(
        P1_U3170) );
  AND2_X1 U24033 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n21136), .ZN(
        P1_U3171) );
  AND2_X1 U24034 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n21136), .ZN(
        P1_U3172) );
  AND2_X1 U24035 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n21136), .ZN(
        P1_U3173) );
  AND2_X1 U24036 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n21136), .ZN(
        P1_U3174) );
  AND2_X1 U24037 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n21136), .ZN(
        P1_U3175) );
  AND2_X1 U24038 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n21136), .ZN(
        P1_U3176) );
  INV_X1 U24039 ( .A(P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n21344) );
  NOR2_X1 U24040 ( .A1(n21204), .A2(n21344), .ZN(P1_U3177) );
  AND2_X1 U24041 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n21136), .ZN(
        P1_U3178) );
  AND2_X1 U24042 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n21136), .ZN(
        P1_U3179) );
  AND2_X1 U24043 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n21136), .ZN(
        P1_U3180) );
  AND2_X1 U24044 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n21136), .ZN(
        P1_U3181) );
  AND2_X1 U24045 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n21136), .ZN(
        P1_U3182) );
  INV_X1 U24046 ( .A(P1_DATAWIDTH_REG_12__SCAN_IN), .ZN(n21255) );
  NOR2_X1 U24047 ( .A1(n21204), .A2(n21255), .ZN(P1_U3183) );
  AND2_X1 U24048 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n21136), .ZN(
        P1_U3184) );
  AND2_X1 U24049 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n21136), .ZN(
        P1_U3185) );
  AND2_X1 U24050 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n21136), .ZN(P1_U3186) );
  AND2_X1 U24051 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n21136), .ZN(P1_U3187) );
  AND2_X1 U24052 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n21136), .ZN(P1_U3188) );
  AND2_X1 U24053 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n21136), .ZN(P1_U3189) );
  AND2_X1 U24054 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n21136), .ZN(P1_U3190) );
  AND2_X1 U24055 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n21136), .ZN(P1_U3191) );
  INV_X1 U24056 ( .A(P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n21256) );
  NOR2_X1 U24057 ( .A1(n21204), .A2(n21256), .ZN(P1_U3192) );
  INV_X1 U24058 ( .A(P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n21352) );
  NOR2_X1 U24059 ( .A1(n21204), .A2(n21352), .ZN(P1_U3193) );
  AOI21_X1 U24060 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21142), .A(n21137), 
        .ZN(n21145) );
  NAND2_X1 U24061 ( .A1(n21151), .A2(n21150), .ZN(n21139) );
  OAI21_X1 U24062 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n21141), .A(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21138) );
  AOI21_X1 U24063 ( .B1(HOLD), .B2(n21139), .A(n21138), .ZN(n21140) );
  OAI22_X1 U24064 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21145), .B1(n21214), 
        .B2(n21140), .ZN(P1_U3194) );
  NAND4_X1 U24065 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21142), .A3(
        P1_REQUESTPENDING_REG_SCAN_IN), .A4(n21141), .ZN(n21149) );
  NAND2_X1 U24066 ( .A1(n21142), .A2(n21141), .ZN(n21143) );
  OAI221_X1 U24067 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(
        P1_STATE_REG_1__SCAN_IN), .C1(P1_REQUESTPENDING_REG_SCAN_IN), .C2(
        n21143), .A(n21151), .ZN(n21144) );
  NAND3_X1 U24068 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(HOLD), .A3(n21144), .ZN(
        n21148) );
  AOI211_X1 U24069 ( .C1(n21150), .C2(NA), .A(n21151), .B(n21145), .ZN(n21146)
         );
  INV_X1 U24070 ( .A(n21146), .ZN(n21147) );
  OAI211_X1 U24071 ( .C1(n21150), .C2(n21149), .A(n21148), .B(n21147), .ZN(
        P1_U3196) );
  NAND2_X1 U24072 ( .A1(n21151), .A2(n21214), .ZN(n21182) );
  AOI22_X1 U24073 ( .A1(P1_ADDRESS_REG_0__SCAN_IN), .A2(n21198), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n21193), .ZN(n21152) );
  OAI21_X1 U24074 ( .B1(n21206), .B2(n21179), .A(n21152), .ZN(P1_U3197) );
  INV_X1 U24075 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n21154) );
  AOI22_X1 U24076 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(n21198), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n21193), .ZN(n21153) );
  OAI21_X1 U24077 ( .B1(n21154), .B2(n21179), .A(n21153), .ZN(P1_U3198) );
  INV_X1 U24078 ( .A(n21179), .ZN(n21194) );
  AOI222_X1 U24079 ( .A1(n21194), .A2(P1_REIP_REG_3__SCAN_IN), .B1(
        P1_ADDRESS_REG_2__SCAN_IN), .B2(n21198), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n21193), .ZN(n21155) );
  INV_X1 U24080 ( .A(n21155), .ZN(P1_U3199) );
  AOI22_X1 U24081 ( .A1(P1_ADDRESS_REG_3__SCAN_IN), .A2(n21198), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n21193), .ZN(n21156) );
  OAI21_X1 U24082 ( .B1(n21157), .B2(n21179), .A(n21156), .ZN(P1_U3200) );
  AOI22_X1 U24083 ( .A1(P1_ADDRESS_REG_4__SCAN_IN), .A2(n21198), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n21194), .ZN(n21158) );
  OAI21_X1 U24084 ( .B1(n21160), .B2(n21182), .A(n21158), .ZN(P1_U3201) );
  AOI22_X1 U24085 ( .A1(P1_ADDRESS_REG_5__SCAN_IN), .A2(n21198), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n21193), .ZN(n21159) );
  OAI21_X1 U24086 ( .B1(n21160), .B2(n21179), .A(n21159), .ZN(P1_U3202) );
  AOI22_X1 U24087 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n21198), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n21194), .ZN(n21161) );
  OAI21_X1 U24088 ( .B1(n21162), .B2(n21182), .A(n21161), .ZN(P1_U3203) );
  AOI222_X1 U24089 ( .A1(n21193), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n21198), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n21194), .ZN(n21163) );
  INV_X1 U24090 ( .A(n21163), .ZN(P1_U3204) );
  AOI222_X1 U24091 ( .A1(n21194), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n21198), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n21193), .ZN(n21164) );
  INV_X1 U24092 ( .A(n21164), .ZN(P1_U3205) );
  AOI222_X1 U24093 ( .A1(n21193), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n21198), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n21194), .ZN(n21165) );
  INV_X1 U24094 ( .A(n21165), .ZN(P1_U3206) );
  AOI222_X1 U24095 ( .A1(n21194), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n21198), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n21193), .ZN(n21166) );
  INV_X1 U24096 ( .A(n21166), .ZN(P1_U3207) );
  AOI222_X1 U24097 ( .A1(n21194), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n21198), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n21193), .ZN(n21167) );
  INV_X1 U24098 ( .A(n21167), .ZN(P1_U3208) );
  AOI22_X1 U24099 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(n21198), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n21193), .ZN(n21168) );
  OAI21_X1 U24100 ( .B1(n21169), .B2(n21179), .A(n21168), .ZN(P1_U3209) );
  AOI22_X1 U24101 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n21198), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n21194), .ZN(n21170) );
  OAI21_X1 U24102 ( .B1(n21171), .B2(n21182), .A(n21170), .ZN(P1_U3210) );
  AOI222_X1 U24103 ( .A1(n21194), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n21198), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n21193), .ZN(n21172) );
  INV_X1 U24104 ( .A(n21172), .ZN(P1_U3211) );
  AOI22_X1 U24105 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n21198), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n21193), .ZN(n21173) );
  OAI21_X1 U24106 ( .B1(n21174), .B2(n21179), .A(n21173), .ZN(P1_U3212) );
  AOI22_X1 U24107 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n21198), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n21194), .ZN(n21175) );
  OAI21_X1 U24108 ( .B1(n21176), .B2(n21182), .A(n21175), .ZN(P1_U3213) );
  AOI222_X1 U24109 ( .A1(n21194), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n21198), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n21193), .ZN(n21177) );
  INV_X1 U24110 ( .A(n21177), .ZN(P1_U3214) );
  INV_X1 U24111 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n21180) );
  AOI22_X1 U24112 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n21198), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n21193), .ZN(n21178) );
  OAI21_X1 U24113 ( .B1(n21180), .B2(n21179), .A(n21178), .ZN(P1_U3215) );
  AOI22_X1 U24114 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(n21198), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n21194), .ZN(n21181) );
  OAI21_X1 U24115 ( .B1(n21183), .B2(n21182), .A(n21181), .ZN(P1_U3216) );
  AOI222_X1 U24116 ( .A1(n21194), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n21198), .C1(P1_REIP_REG_22__SCAN_IN), 
        .C2(n21193), .ZN(n21184) );
  INV_X1 U24117 ( .A(n21184), .ZN(P1_U3217) );
  AOI222_X1 U24118 ( .A1(n21194), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n21198), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n21193), .ZN(n21185) );
  INV_X1 U24119 ( .A(n21185), .ZN(P1_U3218) );
  AOI222_X1 U24120 ( .A1(n21194), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n21198), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n21193), .ZN(n21186) );
  INV_X1 U24121 ( .A(n21186), .ZN(P1_U3219) );
  AOI222_X1 U24122 ( .A1(n21194), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n21198), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n21193), .ZN(n21187) );
  INV_X1 U24123 ( .A(n21187), .ZN(P1_U3220) );
  AOI222_X1 U24124 ( .A1(n21194), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n21198), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n21193), .ZN(n21188) );
  INV_X1 U24125 ( .A(n21188), .ZN(P1_U3221) );
  AOI222_X1 U24126 ( .A1(n21194), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n21198), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n21193), .ZN(n21189) );
  INV_X1 U24127 ( .A(n21189), .ZN(P1_U3222) );
  AOI222_X1 U24128 ( .A1(n21194), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n21198), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n21193), .ZN(n21190) );
  INV_X1 U24129 ( .A(n21190), .ZN(P1_U3223) );
  AOI222_X1 U24130 ( .A1(n21194), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n21198), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n21193), .ZN(n21191) );
  INV_X1 U24131 ( .A(n21191), .ZN(P1_U3224) );
  AOI222_X1 U24132 ( .A1(n21193), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n21198), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n21194), .ZN(n21192) );
  INV_X1 U24133 ( .A(n21192), .ZN(P1_U3225) );
  AOI222_X1 U24134 ( .A1(n21194), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n21198), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n21193), .ZN(n21195) );
  INV_X1 U24135 ( .A(n21195), .ZN(P1_U3226) );
  OAI22_X1 U24136 ( .A1(n21198), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n21214), .ZN(n21196) );
  INV_X1 U24137 ( .A(n21196), .ZN(P1_U3458) );
  OAI22_X1 U24138 ( .A1(n21198), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n21214), .ZN(n21197) );
  INV_X1 U24139 ( .A(n21197), .ZN(P1_U3459) );
  OAI22_X1 U24140 ( .A1(n21198), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n21214), .ZN(n21199) );
  INV_X1 U24141 ( .A(n21199), .ZN(P1_U3460) );
  OAI22_X1 U24142 ( .A1(n21198), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n21214), .ZN(n21200) );
  INV_X1 U24143 ( .A(n21200), .ZN(P1_U3461) );
  OAI21_X1 U24144 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n21204), .A(n21202), 
        .ZN(n21201) );
  INV_X1 U24145 ( .A(n21201), .ZN(P1_U3464) );
  OAI21_X1 U24146 ( .B1(n21204), .B2(n21203), .A(n21202), .ZN(P1_U3465) );
  AOI21_X1 U24147 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n21205) );
  OAI22_X1 U24148 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(n21206), .B1(
        P1_REIP_REG_1__SCAN_IN), .B2(n21205), .ZN(n21208) );
  INV_X1 U24149 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21207) );
  AOI22_X1 U24150 ( .A1(n21212), .A2(n21208), .B1(n21207), .B2(n21209), .ZN(
        P1_U3481) );
  NOR2_X1 U24151 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .ZN(n21211) );
  INV_X1 U24152 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21210) );
  AOI22_X1 U24153 ( .A1(n21212), .A2(n21211), .B1(n21210), .B2(n21209), .ZN(
        P1_U3482) );
  AOI22_X1 U24154 ( .A1(n21214), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21213), 
        .B2(n21198), .ZN(P1_U3483) );
  OAI211_X1 U24155 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n21216), .A(n21215), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n21217) );
  OAI21_X1 U24156 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n21218), .A(n21217), 
        .ZN(n21224) );
  AOI211_X1 U24157 ( .C1(n20473), .C2(n21221), .A(n21220), .B(n21219), .ZN(
        n21223) );
  NAND2_X1 U24158 ( .A1(n21223), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n21222) );
  OAI21_X1 U24159 ( .B1(n21224), .B2(n21223), .A(n21222), .ZN(P1_U3485) );
  MUX2_X1 U24160 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(P1_M_IO_N_REG_SCAN_IN), 
        .S(n21198), .Z(P1_U3486) );
  INV_X1 U24161 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n21359) );
  NAND4_X1 U24162 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(P1_EAX_REG_22__SCAN_IN), 
        .A3(n21359), .A4(n21368), .ZN(n21229) );
  NAND4_X1 U24163 ( .A1(P2_EAX_REG_28__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_2__0__SCAN_IN), .A3(P1_UWORD_REG_4__SCAN_IN), .A4(
        n21365), .ZN(n21225) );
  NOR3_X1 U24164 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n21225), .A3(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n21226) );
  NAND3_X1 U24165 ( .A1(n21226), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A3(
        P2_EBX_REG_9__SCAN_IN), .ZN(n21228) );
  INV_X1 U24166 ( .A(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n21350) );
  NAND4_X1 U24167 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P1_LWORD_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_2__SCAN_IN), .A4(
        n21350), .ZN(n21227) );
  NOR3_X1 U24168 ( .A1(n21229), .A2(n21228), .A3(n21227), .ZN(n21381) );
  NAND4_X1 U24169 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_9__3__SCAN_IN), .A3(P3_EBX_REG_24__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n21244) );
  NOR4_X1 U24170 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        n21247), .ZN(n21232) );
  NOR4_X1 U24171 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n21253), .A3(
        n21252), .A4(n21250), .ZN(n21231) );
  INV_X1 U24172 ( .A(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n21272) );
  NOR3_X1 U24173 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A3(n21272), .ZN(n21230) );
  NAND4_X1 U24174 ( .A1(n21232), .A2(n21231), .A3(P1_DATAO_REG_31__SCAN_IN), 
        .A4(n21230), .ZN(n21243) );
  NOR4_X1 U24175 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_EBX_REG_15__SCAN_IN), .A3(n15014), .A4(n21279), .ZN(n21236) );
  INV_X1 U24176 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n21281) );
  NOR4_X1 U24177 ( .A1(P2_CODEFETCH_REG_SCAN_IN), .A2(n12545), .A3(n21281), 
        .A4(n21286), .ZN(n21235) );
  INV_X1 U24178 ( .A(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n21296) );
  NOR4_X1 U24179 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A3(n21296), .A4(n21285), .ZN(n21234) );
  NOR4_X1 U24180 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P1_DATAO_REG_12__SCAN_IN), .A3(P2_LWORD_REG_11__SCAN_IN), .A4(n21299), 
        .ZN(n21233) );
  NAND4_X1 U24181 ( .A1(n21236), .A2(n21235), .A3(n21234), .A4(n21233), .ZN(
        n21242) );
  INV_X1 U24182 ( .A(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n21332) );
  NOR4_X1 U24183 ( .A1(DATAI_30_), .A2(n21332), .A3(n14148), .A4(n21334), .ZN(
        n21240) );
  NOR4_X1 U24184 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(
        P2_UWORD_REG_1__SCAN_IN), .A3(P3_FLUSH_REG_SCAN_IN), .A4(
        P3_DATAO_REG_27__SCAN_IN), .ZN(n21239) );
  NOR4_X1 U24185 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_REIP_REG_3__SCAN_IN), .A3(P3_DATAO_REG_3__SCAN_IN), .A4(n21323), 
        .ZN(n21238) );
  NOR4_X1 U24186 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(P3_DATAO_REG_15__SCAN_IN), 
        .A3(n21320), .A4(n21312), .ZN(n21237) );
  NAND4_X1 U24187 ( .A1(n21240), .A2(n21239), .A3(n21238), .A4(n21237), .ZN(
        n21241) );
  NOR4_X1 U24188 ( .A1(n21244), .A2(n21243), .A3(n21242), .A4(n21241), .ZN(
        n21380) );
  INV_X1 U24189 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n21246) );
  AOI22_X1 U24190 ( .A1(n21247), .A2(keyinput43), .B1(n21246), .B2(keyinput3), 
        .ZN(n21245) );
  OAI221_X1 U24191 ( .B1(n21247), .B2(keyinput43), .C1(n21246), .C2(keyinput3), 
        .A(n21245), .ZN(n21260) );
  INV_X1 U24192 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n21249) );
  AOI22_X1 U24193 ( .A1(n21250), .A2(keyinput33), .B1(n21249), .B2(keyinput30), 
        .ZN(n21248) );
  OAI221_X1 U24194 ( .B1(n21250), .B2(keyinput33), .C1(n21249), .C2(keyinput30), .A(n21248), .ZN(n21259) );
  AOI22_X1 U24195 ( .A1(n21253), .A2(keyinput39), .B1(keyinput29), .B2(n21252), 
        .ZN(n21251) );
  OAI221_X1 U24196 ( .B1(n21253), .B2(keyinput39), .C1(n21252), .C2(keyinput29), .A(n21251), .ZN(n21258) );
  AOI22_X1 U24197 ( .A1(n21256), .A2(keyinput48), .B1(n21255), .B2(keyinput38), 
        .ZN(n21254) );
  OAI221_X1 U24198 ( .B1(n21256), .B2(keyinput48), .C1(n21255), .C2(keyinput38), .A(n21254), .ZN(n21257) );
  NOR4_X1 U24199 ( .A1(n21260), .A2(n21259), .A3(n21258), .A4(n21257), .ZN(
        n21310) );
  INV_X1 U24200 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n21263) );
  AOI22_X1 U24201 ( .A1(n21263), .A2(keyinput36), .B1(keyinput20), .B2(n21262), 
        .ZN(n21261) );
  OAI221_X1 U24202 ( .B1(n21263), .B2(keyinput36), .C1(n21262), .C2(keyinput20), .A(n21261), .ZN(n21276) );
  INV_X1 U24203 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n21265) );
  AOI22_X1 U24204 ( .A1(n21266), .A2(keyinput59), .B1(n21265), .B2(keyinput37), 
        .ZN(n21264) );
  OAI221_X1 U24205 ( .B1(n21266), .B2(keyinput59), .C1(n21265), .C2(keyinput37), .A(n21264), .ZN(n21275) );
  AOI22_X1 U24206 ( .A1(n21269), .A2(keyinput19), .B1(keyinput26), .B2(n21268), 
        .ZN(n21267) );
  OAI221_X1 U24207 ( .B1(n21269), .B2(keyinput19), .C1(n21268), .C2(keyinput26), .A(n21267), .ZN(n21274) );
  AOI22_X1 U24208 ( .A1(n21272), .A2(keyinput50), .B1(n21271), .B2(keyinput9), 
        .ZN(n21270) );
  OAI221_X1 U24209 ( .B1(n21272), .B2(keyinput50), .C1(n21271), .C2(keyinput9), 
        .A(n21270), .ZN(n21273) );
  NOR4_X1 U24210 ( .A1(n21276), .A2(n21275), .A3(n21274), .A4(n21273), .ZN(
        n21309) );
  AOI22_X1 U24211 ( .A1(n21279), .A2(keyinput60), .B1(keyinput0), .B2(n21278), 
        .ZN(n21277) );
  OAI221_X1 U24212 ( .B1(n21279), .B2(keyinput60), .C1(n21278), .C2(keyinput0), 
        .A(n21277), .ZN(n21290) );
  AOI22_X1 U24213 ( .A1(n15014), .A2(keyinput2), .B1(n21281), .B2(keyinput52), 
        .ZN(n21280) );
  OAI221_X1 U24214 ( .B1(n15014), .B2(keyinput2), .C1(n21281), .C2(keyinput52), 
        .A(n21280), .ZN(n21289) );
  AOI22_X1 U24215 ( .A1(n21283), .A2(keyinput42), .B1(n12545), .B2(keyinput53), 
        .ZN(n21282) );
  OAI221_X1 U24216 ( .B1(n21283), .B2(keyinput42), .C1(n12545), .C2(keyinput53), .A(n21282), .ZN(n21288) );
  AOI22_X1 U24217 ( .A1(n21286), .A2(keyinput46), .B1(keyinput35), .B2(n21285), 
        .ZN(n21284) );
  OAI221_X1 U24218 ( .B1(n21286), .B2(keyinput46), .C1(n21285), .C2(keyinput35), .A(n21284), .ZN(n21287) );
  NOR4_X1 U24219 ( .A1(n21290), .A2(n21289), .A3(n21288), .A4(n21287), .ZN(
        n21308) );
  AOI22_X1 U24220 ( .A1(n21293), .A2(keyinput34), .B1(keyinput24), .B2(n21292), 
        .ZN(n21291) );
  OAI221_X1 U24221 ( .B1(n21293), .B2(keyinput34), .C1(n21292), .C2(keyinput24), .A(n21291), .ZN(n21306) );
  AOI22_X1 U24222 ( .A1(n21296), .A2(keyinput28), .B1(keyinput56), .B2(n21295), 
        .ZN(n21294) );
  OAI221_X1 U24223 ( .B1(n21296), .B2(keyinput28), .C1(n21295), .C2(keyinput56), .A(n21294), .ZN(n21305) );
  AOI22_X1 U24224 ( .A1(n21299), .A2(keyinput62), .B1(keyinput47), .B2(n21298), 
        .ZN(n21297) );
  OAI221_X1 U24225 ( .B1(n21299), .B2(keyinput62), .C1(n21298), .C2(keyinput47), .A(n21297), .ZN(n21304) );
  INV_X1 U24226 ( .A(DATAI_30_), .ZN(n21301) );
  AOI22_X1 U24227 ( .A1(n21302), .A2(keyinput40), .B1(keyinput31), .B2(n21301), 
        .ZN(n21300) );
  OAI221_X1 U24228 ( .B1(n21302), .B2(keyinput40), .C1(n21301), .C2(keyinput31), .A(n21300), .ZN(n21303) );
  NOR4_X1 U24229 ( .A1(n21306), .A2(n21305), .A3(n21304), .A4(n21303), .ZN(
        n21307) );
  NAND4_X1 U24230 ( .A1(n21310), .A2(n21309), .A3(n21308), .A4(n21307), .ZN(
        n21379) );
  AOI22_X1 U24231 ( .A1(n21313), .A2(keyinput16), .B1(n21312), .B2(keyinput18), 
        .ZN(n21311) );
  OAI221_X1 U24232 ( .B1(n21313), .B2(keyinput16), .C1(n21312), .C2(keyinput18), .A(n21311), .ZN(n21317) );
  XOR2_X1 U24233 ( .A(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B(keyinput6), .Z(
        n21316) );
  XNOR2_X1 U24234 ( .A(n21314), .B(keyinput54), .ZN(n21315) );
  OR3_X1 U24235 ( .A1(n21317), .A2(n21316), .A3(n21315), .ZN(n21326) );
  AOI22_X1 U24236 ( .A1(n21320), .A2(keyinput5), .B1(keyinput13), .B2(n21319), 
        .ZN(n21318) );
  OAI221_X1 U24237 ( .B1(n21320), .B2(keyinput5), .C1(n21319), .C2(keyinput13), 
        .A(n21318), .ZN(n21325) );
  AOI22_X1 U24238 ( .A1(n21323), .A2(keyinput12), .B1(n21322), .B2(keyinput7), 
        .ZN(n21321) );
  OAI221_X1 U24239 ( .B1(n21323), .B2(keyinput12), .C1(n21322), .C2(keyinput7), 
        .A(n21321), .ZN(n21324) );
  NOR3_X1 U24240 ( .A1(n21326), .A2(n21325), .A3(n21324), .ZN(n21377) );
  INV_X1 U24241 ( .A(P3_DATAO_REG_27__SCAN_IN), .ZN(n21329) );
  AOI22_X1 U24242 ( .A1(n21329), .A2(keyinput17), .B1(keyinput21), .B2(n21328), 
        .ZN(n21327) );
  OAI221_X1 U24243 ( .B1(n21329), .B2(keyinput17), .C1(n21328), .C2(keyinput21), .A(n21327), .ZN(n21341) );
  AOI22_X1 U24244 ( .A1(n21332), .A2(keyinput44), .B1(keyinput58), .B2(n21331), 
        .ZN(n21330) );
  OAI221_X1 U24245 ( .B1(n21332), .B2(keyinput44), .C1(n21331), .C2(keyinput58), .A(n21330), .ZN(n21340) );
  AOI22_X1 U24246 ( .A1(n21334), .A2(keyinput57), .B1(n14148), .B2(keyinput27), 
        .ZN(n21333) );
  OAI221_X1 U24247 ( .B1(n21334), .B2(keyinput57), .C1(n14148), .C2(keyinput27), .A(n21333), .ZN(n21339) );
  XOR2_X1 U24248 ( .A(n21335), .B(keyinput49), .Z(n21337) );
  XNOR2_X1 U24249 ( .A(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B(keyinput25), .ZN(
        n21336) );
  NAND2_X1 U24250 ( .A1(n21337), .A2(n21336), .ZN(n21338) );
  NOR4_X1 U24251 ( .A1(n21341), .A2(n21340), .A3(n21339), .A4(n21338), .ZN(
        n21376) );
  INV_X1 U24252 ( .A(P1_UWORD_REG_4__SCAN_IN), .ZN(n21343) );
  AOI22_X1 U24253 ( .A1(n21344), .A2(keyinput41), .B1(keyinput8), .B2(n21343), 
        .ZN(n21342) );
  OAI221_X1 U24254 ( .B1(n21344), .B2(keyinput41), .C1(n21343), .C2(keyinput8), 
        .A(n21342), .ZN(n21357) );
  AOI22_X1 U24255 ( .A1(n21347), .A2(keyinput61), .B1(n21346), .B2(keyinput51), 
        .ZN(n21345) );
  OAI221_X1 U24256 ( .B1(n21347), .B2(keyinput61), .C1(n21346), .C2(keyinput51), .A(n21345), .ZN(n21356) );
  AOI22_X1 U24257 ( .A1(n21350), .A2(keyinput32), .B1(keyinput22), .B2(n21349), 
        .ZN(n21348) );
  OAI221_X1 U24258 ( .B1(n21350), .B2(keyinput32), .C1(n21349), .C2(keyinput22), .A(n21348), .ZN(n21355) );
  INV_X1 U24259 ( .A(P1_LWORD_REG_12__SCAN_IN), .ZN(n21353) );
  AOI22_X1 U24260 ( .A1(n21353), .A2(keyinput45), .B1(keyinput55), .B2(n21352), 
        .ZN(n21351) );
  OAI221_X1 U24261 ( .B1(n21353), .B2(keyinput45), .C1(n21352), .C2(keyinput55), .A(n21351), .ZN(n21354) );
  NOR4_X1 U24262 ( .A1(n21357), .A2(n21356), .A3(n21355), .A4(n21354), .ZN(
        n21375) );
  AOI22_X1 U24263 ( .A1(n21360), .A2(keyinput23), .B1(n21359), .B2(keyinput15), 
        .ZN(n21358) );
  OAI221_X1 U24264 ( .B1(n21360), .B2(keyinput23), .C1(n21359), .C2(keyinput15), .A(n21358), .ZN(n21373) );
  INV_X1 U24265 ( .A(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n21363) );
  INV_X1 U24266 ( .A(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n21362) );
  AOI22_X1 U24267 ( .A1(n21363), .A2(keyinput63), .B1(keyinput11), .B2(n21362), 
        .ZN(n21361) );
  OAI221_X1 U24268 ( .B1(n21363), .B2(keyinput63), .C1(n21362), .C2(keyinput11), .A(n21361), .ZN(n21372) );
  AOI22_X1 U24269 ( .A1(n21366), .A2(keyinput14), .B1(keyinput4), .B2(n21365), 
        .ZN(n21364) );
  OAI221_X1 U24270 ( .B1(n21366), .B2(keyinput14), .C1(n21365), .C2(keyinput4), 
        .A(n21364), .ZN(n21371) );
  AOI22_X1 U24271 ( .A1(n21369), .A2(keyinput1), .B1(keyinput10), .B2(n21368), 
        .ZN(n21367) );
  OAI221_X1 U24272 ( .B1(n21369), .B2(keyinput1), .C1(n21368), .C2(keyinput10), 
        .A(n21367), .ZN(n21370) );
  NOR4_X1 U24273 ( .A1(n21373), .A2(n21372), .A3(n21371), .A4(n21370), .ZN(
        n21374) );
  NAND4_X1 U24274 ( .A1(n21377), .A2(n21376), .A3(n21375), .A4(n21374), .ZN(
        n21378) );
  AOI211_X1 U24275 ( .C1(n21381), .C2(n21380), .A(n21379), .B(n21378), .ZN(
        n21392) );
  INV_X1 U24276 ( .A(n21382), .ZN(n21390) );
  AOI22_X1 U24277 ( .A1(n21386), .A2(n21385), .B1(n21384), .B2(n21383), .ZN(
        n21388) );
  NAND3_X1 U24278 ( .A1(n21390), .A2(n21388), .A3(n21387), .ZN(n21389) );
  OAI21_X1 U24279 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n21390), .A(
        n21389), .ZN(n21391) );
  XNOR2_X1 U24280 ( .A(n21392), .B(n21391), .ZN(P1_U3478) );
  INV_X1 U11034 ( .A(n17980), .ZN(n17948) );
  NAND2_X2 U15576 ( .A1(n12285), .A2(n12284), .ZN(n12407) );
  AND3_X1 U15603 ( .A1(n12319), .A2(n12318), .A3(n12411), .ZN(n12380) );
  AND2_X1 U15566 ( .A1(n13968), .A2(n12276), .ZN(n12585) );
  INV_X2 U11194 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10441) );
  CLKBUF_X1 U11041 ( .A(n16829), .Z(n9570) );
  CLKBUF_X2 U11043 ( .A(n12469), .Z(n13043) );
  CLKBUF_X1 U11045 ( .A(n10479), .Z(n10768) );
  CLKBUF_X1 U11055 ( .A(n12426), .Z(n12427) );
  CLKBUF_X1 U11087 ( .A(n12421), .Z(n20626) );
  NOR3_X1 U11096 ( .A1(n15342), .A2(n15335), .A3(n10381), .ZN(n15336) );
  CLKBUF_X1 U11103 ( .A(n14537), .Z(n15158) );
  CLKBUF_X1 U11111 ( .A(n17349), .Z(n17348) );
  OR2_X1 U11179 ( .A1(n20627), .A2(n12403), .ZN(n21393) );
  OR2_X1 U11377 ( .A1(n20627), .A2(n20626), .ZN(n21394) );
endmodule

