

module b21_C_SARLock_k_64_5 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, 
        ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, 
        ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, 
        ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, 
        U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, 
        P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, 
        P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, 
        P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, 
        P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, 
        P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, 
        P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, 
        P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, 
        P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, 
        P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, 
        P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, 
        P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, 
        P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, 
        P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, 
        P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, 
        P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, 
        P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, 
        P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, 
        P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, 
        P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, 
        P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, 
        P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, 
        P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, 
        P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, 
        P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, 
        P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, 
        P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, 
        P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, 
        P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, 
        P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, 
        P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, 
        P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, 
        P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, 
        P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, 
        P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, 
        P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, 
        P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, 
        P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167;

  AND2_X1 U4816 ( .A1(n6203), .A2(n6343), .ZN(n8953) );
  INV_X1 U4817 ( .A(n9425), .ZN(n8539) );
  INV_X1 U4819 ( .A(n4311), .ZN(n6738) );
  INV_X2 U4820 ( .A(n6727), .ZN(n8323) );
  CLKBUF_X2 U4821 ( .A(n6528), .Z(n6716) );
  BUF_X4 U4822 ( .A(n8327), .Z(n4311) );
  INV_X2 U4823 ( .A(n6175), .ZN(n5648) );
  INV_X1 U4824 ( .A(n5558), .ZN(n4613) );
  NAND2_X2 U4825 ( .A1(n4701), .A2(n6518), .ZN(n6528) );
  INV_X1 U4826 ( .A(n7015), .ZN(n4701) );
  OR2_X1 U4827 ( .A1(n8219), .A2(n8034), .ZN(n4700) );
  OAI21_X1 U4828 ( .B1(n9044), .B2(n4757), .A(n4322), .ZN(n8989) );
  INV_X1 U4829 ( .A(n6032), .ZN(n6057) );
  AND2_X1 U4830 ( .A1(n9109), .A2(n8713), .ZN(n6349) );
  AND2_X1 U4831 ( .A1(n7806), .A2(n9930), .ZN(n8650) );
  NAND2_X1 U4832 ( .A1(n5707), .A2(n6799), .ZN(n5685) );
  INV_X1 U4833 ( .A(n7640), .ZN(n10076) );
  CLKBUF_X2 U4835 ( .A(n5102), .Z(n5459) );
  NOR2_X1 U4836 ( .A1(n5022), .A2(n9708), .ZN(n5086) );
  INV_X1 U4837 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9695) );
  NAND2_X1 U4838 ( .A1(n5010), .A2(n5003), .ZN(n6948) );
  NAND2_X1 U4839 ( .A1(n5468), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5469) );
  NAND2_X1 U4840 ( .A1(n5975), .A2(n5974), .ZN(n9135) );
  NAND2_X1 U4841 ( .A1(n5997), .A2(n5996), .ZN(n9124) );
  OAI211_X2 U4842 ( .C1(n6809), .C2(n5685), .A(n5585), .B(n5584), .ZN(n7546)
         );
  AND4_X1 U4843 ( .A1(n5149), .A2(n5148), .A3(n5147), .A4(n5146), .ZN(n8431)
         );
  INV_X1 U4844 ( .A(n9437), .ZN(n9431) );
  NAND2_X1 U4845 ( .A1(n6094), .A2(n6093), .ZN(n9109) );
  NAND2_X1 U4846 ( .A1(n8558), .A2(n4701), .ZN(n8327) );
  BUF_X2 U4847 ( .A(n4886), .Z(n4310) );
  OAI21_X2 U4848 ( .B1(P2_ADDR_REG_19__SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        n4882), .ZN(n4886) );
  INV_X1 U4849 ( .A(n8858), .ZN(n7634) );
  BUF_X1 U4850 ( .A(n9251), .Z(n9320) );
  NAND2_X1 U4851 ( .A1(n6189), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5585) );
  NAND2_X1 U4852 ( .A1(n6516), .A2(n9930), .ZN(n8558) );
  OAI21_X2 U4853 ( .B1(n5220), .B2(n4809), .A(n4806), .ZN(n4941) );
  AOI21_X2 U4854 ( .B1(n9370), .B2(n9360), .A(n9359), .ZN(n9361) );
  INV_X1 U4855 ( .A(n7745), .ZN(n6200) );
  XNOR2_X2 U4856 ( .A(n5572), .B(n5571), .ZN(n7745) );
  NAND2_X2 U4857 ( .A1(n6014), .A2(n6013), .ZN(n9119) );
  NAND2_X1 U4858 ( .A1(n4439), .A2(n4436), .ZN(n4435) );
  OR2_X1 U4859 ( .A1(n6365), .A2(n4440), .ZN(n4439) );
  NAND2_X1 U4860 ( .A1(n4837), .A2(n4836), .ZN(n9594) );
  NAND2_X1 U4861 ( .A1(n4389), .A2(n5377), .ZN(n9460) );
  NAND2_X1 U4862 ( .A1(n6165), .A2(n6164), .ZN(n9097) );
  AND2_X1 U4863 ( .A1(n4370), .A2(n4841), .ZN(n4836) );
  INV_X1 U4864 ( .A(n6350), .ZN(n6357) );
  AND2_X1 U4865 ( .A1(n9101), .A2(n6154), .ZN(n6350) );
  NAND2_X1 U4866 ( .A1(n4546), .A2(n4544), .ZN(n9517) );
  NAND2_X1 U4867 ( .A1(n6162), .A2(n6161), .ZN(n6182) );
  NAND2_X1 U4868 ( .A1(n8211), .A2(n4870), .ZN(n9545) );
  NAND2_X1 U4869 ( .A1(n4800), .A2(n4798), .ZN(n6162) );
  NAND2_X1 U4870 ( .A1(n5389), .A2(n5388), .ZN(n9612) );
  NAND2_X1 U4871 ( .A1(n6031), .A2(n6030), .ZN(n9113) );
  XNOR2_X1 U4872 ( .A(n5431), .B(n5430), .ZN(n8320) );
  NAND2_X1 U4873 ( .A1(n5986), .A2(n5985), .ZN(n9127) );
  NAND2_X1 U4874 ( .A1(n4740), .A2(n4337), .ZN(n8285) );
  AOI21_X1 U4875 ( .B1(n4833), .B2(n9573), .A(n4831), .ZN(n4830) );
  NAND2_X1 U4876 ( .A1(n5959), .A2(n5958), .ZN(n9141) );
  OR2_X1 U4877 ( .A1(n9746), .A2(n9749), .ZN(n9744) );
  AND2_X1 U4878 ( .A1(n6578), .A2(n6577), .ZN(n6579) );
  NAND2_X1 U4879 ( .A1(n5044), .A2(n5043), .ZN(n9644) );
  NAND2_X1 U4880 ( .A1(n5318), .A2(n5317), .ZN(n9647) );
  NAND2_X1 U4881 ( .A1(n5306), .A2(n5305), .ZN(n9654) );
  NAND2_X1 U4882 ( .A1(n7483), .A2(n5187), .ZN(n7582) );
  OAI211_X1 U4883 ( .C1(n7003), .C2(n4675), .A(n4674), .B(n9225), .ZN(n9227)
         );
  NAND2_X1 U4884 ( .A1(n5223), .A2(n5222), .ZN(n6600) );
  NAND2_X1 U4885 ( .A1(n5733), .A2(n5732), .ZN(n7957) );
  AND2_X1 U4886 ( .A1(n8422), .A2(n8429), .ZN(n8569) );
  AND2_X1 U4887 ( .A1(n6925), .A2(n6924), .ZN(n9876) );
  INV_X1 U4888 ( .A(n8434), .ZN(n9967) );
  NOR2_X1 U4889 ( .A1(n6749), .A2(n6758), .ZN(n9322) );
  AND2_X1 U4890 ( .A1(n7019), .A2(n5098), .ZN(n7131) );
  NAND2_X1 U4891 ( .A1(n4572), .A2(n4571), .ZN(n9925) );
  NAND2_X1 U4892 ( .A1(n7344), .A2(n8372), .ZN(n8564) );
  INV_X1 U4893 ( .A(n8556), .ZN(n8536) );
  NAND2_X1 U4894 ( .A1(n6236), .A2(n7667), .ZN(n8700) );
  NAND2_X1 U4895 ( .A1(n8377), .A2(n8378), .ZN(n8565) );
  INV_X1 U4896 ( .A(n7287), .ZN(n9355) );
  INV_X1 U4897 ( .A(n7438), .ZN(n9354) );
  INV_X1 U4898 ( .A(n8859), .ZN(n7555) );
  INV_X2 U4899 ( .A(n6544), .ZN(n6727) );
  INV_X1 U4900 ( .A(n6544), .ZN(n4312) );
  INV_X1 U4901 ( .A(n7546), .ZN(n10052) );
  XNOR2_X2 U4902 ( .A(n6529), .B(n4393), .ZN(n7018) );
  NAND2_X1 U4903 ( .A1(n5115), .A2(n4541), .ZN(n9230) );
  AND4_X1 U4904 ( .A1(n5162), .A2(n5161), .A3(n5160), .A4(n5159), .ZN(n8438)
         );
  INV_X1 U4905 ( .A(n7202), .ZN(n9357) );
  AND4_X1 U4906 ( .A1(n5121), .A2(n5120), .A3(n5119), .A4(n5118), .ZN(n7287)
         );
  NAND2_X1 U4907 ( .A1(n4819), .A2(n4903), .ZN(n5138) );
  AND2_X2 U4908 ( .A1(n7015), .A2(n6518), .ZN(n6544) );
  INV_X1 U4909 ( .A(n6518), .ZN(n6765) );
  NAND4_X1 U4910 ( .A1(n5091), .A2(n5090), .A3(n5089), .A4(n5088), .ZN(n6526)
         );
  AND4_X1 U4911 ( .A1(n5061), .A2(n5060), .A3(n5059), .A4(n5058), .ZN(n7202)
         );
  OAI211_X1 U4912 ( .C1(n5165), .C2(n6811), .A(n5070), .B(n5069), .ZN(n7010)
         );
  NAND2_X1 U4913 ( .A1(n4820), .A2(n4900), .ZN(n5122) );
  INV_X4 U4914 ( .A(n5140), .ZN(n6769) );
  INV_X1 U4915 ( .A(n5114), .ZN(n5165) );
  INV_X2 U4916 ( .A(n5685), .ZN(n6188) );
  BUF_X2 U4917 ( .A(n5622), .Z(n6166) );
  NAND2_X1 U4918 ( .A1(n5557), .A2(n5558), .ZN(n6175) );
  INV_X1 U4919 ( .A(n5707), .ZN(n5863) );
  XNOR2_X1 U4920 ( .A(n5474), .B(n5473), .ZN(n8242) );
  AND2_X1 U4921 ( .A1(n5022), .A2(n5020), .ZN(n5102) );
  NAND2_X1 U4922 ( .A1(n5466), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5470) );
  CLKBUF_X3 U4923 ( .A(n5087), .Z(n6817) );
  XNOR2_X1 U4924 ( .A(n5042), .B(n5041), .ZN(n9930) );
  AND2_X1 U4925 ( .A1(n5022), .A2(n9708), .ZN(n5087) );
  NAND2_X1 U4926 ( .A1(n5482), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5474) );
  NAND2_X1 U4927 ( .A1(n5017), .A2(n5018), .ZN(n9708) );
  XNOR2_X1 U4928 ( .A(n5478), .B(n5477), .ZN(n8034) );
  NAND2_X1 U4929 ( .A1(n5579), .A2(n5578), .ZN(n8663) );
  NAND2_X1 U4930 ( .A1(n5476), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5478) );
  NAND2_X1 U4931 ( .A1(n5583), .A2(n5582), .ZN(n8687) );
  MUX2_X1 U4932 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5014), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5017) );
  XNOR2_X1 U4933 ( .A(n5019), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5022) );
  MUX2_X1 U4934 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5009), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n5010) );
  NAND2_X1 U4935 ( .A1(n5018), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5019) );
  AND2_X1 U4936 ( .A1(n5047), .A2(n5037), .ZN(n5280) );
  NAND2_X2 U4937 ( .A1(n6799), .A2(P1_U3084), .ZN(n9704) );
  AND3_X1 U4939 ( .A1(n4990), .A2(n4989), .A3(n4988), .ZN(n4997) );
  NAND2_X2 U4940 ( .A1(n4884), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4885) );
  NAND2_X1 U4941 ( .A1(n4883), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4884) );
  AND2_X1 U4942 ( .A1(n5110), .A2(n4999), .ZN(n4873) );
  AND4_X1 U4943 ( .A1(n4994), .A2(n4993), .A3(n4992), .A4(n4991), .ZN(n4996)
         );
  INV_X1 U4944 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5238) );
  NOR2_X1 U4945 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n4991) );
  NOR2_X1 U4946 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n4992) );
  NOR2_X1 U4947 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5034) );
  NOR2_X1 U4948 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n4993) );
  NOR2_X1 U4949 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n4988) );
  INV_X1 U4950 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5110) );
  INV_X4 U4951 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U4952 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5821) );
  INV_X4 U4953 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U4954 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4882) );
  INV_X1 U4955 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4883) );
  INV_X1 U4956 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5687) );
  AND2_X1 U4957 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5129) );
  NOR2_X2 U4958 ( .A1(n8232), .A2(n9172), .ZN(n8282) );
  OAI21_X1 U4959 ( .B1(n9445), .B2(n8593), .A(n4847), .ZN(n9432) );
  NOR2_X2 U4960 ( .A1(n9113), .A2(n8956), .ZN(n6342) );
  NOR2_X2 U4961 ( .A1(n9564), .A2(n9654), .ZN(n9563) );
  XNOR2_X2 U4962 ( .A(n6049), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8941) );
  NAND2_X2 U4963 ( .A1(n6015), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6049) );
  AOI21_X1 U4964 ( .B1(n4802), .B2(n4804), .A(n4799), .ZN(n4798) );
  INV_X1 U4965 ( .A(n6157), .ZN(n4799) );
  AND2_X1 U4966 ( .A1(n5558), .A2(n5559), .ZN(n5622) );
  INV_X1 U4967 ( .A(n4644), .ZN(n4642) );
  NAND2_X1 U4968 ( .A1(n9038), .A2(n8673), .ZN(n4648) );
  NOR2_X1 U4969 ( .A1(n6677), .A2(n9306), .ZN(n4689) );
  NAND2_X1 U4970 ( .A1(n4851), .A2(n4850), .ZN(n9487) );
  AOI21_X1 U4971 ( .B1(n4852), .B2(n4858), .A(n4350), .ZN(n4850) );
  NAND2_X1 U4972 ( .A1(n5339), .A2(n4852), .ZN(n4851) );
  OAI21_X1 U4973 ( .B1(n6296), .B2(n4878), .A(n6295), .ZN(n6311) );
  OR2_X1 U4974 ( .A1(n7756), .A2(n7555), .ZN(n6245) );
  NAND2_X1 U4975 ( .A1(n4932), .A2(n6424), .ZN(n4935) );
  INV_X1 U4976 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n4918) );
  NAND2_X1 U4977 ( .A1(n4914), .A2(n4913), .ZN(n4917) );
  INV_X1 U4978 ( .A(n6349), .ZN(n6152) );
  NOR2_X1 U4979 ( .A1(n8083), .A2(n4460), .ZN(n4459) );
  INV_X1 U4980 ( .A(n4461), .ZN(n4460) );
  AND2_X1 U4981 ( .A1(n7722), .A2(n7721), .ZN(n7854) );
  NAND2_X1 U4982 ( .A1(n5707), .A2(n5400), .ZN(n5684) );
  NAND2_X1 U4983 ( .A1(n6200), .A2(n6226), .ZN(n7331) );
  OR2_X1 U4984 ( .A1(n8083), .A2(n8852), .ZN(n4637) );
  NOR2_X1 U4985 ( .A1(n7991), .A2(n4635), .ZN(n4634) );
  INV_X1 U4986 ( .A(n4637), .ZN(n4635) );
  NAND2_X1 U4987 ( .A1(n9261), .A2(n6669), .ZN(n6675) );
  OR2_X1 U4988 ( .A1(n9583), .A2(n8410), .ZN(n8639) );
  OR2_X1 U4989 ( .A1(n9596), .A2(n9438), .ZN(n8541) );
  NAND2_X1 U4990 ( .A1(n9436), .A2(n9450), .ZN(n4846) );
  OR2_X1 U4991 ( .A1(n9634), .A2(n9538), .ZN(n8511) );
  OAI211_X1 U4992 ( .C1(n4830), .C2(n4543), .A(n8502), .B(n4542), .ZN(n4552)
         );
  INV_X1 U4993 ( .A(n9547), .ZN(n4543) );
  NAND2_X1 U4994 ( .A1(n4833), .A2(n9547), .ZN(n4542) );
  NAND2_X1 U4995 ( .A1(n4830), .A2(n8502), .ZN(n4553) );
  NOR2_X1 U4996 ( .A1(n9637), .A2(n4527), .ZN(n4526) );
  INV_X1 U4997 ( .A(n4528), .ZN(n4527) );
  NOR2_X1 U4998 ( .A1(n6187), .A2(SI_30_), .ZN(n4770) );
  OR2_X1 U4999 ( .A1(n4774), .A2(n6163), .ZN(n4767) );
  NAND2_X1 U5000 ( .A1(n6182), .A2(n6187), .ZN(n4774) );
  NAND2_X1 U5001 ( .A1(n5433), .A2(n5432), .ZN(n5447) );
  AOI21_X1 U5002 ( .B1(n4783), .B2(n4781), .A(n4780), .ZN(n4779) );
  INV_X1 U5003 ( .A(n5413), .ZN(n4780) );
  INV_X1 U5004 ( .A(n4785), .ZN(n4781) );
  NAND2_X1 U5005 ( .A1(n5369), .A2(n5368), .ZN(n5383) );
  AND2_X1 U5006 ( .A1(n4956), .A2(n4955), .ZN(n5268) );
  NAND2_X1 U5007 ( .A1(n4515), .A2(n4944), .ZN(n5279) );
  NAND2_X1 U5008 ( .A1(n4941), .A2(n4520), .ZN(n4515) );
  NAND2_X1 U5009 ( .A1(n4928), .A2(n4927), .ZN(n5220) );
  NAND2_X1 U5010 ( .A1(n5164), .A2(n4909), .ZN(n4816) );
  INV_X1 U5011 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4998) );
  INV_X1 U5012 ( .A(n10046), .ZN(n6374) );
  OR2_X1 U5013 ( .A1(n7045), .A2(n7044), .ZN(n4481) );
  NAND2_X1 U5014 ( .A1(n4663), .A2(n4668), .ZN(n4662) );
  INV_X1 U5015 ( .A(n4666), .ZN(n4663) );
  AOI21_X1 U5016 ( .B1(n8953), .B2(n4669), .A(n4667), .ZN(n4666) );
  INV_X1 U5017 ( .A(n8988), .ZN(n8954) );
  OR2_X1 U5018 ( .A1(n9127), .A2(n8843), .ZN(n8675) );
  NAND2_X1 U5019 ( .A1(n4356), .A2(n4648), .ZN(n4644) );
  OR2_X1 U5020 ( .A1(n9155), .A2(n9071), .ZN(n8671) );
  NAND2_X1 U5021 ( .A1(n7981), .A2(n6133), .ZN(n4739) );
  OR2_X1 U5022 ( .A1(n10087), .A2(n6226), .ZN(n7538) );
  NAND2_X1 U5023 ( .A1(n5550), .A2(n4766), .ZN(n4765) );
  INV_X1 U5024 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5550) );
  NAND2_X1 U5025 ( .A1(n5553), .A2(n5556), .ZN(n5558) );
  MUX2_X1 U5026 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5555), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n5556) );
  OR2_X1 U5027 ( .A1(n4725), .A2(n9315), .ZN(n4721) );
  NAND2_X1 U5028 ( .A1(n5456), .A2(n5455), .ZN(n9591) );
  AND2_X1 U5029 ( .A1(n5425), .A2(n5458), .ZN(n9434) );
  OR2_X1 U5030 ( .A1(n9624), .A2(n9505), .ZN(n8412) );
  AND2_X1 U5031 ( .A1(n9624), .A2(n9339), .ZN(n5364) );
  AOI21_X1 U5032 ( .B1(n4857), .B2(n4855), .A(n4345), .ZN(n4854) );
  INV_X1 U5033 ( .A(n4872), .ZN(n4855) );
  OR2_X1 U5034 ( .A1(n9637), .A2(n9549), .ZN(n9518) );
  NOR2_X1 U5035 ( .A1(n9637), .A2(n9342), .ZN(n5338) );
  AND2_X1 U5036 ( .A1(n9644), .A2(n9343), .ZN(n5324) );
  NAND2_X1 U5037 ( .A1(n9558), .A2(n9537), .ZN(n4390) );
  AND2_X1 U5038 ( .A1(n4867), .A2(n4866), .ZN(n4865) );
  AND2_X1 U5039 ( .A1(n5485), .A2(n5001), .ZN(n4866) );
  INV_X1 U5040 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5001) );
  NOR4_X1 U5041 ( .A1(n6240), .A2(n6234), .A3(n6233), .A4(n6254), .ZN(n6243)
         );
  NAND2_X1 U5042 ( .A1(n4495), .A2(n4492), .ZN(n6329) );
  NAND2_X1 U5043 ( .A1(n4493), .A2(n4453), .ZN(n4492) );
  OAI21_X1 U5044 ( .B1(n4447), .B2(n4445), .A(n4443), .ZN(n4442) );
  OR2_X1 U5045 ( .A1(n6338), .A2(n4446), .ZN(n4445) );
  AOI21_X1 U5046 ( .B1(n6319), .B2(n4448), .A(n4346), .ZN(n4447) );
  NOR2_X1 U5047 ( .A1(n6336), .A2(n4444), .ZN(n4443) );
  INV_X1 U5048 ( .A(n4803), .ZN(n4802) );
  OAI21_X1 U5049 ( .B1(n5446), .B2(n4804), .A(n6155), .ZN(n4803) );
  OR2_X1 U5050 ( .A1(n6193), .A2(n6192), .ZN(n6368) );
  OR2_X1 U5051 ( .A1(n9097), .A2(n8685), .ZN(n6363) );
  AND3_X1 U5052 ( .A1(n5687), .A2(n5749), .A3(n5821), .ZN(n5545) );
  NOR2_X1 U5053 ( .A1(n4686), .A2(n4682), .ZN(n4681) );
  INV_X1 U5054 ( .A(n9281), .ZN(n4682) );
  INV_X1 U5055 ( .A(n9244), .ZN(n4686) );
  NAND2_X1 U5056 ( .A1(n9244), .A2(n4685), .ZN(n4684) );
  INV_X1 U5057 ( .A(n6697), .ZN(n4685) );
  OAI21_X1 U5058 ( .B1(n4400), .B2(n4319), .A(n4398), .ZN(n4397) );
  AOI21_X1 U5059 ( .B1(n8524), .B2(n8528), .A(n9607), .ZN(n4400) );
  OAI21_X1 U5060 ( .B1(n8524), .B2(n9337), .A(n4399), .ZN(n4398) );
  INV_X1 U5061 ( .A(n4793), .ZN(n4792) );
  INV_X1 U5062 ( .A(n5268), .ZN(n4797) );
  NAND2_X1 U5063 ( .A1(n4924), .A2(n6484), .ZN(n4927) );
  NAND2_X1 U5064 ( .A1(n4583), .A2(n4586), .ZN(n4582) );
  OR2_X1 U5065 ( .A1(n8775), .A2(n8774), .ZN(n4609) );
  NAND2_X1 U5066 ( .A1(n4441), .A2(n4453), .ZN(n4440) );
  INV_X1 U5067 ( .A(n6364), .ZN(n4441) );
  NAND2_X1 U5068 ( .A1(n6371), .A2(n6370), .ZN(n4438) );
  OAI21_X1 U5069 ( .B1(n6219), .B2(n10027), .A(n7820), .ZN(n6218) );
  AND2_X1 U5070 ( .A1(n5747), .A2(n5746), .ZN(n5786) );
  INV_X1 U5071 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5547) );
  NAND4_X1 U5072 ( .A1(n5545), .A2(n5544), .A3(n5543), .A4(n5542), .ZN(n5546)
         );
  NOR2_X1 U5073 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5544) );
  NOR2_X1 U5074 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5543) );
  NOR2_X1 U5075 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5542) );
  NAND2_X1 U5076 ( .A1(n4484), .A2(n4483), .ZN(n4482) );
  NAND2_X1 U5077 ( .A1(n8885), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4483) );
  NAND2_X1 U5078 ( .A1(n8682), .A2(n4474), .ZN(n4473) );
  NAND2_X1 U5079 ( .A1(n8943), .A2(n8956), .ZN(n4668) );
  INV_X1 U5080 ( .A(n6146), .ZN(n4755) );
  AND2_X1 U5081 ( .A1(n9135), .A2(n8778), .ZN(n6323) );
  INV_X1 U5082 ( .A(n6323), .ZN(n8991) );
  AND2_X1 U5083 ( .A1(n6142), .A2(n4748), .ZN(n4747) );
  NAND2_X1 U5084 ( .A1(n9082), .A2(n4749), .ZN(n4748) );
  INV_X1 U5085 ( .A(n9082), .ZN(n4750) );
  OR2_X1 U5086 ( .A1(n9149), .A2(n9050), .ZN(n6318) );
  NOR2_X1 U5087 ( .A1(n9161), .A2(n9167), .ZN(n4469) );
  INV_X1 U5088 ( .A(n4628), .ZN(n4622) );
  OR2_X1 U5089 ( .A1(n8264), .A2(n8155), .ZN(n6289) );
  AND2_X1 U5090 ( .A1(n8040), .A2(n8075), .ZN(n6270) );
  NOR2_X1 U5091 ( .A1(n8040), .A2(n7986), .ZN(n4461) );
  NOR2_X1 U5092 ( .A1(n7631), .A2(n6125), .ZN(n4743) );
  OR2_X1 U5093 ( .A1(n10022), .A2(n7634), .ZN(n6249) );
  OR2_X1 U5094 ( .A1(n8068), .A2(n8074), .ZN(n4636) );
  INV_X1 U5095 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5749) );
  AND2_X1 U5096 ( .A1(n4432), .A2(n4431), .ZN(n4731) );
  INV_X1 U5097 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4432) );
  INV_X1 U5098 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n4431) );
  NOR2_X1 U5099 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4730) );
  MUX2_X1 U5100 ( .A(n8545), .B(n8556), .S(n9591), .Z(n8549) );
  NAND2_X1 U5101 ( .A1(n9372), .A2(n9373), .ZN(n9375) );
  NOR2_X1 U5102 ( .A1(n8539), .A2(n4828), .ZN(n4827) );
  INV_X1 U5103 ( .A(n8541), .ZN(n4828) );
  NAND2_X1 U5104 ( .A1(n5519), .A2(n8541), .ZN(n4826) );
  OR2_X1 U5105 ( .A1(n9591), .A2(n9418), .ZN(n8405) );
  OR2_X1 U5106 ( .A1(n9601), .A2(n9450), .ZN(n8626) );
  INV_X1 U5107 ( .A(n8413), .ZN(n4560) );
  NOR2_X1 U5108 ( .A1(n9475), .A2(n4563), .ZN(n4562) );
  INV_X1 U5109 ( .A(n8412), .ZN(n4563) );
  AND2_X1 U5110 ( .A1(n4854), .A2(n4365), .ZN(n4852) );
  NAND2_X1 U5111 ( .A1(n4549), .A2(n4551), .ZN(n4545) );
  AOI21_X1 U5112 ( .B1(n4552), .B2(n4553), .A(n4550), .ZN(n4549) );
  INV_X1 U5113 ( .A(n5296), .ZN(n4861) );
  AND2_X1 U5114 ( .A1(n8481), .A2(n8480), .ZN(n8585) );
  NAND2_X1 U5115 ( .A1(n7969), .A2(n4568), .ZN(n4567) );
  NOR2_X1 U5116 ( .A1(n8115), .A2(n4569), .ZN(n4568) );
  INV_X1 U5117 ( .A(n8472), .ZN(n4569) );
  OR2_X1 U5118 ( .A1(n9761), .A2(n7772), .ZN(n8487) );
  OR2_X1 U5119 ( .A1(n7707), .A2(n7736), .ZN(n8466) );
  OR2_X1 U5120 ( .A1(n7498), .A2(n7589), .ZN(n8451) );
  AND2_X1 U5121 ( .A1(n8372), .A2(n8377), .ZN(n4401) );
  NAND2_X1 U5122 ( .A1(n9357), .A2(n7368), .ZN(n8378) );
  OR2_X1 U5123 ( .A1(n5350), .A2(n5100), .ZN(n5107) );
  NAND2_X1 U5124 ( .A1(n4554), .A2(n4555), .ZN(n9416) );
  AOI21_X1 U5125 ( .B1(n9448), .B2(n4558), .A(n4556), .ZN(n4555) );
  NAND2_X1 U5126 ( .A1(n9447), .A2(n4558), .ZN(n4554) );
  INV_X1 U5127 ( .A(n8626), .ZN(n4556) );
  NOR2_X1 U5128 ( .A1(n4324), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n4867) );
  OAI22_X1 U5129 ( .A1(n4773), .A2(n4380), .B1(n6182), .B2(n4772), .ZN(n4771)
         );
  INV_X1 U5130 ( .A(n6187), .ZN(n4772) );
  INV_X1 U5131 ( .A(n6182), .ZN(n4773) );
  NAND2_X1 U5132 ( .A1(n6160), .A2(n6159), .ZN(n6163) );
  INV_X1 U5133 ( .A(n4783), .ZN(n4782) );
  AND2_X1 U5134 ( .A1(n5415), .A2(n5404), .ZN(n5413) );
  NOR2_X1 U5135 ( .A1(n5398), .A2(n4786), .ZN(n4785) );
  INV_X1 U5136 ( .A(n5381), .ZN(n4786) );
  AOI21_X1 U5137 ( .B1(n4785), .B2(n5382), .A(n4784), .ZN(n4783) );
  INV_X1 U5138 ( .A(n5397), .ZN(n4784) );
  INV_X1 U5139 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5485) );
  AND2_X1 U5140 ( .A1(n5368), .A2(n4987), .ZN(n5366) );
  INV_X1 U5141 ( .A(n5340), .ZN(n4815) );
  NAND2_X1 U5142 ( .A1(n4937), .A2(n4936), .ZN(n4940) );
  INV_X1 U5143 ( .A(SI_13_), .ZN(n4936) );
  INV_X1 U5144 ( .A(n4931), .ZN(n4812) );
  NOR2_X1 U5145 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5203) );
  INV_X1 U5146 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5166) );
  OAI21_X1 U5147 ( .B1(n4503), .B2(n4508), .A(n4504), .ZN(n5202) );
  AOI21_X1 U5148 ( .B1(n4507), .B2(n4509), .A(n4505), .ZN(n4504) );
  INV_X1 U5149 ( .A(n4923), .ZN(n4505) );
  OAI211_X1 U5150 ( .C1(n4310), .C2(P1_DATAO_REG_5__SCAN_IN), .A(n4524), .B(
        n4523), .ZN(n4904) );
  NAND2_X1 U5151 ( .A1(n4672), .A2(n6797), .ZN(n4524) );
  NOR2_X2 U5152 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5064) );
  INV_X1 U5153 ( .A(n6115), .ZN(n7226) );
  XNOR2_X1 U5154 ( .A(n7546), .B(n6032), .ZN(n5589) );
  NAND2_X1 U5155 ( .A1(n9181), .A2(n10027), .ZN(n6196) );
  NAND2_X1 U5156 ( .A1(n8775), .A2(n8774), .ZN(n4608) );
  NAND2_X1 U5157 ( .A1(n8773), .A2(n4609), .ZN(n4607) );
  INV_X1 U5158 ( .A(n5843), .ZN(n4597) );
  INV_X1 U5159 ( .A(n8258), .ZN(n4600) );
  OR2_X1 U5160 ( .A1(n6173), .A2(n10110), .ZN(n5604) );
  INV_X1 U5161 ( .A(n5622), .ZN(n5956) );
  AND3_X1 U5162 ( .A1(n5594), .A2(n5593), .A3(n4614), .ZN(n7548) );
  OAI21_X1 U5163 ( .B1(n4323), .B2(n4612), .A(n4613), .ZN(n4614) );
  NOR2_X1 U5164 ( .A1(n7120), .A2(n4372), .ZN(n7123) );
  OR2_X1 U5165 ( .A1(n7123), .A2(n7122), .ZN(n4487) );
  OR2_X1 U5166 ( .A1(n8270), .A2(n8269), .ZN(n4484) );
  XNOR2_X1 U5167 ( .A(n4482), .B(n8900), .ZN(n8886) );
  INV_X1 U5168 ( .A(n6342), .ZN(n8926) );
  AND2_X1 U5169 ( .A1(n4669), .A2(n4668), .ZN(n4664) );
  NAND2_X1 U5170 ( .A1(n8952), .A2(n6203), .ZN(n4761) );
  NAND2_X1 U5171 ( .A1(n4761), .A2(n4759), .ZN(n4881) );
  OR2_X1 U5172 ( .A1(n9119), .A2(n8842), .ZN(n4669) );
  OR2_X1 U5173 ( .A1(n9127), .A2(n9003), .ZN(n8964) );
  AOI21_X1 U5174 ( .B1(n4315), .B2(n4641), .A(n4352), .ZN(n4640) );
  INV_X1 U5175 ( .A(n4645), .ZN(n4641) );
  NAND2_X1 U5176 ( .A1(n6146), .A2(n9044), .ZN(n9020) );
  AND2_X1 U5177 ( .A1(n4648), .A2(n9056), .ZN(n4645) );
  AOI21_X1 U5178 ( .B1(n8670), .B2(n8669), .A(n8668), .ZN(n9076) );
  NOR2_X1 U5179 ( .A1(n9161), .A2(n8846), .ZN(n8668) );
  AND2_X1 U5180 ( .A1(n8288), .A2(n8223), .ZN(n4628) );
  NOR2_X1 U5181 ( .A1(n4625), .A2(n4627), .ZN(n4624) );
  INV_X1 U5182 ( .A(n8290), .ZN(n4625) );
  NAND2_X1 U5183 ( .A1(n4632), .A2(n4630), .ZN(n8159) );
  NOR2_X1 U5184 ( .A1(n4631), .A2(n6135), .ZN(n4630) );
  NAND2_X1 U5185 ( .A1(n4739), .A2(n4344), .ZN(n8057) );
  AOI21_X1 U5186 ( .B1(n4634), .B2(n8074), .A(n4347), .ZN(n4633) );
  AND2_X1 U5187 ( .A1(n6131), .A2(n6134), .ZN(n7991) );
  NAND2_X1 U5188 ( .A1(n5790), .A2(n5789), .ZN(n8083) );
  AND2_X1 U5189 ( .A1(n7982), .A2(n6281), .ZN(n8074) );
  NAND2_X1 U5190 ( .A1(n7858), .A2(n4618), .ZN(n4617) );
  NAND2_X1 U5191 ( .A1(n7854), .A2(n4619), .ZN(n4618) );
  OR2_X1 U5194 ( .A1(n7725), .A2(n7851), .ZN(n7866) );
  OAI211_X1 U5195 ( .C1(n6803), .C2(n5685), .A(n5641), .B(n5640), .ZN(n7756)
         );
  INV_X1 U5196 ( .A(n9053), .ZN(n9068) );
  INV_X1 U5197 ( .A(n9084), .ZN(n9049) );
  INV_X1 U5198 ( .A(n9070), .ZN(n9051) );
  NAND2_X1 U5199 ( .A1(n5949), .A2(n5948), .ZN(n9146) );
  AND2_X1 U5200 ( .A1(n8225), .A2(n10087), .ZN(n9170) );
  INV_X1 U5201 ( .A(n10022), .ZN(n7562) );
  OR2_X1 U5202 ( .A1(n6374), .A2(n6108), .ZN(n10095) );
  AND2_X1 U5203 ( .A1(n6073), .A2(n6072), .ZN(n10034) );
  NAND2_X1 U5204 ( .A1(n7038), .A2(n10045), .ZN(n10035) );
  XNOR2_X1 U5205 ( .A(n5552), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5559) );
  NAND2_X1 U5206 ( .A1(n5553), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5552) );
  OAI21_X1 U5207 ( .B1(n5581), .B2(n5554), .A(P2_IR_REG_28__SCAN_IN), .ZN(
        n4477) );
  NAND2_X1 U5208 ( .A1(n4611), .A2(n4476), .ZN(n4610) );
  INV_X1 U5209 ( .A(n4765), .ZN(n4611) );
  NOR2_X1 U5210 ( .A1(n6061), .A2(n4765), .ZN(n5581) );
  OR2_X1 U5211 ( .A1(n5567), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n6068) );
  XNOR2_X1 U5212 ( .A(n5568), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6226) );
  AND2_X1 U5213 ( .A1(n5826), .A2(n5861), .ZN(n7940) );
  AND2_X1 U5214 ( .A1(n5674), .A2(n5658), .ZN(n7091) );
  XNOR2_X1 U5215 ( .A(n4479), .B(P2_IR_REG_1__SCAN_IN), .ZN(n7033) );
  NAND2_X1 U5216 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4479) );
  INV_X1 U5217 ( .A(n6564), .ZN(n4694) );
  INV_X1 U5218 ( .A(n6556), .ZN(n4698) );
  AND2_X1 U5219 ( .A1(n6550), .A2(n6549), .ZN(n9225) );
  NAND2_X1 U5220 ( .A1(n6666), .A2(n6665), .ZN(n9261) );
  NOR2_X1 U5221 ( .A1(n9271), .A2(n4708), .ZN(n4707) );
  INV_X1 U5222 ( .A(n9216), .ZN(n4708) );
  NOR2_X1 U5223 ( .A1(n9271), .A2(n6715), .ZN(n4706) );
  AND2_X1 U5224 ( .A1(n9294), .A2(n4712), .ZN(n4704) );
  OR2_X1 U5225 ( .A1(n6548), .A2(n6547), .ZN(n6550) );
  AND2_X1 U5226 ( .A1(n4702), .A2(n4699), .ZN(n6520) );
  NAND2_X1 U5227 ( .A1(n6696), .A2(n9281), .ZN(n9284) );
  INV_X1 U5228 ( .A(n7681), .ZN(n4383) );
  NAND2_X1 U5229 ( .A1(n6539), .A2(n6538), .ZN(n6991) );
  OR2_X1 U5230 ( .A1(n6675), .A2(n6676), .ZN(n9304) );
  INV_X1 U5231 ( .A(n5086), .ZN(n5350) );
  INV_X1 U5232 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4999) );
  NAND2_X1 U5233 ( .A1(n6841), .A2(n9831), .ZN(n6844) );
  OR2_X1 U5234 ( .A1(n6939), .A2(n6938), .ZN(n4419) );
  NOR2_X1 U5235 ( .A1(n7248), .A2(n4425), .ZN(n7250) );
  AND2_X1 U5236 ( .A1(n7249), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4425) );
  XNOR2_X1 U5237 ( .A(n9375), .B(n9374), .ZN(n9885) );
  NOR2_X1 U5238 ( .A1(n9885), .A2(n9884), .ZN(n9883) );
  NAND2_X1 U5239 ( .A1(n8346), .A2(n8345), .ZN(n9410) );
  NAND2_X1 U5240 ( .A1(n4557), .A2(n8593), .ZN(n4559) );
  INV_X1 U5241 ( .A(n4559), .ZN(n9446) );
  INV_X1 U5242 ( .A(n4561), .ZN(n9473) );
  AND2_X1 U5243 ( .A1(n8412), .A2(n8351), .ZN(n9489) );
  AND4_X1 U5244 ( .A1(n5026), .A2(n5025), .A3(n5024), .A4(n5023), .ZN(n9505)
         );
  AND2_X1 U5245 ( .A1(n8515), .A2(n8508), .ZN(n9503) );
  NAND2_X1 U5246 ( .A1(n4872), .A2(n5338), .ZN(n4859) );
  INV_X1 U5247 ( .A(n8365), .ZN(n4831) );
  INV_X1 U5248 ( .A(n9574), .ZN(n4832) );
  AND2_X1 U5249 ( .A1(n8500), .A2(n8502), .ZN(n9547) );
  OR2_X1 U5250 ( .A1(n8206), .A2(n9551), .ZN(n4870) );
  NAND2_X1 U5251 ( .A1(n4832), .A2(n9561), .ZN(n4835) );
  AND2_X1 U5252 ( .A1(n4570), .A2(n8481), .ZN(n9574) );
  INV_X1 U5253 ( .A(n4835), .ZN(n9571) );
  AOI21_X1 U5254 ( .B1(n7582), .B2(n5201), .A(n5200), .ZN(n7597) );
  AND2_X1 U5255 ( .A1(n5141), .A2(n5128), .ZN(n4862) );
  INV_X1 U5256 ( .A(n8569), .ZN(n5141) );
  NAND2_X1 U5257 ( .A1(n7021), .A2(n5507), .ZN(n8380) );
  OR2_X1 U5258 ( .A1(n6767), .A2(n6951), .ZN(n9550) );
  INV_X1 U5259 ( .A(n7018), .ZN(n7023) );
  AND2_X1 U5260 ( .A1(n6526), .A2(n6519), .ZN(n7020) );
  NAND2_X1 U5261 ( .A1(n9591), .A2(n9670), .ZN(n4539) );
  INV_X1 U5262 ( .A(n9592), .ZN(n4540) );
  INV_X1 U5263 ( .A(n9512), .ZN(n9629) );
  NAND2_X1 U5264 ( .A1(n5328), .A2(n5327), .ZN(n9637) );
  OR2_X1 U5265 ( .A1(n6807), .A2(n5165), .ZN(n4571) );
  NOR2_X1 U5266 ( .A1(n4334), .A2(n4573), .ZN(n4572) );
  NOR2_X1 U5267 ( .A1(n5140), .A2(n6808), .ZN(n4573) );
  OR2_X1 U5268 ( .A1(n8556), .A2(n8647), .ZN(n7210) );
  AND3_X1 U5269 ( .A1(n4771), .A2(n4769), .A3(n4767), .ZN(n9203) );
  XNOR2_X1 U5270 ( .A(n6156), .B(n6155), .ZN(n9209) );
  NAND2_X1 U5271 ( .A1(n4801), .A2(n5448), .ZN(n6156) );
  NAND2_X1 U5272 ( .A1(n5003), .A2(n5005), .ZN(n5006) );
  NOR2_X1 U5273 ( .A1(n5004), .A2(n9695), .ZN(n5005) );
  XNOR2_X1 U5274 ( .A(n4522), .B(n5268), .ZN(n7240) );
  INV_X1 U5275 ( .A(n4517), .ZN(n4516) );
  OAI21_X1 U5276 ( .B1(n4520), .B2(n4518), .A(n4950), .ZN(n4517) );
  NOR2_X1 U5277 ( .A1(n5207), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5236) );
  INV_X1 U5278 ( .A(n4506), .ZN(n5188) );
  AOI21_X1 U5279 ( .B1(n4816), .B2(n4510), .A(n4509), .ZN(n4506) );
  XNOR2_X1 U5280 ( .A(n5172), .B(n5171), .ZN(n6823) );
  CLKBUF_X1 U5281 ( .A(n5011), .Z(n6799) );
  OR2_X1 U5282 ( .A1(n7312), .A2(n7313), .ZN(n7310) );
  INV_X1 U5283 ( .A(n9071), .ZN(n8807) );
  NAND2_X1 U5284 ( .A1(n7234), .A2(n7235), .ZN(n7233) );
  INV_X1 U5285 ( .A(n10002), .ZN(n8836) );
  NAND2_X1 U5286 ( .A1(n5865), .A2(n5864), .ZN(n8833) );
  NAND2_X1 U5287 ( .A1(n4501), .A2(n6374), .ZN(n4500) );
  NAND4_X1 U5288 ( .A1(n5724), .A2(n5723), .A3(n5722), .A4(n5721), .ZN(n8856)
         );
  NOR2_X1 U5289 ( .A1(n7076), .A2(n4330), .ZN(n7045) );
  AND2_X1 U5290 ( .A1(n5713), .A2(n5712), .ZN(n7180) );
  AOI21_X1 U5291 ( .B1(n8692), .B2(n9084), .A(n8691), .ZN(n9103) );
  NAND2_X1 U5292 ( .A1(n8690), .A2(n8689), .ZN(n8691) );
  OAI21_X1 U5293 ( .B1(n4658), .B2(n8677), .A(n4651), .ZN(n4650) );
  OR2_X1 U5294 ( .A1(n8951), .A2(n4655), .ZN(n4654) );
  NAND2_X1 U5295 ( .A1(n9079), .A2(n10018), .ZN(n9094) );
  INV_X1 U5296 ( .A(n4721), .ZN(n4718) );
  NOR2_X1 U5297 ( .A1(n4722), .A2(n9315), .ZN(n4720) );
  INV_X1 U5298 ( .A(n4723), .ZN(n4722) );
  AOI21_X1 U5299 ( .B1(n4727), .B2(n4726), .A(n4724), .ZN(n4723) );
  OAI21_X1 U5300 ( .B1(n4721), .B2(n4717), .A(n4375), .ZN(n4716) );
  INV_X1 U5301 ( .A(n4727), .ZN(n4717) );
  INV_X1 U5302 ( .A(n6529), .ZN(n7134) );
  AND2_X1 U5303 ( .A1(n8652), .A2(n4364), .ZN(n4411) );
  NAND2_X1 U5304 ( .A1(n9903), .A2(n9902), .ZN(n9901) );
  INV_X1 U5305 ( .A(n4840), .ZN(n9426) );
  AOI21_X1 U5306 ( .B1(n9445), .B2(n4845), .A(n4842), .ZN(n4840) );
  NAND2_X1 U5307 ( .A1(n9460), .A2(n4838), .ZN(n4837) );
  AOI21_X1 U5308 ( .B1(n4843), .B2(n4844), .A(n8539), .ZN(n4841) );
  INV_X1 U5309 ( .A(n8350), .ZN(n9619) );
  INV_X1 U5310 ( .A(n9568), .ZN(n9941) );
  NAND2_X1 U5311 ( .A1(n4452), .A2(n4450), .ZN(n6252) );
  NAND2_X1 U5312 ( .A1(n6228), .A2(n4453), .ZN(n4452) );
  NAND2_X1 U5313 ( .A1(n4451), .A2(n6372), .ZN(n4450) );
  NAND2_X1 U5314 ( .A1(n6245), .A2(n6249), .ZN(n4451) );
  NAND2_X1 U5315 ( .A1(n6244), .A2(n6250), .ZN(n6258) );
  NOR2_X1 U5316 ( .A1(n6276), .A2(n4453), .ZN(n4427) );
  OR2_X1 U5317 ( .A1(n6273), .A2(n6274), .ZN(n4428) );
  OR2_X1 U5318 ( .A1(n6294), .A2(n6293), .ZN(n4878) );
  NAND2_X1 U5319 ( .A1(n4494), .A2(n6318), .ZN(n4493) );
  OR2_X1 U5320 ( .A1(n8495), .A2(n8494), .ZN(n4409) );
  AND2_X1 U5321 ( .A1(n6324), .A2(n4453), .ZN(n4444) );
  AND2_X1 U5322 ( .A1(n6330), .A2(n6318), .ZN(n4491) );
  NOR2_X1 U5323 ( .A1(n4449), .A2(n6145), .ZN(n4448) );
  INV_X1 U5324 ( .A(n6333), .ZN(n4449) );
  OR2_X1 U5325 ( .A1(n6323), .A2(n4453), .ZN(n4446) );
  OAI211_X1 U5326 ( .C1(n4407), .C2(n8503), .A(n8502), .B(n8501), .ZN(n4406)
         );
  NAND2_X1 U5327 ( .A1(n4405), .A2(n4403), .ZN(n8514) );
  NAND2_X1 U5328 ( .A1(n4404), .A2(n8556), .ZN(n4403) );
  NAND2_X1 U5329 ( .A1(n4406), .A2(n8536), .ZN(n4405) );
  OAI21_X1 U5330 ( .B1(n4407), .B2(n8505), .A(n8504), .ZN(n4404) );
  NAND2_X1 U5331 ( .A1(n6335), .A2(n4442), .ZN(n6340) );
  NOR2_X1 U5332 ( .A1(n8526), .A2(n8536), .ZN(n4399) );
  INV_X1 U5333 ( .A(n5448), .ZN(n4804) );
  NOR2_X1 U5334 ( .A1(n9096), .A2(n8913), .ZN(n6364) );
  INV_X1 U5335 ( .A(SI_12_), .ZN(n6424) );
  AND2_X1 U5336 ( .A1(n8682), .A2(n8839), .ZN(n6359) );
  NOR2_X1 U5337 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5564) );
  INV_X1 U5338 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4458) );
  OR2_X1 U5339 ( .A1(n6676), .A2(n4688), .ZN(n4687) );
  INV_X1 U5340 ( .A(n9306), .ZN(n4688) );
  INV_X1 U5341 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n4951) );
  INV_X1 U5342 ( .A(SI_9_), .ZN(n4919) );
  INV_X1 U5343 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n4912) );
  AND2_X1 U5344 ( .A1(n9207), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n4612) );
  NOR2_X1 U5345 ( .A1(n9712), .A2(n4478), .ZN(n9710) );
  NAND2_X1 U5346 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n4478) );
  NAND2_X1 U5347 ( .A1(n4759), .A2(n6341), .ZN(n4758) );
  INV_X1 U5348 ( .A(n6359), .ZN(n6202) );
  NAND2_X1 U5349 ( .A1(n4662), .A2(n8924), .ZN(n4661) );
  NOR2_X1 U5350 ( .A1(n4329), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n5569) );
  NOR2_X1 U5351 ( .A1(n5867), .A2(n8827), .ZN(n5853) );
  NAND2_X1 U5352 ( .A1(n8153), .A2(n6303), .ZN(n4740) );
  INV_X1 U5353 ( .A(n6293), .ZN(n6303) );
  OR2_X1 U5354 ( .A1(n8833), .A2(n8228), .ZN(n6305) );
  INV_X1 U5355 ( .A(n4633), .ZN(n4631) );
  INV_X1 U5356 ( .A(n7559), .ZN(n4462) );
  AND2_X1 U5357 ( .A1(n10062), .A2(n10076), .ZN(n4463) );
  AND2_X1 U5358 ( .A1(n8702), .A2(n4466), .ZN(n7637) );
  NOR2_X1 U5359 ( .A1(n7559), .A2(n6119), .ZN(n4466) );
  AND2_X1 U5360 ( .A1(n7745), .A2(n10027), .ZN(n6108) );
  INV_X1 U5361 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4753) );
  INV_X1 U5362 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4456) );
  OAI21_X1 U5363 ( .B1(n6068), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6087) );
  INV_X1 U5364 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6086) );
  AND2_X1 U5365 ( .A1(n5656), .A2(n5540), .ZN(n4874) );
  INV_X1 U5366 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5656) );
  OR2_X1 U5367 ( .A1(n6555), .A2(n6554), .ZN(n6556) );
  AND2_X1 U5368 ( .A1(n4684), .A2(n6705), .ZN(n4683) );
  NOR2_X2 U5369 ( .A1(n6517), .A2(n6528), .ZN(n8324) );
  NOR2_X1 U5370 ( .A1(n6516), .A2(n6746), .ZN(n6517) );
  AND2_X1 U5371 ( .A1(n8539), .A2(n8538), .ZN(n4396) );
  INV_X1 U5372 ( .A(n9477), .ZN(n5395) );
  NOR2_X1 U5373 ( .A1(n9644), .A2(n9647), .ZN(n4528) );
  AND3_X1 U5374 ( .A1(n4532), .A2(n9783), .A3(n4531), .ZN(n4536) );
  NOR2_X1 U5375 ( .A1(n9478), .A2(n9612), .ZN(n9451) );
  NOR2_X1 U5376 ( .A1(n9506), .A2(n9624), .ZN(n9494) );
  AND2_X1 U5377 ( .A1(n9563), .A2(n4325), .ZN(n9523) );
  OR2_X1 U5378 ( .A1(n7358), .A2(n7357), .ZN(n7360) );
  NAND2_X1 U5379 ( .A1(n8555), .A2(n9497), .ZN(n8556) );
  AND2_X1 U5380 ( .A1(n6157), .A2(n5453), .ZN(n6155) );
  NOR2_X1 U5381 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n5002) );
  AND2_X1 U5382 ( .A1(n5448), .A2(n5438), .ZN(n5446) );
  XNOR2_X1 U5383 ( .A(n5470), .B(P1_IR_REG_21__SCAN_IN), .ZN(n5506) );
  OAI21_X1 U5384 ( .B1(n5031), .B2(n5030), .A(n4968), .ZN(n5326) );
  AND2_X1 U5385 ( .A1(n4972), .A2(n4971), .ZN(n5325) );
  INV_X1 U5386 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5299) );
  AOI21_X1 U5387 ( .B1(n4791), .B2(n4790), .A(n4376), .ZN(n4789) );
  AOI21_X1 U5388 ( .B1(n4796), .B2(n4795), .A(n4794), .ZN(n4793) );
  INV_X1 U5389 ( .A(n4956), .ZN(n4794) );
  INV_X1 U5390 ( .A(n4950), .ZN(n4795) );
  INV_X1 U5391 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5038) );
  NOR2_X1 U5392 ( .A1(n4945), .A2(n4521), .ZN(n4520) );
  INV_X1 U5393 ( .A(n4940), .ZN(n4521) );
  NAND2_X1 U5394 ( .A1(n4519), .A2(n4944), .ZN(n4518) );
  INV_X1 U5395 ( .A(n5278), .ZN(n4519) );
  AOI21_X1 U5396 ( .B1(n4808), .B2(n4810), .A(n4807), .ZN(n4806) );
  INV_X1 U5397 ( .A(n5261), .ZN(n4807) );
  INV_X1 U5398 ( .A(n5171), .ZN(n4511) );
  AOI21_X1 U5399 ( .B1(n4513), .B2(n5150), .A(n4355), .ZN(n4512) );
  INV_X1 U5400 ( .A(n4906), .ZN(n4513) );
  OAI211_X1 U5401 ( .C1(n4310), .C2(P1_DATAO_REG_3__SCAN_IN), .A(n4575), .B(
        n4574), .ZN(n4898) );
  NAND2_X1 U5402 ( .A1(n4672), .A2(n6793), .ZN(n4575) );
  OAI211_X1 U5403 ( .C1(n4310), .C2(P1_DATAO_REG_2__SCAN_IN), .A(n4671), .B(
        n4670), .ZN(n4893) );
  NAND2_X1 U5404 ( .A1(n4672), .A2(n6794), .ZN(n4671) );
  NAND2_X1 U5405 ( .A1(n5597), .A2(n5094), .ZN(n4890) );
  NAND2_X1 U5406 ( .A1(n5820), .A2(n4598), .ZN(n8255) );
  NOR2_X1 U5407 ( .A1(n7514), .A2(n4592), .ZN(n4591) );
  INV_X1 U5408 ( .A(n5683), .ZN(n4592) );
  AND2_X1 U5409 ( .A1(n5957), .A2(n4582), .ZN(n4581) );
  INV_X1 U5410 ( .A(n8728), .ZN(n4586) );
  AND2_X1 U5411 ( .A1(n4584), .A2(n8729), .ZN(n4583) );
  NAND2_X1 U5412 ( .A1(n8728), .A2(n4585), .ZN(n4584) );
  INV_X1 U5413 ( .A(n5915), .ZN(n4585) );
  NAND2_X1 U5414 ( .A1(n8035), .A2(n8038), .ZN(n4579) );
  OR2_X1 U5415 ( .A1(n5960), .A2(n8799), .ZN(n5978) );
  NAND2_X1 U5416 ( .A1(n5784), .A2(n5783), .ZN(n8036) );
  NOR2_X1 U5417 ( .A1(n5668), .A2(n5667), .ZN(n5694) );
  INV_X1 U5418 ( .A(n4609), .ZN(n4603) );
  NOR2_X1 U5419 ( .A1(n8750), .A2(n4606), .ZN(n4605) );
  INV_X1 U5420 ( .A(n4608), .ZN(n4606) );
  NAND2_X1 U5421 ( .A1(n8255), .A2(n5843), .ZN(n8761) );
  NOR2_X1 U5422 ( .A1(n4502), .A2(n6200), .ZN(n4501) );
  INV_X1 U5423 ( .A(n7332), .ZN(n4502) );
  NAND2_X1 U5424 ( .A1(n4438), .A2(n4437), .ZN(n4436) );
  NOR2_X1 U5425 ( .A1(n6369), .A2(n4453), .ZN(n4437) );
  AND2_X1 U5426 ( .A1(n4487), .A2(n4486), .ZN(n7178) );
  NAND2_X1 U5427 ( .A1(n7148), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4486) );
  NOR2_X1 U5428 ( .A1(n7178), .A2(n7177), .ZN(n7176) );
  NOR2_X1 U5429 ( .A1(n7649), .A2(n4489), .ZN(n7653) );
  AND2_X1 U5430 ( .A1(n7650), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4489) );
  NAND2_X1 U5431 ( .A1(n7653), .A2(n7652), .ZN(n7782) );
  OR2_X1 U5432 ( .A1(n5806), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5807) );
  NAND2_X1 U5433 ( .A1(n7782), .A2(n4488), .ZN(n7786) );
  OR2_X1 U5434 ( .A1(n7783), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4488) );
  NAND2_X1 U5435 ( .A1(n7786), .A2(n7785), .ZN(n7939) );
  INV_X1 U5436 ( .A(n4482), .ZN(n8894) );
  NAND2_X1 U5437 ( .A1(n6191), .A2(n6190), .ZN(n6193) );
  AND2_X1 U5438 ( .A1(n4769), .A2(n6188), .ZN(n4768) );
  NOR2_X1 U5439 ( .A1(n9097), .A2(n4471), .ZN(n4470) );
  NAND2_X1 U5440 ( .A1(n4472), .A2(n8943), .ZN(n4471) );
  INV_X1 U5441 ( .A(n4473), .ZN(n4472) );
  NOR2_X1 U5442 ( .A1(n8938), .A2(n9109), .ZN(n8931) );
  NAND2_X1 U5443 ( .A1(n8840), .A2(n9070), .ZN(n8690) );
  NAND2_X1 U5444 ( .A1(n4656), .A2(n8677), .ZN(n4655) );
  INV_X1 U5445 ( .A(n4661), .ZN(n4656) );
  NAND2_X1 U5446 ( .A1(n4658), .A2(n4652), .ZN(n4651) );
  NAND2_X1 U5447 ( .A1(n4661), .A2(n8683), .ZN(n4652) );
  AOI21_X1 U5448 ( .B1(n4662), .B2(n4660), .A(n4659), .ZN(n4658) );
  NOR2_X1 U5449 ( .A1(n9109), .A2(n8840), .ZN(n4659) );
  NOR2_X1 U5450 ( .A1(n8927), .A2(n4664), .ZN(n4660) );
  NOR2_X1 U5451 ( .A1(n8969), .A2(n9119), .ZN(n8957) );
  OR2_X1 U5452 ( .A1(n5999), .A2(n5998), .ZN(n6016) );
  INV_X1 U5453 ( .A(n8841), .ZN(n8956) );
  NAND2_X1 U5454 ( .A1(n4756), .A2(n4755), .ZN(n4754) );
  NAND2_X1 U5455 ( .A1(n9020), .A2(n4756), .ZN(n8992) );
  NOR2_X1 U5456 ( .A1(n9008), .A2(n9127), .ZN(n8983) );
  NOR2_X1 U5457 ( .A1(n9026), .A2(n9135), .ZN(n8678) );
  NAND2_X1 U5458 ( .A1(n5934), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5952) );
  INV_X1 U5459 ( .A(n5936), .ZN(n5934) );
  NAND2_X1 U5460 ( .A1(n4746), .A2(n4744), .ZN(n9046) );
  AOI21_X1 U5461 ( .B1(n4747), .B2(n4750), .A(n4745), .ZN(n4744) );
  INV_X1 U5462 ( .A(n6318), .ZN(n4745) );
  NAND2_X1 U5463 ( .A1(n8282), .A2(n4321), .ZN(n9058) );
  NAND2_X1 U5464 ( .A1(n8282), .A2(n4317), .ZN(n9086) );
  NAND2_X1 U5465 ( .A1(n6140), .A2(n6315), .ZN(n9081) );
  NAND2_X1 U5466 ( .A1(n9081), .A2(n9082), .ZN(n9080) );
  OR2_X1 U5467 ( .A1(n5922), .A2(n6488), .ZN(n5936) );
  AND2_X1 U5468 ( .A1(n6141), .A2(n9064), .ZN(n9082) );
  NAND2_X1 U5469 ( .A1(n8282), .A2(n4469), .ZN(n9088) );
  AOI21_X1 U5470 ( .B1(n4622), .B2(n4624), .A(n4348), .ZN(n4621) );
  INV_X1 U5471 ( .A(n4624), .ZN(n4623) );
  OR2_X1 U5472 ( .A1(n5889), .A2(n8313), .ZN(n5906) );
  AND2_X1 U5473 ( .A1(n8282), .A2(n8292), .ZN(n8299) );
  OR2_X1 U5474 ( .A1(n8162), .A2(n8833), .ZN(n8232) );
  INV_X1 U5475 ( .A(n8848), .ZN(n8828) );
  NAND2_X1 U5476 ( .A1(n8057), .A2(n6289), .ZN(n8153) );
  NAND2_X1 U5477 ( .A1(n5791), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5831) );
  INV_X1 U5478 ( .A(n5792), .ZN(n5791) );
  AND2_X1 U5479 ( .A1(n7889), .A2(n4362), .ZN(n8061) );
  INV_X1 U5480 ( .A(n6270), .ZN(n8071) );
  NAND2_X1 U5481 ( .A1(n7889), .A2(n10089), .ZN(n8018) );
  NAND2_X1 U5482 ( .A1(n7889), .A2(n4461), .ZN(n8078) );
  NAND2_X1 U5483 ( .A1(n4617), .A2(n7878), .ZN(n4868) );
  INV_X1 U5484 ( .A(n5736), .ZN(n5735) );
  CLKBUF_X1 U5485 ( .A(n7882), .Z(n8009) );
  INV_X1 U5486 ( .A(n8853), .ZN(n8075) );
  NOR2_X1 U5487 ( .A1(n7866), .A2(n7957), .ZN(n7889) );
  NAND2_X1 U5488 ( .A1(n4357), .A2(n6260), .ZN(n4742) );
  NAND2_X1 U5489 ( .A1(n8702), .A2(n4464), .ZN(n7797) );
  NOR2_X1 U5490 ( .A1(n4465), .A2(n7559), .ZN(n4464) );
  NAND2_X1 U5491 ( .A1(n10062), .A2(n10076), .ZN(n4465) );
  AND2_X1 U5492 ( .A1(n6206), .A2(n4733), .ZN(n4732) );
  NOR2_X1 U5493 ( .A1(n4737), .A2(n4738), .ZN(n4735) );
  NAND2_X1 U5494 ( .A1(n8702), .A2(n10062), .ZN(n7753) );
  OAI211_X1 U5495 ( .C1(n6811), .C2(n5685), .A(n5611), .B(n5610), .ZN(n6116)
         );
  AND2_X1 U5496 ( .A1(n8704), .A2(n10058), .ZN(n8702) );
  AND3_X1 U5497 ( .A1(n4880), .A2(n5627), .A3(n5626), .ZN(n8699) );
  OR2_X1 U5498 ( .A1(n6173), .A2(n7050), .ZN(n5626) );
  AND2_X1 U5499 ( .A1(n10034), .A2(n10040), .ZN(n6084) );
  AND2_X1 U5500 ( .A1(n4639), .A2(n4359), .ZN(n9138) );
  NAND2_X1 U5501 ( .A1(n4636), .A2(n4634), .ZN(n8056) );
  NAND2_X1 U5502 ( .A1(n4636), .A2(n4637), .ZN(n7992) );
  NAND2_X1 U5503 ( .A1(n5771), .A2(n5770), .ZN(n8040) );
  INV_X1 U5504 ( .A(n7756), .ZN(n10071) );
  INV_X1 U5505 ( .A(n9181), .ZN(n10097) );
  AND2_X1 U5506 ( .A1(n7543), .A2(n7542), .ZN(n7574) );
  AND3_X1 U5507 ( .A1(n4752), .A2(n4314), .A3(n4751), .ZN(n6064) );
  INV_X1 U5508 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6069) );
  AND2_X1 U5509 ( .A1(n5751), .A2(n5766), .ZN(n7268) );
  INV_X1 U5510 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5746) );
  AND2_X1 U5511 ( .A1(n5711), .A2(n5710), .ZN(n5747) );
  AND2_X1 U5512 ( .A1(n4730), .A2(n4731), .ZN(n5638) );
  NAND2_X1 U5513 ( .A1(n4729), .A2(n4728), .ZN(n4727) );
  INV_X1 U5514 ( .A(n9319), .ZN(n4728) );
  INV_X1 U5515 ( .A(n9318), .ZN(n4729) );
  INV_X1 U5516 ( .A(n5372), .ZN(n5370) );
  NAND2_X1 U5517 ( .A1(n4724), .A2(n4726), .ZN(n4725) );
  NAND2_X1 U5518 ( .A1(n4694), .A2(n7415), .ZN(n4691) );
  INV_X1 U5519 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5180) );
  NAND2_X1 U5520 ( .A1(n5370), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5390) );
  INV_X1 U5521 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5193) );
  NOR2_X1 U5522 ( .A1(n5194), .A2(n5193), .ZN(n5212) );
  OR2_X1 U5523 ( .A1(n5330), .A2(n5329), .ZN(n5344) );
  AND2_X1 U5524 ( .A1(n5212), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5224) );
  AND2_X1 U5525 ( .A1(n6753), .A2(n9951), .ZN(n6895) );
  NOR2_X1 U5526 ( .A1(n5144), .A2(n5143), .ZN(n5157) );
  OR2_X1 U5527 ( .A1(n6751), .A2(n6748), .ZN(n6758) );
  AND4_X1 U5528 ( .A1(n5463), .A2(n5462), .A3(n5461), .A4(n5460), .ZN(n9418)
         );
  NAND2_X1 U5529 ( .A1(n6877), .A2(n6950), .ZN(n6876) );
  OR2_X1 U5530 ( .A1(n6954), .A2(n6840), .ZN(n6956) );
  NOR2_X1 U5531 ( .A1(n6921), .A2(n6920), .ZN(n9843) );
  NOR2_X1 U5532 ( .A1(n6932), .A2(n4421), .ZN(n9846) );
  NOR2_X1 U5533 ( .A1(n6842), .A2(n4422), .ZN(n4421) );
  INV_X1 U5534 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n4422) );
  NAND2_X1 U5535 ( .A1(n9846), .A2(n9847), .ZN(n9845) );
  NAND2_X1 U5536 ( .A1(n9845), .A2(n4420), .ZN(n9861) );
  OR2_X1 U5537 ( .A1(n6934), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4420) );
  NAND2_X1 U5538 ( .A1(n9861), .A2(n9860), .ZN(n9859) );
  AND2_X1 U5539 ( .A1(n4419), .A2(n4418), .ZN(n6983) );
  NAND2_X1 U5540 ( .A1(n6982), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4418) );
  NAND2_X1 U5541 ( .A1(n6983), .A2(n6984), .ZN(n7165) );
  NAND2_X1 U5542 ( .A1(n7165), .A2(n4417), .ZN(n7169) );
  OR2_X1 U5543 ( .A1(n7166), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4417) );
  NOR2_X1 U5544 ( .A1(n7250), .A2(n7251), .ZN(n7610) );
  NOR2_X1 U5545 ( .A1(n7610), .A2(n4424), .ZN(n9371) );
  AND2_X1 U5546 ( .A1(n7611), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4424) );
  AOI21_X1 U5547 ( .B1(n9776), .B2(n7617), .A(n7616), .ZN(n7620) );
  NOR2_X1 U5548 ( .A1(n9883), .A2(n9376), .ZN(n9897) );
  INV_X1 U5549 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5302) );
  NOR2_X1 U5550 ( .A1(n9909), .A2(n4416), .ZN(n9379) );
  AND2_X1 U5551 ( .A1(n9914), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4416) );
  NAND2_X1 U5552 ( .A1(n5483), .A2(n4339), .ZN(n5008) );
  NOR2_X1 U5553 ( .A1(n9379), .A2(n9380), .ZN(n9388) );
  OAI21_X1 U5554 ( .B1(n5519), .B2(n4827), .A(n4826), .ZN(n4825) );
  OR2_X1 U5555 ( .A1(n9416), .A2(n4829), .ZN(n4824) );
  NAND2_X1 U5556 ( .A1(n8596), .A2(n8541), .ZN(n4829) );
  NOR2_X1 U5557 ( .A1(n9414), .A2(n9591), .ZN(n9408) );
  INV_X1 U5558 ( .A(n4843), .ZN(n4842) );
  AOI22_X1 U5559 ( .A1(n9431), .A2(n4846), .B1(n4845), .B2(n8593), .ZN(n4843)
         );
  NOR2_X1 U5560 ( .A1(n4842), .A2(n4839), .ZN(n4838) );
  NAND2_X1 U5561 ( .A1(n9451), .A2(n4848), .ZN(n9452) );
  NOR2_X1 U5562 ( .A1(n9601), .A2(n9452), .ZN(n9433) );
  NAND2_X1 U5563 ( .A1(n4848), .A2(n9465), .ZN(n4847) );
  AND4_X1 U5564 ( .A1(n5429), .A2(n5428), .A3(n5427), .A4(n5426), .ZN(n9450)
         );
  NAND2_X1 U5565 ( .A1(n4561), .A2(n4343), .ZN(n9467) );
  NAND2_X1 U5566 ( .A1(n9494), .A2(n8350), .ZN(n9478) );
  NAND2_X1 U5567 ( .A1(n9472), .A2(n4879), .ZN(n4389) );
  AND2_X1 U5568 ( .A1(n5013), .A2(n5012), .ZN(n6713) );
  NOR2_X1 U5569 ( .A1(n4877), .A2(n9298), .ZN(n5359) );
  AND4_X1 U5570 ( .A1(n5363), .A2(n5362), .A3(n5361), .A4(n5360), .ZN(n9522)
         );
  AND2_X1 U5571 ( .A1(n4545), .A2(n4363), .ZN(n4544) );
  NAND2_X1 U5572 ( .A1(n4832), .A2(n4549), .ZN(n4546) );
  INV_X1 U5573 ( .A(n4552), .ZN(n4551) );
  INV_X1 U5574 ( .A(n4553), .ZN(n4548) );
  OAI21_X1 U5575 ( .B1(n4832), .B2(n4551), .A(n4549), .ZN(n9540) );
  NAND2_X1 U5576 ( .A1(n9563), .A2(n4526), .ZN(n9531) );
  AND2_X1 U5577 ( .A1(n5319), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5321) );
  AOI21_X1 U5578 ( .B1(n8129), .B2(n4860), .A(n5312), .ZN(n8210) );
  NOR2_X1 U5579 ( .A1(n4861), .A2(n4331), .ZN(n4860) );
  NAND2_X1 U5580 ( .A1(n9563), .A2(n8206), .ZN(n9553) );
  AND4_X1 U5581 ( .A1(n5277), .A2(n5276), .A3(n5275), .A4(n5274), .ZN(n9570)
         );
  OR2_X1 U5582 ( .A1(n5285), .A2(n5272), .ZN(n5308) );
  NOR2_X1 U5583 ( .A1(n8132), .A2(n8133), .ZN(n4566) );
  INV_X1 U5584 ( .A(n4567), .ZN(n8134) );
  NOR2_X1 U5585 ( .A1(n5254), .A2(n5051), .ZN(n5284) );
  AOI21_X1 U5586 ( .B1(n9749), .B2(n5250), .A(n7813), .ZN(n4864) );
  NOR2_X1 U5587 ( .A1(n4534), .A2(n7604), .ZN(n7973) );
  NAND2_X1 U5588 ( .A1(n4536), .A2(n4535), .ZN(n4534) );
  NAND2_X1 U5589 ( .A1(n9744), .A2(n5250), .ZN(n7896) );
  OR2_X1 U5590 ( .A1(n5252), .A2(n5251), .ZN(n5254) );
  AND2_X1 U5591 ( .A1(n8470), .A2(n8366), .ZN(n8581) );
  NAND2_X1 U5592 ( .A1(n4533), .A2(n4536), .ZN(n9763) );
  NAND2_X1 U5593 ( .A1(n5224), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5244) );
  INV_X1 U5594 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5243) );
  NAND2_X1 U5595 ( .A1(n4533), .A2(n4537), .ZN(n9762) );
  NOR2_X1 U5596 ( .A1(n6600), .A2(n7707), .ZN(n4537) );
  AND4_X1 U5597 ( .A1(n5217), .A2(n5216), .A3(n5215), .A4(n5214), .ZN(n7736)
         );
  NAND2_X1 U5598 ( .A1(n4821), .A2(n5179), .ZN(n7498) );
  NAND2_X1 U5599 ( .A1(n6823), .A2(n5454), .ZN(n4821) );
  NAND2_X1 U5600 ( .A1(n7395), .A2(n5170), .ZN(n7484) );
  NAND2_X1 U5601 ( .A1(n7397), .A2(n7396), .ZN(n7395) );
  AND4_X1 U5602 ( .A1(n5186), .A2(n5185), .A3(n5184), .A4(n5183), .ZN(n7589)
         );
  NOR2_X1 U5603 ( .A1(n7360), .A2(n9925), .ZN(n7443) );
  AND2_X1 U5604 ( .A1(n7443), .A2(n9967), .ZN(n7445) );
  NAND2_X1 U5605 ( .A1(n7282), .A2(n5142), .ZN(n7435) );
  NAND2_X1 U5606 ( .A1(n7347), .A2(n8566), .ZN(n7349) );
  NAND2_X1 U5607 ( .A1(n7455), .A2(n7132), .ZN(n7358) );
  NAND2_X1 U5608 ( .A1(n7131), .A2(n8565), .ZN(n7130) );
  OR2_X1 U5609 ( .A1(n5526), .A2(n5103), .ZN(n5105) );
  INV_X1 U5610 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n5097) );
  NAND2_X1 U5611 ( .A1(n5140), .A2(n9709), .ZN(n5096) );
  NAND2_X1 U5612 ( .A1(n5283), .A2(n5282), .ZN(n9662) );
  NAND2_X1 U5613 ( .A1(n5050), .A2(n5049), .ZN(n9669) );
  AOI22_X1 U5614 ( .A1(n5113), .A2(n5114), .B1(n6909), .B2(n6769), .ZN(n4541)
         );
  INV_X1 U5615 ( .A(n9670), .ZN(n9973) );
  XNOR2_X1 U5616 ( .A(n6183), .B(SI_30_), .ZN(n9206) );
  XNOR2_X1 U5617 ( .A(n5447), .B(n5446), .ZN(n8309) );
  NAND2_X1 U5618 ( .A1(n4777), .A2(n4775), .ZN(n5431) );
  AOI21_X1 U5619 ( .B1(n4779), .B2(n4782), .A(n4776), .ZN(n4775) );
  INV_X1 U5620 ( .A(n5415), .ZN(n4776) );
  AND2_X1 U5621 ( .A1(n5432), .A2(n5419), .ZN(n5430) );
  NAND2_X1 U5622 ( .A1(n5383), .A2(n4785), .ZN(n4778) );
  NAND2_X1 U5623 ( .A1(n4676), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5480) );
  INV_X1 U5624 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5479) );
  XNOR2_X1 U5625 ( .A(n5399), .B(n5398), .ZN(n8214) );
  NAND2_X1 U5626 ( .A1(n4787), .A2(n5381), .ZN(n5399) );
  INV_X1 U5627 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5471) );
  NAND2_X1 U5628 ( .A1(n4805), .A2(n4808), .ZN(n5262) );
  NAND2_X1 U5629 ( .A1(n5220), .A2(n4811), .ZN(n4805) );
  AND2_X1 U5630 ( .A1(n5263), .A2(n5240), .ZN(n7249) );
  NAND2_X1 U5631 ( .A1(n4813), .A2(n4931), .ZN(n5234) );
  NAND2_X1 U5632 ( .A1(n4814), .A2(n5219), .ZN(n4813) );
  INV_X1 U5633 ( .A(n5220), .ZN(n4814) );
  OR3_X1 U5634 ( .A1(n5205), .A2(P1_IR_REG_7__SCAN_IN), .A3(n5204), .ZN(n5207)
         );
  INV_X1 U5635 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5176) );
  NOR2_X1 U5636 ( .A1(n5067), .A2(n5000), .ZN(n6851) );
  XNOR2_X1 U5637 ( .A(n4423), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6849) );
  NAND2_X1 U5638 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4423) );
  AND2_X1 U5639 ( .A1(n6046), .A2(n6043), .ZN(n8711) );
  NAND2_X1 U5640 ( .A1(n5820), .A2(n5819), .ZN(n8257) );
  NAND2_X1 U5641 ( .A1(n5829), .A2(n5828), .ZN(n8264) );
  NAND2_X1 U5642 ( .A1(n5916), .A2(n5915), .ZN(n8730) );
  NAND2_X1 U5643 ( .A1(n4590), .A2(n4589), .ZN(n4588) );
  INV_X1 U5644 ( .A(n6112), .ZN(n4589) );
  NAND2_X1 U5645 ( .A1(n9109), .A2(n8834), .ZN(n4590) );
  AND2_X1 U5646 ( .A1(n5600), .A2(n5591), .ZN(n7106) );
  MUX2_X1 U5647 ( .A(n5599), .B(n6032), .S(n7467), .Z(n7107) );
  NAND2_X1 U5648 ( .A1(n4607), .A2(n4608), .ZN(n8751) );
  NAND2_X1 U5649 ( .A1(n4607), .A2(n4605), .ZN(n8753) );
  OAI211_X1 U5650 ( .C1(n6807), .C2(n5685), .A(n5660), .B(n5659), .ZN(n10022)
         );
  OAI21_X1 U5651 ( .B1(n5820), .B2(n4596), .A(n4593), .ZN(n8312) );
  AND2_X1 U5652 ( .A1(n4594), .A2(n5882), .ZN(n4593) );
  NAND2_X1 U5653 ( .A1(n4595), .A2(n4599), .ZN(n4594) );
  OAI21_X1 U5654 ( .B1(n8722), .B2(n8720), .A(n8719), .ZN(n5984) );
  OR2_X1 U5655 ( .A1(n5629), .A2(n5628), .ZN(n4578) );
  INV_X1 U5656 ( .A(n7224), .ZN(n4577) );
  NAND2_X1 U5657 ( .A1(n7548), .A2(n10047), .ZN(n7461) );
  OAI21_X1 U5658 ( .B1(n5916), .B2(n4586), .A(n4583), .ZN(n8739) );
  NAND2_X1 U5659 ( .A1(n7476), .A2(n7477), .ZN(n7475) );
  OAI21_X1 U5660 ( .B1(n8773), .B2(n4604), .A(n4601), .ZN(n8816) );
  AOI21_X1 U5661 ( .B1(n4605), .B2(n4603), .A(n4602), .ZN(n4601) );
  INV_X1 U5662 ( .A(n4605), .ZN(n4604) );
  INV_X1 U5663 ( .A(n6012), .ZN(n4602) );
  AND2_X1 U5664 ( .A1(n6107), .A2(n6091), .ZN(n10002) );
  NOR2_X1 U5665 ( .A1(n8800), .A2(n9053), .ZN(n8821) );
  INV_X1 U5666 ( .A(n8699), .ZN(n8860) );
  OR2_X1 U5667 ( .A1(n6175), .A2(n5601), .ZN(n5603) );
  OR2_X1 U5668 ( .A1(n6018), .A2(n8705), .ZN(n5602) );
  OR2_X1 U5669 ( .A1(n5956), .A2(n7032), .ZN(n5561) );
  OR2_X1 U5670 ( .A1(n6018), .A2(n7111), .ZN(n5560) );
  OR2_X1 U5671 ( .A1(n6173), .A2(n10108), .ZN(n5562) );
  INV_X1 U5672 ( .A(n7548), .ZN(n8863) );
  INV_X2 U5673 ( .A(P2_U3966), .ZN(n8862) );
  NOR2_X1 U5674 ( .A1(n7078), .A2(n7077), .ZN(n7076) );
  INV_X1 U5675 ( .A(n4481), .ZN(n7088) );
  NAND2_X1 U5676 ( .A1(n7091), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4480) );
  INV_X1 U5677 ( .A(n4487), .ZN(n7147) );
  OR2_X1 U5678 ( .A1(n8872), .A2(n8871), .ZN(n8873) );
  INV_X1 U5679 ( .A(n10011), .ZN(n10007) );
  AND2_X1 U5680 ( .A1(n8873), .A2(n4490), .ZN(n7267) );
  NAND2_X1 U5681 ( .A1(n7268), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4490) );
  NAND2_X1 U5682 ( .A1(n7267), .A2(n7266), .ZN(n7531) );
  INV_X1 U5683 ( .A(n9714), .ZN(n10013) );
  NOR2_X1 U5684 ( .A1(n8267), .A2(n4485), .ZN(n8270) );
  AND2_X1 U5685 ( .A1(n8271), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4485) );
  INV_X1 U5686 ( .A(n4484), .ZN(n8884) );
  INV_X1 U5687 ( .A(n6193), .ZN(n9096) );
  NAND2_X1 U5688 ( .A1(n4657), .A2(n4662), .ZN(n8925) );
  NAND2_X1 U5689 ( .A1(n8951), .A2(n4664), .ZN(n4657) );
  NAND2_X1 U5690 ( .A1(n4761), .A2(n6343), .ZN(n8945) );
  INV_X1 U5691 ( .A(n9113), .ZN(n8943) );
  NAND2_X1 U5692 ( .A1(n4665), .A2(n4669), .ZN(n8937) );
  AND2_X1 U5693 ( .A1(n5576), .A2(n5575), .ZN(n8974) );
  NAND2_X1 U5694 ( .A1(n9020), .A2(n6331), .ZN(n9001) );
  NAND2_X1 U5695 ( .A1(n4639), .A2(n4640), .ZN(n9005) );
  NAND2_X1 U5696 ( .A1(n4643), .A2(n4644), .ZN(n9019) );
  NAND2_X1 U5697 ( .A1(n9057), .A2(n4645), .ZN(n4643) );
  AND2_X1 U5698 ( .A1(n4646), .A2(n4649), .ZN(n9036) );
  NAND2_X1 U5699 ( .A1(n9057), .A2(n9056), .ZN(n4646) );
  NAND2_X1 U5700 ( .A1(n4626), .A2(n4624), .ZN(n8298) );
  AND2_X1 U5701 ( .A1(n4626), .A2(n4629), .ZN(n8291) );
  NAND2_X1 U5702 ( .A1(n8224), .A2(n4628), .ZN(n4626) );
  AND2_X1 U5703 ( .A1(n8224), .A2(n8223), .ZN(n8289) );
  NAND2_X1 U5704 ( .A1(n5851), .A2(n5850), .ZN(n9172) );
  NAND2_X1 U5705 ( .A1(n4739), .A2(n6134), .ZN(n8059) );
  NAND2_X1 U5706 ( .A1(n4632), .A2(n4633), .ZN(n8157) );
  INV_X1 U5707 ( .A(n8916), .ZN(n9043) );
  INV_X1 U5708 ( .A(n4617), .ZN(n7879) );
  NAND2_X1 U5709 ( .A1(n4616), .A2(n5715), .ZN(n7851) );
  NAND2_X1 U5710 ( .A1(n6823), .A2(n6188), .ZN(n4616) );
  NAND2_X1 U5711 ( .A1(n7629), .A2(n6124), .ZN(n7792) );
  INV_X1 U5712 ( .A(n6116), .ZN(n10058) );
  OR2_X1 U5713 ( .A1(n10035), .A2(n7538), .ZN(n10025) );
  INV_X1 U5714 ( .A(n9094), .ZN(n9006) );
  INV_X1 U5715 ( .A(n9063), .ZN(n9092) );
  AND2_X2 U5716 ( .A1(n7574), .A2(n7544), .ZN(n10119) );
  AND2_X1 U5717 ( .A1(n9104), .A2(n9103), .ZN(n9105) );
  AND2_X2 U5718 ( .A1(n7574), .A2(n7573), .ZN(n10105) );
  AND2_X1 U5719 ( .A1(n6376), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10045) );
  INV_X1 U5720 ( .A(n10039), .ZN(n10042) );
  NOR2_X1 U5721 ( .A1(n4764), .A2(n4765), .ZN(n4762) );
  NAND2_X1 U5722 ( .A1(n4476), .A2(n5551), .ZN(n4764) );
  NAND2_X1 U5724 ( .A1(n4477), .A2(n4475), .ZN(n5579) );
  NAND2_X1 U5725 ( .A1(n4476), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4475) );
  NAND2_X1 U5726 ( .A1(n6063), .A2(n4328), .ZN(n8222) );
  INV_X1 U5727 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7849) );
  XNOR2_X1 U5728 ( .A(n5566), .B(n5565), .ZN(n7847) );
  NAND2_X1 U5729 ( .A1(n6068), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5566) );
  INV_X1 U5730 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7819) );
  INV_X1 U5731 ( .A(n6226), .ZN(n7820) );
  INV_X1 U5732 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7744) );
  INV_X1 U5733 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7662) );
  INV_X1 U5734 ( .A(n8974), .ZN(n10027) );
  INV_X1 U5735 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7341) );
  INV_X1 U5736 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7259) );
  INV_X1 U5737 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7158) );
  INV_X1 U5738 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7113) );
  INV_X1 U5739 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7000) );
  INV_X1 U5740 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6889) );
  INV_X1 U5741 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6875) );
  INV_X1 U5742 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6827) );
  INV_X1 U5743 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6798) );
  OAI21_X1 U5744 ( .B1(n7191), .B2(n4694), .A(n4693), .ZN(n7301) );
  AOI21_X1 U5745 ( .B1(n4697), .B2(n6564), .A(n4696), .ZN(n4693) );
  INV_X1 U5746 ( .A(n4316), .ZN(n4697) );
  AND2_X1 U5747 ( .A1(n9291), .A2(n9294), .ZN(n4713) );
  NAND2_X1 U5748 ( .A1(n9303), .A2(n9306), .ZN(n4690) );
  AND2_X1 U5749 ( .A1(n8332), .A2(n9322), .ZN(n4386) );
  OR2_X1 U5750 ( .A1(n6534), .A2(n6533), .ZN(n6535) );
  NAND2_X1 U5751 ( .A1(n9284), .A2(n6697), .ZN(n9243) );
  NAND2_X1 U5752 ( .A1(n8102), .A2(n8106), .ZN(n8173) );
  INV_X1 U5753 ( .A(n9925), .ZN(n7386) );
  NAND2_X1 U5754 ( .A1(n4679), .A2(n4373), .ZN(n4387) );
  NAND2_X1 U5755 ( .A1(n4707), .A2(n4712), .ZN(n4705) );
  AND2_X1 U5756 ( .A1(n4369), .A2(n4709), .ZN(n9272) );
  OR2_X1 U5757 ( .A1(n9294), .A2(n4712), .ZN(n4710) );
  OR2_X1 U5758 ( .A1(n9291), .A2(n4712), .ZN(n4711) );
  NAND2_X1 U5759 ( .A1(n6590), .A2(n6589), .ZN(n7680) );
  NAND2_X1 U5760 ( .A1(n5192), .A2(n5191), .ZN(n7698) );
  AND2_X1 U5761 ( .A1(n5353), .A2(n5352), .ZN(n9538) );
  AND4_X1 U5762 ( .A1(n5249), .A2(n5248), .A3(n5247), .A4(n5246), .ZN(n7772)
         );
  NAND2_X1 U5763 ( .A1(n6761), .A2(n6756), .ZN(n9325) );
  NAND2_X1 U5764 ( .A1(n8105), .A2(n8104), .ZN(n8102) );
  NAND2_X1 U5765 ( .A1(n6655), .A2(n6654), .ZN(n8106) );
  NAND2_X1 U5766 ( .A1(n6896), .A2(n6755), .ZN(n9329) );
  INV_X1 U5767 ( .A(n7772), .ZN(n9348) );
  NAND2_X1 U5768 ( .A1(n5085), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5073) );
  AND2_X1 U5769 ( .A1(n5137), .A2(n5136), .ZN(n9819) );
  OR2_X1 U5770 ( .A1(n9829), .A2(n9828), .ZN(n9831) );
  NOR2_X1 U5771 ( .A1(n6927), .A2(n9875), .ZN(n6929) );
  INV_X1 U5772 ( .A(n4419), .ZN(n6981) );
  AOI21_X1 U5773 ( .B1(n9789), .B2(n7162), .A(n7161), .ZN(n7164) );
  XNOR2_X1 U5774 ( .A(n9371), .B(n7618), .ZN(n7613) );
  NAND2_X1 U5775 ( .A1(n9901), .A2(n4382), .ZN(n9918) );
  AOI21_X1 U5776 ( .B1(n9392), .B2(n9391), .A(n9390), .ZN(n9393) );
  XNOR2_X1 U5777 ( .A(n4414), .B(n4413), .ZN(n9398) );
  INV_X1 U5778 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n4413) );
  OR2_X1 U5779 ( .A1(n9388), .A2(n4415), .ZN(n4414) );
  AND2_X1 U5780 ( .A1(n9389), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4415) );
  NAND2_X1 U5781 ( .A1(n8343), .A2(n8342), .ZN(n9583) );
  INV_X1 U5782 ( .A(n9410), .ZN(n9590) );
  NAND2_X1 U5783 ( .A1(n4559), .A2(n4558), .ZN(n9440) );
  NAND2_X1 U5784 ( .A1(n9488), .A2(n8412), .ZN(n9474) );
  INV_X1 U5785 ( .A(n6713), .ZN(n9624) );
  AND2_X1 U5786 ( .A1(n5358), .A2(n5357), .ZN(n9512) );
  OR2_X1 U5787 ( .A1(n5339), .A2(n4858), .ZN(n4853) );
  NAND2_X1 U5788 ( .A1(n4856), .A2(n4872), .ZN(n9516) );
  OR2_X1 U5789 ( .A1(n5339), .A2(n5338), .ZN(n4856) );
  INV_X1 U5790 ( .A(n5339), .ZN(n9530) );
  OAI21_X1 U5791 ( .B1(n4832), .B2(n4834), .A(n4830), .ZN(n9546) );
  NAND2_X1 U5792 ( .A1(n4835), .A2(n4833), .ZN(n8201) );
  AND2_X1 U5793 ( .A1(n8129), .A2(n5296), .ZN(n9562) );
  AND2_X1 U5794 ( .A1(n9945), .A2(n5534), .ZN(n9940) );
  NAND2_X1 U5795 ( .A1(n7504), .A2(n9949), .ZN(n9945) );
  OAI21_X1 U5796 ( .B1(n9593), .B2(n9672), .A(n4394), .ZN(n9676) );
  NOR2_X1 U5797 ( .A1(n4540), .A2(n9975), .ZN(n4395) );
  NAND2_X1 U5798 ( .A1(n4354), .A2(n4539), .ZN(n4538) );
  INV_X1 U5799 ( .A(n9957), .ZN(n9958) );
  NOR2_X1 U5800 ( .A1(n8653), .A2(P1_U3084), .ZN(n9951) );
  AND2_X1 U5801 ( .A1(n4865), .A2(n4392), .ZN(n4391) );
  AND2_X1 U5802 ( .A1(n5004), .A2(n5015), .ZN(n4392) );
  INV_X1 U5803 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5015) );
  INV_X1 U5804 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7846) );
  INV_X1 U5805 ( .A(n6516), .ZN(n8555) );
  INV_X1 U5806 ( .A(n8640), .ZN(n8602) );
  INV_X1 U5807 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7804) );
  INV_X1 U5808 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7663) );
  INV_X1 U5809 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7342) );
  INV_X1 U5810 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7159) );
  INV_X1 U5811 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n7128) );
  INV_X1 U5812 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7001) );
  INV_X1 U5813 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6887) );
  INV_X1 U5814 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6804) );
  NAND2_X1 U5815 ( .A1(n4620), .A2(n4906), .ZN(n5151) );
  NAND2_X1 U5816 ( .A1(n5138), .A2(n5139), .ZN(n4620) );
  INV_X1 U5817 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6806) );
  NOR2_X1 U5818 ( .A1(n7932), .A2(n10159), .ZN(n10148) );
  AOI21_X1 U5819 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10146), .ZN(n10145) );
  NOR2_X1 U5820 ( .A1(n10145), .A2(n10144), .ZN(n10143) );
  INV_X1 U5821 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8910) );
  NAND2_X1 U5822 ( .A1(n7233), .A2(n5617), .ZN(n7225) );
  NOR2_X1 U5823 ( .A1(n9103), .A2(n9017), .ZN(n8693) );
  AOI21_X1 U5824 ( .B1(n4720), .B2(n6745), .A(n4716), .ZN(n4715) );
  INV_X1 U5825 ( .A(n4720), .ZN(n4719) );
  NAND2_X1 U5826 ( .A1(n4410), .A2(n8660), .ZN(P1_U3240) );
  AOI211_X1 U5827 ( .C1(n9759), .C2(n9424), .A(n9423), .B(n9422), .ZN(n9430)
         );
  NAND2_X1 U5828 ( .A1(n4565), .A2(n4564), .ZN(P1_U3520) );
  NAND2_X1 U5829 ( .A1(n9981), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n4564) );
  NAND2_X1 U5830 ( .A1(n9676), .A2(n9983), .ZN(n4565) );
  INV_X1 U5831 ( .A(n6519), .ZN(n6524) );
  AND4_X1 U5832 ( .A1(n5564), .A2(n5549), .A3(n5548), .A4(n6069), .ZN(n4314)
         );
  NAND2_X1 U5833 ( .A1(n4763), .A2(n4762), .ZN(n5553) );
  NOR2_X1 U5834 ( .A1(n9021), .A2(n4642), .ZN(n4315) );
  INV_X1 U5835 ( .A(n4796), .ZN(n4790) );
  INV_X1 U5836 ( .A(n9607), .ZN(n4848) );
  NOR2_X1 U5837 ( .A1(n6565), .A2(n4698), .ZN(n4316) );
  AND2_X1 U5838 ( .A1(n4469), .A2(n4468), .ZN(n4317) );
  INV_X1 U5839 ( .A(n6744), .ZN(n4724) );
  OR2_X1 U5840 ( .A1(n4354), .A2(n9578), .ZN(n4318) );
  INV_X1 U5841 ( .A(n4858), .ZN(n4857) );
  NAND2_X1 U5842 ( .A1(n9515), .A2(n4859), .ZN(n4858) );
  OR2_X1 U5843 ( .A1(n9337), .A2(n8556), .ZN(n4319) );
  AND2_X1 U5844 ( .A1(n6151), .A2(n4758), .ZN(n4320) );
  NAND2_X1 U5845 ( .A1(n5903), .A2(n5902), .ZN(n9161) );
  AND2_X1 U5846 ( .A1(n9155), .A2(n8807), .ZN(n6314) );
  AND2_X1 U5847 ( .A1(n4317), .A2(n4467), .ZN(n4321) );
  AND2_X1 U5848 ( .A1(n6148), .A2(n4754), .ZN(n4322) );
  AND2_X1 U5849 ( .A1(n5557), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n4323) );
  NOR2_X1 U5850 ( .A1(n9612), .A2(n5395), .ZN(n5396) );
  OR2_X1 U5851 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n4324) );
  OR2_X1 U5852 ( .A1(n8170), .A2(n8171), .ZN(n4679) );
  AND2_X1 U5853 ( .A1(n4526), .A2(n4525), .ZN(n4325) );
  NAND2_X1 U5854 ( .A1(n4825), .A2(n9747), .ZN(n4326) );
  NAND2_X1 U5855 ( .A1(n5242), .A2(n5241), .ZN(n9761) );
  INV_X1 U5856 ( .A(n9761), .ZN(n4532) );
  INV_X1 U5857 ( .A(n5085), .ZN(n5526) );
  AND2_X1 U5858 ( .A1(n6312), .A2(n6315), .ZN(n4327) );
  OR2_X1 U5859 ( .A1(n4454), .A2(n4457), .ZN(n4328) );
  NAND2_X1 U5860 ( .A1(n4751), .A2(n4752), .ZN(n4329) );
  NAND2_X1 U5861 ( .A1(n5271), .A2(n5270), .ZN(n5294) );
  AND2_X1 U5862 ( .A1(n8349), .A2(n5518), .ZN(n8593) );
  AOI21_X1 U5863 ( .B1(n5278), .B2(n4950), .A(n4797), .ZN(n4796) );
  NAND2_X1 U5864 ( .A1(n8588), .A2(n8357), .ZN(n4834) );
  AND2_X1 U5865 ( .A1(n5483), .A2(n5485), .ZN(n5475) );
  AOI21_X1 U5866 ( .B1(n9209), .B2(n6188), .A(n4869), .ZN(n8682) );
  INV_X1 U5867 ( .A(n8682), .ZN(n9101) );
  AND2_X1 U5868 ( .A1(n7047), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4330) );
  AND2_X1 U5869 ( .A1(n9654), .A2(n9344), .ZN(n4331) );
  INV_X1 U5870 ( .A(n7415), .ZN(n4696) );
  NAND3_X1 U5871 ( .A1(n5083), .A2(n5082), .A3(n5081), .ZN(n5084) );
  INV_X1 U5872 ( .A(n5084), .ZN(n4393) );
  INV_X1 U5873 ( .A(n6315), .ZN(n4749) );
  INV_X1 U5874 ( .A(n6119), .ZN(n10062) );
  AND2_X1 U5875 ( .A1(n9146), .A2(n9069), .ZN(n4332) );
  AND2_X1 U5876 ( .A1(n4853), .A2(n4854), .ZN(n4333) );
  NAND4_X1 U5877 ( .A1(n5605), .A2(n5604), .A3(n5603), .A4(n5602), .ZN(n6115)
         );
  NAND4_X1 U5878 ( .A1(n5637), .A2(n5636), .A3(n5635), .A4(n5634), .ZN(n8859)
         );
  INV_X1 U5879 ( .A(n7855), .ZN(n4619) );
  INV_X1 U5880 ( .A(n9464), .ZN(n4839) );
  NAND2_X1 U5881 ( .A1(n5920), .A2(n5919), .ZN(n9155) );
  INV_X1 U5882 ( .A(n9155), .ZN(n4468) );
  NAND2_X1 U5883 ( .A1(n7226), .A2(n6116), .ZN(n7667) );
  INV_X1 U5884 ( .A(n7667), .ZN(n4738) );
  AND2_X1 U5885 ( .A1(n8344), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n4334) );
  XNOR2_X1 U5886 ( .A(n5464), .B(n8596), .ZN(n9593) );
  NAND2_X1 U5887 ( .A1(n9243), .A2(n9244), .ZN(n9242) );
  NAND2_X1 U5888 ( .A1(n6675), .A2(n6676), .ZN(n9303) );
  AND2_X1 U5889 ( .A1(n4481), .A2(n4480), .ZN(n4335) );
  INV_X1 U5890 ( .A(n9465), .ZN(n9337) );
  AND4_X1 U5891 ( .A1(n5412), .A2(n5411), .A3(n5410), .A4(n5409), .ZN(n9465)
         );
  AND2_X1 U5892 ( .A1(n7486), .A2(n5170), .ZN(n4336) );
  AND2_X1 U5893 ( .A1(n6295), .A2(n6305), .ZN(n4337) );
  NOR2_X1 U5894 ( .A1(n6044), .A2(n8709), .ZN(n4338) );
  INV_X1 U5895 ( .A(n9612), .ZN(n9463) );
  AND2_X1 U5896 ( .A1(n4867), .A2(n5485), .ZN(n4339) );
  AND2_X1 U5897 ( .A1(n4690), .A2(n9304), .ZN(n4340) );
  OR2_X1 U5898 ( .A1(n9473), .A2(n8413), .ZN(n4341) );
  NAND2_X1 U5899 ( .A1(n5888), .A2(n5887), .ZN(n9167) );
  OR2_X1 U5900 ( .A1(n9446), .A2(n8347), .ZN(n4342) );
  AND2_X1 U5901 ( .A1(n4839), .A2(n4560), .ZN(n4343) );
  INV_X1 U5902 ( .A(n4845), .ZN(n4844) );
  AND2_X1 U5903 ( .A1(n4846), .A2(n4847), .ZN(n4845) );
  INV_X1 U5904 ( .A(n4811), .ZN(n4810) );
  NOR2_X1 U5905 ( .A1(n5233), .A2(n4812), .ZN(n4811) );
  AOI21_X1 U5906 ( .B1(n4832), .B2(n4548), .A(n4551), .ZN(n4547) );
  AND2_X1 U5907 ( .A1(n6135), .A2(n6134), .ZN(n4344) );
  INV_X1 U5908 ( .A(n8924), .ZN(n8927) );
  NAND2_X1 U5909 ( .A1(n6150), .A2(n6152), .ZN(n8924) );
  NAND2_X1 U5910 ( .A1(n8626), .A2(n8537), .ZN(n9437) );
  NAND2_X1 U5911 ( .A1(n8541), .A2(n8542), .ZN(n9425) );
  AND2_X1 U5912 ( .A1(n9634), .A2(n9341), .ZN(n4345) );
  INV_X1 U5913 ( .A(n9097), .ZN(n8919) );
  OR2_X1 U5914 ( .A1(n6321), .A2(n6320), .ZN(n4346) );
  NAND2_X1 U5915 ( .A1(n8926), .A2(n6351), .ZN(n8944) );
  INV_X1 U5916 ( .A(n8944), .ZN(n4667) );
  AND2_X1 U5917 ( .A1(n9179), .A2(n8851), .ZN(n4347) );
  NAND2_X1 U5918 ( .A1(n5810), .A2(n5809), .ZN(n9179) );
  NAND2_X1 U5919 ( .A1(n5406), .A2(n5405), .ZN(n9607) );
  INV_X1 U5920 ( .A(n4599), .ZN(n4598) );
  NAND2_X1 U5921 ( .A1(n4600), .A2(n5819), .ZN(n4599) );
  NOR2_X1 U5922 ( .A1(n9167), .A2(n8847), .ZN(n4348) );
  INV_X1 U5923 ( .A(n4809), .ZN(n4808) );
  OAI21_X1 U5924 ( .B1(n5219), .B2(n4810), .A(n4935), .ZN(n4809) );
  AND2_X1 U5925 ( .A1(n9236), .A2(n4687), .ZN(n4349) );
  INV_X1 U5926 ( .A(n4508), .ZN(n4507) );
  OAI21_X1 U5927 ( .B1(n4510), .B2(n4509), .A(n4876), .ZN(n4508) );
  NOR2_X1 U5928 ( .A1(n9629), .A2(n9340), .ZN(n4350) );
  NOR2_X1 U5929 ( .A1(n6616), .A2(n7762), .ZN(n4351) );
  AND2_X1 U5930 ( .A1(n9431), .A2(n5518), .ZN(n4558) );
  INV_X1 U5931 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5477) );
  NOR2_X1 U5932 ( .A1(n9141), .A2(n8844), .ZN(n4352) );
  INV_X1 U5933 ( .A(n4885), .ZN(n4672) );
  INV_X1 U5934 ( .A(n5396), .ZN(n4849) );
  NAND2_X1 U5935 ( .A1(n5547), .A2(n4753), .ZN(n4353) );
  INV_X1 U5936 ( .A(n4757), .ZN(n4756) );
  OR2_X1 U5937 ( .A1(n8674), .A2(n6320), .ZN(n4757) );
  INV_X1 U5938 ( .A(n4596), .ZN(n4595) );
  OR2_X1 U5939 ( .A1(n5883), .A2(n4597), .ZN(n4596) );
  INV_X1 U5940 ( .A(n8593), .ZN(n9448) );
  AND2_X1 U5941 ( .A1(n4823), .A2(n5533), .ZN(n4354) );
  INV_X1 U5942 ( .A(n4834), .ZN(n4833) );
  AND2_X1 U5943 ( .A1(n4908), .A2(SI_6_), .ZN(n4355) );
  INV_X1 U5944 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n4476) );
  OR2_X1 U5945 ( .A1(n4332), .A2(n4647), .ZN(n4356) );
  INV_X1 U5946 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6797) );
  INV_X1 U5947 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5004) );
  OR2_X1 U5948 ( .A1(n7855), .A2(n6254), .ZN(n4357) );
  AND2_X1 U5949 ( .A1(n5519), .A2(n8539), .ZN(n4358) );
  AND2_X1 U5950 ( .A1(n4640), .A2(n8674), .ZN(n4359) );
  OR2_X1 U5951 ( .A1(n6317), .A2(n6313), .ZN(n4360) );
  AND3_X1 U5952 ( .A1(n4874), .A2(n4456), .A3(n4766), .ZN(n4361) );
  AND2_X1 U5953 ( .A1(n4459), .A2(n7997), .ZN(n4362) );
  AND2_X1 U5954 ( .A1(n5354), .A2(n9518), .ZN(n4363) );
  OR2_X1 U5955 ( .A1(n8648), .A2(n8647), .ZN(n4364) );
  OR2_X1 U5956 ( .A1(n9512), .A2(n9522), .ZN(n4365) );
  INV_X1 U5957 ( .A(n7748), .ZN(n4737) );
  AOI22_X1 U5958 ( .A1(n6222), .A2(n8974), .B1(n6221), .B2(n6220), .ZN(n6373)
         );
  AND2_X1 U5959 ( .A1(n4679), .A2(n8104), .ZN(n4366) );
  NOR2_X1 U5960 ( .A1(n4792), .A2(n4959), .ZN(n4791) );
  OR2_X1 U5961 ( .A1(n4707), .A2(n4706), .ZN(n4367) );
  AND2_X1 U5962 ( .A1(n4679), .A2(n6654), .ZN(n4368) );
  NAND2_X1 U5963 ( .A1(n4704), .A2(n9291), .ZN(n4369) );
  OR2_X1 U5964 ( .A1(n4842), .A2(n4849), .ZN(n4370) );
  AND2_X1 U5965 ( .A1(n4408), .A2(n8498), .ZN(n4371) );
  INV_X1 U5966 ( .A(n4760), .ZN(n4759) );
  NAND2_X1 U5967 ( .A1(n4667), .A2(n6343), .ZN(n4760) );
  INV_X1 U5968 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4766) );
  NAND2_X1 U5969 ( .A1(n4384), .A2(n4383), .ZN(n7678) );
  INV_X1 U5970 ( .A(n6745), .ZN(n4726) );
  NAND2_X1 U5971 ( .A1(n5844), .A2(n5547), .ZN(n5847) );
  AND2_X1 U5972 ( .A1(n7121), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4372) );
  NAND2_X1 U5973 ( .A1(n4579), .A2(n8036), .ZN(n8047) );
  AND2_X1 U5974 ( .A1(n8170), .A2(n8171), .ZN(n4373) );
  NOR2_X1 U5975 ( .A1(n5686), .A2(n5546), .ZN(n5844) );
  NAND2_X1 U5976 ( .A1(n4740), .A2(n6305), .ZN(n8226) );
  INV_X1 U5977 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5235) );
  INV_X1 U5978 ( .A(n9109), .ZN(n4474) );
  OR2_X1 U5979 ( .A1(n5294), .A2(n9570), .ZN(n8481) );
  AND2_X1 U5980 ( .A1(n9518), .A2(n8501), .ZN(n9536) );
  INV_X1 U5981 ( .A(n9536), .ZN(n4550) );
  NAND2_X1 U5982 ( .A1(n5421), .A2(n5420), .ZN(n9601) );
  NAND2_X1 U5983 ( .A1(n9563), .A2(n4528), .ZN(n4529) );
  AND2_X1 U5984 ( .A1(n6735), .A2(n6734), .ZN(n6745) );
  INV_X1 U5985 ( .A(n9596), .ZN(n9415) );
  NAND2_X1 U5986 ( .A1(n5440), .A2(n5439), .ZN(n9596) );
  AND2_X1 U5987 ( .A1(n7969), .A2(n8472), .ZN(n4374) );
  AND2_X1 U5988 ( .A1(n6763), .A2(n6764), .ZN(n4375) );
  AND2_X1 U5989 ( .A1(n4958), .A2(SI_17_), .ZN(n4376) );
  NAND2_X1 U5990 ( .A1(n4567), .A2(n4566), .ZN(n4570) );
  AND2_X1 U5991 ( .A1(n9109), .A2(n10002), .ZN(n4377) );
  INV_X1 U5992 ( .A(n4649), .ZN(n4647) );
  NAND2_X1 U5993 ( .A1(n9149), .A2(n8845), .ZN(n4649) );
  NAND2_X1 U5994 ( .A1(n4402), .A2(n8377), .ZN(n7203) );
  NAND2_X1 U5995 ( .A1(n5266), .A2(n5265), .ZN(n7904) );
  INV_X1 U5996 ( .A(n7904), .ZN(n4535) );
  NAND2_X1 U5997 ( .A1(n5933), .A2(n5932), .ZN(n9149) );
  INV_X1 U5998 ( .A(n9149), .ZN(n4467) );
  AND2_X1 U5999 ( .A1(n7191), .A2(n6556), .ZN(n4378) );
  NAND2_X1 U6000 ( .A1(n7889), .A2(n4459), .ZN(n4379) );
  NAND2_X1 U6001 ( .A1(n5343), .A2(n5342), .ZN(n9634) );
  INV_X1 U6002 ( .A(n9634), .ZN(n4525) );
  INV_X1 U6003 ( .A(n7604), .ZN(n4533) );
  AND2_X1 U6004 ( .A1(n6187), .A2(SI_30_), .ZN(n4380) );
  NAND2_X1 U6005 ( .A1(n6579), .A2(n6580), .ZN(n7424) );
  NAND2_X1 U6006 ( .A1(n7475), .A2(n5683), .ZN(n7513) );
  AND2_X1 U6007 ( .A1(n6110), .A2(n6097), .ZN(n8834) );
  AND2_X1 U6008 ( .A1(n8344), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n4381) );
  NAND2_X1 U6009 ( .A1(n7349), .A2(n5128), .ZN(n7283) );
  NAND2_X1 U6010 ( .A1(n7395), .A2(n4336), .ZN(n7483) );
  NAND2_X1 U6011 ( .A1(n6123), .A2(n6122), .ZN(n7629) );
  NAND2_X1 U6012 ( .A1(n5541), .A2(n4874), .ZN(n5686) );
  INV_X1 U6013 ( .A(n4629), .ZN(n4627) );
  NAND2_X1 U6014 ( .A1(n9172), .A2(n8848), .ZN(n4629) );
  AND2_X1 U6015 ( .A1(n9224), .A2(n6543), .ZN(n7003) );
  AND2_X1 U6016 ( .A1(n7025), .A2(n7806), .ZN(n9764) );
  NAND2_X1 U6017 ( .A1(n5211), .A2(n5210), .ZN(n7707) );
  INV_X1 U6018 ( .A(n7707), .ZN(n4531) );
  NAND2_X1 U6019 ( .A1(n7020), .A2(n7018), .ZN(n7019) );
  OR2_X1 U6020 ( .A1(n6542), .A2(n6541), .ZN(n9224) );
  NAND2_X1 U6021 ( .A1(n7349), .A2(n4862), .ZN(n7282) );
  OR2_X1 U6022 ( .A1(n9364), .A2(n9363), .ZN(n4382) );
  INV_X1 U6023 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n4615) );
  INV_X1 U6024 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n4818) );
  AOI21_X2 U6025 ( .B1(n8004), .B2(n5454), .A(n4381), .ZN(n8350) );
  INV_X1 U6026 ( .A(n8524), .ZN(n8527) );
  NAND2_X1 U6027 ( .A1(n4412), .A2(n4411), .ZN(n4410) );
  OAI21_X1 U6028 ( .B1(n8540), .B2(n4397), .A(n4396), .ZN(n8544) );
  INV_X4 U6029 ( .A(n5011), .ZN(n5400) );
  OAI21_X1 U6030 ( .B1(n5341), .B2(n4815), .A(n4976), .ZN(n5356) );
  OAI22_X1 U6031 ( .A1(n8553), .A2(n8554), .B1(n8552), .B2(n8551), .ZN(n8563)
         );
  INV_X4 U6032 ( .A(n6528), .ZN(n8329) );
  INV_X1 U6033 ( .A(n7680), .ZN(n4384) );
  NOR2_X1 U6034 ( .A1(n9253), .A2(n9252), .ZN(n9251) );
  NOR2_X1 U6035 ( .A1(n9317), .A2(n4725), .ZN(n8341) );
  NAND2_X1 U6036 ( .A1(n9235), .A2(n9280), .ZN(n6696) );
  NAND2_X1 U6037 ( .A1(n6655), .A2(n4368), .ZN(n4677) );
  NAND2_X1 U6038 ( .A1(n5475), .A2(n5477), .ZN(n4676) );
  OAI21_X1 U6039 ( .B1(n7835), .B2(n7832), .A(n7831), .ZN(n6650) );
  NAND3_X2 U6040 ( .A1(n8093), .A2(n6653), .A3(n8090), .ZN(n8105) );
  OAI211_X1 U6041 ( .C1(n8341), .C2(n8340), .A(n4385), .B(n8339), .ZN(P1_U3218) );
  NAND2_X1 U6042 ( .A1(n8341), .A2(n4386), .ZN(n4385) );
  NAND3_X1 U6043 ( .A1(n4316), .A2(n7191), .A3(n7415), .ZN(n4692) );
  OAI21_X2 U6044 ( .B1(n8684), .B2(n6350), .A(n6202), .ZN(n6179) );
  AOI21_X1 U6045 ( .B1(n6194), .B2(n6217), .A(n6364), .ZN(n6195) );
  NAND4_X1 U6046 ( .A1(n6375), .A2(n4435), .A3(n4499), .A4(n6373), .ZN(n4434)
         );
  NAND2_X1 U6047 ( .A1(n4514), .A2(n4512), .ZN(n5164) );
  NAND2_X1 U6048 ( .A1(n4788), .A2(n4789), .ZN(n5314) );
  NAND2_X1 U6049 ( .A1(n5367), .A2(n5366), .ZN(n5369) );
  OAI211_X1 U6050 ( .C1(n4435), .C2(n4498), .A(n4434), .B(n7952), .ZN(n4433)
         );
  NAND2_X1 U6051 ( .A1(n4433), .A2(n6381), .ZN(n6515) );
  NAND2_X1 U6052 ( .A1(n4778), .A2(n4783), .ZN(n5414) );
  OAI21_X1 U6053 ( .B1(n5356), .B2(n5355), .A(n4981), .ZN(n5367) );
  NAND2_X1 U6054 ( .A1(n4973), .A2(n4972), .ZN(n5341) );
  NAND2_X1 U6055 ( .A1(n7424), .A2(n6586), .ZN(n6590) );
  NAND2_X1 U6056 ( .A1(n6534), .A2(n6533), .ZN(n7004) );
  NAND2_X2 U6057 ( .A1(n7192), .A2(n7193), .ZN(n7191) );
  NAND2_X1 U6058 ( .A1(n6631), .A2(n6630), .ZN(n7835) );
  NAND2_X1 U6059 ( .A1(n4695), .A2(n6564), .ZN(n6574) );
  NAND3_X1 U6060 ( .A1(n4678), .A2(n4677), .A3(n4387), .ZN(n9260) );
  NAND2_X2 U6061 ( .A1(n9293), .A2(n9292), .ZN(n9291) );
  NOR2_X2 U6062 ( .A1(n5365), .A2(n5364), .ZN(n9472) );
  OAI21_X2 U6063 ( .B1(n9545), .B2(n5324), .A(n4390), .ZN(n5339) );
  NAND3_X1 U6064 ( .A1(n7282), .A2(n5142), .A3(n5155), .ZN(n7433) );
  NAND2_X1 U6065 ( .A1(n4391), .A2(n5483), .ZN(n5018) );
  AND3_X1 U6066 ( .A1(n5483), .A2(n5004), .A3(n4865), .ZN(n5016) );
  NAND2_X1 U6067 ( .A1(n5483), .A2(n4865), .ZN(n5003) );
  NAND4_X1 U6068 ( .A1(n5071), .A2(n5073), .A3(n5072), .A4(n5074), .ZN(n6529)
         );
  NOR2_X2 U6069 ( .A1(n4538), .A2(n4395), .ZN(n4394) );
  NAND2_X1 U6070 ( .A1(n4401), .A2(n4402), .ZN(n7345) );
  NAND2_X1 U6071 ( .A1(n8380), .A2(n5508), .ZN(n4402) );
  NAND3_X1 U6072 ( .A1(n8496), .A2(n8497), .A3(n4371), .ZN(n4407) );
  OR2_X1 U6073 ( .A1(n8493), .A2(n4409), .ZN(n4408) );
  NAND3_X1 U6074 ( .A1(n8646), .A2(n8647), .A3(n8645), .ZN(n4412) );
  NAND2_X1 U6075 ( .A1(n7022), .A2(n7023), .ZN(n7021) );
  XNOR2_X1 U6076 ( .A(n5075), .B(n5076), .ZN(n6809) );
  XNOR2_X1 U6077 ( .A(n4890), .B(n4889), .ZN(n5075) );
  MUX2_X1 U6078 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n7219), .S(n6849), .Z(n6877)
         );
  NAND2_X1 U6079 ( .A1(n4430), .A2(n4426), .ZN(n6284) );
  OAI21_X1 U6080 ( .B1(n4429), .B2(n4428), .A(n4427), .ZN(n4426) );
  NOR2_X1 U6081 ( .A1(n6272), .A2(n6268), .ZN(n4429) );
  NAND2_X1 U6082 ( .A1(n6277), .A2(n4453), .ZN(n4430) );
  NAND3_X1 U6083 ( .A1(n4731), .A2(n4730), .A3(n4458), .ZN(n5655) );
  NAND4_X1 U6085 ( .A1(n4314), .A2(n5541), .A3(n4874), .A4(n4456), .ZN(n4455)
         );
  NAND3_X1 U6086 ( .A1(n4314), .A2(n5541), .A3(n4361), .ZN(n4454) );
  OR2_X2 U6087 ( .A1(n4455), .A2(n4457), .ZN(n6061) );
  INV_X1 U6088 ( .A(n4752), .ZN(n4457) );
  NAND2_X2 U6089 ( .A1(n8687), .A2(n8663), .ZN(n5707) );
  INV_X1 U6090 ( .A(n5655), .ZN(n5541) );
  NAND4_X1 U6091 ( .A1(n8702), .A2(n4463), .A3(n7801), .A4(n4462), .ZN(n7725)
         );
  NAND2_X1 U6092 ( .A1(n8957), .A2(n4470), .ZN(n8917) );
  NAND2_X1 U6093 ( .A1(n8957), .A2(n8943), .ZN(n8938) );
  NOR2_X1 U6094 ( .A1(n8938), .A2(n4473), .ZN(n8918) );
  MUX2_X1 U6095 ( .A(n7032), .B(P2_REG2_REG_1__SCAN_IN), .S(n7033), .Z(n9712)
         );
  NAND2_X1 U6096 ( .A1(n6329), .A2(n4491), .ZN(n6319) );
  OAI21_X1 U6097 ( .B1(n6316), .B2(n4360), .A(n9064), .ZN(n4494) );
  NAND2_X1 U6098 ( .A1(n4496), .A2(n6372), .ZN(n4495) );
  NAND3_X1 U6099 ( .A1(n4497), .A2(n6328), .A3(n9064), .ZN(n4496) );
  OAI21_X1 U6100 ( .B1(n6316), .B2(n4749), .A(n6141), .ZN(n4497) );
  NAND3_X1 U6101 ( .A1(n4499), .A2(n6375), .A3(n4500), .ZN(n4498) );
  OR2_X1 U6102 ( .A1(n6373), .A2(n7745), .ZN(n4499) );
  INV_X1 U6103 ( .A(n4816), .ZN(n4503) );
  NAND2_X1 U6104 ( .A1(n4816), .A2(n4911), .ZN(n5172) );
  INV_X1 U6105 ( .A(n4917), .ZN(n4509) );
  AND2_X1 U6106 ( .A1(n4511), .A2(n4911), .ZN(n4510) );
  NAND3_X1 U6107 ( .A1(n5139), .A2(n5150), .A3(n5138), .ZN(n4514) );
  NAND2_X1 U6108 ( .A1(n4941), .A2(n4940), .ZN(n5046) );
  OAI21_X1 U6109 ( .B1(n4941), .B2(n4518), .A(n4516), .ZN(n4522) );
  NAND2_X2 U6110 ( .A1(n4886), .A2(n4885), .ZN(n5011) );
  NAND3_X1 U6111 ( .A1(n4310), .A2(n4885), .A3(n6806), .ZN(n4523) );
  INV_X1 U6112 ( .A(n4529), .ZN(n9552) );
  NOR2_X2 U6113 ( .A1(n4530), .A2(n5134), .ZN(n5483) );
  NAND2_X2 U6114 ( .A1(n5000), .A2(n4873), .ZN(n5134) );
  NAND4_X1 U6115 ( .A1(n4997), .A2(n4996), .A3(n5034), .A4(n4995), .ZN(n4530)
         );
  NOR2_X1 U6116 ( .A1(n7604), .A2(n7707), .ZN(n7737) );
  INV_X1 U6117 ( .A(n9447), .ZN(n4557) );
  NAND2_X1 U6118 ( .A1(n9488), .A2(n4562), .ZN(n4561) );
  XNOR2_X1 U6119 ( .A(n5138), .B(n5139), .ZN(n6807) );
  NAND3_X1 U6120 ( .A1(n4310), .A2(n4885), .A3(n4897), .ZN(n4574) );
  NAND2_X1 U6121 ( .A1(n4576), .A2(n4578), .ZN(n7312) );
  NAND3_X1 U6122 ( .A1(n7233), .A2(n5617), .A3(n4577), .ZN(n4576) );
  NAND2_X1 U6123 ( .A1(n7105), .A2(n5600), .ZN(n7234) );
  NAND3_X1 U6124 ( .A1(n4579), .A2(n8036), .A3(n5798), .ZN(n5804) );
  NAND2_X1 U6125 ( .A1(n4580), .A2(n4581), .ZN(n8742) );
  NAND2_X1 U6126 ( .A1(n5916), .A2(n4583), .ZN(n4580) );
  OAI21_X1 U6127 ( .B1(n6113), .B2(n9109), .A(n4587), .ZN(P2_U3222) );
  AOI21_X1 U6128 ( .B1(n6095), .B2(n4377), .A(n4588), .ZN(n4587) );
  NAND2_X1 U6129 ( .A1(n7475), .A2(n4591), .ZN(n5706) );
  NOR2_X1 U6130 ( .A1(n6061), .A2(n4610), .ZN(n5577) );
  NAND2_X2 U6131 ( .A1(n4613), .A2(n9207), .ZN(n6018) );
  NAND2_X2 U6132 ( .A1(n4613), .A2(n5557), .ZN(n6173) );
  INV_X1 U6133 ( .A(n6018), .ZN(n6099) );
  INV_X1 U6134 ( .A(n5686), .ZN(n4751) );
  NAND2_X1 U6135 ( .A1(n5576), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5572) );
  AND2_X4 U6136 ( .A1(n10046), .A2(n7745), .ZN(n9181) );
  OAI21_X1 U6137 ( .B1(n8224), .B2(n4623), .A(n4621), .ZN(n8670) );
  NAND2_X1 U6138 ( .A1(n8068), .A2(n4634), .ZN(n4632) );
  INV_X1 U6139 ( .A(n9057), .ZN(n4638) );
  NAND2_X1 U6140 ( .A1(n4638), .A2(n4315), .ZN(n4639) );
  OR2_X1 U6141 ( .A1(n8951), .A2(n8953), .ZN(n4665) );
  NAND3_X1 U6142 ( .A1(n4654), .A2(n4653), .A3(n4650), .ZN(n9106) );
  NAND3_X1 U6143 ( .A1(n8951), .A2(n4658), .A3(n8683), .ZN(n4653) );
  NAND3_X1 U6144 ( .A1(n4310), .A2(n4885), .A3(n6810), .ZN(n4670) );
  NAND2_X1 U6145 ( .A1(n6991), .A2(n4673), .ZN(n4674) );
  AND2_X1 U6146 ( .A1(n9224), .A2(n7004), .ZN(n4673) );
  NAND2_X1 U6147 ( .A1(n6991), .A2(n7004), .ZN(n7007) );
  INV_X1 U6148 ( .A(n9224), .ZN(n4675) );
  NAND2_X1 U6149 ( .A1(n8105), .A2(n4366), .ZN(n4678) );
  NAND2_X1 U6150 ( .A1(n6696), .A2(n4681), .ZN(n4680) );
  NAND2_X1 U6151 ( .A1(n4680), .A2(n4683), .ZN(n6709) );
  OAI21_X2 U6152 ( .B1(n6675), .B2(n4689), .A(n4349), .ZN(n9235) );
  NAND2_X1 U6153 ( .A1(n4692), .A2(n4691), .ZN(n6570) );
  NAND2_X1 U6154 ( .A1(n7191), .A2(n4316), .ZN(n4695) );
  NAND2_X1 U6155 ( .A1(n6765), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n4702) );
  NAND3_X1 U6156 ( .A1(n4701), .A2(n6518), .A3(n6519), .ZN(n4699) );
  OR2_X2 U6157 ( .A1(n8242), .A2(n4700), .ZN(n6518) );
  NAND2_X1 U6158 ( .A1(n4703), .A2(n4705), .ZN(n9270) );
  NAND3_X1 U6159 ( .A1(n9291), .A2(n4367), .A3(n9294), .ZN(n4703) );
  NAND3_X1 U6160 ( .A1(n4711), .A2(n4710), .A3(n9216), .ZN(n4709) );
  OR2_X1 U6161 ( .A1(n4713), .A2(n4712), .ZN(n9215) );
  INV_X1 U6162 ( .A(n6715), .ZN(n4712) );
  NAND2_X1 U6163 ( .A1(n9320), .A2(n4718), .ZN(n4714) );
  NOR2_X1 U6164 ( .A1(n9251), .A2(n4727), .ZN(n9317) );
  OAI211_X1 U6165 ( .C1(n9320), .C2(n4719), .A(n4714), .B(n4715), .ZN(P1_U3212) );
  NAND2_X1 U6166 ( .A1(n7666), .A2(n4735), .ZN(n4734) );
  NAND2_X1 U6167 ( .A1(n7675), .A2(n7748), .ZN(n4733) );
  NAND2_X1 U6168 ( .A1(n4734), .A2(n4732), .ZN(n7563) );
  NAND2_X1 U6169 ( .A1(n4736), .A2(n6231), .ZN(n7665) );
  NAND2_X1 U6170 ( .A1(n7666), .A2(n7667), .ZN(n4736) );
  NAND2_X1 U6171 ( .A1(n6123), .A2(n4743), .ZN(n4741) );
  NAND2_X1 U6172 ( .A1(n4741), .A2(n4742), .ZN(n7715) );
  NAND2_X1 U6173 ( .A1(n6140), .A2(n4747), .ZN(n4746) );
  NOR2_X2 U6174 ( .A1(n5546), .A2(n4353), .ZN(n4752) );
  OAI21_X1 U6175 ( .B1(n8952), .B2(n4760), .A(n4320), .ZN(n6153) );
  INV_X1 U6176 ( .A(n6061), .ZN(n4763) );
  NAND2_X1 U6177 ( .A1(n6163), .A2(n6182), .ZN(n6183) );
  NAND2_X1 U6178 ( .A1(n6163), .A2(n4770), .ZN(n4769) );
  NAND3_X1 U6179 ( .A1(n4771), .A2(n4768), .A3(n4767), .ZN(n6191) );
  NAND2_X1 U6180 ( .A1(n5383), .A2(n4779), .ZN(n4777) );
  OR2_X1 U6181 ( .A1(n5383), .A2(n5382), .ZN(n4787) );
  NAND2_X1 U6182 ( .A1(n5279), .A2(n4791), .ZN(n4788) );
  OAI21_X1 U6183 ( .B1(n5279), .B2(n4790), .A(n4793), .ZN(n5298) );
  NAND2_X1 U6184 ( .A1(n5447), .A2(n4802), .ZN(n4800) );
  NAND2_X1 U6185 ( .A1(n5447), .A2(n5446), .ZN(n4801) );
  NAND2_X1 U6186 ( .A1(n5075), .A2(n5076), .ZN(n4892) );
  OAI21_X1 U6187 ( .B1(n5011), .B2(n4818), .A(n4817), .ZN(n5076) );
  NAND2_X1 U6188 ( .A1(n5011), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4817) );
  NAND2_X1 U6189 ( .A1(n5122), .A2(n5123), .ZN(n4819) );
  NAND2_X1 U6190 ( .A1(n5108), .A2(n5109), .ZN(n4820) );
  NAND2_X1 U6191 ( .A1(n9416), .A2(n8539), .ZN(n9420) );
  NAND2_X1 U6192 ( .A1(n4824), .A2(n4822), .ZN(n4823) );
  AOI21_X1 U6193 ( .B1(n9416), .B2(n4358), .A(n4326), .ZN(n4822) );
  NAND3_X1 U6194 ( .A1(n4310), .A2(n4885), .A3(n4887), .ZN(n5094) );
  NOR2_X1 U6195 ( .A1(n9571), .A2(n5516), .ZN(n8202) );
  NAND2_X1 U6196 ( .A1(n5086), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5061) );
  AOI21_X1 U6197 ( .B1(n9460), .B2(n9464), .A(n5396), .ZN(n9445) );
  NAND2_X1 U6198 ( .A1(n4863), .A2(n4864), .ZN(n7966) );
  NAND2_X1 U6199 ( .A1(n9746), .A2(n5250), .ZN(n4863) );
  CLKBUF_X1 U6200 ( .A(n9235), .Z(n9279) );
  NOR2_X1 U6201 ( .A1(n5032), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5035) );
  AOI21_X2 U6202 ( .B1(n7678), .B2(n6617), .A(n4351), .ZN(n7768) );
  NAND2_X1 U6203 ( .A1(n6570), .A2(n7298), .ZN(n6580) );
  OR2_X2 U6204 ( .A1(n6650), .A2(n6649), .ZN(n8090) );
  OR2_X1 U6205 ( .A1(n8242), .A2(n5488), .ZN(n9950) );
  CLKBUF_X1 U6206 ( .A(n5506), .Z(n8640) );
  XNOR2_X1 U6207 ( .A(n6532), .B(n6551), .ZN(n6533) );
  INV_X1 U6208 ( .A(n6709), .ZN(n6712) );
  NAND2_X1 U6209 ( .A1(n6709), .A2(n6710), .ZN(n9293) );
  INV_X2 U6210 ( .A(n5684), .ZN(n6189) );
  OR2_X1 U6211 ( .A1(n5684), .A2(n6794), .ZN(n5611) );
  OR2_X1 U6212 ( .A1(n5577), .A2(n5554), .ZN(n5555) );
  NAND2_X1 U6213 ( .A1(n6139), .A2(n4327), .ZN(n6140) );
  XNOR2_X1 U6214 ( .A(n5472), .B(n5471), .ZN(n7806) );
  AND4_X2 U6215 ( .A1(n5133), .A2(n5132), .A3(n5131), .A4(n5130), .ZN(n7438)
         );
  NAND2_X1 U6216 ( .A1(n7130), .A2(n5099), .ZN(n7201) );
  INV_X1 U6217 ( .A(n5781), .ZN(n5784) );
  NAND2_X1 U6218 ( .A1(n5086), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5089) );
  INV_X1 U6219 ( .A(n5559), .ZN(n5557) );
  OR2_X1 U6220 ( .A1(n5016), .A2(n9695), .ZN(n5014) );
  NOR2_X1 U6221 ( .A1(n9270), .A2(n6721), .ZN(n9253) );
  NAND2_X1 U6222 ( .A1(n6263), .A2(n6262), .ZN(n7722) );
  INV_X1 U6223 ( .A(n7486), .ZN(n8575) );
  NAND2_X1 U6224 ( .A1(n8451), .A2(n8458), .ZN(n7486) );
  AND2_X2 U6225 ( .A1(n6973), .A2(n6914), .ZN(n9983) );
  AND2_X1 U6226 ( .A1(n6189), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n4869) );
  AND2_X1 U6227 ( .A1(n6747), .A2(n6951), .ZN(n9754) );
  AND2_X1 U6228 ( .A1(n5299), .A2(n5302), .ZN(n4871) );
  OR2_X1 U6229 ( .A1(n9535), .A2(n9549), .ZN(n4872) );
  INV_X1 U6230 ( .A(n7631), .ZN(n6122) );
  AND2_X1 U6231 ( .A1(n6762), .A2(n9949), .ZN(n9332) );
  NAND2_X1 U6232 ( .A1(n5521), .A2(n5520), .ZN(n9747) );
  AND2_X1 U6233 ( .A1(n4927), .A2(n4926), .ZN(n4875) );
  AND2_X1 U6234 ( .A1(n4923), .A2(n4922), .ZN(n4876) );
  AND4_X1 U6235 ( .A1(n5444), .A2(n5443), .A3(n5442), .A4(n5441), .ZN(n9438)
         );
  INV_X1 U6236 ( .A(n8846), .ZN(n8667) );
  OR2_X2 U6237 ( .A1(n9246), .A2(n5344), .ZN(n4877) );
  OR2_X1 U6238 ( .A1(n8350), .A2(n9491), .ZN(n4879) );
  INV_X1 U6239 ( .A(n9515), .ZN(n5354) );
  AND2_X1 U6240 ( .A1(n5625), .A2(n5624), .ZN(n4880) );
  NAND2_X1 U6241 ( .A1(n6254), .A2(n4453), .ZN(n6255) );
  NAND2_X1 U6242 ( .A1(n4619), .A2(n6255), .ZN(n6256) );
  AOI21_X1 U6243 ( .B1(n6258), .B2(n6257), .A(n6256), .ZN(n6267) );
  INV_X1 U6244 ( .A(n8288), .ZN(n6295) );
  NOR2_X1 U6245 ( .A1(n6350), .A2(n6349), .ZN(n6354) );
  AOI21_X1 U6246 ( .B1(n6367), .B2(n6363), .A(n6362), .ZN(n6365) );
  INV_X1 U6247 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5540) );
  OR2_X1 U6248 ( .A1(n5509), .A2(n8429), .ZN(n5510) );
  INV_X1 U6249 ( .A(n8156), .ZN(n6135) );
  NAND2_X1 U6250 ( .A1(n5084), .A2(n8329), .ZN(n6531) );
  AOI21_X1 U6251 ( .B1(n8428), .B2(n8373), .A(n8604), .ZN(n7400) );
  INV_X1 U6252 ( .A(n5066), .ZN(n5000) );
  AND2_X1 U6253 ( .A1(n8861), .A2(n6196), .ZN(n5590) );
  INV_X1 U6254 ( .A(n5782), .ZN(n5783) );
  INV_X1 U6255 ( .A(SI_10_), .ZN(n6484) );
  OR2_X1 U6256 ( .A1(n7185), .A2(n6197), .ZN(n6198) );
  INV_X1 U6257 ( .A(n5978), .ZN(n5976) );
  INV_X1 U6258 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8827) );
  INV_X1 U6259 ( .A(n5906), .ZN(n5904) );
  NAND2_X1 U6260 ( .A1(n8699), .A2(n6119), .ZN(n7748) );
  INV_X1 U6261 ( .A(n8327), .ZN(n6551) );
  INV_X1 U6262 ( .A(n6993), .ZN(n6538) );
  INV_X1 U6263 ( .A(n8571), .ZN(n5155) );
  OAI22_X1 U6264 ( .A1(n9438), .A2(n5531), .B1(n5530), .B2(n5529), .ZN(n5532)
         );
  NAND2_X1 U6265 ( .A1(n5431), .A2(n5430), .ZN(n5433) );
  INV_X1 U6266 ( .A(n5313), .ZN(n4960) );
  INV_X1 U6267 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5037) );
  NAND2_X1 U6268 ( .A1(n5202), .A2(n4875), .ZN(n4928) );
  INV_X1 U6269 ( .A(n6016), .ZN(n6015) );
  OR2_X1 U6270 ( .A1(n6049), .A2(n6048), .ZN(n6098) );
  NAND2_X1 U6271 ( .A1(n5976), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5988) );
  OR3_X1 U6272 ( .A1(n5831), .A2(n7655), .A3(n5830), .ZN(n5867) );
  OR2_X1 U6273 ( .A1(n5952), .A2(n8745), .ZN(n5960) );
  NAND2_X1 U6274 ( .A1(n5904), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5922) );
  INV_X1 U6275 ( .A(n7722), .ZN(n6126) );
  AND2_X1 U6276 ( .A1(n7564), .A2(n6245), .ZN(n6206) );
  INV_X1 U6277 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5143) );
  AND2_X2 U6278 ( .A1(n7806), .A2(n5506), .ZN(n7015) );
  AND2_X1 U6279 ( .A1(n8610), .A2(n8608), .ZN(n8571) );
  NAND2_X1 U6280 ( .A1(n5007), .A2(n5006), .ZN(n5522) );
  XNOR2_X1 U6281 ( .A(n4929), .B(SI_11_), .ZN(n5219) );
  INV_X1 U6282 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5718) );
  AND2_X1 U6283 ( .A1(n5881), .A2(n8759), .ZN(n5882) );
  NAND2_X1 U6284 ( .A1(n5735), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5775) );
  INV_X1 U6285 ( .A(n8821), .ZN(n9995) );
  INV_X1 U6286 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5667) );
  AND3_X1 U6287 ( .A1(n6178), .A2(n6177), .A3(n6176), .ZN(n6192) );
  AND2_X1 U6288 ( .A1(n6050), .A2(n6098), .ZN(n8932) );
  INV_X1 U6289 ( .A(n6173), .ZN(n5980) );
  INV_X1 U6290 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7655) );
  AND2_X1 U6291 ( .A1(n8274), .A2(n8273), .ZN(n8275) );
  AOI21_X1 U6292 ( .B1(n10034), .B2(n10043), .A(n10044), .ZN(n7541) );
  INV_X1 U6293 ( .A(n8957), .ZN(n8940) );
  INV_X1 U6294 ( .A(n8842), .ZN(n8968) );
  INV_X1 U6295 ( .A(n8843), .ZN(n9003) );
  INV_X1 U6296 ( .A(n6314), .ZN(n9064) );
  INV_X1 U6297 ( .A(n8847), .ZN(n8766) );
  INV_X1 U6298 ( .A(n6206), .ZN(n7747) );
  INV_X1 U6299 ( .A(n8674), .ZN(n9004) );
  INV_X1 U6300 ( .A(n10095), .ZN(n9180) );
  NAND2_X1 U6301 ( .A1(n8663), .A2(n7041), .ZN(n9053) );
  NOR2_X1 U6302 ( .A1(n5390), .A2(n9254), .ZN(n5407) );
  INV_X1 U6303 ( .A(n9308), .ZN(n9326) );
  NAND2_X1 U6304 ( .A1(n5321), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5330) );
  NOR2_X1 U6305 ( .A1(n5308), .A2(n5307), .ZN(n5319) );
  INV_X1 U6306 ( .A(n6943), .ZN(n6982) );
  AND2_X1 U6307 ( .A1(n8555), .A2(n8602), .ZN(n7025) );
  INV_X1 U6308 ( .A(n9342), .ZN(n9549) );
  INV_X1 U6309 ( .A(n9930), .ZN(n9497) );
  INV_X1 U6310 ( .A(n7806), .ZN(n8647) );
  AND2_X1 U6311 ( .A1(n8487), .A2(n8486), .ZN(n9749) );
  AND2_X1 U6312 ( .A1(n7017), .A2(n7016), .ZN(n7493) );
  INV_X1 U6313 ( .A(n9747), .ZN(n9572) );
  AND2_X1 U6314 ( .A1(n4940), .A2(n4939), .ZN(n5261) );
  AOI21_X1 U6315 ( .B1(n8816), .B2(n6045), .A(n4338), .ZN(n8710) );
  INV_X1 U6316 ( .A(n8855), .ZN(n9994) );
  OR2_X1 U6317 ( .A1(n5719), .A2(n5718), .ZN(n5736) );
  AND2_X1 U6318 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5649) );
  INV_X1 U6319 ( .A(n8856), .ZN(n7517) );
  AND2_X1 U6320 ( .A1(n8740), .A2(n5947), .ZN(n8785) );
  INV_X1 U6321 ( .A(n8818), .ZN(n9998) );
  AND2_X1 U6322 ( .A1(n8709), .A2(n6029), .ZN(n8815) );
  INV_X1 U6323 ( .A(n6192), .ZN(n8913) );
  INV_X1 U6324 ( .A(n10008), .ZN(n9725) );
  AND2_X1 U6325 ( .A1(n7046), .A2(n7043), .ZN(n10008) );
  INV_X1 U6326 ( .A(n8683), .ZN(n8677) );
  NAND2_X1 U6327 ( .A1(n7332), .A2(n7331), .ZN(n9084) );
  NOR2_X1 U6328 ( .A1(n10041), .A2(n6084), .ZN(n7544) );
  INV_X1 U6329 ( .A(n9170), .ZN(n10101) );
  INV_X1 U6330 ( .A(n9332), .ZN(n9313) );
  AND4_X1 U6331 ( .A1(n5376), .A2(n5375), .A3(n5374), .A4(n5373), .ZN(n9491)
         );
  INV_X1 U6332 ( .A(n5459), .ZN(n5346) );
  AND2_X1 U6333 ( .A1(n9803), .A2(n6847), .ZN(n9862) );
  INV_X1 U6334 ( .A(n9879), .ZN(n9917) );
  INV_X1 U6335 ( .A(n9922), .ZN(n9854) );
  AND2_X1 U6336 ( .A1(n7025), .A2(n8647), .ZN(n9926) );
  INV_X1 U6337 ( .A(n9550), .ZN(n9751) );
  AND2_X1 U6338 ( .A1(n8472), .A2(n8387), .ZN(n8583) );
  INV_X1 U6339 ( .A(n9949), .ZN(n9759) );
  AND2_X1 U6340 ( .A1(n8454), .A2(n8452), .ZN(n8576) );
  AND2_X1 U6341 ( .A1(n9945), .A2(n7356), .ZN(n9768) );
  INV_X1 U6342 ( .A(n9764), .ZN(n9975) );
  AND2_X1 U6343 ( .A1(n7493), .A2(n7210), .ZN(n9672) );
  AND2_X1 U6344 ( .A1(n6895), .A2(n6750), .ZN(n6973) );
  AND2_X1 U6345 ( .A1(n5315), .A2(n5304), .ZN(n9914) );
  AND2_X1 U6346 ( .A1(n5189), .A2(n5178), .ZN(n9853) );
  OR3_X1 U6347 ( .A1(n8006), .A2(n8215), .A3(n8222), .ZN(n7038) );
  INV_X1 U6348 ( .A(n9124), .ZN(n8758) );
  NAND2_X1 U6349 ( .A1(n7102), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10006) );
  INV_X1 U6350 ( .A(n8834), .ZN(n10000) );
  NAND2_X1 U6351 ( .A1(n9079), .A2(n10021), .ZN(n9063) );
  INV_X1 U6352 ( .A(n10119), .ZN(n10117) );
  INV_X1 U6353 ( .A(n10105), .ZN(n10103) );
  NOR2_X1 U6354 ( .A1(n10035), .A2(n10034), .ZN(n10039) );
  AND2_X1 U6355 ( .A1(n8006), .A2(n8222), .ZN(n10041) );
  XNOR2_X1 U6356 ( .A(n6070), .B(n6069), .ZN(n8006) );
  INV_X1 U6357 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7309) );
  INV_X1 U6358 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6870) );
  INV_X1 U6359 ( .A(n9637), .ZN(n9535) );
  INV_X1 U6360 ( .A(n9322), .ZN(n9315) );
  INV_X1 U6361 ( .A(n9438), .ZN(n9335) );
  AND4_X1 U6362 ( .A1(n5394), .A2(n5393), .A3(n5392), .A4(n5391), .ZN(n9477)
         );
  OR2_X1 U6363 ( .A1(n6846), .A2(n6845), .ZN(n9879) );
  NAND2_X1 U6364 ( .A1(n9945), .A2(n9926), .ZN(n9568) );
  NAND2_X1 U6365 ( .A1(n9945), .A2(n9924), .ZN(n9582) );
  OR2_X1 U6366 ( .A1(n7210), .A2(n5505), .ZN(n9949) );
  NAND2_X1 U6367 ( .A1(n6973), .A2(n6972), .ZN(n9987) );
  INV_X1 U6368 ( .A(n9983), .ZN(n9981) );
  AND2_X1 U6369 ( .A1(n9951), .A2(n9950), .ZN(n9957) );
  INV_X1 U6370 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7843) );
  INV_X1 U6371 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7260) );
  INV_X1 U6372 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6873) );
  NOR2_X1 U6373 ( .A1(n10161), .A2(n10160), .ZN(n10159) );
  NOR2_X1 U6374 ( .A1(n10148), .A2(n10147), .ZN(n10146) );
  NOR2_X1 U6375 ( .A1(n7038), .A2(n6771), .ZN(P2_U3966) );
  INV_X1 U6376 ( .A(n9358), .ZN(P1_U4006) );
  AND2_X1 U6377 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4887) );
  AND2_X1 U6378 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4888) );
  NAND2_X1 U6379 ( .A1(n5011), .A2(n4888), .ZN(n5597) );
  INV_X1 U6380 ( .A(SI_1_), .ZN(n4889) );
  NAND2_X1 U6381 ( .A1(n4890), .A2(SI_1_), .ZN(n4891) );
  NAND2_X1 U6382 ( .A1(n4892), .A2(n4891), .ZN(n5062) );
  INV_X1 U6383 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6794) );
  INV_X1 U6384 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6810) );
  XNOR2_X1 U6385 ( .A(n4893), .B(SI_2_), .ZN(n5063) );
  NAND2_X1 U6386 ( .A1(n5062), .A2(n5063), .ZN(n4896) );
  INV_X1 U6387 ( .A(n4893), .ZN(n4894) );
  NAND2_X1 U6388 ( .A1(n4894), .A2(SI_2_), .ZN(n4895) );
  NAND2_X1 U6389 ( .A1(n4896), .A2(n4895), .ZN(n5108) );
  INV_X1 U6390 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6793) );
  INV_X1 U6391 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n4897) );
  XNOR2_X1 U6392 ( .A(n4898), .B(SI_3_), .ZN(n5109) );
  INV_X1 U6393 ( .A(n4898), .ZN(n4899) );
  NAND2_X1 U6394 ( .A1(n4899), .A2(SI_3_), .ZN(n4900) );
  INV_X1 U6395 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6795) );
  INV_X1 U6396 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6802) );
  MUX2_X1 U6397 ( .A(n6795), .B(n6802), .S(n5400), .Z(n4901) );
  XNOR2_X1 U6398 ( .A(n4901), .B(SI_4_), .ZN(n5123) );
  INV_X1 U6399 ( .A(n4901), .ZN(n4902) );
  NAND2_X1 U6400 ( .A1(n4902), .A2(SI_4_), .ZN(n4903) );
  XNOR2_X1 U6401 ( .A(n4904), .B(SI_5_), .ZN(n5139) );
  INV_X1 U6402 ( .A(n4904), .ZN(n4905) );
  NAND2_X1 U6403 ( .A1(n4905), .A2(SI_5_), .ZN(n4906) );
  MUX2_X1 U6404 ( .A(n6798), .B(n6804), .S(n5400), .Z(n4907) );
  XNOR2_X1 U6405 ( .A(n4907), .B(SI_6_), .ZN(n5150) );
  INV_X1 U6406 ( .A(n4907), .ZN(n4908) );
  MUX2_X1 U6407 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n5400), .Z(n4910) );
  XNOR2_X1 U6408 ( .A(n4910), .B(SI_7_), .ZN(n5163) );
  INV_X1 U6409 ( .A(n5163), .ZN(n4909) );
  NAND2_X1 U6410 ( .A1(n4910), .A2(SI_7_), .ZN(n4911) );
  MUX2_X1 U6411 ( .A(n6827), .B(n4912), .S(n5400), .Z(n4914) );
  INV_X1 U6412 ( .A(SI_8_), .ZN(n4913) );
  INV_X1 U6413 ( .A(n4914), .ZN(n4915) );
  NAND2_X1 U6414 ( .A1(n4915), .A2(SI_8_), .ZN(n4916) );
  NAND2_X1 U6415 ( .A1(n4917), .A2(n4916), .ZN(n5171) );
  MUX2_X1 U6416 ( .A(n6870), .B(n4918), .S(n5400), .Z(n4920) );
  NAND2_X1 U6417 ( .A1(n4920), .A2(n4919), .ZN(n4923) );
  INV_X1 U6418 ( .A(n4920), .ZN(n4921) );
  NAND2_X1 U6419 ( .A1(n4921), .A2(SI_9_), .ZN(n4922) );
  MUX2_X1 U6420 ( .A(n6875), .B(n6873), .S(n5400), .Z(n4924) );
  INV_X1 U6421 ( .A(n4924), .ZN(n4925) );
  NAND2_X1 U6422 ( .A1(n4925), .A2(SI_10_), .ZN(n4926) );
  MUX2_X1 U6423 ( .A(n6889), .B(n6887), .S(n5400), .Z(n4929) );
  INV_X1 U6424 ( .A(n4929), .ZN(n4930) );
  NAND2_X1 U6425 ( .A1(n4930), .A2(SI_11_), .ZN(n4931) );
  MUX2_X1 U6426 ( .A(n7000), .B(n7001), .S(n5400), .Z(n4932) );
  INV_X1 U6427 ( .A(n4932), .ZN(n4933) );
  NAND2_X1 U6428 ( .A1(n4933), .A2(SI_12_), .ZN(n4934) );
  NAND2_X1 U6429 ( .A1(n4935), .A2(n4934), .ZN(n5233) );
  MUX2_X1 U6430 ( .A(n7113), .B(n7128), .S(n5400), .Z(n4937) );
  INV_X1 U6431 ( .A(n4937), .ZN(n4938) );
  NAND2_X1 U6432 ( .A1(n4938), .A2(SI_13_), .ZN(n4939) );
  MUX2_X1 U6433 ( .A(n7158), .B(n7159), .S(n5400), .Z(n4942) );
  XNOR2_X1 U6434 ( .A(n4942), .B(SI_14_), .ZN(n5045) );
  INV_X1 U6435 ( .A(n5045), .ZN(n4945) );
  INV_X1 U6436 ( .A(n4942), .ZN(n4943) );
  NAND2_X1 U6437 ( .A1(n4943), .A2(SI_14_), .ZN(n4944) );
  MUX2_X1 U6438 ( .A(n7259), .B(n7260), .S(n5400), .Z(n4947) );
  INV_X1 U6439 ( .A(SI_15_), .ZN(n4946) );
  NAND2_X1 U6440 ( .A1(n4947), .A2(n4946), .ZN(n4950) );
  INV_X1 U6441 ( .A(n4947), .ZN(n4948) );
  NAND2_X1 U6442 ( .A1(n4948), .A2(SI_15_), .ZN(n4949) );
  NAND2_X1 U6443 ( .A1(n4950), .A2(n4949), .ZN(n5278) );
  MUX2_X1 U6444 ( .A(n7309), .B(n4951), .S(n5400), .Z(n4953) );
  INV_X1 U6445 ( .A(SI_16_), .ZN(n4952) );
  NAND2_X1 U6446 ( .A1(n4953), .A2(n4952), .ZN(n4956) );
  INV_X1 U6447 ( .A(n4953), .ZN(n4954) );
  NAND2_X1 U6448 ( .A1(n4954), .A2(SI_16_), .ZN(n4955) );
  MUX2_X1 U6449 ( .A(n7341), .B(n7342), .S(n5400), .Z(n4957) );
  XNOR2_X1 U6450 ( .A(n4957), .B(SI_17_), .ZN(n5297) );
  INV_X1 U6451 ( .A(n5297), .ZN(n4959) );
  INV_X1 U6452 ( .A(n4957), .ZN(n4958) );
  MUX2_X1 U6453 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5400), .Z(n4961) );
  XNOR2_X1 U6454 ( .A(n4961), .B(SI_18_), .ZN(n5313) );
  NAND2_X1 U6455 ( .A1(n5314), .A2(n4960), .ZN(n4963) );
  NAND2_X1 U6456 ( .A1(n4961), .A2(SI_18_), .ZN(n4962) );
  NAND2_X1 U6457 ( .A1(n4963), .A2(n4962), .ZN(n5031) );
  MUX2_X1 U6458 ( .A(n7662), .B(n7663), .S(n5400), .Z(n4965) );
  INV_X1 U6459 ( .A(SI_19_), .ZN(n4964) );
  NAND2_X1 U6460 ( .A1(n4965), .A2(n4964), .ZN(n4968) );
  INV_X1 U6461 ( .A(n4965), .ZN(n4966) );
  NAND2_X1 U6462 ( .A1(n4966), .A2(SI_19_), .ZN(n4967) );
  NAND2_X1 U6463 ( .A1(n4968), .A2(n4967), .ZN(n5030) );
  MUX2_X1 U6464 ( .A(n7744), .B(n7804), .S(n5400), .Z(n4969) );
  INV_X1 U6465 ( .A(SI_20_), .ZN(n6475) );
  NAND2_X1 U6466 ( .A1(n4969), .A2(n6475), .ZN(n4972) );
  INV_X1 U6467 ( .A(n4969), .ZN(n4970) );
  NAND2_X1 U6468 ( .A1(n4970), .A2(SI_20_), .ZN(n4971) );
  NAND2_X1 U6469 ( .A1(n5326), .A2(n5325), .ZN(n4973) );
  MUX2_X1 U6470 ( .A(n7819), .B(n7843), .S(n5400), .Z(n4974) );
  XNOR2_X1 U6471 ( .A(n4974), .B(SI_21_), .ZN(n5340) );
  INV_X1 U6472 ( .A(n4974), .ZN(n4975) );
  NAND2_X1 U6473 ( .A1(n4975), .A2(SI_21_), .ZN(n4976) );
  MUX2_X1 U6474 ( .A(n7849), .B(n7846), .S(n5400), .Z(n4978) );
  INV_X1 U6475 ( .A(SI_22_), .ZN(n4977) );
  NAND2_X1 U6476 ( .A1(n4978), .A2(n4977), .ZN(n4981) );
  INV_X1 U6477 ( .A(n4978), .ZN(n4979) );
  NAND2_X1 U6478 ( .A1(n4979), .A2(SI_22_), .ZN(n4980) );
  NAND2_X1 U6479 ( .A1(n4981), .A2(n4980), .ZN(n5355) );
  INV_X1 U6480 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n4983) );
  INV_X1 U6481 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n4982) );
  MUX2_X1 U6482 ( .A(n4983), .B(n4982), .S(n5400), .Z(n4985) );
  INV_X1 U6483 ( .A(SI_23_), .ZN(n4984) );
  NAND2_X1 U6484 ( .A1(n4985), .A2(n4984), .ZN(n5368) );
  INV_X1 U6485 ( .A(n4985), .ZN(n4986) );
  NAND2_X1 U6486 ( .A1(n4986), .A2(SI_23_), .ZN(n4987) );
  XNOR2_X1 U6487 ( .A(n5367), .B(n5366), .ZN(n7951) );
  NAND2_X1 U6488 ( .A1(n5235), .A2(n5238), .ZN(n5032) );
  INV_X1 U6489 ( .A(n5032), .ZN(n4990) );
  NOR2_X1 U6490 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n4989) );
  NOR2_X1 U6491 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n4994) );
  NOR2_X1 U6492 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n4995) );
  NAND2_X1 U6493 ( .A1(n5064), .A2(n4998), .ZN(n5066) );
  NOR2_X1 U6494 ( .A1(n5016), .A2(n5002), .ZN(n5007) );
  NAND2_X1 U6495 ( .A1(n5008), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5009) );
  NAND2_X2 U6496 ( .A1(n5522), .A2(n6948), .ZN(n5080) );
  AND2_X2 U6497 ( .A1(n5080), .A2(n5400), .ZN(n5114) );
  INV_X2 U6498 ( .A(n5165), .ZN(n5454) );
  NAND2_X1 U6499 ( .A1(n7951), .A2(n5454), .ZN(n5013) );
  AND2_X2 U6500 ( .A1(n5080), .A2(n6799), .ZN(n5078) );
  BUF_X4 U6501 ( .A(n5078), .Z(n8344) );
  NAND2_X1 U6502 ( .A1(n8344), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5012) );
  NAND2_X1 U6503 ( .A1(n6816), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5026) );
  INV_X1 U6504 ( .A(n5022), .ZN(n9703) );
  AND2_X2 U6505 ( .A1(n9703), .A2(n9708), .ZN(n5085) );
  INV_X2 U6506 ( .A(n5526), .ZN(n6818) );
  NAND2_X1 U6507 ( .A1(n6818), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5025) );
  INV_X1 U6508 ( .A(n9708), .ZN(n5020) );
  INV_X1 U6509 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9218) );
  INV_X1 U6510 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9246) );
  NAND2_X1 U6511 ( .A1(n5129), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5144) );
  NAND2_X1 U6512 ( .A1(n5157), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5181) );
  OR2_X2 U6513 ( .A1(n5181), .A2(n5180), .ZN(n5194) );
  OR2_X2 U6514 ( .A1(n5244), .A2(n5243), .ZN(n5252) );
  INV_X1 U6515 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5251) );
  INV_X1 U6516 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5051) );
  NAND2_X1 U6517 ( .A1(n5284), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5285) );
  INV_X1 U6518 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5272) );
  INV_X1 U6519 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5307) );
  INV_X1 U6520 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5329) );
  INV_X1 U6521 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9298) );
  INV_X1 U6522 ( .A(n5359), .ZN(n5021) );
  NAND2_X1 U6523 ( .A1(n5359), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5372) );
  AOI21_X1 U6524 ( .B1(n9218), .B2(n5021), .A(n5370), .ZN(n9495) );
  NAND2_X1 U6525 ( .A1(n5459), .A2(n9495), .ZN(n5024) );
  NAND2_X1 U6526 ( .A1(n6817), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5023) );
  OR2_X1 U6527 ( .A1(n5321), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5027) );
  NAND2_X1 U6528 ( .A1(n5330), .A2(n5027), .ZN(n9554) );
  INV_X4 U6529 ( .A(n5350), .ZN(n6816) );
  AOI22_X1 U6530 ( .A1(n6816), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n6818), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n5029) );
  NAND2_X1 U6531 ( .A1(n6817), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5028) );
  OAI211_X1 U6532 ( .C1(n9554), .C2(n5346), .A(n5029), .B(n5028), .ZN(n9343)
         );
  INV_X1 U6533 ( .A(n9343), .ZN(n9537) );
  XNOR2_X1 U6534 ( .A(n5031), .B(n5030), .ZN(n7661) );
  NAND2_X1 U6535 ( .A1(n7661), .A2(n5454), .ZN(n5044) );
  NOR2_X1 U6536 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5033) );
  NAND4_X1 U6537 ( .A1(n5035), .A2(n5034), .A3(n5033), .A4(n5203), .ZN(n5036)
         );
  NOR2_X2 U6538 ( .A1(n5134), .A2(n5036), .ZN(n5047) );
  NAND2_X1 U6539 ( .A1(n5280), .A2(n5038), .ZN(n5269) );
  INV_X1 U6540 ( .A(n5269), .ZN(n5040) );
  INV_X1 U6541 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5039) );
  NAND3_X1 U6542 ( .A1(n5040), .A2(n5039), .A3(n4871), .ZN(n5465) );
  NAND2_X1 U6543 ( .A1(n5465), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5042) );
  INV_X1 U6544 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5041) );
  CLKBUF_X3 U6545 ( .A(n5080), .Z(n5140) );
  AOI22_X1 U6546 ( .A1(n8344), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9497), .B2(
        n6769), .ZN(n5043) );
  INV_X1 U6547 ( .A(n9644), .ZN(n9558) );
  XNOR2_X1 U6548 ( .A(n5046), .B(n5045), .ZN(n7157) );
  NAND2_X1 U6549 ( .A1(n7157), .A2(n5454), .ZN(n5050) );
  OR2_X1 U6550 ( .A1(n5047), .A2(n9695), .ZN(n5048) );
  XNOR2_X1 U6551 ( .A(n5048), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7618) );
  AOI22_X1 U6552 ( .A1(n8344), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6769), .B2(
        n7618), .ZN(n5049) );
  NAND2_X1 U6553 ( .A1(n6816), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5056) );
  AND2_X1 U6554 ( .A1(n5254), .A2(n5051), .ZN(n5052) );
  NOR2_X1 U6555 ( .A1(n5284), .A2(n5052), .ZN(n8098) );
  NAND2_X1 U6556 ( .A1(n5459), .A2(n8098), .ZN(n5055) );
  NAND2_X1 U6557 ( .A1(n6818), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5054) );
  NAND2_X1 U6558 ( .A1(n6817), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5053) );
  NAND4_X1 U6559 ( .A1(n5056), .A2(n5055), .A3(n5054), .A4(n5053), .ZN(n9347)
         );
  AND2_X1 U6560 ( .A1(n9669), .A2(n9347), .ZN(n5260) );
  INV_X1 U6561 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n5057) );
  NAND2_X1 U6562 ( .A1(n5102), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5060) );
  NAND2_X1 U6563 ( .A1(n5085), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5059) );
  NAND2_X1 U6564 ( .A1(n5087), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5058) );
  XNOR2_X1 U6565 ( .A(n5062), .B(n5063), .ZN(n6811) );
  NAND2_X1 U6566 ( .A1(n5078), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5070) );
  NOR2_X1 U6567 ( .A1(n5064), .A2(n9695), .ZN(n5065) );
  MUX2_X1 U6568 ( .A(n9695), .B(n5065), .S(P1_IR_REG_2__SCAN_IN), .Z(n5067) );
  INV_X1 U6569 ( .A(n4313), .ZN(n5068) );
  OR2_X1 U6570 ( .A1(n5140), .A2(n5068), .ZN(n5069) );
  NAND2_X1 U6571 ( .A1(n7202), .A2(n7010), .ZN(n8377) );
  INV_X2 U6572 ( .A(n7010), .ZN(n7368) );
  NAND2_X1 U6573 ( .A1(n5086), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5074) );
  NAND2_X1 U6574 ( .A1(n5087), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5072) );
  NAND2_X1 U6575 ( .A1(n5102), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5071) );
  INV_X1 U6576 ( .A(n6809), .ZN(n5077) );
  NAND2_X1 U6577 ( .A1(n5114), .A2(n5077), .ZN(n5083) );
  NAND2_X1 U6578 ( .A1(n5078), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5082) );
  INV_X1 U6579 ( .A(n6849), .ZN(n5079) );
  OR2_X1 U6580 ( .A1(n5080), .A2(n5079), .ZN(n5081) );
  NAND2_X1 U6581 ( .A1(n5085), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5091) );
  NAND2_X1 U6582 ( .A1(n5102), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5090) );
  NAND2_X1 U6583 ( .A1(n5087), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5088) );
  INV_X1 U6584 ( .A(SI_0_), .ZN(n5093) );
  INV_X1 U6585 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5092) );
  OAI21_X1 U6586 ( .B1(n6799), .B2(n5093), .A(n5092), .ZN(n5095) );
  AND2_X1 U6587 ( .A1(n5095), .A2(n5094), .ZN(n9709) );
  OAI21_X2 U6588 ( .B1(n5140), .B2(n5097), .A(n5096), .ZN(n6519) );
  NAND2_X1 U6589 ( .A1(n6529), .A2(n5084), .ZN(n5098) );
  NAND2_X1 U6590 ( .A1(n7202), .A2(n7368), .ZN(n5099) );
  INV_X1 U6591 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n5100) );
  INV_X1 U6592 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5101) );
  NAND2_X1 U6593 ( .A1(n5102), .A2(n5101), .ZN(n5106) );
  INV_X1 U6594 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5103) );
  NAND2_X1 U6595 ( .A1(n6817), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5104) );
  AND4_X2 U6596 ( .A1(n5107), .A2(n5106), .A3(n5105), .A4(n5104), .ZN(n7350)
         );
  INV_X1 U6597 ( .A(n7350), .ZN(n9356) );
  NAND2_X1 U6598 ( .A1(n8344), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5115) );
  XNOR2_X1 U6599 ( .A(n5108), .B(n5109), .ZN(n6801) );
  INV_X1 U6600 ( .A(n6801), .ZN(n5113) );
  NAND2_X1 U6601 ( .A1(n5066), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5111) );
  NAND2_X1 U6602 ( .A1(n5111), .A2(n5110), .ZN(n5124) );
  OR2_X1 U6603 ( .A1(n5111), .A2(n5110), .ZN(n5112) );
  AND2_X1 U6604 ( .A1(n5124), .A2(n5112), .ZN(n6909) );
  INV_X2 U6605 ( .A(n9230), .ZN(n7455) );
  NAND2_X1 U6606 ( .A1(n9356), .A2(n7455), .ZN(n7344) );
  NAND2_X1 U6607 ( .A1(n7350), .A2(n9230), .ZN(n8372) );
  NAND2_X1 U6608 ( .A1(n7201), .A2(n8564), .ZN(n7200) );
  NAND2_X1 U6609 ( .A1(n7350), .A2(n7455), .ZN(n5116) );
  NAND2_X1 U6610 ( .A1(n7200), .A2(n5116), .ZN(n7347) );
  NAND2_X1 U6611 ( .A1(n6816), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5121) );
  NOR2_X1 U6612 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5117) );
  NOR2_X1 U6613 ( .A1(n5129), .A2(n5117), .ZN(n7190) );
  NAND2_X1 U6614 ( .A1(n5459), .A2(n7190), .ZN(n5120) );
  NAND2_X1 U6615 ( .A1(n6818), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5119) );
  NAND2_X1 U6616 ( .A1(n6817), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5118) );
  XNOR2_X1 U6617 ( .A(n5123), .B(n5122), .ZN(n6803) );
  NAND2_X1 U6618 ( .A1(n5078), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5127) );
  NAND2_X1 U6619 ( .A1(n5124), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5125) );
  XNOR2_X1 U6620 ( .A(n5125), .B(P1_IR_REG_4__SCAN_IN), .ZN(n6955) );
  NAND2_X1 U6621 ( .A1(n6769), .A2(n6955), .ZN(n5126) );
  OAI211_X1 U6622 ( .C1(n5165), .C2(n6803), .A(n5127), .B(n5126), .ZN(n7357)
         );
  NAND2_X1 U6623 ( .A1(n7287), .A2(n7357), .ZN(n7285) );
  INV_X1 U6624 ( .A(n7357), .ZN(n9961) );
  NAND2_X1 U6625 ( .A1(n9355), .A2(n9961), .ZN(n8420) );
  NAND2_X1 U6626 ( .A1(n7285), .A2(n8420), .ZN(n8566) );
  NAND2_X1 U6627 ( .A1(n7287), .A2(n9961), .ZN(n5128) );
  OAI21_X1 U6628 ( .B1(n5129), .B2(P1_REG3_REG_5__SCAN_IN), .A(n5144), .ZN(
        n9928) );
  INV_X1 U6629 ( .A(n9928), .ZN(n7383) );
  NAND2_X1 U6630 ( .A1(n5459), .A2(n7383), .ZN(n5133) );
  NAND2_X1 U6631 ( .A1(n6816), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5132) );
  NAND2_X1 U6632 ( .A1(n6818), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5131) );
  NAND2_X1 U6633 ( .A1(n6817), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5130) );
  NAND2_X1 U6634 ( .A1(n5134), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5135) );
  MUX2_X1 U6635 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5135), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5137) );
  NOR2_X1 U6636 ( .A1(n5134), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5167) );
  INV_X1 U6637 ( .A(n5167), .ZN(n5136) );
  INV_X1 U6638 ( .A(n9819), .ZN(n6808) );
  NAND2_X1 U6639 ( .A1(n7438), .A2(n9925), .ZN(n8422) );
  NAND2_X1 U6640 ( .A1(n9354), .A2(n7386), .ZN(n8429) );
  NAND2_X1 U6641 ( .A1(n9354), .A2(n9925), .ZN(n5142) );
  NAND2_X1 U6642 ( .A1(n6816), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5149) );
  AND2_X1 U6643 ( .A1(n5144), .A2(n5143), .ZN(n5145) );
  NOR2_X1 U6644 ( .A1(n5157), .A2(n5145), .ZN(n7446) );
  NAND2_X1 U6645 ( .A1(n5459), .A2(n7446), .ZN(n5148) );
  NAND2_X1 U6646 ( .A1(n6818), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5147) );
  NAND2_X1 U6647 ( .A1(n6817), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5146) );
  XNOR2_X1 U6648 ( .A(n5151), .B(n5150), .ZN(n6805) );
  OR2_X1 U6649 ( .A1(n6805), .A2(n5165), .ZN(n5154) );
  OR2_X1 U6650 ( .A1(n5167), .A2(n9695), .ZN(n5152) );
  XNOR2_X1 U6651 ( .A(n5152), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6933) );
  AOI22_X1 U6652 ( .A1(n8344), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6769), .B2(
        n6933), .ZN(n5153) );
  NAND2_X1 U6653 ( .A1(n5154), .A2(n5153), .ZN(n8434) );
  NAND2_X1 U6654 ( .A1(n8431), .A2(n8434), .ZN(n8610) );
  INV_X1 U6655 ( .A(n8431), .ZN(n9353) );
  NAND2_X1 U6656 ( .A1(n9353), .A2(n9967), .ZN(n8608) );
  NAND2_X1 U6657 ( .A1(n8431), .A2(n9967), .ZN(n5156) );
  NAND2_X1 U6658 ( .A1(n7433), .A2(n5156), .ZN(n7397) );
  NAND2_X1 U6659 ( .A1(n6816), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5162) );
  OR2_X1 U6660 ( .A1(n5157), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5158) );
  AND2_X1 U6661 ( .A1(n5181), .A2(n5158), .ZN(n7505) );
  NAND2_X1 U6662 ( .A1(n5459), .A2(n7505), .ZN(n5161) );
  NAND2_X1 U6663 ( .A1(n6818), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5160) );
  NAND2_X1 U6664 ( .A1(n6817), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5159) );
  XNOR2_X1 U6665 ( .A(n5164), .B(n5163), .ZN(n6812) );
  NAND2_X1 U6666 ( .A1(n6812), .A2(n5454), .ZN(n5169) );
  NAND2_X1 U6667 ( .A1(n5167), .A2(n5166), .ZN(n5205) );
  NAND2_X1 U6668 ( .A1(n5205), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5174) );
  XNOR2_X1 U6669 ( .A(n5174), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6934) );
  AOI22_X1 U6670 ( .A1(n8344), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6769), .B2(
        n6934), .ZN(n5168) );
  NAND2_X1 U6671 ( .A1(n5169), .A2(n5168), .ZN(n8441) );
  OR2_X1 U6672 ( .A1(n8438), .A2(n8441), .ZN(n8430) );
  NAND2_X1 U6673 ( .A1(n8441), .A2(n8438), .ZN(n8425) );
  NAND2_X1 U6674 ( .A1(n8430), .A2(n8425), .ZN(n7396) );
  INV_X1 U6675 ( .A(n8441), .ZN(n8436) );
  NAND2_X1 U6676 ( .A1(n8436), .A2(n8438), .ZN(n5170) );
  INV_X1 U6677 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5173) );
  NAND2_X1 U6678 ( .A1(n5174), .A2(n5173), .ZN(n5175) );
  NAND2_X1 U6679 ( .A1(n5175), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5177) );
  NAND2_X1 U6680 ( .A1(n5177), .A2(n5176), .ZN(n5189) );
  OR2_X1 U6681 ( .A1(n5177), .A2(n5176), .ZN(n5178) );
  AOI22_X1 U6682 ( .A1(n8344), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6769), .B2(
        n9853), .ZN(n5179) );
  NAND2_X1 U6683 ( .A1(n6816), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5186) );
  NAND2_X1 U6684 ( .A1(n5181), .A2(n5180), .ZN(n5182) );
  AND2_X1 U6685 ( .A1(n5194), .A2(n5182), .ZN(n7497) );
  NAND2_X1 U6686 ( .A1(n5459), .A2(n7497), .ZN(n5185) );
  NAND2_X1 U6687 ( .A1(n6818), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5184) );
  NAND2_X1 U6688 ( .A1(n6817), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5183) );
  NAND2_X1 U6689 ( .A1(n7498), .A2(n7589), .ZN(n8458) );
  INV_X1 U6690 ( .A(n7589), .ZN(n9351) );
  NAND2_X1 U6691 ( .A1(n7498), .A2(n9351), .ZN(n5187) );
  XNOR2_X1 U6692 ( .A(n5188), .B(n4876), .ZN(n6830) );
  NAND2_X1 U6693 ( .A1(n6830), .A2(n5454), .ZN(n5192) );
  NAND2_X1 U6694 ( .A1(n5189), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5190) );
  XNOR2_X1 U6695 ( .A(n5190), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9874) );
  AOI22_X1 U6696 ( .A1(n8344), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6769), .B2(
        n9874), .ZN(n5191) );
  AND2_X1 U6697 ( .A1(n5194), .A2(n5193), .ZN(n5195) );
  NOR2_X1 U6698 ( .A1(n5212), .A2(n5195), .ZN(n7684) );
  NAND2_X1 U6699 ( .A1(n5459), .A2(n7684), .ZN(n5199) );
  NAND2_X1 U6700 ( .A1(n6816), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5198) );
  NAND2_X1 U6701 ( .A1(n6818), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5197) );
  NAND2_X1 U6702 ( .A1(n6817), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5196) );
  NAND4_X1 U6703 ( .A1(n5199), .A2(n5198), .A3(n5197), .A4(n5196), .ZN(n9350)
         );
  OR2_X1 U6704 ( .A1(n7698), .A2(n9350), .ZN(n5201) );
  AND2_X1 U6705 ( .A1(n7698), .A2(n9350), .ZN(n5200) );
  XNOR2_X1 U6706 ( .A(n5202), .B(n4875), .ZN(n6872) );
  NAND2_X1 U6707 ( .A1(n6872), .A2(n5454), .ZN(n5211) );
  INV_X1 U6708 ( .A(n5203), .ZN(n5204) );
  NAND2_X1 U6709 ( .A1(n5207), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5206) );
  MUX2_X1 U6710 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5206), .S(
        P1_IR_REG_10__SCAN_IN), .Z(n5209) );
  INV_X1 U6711 ( .A(n5236), .ZN(n5208) );
  NAND2_X1 U6712 ( .A1(n5209), .A2(n5208), .ZN(n6943) );
  AOI22_X1 U6713 ( .A1(n8344), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6769), .B2(
        n6982), .ZN(n5210) );
  NAND2_X1 U6714 ( .A1(n6816), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5217) );
  NAND2_X1 U6715 ( .A1(n6818), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5216) );
  NOR2_X1 U6716 ( .A1(n5212), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5213) );
  OR2_X1 U6717 ( .A1(n5224), .A2(n5213), .ZN(n7694) );
  INV_X1 U6718 ( .A(n7694), .ZN(n7605) );
  NAND2_X1 U6719 ( .A1(n5459), .A2(n7605), .ZN(n5215) );
  NAND2_X1 U6720 ( .A1(n6817), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5214) );
  NAND2_X1 U6721 ( .A1(n7707), .A2(n7736), .ZN(n8456) );
  NAND2_X1 U6722 ( .A1(n8466), .A2(n8456), .ZN(n8578) );
  NAND2_X1 U6723 ( .A1(n7597), .A2(n8578), .ZN(n7596) );
  INV_X1 U6724 ( .A(n7736), .ZN(n9349) );
  OR2_X1 U6725 ( .A1(n7707), .A2(n9349), .ZN(n5218) );
  NAND2_X1 U6726 ( .A1(n7596), .A2(n5218), .ZN(n7731) );
  XNOR2_X1 U6727 ( .A(n5220), .B(n5219), .ZN(n5765) );
  NAND2_X1 U6728 ( .A1(n5765), .A2(n5454), .ZN(n5223) );
  OR2_X1 U6729 ( .A1(n5236), .A2(n9695), .ZN(n5221) );
  XNOR2_X1 U6730 ( .A(n5221), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7166) );
  AOI22_X1 U6731 ( .A1(n8344), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6769), .B2(
        n7166), .ZN(n5222) );
  NAND2_X1 U6732 ( .A1(n6816), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5229) );
  OR2_X1 U6733 ( .A1(n5224), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5225) );
  AND2_X1 U6734 ( .A1(n5244), .A2(n5225), .ZN(n7774) );
  NAND2_X1 U6735 ( .A1(n5459), .A2(n7774), .ZN(n5228) );
  NAND2_X1 U6736 ( .A1(n6818), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5227) );
  NAND2_X1 U6737 ( .A1(n6817), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5226) );
  NAND4_X1 U6738 ( .A1(n5229), .A2(n5228), .A3(n5227), .A4(n5226), .ZN(n9753)
         );
  NAND2_X1 U6739 ( .A1(n6600), .A2(n9753), .ZN(n5230) );
  NAND2_X1 U6740 ( .A1(n7731), .A2(n5230), .ZN(n5232) );
  OR2_X1 U6741 ( .A1(n6600), .A2(n9753), .ZN(n5231) );
  NAND2_X1 U6742 ( .A1(n5232), .A2(n5231), .ZN(n9746) );
  XNOR2_X1 U6743 ( .A(n5234), .B(n5233), .ZN(n6999) );
  NAND2_X1 U6744 ( .A1(n6999), .A2(n5454), .ZN(n5242) );
  NAND2_X1 U6745 ( .A1(n5236), .A2(n5235), .ZN(n5237) );
  NAND2_X1 U6746 ( .A1(n5237), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5239) );
  NAND2_X1 U6747 ( .A1(n5239), .A2(n5238), .ZN(n5263) );
  OR2_X1 U6748 ( .A1(n5239), .A2(n5238), .ZN(n5240) );
  AOI22_X1 U6749 ( .A1(n8344), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6769), .B2(
        n7249), .ZN(n5241) );
  NAND2_X1 U6750 ( .A1(n5244), .A2(n5243), .ZN(n5245) );
  AND2_X1 U6751 ( .A1(n5252), .A2(n5245), .ZN(n9760) );
  NAND2_X1 U6752 ( .A1(n5459), .A2(n9760), .ZN(n5249) );
  NAND2_X1 U6753 ( .A1(n6818), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5248) );
  NAND2_X1 U6754 ( .A1(n6816), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5247) );
  NAND2_X1 U6755 ( .A1(n6817), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5246) );
  NAND2_X1 U6756 ( .A1(n9761), .A2(n7772), .ZN(n8486) );
  NAND2_X1 U6757 ( .A1(n9761), .A2(n9348), .ZN(n5250) );
  NAND2_X1 U6758 ( .A1(n5252), .A2(n5251), .ZN(n5253) );
  AND2_X1 U6759 ( .A1(n5254), .A2(n5253), .ZN(n7903) );
  NAND2_X1 U6760 ( .A1(n5459), .A2(n7903), .ZN(n5258) );
  NAND2_X1 U6761 ( .A1(n6816), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5257) );
  NAND2_X1 U6762 ( .A1(n6818), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5256) );
  NAND2_X1 U6763 ( .A1(n6817), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5255) );
  NAND4_X1 U6764 ( .A1(n5258), .A2(n5257), .A3(n5256), .A4(n5255), .ZN(n9752)
         );
  INV_X1 U6765 ( .A(n7966), .ZN(n5259) );
  NOR2_X1 U6766 ( .A1(n5260), .A2(n5259), .ZN(n5267) );
  XNOR2_X1 U6767 ( .A(n5262), .B(n5261), .ZN(n7112) );
  NAND2_X1 U6768 ( .A1(n7112), .A2(n5454), .ZN(n5266) );
  NAND2_X1 U6769 ( .A1(n5263), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5264) );
  XNOR2_X1 U6770 ( .A(n5264), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7611) );
  AOI22_X1 U6771 ( .A1(n8344), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6769), .B2(
        n7611), .ZN(n5265) );
  OAI21_X1 U6772 ( .B1(n7896), .B2(n9752), .A(n7904), .ZN(n7967) );
  NAND2_X1 U6773 ( .A1(n5267), .A2(n7967), .ZN(n8113) );
  OR2_X1 U6774 ( .A1(n9669), .A2(n9347), .ZN(n8114) );
  NAND2_X1 U6775 ( .A1(n7240), .A2(n5454), .ZN(n5271) );
  NAND2_X1 U6776 ( .A1(n5269), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5300) );
  XNOR2_X1 U6777 ( .A(n5300), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9900) );
  AOI22_X1 U6778 ( .A1(n8344), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6769), .B2(
        n9900), .ZN(n5270) );
  NAND2_X1 U6779 ( .A1(n5285), .A2(n5272), .ZN(n5273) );
  AND2_X1 U6780 ( .A1(n5308), .A2(n5273), .ZN(n8179) );
  NAND2_X1 U6781 ( .A1(n8179), .A2(n5459), .ZN(n5277) );
  NAND2_X1 U6782 ( .A1(n6816), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5276) );
  NAND2_X1 U6783 ( .A1(n6818), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5275) );
  NAND2_X1 U6784 ( .A1(n6817), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5274) );
  NAND2_X1 U6785 ( .A1(n5294), .A2(n9570), .ZN(n8480) );
  INV_X1 U6786 ( .A(n8585), .ZN(n8132) );
  XNOR2_X1 U6787 ( .A(n5279), .B(n5278), .ZN(n7258) );
  NAND2_X1 U6788 ( .A1(n7258), .A2(n5454), .ZN(n5283) );
  OR2_X1 U6789 ( .A1(n5280), .A2(n9695), .ZN(n5281) );
  XNOR2_X1 U6790 ( .A(n5281), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9888) );
  AOI22_X1 U6791 ( .A1(n8344), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6769), .B2(
        n9888), .ZN(n5282) );
  INV_X1 U6792 ( .A(n9662), .ZN(n8119) );
  NAND2_X1 U6793 ( .A1(n6816), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5290) );
  OR2_X1 U6794 ( .A1(n5284), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5286) );
  AND2_X1 U6795 ( .A1(n5286), .A2(n5285), .ZN(n8117) );
  NAND2_X1 U6796 ( .A1(n5459), .A2(n8117), .ZN(n5289) );
  NAND2_X1 U6797 ( .A1(n6818), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5288) );
  NAND2_X1 U6798 ( .A1(n6817), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5287) );
  NAND4_X1 U6799 ( .A1(n5290), .A2(n5289), .A3(n5288), .A4(n5287), .ZN(n9346)
         );
  INV_X1 U6800 ( .A(n9346), .ZN(n8175) );
  NAND2_X1 U6801 ( .A1(n8119), .A2(n8175), .ZN(n8126) );
  AND2_X1 U6802 ( .A1(n8132), .A2(n8126), .ZN(n5292) );
  AND2_X1 U6803 ( .A1(n8114), .A2(n5292), .ZN(n5291) );
  NAND2_X1 U6804 ( .A1(n8113), .A2(n5291), .ZN(n8129) );
  INV_X1 U6805 ( .A(n5292), .ZN(n5293) );
  NAND2_X1 U6806 ( .A1(n9662), .A2(n9346), .ZN(n8124) );
  OR2_X1 U6807 ( .A1(n5293), .A2(n8124), .ZN(n8128) );
  INV_X1 U6808 ( .A(n9570), .ZN(n9345) );
  NAND2_X1 U6809 ( .A1(n5294), .A2(n9345), .ZN(n5295) );
  AND2_X1 U6810 ( .A1(n8128), .A2(n5295), .ZN(n5296) );
  XNOR2_X1 U6811 ( .A(n5298), .B(n5297), .ZN(n7340) );
  NAND2_X1 U6812 ( .A1(n7340), .A2(n5454), .ZN(n5306) );
  NAND2_X1 U6813 ( .A1(n5300), .A2(n5299), .ZN(n5301) );
  NAND2_X1 U6814 ( .A1(n5301), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5303) );
  NAND2_X1 U6815 ( .A1(n5303), .A2(n5302), .ZN(n5315) );
  OR2_X1 U6816 ( .A1(n5303), .A2(n5302), .ZN(n5304) );
  AOI22_X1 U6817 ( .A1(n8344), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6769), .B2(
        n9914), .ZN(n5305) );
  AND2_X1 U6818 ( .A1(n5308), .A2(n5307), .ZN(n5309) );
  OR2_X1 U6819 ( .A1(n5309), .A2(n5319), .ZN(n9565) );
  AOI22_X1 U6820 ( .A1(n6817), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n6818), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n5311) );
  NAND2_X1 U6821 ( .A1(n6816), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5310) );
  OAI211_X1 U6822 ( .C1(n9565), .C2(n5346), .A(n5311), .B(n5310), .ZN(n9344)
         );
  NOR2_X1 U6823 ( .A1(n9654), .A2(n9344), .ZN(n5312) );
  XNOR2_X1 U6824 ( .A(n5314), .B(n5313), .ZN(n7578) );
  NAND2_X1 U6825 ( .A1(n7578), .A2(n5454), .ZN(n5318) );
  NAND2_X1 U6826 ( .A1(n5315), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5316) );
  XNOR2_X1 U6827 ( .A(n5316), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9389) );
  AOI22_X1 U6828 ( .A1(n8344), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6769), .B2(
        n9389), .ZN(n5317) );
  NOR2_X1 U6829 ( .A1(n5319), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5320) );
  OR2_X1 U6830 ( .A1(n5321), .A2(n5320), .ZN(n9310) );
  AOI22_X1 U6831 ( .A1(n6816), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n6818), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n5323) );
  NAND2_X1 U6832 ( .A1(n6817), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5322) );
  OAI211_X1 U6833 ( .C1(n9310), .C2(n5346), .A(n5323), .B(n5322), .ZN(n9577)
         );
  INV_X1 U6834 ( .A(n9577), .ZN(n9551) );
  OR2_X1 U6835 ( .A1(n9647), .A2(n9551), .ZN(n8499) );
  NAND2_X1 U6836 ( .A1(n9647), .A2(n9551), .ZN(n8365) );
  NAND2_X1 U6837 ( .A1(n8499), .A2(n8365), .ZN(n8209) );
  NAND2_X1 U6838 ( .A1(n8210), .A2(n8209), .ZN(n8211) );
  INV_X1 U6839 ( .A(n9647), .ZN(n8206) );
  XNOR2_X1 U6840 ( .A(n5326), .B(n5325), .ZN(n7743) );
  NAND2_X1 U6841 ( .A1(n7743), .A2(n5454), .ZN(n5328) );
  NAND2_X1 U6842 ( .A1(n8344), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5327) );
  NAND2_X1 U6843 ( .A1(n5330), .A2(n5329), .ZN(n5331) );
  AND2_X1 U6844 ( .A1(n5344), .A2(n5331), .ZN(n9533) );
  NAND2_X1 U6845 ( .A1(n9533), .A2(n5459), .ZN(n5337) );
  INV_X1 U6846 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n5334) );
  NAND2_X1 U6847 ( .A1(n6818), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5333) );
  NAND2_X1 U6848 ( .A1(n6817), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5332) );
  OAI211_X1 U6849 ( .C1(n5350), .C2(n5334), .A(n5333), .B(n5332), .ZN(n5335)
         );
  INV_X1 U6850 ( .A(n5335), .ZN(n5336) );
  NAND2_X1 U6851 ( .A1(n5337), .A2(n5336), .ZN(n9342) );
  XNOR2_X1 U6852 ( .A(n5341), .B(n5340), .ZN(n7818) );
  NAND2_X1 U6853 ( .A1(n7818), .A2(n5454), .ZN(n5343) );
  NAND2_X1 U6854 ( .A1(n8344), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5342) );
  NAND2_X1 U6855 ( .A1(n5344), .A2(n9246), .ZN(n5345) );
  NAND2_X1 U6856 ( .A1(n5345), .A2(n4877), .ZN(n9524) );
  OR2_X1 U6857 ( .A1(n9524), .A2(n5346), .ZN(n5353) );
  INV_X1 U6858 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n5349) );
  NAND2_X1 U6859 ( .A1(n6817), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5348) );
  NAND2_X1 U6860 ( .A1(n6818), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5347) );
  OAI211_X1 U6861 ( .C1(n5350), .C2(n5349), .A(n5348), .B(n5347), .ZN(n5351)
         );
  INV_X1 U6862 ( .A(n5351), .ZN(n5352) );
  NAND2_X1 U6863 ( .A1(n9634), .A2(n9538), .ZN(n8506) );
  NAND2_X1 U6864 ( .A1(n8511), .A2(n8506), .ZN(n9515) );
  INV_X1 U6865 ( .A(n9538), .ZN(n9341) );
  XNOR2_X1 U6866 ( .A(n5356), .B(n5355), .ZN(n7845) );
  NAND2_X1 U6867 ( .A1(n7845), .A2(n5454), .ZN(n5358) );
  NAND2_X1 U6868 ( .A1(n8344), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5357) );
  NAND2_X1 U6869 ( .A1(n6816), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5363) );
  AOI21_X1 U6870 ( .B1(n9298), .B2(n4877), .A(n5359), .ZN(n9509) );
  NAND2_X1 U6871 ( .A1(n5459), .A2(n9509), .ZN(n5362) );
  NAND2_X1 U6872 ( .A1(n5085), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5361) );
  NAND2_X1 U6873 ( .A1(n6817), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5360) );
  INV_X1 U6874 ( .A(n9522), .ZN(n9340) );
  AOI21_X1 U6875 ( .B1(n6713), .B2(n9505), .A(n9487), .ZN(n5365) );
  INV_X1 U6876 ( .A(n9505), .ZN(n9339) );
  INV_X1 U6877 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8005) );
  INV_X1 U6878 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8032) );
  MUX2_X1 U6879 ( .A(n8005), .B(n8032), .S(n5400), .Z(n5379) );
  XNOR2_X1 U6880 ( .A(n5379), .B(SI_24_), .ZN(n5378) );
  XNOR2_X1 U6881 ( .A(n5383), .B(n5378), .ZN(n8004) );
  NAND2_X1 U6882 ( .A1(n6816), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5376) );
  INV_X1 U6883 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9273) );
  INV_X1 U6884 ( .A(n5390), .ZN(n5371) );
  AOI21_X1 U6885 ( .B1(n9273), .B2(n5372), .A(n5371), .ZN(n9481) );
  NAND2_X1 U6886 ( .A1(n5459), .A2(n9481), .ZN(n5375) );
  NAND2_X1 U6887 ( .A1(n6818), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5374) );
  NAND2_X1 U6888 ( .A1(n6817), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5373) );
  INV_X1 U6889 ( .A(n9491), .ZN(n9338) );
  NAND2_X1 U6890 ( .A1(n8350), .A2(n9491), .ZN(n5377) );
  INV_X1 U6891 ( .A(n5378), .ZN(n5382) );
  INV_X1 U6892 ( .A(n5379), .ZN(n5380) );
  NAND2_X1 U6893 ( .A1(n5380), .A2(SI_24_), .ZN(n5381) );
  INV_X1 U6894 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8216) );
  INV_X1 U6895 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8217) );
  MUX2_X1 U6896 ( .A(n8216), .B(n8217), .S(n5400), .Z(n5385) );
  INV_X1 U6897 ( .A(SI_25_), .ZN(n5384) );
  NAND2_X1 U6898 ( .A1(n5385), .A2(n5384), .ZN(n5397) );
  INV_X1 U6899 ( .A(n5385), .ZN(n5386) );
  NAND2_X1 U6900 ( .A1(n5386), .A2(SI_25_), .ZN(n5387) );
  NAND2_X1 U6901 ( .A1(n5397), .A2(n5387), .ZN(n5398) );
  NAND2_X1 U6902 ( .A1(n8214), .A2(n5454), .ZN(n5389) );
  NAND2_X1 U6903 ( .A1(n8344), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5388) );
  NAND2_X1 U6904 ( .A1(n6816), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5394) );
  INV_X1 U6905 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9254) );
  AOI21_X1 U6906 ( .B1(n9254), .B2(n5390), .A(n5407), .ZN(n9461) );
  NAND2_X1 U6907 ( .A1(n5459), .A2(n9461), .ZN(n5393) );
  NAND2_X1 U6908 ( .A1(n5085), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5392) );
  NAND2_X1 U6909 ( .A1(n6817), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5391) );
  OR2_X2 U6910 ( .A1(n9612), .A2(n9477), .ZN(n8528) );
  NAND2_X1 U6911 ( .A1(n9612), .A2(n9477), .ZN(n8530) );
  NAND2_X1 U6912 ( .A1(n8528), .A2(n8530), .ZN(n9464) );
  INV_X1 U6913 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8221) );
  INV_X1 U6914 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8240) );
  MUX2_X1 U6915 ( .A(n8221), .B(n8240), .S(n5400), .Z(n5402) );
  INV_X1 U6916 ( .A(SI_26_), .ZN(n5401) );
  NAND2_X1 U6917 ( .A1(n5402), .A2(n5401), .ZN(n5415) );
  INV_X1 U6918 ( .A(n5402), .ZN(n5403) );
  NAND2_X1 U6919 ( .A1(n5403), .A2(SI_26_), .ZN(n5404) );
  XNOR2_X1 U6920 ( .A(n5414), .B(n5413), .ZN(n8220) );
  NAND2_X1 U6921 ( .A1(n8220), .A2(n5454), .ZN(n5406) );
  NAND2_X1 U6922 ( .A1(n8344), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5405) );
  NAND2_X1 U6923 ( .A1(n6816), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5412) );
  NAND2_X1 U6924 ( .A1(n5407), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5423) );
  OAI21_X1 U6925 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(n5407), .A(n5423), .ZN(
        n5408) );
  INV_X1 U6926 ( .A(n5408), .ZN(n9455) );
  NAND2_X1 U6927 ( .A1(n5459), .A2(n9455), .ZN(n5411) );
  NAND2_X1 U6928 ( .A1(n5085), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5410) );
  NAND2_X1 U6929 ( .A1(n6817), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5409) );
  OR2_X1 U6930 ( .A1(n9607), .A2(n9465), .ZN(n8349) );
  NAND2_X1 U6931 ( .A1(n9607), .A2(n9465), .ZN(n5518) );
  INV_X1 U6932 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8321) );
  INV_X1 U6933 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8245) );
  MUX2_X1 U6934 ( .A(n8321), .B(n8245), .S(n5400), .Z(n5417) );
  INV_X1 U6935 ( .A(SI_27_), .ZN(n5416) );
  NAND2_X1 U6936 ( .A1(n5417), .A2(n5416), .ZN(n5432) );
  INV_X1 U6937 ( .A(n5417), .ZN(n5418) );
  NAND2_X1 U6938 ( .A1(n5418), .A2(SI_27_), .ZN(n5419) );
  NAND2_X1 U6939 ( .A1(n8320), .A2(n5454), .ZN(n5421) );
  NAND2_X1 U6940 ( .A1(n8344), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5420) );
  NAND2_X1 U6941 ( .A1(n5085), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5429) );
  NAND2_X1 U6942 ( .A1(n6816), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5428) );
  INV_X1 U6943 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5422) );
  NAND2_X1 U6944 ( .A1(n5422), .A2(n5423), .ZN(n5425) );
  INV_X1 U6945 ( .A(n5423), .ZN(n5424) );
  NAND2_X1 U6946 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n5424), .ZN(n5458) );
  NAND2_X1 U6947 ( .A1(n5459), .A2(n9434), .ZN(n5427) );
  NAND2_X1 U6948 ( .A1(n6817), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5426) );
  NAND2_X1 U6949 ( .A1(n9601), .A2(n9450), .ZN(n8537) );
  INV_X1 U6950 ( .A(n9601), .ZN(n9436) );
  INV_X1 U6951 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8662) );
  INV_X1 U6952 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n5434) );
  MUX2_X1 U6953 ( .A(n8662), .B(n5434), .S(n5400), .Z(n5436) );
  INV_X1 U6954 ( .A(SI_28_), .ZN(n5435) );
  NAND2_X1 U6955 ( .A1(n5436), .A2(n5435), .ZN(n5448) );
  INV_X1 U6956 ( .A(n5436), .ZN(n5437) );
  NAND2_X1 U6957 ( .A1(n5437), .A2(SI_28_), .ZN(n5438) );
  NAND2_X1 U6958 ( .A1(n8309), .A2(n5454), .ZN(n5440) );
  NAND2_X1 U6959 ( .A1(n8344), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5439) );
  NAND2_X1 U6960 ( .A1(n6816), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5444) );
  NAND2_X1 U6961 ( .A1(n5085), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5443) );
  XNOR2_X1 U6962 ( .A(n5458), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n9424) );
  NAND2_X1 U6963 ( .A1(n5459), .A2(n9424), .ZN(n5442) );
  NAND2_X1 U6964 ( .A1(n6817), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5441) );
  NAND2_X1 U6965 ( .A1(n9596), .A2(n9438), .ZN(n8542) );
  NAND2_X1 U6966 ( .A1(n9596), .A2(n9335), .ZN(n5445) );
  NAND2_X1 U6967 ( .A1(n9594), .A2(n5445), .ZN(n5464) );
  INV_X1 U6968 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9705) );
  INV_X1 U6969 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n5449) );
  MUX2_X1 U6970 ( .A(n9705), .B(n5449), .S(n6799), .Z(n5451) );
  INV_X1 U6971 ( .A(SI_29_), .ZN(n5450) );
  NAND2_X1 U6972 ( .A1(n5451), .A2(n5450), .ZN(n6157) );
  INV_X1 U6973 ( .A(n5451), .ZN(n5452) );
  NAND2_X1 U6974 ( .A1(n5452), .A2(SI_29_), .ZN(n5453) );
  NAND2_X1 U6975 ( .A1(n9209), .A2(n5454), .ZN(n5456) );
  NAND2_X1 U6976 ( .A1(n8344), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n5455) );
  NAND2_X1 U6977 ( .A1(n6816), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5463) );
  NAND2_X1 U6978 ( .A1(n5085), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5462) );
  INV_X1 U6979 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5457) );
  NOR2_X1 U6980 ( .A1(n5458), .A2(n5457), .ZN(n5535) );
  NAND2_X1 U6981 ( .A1(n5459), .A2(n5535), .ZN(n5461) );
  NAND2_X1 U6982 ( .A1(n6817), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5460) );
  NAND2_X1 U6983 ( .A1(n9591), .A2(n9418), .ZN(n8633) );
  NAND2_X1 U6984 ( .A1(n8405), .A2(n8633), .ZN(n8596) );
  OAI21_X2 U6985 ( .B1(n5465), .B2(P1_IR_REG_19__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5472) );
  NAND2_X1 U6986 ( .A1(n5472), .A2(n5471), .ZN(n5466) );
  INV_X1 U6987 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5467) );
  NAND2_X1 U6988 ( .A1(n5470), .A2(n5467), .ZN(n5468) );
  XNOR2_X2 U6989 ( .A(n5469), .B(P1_IR_REG_22__SCAN_IN), .ZN(n6516) );
  NAND2_X1 U6990 ( .A1(n6516), .A2(n8640), .ZN(n6767) );
  OR2_X1 U6991 ( .A1(n6767), .A2(n8650), .ZN(n6753) );
  NAND2_X1 U6992 ( .A1(n5480), .A2(n5479), .ZN(n5482) );
  INV_X1 U6993 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5473) );
  INV_X1 U6994 ( .A(n5475), .ZN(n5476) );
  OR2_X1 U6995 ( .A1(n5480), .A2(n5479), .ZN(n5481) );
  NAND2_X1 U6996 ( .A1(n5482), .A2(n5481), .ZN(n8219) );
  INV_X1 U6997 ( .A(n5483), .ZN(n5484) );
  NAND2_X1 U6998 ( .A1(n5484), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5486) );
  XNOR2_X1 U6999 ( .A(n5486), .B(n5485), .ZN(n7954) );
  NAND2_X1 U7000 ( .A1(n6518), .A2(n7954), .ZN(n8653) );
  NAND3_X1 U7001 ( .A1(n8219), .A2(P1_B_REG_SCAN_IN), .A3(n8034), .ZN(n5487)
         );
  OAI21_X1 U7002 ( .B1(P1_B_REG_SCAN_IN), .B2(n8034), .A(n5487), .ZN(n5488) );
  INV_X1 U7003 ( .A(n8242), .ZN(n5490) );
  INV_X1 U7004 ( .A(n8034), .ZN(n5489) );
  OAI22_X1 U7005 ( .A1(n9950), .A2(P1_D_REG_0__SCAN_IN), .B1(n5490), .B2(n5489), .ZN(n6970) );
  INV_X1 U7006 ( .A(n9950), .ZN(n5501) );
  NOR4_X1 U7007 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n5499) );
  NOR4_X1 U7008 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5498) );
  INV_X1 U7009 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n9952) );
  INV_X1 U7010 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n9953) );
  INV_X1 U7011 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n9956) );
  INV_X1 U7012 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n9955) );
  NAND4_X1 U7013 ( .A1(n9952), .A2(n9953), .A3(n9956), .A4(n9955), .ZN(n5496)
         );
  NOR4_X1 U7014 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n5494) );
  NOR4_X1 U7015 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n5493) );
  NOR4_X1 U7016 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5492) );
  NOR4_X1 U7017 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n5491) );
  NAND4_X1 U7018 ( .A1(n5494), .A2(n5493), .A3(n5492), .A4(n5491), .ZN(n5495)
         );
  NOR4_X1 U7019 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        n5496), .A4(n5495), .ZN(n5497) );
  NAND3_X1 U7020 ( .A1(n5499), .A2(n5498), .A3(n5497), .ZN(n5500) );
  NAND2_X1 U7021 ( .A1(n5501), .A2(n5500), .ZN(n6912) );
  NAND2_X1 U7022 ( .A1(n6970), .A2(n6912), .ZN(n5503) );
  NAND2_X1 U7023 ( .A1(n8242), .A2(n8219), .ZN(n5502) );
  OAI21_X1 U7024 ( .B1(n9950), .B2(P1_D_REG_1__SCAN_IN), .A(n5502), .ZN(n6913)
         );
  NOR2_X1 U7025 ( .A1(n5503), .A2(n6913), .ZN(n5504) );
  NAND2_X1 U7026 ( .A1(n6895), .A2(n5504), .ZN(n7504) );
  NAND2_X1 U7027 ( .A1(n9951), .A2(n8602), .ZN(n5505) );
  OR2_X1 U7028 ( .A1(n8558), .A2(n4701), .ZN(n8659) );
  AND2_X1 U7029 ( .A1(n8659), .A2(n4311), .ZN(n9924) );
  NOR2_X1 U7030 ( .A1(n6526), .A2(n6524), .ZN(n7022) );
  NAND2_X1 U7031 ( .A1(n7134), .A2(n5084), .ZN(n5507) );
  INV_X1 U7032 ( .A(n8565), .ZN(n5508) );
  AND2_X1 U7033 ( .A1(n7344), .A2(n8420), .ZN(n8605) );
  NAND2_X1 U7034 ( .A1(n7345), .A2(n8605), .ZN(n8428) );
  AND2_X1 U7035 ( .A1(n8422), .A2(n7285), .ZN(n8427) );
  AND2_X1 U7036 ( .A1(n8427), .A2(n8610), .ZN(n8373) );
  INV_X1 U7037 ( .A(n8610), .ZN(n5509) );
  NAND2_X1 U7038 ( .A1(n5510), .A2(n8608), .ZN(n8604) );
  INV_X1 U7039 ( .A(n7396), .ZN(n8574) );
  NAND2_X1 U7040 ( .A1(n7400), .A2(n8574), .ZN(n7399) );
  INV_X1 U7041 ( .A(n8425), .ZN(n7487) );
  NOR2_X1 U7042 ( .A1(n7486), .A2(n7487), .ZN(n5511) );
  NAND2_X1 U7043 ( .A1(n7399), .A2(n5511), .ZN(n7489) );
  NAND2_X1 U7044 ( .A1(n7489), .A2(n8451), .ZN(n7586) );
  INV_X1 U7045 ( .A(n9350), .ZN(n7691) );
  OR2_X1 U7046 ( .A1(n7698), .A2(n7691), .ZN(n8454) );
  NAND2_X1 U7047 ( .A1(n7698), .A2(n7691), .ZN(n8452) );
  NAND2_X1 U7048 ( .A1(n7586), .A2(n8576), .ZN(n7591) );
  NAND2_X1 U7049 ( .A1(n7591), .A2(n8454), .ZN(n7601) );
  INV_X1 U7050 ( .A(n8578), .ZN(n7600) );
  NAND2_X1 U7051 ( .A1(n7601), .A2(n7600), .ZN(n7599) );
  NAND2_X1 U7052 ( .A1(n7599), .A2(n8466), .ZN(n7733) );
  XNOR2_X1 U7053 ( .A(n6600), .B(n9753), .ZN(n8579) );
  NAND2_X1 U7054 ( .A1(n7733), .A2(n8579), .ZN(n7732) );
  INV_X1 U7055 ( .A(n9753), .ZN(n8367) );
  OR2_X1 U7056 ( .A1(n6600), .A2(n8367), .ZN(n5512) );
  NAND2_X1 U7057 ( .A1(n7732), .A2(n5512), .ZN(n9750) );
  NAND2_X1 U7058 ( .A1(n9750), .A2(n9749), .ZN(n9748) );
  INV_X1 U7059 ( .A(n5512), .ZN(n5513) );
  NAND2_X1 U7060 ( .A1(n8486), .A2(n5513), .ZN(n5514) );
  AND2_X1 U7061 ( .A1(n5514), .A2(n8487), .ZN(n8471) );
  NAND2_X1 U7062 ( .A1(n9748), .A2(n8471), .ZN(n7898) );
  INV_X1 U7063 ( .A(n9752), .ZN(n7813) );
  OR2_X1 U7064 ( .A1(n7904), .A2(n7813), .ZN(n8470) );
  NAND2_X1 U7065 ( .A1(n7904), .A2(n7813), .ZN(n8366) );
  NAND2_X1 U7066 ( .A1(n7898), .A2(n8581), .ZN(n7897) );
  NAND2_X1 U7067 ( .A1(n7897), .A2(n8470), .ZN(n7970) );
  INV_X1 U7068 ( .A(n9347), .ZN(n7838) );
  OR2_X1 U7069 ( .A1(n9669), .A2(n7838), .ZN(n8472) );
  NAND2_X1 U7070 ( .A1(n9669), .A2(n7838), .ZN(n8387) );
  NAND2_X1 U7071 ( .A1(n7970), .A2(n8583), .ZN(n7969) );
  OR2_X1 U7072 ( .A1(n9662), .A2(n8175), .ZN(n8478) );
  NAND2_X1 U7073 ( .A1(n9662), .A2(n8175), .ZN(n8489) );
  NAND2_X1 U7074 ( .A1(n8478), .A2(n8489), .ZN(n8115) );
  INV_X1 U7075 ( .A(n8489), .ZN(n8133) );
  INV_X1 U7076 ( .A(n9344), .ZN(n5515) );
  OR2_X1 U7077 ( .A1(n9654), .A2(n5515), .ZN(n8357) );
  NAND2_X1 U7078 ( .A1(n9654), .A2(n5515), .ZN(n8364) );
  NAND2_X1 U7079 ( .A1(n8357), .A2(n8364), .ZN(n9573) );
  INV_X1 U7080 ( .A(n8357), .ZN(n5516) );
  INV_X1 U7081 ( .A(n8209), .ZN(n8588) );
  OR2_X1 U7082 ( .A1(n9644), .A2(n9537), .ZN(n8500) );
  NAND2_X1 U7083 ( .A1(n9644), .A2(n9537), .ZN(n8502) );
  INV_X1 U7084 ( .A(n8502), .ZN(n8362) );
  NAND2_X1 U7085 ( .A1(n9637), .A2(n9549), .ZN(n8501) );
  NAND2_X1 U7086 ( .A1(n9517), .A2(n8506), .ZN(n9502) );
  OR2_X1 U7087 ( .A1(n9629), .A2(n9522), .ZN(n8515) );
  NAND2_X1 U7088 ( .A1(n9629), .A2(n9522), .ZN(n8508) );
  INV_X1 U7089 ( .A(n8508), .ZN(n5517) );
  AOI21_X1 U7090 ( .B1(n9502), .B2(n9503), .A(n5517), .ZN(n9490) );
  NAND2_X1 U7091 ( .A1(n9624), .A2(n9505), .ZN(n8351) );
  NAND2_X1 U7092 ( .A1(n9490), .A2(n9489), .ZN(n9488) );
  XNOR2_X1 U7093 ( .A(n9619), .B(n9491), .ZN(n9475) );
  AND2_X1 U7094 ( .A1(n9619), .A2(n9491), .ZN(n8413) );
  NAND2_X1 U7095 ( .A1(n9467), .A2(n8528), .ZN(n9447) );
  INV_X1 U7096 ( .A(n5518), .ZN(n8347) );
  INV_X1 U7097 ( .A(n8596), .ZN(n5519) );
  NAND2_X1 U7098 ( .A1(n6516), .A2(n9497), .ZN(n5521) );
  NAND2_X1 U7099 ( .A1(n8640), .A2(n8647), .ZN(n5520) );
  INV_X1 U7100 ( .A(n6767), .ZN(n6747) );
  INV_X1 U7101 ( .A(n5522), .ZN(n6951) );
  INV_X1 U7102 ( .A(n9754), .ZN(n5531) );
  INV_X1 U7103 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n5525) );
  NAND2_X1 U7104 ( .A1(n6816), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n5524) );
  NAND2_X1 U7105 ( .A1(n6817), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5523) );
  OAI211_X1 U7106 ( .C1(n5526), .C2(n5525), .A(n5524), .B(n5523), .ZN(n9333)
         );
  INV_X1 U7107 ( .A(n9333), .ZN(n5530) );
  INV_X1 U7108 ( .A(P1_B_REG_SCAN_IN), .ZN(n5527) );
  NOR2_X1 U7109 ( .A1(n6948), .A2(n5527), .ZN(n5528) );
  NOR2_X1 U7110 ( .A1(n9550), .A2(n5528), .ZN(n9404) );
  INV_X1 U7111 ( .A(n9404), .ZN(n5529) );
  INV_X1 U7112 ( .A(n5532), .ZN(n5533) );
  INV_X2 U7113 ( .A(n9945), .ZN(n9578) );
  NOR2_X1 U7114 ( .A1(n5084), .A2(n6519), .ZN(n7133) );
  AND2_X1 U7115 ( .A1(n7133), .A2(n7368), .ZN(n7132) );
  NAND2_X1 U7116 ( .A1(n7445), .A2(n8436), .ZN(n7495) );
  OR2_X1 U7117 ( .A1(n7495), .A2(n7498), .ZN(n7583) );
  OR2_X1 U7118 ( .A1(n7583), .A2(n7698), .ZN(n7604) );
  INV_X1 U7119 ( .A(n6600), .ZN(n9783) );
  INV_X1 U7120 ( .A(n9669), .ZN(n8101) );
  NAND2_X1 U7121 ( .A1(n7973), .A2(n8101), .ZN(n8116) );
  NOR2_X2 U7122 ( .A1(n8116), .A2(n9662), .ZN(n8138) );
  INV_X1 U7123 ( .A(n5294), .ZN(n8176) );
  NAND2_X1 U7124 ( .A1(n8138), .A2(n8176), .ZN(n9564) );
  NAND2_X1 U7125 ( .A1(n9523), .A2(n9512), .ZN(n9506) );
  NAND2_X1 U7126 ( .A1(n9433), .A2(n9415), .ZN(n9414) );
  AOI21_X1 U7127 ( .B1(n9591), .B2(n9414), .A(n9408), .ZN(n9592) );
  AND2_X1 U7128 ( .A1(n8650), .A2(n7025), .ZN(n5534) );
  INV_X1 U7129 ( .A(n9591), .ZN(n5537) );
  AOI22_X1 U7130 ( .A1(n9578), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n5535), .B2(
        n9759), .ZN(n5536) );
  OAI21_X1 U7131 ( .B1(n5537), .B2(n9568), .A(n5536), .ZN(n5538) );
  AOI21_X1 U7132 ( .B1(n9592), .B2(n9940), .A(n5538), .ZN(n5539) );
  OAI211_X1 U7133 ( .C1(n9593), .C2(n9582), .A(n4318), .B(n5539), .ZN(P1_U3355) );
  NOR2_X1 U7134 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5549) );
  NOR2_X1 U7135 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5548) );
  INV_X1 U7136 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5551) );
  INV_X1 U7137 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5554) );
  NAND2_X1 U7138 ( .A1(n5648), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5563) );
  INV_X1 U7139 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10108) );
  INV_X1 U7140 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7032) );
  INV_X1 U7141 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7111) );
  NAND4_X2 U7142 ( .A1(n5563), .A2(n5562), .A3(n5561), .A4(n5560), .ZN(n8861)
         );
  NAND2_X1 U7143 ( .A1(n5569), .A2(n5564), .ZN(n5567) );
  INV_X1 U7144 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5565) );
  NAND2_X1 U7145 ( .A1(n5567), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5568) );
  AND2_X2 U7146 ( .A1(n7847), .A2(n7820), .ZN(n10046) );
  INV_X1 U7147 ( .A(n5569), .ZN(n5570) );
  NAND2_X1 U7148 ( .A1(n5570), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5574) );
  INV_X1 U7149 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5573) );
  NAND2_X1 U7150 ( .A1(n5574), .A2(n5573), .ZN(n5576) );
  INV_X1 U7151 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5571) );
  OR2_X1 U7152 ( .A1(n5574), .A2(n5573), .ZN(n5575) );
  INV_X1 U7153 ( .A(n5590), .ZN(n5588) );
  INV_X1 U7154 ( .A(n5577), .ZN(n5578) );
  NAND2_X1 U7155 ( .A1(n4328), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5580) );
  MUX2_X1 U7156 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5580), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5583) );
  INV_X1 U7157 ( .A(n5581), .ZN(n5582) );
  NAND2_X1 U7158 ( .A1(n5863), .A2(n7033), .ZN(n5584) );
  NAND2_X1 U7159 ( .A1(n7820), .A2(n8974), .ZN(n5586) );
  AND3_X4 U7160 ( .A1(n6374), .A2(n7331), .A3(n5586), .ZN(n6032) );
  INV_X1 U7161 ( .A(n5589), .ZN(n5587) );
  NAND2_X1 U7162 ( .A1(n5588), .A2(n5587), .ZN(n5600) );
  NAND2_X1 U7163 ( .A1(n5590), .A2(n5589), .ZN(n5591) );
  NAND2_X1 U7164 ( .A1(n6166), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5594) );
  INV_X1 U7165 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10106) );
  INV_X1 U7166 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5592) );
  OR2_X1 U7167 ( .A1(n6175), .A2(n5592), .ZN(n5593) );
  NAND2_X1 U7168 ( .A1(n8863), .A2(n6196), .ZN(n5599) );
  INV_X1 U7169 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10016) );
  NAND2_X1 U7170 ( .A1(n6799), .A2(SI_0_), .ZN(n5596) );
  INV_X1 U7171 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5595) );
  NAND2_X1 U7172 ( .A1(n5596), .A2(n5595), .ZN(n5598) );
  NAND2_X1 U7173 ( .A1(n5598), .A2(n5597), .ZN(n9213) );
  MUX2_X1 U7174 ( .A(n10016), .B(n9213), .S(n5707), .Z(n7467) );
  NAND2_X1 U7175 ( .A1(n7106), .A2(n7107), .ZN(n7105) );
  NAND2_X1 U7176 ( .A1(n6166), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5605) );
  INV_X1 U7177 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10110) );
  INV_X1 U7178 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5601) );
  INV_X1 U7179 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n8705) );
  AND2_X1 U7180 ( .A1(n6115), .A2(n6196), .ZN(n5612) );
  NOR2_X1 U7181 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5608) );
  INV_X1 U7182 ( .A(n5608), .ZN(n5606) );
  NAND2_X1 U7183 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5606), .ZN(n5607) );
  INV_X1 U7184 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6478) );
  MUX2_X1 U7185 ( .A(n5607), .B(P2_IR_REG_31__SCAN_IN), .S(n6478), .Z(n5609)
         );
  NAND2_X1 U7186 ( .A1(n6478), .A2(n5608), .ZN(n5618) );
  AND2_X1 U7187 ( .A1(n5609), .A2(n5618), .ZN(n9730) );
  NAND2_X1 U7188 ( .A1(n5863), .A2(n9730), .ZN(n5610) );
  XNOR2_X1 U7189 ( .A(n6116), .B(n6032), .ZN(n5613) );
  NAND2_X1 U7190 ( .A1(n5612), .A2(n5613), .ZN(n5616) );
  INV_X1 U7191 ( .A(n5612), .ZN(n5615) );
  INV_X1 U7192 ( .A(n5613), .ZN(n5614) );
  NAND2_X1 U7193 ( .A1(n5615), .A2(n5614), .ZN(n5617) );
  AND2_X1 U7194 ( .A1(n5616), .A2(n5617), .ZN(n7235) );
  NAND2_X1 U7195 ( .A1(n6189), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5621) );
  NAND2_X1 U7196 ( .A1(n5618), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5619) );
  XNOR2_X1 U7197 ( .A(n5619), .B(P2_IR_REG_3__SCAN_IN), .ZN(n7049) );
  NAND2_X1 U7198 ( .A1(n5863), .A2(n7049), .ZN(n5620) );
  OAI211_X1 U7199 ( .C1(n6801), .C2(n5685), .A(n5621), .B(n5620), .ZN(n6119)
         );
  XNOR2_X1 U7200 ( .A(n6119), .B(n6057), .ZN(n5629) );
  NAND2_X1 U7201 ( .A1(n5622), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5625) );
  INV_X1 U7202 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5623) );
  OR2_X1 U7203 ( .A1(n6175), .A2(n5623), .ZN(n5624) );
  OR2_X1 U7204 ( .A1(n6018), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5627) );
  INV_X1 U7205 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7050) );
  NAND2_X1 U7206 ( .A1(n8860), .A2(n7336), .ZN(n5628) );
  XNOR2_X1 U7207 ( .A(n5629), .B(n5628), .ZN(n7224) );
  NAND2_X1 U7208 ( .A1(n5648), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5637) );
  INV_X1 U7209 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7048) );
  OR2_X1 U7210 ( .A1(n6173), .A2(n7048), .ZN(n5636) );
  INV_X1 U7211 ( .A(n5649), .ZN(n5632) );
  INV_X1 U7212 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7229) );
  INV_X1 U7213 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5630) );
  NAND2_X1 U7214 ( .A1(n7229), .A2(n5630), .ZN(n5631) );
  NAND2_X1 U7215 ( .A1(n5632), .A2(n5631), .ZN(n7314) );
  OR2_X1 U7216 ( .A1(n6018), .A2(n7314), .ZN(n5635) );
  INV_X1 U7217 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n5633) );
  OR2_X1 U7218 ( .A1(n5956), .A2(n5633), .ZN(n5634) );
  AND2_X1 U7219 ( .A1(n8859), .A2(n7336), .ZN(n5642) );
  NAND2_X1 U7220 ( .A1(n6189), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5641) );
  OR2_X1 U7221 ( .A1(n5638), .A2(n5554), .ZN(n5639) );
  XNOR2_X1 U7222 ( .A(n5639), .B(P2_IR_REG_4__SCAN_IN), .ZN(n7047) );
  NAND2_X1 U7223 ( .A1(n5863), .A2(n7047), .ZN(n5640) );
  XNOR2_X1 U7224 ( .A(n7756), .B(n6032), .ZN(n5643) );
  NAND2_X1 U7225 ( .A1(n5642), .A2(n5643), .ZN(n5646) );
  INV_X1 U7226 ( .A(n5642), .ZN(n5645) );
  INV_X1 U7227 ( .A(n5643), .ZN(n5644) );
  NAND2_X1 U7228 ( .A1(n5645), .A2(n5644), .ZN(n5647) );
  NAND2_X1 U7229 ( .A1(n5646), .A2(n5647), .ZN(n7313) );
  NAND2_X1 U7230 ( .A1(n7310), .A2(n5647), .ZN(n7388) );
  NAND2_X1 U7231 ( .A1(n5648), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5654) );
  INV_X1 U7232 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7054) );
  OR2_X1 U7233 ( .A1(n6173), .A2(n7054), .ZN(n5653) );
  NAND2_X1 U7234 ( .A1(n5649), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5668) );
  OAI21_X1 U7235 ( .B1(n5649), .B2(P2_REG3_REG_5__SCAN_IN), .A(n5668), .ZN(
        n10024) );
  OR2_X1 U7236 ( .A1(n6018), .A2(n10024), .ZN(n5652) );
  INV_X1 U7237 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n5650) );
  OR2_X1 U7238 ( .A1(n5956), .A2(n5650), .ZN(n5651) );
  NAND4_X1 U7239 ( .A1(n5654), .A2(n5653), .A3(n5652), .A4(n5651), .ZN(n8858)
         );
  AND2_X1 U7240 ( .A1(n8858), .A2(n7336), .ZN(n5661) );
  NAND2_X1 U7241 ( .A1(n6189), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5660) );
  NAND2_X1 U7242 ( .A1(n5655), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5657) );
  NAND2_X1 U7243 ( .A1(n5657), .A2(n5656), .ZN(n5674) );
  OR2_X1 U7244 ( .A1(n5657), .A2(n5656), .ZN(n5658) );
  NAND2_X1 U7245 ( .A1(n5863), .A2(n7091), .ZN(n5659) );
  XNOR2_X1 U7246 ( .A(n10022), .B(n6032), .ZN(n5662) );
  NAND2_X1 U7247 ( .A1(n5661), .A2(n5662), .ZN(n5665) );
  INV_X1 U7248 ( .A(n5661), .ZN(n5664) );
  INV_X1 U7249 ( .A(n5662), .ZN(n5663) );
  NAND2_X1 U7250 ( .A1(n5664), .A2(n5663), .ZN(n5666) );
  AND2_X1 U7251 ( .A1(n5665), .A2(n5666), .ZN(n7389) );
  NAND2_X1 U7252 ( .A1(n7388), .A2(n7389), .ZN(n7387) );
  NAND2_X1 U7253 ( .A1(n7387), .A2(n5666), .ZN(n7476) );
  NAND2_X1 U7254 ( .A1(n5648), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5673) );
  INV_X1 U7255 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7094) );
  OR2_X1 U7256 ( .A1(n6173), .A2(n7094), .ZN(n5672) );
  AND2_X1 U7257 ( .A1(n5668), .A2(n5667), .ZN(n5669) );
  OR2_X1 U7258 ( .A1(n5669), .A2(n5694), .ZN(n7635) );
  OR2_X1 U7259 ( .A1(n6018), .A2(n7635), .ZN(n5671) );
  INV_X1 U7260 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7636) );
  OR2_X1 U7261 ( .A1(n5956), .A2(n7636), .ZN(n5670) );
  NAND4_X1 U7262 ( .A1(n5673), .A2(n5672), .A3(n5671), .A4(n5670), .ZN(n8857)
         );
  AND2_X1 U7263 ( .A1(n8857), .A2(n7336), .ZN(n5678) );
  NAND2_X1 U7264 ( .A1(n6189), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n5677) );
  NAND2_X1 U7265 ( .A1(n5674), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5675) );
  XNOR2_X1 U7266 ( .A(n5675), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7121) );
  NAND2_X1 U7267 ( .A1(n5863), .A2(n7121), .ZN(n5676) );
  OAI211_X1 U7268 ( .C1(n6805), .C2(n5685), .A(n5677), .B(n5676), .ZN(n7640)
         );
  XNOR2_X1 U7269 ( .A(n7640), .B(n6032), .ZN(n5679) );
  NAND2_X1 U7270 ( .A1(n5678), .A2(n5679), .ZN(n5682) );
  INV_X1 U7271 ( .A(n5678), .ZN(n5681) );
  INV_X1 U7272 ( .A(n5679), .ZN(n5680) );
  NAND2_X1 U7273 ( .A1(n5681), .A2(n5680), .ZN(n5683) );
  AND2_X1 U7274 ( .A1(n5682), .A2(n5683), .ZN(n7477) );
  INV_X1 U7275 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6815) );
  NAND2_X1 U7276 ( .A1(n6188), .A2(n6812), .ZN(n5692) );
  NAND2_X1 U7277 ( .A1(n5686), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5688) );
  MUX2_X1 U7278 ( .A(n5688), .B(P2_IR_REG_31__SCAN_IN), .S(n5687), .Z(n5690)
         );
  NOR2_X1 U7279 ( .A1(n5686), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5711) );
  INV_X1 U7280 ( .A(n5711), .ZN(n5689) );
  NAND2_X1 U7281 ( .A1(n5690), .A2(n5689), .ZN(n7127) );
  INV_X1 U7282 ( .A(n7127), .ZN(n7148) );
  NAND2_X1 U7283 ( .A1(n5863), .A2(n7148), .ZN(n5691) );
  OAI211_X1 U7284 ( .C1(n5917), .C2(n6815), .A(n5692), .B(n5691), .ZN(n7822)
         );
  XNOR2_X1 U7285 ( .A(n7822), .B(n6057), .ZN(n5702) );
  NAND2_X1 U7286 ( .A1(n5980), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5700) );
  INV_X1 U7287 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n5693) );
  OR2_X1 U7288 ( .A1(n5956), .A2(n5693), .ZN(n5699) );
  NAND2_X1 U7289 ( .A1(n5694), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5719) );
  OR2_X1 U7290 ( .A1(n5694), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5695) );
  NAND2_X1 U7291 ( .A1(n5719), .A2(n5695), .ZN(n7515) );
  OR2_X1 U7292 ( .A1(n6018), .A2(n7515), .ZN(n5698) );
  INV_X1 U7293 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n5696) );
  OR2_X1 U7294 ( .A1(n6175), .A2(n5696), .ZN(n5697) );
  NAND4_X1 U7295 ( .A1(n5700), .A2(n5699), .A3(n5698), .A4(n5697), .ZN(n9997)
         );
  NAND2_X1 U7296 ( .A1(n9997), .A2(n7336), .ZN(n5701) );
  XNOR2_X1 U7297 ( .A(n5702), .B(n5701), .ZN(n7514) );
  INV_X1 U7298 ( .A(n5701), .ZN(n5704) );
  INV_X1 U7299 ( .A(n5702), .ZN(n5703) );
  NAND2_X1 U7300 ( .A1(n5704), .A2(n5703), .ZN(n5705) );
  NAND2_X1 U7301 ( .A1(n5706), .A2(n5705), .ZN(n9992) );
  NOR2_X1 U7302 ( .A1(n5711), .A2(n5554), .ZN(n5708) );
  MUX2_X1 U7303 ( .A(n5554), .B(n5708), .S(P2_IR_REG_8__SCAN_IN), .Z(n5709) );
  INV_X1 U7304 ( .A(n5709), .ZN(n5713) );
  INV_X1 U7305 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5710) );
  INV_X1 U7306 ( .A(n5747), .ZN(n5712) );
  INV_X1 U7307 ( .A(n7180), .ZN(n6825) );
  OAI22_X1 U7308 ( .A1(n5917), .A2(n6827), .B1(n5805), .B2(n6825), .ZN(n5714)
         );
  INV_X1 U7309 ( .A(n5714), .ZN(n5715) );
  XNOR2_X1 U7310 ( .A(n7851), .B(n6032), .ZN(n5727) );
  NAND2_X1 U7311 ( .A1(n6166), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5724) );
  INV_X1 U7312 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n5716) );
  OR2_X1 U7313 ( .A1(n6173), .A2(n5716), .ZN(n5723) );
  INV_X1 U7314 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5717) );
  OR2_X1 U7315 ( .A1(n6175), .A2(n5717), .ZN(n5722) );
  NAND2_X1 U7316 ( .A1(n5719), .A2(n5718), .ZN(n5720) );
  NAND2_X1 U7317 ( .A1(n5736), .A2(n5720), .ZN(n10005) );
  OR2_X1 U7318 ( .A1(n6018), .A2(n10005), .ZN(n5721) );
  NAND2_X1 U7319 ( .A1(n8856), .A2(n7336), .ZN(n5725) );
  XNOR2_X1 U7320 ( .A(n5727), .B(n5725), .ZN(n9991) );
  NAND2_X1 U7321 ( .A1(n9992), .A2(n9991), .ZN(n5729) );
  INV_X1 U7322 ( .A(n5725), .ZN(n5726) );
  NAND2_X1 U7323 ( .A1(n5727), .A2(n5726), .ZN(n5728) );
  NAND2_X1 U7324 ( .A1(n5729), .A2(n5728), .ZN(n6781) );
  NAND2_X1 U7325 ( .A1(n6830), .A2(n6188), .ZN(n5733) );
  OR2_X1 U7326 ( .A1(n5747), .A2(n5554), .ZN(n5730) );
  XNOR2_X1 U7327 ( .A(n5730), .B(n5746), .ZN(n7272) );
  OAI22_X1 U7328 ( .A1(n5917), .A2(n6870), .B1(n5805), .B2(n7272), .ZN(n5731)
         );
  INV_X1 U7329 ( .A(n5731), .ZN(n5732) );
  XNOR2_X1 U7330 ( .A(n7957), .B(n6057), .ZN(n5742) );
  NAND2_X1 U7331 ( .A1(n5648), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5741) );
  INV_X1 U7332 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7271) );
  OR2_X1 U7333 ( .A1(n6173), .A2(n7271), .ZN(n5740) );
  INV_X1 U7334 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n5734) );
  OR2_X1 U7335 ( .A1(n5956), .A2(n5734), .ZN(n5739) );
  INV_X1 U7336 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6786) );
  NAND2_X1 U7337 ( .A1(n5736), .A2(n6786), .ZN(n5737) );
  NAND2_X1 U7338 ( .A1(n5775), .A2(n5737), .ZN(n7867) );
  OR2_X1 U7339 ( .A1(n6018), .A2(n7867), .ZN(n5738) );
  NAND4_X1 U7340 ( .A1(n5741), .A2(n5740), .A3(n5739), .A4(n5738), .ZN(n8855)
         );
  NAND2_X1 U7341 ( .A1(n8855), .A2(n7336), .ZN(n5743) );
  NAND2_X1 U7342 ( .A1(n5742), .A2(n5743), .ZN(n6782) );
  NAND2_X1 U7343 ( .A1(n6781), .A2(n6782), .ZN(n6780) );
  INV_X1 U7344 ( .A(n5742), .ZN(n5745) );
  INV_X1 U7345 ( .A(n5743), .ZN(n5744) );
  NAND2_X1 U7346 ( .A1(n5745), .A2(n5744), .ZN(n6784) );
  NAND2_X1 U7347 ( .A1(n6780), .A2(n6784), .ZN(n6773) );
  NAND2_X1 U7348 ( .A1(n6872), .A2(n6188), .ZN(n5754) );
  NOR2_X1 U7349 ( .A1(n5786), .A2(n5554), .ZN(n5748) );
  NAND2_X1 U7350 ( .A1(n5748), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n5751) );
  INV_X1 U7351 ( .A(n5748), .ZN(n5750) );
  NAND2_X1 U7352 ( .A1(n5750), .A2(n5749), .ZN(n5766) );
  INV_X1 U7353 ( .A(n7268), .ZN(n8865) );
  OAI22_X1 U7354 ( .A1(n5917), .A2(n6875), .B1(n5805), .B2(n8865), .ZN(n5752)
         );
  INV_X1 U7355 ( .A(n5752), .ZN(n5753) );
  NAND2_X1 U7356 ( .A1(n5754), .A2(n5753), .ZN(n7986) );
  XNOR2_X1 U7357 ( .A(n7986), .B(n6032), .ZN(n5762) );
  NAND2_X1 U7358 ( .A1(n6166), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5759) );
  INV_X1 U7359 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7269) );
  OR2_X1 U7360 ( .A1(n6173), .A2(n7269), .ZN(n5758) );
  INV_X1 U7361 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5755) );
  OR2_X1 U7362 ( .A1(n6175), .A2(n5755), .ZN(n5757) );
  INV_X1 U7363 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5773) );
  XNOR2_X1 U7364 ( .A(n5775), .B(n5773), .ZN(n7887) );
  OR2_X1 U7365 ( .A1(n6018), .A2(n7887), .ZN(n5756) );
  NAND4_X1 U7366 ( .A1(n5759), .A2(n5758), .A3(n5757), .A4(n5756), .ZN(n8854)
         );
  NAND2_X1 U7367 ( .A1(n8854), .A2(n7336), .ZN(n5760) );
  XNOR2_X1 U7368 ( .A(n5762), .B(n5760), .ZN(n6772) );
  NAND2_X1 U7369 ( .A1(n6773), .A2(n6772), .ZN(n5764) );
  INV_X1 U7370 ( .A(n5760), .ZN(n5761) );
  NAND2_X1 U7371 ( .A1(n5762), .A2(n5761), .ZN(n5763) );
  NAND2_X1 U7372 ( .A1(n5764), .A2(n5763), .ZN(n5781) );
  NAND2_X1 U7373 ( .A1(n5765), .A2(n6188), .ZN(n5771) );
  NAND2_X1 U7374 ( .A1(n5766), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5768) );
  INV_X1 U7375 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5767) );
  XNOR2_X1 U7376 ( .A(n5768), .B(n5767), .ZN(n7530) );
  OAI22_X1 U7377 ( .A1(n5917), .A2(n6889), .B1(n5805), .B2(n7530), .ZN(n5769)
         );
  INV_X1 U7378 ( .A(n5769), .ZN(n5770) );
  XNOR2_X1 U7379 ( .A(n8040), .B(n6032), .ZN(n5782) );
  NAND2_X1 U7380 ( .A1(n5781), .A2(n5782), .ZN(n8035) );
  NAND2_X1 U7381 ( .A1(n5648), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5780) );
  INV_X1 U7382 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7273) );
  OR2_X1 U7383 ( .A1(n6173), .A2(n7273), .ZN(n5779) );
  INV_X1 U7384 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n8016) );
  OR2_X1 U7385 ( .A1(n5956), .A2(n8016), .ZN(n5778) );
  INV_X1 U7386 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5772) );
  OAI21_X1 U7387 ( .B1(n5775), .B2(n5773), .A(n5772), .ZN(n5776) );
  NAND2_X1 U7388 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_REG3_REG_11__SCAN_IN), 
        .ZN(n5774) );
  OR2_X2 U7389 ( .A1(n5775), .A2(n5774), .ZN(n5792) );
  NAND2_X1 U7390 ( .A1(n5776), .A2(n5792), .ZN(n8043) );
  OR2_X1 U7391 ( .A1(n6018), .A2(n8043), .ZN(n5777) );
  NAND4_X1 U7392 ( .A1(n5780), .A2(n5779), .A3(n5778), .A4(n5777), .ZN(n8853)
         );
  NAND2_X1 U7393 ( .A1(n8853), .A2(n7336), .ZN(n8038) );
  NAND2_X1 U7394 ( .A1(n6999), .A2(n6188), .ZN(n5790) );
  NOR2_X1 U7395 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5785) );
  NAND2_X1 U7396 ( .A1(n5786), .A2(n5785), .ZN(n5806) );
  NAND2_X1 U7397 ( .A1(n5806), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5787) );
  XNOR2_X1 U7398 ( .A(n5787), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7650) );
  INV_X1 U7399 ( .A(n7650), .ZN(n7645) );
  OAI22_X1 U7400 ( .A1(n5917), .A2(n7000), .B1(n5805), .B2(n7645), .ZN(n5788)
         );
  INV_X1 U7401 ( .A(n5788), .ZN(n5789) );
  XNOR2_X1 U7402 ( .A(n8083), .B(n6057), .ZN(n5799) );
  NAND2_X1 U7403 ( .A1(n5648), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5797) );
  INV_X1 U7404 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7523) );
  OR2_X1 U7405 ( .A1(n6173), .A2(n7523), .ZN(n5796) );
  INV_X1 U7406 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8081) );
  OR2_X1 U7407 ( .A1(n5956), .A2(n8081), .ZN(n5795) );
  INV_X1 U7408 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7526) );
  NAND2_X1 U7409 ( .A1(n5792), .A2(n7526), .ZN(n5793) );
  NAND2_X1 U7410 ( .A1(n5831), .A2(n5793), .ZN(n8080) );
  OR2_X1 U7411 ( .A1(n6018), .A2(n8080), .ZN(n5794) );
  NAND4_X1 U7412 ( .A1(n5797), .A2(n5796), .A3(n5795), .A4(n5794), .ZN(n8852)
         );
  NAND2_X1 U7413 ( .A1(n8852), .A2(n7336), .ZN(n5800) );
  XNOR2_X1 U7414 ( .A(n5799), .B(n5800), .ZN(n8048) );
  INV_X1 U7415 ( .A(n8048), .ZN(n5798) );
  INV_X1 U7416 ( .A(n5799), .ZN(n5802) );
  INV_X1 U7417 ( .A(n5800), .ZN(n5801) );
  NAND2_X1 U7418 ( .A1(n5802), .A2(n5801), .ZN(n5803) );
  NAND2_X1 U7419 ( .A1(n5804), .A2(n5803), .ZN(n8146) );
  NAND2_X1 U7420 ( .A1(n7112), .A2(n6188), .ZN(n5810) );
  NAND2_X1 U7421 ( .A1(n5807), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5822) );
  XNOR2_X1 U7422 ( .A(n5822), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7783) );
  INV_X1 U7423 ( .A(n7783), .ZN(n7646) );
  OAI22_X1 U7424 ( .A1(n5917), .A2(n7113), .B1(n5805), .B2(n7646), .ZN(n5808)
         );
  INV_X1 U7425 ( .A(n5808), .ZN(n5809) );
  XNOR2_X1 U7426 ( .A(n9179), .B(n6032), .ZN(n5818) );
  NAND2_X1 U7427 ( .A1(n5648), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5815) );
  INV_X1 U7428 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5811) );
  OR2_X1 U7429 ( .A1(n6173), .A2(n5811), .ZN(n5814) );
  INV_X1 U7430 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7998) );
  OR2_X1 U7431 ( .A1(n5956), .A2(n7998), .ZN(n5813) );
  XNOR2_X1 U7432 ( .A(n5831), .B(n7655), .ZN(n8149) );
  OR2_X1 U7433 ( .A1(n6018), .A2(n8149), .ZN(n5812) );
  NAND4_X1 U7434 ( .A1(n5815), .A2(n5814), .A3(n5813), .A4(n5812), .ZN(n8851)
         );
  NAND2_X1 U7435 ( .A1(n8851), .A2(n7336), .ZN(n5816) );
  XNOR2_X1 U7436 ( .A(n5818), .B(n5816), .ZN(n8145) );
  NAND2_X1 U7437 ( .A1(n8146), .A2(n8145), .ZN(n5820) );
  INV_X1 U7438 ( .A(n5816), .ZN(n5817) );
  NAND2_X1 U7439 ( .A1(n5818), .A2(n5817), .ZN(n5819) );
  NAND2_X1 U7440 ( .A1(n7157), .A2(n6188), .ZN(n5829) );
  AOI21_X1 U7441 ( .B1(n5822), .B2(n5821), .A(n5554), .ZN(n5823) );
  NAND2_X1 U7442 ( .A1(n5823), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n5826) );
  INV_X1 U7443 ( .A(n5823), .ZN(n5825) );
  INV_X1 U7444 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5824) );
  NAND2_X1 U7445 ( .A1(n5825), .A2(n5824), .ZN(n5861) );
  INV_X1 U7446 ( .A(n7940), .ZN(n7943) );
  OAI22_X1 U7447 ( .A1(n5917), .A2(n7158), .B1(n5805), .B2(n7943), .ZN(n5827)
         );
  INV_X1 U7448 ( .A(n5827), .ZN(n5828) );
  XNOR2_X1 U7449 ( .A(n8264), .B(n6057), .ZN(n5838) );
  NAND2_X1 U7450 ( .A1(n6166), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5837) );
  INV_X1 U7451 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5830) );
  OAI21_X1 U7452 ( .B1(n5831), .B2(n7655), .A(n5830), .ZN(n5832) );
  NAND2_X1 U7453 ( .A1(n5832), .A2(n5867), .ZN(n8262) );
  OR2_X1 U7454 ( .A1(n6018), .A2(n8262), .ZN(n5836) );
  INV_X1 U7455 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7779) );
  OR2_X1 U7456 ( .A1(n6173), .A2(n7779), .ZN(n5835) );
  INV_X1 U7457 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n5833) );
  OR2_X1 U7458 ( .A1(n6175), .A2(n5833), .ZN(n5834) );
  NAND4_X1 U7459 ( .A1(n5837), .A2(n5836), .A3(n5835), .A4(n5834), .ZN(n8850)
         );
  NAND2_X1 U7460 ( .A1(n8850), .A2(n7336), .ZN(n5839) );
  NAND2_X1 U7461 ( .A1(n5838), .A2(n5839), .ZN(n5843) );
  INV_X1 U7462 ( .A(n5838), .ZN(n5841) );
  INV_X1 U7463 ( .A(n5839), .ZN(n5840) );
  NAND2_X1 U7464 ( .A1(n5841), .A2(n5840), .ZN(n5842) );
  NAND2_X1 U7465 ( .A1(n5843), .A2(n5842), .ZN(n8258) );
  NAND2_X1 U7466 ( .A1(n7240), .A2(n6188), .ZN(n5851) );
  NOR2_X1 U7467 ( .A1(n5844), .A2(n5554), .ZN(n5845) );
  MUX2_X1 U7468 ( .A(n5554), .B(n5845), .S(P2_IR_REG_16__SCAN_IN), .Z(n5846)
         );
  INV_X1 U7469 ( .A(n5846), .ZN(n5848) );
  AND2_X1 U7470 ( .A1(n5848), .A2(n5847), .ZN(n8271) );
  INV_X1 U7471 ( .A(n8271), .ZN(n7308) );
  OAI22_X1 U7472 ( .A1(n5917), .A2(n7309), .B1(n5805), .B2(n7308), .ZN(n5849)
         );
  INV_X1 U7473 ( .A(n5849), .ZN(n5850) );
  XNOR2_X1 U7474 ( .A(n9172), .B(n6057), .ZN(n5877) );
  NAND2_X1 U7475 ( .A1(n6166), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5860) );
  INV_X1 U7476 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n5852) );
  OR2_X1 U7477 ( .A1(n6173), .A2(n5852), .ZN(n5859) );
  NAND2_X1 U7478 ( .A1(n5853), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5889) );
  INV_X1 U7479 ( .A(n5853), .ZN(n5869) );
  INV_X1 U7480 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5854) );
  NAND2_X1 U7481 ( .A1(n5869), .A2(n5854), .ZN(n5855) );
  NAND2_X1 U7482 ( .A1(n5889), .A2(n5855), .ZN(n8769) );
  OR2_X1 U7483 ( .A1(n6018), .A2(n8769), .ZN(n5858) );
  INV_X1 U7484 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n5856) );
  OR2_X1 U7485 ( .A1(n6175), .A2(n5856), .ZN(n5857) );
  NAND4_X1 U7486 ( .A1(n5860), .A2(n5859), .A3(n5858), .A4(n5857), .ZN(n8848)
         );
  NAND2_X1 U7487 ( .A1(n8848), .A2(n7336), .ZN(n5878) );
  NAND2_X1 U7488 ( .A1(n5877), .A2(n5878), .ZN(n8760) );
  NAND2_X1 U7489 ( .A1(n7258), .A2(n6188), .ZN(n5865) );
  NAND2_X1 U7490 ( .A1(n5861), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5862) );
  XNOR2_X1 U7491 ( .A(n5862), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8183) );
  AOI22_X1 U7492 ( .A1(n6189), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5863), .B2(
        n8183), .ZN(n5864) );
  XNOR2_X1 U7493 ( .A(n8833), .B(n6032), .ZN(n5875) );
  INV_X1 U7494 ( .A(n5875), .ZN(n8762) );
  NAND2_X1 U7495 ( .A1(n5648), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5873) );
  INV_X1 U7496 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n5866) );
  OR2_X1 U7497 ( .A1(n6173), .A2(n5866), .ZN(n5872) );
  INV_X1 U7498 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8164) );
  OR2_X1 U7499 ( .A1(n5956), .A2(n8164), .ZN(n5871) );
  NAND2_X1 U7500 ( .A1(n5867), .A2(n8827), .ZN(n5868) );
  NAND2_X1 U7501 ( .A1(n5869), .A2(n5868), .ZN(n8831) );
  OR2_X1 U7502 ( .A1(n6018), .A2(n8831), .ZN(n5870) );
  NAND4_X1 U7503 ( .A1(n5873), .A2(n5872), .A3(n5871), .A4(n5870), .ZN(n8849)
         );
  AND2_X1 U7504 ( .A1(n8849), .A2(n7336), .ZN(n5876) );
  INV_X1 U7505 ( .A(n5876), .ZN(n8825) );
  NAND2_X1 U7506 ( .A1(n8762), .A2(n8825), .ZN(n5874) );
  NAND2_X1 U7507 ( .A1(n8760), .A2(n5874), .ZN(n5883) );
  NAND3_X1 U7508 ( .A1(n8760), .A2(n5876), .A3(n5875), .ZN(n5881) );
  INV_X1 U7509 ( .A(n5877), .ZN(n5880) );
  INV_X1 U7510 ( .A(n5878), .ZN(n5879) );
  NAND2_X1 U7511 ( .A1(n5880), .A2(n5879), .ZN(n8759) );
  NAND2_X1 U7512 ( .A1(n7340), .A2(n6188), .ZN(n5888) );
  NAND2_X1 U7513 ( .A1(n5847), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5884) );
  MUX2_X1 U7514 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5884), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n5885) );
  AND2_X1 U7515 ( .A1(n5885), .A2(n4329), .ZN(n8885) );
  INV_X1 U7516 ( .A(n8885), .ZN(n8880) );
  OAI22_X1 U7517 ( .A1(n5917), .A2(n7341), .B1(n5805), .B2(n8880), .ZN(n5886)
         );
  INV_X1 U7518 ( .A(n5886), .ZN(n5887) );
  XNOR2_X1 U7519 ( .A(n9167), .B(n6032), .ZN(n5897) );
  NAND2_X1 U7520 ( .A1(n5648), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5894) );
  INV_X1 U7521 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8881) );
  OR2_X1 U7522 ( .A1(n6173), .A2(n8881), .ZN(n5893) );
  INV_X1 U7523 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8313) );
  NAND2_X1 U7524 ( .A1(n5889), .A2(n8313), .ZN(n5890) );
  NAND2_X1 U7525 ( .A1(n5906), .A2(n5890), .ZN(n8316) );
  OR2_X1 U7526 ( .A1(n6018), .A2(n8316), .ZN(n5892) );
  INV_X1 U7527 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8293) );
  OR2_X1 U7528 ( .A1(n5956), .A2(n8293), .ZN(n5891) );
  NAND4_X1 U7529 ( .A1(n5894), .A2(n5893), .A3(n5892), .A4(n5891), .ZN(n8847)
         );
  NAND2_X1 U7530 ( .A1(n8847), .A2(n7336), .ZN(n5895) );
  XNOR2_X1 U7531 ( .A(n5897), .B(n5895), .ZN(n8311) );
  NAND2_X1 U7532 ( .A1(n8312), .A2(n8311), .ZN(n5899) );
  INV_X1 U7533 ( .A(n5895), .ZN(n5896) );
  NAND2_X1 U7534 ( .A1(n5897), .A2(n5896), .ZN(n5898) );
  NAND2_X1 U7535 ( .A1(n5899), .A2(n5898), .ZN(n8805) );
  NAND2_X1 U7536 ( .A1(n7578), .A2(n6188), .ZN(n5903) );
  INV_X1 U7537 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7581) );
  NAND2_X1 U7538 ( .A1(n4329), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5900) );
  XNOR2_X1 U7539 ( .A(n5900), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8890) );
  INV_X1 U7540 ( .A(n8890), .ZN(n8900) );
  OAI22_X1 U7541 ( .A1(n5917), .A2(n7581), .B1(n5805), .B2(n8900), .ZN(n5901)
         );
  INV_X1 U7542 ( .A(n5901), .ZN(n5902) );
  XNOR2_X1 U7543 ( .A(n9161), .B(n6032), .ZN(n5914) );
  NAND2_X1 U7544 ( .A1(n5648), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5911) );
  INV_X1 U7545 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8899) );
  OR2_X1 U7546 ( .A1(n6173), .A2(n8899), .ZN(n5910) );
  INV_X1 U7547 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5905) );
  NAND2_X1 U7548 ( .A1(n5906), .A2(n5905), .ZN(n5907) );
  NAND2_X1 U7549 ( .A1(n5922), .A2(n5907), .ZN(n8810) );
  OR2_X1 U7550 ( .A1(n6018), .A2(n8810), .ZN(n5909) );
  INV_X1 U7551 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8302) );
  OR2_X1 U7552 ( .A1(n5956), .A2(n8302), .ZN(n5908) );
  NAND4_X1 U7553 ( .A1(n5911), .A2(n5910), .A3(n5909), .A4(n5908), .ZN(n8846)
         );
  NAND2_X1 U7554 ( .A1(n8846), .A2(n7336), .ZN(n5912) );
  XNOR2_X1 U7555 ( .A(n5914), .B(n5912), .ZN(n8806) );
  NAND2_X1 U7556 ( .A1(n8805), .A2(n8806), .ZN(n5916) );
  INV_X1 U7557 ( .A(n5912), .ZN(n5913) );
  NAND2_X1 U7558 ( .A1(n5914), .A2(n5913), .ZN(n5915) );
  NAND2_X1 U7559 ( .A1(n7661), .A2(n6188), .ZN(n5920) );
  OAI22_X1 U7560 ( .A1(n5917), .A2(n7662), .B1(n10027), .B2(n5805), .ZN(n5918)
         );
  INV_X1 U7561 ( .A(n5918), .ZN(n5919) );
  XNOR2_X1 U7562 ( .A(n9155), .B(n6057), .ZN(n5928) );
  NAND2_X1 U7563 ( .A1(n5648), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5927) );
  INV_X1 U7564 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n5921) );
  OR2_X1 U7565 ( .A1(n6173), .A2(n5921), .ZN(n5926) );
  INV_X1 U7566 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n9078) );
  OR2_X1 U7567 ( .A1(n5956), .A2(n9078), .ZN(n5925) );
  INV_X1 U7568 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6488) );
  NAND2_X1 U7569 ( .A1(n5922), .A2(n6488), .ZN(n5923) );
  NAND2_X1 U7570 ( .A1(n5936), .A2(n5923), .ZN(n9077) );
  OR2_X1 U7571 ( .A1(n6018), .A2(n9077), .ZN(n5924) );
  NAND4_X1 U7572 ( .A1(n5927), .A2(n5926), .A3(n5925), .A4(n5924), .ZN(n9071)
         );
  NAND2_X1 U7573 ( .A1(n9071), .A2(n6196), .ZN(n5929) );
  NAND2_X1 U7574 ( .A1(n5928), .A2(n5929), .ZN(n8728) );
  INV_X1 U7575 ( .A(n5928), .ZN(n5931) );
  INV_X1 U7576 ( .A(n5929), .ZN(n5930) );
  NAND2_X1 U7577 ( .A1(n5931), .A2(n5930), .ZN(n8729) );
  NAND2_X1 U7578 ( .A1(n7743), .A2(n6188), .ZN(n5933) );
  NAND2_X1 U7579 ( .A1(n6189), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5932) );
  XNOR2_X1 U7580 ( .A(n9149), .B(n6032), .ZN(n5943) );
  NAND2_X1 U7581 ( .A1(n5980), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5942) );
  INV_X1 U7582 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n5935) );
  NAND2_X1 U7583 ( .A1(n5936), .A2(n5935), .ZN(n5937) );
  NAND2_X1 U7584 ( .A1(n5952), .A2(n5937), .ZN(n8786) );
  OR2_X1 U7585 ( .A1(n8786), .A2(n6018), .ZN(n5941) );
  INV_X1 U7586 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n6490) );
  OR2_X1 U7587 ( .A1(n6175), .A2(n6490), .ZN(n5940) );
  INV_X1 U7588 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n5938) );
  OR2_X1 U7589 ( .A1(n5956), .A2(n5938), .ZN(n5939) );
  NAND4_X1 U7590 ( .A1(n5942), .A2(n5941), .A3(n5940), .A4(n5939), .ZN(n8845)
         );
  AND2_X1 U7591 ( .A1(n8845), .A2(n7336), .ZN(n5944) );
  NAND2_X1 U7592 ( .A1(n5943), .A2(n5944), .ZN(n8740) );
  INV_X1 U7593 ( .A(n5943), .ZN(n5946) );
  INV_X1 U7594 ( .A(n5944), .ZN(n5945) );
  NAND2_X1 U7595 ( .A1(n5946), .A2(n5945), .ZN(n5947) );
  NAND2_X1 U7596 ( .A1(n7818), .A2(n6188), .ZN(n5949) );
  NAND2_X1 U7597 ( .A1(n6189), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5948) );
  XNOR2_X1 U7598 ( .A(n9146), .B(n6032), .ZN(n5966) );
  INV_X1 U7599 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n9040) );
  NAND2_X1 U7600 ( .A1(n5648), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5951) );
  NAND2_X1 U7601 ( .A1(n5980), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5950) );
  AND2_X1 U7602 ( .A1(n5951), .A2(n5950), .ZN(n5955) );
  INV_X1 U7603 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8745) );
  NAND2_X1 U7604 ( .A1(n5952), .A2(n8745), .ZN(n5953) );
  NAND2_X1 U7605 ( .A1(n5960), .A2(n5953), .ZN(n9039) );
  OR2_X1 U7606 ( .A1(n9039), .A2(n6018), .ZN(n5954) );
  OAI211_X1 U7607 ( .C1(n5956), .C2(n9040), .A(n5955), .B(n5954), .ZN(n9069)
         );
  NAND2_X1 U7608 ( .A1(n9069), .A2(n7336), .ZN(n5964) );
  XNOR2_X1 U7609 ( .A(n5966), .B(n5964), .ZN(n8744) );
  AND2_X1 U7610 ( .A1(n8785), .A2(n8744), .ZN(n5957) );
  NAND2_X1 U7611 ( .A1(n7845), .A2(n6188), .ZN(n5959) );
  NAND2_X1 U7612 ( .A1(n6189), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5958) );
  XNOR2_X1 U7613 ( .A(n9141), .B(n6032), .ZN(n8796) );
  INV_X1 U7614 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8799) );
  NAND2_X1 U7615 ( .A1(n5960), .A2(n8799), .ZN(n5961) );
  NAND2_X1 U7616 ( .A1(n5978), .A2(n5961), .ZN(n9029) );
  AOI22_X1 U7617 ( .A1(n5980), .A2(P2_REG1_REG_22__SCAN_IN), .B1(n5648), .B2(
        P2_REG0_REG_22__SCAN_IN), .ZN(n5963) );
  NAND2_X1 U7618 ( .A1(n6166), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5962) );
  OAI211_X1 U7619 ( .C1(n9029), .C2(n6018), .A(n5963), .B(n5962), .ZN(n8844)
         );
  AND2_X1 U7620 ( .A1(n8844), .A2(n7336), .ZN(n8795) );
  INV_X1 U7621 ( .A(n5964), .ZN(n5965) );
  AND2_X1 U7622 ( .A1(n5966), .A2(n5965), .ZN(n8793) );
  AOI21_X1 U7623 ( .B1(n8796), .B2(n8795), .A(n8793), .ZN(n5968) );
  INV_X1 U7624 ( .A(n8744), .ZN(n5967) );
  OR2_X1 U7625 ( .A1(n5967), .A2(n8740), .ZN(n8741) );
  AND2_X1 U7626 ( .A1(n5968), .A2(n8741), .ZN(n5969) );
  NAND2_X1 U7627 ( .A1(n8742), .A2(n5969), .ZN(n5973) );
  INV_X1 U7628 ( .A(n8796), .ZN(n5971) );
  INV_X1 U7629 ( .A(n8795), .ZN(n5970) );
  NAND2_X1 U7630 ( .A1(n5971), .A2(n5970), .ZN(n5972) );
  NAND2_X1 U7631 ( .A1(n5973), .A2(n5972), .ZN(n8722) );
  NAND2_X1 U7632 ( .A1(n7951), .A2(n6188), .ZN(n5975) );
  NAND2_X1 U7633 ( .A1(n6189), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5974) );
  XNOR2_X1 U7634 ( .A(n9135), .B(n6057), .ZN(n8720) );
  INV_X1 U7635 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n6418) );
  INV_X1 U7636 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n5977) );
  NAND2_X1 U7637 ( .A1(n5978), .A2(n5977), .ZN(n5979) );
  NAND2_X1 U7638 ( .A1(n5988), .A2(n5979), .ZN(n9009) );
  OR2_X1 U7639 ( .A1(n9009), .A2(n6018), .ZN(n5982) );
  AOI22_X1 U7640 ( .A1(n5980), .A2(P2_REG1_REG_23__SCAN_IN), .B1(n6166), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n5981) );
  OAI211_X1 U7641 ( .C1(n6175), .C2(n6418), .A(n5982), .B(n5981), .ZN(n8997)
         );
  NAND2_X1 U7642 ( .A1(n8997), .A2(n7336), .ZN(n8719) );
  NAND2_X1 U7643 ( .A1(n8722), .A2(n8720), .ZN(n5983) );
  NAND2_X1 U7644 ( .A1(n5984), .A2(n5983), .ZN(n8773) );
  NAND2_X1 U7645 ( .A1(n8004), .A2(n6188), .ZN(n5986) );
  NAND2_X1 U7646 ( .A1(n6189), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5985) );
  XNOR2_X1 U7647 ( .A(n9127), .B(n6057), .ZN(n8775) );
  INV_X1 U7648 ( .A(n5988), .ZN(n5987) );
  NAND2_X1 U7649 ( .A1(n5987), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5999) );
  INV_X1 U7650 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8777) );
  NAND2_X1 U7651 ( .A1(n5988), .A2(n8777), .ZN(n5989) );
  NAND2_X1 U7652 ( .A1(n5999), .A2(n5989), .ZN(n8984) );
  OR2_X1 U7653 ( .A1(n8984), .A2(n6018), .ZN(n5995) );
  INV_X1 U7654 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n5992) );
  NAND2_X1 U7655 ( .A1(n5648), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5991) );
  NAND2_X1 U7656 ( .A1(n6166), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5990) );
  OAI211_X1 U7657 ( .C1(n6173), .C2(n5992), .A(n5991), .B(n5990), .ZN(n5993)
         );
  INV_X1 U7658 ( .A(n5993), .ZN(n5994) );
  NAND2_X1 U7659 ( .A1(n5995), .A2(n5994), .ZN(n8843) );
  NAND2_X1 U7660 ( .A1(n8843), .A2(n7336), .ZN(n8774) );
  NAND2_X1 U7661 ( .A1(n8214), .A2(n6188), .ZN(n5997) );
  NAND2_X1 U7662 ( .A1(n6189), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5996) );
  XNOR2_X1 U7663 ( .A(n9124), .B(n6032), .ZN(n6007) );
  INV_X1 U7664 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5998) );
  NAND2_X1 U7665 ( .A1(n5999), .A2(n5998), .ZN(n6000) );
  AND2_X1 U7666 ( .A1(n6016), .A2(n6000), .ZN(n8972) );
  NAND2_X1 U7667 ( .A1(n8972), .A2(n6099), .ZN(n6006) );
  INV_X1 U7668 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n6003) );
  NAND2_X1 U7669 ( .A1(n5648), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6002) );
  NAND2_X1 U7670 ( .A1(n6166), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6001) );
  OAI211_X1 U7671 ( .C1(n6173), .C2(n6003), .A(n6002), .B(n6001), .ZN(n6004)
         );
  INV_X1 U7672 ( .A(n6004), .ZN(n6005) );
  NAND2_X1 U7673 ( .A1(n6006), .A2(n6005), .ZN(n8988) );
  AND2_X1 U7674 ( .A1(n8988), .A2(n7336), .ZN(n6008) );
  NAND2_X1 U7675 ( .A1(n6007), .A2(n6008), .ZN(n6012) );
  INV_X1 U7676 ( .A(n6007), .ZN(n6010) );
  INV_X1 U7677 ( .A(n6008), .ZN(n6009) );
  NAND2_X1 U7678 ( .A1(n6010), .A2(n6009), .ZN(n6011) );
  NAND2_X1 U7679 ( .A1(n6012), .A2(n6011), .ZN(n8750) );
  NAND2_X1 U7680 ( .A1(n8220), .A2(n6188), .ZN(n6014) );
  NAND2_X1 U7681 ( .A1(n6189), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6013) );
  XNOR2_X1 U7682 ( .A(n9119), .B(n6032), .ZN(n6025) );
  INV_X1 U7683 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8817) );
  NAND2_X1 U7684 ( .A1(n6016), .A2(n8817), .ZN(n6017) );
  NAND2_X1 U7685 ( .A1(n6049), .A2(n6017), .ZN(n8958) );
  OR2_X1 U7686 ( .A1(n8958), .A2(n6018), .ZN(n6024) );
  INV_X1 U7687 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n6021) );
  NAND2_X1 U7688 ( .A1(n5648), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6020) );
  NAND2_X1 U7689 ( .A1(n6166), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6019) );
  OAI211_X1 U7690 ( .C1(n6173), .C2(n6021), .A(n6020), .B(n6019), .ZN(n6022)
         );
  INV_X1 U7691 ( .A(n6022), .ZN(n6023) );
  NAND2_X1 U7692 ( .A1(n6024), .A2(n6023), .ZN(n8842) );
  AND2_X1 U7693 ( .A1(n8842), .A2(n7336), .ZN(n6026) );
  NAND2_X1 U7694 ( .A1(n6025), .A2(n6026), .ZN(n8709) );
  INV_X1 U7695 ( .A(n6025), .ZN(n6028) );
  INV_X1 U7696 ( .A(n6026), .ZN(n6027) );
  NAND2_X1 U7697 ( .A1(n6028), .A2(n6027), .ZN(n6029) );
  NAND2_X1 U7698 ( .A1(n8320), .A2(n6188), .ZN(n6031) );
  NAND2_X1 U7699 ( .A1(n6189), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6030) );
  XNOR2_X1 U7700 ( .A(n9113), .B(n6032), .ZN(n6039) );
  NAND2_X1 U7701 ( .A1(n8941), .A2(n6099), .ZN(n6038) );
  INV_X1 U7702 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n6035) );
  NAND2_X1 U7703 ( .A1(n6166), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6034) );
  NAND2_X1 U7704 ( .A1(n5648), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6033) );
  OAI211_X1 U7705 ( .C1(n6173), .C2(n6035), .A(n6034), .B(n6033), .ZN(n6036)
         );
  INV_X1 U7706 ( .A(n6036), .ZN(n6037) );
  NAND2_X1 U7707 ( .A1(n6038), .A2(n6037), .ZN(n8841) );
  AND2_X1 U7708 ( .A1(n8841), .A2(n6196), .ZN(n6040) );
  NAND2_X1 U7709 ( .A1(n6039), .A2(n6040), .ZN(n6046) );
  INV_X1 U7710 ( .A(n6039), .ZN(n6042) );
  INV_X1 U7711 ( .A(n6040), .ZN(n6041) );
  NAND2_X1 U7712 ( .A1(n6042), .A2(n6041), .ZN(n6043) );
  AND2_X1 U7713 ( .A1(n8815), .A2(n8711), .ZN(n6045) );
  INV_X1 U7714 ( .A(n8711), .ZN(n6044) );
  NAND2_X1 U7715 ( .A1(n8710), .A2(n6046), .ZN(n6060) );
  INV_X1 U7716 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8714) );
  INV_X1 U7717 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6047) );
  OAI21_X1 U7718 ( .B1(n6049), .B2(n8714), .A(n6047), .ZN(n6050) );
  NAND2_X1 U7719 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n6048) );
  NAND2_X1 U7720 ( .A1(n8932), .A2(n6099), .ZN(n6056) );
  INV_X1 U7721 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6053) );
  NAND2_X1 U7722 ( .A1(n5648), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6052) );
  NAND2_X1 U7723 ( .A1(n6166), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6051) );
  OAI211_X1 U7724 ( .C1(n6173), .C2(n6053), .A(n6052), .B(n6051), .ZN(n6054)
         );
  INV_X1 U7725 ( .A(n6054), .ZN(n6055) );
  NAND2_X1 U7726 ( .A1(n6056), .A2(n6055), .ZN(n8840) );
  XNOR2_X1 U7727 ( .A(n8840), .B(n6057), .ZN(n6058) );
  NAND2_X1 U7728 ( .A1(n6058), .A2(n7336), .ZN(n6059) );
  XNOR2_X1 U7729 ( .A(n6060), .B(n6059), .ZN(n6095) );
  INV_X1 U7730 ( .A(n6095), .ZN(n6092) );
  NAND2_X1 U7731 ( .A1(n6061), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6062) );
  MUX2_X1 U7732 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6062), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6063) );
  INV_X1 U7733 ( .A(n8222), .ZN(n6073) );
  NOR2_X1 U7734 ( .A1(n6064), .A2(n5554), .ZN(n6065) );
  MUX2_X1 U7735 ( .A(n5554), .B(n6065), .S(P2_IR_REG_25__SCAN_IN), .Z(n6066)
         );
  INV_X1 U7736 ( .A(n6066), .ZN(n6067) );
  NAND2_X1 U7737 ( .A1(n6067), .A2(n6061), .ZN(n8215) );
  NAND2_X1 U7738 ( .A1(n6087), .A2(n6086), .ZN(n6089) );
  NAND2_X1 U7739 ( .A1(n6089), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6070) );
  INV_X1 U7740 ( .A(P2_B_REG_SCAN_IN), .ZN(n8686) );
  XOR2_X1 U7741 ( .A(n8006), .B(n8686), .Z(n6071) );
  NAND2_X1 U7742 ( .A1(n8215), .A2(n6071), .ZN(n6072) );
  INV_X1 U7743 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10043) );
  AND2_X1 U7744 ( .A1(n8222), .A2(n8215), .ZN(n10044) );
  NOR4_X1 U7745 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n6077) );
  NOR4_X1 U7746 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n6076) );
  NOR4_X1 U7747 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n6075) );
  NOR4_X1 U7748 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n6074) );
  NAND4_X1 U7749 ( .A1(n6077), .A2(n6076), .A3(n6075), .A4(n6074), .ZN(n6083)
         );
  NOR2_X1 U7750 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .ZN(
        n6081) );
  NOR4_X1 U7751 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n6080) );
  NOR4_X1 U7752 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n6079) );
  NOR4_X1 U7753 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_30__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6078) );
  NAND4_X1 U7754 ( .A1(n6081), .A2(n6080), .A3(n6079), .A4(n6078), .ZN(n6082)
         );
  OAI21_X1 U7755 ( .B1(n6083), .B2(n6082), .A(n10034), .ZN(n7324) );
  INV_X1 U7756 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10040) );
  AND2_X1 U7757 ( .A1(n7324), .A2(n7544), .ZN(n6085) );
  NAND2_X1 U7758 ( .A1(n7541), .A2(n6085), .ZN(n6096) );
  INV_X1 U7759 ( .A(n6096), .ZN(n6107) );
  OR2_X1 U7760 ( .A1(n6087), .A2(n6086), .ZN(n6088) );
  NAND2_X1 U7761 ( .A1(n6089), .A2(n6088), .ZN(n6376) );
  INV_X1 U7762 ( .A(n7847), .ZN(n7327) );
  NAND2_X1 U7763 ( .A1(n7327), .A2(n6226), .ZN(n7326) );
  NAND2_X1 U7764 ( .A1(n10095), .A2(n7326), .ZN(n6090) );
  NOR2_X1 U7765 ( .A1(n10035), .A2(n6090), .ZN(n6091) );
  NAND2_X1 U7766 ( .A1(n6092), .A2(n10002), .ZN(n6113) );
  NAND2_X1 U7767 ( .A1(n8309), .A2(n6188), .ZN(n6094) );
  NAND2_X1 U7768 ( .A1(n6189), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6093) );
  NAND3_X1 U7769 ( .A1(n7847), .A2(n8974), .A3(n7745), .ZN(n10087) );
  NAND2_X1 U7770 ( .A1(n6096), .A2(n7538), .ZN(n6110) );
  NOR2_X1 U7771 ( .A1(n10035), .A2(n10095), .ZN(n6097) );
  NOR2_X2 U7772 ( .A1(n8663), .A2(n7326), .ZN(n9070) );
  INV_X1 U7773 ( .A(n6098), .ZN(n8680) );
  NAND2_X1 U7774 ( .A1(n8680), .A2(n6099), .ZN(n6105) );
  INV_X1 U7775 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6102) );
  NAND2_X1 U7776 ( .A1(n6166), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6101) );
  NAND2_X1 U7777 ( .A1(n5648), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6100) );
  OAI211_X1 U7778 ( .C1(n6173), .C2(n6102), .A(n6101), .B(n6100), .ZN(n6103)
         );
  INV_X1 U7779 ( .A(n6103), .ZN(n6104) );
  NAND2_X1 U7780 ( .A1(n6105), .A2(n6104), .ZN(n8839) );
  INV_X1 U7781 ( .A(n7326), .ZN(n7041) );
  AOI22_X1 U7782 ( .A1(n8841), .A2(n9070), .B1(n8839), .B2(n9068), .ZN(n8929)
         );
  INV_X1 U7783 ( .A(n6108), .ZN(n6106) );
  NOR2_X1 U7784 ( .A1(n10035), .A2(n6106), .ZN(n6378) );
  NAND2_X1 U7785 ( .A1(n6107), .A2(n6378), .ZN(n8800) );
  OR2_X1 U7786 ( .A1(n7326), .A2(n6108), .ZN(n7321) );
  AND3_X1 U7787 ( .A1(n7038), .A2(n6376), .A3(n7321), .ZN(n6109) );
  NAND2_X1 U7788 ( .A1(n6110), .A2(n6109), .ZN(n7102) );
  INV_X1 U7789 ( .A(n10006), .ZN(n8789) );
  AOI22_X1 U7790 ( .A1(n8932), .A2(n8789), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n6111) );
  OAI21_X1 U7791 ( .B1(n8929), .B2(n8800), .A(n6111), .ZN(n6112) );
  INV_X1 U7792 ( .A(n8861), .ZN(n8696) );
  NAND2_X1 U7793 ( .A1(n8696), .A2(n7546), .ZN(n6204) );
  INV_X1 U7794 ( .A(n7467), .ZN(n10047) );
  NAND2_X1 U7795 ( .A1(n6204), .A2(n7461), .ZN(n6114) );
  NAND2_X1 U7796 ( .A1(n8861), .A2(n10052), .ZN(n7460) );
  NAND2_X1 U7797 ( .A1(n6114), .A2(n7460), .ZN(n6224) );
  INV_X1 U7798 ( .A(n6224), .ZN(n6118) );
  NAND2_X1 U7799 ( .A1(n6115), .A2(n10058), .ZN(n6236) );
  INV_X1 U7800 ( .A(n8700), .ZN(n6117) );
  NAND2_X1 U7801 ( .A1(n6118), .A2(n6117), .ZN(n7666) );
  NAND2_X1 U7802 ( .A1(n8860), .A2(n10062), .ZN(n6246) );
  AND2_X1 U7803 ( .A1(n7748), .A2(n6246), .ZN(n6231) );
  NAND2_X1 U7804 ( .A1(n7555), .A2(n7756), .ZN(n7564) );
  NAND2_X1 U7805 ( .A1(n7634), .A2(n10022), .ZN(n6232) );
  NAND2_X1 U7806 ( .A1(n7564), .A2(n6232), .ZN(n6228) );
  INV_X1 U7807 ( .A(n6228), .ZN(n6120) );
  NAND2_X1 U7808 ( .A1(n7563), .A2(n6120), .ZN(n6121) );
  NAND2_X1 U7809 ( .A1(n6121), .A2(n6249), .ZN(n7632) );
  INV_X1 U7810 ( .A(n7632), .ZN(n6123) );
  NOR2_X1 U7811 ( .A1(n8857), .A2(n10076), .ZN(n6254) );
  INV_X1 U7812 ( .A(n6254), .ZN(n6124) );
  NAND2_X1 U7813 ( .A1(n8857), .A2(n10076), .ZN(n6250) );
  NAND2_X1 U7814 ( .A1(n6124), .A2(n6250), .ZN(n7631) );
  INV_X1 U7815 ( .A(n9997), .ZN(n7720) );
  NAND2_X1 U7816 ( .A1(n7720), .A2(n7822), .ZN(n6259) );
  INV_X1 U7817 ( .A(n7822), .ZN(n7801) );
  NAND2_X1 U7818 ( .A1(n9997), .A2(n7801), .ZN(n6260) );
  NAND2_X1 U7819 ( .A1(n6259), .A2(n6260), .ZN(n7855) );
  INV_X1 U7820 ( .A(n6260), .ZN(n6125) );
  NAND2_X1 U7821 ( .A1(n7517), .A2(n7851), .ZN(n6263) );
  INV_X1 U7822 ( .A(n7851), .ZN(n10084) );
  NAND2_X1 U7823 ( .A1(n10084), .A2(n8856), .ZN(n6262) );
  NAND2_X1 U7824 ( .A1(n7715), .A2(n6126), .ZN(n7714) );
  NAND2_X1 U7825 ( .A1(n7714), .A2(n6263), .ZN(n7850) );
  NAND2_X1 U7826 ( .A1(n7957), .A2(n9994), .ZN(n6264) );
  INV_X1 U7827 ( .A(n6264), .ZN(n6273) );
  NOR2_X1 U7828 ( .A1(n7957), .A2(n9994), .ZN(n6268) );
  INV_X1 U7829 ( .A(n6268), .ZN(n6275) );
  OAI21_X1 U7830 ( .B1(n7850), .B2(n6273), .A(n6275), .ZN(n7882) );
  INV_X1 U7831 ( .A(n8854), .ZN(n6129) );
  AND2_X1 U7832 ( .A1(n7986), .A2(n6129), .ZN(n6274) );
  INV_X1 U7833 ( .A(n6274), .ZN(n8008) );
  INV_X1 U7834 ( .A(n8852), .ZN(n7985) );
  NAND2_X1 U7835 ( .A1(n8083), .A2(n7985), .ZN(n6281) );
  AND2_X1 U7836 ( .A1(n8071), .A2(n6281), .ZN(n6128) );
  AND2_X1 U7837 ( .A1(n8008), .A2(n6128), .ZN(n6127) );
  NAND2_X1 U7838 ( .A1(n7882), .A2(n6127), .ZN(n7981) );
  INV_X1 U7839 ( .A(n6128), .ZN(n6130) );
  OR2_X1 U7840 ( .A1(n8040), .A2(n8075), .ZN(n6278) );
  NOR2_X1 U7841 ( .A1(n7986), .A2(n6129), .ZN(n6269) );
  INV_X1 U7842 ( .A(n6269), .ZN(n8010) );
  NAND2_X1 U7843 ( .A1(n6278), .A2(n8010), .ZN(n6276) );
  INV_X1 U7844 ( .A(n6276), .ZN(n8069) );
  OR2_X1 U7845 ( .A1(n6130), .A2(n8069), .ZN(n7980) );
  INV_X1 U7846 ( .A(n8851), .ZN(n8077) );
  NOR2_X1 U7847 ( .A1(n9179), .A2(n8077), .ZN(n6285) );
  INV_X1 U7848 ( .A(n6285), .ZN(n6131) );
  AND2_X1 U7849 ( .A1(n9179), .A2(n8077), .ZN(n6286) );
  INV_X1 U7850 ( .A(n6286), .ZN(n6134) );
  OR2_X1 U7851 ( .A1(n8083), .A2(n7985), .ZN(n7982) );
  AND2_X1 U7852 ( .A1(n7991), .A2(n7982), .ZN(n6132) );
  AND2_X1 U7853 ( .A1(n7980), .A2(n6132), .ZN(n6133) );
  INV_X1 U7854 ( .A(n8850), .ZN(n8155) );
  NAND2_X1 U7855 ( .A1(n8264), .A2(n8155), .ZN(n6290) );
  NAND2_X1 U7856 ( .A1(n6289), .A2(n6290), .ZN(n8156) );
  INV_X1 U7857 ( .A(n8849), .ZN(n8228) );
  AND2_X1 U7858 ( .A1(n8833), .A2(n8228), .ZN(n6293) );
  OR2_X1 U7859 ( .A1(n9172), .A2(n8828), .ZN(n6297) );
  NAND2_X1 U7860 ( .A1(n9172), .A2(n8828), .ZN(n8284) );
  NAND2_X1 U7861 ( .A1(n6297), .A2(n8284), .ZN(n8288) );
  NOR2_X1 U7862 ( .A1(n9167), .A2(n8766), .ZN(n6300) );
  INV_X1 U7863 ( .A(n6300), .ZN(n6304) );
  NAND2_X1 U7864 ( .A1(n9167), .A2(n8766), .ZN(n6302) );
  NAND2_X1 U7865 ( .A1(n6304), .A2(n6302), .ZN(n8290) );
  INV_X1 U7866 ( .A(n8284), .ZN(n6136) );
  NOR2_X1 U7867 ( .A1(n8290), .A2(n6136), .ZN(n6137) );
  NAND2_X1 U7868 ( .A1(n8285), .A2(n6137), .ZN(n6138) );
  NAND2_X1 U7869 ( .A1(n6138), .A2(n6304), .ZN(n8305) );
  INV_X1 U7870 ( .A(n8305), .ZN(n6139) );
  OR2_X1 U7871 ( .A1(n9161), .A2(n8667), .ZN(n6312) );
  NAND2_X1 U7872 ( .A1(n9161), .A2(n8667), .ZN(n6315) );
  NOR2_X1 U7873 ( .A1(n9155), .A2(n8807), .ZN(n6317) );
  INV_X1 U7874 ( .A(n6317), .ZN(n6141) );
  INV_X1 U7875 ( .A(n8845), .ZN(n9050) );
  NAND2_X1 U7876 ( .A1(n9149), .A2(n9050), .ZN(n6328) );
  NAND2_X1 U7877 ( .A1(n6318), .A2(n6328), .ZN(n9056) );
  NOR2_X1 U7878 ( .A1(n9056), .A2(n6314), .ZN(n6142) );
  INV_X1 U7879 ( .A(n9046), .ZN(n6144) );
  INV_X1 U7880 ( .A(n9069), .ZN(n8673) );
  XNOR2_X1 U7881 ( .A(n9146), .B(n8673), .ZN(n9047) );
  INV_X1 U7882 ( .A(n9047), .ZN(n6143) );
  NAND2_X1 U7883 ( .A1(n6144), .A2(n6143), .ZN(n9044) );
  INV_X1 U7884 ( .A(n8844), .ZN(n9052) );
  NOR2_X1 U7885 ( .A1(n9141), .A2(n9052), .ZN(n6320) );
  INV_X1 U7886 ( .A(n6320), .ZN(n6331) );
  NAND2_X1 U7887 ( .A1(n9141), .A2(n9052), .ZN(n6333) );
  NAND2_X1 U7888 ( .A1(n6331), .A2(n6333), .ZN(n9018) );
  NAND2_X1 U7889 ( .A1(n9146), .A2(n8673), .ZN(n9022) );
  INV_X1 U7890 ( .A(n9022), .ZN(n6145) );
  NOR2_X1 U7891 ( .A1(n9018), .A2(n6145), .ZN(n6146) );
  INV_X1 U7892 ( .A(n8997), .ZN(n8778) );
  NOR2_X1 U7893 ( .A1(n9135), .A2(n8778), .ZN(n6321) );
  INV_X1 U7894 ( .A(n6321), .ZN(n6147) );
  NAND2_X1 U7895 ( .A1(n6147), .A2(n8991), .ZN(n8674) );
  NAND2_X1 U7896 ( .A1(n9127), .A2(n9003), .ZN(n6322) );
  NAND2_X1 U7897 ( .A1(n8964), .A2(n6322), .ZN(n8980) );
  NOR2_X1 U7898 ( .A1(n8980), .A2(n6323), .ZN(n6148) );
  OR2_X1 U7899 ( .A1(n9124), .A2(n8954), .ZN(n6337) );
  NAND2_X1 U7900 ( .A1(n6337), .A2(n8964), .ZN(n6223) );
  INV_X1 U7901 ( .A(n6223), .ZN(n6327) );
  NAND2_X1 U7902 ( .A1(n8989), .A2(n6327), .ZN(n6149) );
  NAND2_X1 U7903 ( .A1(n9124), .A2(n8954), .ZN(n6325) );
  NAND2_X1 U7904 ( .A1(n6149), .A2(n6325), .ZN(n8952) );
  NOR2_X1 U7905 ( .A1(n9119), .A2(n8968), .ZN(n6341) );
  INV_X1 U7906 ( .A(n6341), .ZN(n6203) );
  NAND2_X1 U7907 ( .A1(n9119), .A2(n8968), .ZN(n6343) );
  NAND2_X1 U7908 ( .A1(n9113), .A2(n8956), .ZN(n6351) );
  INV_X1 U7909 ( .A(n8840), .ZN(n8713) );
  NOR2_X1 U7910 ( .A1(n9109), .A2(n8713), .ZN(n6358) );
  INV_X1 U7911 ( .A(n6358), .ZN(n6150) );
  NOR2_X1 U7912 ( .A1(n6342), .A2(n8924), .ZN(n6151) );
  NAND2_X1 U7913 ( .A1(n6153), .A2(n6152), .ZN(n8684) );
  INV_X1 U7914 ( .A(n8839), .ZN(n6154) );
  INV_X1 U7915 ( .A(n6179), .ZN(n6181) );
  INV_X1 U7916 ( .A(n6162), .ZN(n6160) );
  INV_X1 U7917 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9701) );
  INV_X1 U7918 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n6158) );
  MUX2_X1 U7919 ( .A(n9701), .B(n6158), .S(n6799), .Z(n6161) );
  INV_X1 U7920 ( .A(n6161), .ZN(n6159) );
  NAND2_X1 U7921 ( .A1(n9206), .A2(n6188), .ZN(n6165) );
  NAND2_X1 U7922 ( .A1(n6189), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n6164) );
  NAND2_X1 U7923 ( .A1(n6166), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6171) );
  INV_X1 U7924 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n6167) );
  OR2_X1 U7925 ( .A1(n6173), .A2(n6167), .ZN(n6170) );
  INV_X1 U7926 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n6168) );
  OR2_X1 U7927 ( .A1(n6175), .A2(n6168), .ZN(n6169) );
  AND3_X1 U7928 ( .A1(n6171), .A2(n6170), .A3(n6169), .ZN(n8685) );
  INV_X1 U7929 ( .A(n6363), .ZN(n6201) );
  NAND2_X1 U7930 ( .A1(n6166), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6178) );
  INV_X1 U7931 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n6172) );
  OR2_X1 U7932 ( .A1(n6173), .A2(n6172), .ZN(n6177) );
  INV_X1 U7933 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n6174) );
  OR2_X1 U7934 ( .A1(n6175), .A2(n6174), .ZN(n6176) );
  OAI22_X1 U7935 ( .A1(n6179), .A2(n6201), .B1(n7820), .B2(n8913), .ZN(n6180)
         );
  OAI21_X1 U7936 ( .B1(n6181), .B2(n9097), .A(n6180), .ZN(n6194) );
  INV_X1 U7937 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6185) );
  INV_X1 U7938 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6184) );
  MUX2_X1 U7939 ( .A(n6185), .B(n6184), .S(n6799), .Z(n6186) );
  XNOR2_X1 U7940 ( .A(n6186), .B(SI_31_), .ZN(n6187) );
  NAND2_X1 U7941 ( .A1(n6189), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n6190) );
  NAND2_X1 U7942 ( .A1(n9097), .A2(n8685), .ZN(n6366) );
  NAND2_X1 U7943 ( .A1(n6368), .A2(n6366), .ZN(n6362) );
  INV_X1 U7944 ( .A(n6362), .ZN(n6217) );
  XNOR2_X1 U7945 ( .A(n6195), .B(n10027), .ZN(n6199) );
  INV_X1 U7946 ( .A(n6196), .ZN(n7185) );
  INV_X1 U7947 ( .A(n7331), .ZN(n6197) );
  NAND2_X1 U7948 ( .A1(n6199), .A2(n6198), .ZN(n6375) );
  NOR2_X1 U7949 ( .A1(n6364), .A2(n6201), .ZN(n6370) );
  NAND2_X1 U7950 ( .A1(n6202), .A2(n6357), .ZN(n8683) );
  INV_X1 U7951 ( .A(n8980), .ZN(n8990) );
  AND2_X2 U7952 ( .A1(n6337), .A2(n6325), .ZN(n8965) );
  INV_X1 U7953 ( .A(n9056), .ZN(n9065) );
  NAND2_X1 U7954 ( .A1(n6305), .A2(n6303), .ZN(n8160) );
  NAND2_X1 U7955 ( .A1(n8863), .A2(n7467), .ZN(n7320) );
  NAND2_X1 U7956 ( .A1(n7460), .A2(n7320), .ZN(n6238) );
  NOR2_X1 U7957 ( .A1(n8700), .A2(n6238), .ZN(n6205) );
  INV_X1 U7958 ( .A(n6204), .ZN(n6235) );
  NAND4_X1 U7959 ( .A1(n6205), .A2(n6200), .A3(n7461), .A4(n6204), .ZN(n6207)
         );
  INV_X2 U7960 ( .A(n6231), .ZN(n7675) );
  NAND2_X1 U7961 ( .A1(n6232), .A2(n6249), .ZN(n7565) );
  NOR4_X1 U7962 ( .A1(n6207), .A2(n7675), .A3(n7747), .A4(n7565), .ZN(n6208)
         );
  NAND4_X1 U7963 ( .A1(n6208), .A2(n4619), .A3(n6126), .A4(n6122), .ZN(n6209)
         );
  NAND2_X1 U7964 ( .A1(n6278), .A2(n8071), .ZN(n8011) );
  NAND2_X1 U7965 ( .A1(n8010), .A2(n8008), .ZN(n7883) );
  NAND2_X1 U7966 ( .A1(n6275), .A2(n6264), .ZN(n7857) );
  NOR4_X1 U7967 ( .A1(n6209), .A2(n8011), .A3(n7883), .A4(n7857), .ZN(n6210)
         );
  NAND4_X1 U7968 ( .A1(n6135), .A2(n7991), .A3(n8074), .A4(n6210), .ZN(n6211)
         );
  NOR4_X1 U7969 ( .A1(n8290), .A2(n8288), .A3(n8160), .A4(n6211), .ZN(n6212)
         );
  NAND4_X1 U7970 ( .A1(n9065), .A2(n4327), .A3(n9082), .A4(n6212), .ZN(n6213)
         );
  NOR4_X1 U7971 ( .A1(n8674), .A2(n9018), .A3(n9047), .A4(n6213), .ZN(n6214)
         );
  NAND4_X1 U7972 ( .A1(n8953), .A2(n8990), .A3(n8965), .A4(n6214), .ZN(n6215)
         );
  NOR4_X1 U7973 ( .A1(n8683), .A2(n8924), .A3(n8944), .A4(n6215), .ZN(n6216)
         );
  NAND3_X1 U7974 ( .A1(n6370), .A2(n6217), .A3(n6216), .ZN(n6219) );
  OAI21_X1 U7975 ( .B1(n6200), .B2(n7847), .A(n6218), .ZN(n6222) );
  INV_X1 U7976 ( .A(n6218), .ZN(n6221) );
  INV_X1 U7977 ( .A(n6219), .ZN(n6220) );
  NOR2_X1 U7978 ( .A1(n6223), .A2(n6321), .ZN(n6324) );
  OAI21_X1 U7979 ( .B1(n6238), .B2(n7820), .A(n6224), .ZN(n6225) );
  NAND2_X1 U7980 ( .A1(n6225), .A2(n6236), .ZN(n6227) );
  AND2_X1 U7981 ( .A1(n6226), .A2(n8974), .ZN(n7330) );
  NAND2_X1 U7982 ( .A1(n7330), .A2(n7847), .ZN(n6372) );
  NAND3_X1 U7983 ( .A1(n6227), .A2(n6372), .A3(n7667), .ZN(n6230) );
  INV_X1 U7984 ( .A(n6252), .ZN(n6229) );
  AND3_X1 U7985 ( .A1(n6231), .A2(n6230), .A3(n6229), .ZN(n6240) );
  AOI21_X1 U7986 ( .B1(n7564), .B2(n7748), .A(n6252), .ZN(n6234) );
  INV_X1 U7987 ( .A(n6232), .ZN(n6233) );
  NOR2_X1 U7988 ( .A1(n4738), .A2(n6235), .ZN(n6239) );
  INV_X1 U7989 ( .A(n6236), .ZN(n6237) );
  AOI21_X1 U7990 ( .B1(n6239), .B2(n6238), .A(n6237), .ZN(n6242) );
  INV_X1 U7991 ( .A(n6240), .ZN(n6241) );
  OAI22_X1 U7992 ( .A1(n6243), .A2(n4453), .B1(n6242), .B2(n6241), .ZN(n6244)
         );
  INV_X1 U7993 ( .A(n6245), .ZN(n6248) );
  INV_X1 U7994 ( .A(n6246), .ZN(n6247) );
  NOR2_X1 U7995 ( .A1(n6248), .A2(n6247), .ZN(n6251) );
  OAI211_X1 U7996 ( .C1(n6252), .C2(n6251), .A(n6250), .B(n6249), .ZN(n6253)
         );
  NAND2_X1 U7997 ( .A1(n6253), .A2(n4453), .ZN(n6257) );
  MUX2_X1 U7998 ( .A(n6260), .B(n6259), .S(n6372), .Z(n6261) );
  NAND2_X1 U7999 ( .A1(n6261), .A2(n6126), .ZN(n6266) );
  MUX2_X1 U8000 ( .A(n6263), .B(n6262), .S(n6372), .Z(n6265) );
  OAI211_X1 U8001 ( .C1(n6267), .C2(n6266), .A(n6265), .B(n6264), .ZN(n6272)
         );
  NOR2_X1 U8002 ( .A1(n6269), .A2(n6268), .ZN(n6271) );
  AOI211_X1 U8003 ( .C1(n6272), .C2(n6271), .A(n6270), .B(n6274), .ZN(n6277)
         );
  NAND2_X1 U8004 ( .A1(n6281), .A2(n8071), .ZN(n6280) );
  NAND2_X1 U8005 ( .A1(n7982), .A2(n6278), .ZN(n6279) );
  MUX2_X1 U8006 ( .A(n6280), .B(n6279), .S(n4453), .Z(n6283) );
  MUX2_X1 U8007 ( .A(n6281), .B(n7982), .S(n6372), .Z(n6282) );
  OAI21_X1 U8008 ( .B1(n6284), .B2(n6283), .A(n6282), .ZN(n6288) );
  MUX2_X1 U8009 ( .A(n6286), .B(n6285), .S(n6372), .Z(n6287) );
  AOI211_X1 U8010 ( .C1(n6288), .C2(n7991), .A(n6287), .B(n8156), .ZN(n6296)
         );
  NAND2_X1 U8011 ( .A1(n6305), .A2(n6289), .ZN(n6292) );
  INV_X1 U8012 ( .A(n6290), .ZN(n6291) );
  MUX2_X1 U8013 ( .A(n6292), .B(n6291), .S(n6372), .Z(n6294) );
  INV_X1 U8014 ( .A(n6297), .ZN(n6299) );
  NAND2_X1 U8015 ( .A1(n6302), .A2(n8284), .ZN(n6298) );
  MUX2_X1 U8016 ( .A(n6299), .B(n6298), .S(n6372), .Z(n6301) );
  OR2_X1 U8017 ( .A1(n6301), .A2(n6300), .ZN(n6306) );
  INV_X1 U8018 ( .A(n6306), .ZN(n6310) );
  OAI211_X1 U8019 ( .C1(n6306), .C2(n6303), .A(n6315), .B(n6302), .ZN(n6308)
         );
  OAI211_X1 U8020 ( .C1(n6306), .C2(n6305), .A(n6304), .B(n6312), .ZN(n6307)
         );
  MUX2_X1 U8021 ( .A(n6308), .B(n6307), .S(n6372), .Z(n6309) );
  AOI21_X1 U8022 ( .B1(n6311), .B2(n6310), .A(n6309), .ZN(n6316) );
  INV_X1 U8023 ( .A(n6312), .ZN(n6313) );
  INV_X1 U8024 ( .A(n9146), .ZN(n9038) );
  NAND2_X1 U8025 ( .A1(n9038), .A2(n9069), .ZN(n6330) );
  NAND2_X1 U8026 ( .A1(n6325), .A2(n6322), .ZN(n6338) );
  INV_X1 U8027 ( .A(n6325), .ZN(n6326) );
  NOR3_X1 U8028 ( .A1(n6327), .A2(n4453), .A3(n6326), .ZN(n6336) );
  NAND3_X1 U8029 ( .A1(n6329), .A2(n6328), .A3(n9022), .ZN(n6332) );
  NAND3_X1 U8030 ( .A1(n6332), .A2(n6331), .A3(n6330), .ZN(n6334) );
  NAND4_X1 U8031 ( .A1(n6334), .A2(n4453), .A3(n8991), .A4(n6333), .ZN(n6335)
         );
  NAND3_X1 U8032 ( .A1(n6338), .A2(n4453), .A3(n6337), .ZN(n6339) );
  NAND2_X1 U8033 ( .A1(n6340), .A2(n6339), .ZN(n6344) );
  NOR2_X1 U8034 ( .A1(n6342), .A2(n6341), .ZN(n6353) );
  NAND2_X1 U8035 ( .A1(n6351), .A2(n6343), .ZN(n6345) );
  AOI21_X1 U8036 ( .B1(n6344), .B2(n6353), .A(n6345), .ZN(n6348) );
  INV_X1 U8037 ( .A(n6345), .ZN(n6346) );
  AOI21_X1 U8038 ( .B1(n4453), .B2(n8926), .A(n6346), .ZN(n6347) );
  NOR4_X1 U8039 ( .A1(n6348), .A2(n6359), .A3(n6358), .A4(n6347), .ZN(n6356)
         );
  NAND2_X1 U8040 ( .A1(n6351), .A2(n6372), .ZN(n6352) );
  OAI22_X1 U8041 ( .A1(n6354), .A2(n6359), .B1(n6353), .B2(n6352), .ZN(n6355)
         );
  OAI22_X1 U8042 ( .A1(n6356), .A2(n6355), .B1(n4453), .B2(n6354), .ZN(n6361)
         );
  OAI211_X1 U8043 ( .C1(n6359), .C2(n6358), .A(n6372), .B(n6357), .ZN(n6360)
         );
  NAND2_X1 U8044 ( .A1(n6361), .A2(n6360), .ZN(n6367) );
  NAND2_X1 U8045 ( .A1(n6367), .A2(n6366), .ZN(n6371) );
  INV_X1 U8046 ( .A(n6368), .ZN(n6369) );
  OR2_X1 U8047 ( .A1(n7847), .A2(n10027), .ZN(n7332) );
  NOR2_X1 U8048 ( .A1(n6376), .A2(P2_U3152), .ZN(n7952) );
  INV_X1 U8049 ( .A(n8687), .ZN(n6377) );
  NAND3_X1 U8050 ( .A1(n6378), .A2(n9070), .A3(n6377), .ZN(n6380) );
  AOI21_X1 U8051 ( .B1(n7952), .B2(n7847), .A(n8686), .ZN(n6379) );
  NAND2_X1 U8052 ( .A1(n6380), .A2(n6379), .ZN(n6381) );
  NOR2_X1 U8053 ( .A1(keyinput4), .A2(keyinput14), .ZN(n6385) );
  NAND3_X1 U8054 ( .A1(keyinput11), .A2(keyinput34), .A3(keyinput9), .ZN(n6383) );
  NAND3_X1 U8055 ( .A1(keyinput10), .A2(keyinput61), .A3(keyinput56), .ZN(
        n6382) );
  NOR4_X1 U8056 ( .A1(keyinput15), .A2(keyinput49), .A3(n6383), .A4(n6382), 
        .ZN(n6384) );
  NAND4_X1 U8057 ( .A1(keyinput25), .A2(keyinput40), .A3(n6385), .A4(n6384), 
        .ZN(n6386) );
  NOR4_X1 U8058 ( .A1(keyinput37), .A2(keyinput59), .A3(keyinput62), .A4(n6386), .ZN(n6409) );
  NAND2_X1 U8059 ( .A1(keyinput21), .A2(keyinput24), .ZN(n6387) );
  NOR3_X1 U8060 ( .A1(keyinput55), .A2(keyinput18), .A3(n6387), .ZN(n6393) );
  NOR3_X1 U8061 ( .A1(keyinput35), .A2(keyinput8), .A3(keyinput17), .ZN(n6392)
         );
  NAND3_X1 U8062 ( .A1(keyinput22), .A2(keyinput42), .A3(keyinput41), .ZN(
        n6390) );
  INV_X1 U8063 ( .A(keyinput23), .ZN(n6388) );
  NAND3_X1 U8064 ( .A1(keyinput30), .A2(keyinput36), .A3(n6388), .ZN(n6389) );
  NOR4_X1 U8065 ( .A1(keyinput29), .A2(keyinput20), .A3(n6390), .A4(n6389), 
        .ZN(n6391) );
  NAND4_X1 U8066 ( .A1(n6393), .A2(keyinput0), .A3(n6392), .A4(n6391), .ZN(
        n6407) );
  NOR3_X1 U8067 ( .A1(keyinput31), .A2(keyinput26), .A3(keyinput48), .ZN(n6399) );
  INV_X1 U8068 ( .A(keyinput6), .ZN(n6394) );
  NOR4_X1 U8069 ( .A1(keyinput44), .A2(keyinput47), .A3(keyinput5), .A4(n6394), 
        .ZN(n6398) );
  NAND3_X1 U8070 ( .A1(keyinput51), .A2(keyinput39), .A3(keyinput54), .ZN(
        n6396) );
  NAND3_X1 U8071 ( .A1(keyinput63), .A2(keyinput28), .A3(keyinput16), .ZN(
        n6395) );
  NOR4_X1 U8072 ( .A1(keyinput60), .A2(keyinput52), .A3(n6396), .A4(n6395), 
        .ZN(n6397) );
  NAND4_X1 U8073 ( .A1(keyinput58), .A2(n6399), .A3(n6398), .A4(n6397), .ZN(
        n6406) );
  NAND4_X1 U8074 ( .A1(keyinput12), .A2(keyinput27), .A3(keyinput38), .A4(
        keyinput43), .ZN(n6405) );
  NOR2_X1 U8075 ( .A1(keyinput32), .A2(keyinput46), .ZN(n6403) );
  NAND3_X1 U8076 ( .A1(keyinput50), .A2(keyinput19), .A3(keyinput33), .ZN(
        n6401) );
  NAND3_X1 U8077 ( .A1(keyinput7), .A2(keyinput53), .A3(keyinput2), .ZN(n6400)
         );
  NOR4_X1 U8078 ( .A1(keyinput3), .A2(keyinput13), .A3(n6401), .A4(n6400), 
        .ZN(n6402) );
  NAND4_X1 U8079 ( .A1(keyinput45), .A2(keyinput1), .A3(n6403), .A4(n6402), 
        .ZN(n6404) );
  NOR4_X1 U8080 ( .A1(n6407), .A2(n6406), .A3(n6405), .A4(n6404), .ZN(n6408)
         );
  AOI21_X1 U8081 ( .B1(n6409), .B2(n6408), .A(keyinput57), .ZN(n6410) );
  MUX2_X1 U8082 ( .A(n6410), .B(keyinput57), .S(P2_IR_REG_23__SCAN_IN), .Z(
        n6513) );
  INV_X1 U8083 ( .A(keyinput24), .ZN(n6412) );
  AOI22_X1 U8084 ( .A1(n7581), .A2(keyinput18), .B1(P1_ADDR_REG_7__SCAN_IN), 
        .B2(n6412), .ZN(n6411) );
  OAI221_X1 U8085 ( .B1(n7581), .B2(keyinput18), .C1(n6412), .C2(
        P1_ADDR_REG_7__SCAN_IN), .A(n6411), .ZN(n6422) );
  INV_X1 U8086 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n10036) );
  INV_X1 U8087 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n6414) );
  AOI22_X1 U8088 ( .A1(n10036), .A2(keyinput21), .B1(keyinput22), .B2(n6414), 
        .ZN(n6413) );
  OAI221_X1 U8089 ( .B1(n10036), .B2(keyinput21), .C1(n6414), .C2(keyinput22), 
        .A(n6413), .ZN(n6421) );
  INV_X1 U8090 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6855) );
  AOI22_X1 U8091 ( .A1(n6855), .A2(keyinput29), .B1(n9953), .B2(keyinput42), 
        .ZN(n6415) );
  OAI221_X1 U8092 ( .B1(n6855), .B2(keyinput29), .C1(n9953), .C2(keyinput42), 
        .A(n6415), .ZN(n6420) );
  INV_X1 U8093 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n6417) );
  AOI22_X1 U8094 ( .A1(n6418), .A2(keyinput41), .B1(n6417), .B2(keyinput35), 
        .ZN(n6416) );
  OAI221_X1 U8095 ( .B1(n6418), .B2(keyinput41), .C1(n6417), .C2(keyinput35), 
        .A(n6416), .ZN(n6419) );
  NOR4_X1 U8096 ( .A1(n6422), .A2(n6421), .A3(n6420), .A4(n6419), .ZN(n6512)
         );
  AOI22_X1 U8097 ( .A1(n6424), .A2(keyinput4), .B1(n9952), .B2(keyinput40), 
        .ZN(n6423) );
  OAI221_X1 U8098 ( .B1(n6424), .B2(keyinput4), .C1(n9952), .C2(keyinput40), 
        .A(n6423), .ZN(n6430) );
  INV_X1 U8099 ( .A(P1_RD_REG_SCAN_IN), .ZN(n9796) );
  INV_X1 U8100 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7612) );
  AOI22_X1 U8101 ( .A1(n9796), .A2(keyinput31), .B1(keyinput26), .B2(n7612), 
        .ZN(n6425) );
  OAI221_X1 U8102 ( .B1(n9796), .B2(keyinput31), .C1(n7612), .C2(keyinput26), 
        .A(n6425), .ZN(n6429) );
  XNOR2_X1 U8103 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput25), .ZN(n6427) );
  XNOR2_X1 U8104 ( .A(keyinput47), .B(P1_REG0_REG_10__SCAN_IN), .ZN(n6426) );
  NAND2_X1 U8105 ( .A1(n6427), .A2(n6426), .ZN(n6428) );
  NOR3_X1 U8106 ( .A1(n6430), .A2(n6429), .A3(n6428), .ZN(n6463) );
  INV_X1 U8107 ( .A(keyinput48), .ZN(n6432) );
  AOI22_X1 U8108 ( .A1(n7269), .A2(keyinput44), .B1(P1_REG0_REG_31__SCAN_IN), 
        .B2(n6432), .ZN(n6431) );
  OAI221_X1 U8109 ( .B1(n7269), .B2(keyinput44), .C1(n6432), .C2(
        P1_REG0_REG_31__SCAN_IN), .A(n6431), .ZN(n6436) );
  INV_X1 U8110 ( .A(keyinput14), .ZN(n6434) );
  AOI22_X1 U8111 ( .A1(n8245), .A2(keyinput55), .B1(P2_ADDR_REG_18__SCAN_IN), 
        .B2(n6434), .ZN(n6433) );
  OAI221_X1 U8112 ( .B1(n8245), .B2(keyinput55), .C1(n6434), .C2(
        P2_ADDR_REG_18__SCAN_IN), .A(n6433), .ZN(n6435) );
  NOR2_X1 U8113 ( .A1(n6436), .A2(n6435), .ZN(n6462) );
  INV_X1 U8114 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9988) );
  AOI22_X1 U8115 ( .A1(n9988), .A2(keyinput9), .B1(n7341), .B2(keyinput10), 
        .ZN(n6437) );
  OAI221_X1 U8116 ( .B1(n9988), .B2(keyinput9), .C1(n7341), .C2(keyinput10), 
        .A(n6437), .ZN(n6453) );
  XNOR2_X1 U8117 ( .A(P1_REG1_REG_2__SCAN_IN), .B(keyinput5), .ZN(n6439) );
  NAND2_X1 U8118 ( .A1(n8081), .A2(keyinput37), .ZN(n6438) );
  OAI211_X1 U8119 ( .C1(keyinput37), .C2(n8081), .A(n6439), .B(n6438), .ZN(
        n6440) );
  INV_X1 U8120 ( .A(n6440), .ZN(n6446) );
  INV_X1 U8121 ( .A(keyinput50), .ZN(n6442) );
  INV_X1 U8122 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n6441) );
  XNOR2_X1 U8123 ( .A(n6442), .B(n6441), .ZN(n6445) );
  XNOR2_X1 U8124 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput6), .ZN(n6444) );
  XNOR2_X1 U8125 ( .A(P2_IR_REG_9__SCAN_IN), .B(keyinput12), .ZN(n6443) );
  NAND4_X1 U8126 ( .A1(n6446), .A2(n6445), .A3(n6444), .A4(n6443), .ZN(n6452)
         );
  XNOR2_X1 U8127 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(keyinput46), .ZN(n6450) );
  XNOR2_X1 U8128 ( .A(P2_IR_REG_7__SCAN_IN), .B(keyinput34), .ZN(n6449) );
  XNOR2_X1 U8129 ( .A(P2_REG3_REG_7__SCAN_IN), .B(keyinput11), .ZN(n6448) );
  XNOR2_X1 U8130 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput56), .ZN(n6447) );
  NAND4_X1 U8131 ( .A1(n6450), .A2(n6449), .A3(n6448), .A4(n6447), .ZN(n6451)
         );
  NOR3_X1 U8132 ( .A1(n6453), .A2(n6452), .A3(n6451), .ZN(n6461) );
  INV_X1 U8133 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6455) );
  AOI22_X1 U8134 ( .A1(n7526), .A2(keyinput49), .B1(n6455), .B2(keyinput61), 
        .ZN(n6454) );
  OAI221_X1 U8135 ( .B1(n7526), .B2(keyinput49), .C1(n6455), .C2(keyinput61), 
        .A(n6454), .ZN(n6459) );
  INV_X1 U8136 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9959) );
  INV_X1 U8137 ( .A(keyinput59), .ZN(n6457) );
  AOI22_X1 U8138 ( .A1(n9959), .A2(keyinput15), .B1(P1_REG0_REG_30__SCAN_IN), 
        .B2(n6457), .ZN(n6456) );
  OAI221_X1 U8139 ( .B1(n9959), .B2(keyinput15), .C1(n6457), .C2(
        P1_REG0_REG_30__SCAN_IN), .A(n6456), .ZN(n6458) );
  NOR2_X1 U8140 ( .A1(n6459), .A2(n6458), .ZN(n6460) );
  AND4_X1 U8141 ( .A1(n6463), .A2(n6462), .A3(n6461), .A4(n6460), .ZN(n6471)
         );
  INV_X1 U8142 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n10037) );
  OAI22_X1 U8143 ( .A1(n10037), .A2(keyinput62), .B1(n5833), .B2(keyinput13), 
        .ZN(n6464) );
  AOI221_X1 U8144 ( .B1(n10037), .B2(keyinput62), .C1(keyinput13), .C2(n5833), 
        .A(n6464), .ZN(n6470) );
  INV_X1 U8145 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n6466) );
  INV_X1 U8146 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n8029) );
  OAI22_X1 U8147 ( .A1(n6466), .A2(keyinput53), .B1(n8029), .B2(keyinput2), 
        .ZN(n6465) );
  AOI221_X1 U8148 ( .B1(n6466), .B2(keyinput53), .C1(keyinput2), .C2(n8029), 
        .A(n6465), .ZN(n6469) );
  INV_X1 U8149 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n10038) );
  OAI22_X1 U8150 ( .A1(n10038), .A2(keyinput33), .B1(n7273), .B2(keyinput32), 
        .ZN(n6467) );
  AOI221_X1 U8151 ( .B1(n10038), .B2(keyinput33), .C1(keyinput32), .C2(n7273), 
        .A(n6467), .ZN(n6468) );
  AND4_X1 U8152 ( .A1(n6471), .A2(n6470), .A3(n6469), .A4(n6468), .ZN(n6511)
         );
  INV_X1 U8153 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n6473) );
  AOI22_X1 U8154 ( .A1(n6473), .A2(keyinput8), .B1(n9956), .B2(keyinput17), 
        .ZN(n6472) );
  OAI221_X1 U8155 ( .B1(n6473), .B2(keyinput8), .C1(n9956), .C2(keyinput17), 
        .A(n6472), .ZN(n6482) );
  AOI22_X1 U8156 ( .A1(n6475), .A2(keyinput0), .B1(keyinput20), .B2(n6870), 
        .ZN(n6474) );
  OAI221_X1 U8157 ( .B1(n6475), .B2(keyinput0), .C1(n6870), .C2(keyinput20), 
        .A(n6474), .ZN(n6481) );
  INV_X1 U8158 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9360) );
  AOI22_X1 U8159 ( .A1(n9360), .A2(keyinput30), .B1(n9955), .B2(keyinput23), 
        .ZN(n6476) );
  OAI221_X1 U8160 ( .B1(n9360), .B2(keyinput30), .C1(n9955), .C2(keyinput23), 
        .A(n6476), .ZN(n6480) );
  INV_X1 U8161 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7828) );
  AOI22_X1 U8162 ( .A1(n6478), .A2(keyinput36), .B1(keyinput60), .B2(n7828), 
        .ZN(n6477) );
  OAI221_X1 U8163 ( .B1(n6478), .B2(keyinput36), .C1(n7828), .C2(keyinput60), 
        .A(n6477), .ZN(n6479) );
  NOR4_X1 U8164 ( .A1(n6482), .A2(n6481), .A3(n6480), .A4(n6479), .ZN(n6509)
         );
  INV_X1 U8165 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6931) );
  AOI22_X1 U8166 ( .A1(n6931), .A2(keyinput54), .B1(n6484), .B2(keyinput63), 
        .ZN(n6483) );
  OAI221_X1 U8167 ( .B1(n6931), .B2(keyinput54), .C1(n6484), .C2(keyinput63), 
        .A(n6483), .ZN(n6494) );
  INV_X1 U8168 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n6486) );
  AOI22_X1 U8169 ( .A1(n6815), .A2(keyinput51), .B1(keyinput39), .B2(n6486), 
        .ZN(n6485) );
  OAI221_X1 U8170 ( .B1(n6815), .B2(keyinput51), .C1(n6486), .C2(keyinput39), 
        .A(n6485), .ZN(n6493) );
  AOI22_X1 U8171 ( .A1(n6488), .A2(keyinput16), .B1(n7260), .B2(keyinput58), 
        .ZN(n6487) );
  OAI221_X1 U8172 ( .B1(n6488), .B2(keyinput16), .C1(n7260), .C2(keyinput58), 
        .A(n6487), .ZN(n6492) );
  AOI22_X1 U8173 ( .A1(n8817), .A2(keyinput52), .B1(keyinput28), .B2(n6490), 
        .ZN(n6489) );
  OAI221_X1 U8174 ( .B1(n8817), .B2(keyinput52), .C1(n6490), .C2(keyinput28), 
        .A(n6489), .ZN(n6491) );
  NOR4_X1 U8175 ( .A1(n6494), .A2(n6493), .A3(n6492), .A4(n6491), .ZN(n6508)
         );
  INV_X1 U8176 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n6497) );
  INV_X1 U8177 ( .A(keyinput1), .ZN(n6496) );
  OAI22_X1 U8178 ( .A1(n6497), .A2(keyinput45), .B1(n6496), .B2(
        P2_ADDR_REG_5__SCAN_IN), .ZN(n6495) );
  AOI221_X1 U8179 ( .B1(n6497), .B2(keyinput45), .C1(P2_ADDR_REG_5__SCAN_IN), 
        .C2(n6496), .A(n6495), .ZN(n6506) );
  INV_X1 U8180 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n6500) );
  INV_X1 U8181 ( .A(keyinput19), .ZN(n6499) );
  OAI22_X1 U8182 ( .A1(n6500), .A2(keyinput3), .B1(n6499), .B2(
        P2_ADDR_REG_7__SCAN_IN), .ZN(n6498) );
  AOI221_X1 U8183 ( .B1(n6500), .B2(keyinput3), .C1(P2_ADDR_REG_7__SCAN_IN), 
        .C2(n6499), .A(n6498), .ZN(n6505) );
  INV_X1 U8184 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n9954) );
  OAI22_X1 U8185 ( .A1(n9954), .A2(keyinput43), .B1(n9246), .B2(keyinput7), 
        .ZN(n6501) );
  AOI221_X1 U8186 ( .B1(n9954), .B2(keyinput43), .C1(keyinput7), .C2(n9246), 
        .A(n6501), .ZN(n6504) );
  INV_X1 U8187 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6813) );
  OAI22_X1 U8188 ( .A1(n7113), .A2(keyinput27), .B1(n6813), .B2(keyinput38), 
        .ZN(n6502) );
  AOI221_X1 U8189 ( .B1(n7113), .B2(keyinput27), .C1(keyinput38), .C2(n6813), 
        .A(n6502), .ZN(n6503) );
  AND4_X1 U8190 ( .A1(n6506), .A2(n6505), .A3(n6504), .A4(n6503), .ZN(n6507)
         );
  AND3_X1 U8191 ( .A1(n6509), .A2(n6508), .A3(n6507), .ZN(n6510) );
  NAND4_X1 U8192 ( .A1(n6513), .A2(n6512), .A3(n6511), .A4(n6510), .ZN(n6514)
         );
  XNOR2_X1 U8193 ( .A(n6515), .B(n6514), .ZN(P2_U3244) );
  INV_X1 U8194 ( .A(n8650), .ZN(n6746) );
  AOI22_X1 U8195 ( .A1(n9624), .A2(n8323), .B1(n4388), .B2(n9339), .ZN(n9216)
         );
  NAND2_X1 U8196 ( .A1(n6526), .A2(n6544), .ZN(n6521) );
  NAND2_X1 U8197 ( .A1(n6521), .A2(n6520), .ZN(n6892) );
  INV_X1 U8198 ( .A(n6892), .ZN(n6522) );
  NAND2_X1 U8199 ( .A1(n6522), .A2(n4311), .ZN(n6527) );
  INV_X1 U8200 ( .A(n6544), .ZN(n6546) );
  NAND2_X1 U8201 ( .A1(n6765), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n6523) );
  OAI21_X1 U8202 ( .B1(n6524), .B2(n6546), .A(n6523), .ZN(n6525) );
  AOI21_X1 U8203 ( .B1(n6526), .B2(n8324), .A(n6525), .ZN(n6890) );
  NAND2_X1 U8204 ( .A1(n6890), .A2(n6892), .ZN(n6891) );
  NAND2_X1 U8205 ( .A1(n6527), .A2(n6891), .ZN(n6534) );
  NAND2_X1 U8206 ( .A1(n6529), .A2(n6544), .ZN(n6530) );
  NAND2_X1 U8207 ( .A1(n6531), .A2(n6530), .ZN(n6532) );
  NAND2_X1 U8208 ( .A1(n6535), .A2(n7004), .ZN(n6992) );
  INV_X1 U8209 ( .A(n6992), .ZN(n6539) );
  NAND2_X1 U8210 ( .A1(n6529), .A2(n4388), .ZN(n6537) );
  OR2_X1 U8211 ( .A1(n4393), .A2(n6727), .ZN(n6536) );
  NAND2_X1 U8212 ( .A1(n6537), .A2(n6536), .ZN(n6993) );
  OAI22_X1 U8213 ( .A1(n7202), .A2(n4312), .B1(n7368), .B2(n6716), .ZN(n6540)
         );
  XNOR2_X1 U8214 ( .A(n6540), .B(n4311), .ZN(n6542) );
  INV_X2 U8215 ( .A(n8324), .ZN(n6740) );
  OAI22_X1 U8216 ( .A1(n7202), .A2(n6740), .B1(n7368), .B2(n6727), .ZN(n6541)
         );
  NAND2_X1 U8217 ( .A1(n6542), .A2(n6541), .ZN(n6543) );
  OAI22_X1 U8218 ( .A1(n7350), .A2(n6727), .B1(n7455), .B2(n6716), .ZN(n6545)
         );
  XNOR2_X1 U8219 ( .A(n6545), .B(n4311), .ZN(n6548) );
  OAI22_X1 U8220 ( .A1(n7350), .A2(n6740), .B1(n7455), .B2(n6727), .ZN(n6547)
         );
  NAND2_X1 U8221 ( .A1(n6548), .A2(n6547), .ZN(n6549) );
  NAND2_X1 U8222 ( .A1(n9227), .A2(n6550), .ZN(n7192) );
  OAI22_X1 U8223 ( .A1(n7287), .A2(n6727), .B1(n9961), .B2(n6716), .ZN(n6552)
         );
  XNOR2_X1 U8224 ( .A(n6552), .B(n6738), .ZN(n6553) );
  OAI22_X1 U8225 ( .A1(n7287), .A2(n6740), .B1(n9961), .B2(n6727), .ZN(n6554)
         );
  XNOR2_X1 U8226 ( .A(n6553), .B(n6554), .ZN(n7193) );
  INV_X1 U8227 ( .A(n6553), .ZN(n6555) );
  OAI22_X1 U8228 ( .A1(n7438), .A2(n6727), .B1(n7386), .B2(n6716), .ZN(n6557)
         );
  XNOR2_X1 U8229 ( .A(n6557), .B(n6738), .ZN(n6560) );
  OR2_X1 U8230 ( .A1(n7438), .A2(n6740), .ZN(n6559) );
  NAND2_X1 U8231 ( .A1(n9925), .A2(n8323), .ZN(n6558) );
  NAND2_X1 U8232 ( .A1(n6559), .A2(n6558), .ZN(n6561) );
  INV_X1 U8233 ( .A(n6561), .ZN(n7379) );
  AND2_X1 U8234 ( .A1(n6560), .A2(n7379), .ZN(n6565) );
  INV_X1 U8235 ( .A(n6560), .ZN(n7377) );
  NAND2_X1 U8236 ( .A1(n7377), .A2(n6561), .ZN(n6563) );
  OAI22_X1 U8237 ( .A1(n8431), .A2(n6727), .B1(n9967), .B2(n6716), .ZN(n6562)
         );
  XNOR2_X1 U8238 ( .A(n6562), .B(n4311), .ZN(n6567) );
  OAI22_X1 U8239 ( .A1(n8431), .A2(n6740), .B1(n9967), .B2(n6727), .ZN(n6566)
         );
  NAND2_X1 U8240 ( .A1(n6567), .A2(n6566), .ZN(n7414) );
  AND2_X1 U8241 ( .A1(n6563), .A2(n7414), .ZN(n6564) );
  OR2_X1 U8242 ( .A1(n6567), .A2(n6566), .ZN(n7415) );
  OR2_X1 U8243 ( .A1(n8438), .A2(n6740), .ZN(n6569) );
  NAND2_X1 U8244 ( .A1(n8441), .A2(n8323), .ZN(n6568) );
  NAND2_X1 U8245 ( .A1(n6569), .A2(n6568), .ZN(n7298) );
  NAND2_X1 U8246 ( .A1(n8441), .A2(n8329), .ZN(n6571) );
  OAI21_X1 U8247 ( .B1(n8438), .B2(n6727), .A(n6571), .ZN(n6572) );
  XNOR2_X1 U8248 ( .A(n6572), .B(n4311), .ZN(n7299) );
  AND2_X1 U8249 ( .A1(n7415), .A2(n7299), .ZN(n6573) );
  NAND2_X1 U8250 ( .A1(n6574), .A2(n6573), .ZN(n6578) );
  INV_X1 U8251 ( .A(n7299), .ZN(n6576) );
  INV_X1 U8252 ( .A(n7298), .ZN(n6575) );
  OR2_X1 U8253 ( .A1(n6576), .A2(n6575), .ZN(n6577) );
  NAND2_X1 U8254 ( .A1(n7498), .A2(n8329), .ZN(n6582) );
  OR2_X1 U8255 ( .A1(n7589), .A2(n6727), .ZN(n6581) );
  NAND2_X1 U8256 ( .A1(n6582), .A2(n6581), .ZN(n6583) );
  XNOR2_X1 U8257 ( .A(n6583), .B(n6738), .ZN(n7426) );
  NAND2_X1 U8258 ( .A1(n7498), .A2(n8323), .ZN(n6585) );
  OR2_X1 U8259 ( .A1(n7589), .A2(n6740), .ZN(n6584) );
  AND2_X1 U8260 ( .A1(n6585), .A2(n6584), .ZN(n6587) );
  NAND2_X1 U8261 ( .A1(n7426), .A2(n6587), .ZN(n6586) );
  INV_X1 U8262 ( .A(n7426), .ZN(n6588) );
  INV_X1 U8263 ( .A(n6587), .ZN(n7425) );
  NAND2_X1 U8264 ( .A1(n6588), .A2(n7425), .ZN(n6589) );
  NAND2_X1 U8265 ( .A1(n7698), .A2(n8329), .ZN(n6592) );
  NAND2_X1 U8266 ( .A1(n9350), .A2(n8323), .ZN(n6591) );
  NAND2_X1 U8267 ( .A1(n6592), .A2(n6591), .ZN(n6593) );
  XNOR2_X1 U8268 ( .A(n6593), .B(n6738), .ZN(n6595) );
  AND2_X1 U8269 ( .A1(n9350), .A2(n4388), .ZN(n6594) );
  AOI21_X1 U8270 ( .B1(n7698), .B2(n8323), .A(n6594), .ZN(n6596) );
  NAND2_X1 U8271 ( .A1(n6595), .A2(n6596), .ZN(n7688) );
  INV_X1 U8272 ( .A(n6595), .ZN(n6598) );
  INV_X1 U8273 ( .A(n6596), .ZN(n6597) );
  NAND2_X1 U8274 ( .A1(n6598), .A2(n6597), .ZN(n6599) );
  NAND2_X1 U8275 ( .A1(n7688), .A2(n6599), .ZN(n7681) );
  NAND2_X1 U8276 ( .A1(n6600), .A2(n8329), .ZN(n6602) );
  NAND2_X1 U8277 ( .A1(n9753), .A2(n8323), .ZN(n6601) );
  NAND2_X1 U8278 ( .A1(n6602), .A2(n6601), .ZN(n6603) );
  XNOR2_X1 U8279 ( .A(n6603), .B(n6738), .ZN(n6618) );
  AND2_X1 U8280 ( .A1(n9753), .A2(n4388), .ZN(n6604) );
  AOI21_X1 U8281 ( .B1(n6600), .B2(n8323), .A(n6604), .ZN(n6619) );
  XNOR2_X1 U8282 ( .A(n6618), .B(n6619), .ZN(n7766) );
  INV_X1 U8283 ( .A(n7766), .ZN(n6612) );
  NAND2_X1 U8284 ( .A1(n7707), .A2(n8329), .ZN(n6606) );
  NAND2_X1 U8285 ( .A1(n9349), .A2(n8323), .ZN(n6605) );
  NAND2_X1 U8286 ( .A1(n6606), .A2(n6605), .ZN(n6607) );
  XNOR2_X1 U8287 ( .A(n6607), .B(n4311), .ZN(n6615) );
  INV_X1 U8288 ( .A(n6615), .ZN(n6611) );
  NAND2_X1 U8289 ( .A1(n7707), .A2(n8323), .ZN(n6609) );
  NAND2_X1 U8290 ( .A1(n9349), .A2(n4388), .ZN(n6608) );
  NAND2_X1 U8291 ( .A1(n6609), .A2(n6608), .ZN(n6614) );
  INV_X1 U8292 ( .A(n6614), .ZN(n6610) );
  NAND2_X1 U8293 ( .A1(n6611), .A2(n6610), .ZN(n7764) );
  AND2_X1 U8294 ( .A1(n6612), .A2(n7764), .ZN(n6613) );
  AND2_X1 U8295 ( .A1(n7688), .A2(n6613), .ZN(n6617) );
  INV_X1 U8296 ( .A(n6613), .ZN(n6616) );
  NAND2_X1 U8297 ( .A1(n6615), .A2(n6614), .ZN(n7762) );
  INV_X1 U8298 ( .A(n6618), .ZN(n6621) );
  INV_X1 U8299 ( .A(n6619), .ZN(n6620) );
  NAND2_X1 U8300 ( .A1(n6621), .A2(n6620), .ZN(n6622) );
  NAND2_X1 U8301 ( .A1(n7768), .A2(n6622), .ZN(n7807) );
  NAND2_X1 U8302 ( .A1(n9761), .A2(n8329), .ZN(n6624) );
  NAND2_X1 U8303 ( .A1(n9348), .A2(n8323), .ZN(n6623) );
  NAND2_X1 U8304 ( .A1(n6624), .A2(n6623), .ZN(n6625) );
  XNOR2_X1 U8305 ( .A(n6625), .B(n6738), .ZN(n7809) );
  NOR2_X1 U8306 ( .A1(n7772), .A2(n6740), .ZN(n6626) );
  AOI21_X1 U8307 ( .B1(n9761), .B2(n8323), .A(n6626), .ZN(n6628) );
  NAND2_X1 U8308 ( .A1(n7809), .A2(n6628), .ZN(n6627) );
  NAND2_X1 U8309 ( .A1(n7807), .A2(n6627), .ZN(n6631) );
  INV_X1 U8310 ( .A(n7809), .ZN(n6629) );
  INV_X1 U8311 ( .A(n6628), .ZN(n7808) );
  NAND2_X1 U8312 ( .A1(n6629), .A2(n7808), .ZN(n6630) );
  NAND2_X1 U8313 ( .A1(n7904), .A2(n8329), .ZN(n6633) );
  NAND2_X1 U8314 ( .A1(n9752), .A2(n8323), .ZN(n6632) );
  NAND2_X1 U8315 ( .A1(n6633), .A2(n6632), .ZN(n6634) );
  XNOR2_X1 U8316 ( .A(n6634), .B(n4311), .ZN(n6637) );
  NAND2_X1 U8317 ( .A1(n7904), .A2(n8323), .ZN(n6636) );
  NAND2_X1 U8318 ( .A1(n9752), .A2(n4388), .ZN(n6635) );
  NAND2_X1 U8319 ( .A1(n6636), .A2(n6635), .ZN(n6638) );
  AND2_X1 U8320 ( .A1(n6637), .A2(n6638), .ZN(n7832) );
  INV_X1 U8321 ( .A(n6637), .ZN(n6640) );
  INV_X1 U8322 ( .A(n6638), .ZN(n6639) );
  NAND2_X1 U8323 ( .A1(n6640), .A2(n6639), .ZN(n7831) );
  NAND2_X1 U8324 ( .A1(n9669), .A2(n8329), .ZN(n6642) );
  NAND2_X1 U8325 ( .A1(n9347), .A2(n8323), .ZN(n6641) );
  NAND2_X1 U8326 ( .A1(n6642), .A2(n6641), .ZN(n6643) );
  XNOR2_X1 U8327 ( .A(n6643), .B(n6738), .ZN(n6649) );
  NAND2_X1 U8328 ( .A1(n6650), .A2(n6649), .ZN(n8089) );
  NAND2_X1 U8329 ( .A1(n9669), .A2(n8323), .ZN(n6645) );
  NAND2_X1 U8330 ( .A1(n9347), .A2(n4388), .ZN(n6644) );
  NAND2_X1 U8331 ( .A1(n6645), .A2(n6644), .ZN(n8088) );
  NAND2_X2 U8332 ( .A1(n8089), .A2(n8088), .ZN(n8093) );
  NAND2_X1 U8333 ( .A1(n9662), .A2(n8329), .ZN(n6647) );
  NAND2_X1 U8334 ( .A1(n9346), .A2(n8323), .ZN(n6646) );
  NAND2_X1 U8335 ( .A1(n6647), .A2(n6646), .ZN(n6648) );
  XNOR2_X1 U8336 ( .A(n6648), .B(n6738), .ZN(n6653) );
  NAND2_X1 U8337 ( .A1(n9662), .A2(n8323), .ZN(n6652) );
  NAND2_X1 U8338 ( .A1(n9346), .A2(n4388), .ZN(n6651) );
  NAND2_X1 U8339 ( .A1(n6652), .A2(n6651), .ZN(n8104) );
  NAND2_X1 U8340 ( .A1(n8093), .A2(n8090), .ZN(n6655) );
  INV_X1 U8341 ( .A(n6653), .ZN(n6654) );
  NAND2_X1 U8342 ( .A1(n5294), .A2(n8329), .ZN(n6657) );
  OR2_X1 U8343 ( .A1(n9570), .A2(n4312), .ZN(n6656) );
  NAND2_X1 U8344 ( .A1(n6657), .A2(n6656), .ZN(n6658) );
  XNOR2_X1 U8345 ( .A(n6658), .B(n4311), .ZN(n8170) );
  NAND2_X1 U8346 ( .A1(n5294), .A2(n8323), .ZN(n6660) );
  OR2_X1 U8347 ( .A1(n9570), .A2(n6740), .ZN(n6659) );
  NAND2_X1 U8348 ( .A1(n6660), .A2(n6659), .ZN(n8171) );
  INV_X1 U8349 ( .A(n9260), .ZN(n6666) );
  NAND2_X1 U8350 ( .A1(n9654), .A2(n8329), .ZN(n6662) );
  NAND2_X1 U8351 ( .A1(n9344), .A2(n8323), .ZN(n6661) );
  NAND2_X1 U8352 ( .A1(n6662), .A2(n6661), .ZN(n6663) );
  XNOR2_X1 U8353 ( .A(n6663), .B(n6738), .ZN(n6668) );
  AND2_X1 U8354 ( .A1(n9344), .A2(n4388), .ZN(n6664) );
  AOI21_X1 U8355 ( .B1(n9654), .B2(n8323), .A(n6664), .ZN(n6667) );
  XNOR2_X1 U8356 ( .A(n6668), .B(n6667), .ZN(n9263) );
  INV_X1 U8357 ( .A(n9263), .ZN(n6665) );
  NAND2_X1 U8358 ( .A1(n6668), .A2(n6667), .ZN(n6669) );
  NAND2_X1 U8359 ( .A1(n9647), .A2(n8329), .ZN(n6671) );
  NAND2_X1 U8360 ( .A1(n9577), .A2(n8323), .ZN(n6670) );
  NAND2_X1 U8361 ( .A1(n6671), .A2(n6670), .ZN(n6672) );
  XNOR2_X1 U8362 ( .A(n6672), .B(n6738), .ZN(n6676) );
  NAND2_X1 U8363 ( .A1(n9647), .A2(n8323), .ZN(n6674) );
  NAND2_X1 U8364 ( .A1(n9577), .A2(n4388), .ZN(n6673) );
  NAND2_X1 U8365 ( .A1(n6674), .A2(n6673), .ZN(n9306) );
  INV_X1 U8366 ( .A(n6676), .ZN(n6677) );
  NAND2_X1 U8367 ( .A1(n9644), .A2(n8329), .ZN(n6679) );
  NAND2_X1 U8368 ( .A1(n9343), .A2(n8323), .ZN(n6678) );
  NAND2_X1 U8369 ( .A1(n6679), .A2(n6678), .ZN(n6680) );
  XNOR2_X1 U8370 ( .A(n6680), .B(n6738), .ZN(n6682) );
  AND2_X1 U8371 ( .A1(n9343), .A2(n4388), .ZN(n6681) );
  AOI21_X1 U8372 ( .B1(n9644), .B2(n8323), .A(n6681), .ZN(n6683) );
  NAND2_X1 U8373 ( .A1(n6682), .A2(n6683), .ZN(n9280) );
  INV_X1 U8374 ( .A(n6682), .ZN(n6685) );
  INV_X1 U8375 ( .A(n6683), .ZN(n6684) );
  NAND2_X1 U8376 ( .A1(n6685), .A2(n6684), .ZN(n6686) );
  AND2_X1 U8377 ( .A1(n9280), .A2(n6686), .ZN(n9236) );
  NAND2_X1 U8378 ( .A1(n9637), .A2(n8329), .ZN(n6688) );
  NAND2_X1 U8379 ( .A1(n9342), .A2(n8323), .ZN(n6687) );
  NAND2_X1 U8380 ( .A1(n6688), .A2(n6687), .ZN(n6689) );
  XNOR2_X1 U8381 ( .A(n6689), .B(n6738), .ZN(n6691) );
  AND2_X1 U8382 ( .A1(n9342), .A2(n4388), .ZN(n6690) );
  AOI21_X1 U8383 ( .B1(n9637), .B2(n8323), .A(n6690), .ZN(n6692) );
  NAND2_X1 U8384 ( .A1(n6691), .A2(n6692), .ZN(n6697) );
  INV_X1 U8385 ( .A(n6691), .ZN(n6694) );
  INV_X1 U8386 ( .A(n6692), .ZN(n6693) );
  NAND2_X1 U8387 ( .A1(n6694), .A2(n6693), .ZN(n6695) );
  AND2_X1 U8388 ( .A1(n6697), .A2(n6695), .ZN(n9281) );
  NAND2_X1 U8389 ( .A1(n9634), .A2(n8329), .ZN(n6699) );
  NAND2_X1 U8390 ( .A1(n9341), .A2(n8323), .ZN(n6698) );
  NAND2_X1 U8391 ( .A1(n6699), .A2(n6698), .ZN(n6700) );
  XNOR2_X1 U8392 ( .A(n6700), .B(n4311), .ZN(n6702) );
  NOR2_X1 U8393 ( .A1(n9538), .A2(n6740), .ZN(n6701) );
  AOI21_X1 U8394 ( .B1(n9634), .B2(n8323), .A(n6701), .ZN(n6703) );
  XNOR2_X1 U8395 ( .A(n6702), .B(n6703), .ZN(n9244) );
  INV_X1 U8396 ( .A(n6702), .ZN(n6704) );
  NAND2_X1 U8397 ( .A1(n6704), .A2(n6703), .ZN(n6705) );
  OR2_X1 U8398 ( .A1(n9512), .A2(n4312), .ZN(n6707) );
  OR2_X1 U8399 ( .A1(n9522), .A2(n6740), .ZN(n6706) );
  AND2_X1 U8400 ( .A1(n6707), .A2(n6706), .ZN(n6710) );
  OAI22_X1 U8401 ( .A1(n9512), .A2(n6716), .B1(n9522), .B2(n6727), .ZN(n6708)
         );
  XNOR2_X1 U8402 ( .A(n6708), .B(n4311), .ZN(n9292) );
  INV_X1 U8403 ( .A(n6710), .ZN(n6711) );
  NAND2_X2 U8404 ( .A1(n6712), .A2(n6711), .ZN(n9294) );
  OAI22_X1 U8405 ( .A1(n6713), .A2(n6716), .B1(n9505), .B2(n4312), .ZN(n6714)
         );
  XNOR2_X1 U8406 ( .A(n6714), .B(n4311), .ZN(n6715) );
  OAI22_X1 U8407 ( .A1(n8350), .A2(n6716), .B1(n9491), .B2(n6727), .ZN(n6717)
         );
  XOR2_X1 U8408 ( .A(n4311), .B(n6717), .Z(n6719) );
  AOI22_X1 U8409 ( .A1(n9619), .A2(n8323), .B1(n4388), .B2(n9338), .ZN(n6718)
         );
  NAND2_X1 U8410 ( .A1(n6719), .A2(n6718), .ZN(n6720) );
  OAI21_X1 U8411 ( .B1(n6719), .B2(n6718), .A(n6720), .ZN(n9271) );
  INV_X1 U8412 ( .A(n6720), .ZN(n6721) );
  NAND2_X1 U8413 ( .A1(n9612), .A2(n8329), .ZN(n6723) );
  OR2_X1 U8414 ( .A1(n9477), .A2(n6727), .ZN(n6722) );
  NAND2_X1 U8415 ( .A1(n6723), .A2(n6722), .ZN(n6724) );
  XNOR2_X1 U8416 ( .A(n6724), .B(n4311), .ZN(n6726) );
  OAI22_X1 U8417 ( .A1(n9463), .A2(n4312), .B1(n9477), .B2(n6740), .ZN(n6725)
         );
  XNOR2_X1 U8418 ( .A(n6726), .B(n6725), .ZN(n9252) );
  NOR2_X1 U8419 ( .A1(n6726), .A2(n6725), .ZN(n9319) );
  NAND2_X1 U8420 ( .A1(n9607), .A2(n8329), .ZN(n6729) );
  OR2_X1 U8421 ( .A1(n9465), .A2(n4312), .ZN(n6728) );
  NAND2_X1 U8422 ( .A1(n6729), .A2(n6728), .ZN(n6730) );
  XNOR2_X1 U8423 ( .A(n6730), .B(n6738), .ZN(n6732) );
  NOR2_X1 U8424 ( .A1(n9465), .A2(n6740), .ZN(n6731) );
  AOI21_X1 U8425 ( .B1(n9607), .B2(n6544), .A(n6731), .ZN(n6733) );
  XNOR2_X1 U8426 ( .A(n6732), .B(n6733), .ZN(n9318) );
  INV_X1 U8427 ( .A(n6732), .ZN(n6735) );
  INV_X1 U8428 ( .A(n6733), .ZN(n6734) );
  NAND2_X1 U8429 ( .A1(n9601), .A2(n8329), .ZN(n6737) );
  INV_X1 U8430 ( .A(n9450), .ZN(n9336) );
  NAND2_X1 U8431 ( .A1(n9336), .A2(n8323), .ZN(n6736) );
  NAND2_X1 U8432 ( .A1(n6737), .A2(n6736), .ZN(n6739) );
  XNOR2_X1 U8433 ( .A(n6739), .B(n6738), .ZN(n6743) );
  NOR2_X1 U8434 ( .A1(n9450), .A2(n6740), .ZN(n6741) );
  AOI21_X1 U8435 ( .B1(n9601), .B2(n8323), .A(n6741), .ZN(n6742) );
  NAND2_X1 U8436 ( .A1(n6743), .A2(n6742), .ZN(n8335) );
  OAI21_X1 U8437 ( .B1(n6743), .B2(n6742), .A(n8335), .ZN(n6744) );
  AND2_X2 U8438 ( .A1(n7025), .A2(n6746), .ZN(n9670) );
  OR2_X1 U8439 ( .A1(n9670), .A2(n6747), .ZN(n6749) );
  INV_X1 U8440 ( .A(n6970), .ZN(n9694) );
  INV_X1 U8441 ( .A(n6913), .ZN(n9693) );
  NAND3_X1 U8442 ( .A1(n9694), .A2(n9693), .A3(n6912), .ZN(n6751) );
  INV_X1 U8443 ( .A(n9951), .ZN(n6748) );
  OR2_X1 U8444 ( .A1(n7210), .A2(n8640), .ZN(n6750) );
  NAND2_X1 U8445 ( .A1(n6973), .A2(n6751), .ZN(n6896) );
  INV_X1 U8446 ( .A(n8653), .ZN(n6752) );
  NAND2_X1 U8447 ( .A1(n6753), .A2(n6752), .ZN(n6754) );
  NAND2_X1 U8448 ( .A1(n6754), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6755) );
  INV_X1 U8449 ( .A(n6758), .ZN(n6761) );
  NOR2_X1 U8450 ( .A1(n8659), .A2(n6951), .ZN(n6756) );
  OR2_X1 U8451 ( .A1(n8659), .A2(n5522), .ZN(n6757) );
  NOR2_X2 U8452 ( .A1(n6758), .A2(n6757), .ZN(n9308) );
  AOI22_X1 U8453 ( .A1(n9337), .A2(n9308), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n6759) );
  OAI21_X1 U8454 ( .B1(n9438), .B2(n9325), .A(n6759), .ZN(n6760) );
  AOI21_X1 U8455 ( .B1(n9434), .B2(n9329), .A(n6760), .ZN(n6764) );
  NAND2_X1 U8456 ( .A1(n6761), .A2(n9926), .ZN(n6762) );
  NAND2_X1 U8457 ( .A1(n9601), .A2(n9313), .ZN(n6763) );
  NAND2_X1 U8458 ( .A1(n6765), .A2(n7954), .ZN(n6832) );
  OR2_X2 U8459 ( .A1(n6832), .A2(P1_U3084), .ZN(n9358) );
  INV_X1 U8460 ( .A(n7954), .ZN(n6766) );
  OR2_X1 U8461 ( .A1(n6767), .A2(n6766), .ZN(n6768) );
  NAND2_X1 U8462 ( .A1(n6768), .A2(n6832), .ZN(n6846) );
  OR2_X1 U8463 ( .A1(n6846), .A2(n6769), .ZN(n6770) );
  NAND2_X1 U8464 ( .A1(n6770), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U8465 ( .A(n10045), .ZN(n6771) );
  XNOR2_X1 U8466 ( .A(n6773), .B(n6772), .ZN(n6774) );
  NOR2_X1 U8467 ( .A1(n6774), .A2(n8836), .ZN(n6779) );
  AND2_X1 U8468 ( .A1(n8834), .A2(n7986), .ZN(n6778) );
  NOR2_X1 U8469 ( .A1(n10006), .A2(n7887), .ZN(n6777) );
  INV_X1 U8470 ( .A(n8800), .ZN(n8734) );
  NAND2_X1 U8471 ( .A1(n8734), .A2(n9070), .ZN(n8818) );
  NAND2_X1 U8472 ( .A1(n8821), .A2(n8853), .ZN(n6775) );
  NAND2_X1 U8473 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n8864) );
  OAI211_X1 U8474 ( .C1(n8818), .C2(n9994), .A(n6775), .B(n8864), .ZN(n6776)
         );
  OR4_X1 U8475 ( .A1(n6779), .A2(n6778), .A3(n6777), .A4(n6776), .ZN(P2_U3219)
         );
  INV_X1 U8476 ( .A(n6780), .ZN(n6785) );
  AOI21_X1 U8477 ( .B1(n6784), .B2(n6782), .A(n6781), .ZN(n6783) );
  AOI211_X1 U8478 ( .C1(n6785), .C2(n6784), .A(n8836), .B(n6783), .ZN(n6792)
         );
  AND2_X1 U8479 ( .A1(n8834), .A2(n7957), .ZN(n6791) );
  NOR2_X1 U8480 ( .A1(n10006), .A2(n7867), .ZN(n6790) );
  NAND2_X1 U8481 ( .A1(n8821), .A2(n8854), .ZN(n6788) );
  NOR2_X1 U8482 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6786), .ZN(n7154) );
  INV_X1 U8483 ( .A(n7154), .ZN(n6787) );
  OAI211_X1 U8484 ( .C1(n8818), .C2(n7517), .A(n6788), .B(n6787), .ZN(n6789)
         );
  OR4_X1 U8485 ( .A1(n6792), .A2(n6791), .A3(n6790), .A4(n6789), .ZN(P2_U3233)
         );
  NOR2_X1 U8486 ( .A1(n6799), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9210) );
  INV_X2 U8487 ( .A(n9210), .ZN(n8661) );
  NAND2_X1 U8488 ( .A1(n6799), .A2(P2_U3152), .ZN(n9212) );
  INV_X1 U8489 ( .A(n7049), .ZN(n7073) );
  OAI222_X1 U8490 ( .A1(n8661), .A2(n6793), .B1(n9212), .B2(n6801), .C1(
        P2_U3152), .C2(n7073), .ZN(P2_U3355) );
  INV_X1 U8491 ( .A(n9730), .ZN(n7051) );
  OAI222_X1 U8492 ( .A1(n8661), .A2(n6794), .B1(n9212), .B2(n6811), .C1(
        P2_U3152), .C2(n7051), .ZN(P2_U3356) );
  INV_X1 U8493 ( .A(n7047), .ZN(n7085) );
  OAI222_X1 U8494 ( .A1(n8661), .A2(n6795), .B1(n9212), .B2(n6803), .C1(
        P2_U3152), .C2(n7085), .ZN(P2_U3354) );
  INV_X1 U8495 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6796) );
  CLKBUF_X1 U8496 ( .A(n9212), .Z(n8665) );
  INV_X1 U8497 ( .A(n7033), .ZN(n9718) );
  OAI222_X1 U8498 ( .A1(n8661), .A2(n6796), .B1(n8665), .B2(n6809), .C1(
        P2_U3152), .C2(n9718), .ZN(P2_U3357) );
  INV_X1 U8499 ( .A(n7091), .ZN(n7061) );
  OAI222_X1 U8500 ( .A1(n8661), .A2(n6797), .B1(n8665), .B2(n6807), .C1(
        P2_U3152), .C2(n7061), .ZN(P2_U3353) );
  INV_X1 U8501 ( .A(n7121), .ZN(n7099) );
  OAI222_X1 U8502 ( .A1(n8661), .A2(n6798), .B1(n8665), .B2(n6805), .C1(
        P2_U3152), .C2(n7099), .ZN(P2_U3352) );
  NAND2_X1 U8503 ( .A1(n5400), .A2(P1_U3084), .ZN(n9707) );
  INV_X1 U8504 ( .A(n9707), .ZN(n8243) );
  INV_X1 U8505 ( .A(n8243), .ZN(n9699) );
  INV_X1 U8506 ( .A(n9704), .ZN(n9697) );
  AOI22_X1 U8507 ( .A1(n6909), .A2(P1_STATE_REG_SCAN_IN), .B1(n9697), .B2(
        P2_DATAO_REG_3__SCAN_IN), .ZN(n6800) );
  OAI21_X1 U8508 ( .B1(n6801), .B2(n9699), .A(n6800), .ZN(P1_U3350) );
  INV_X1 U8509 ( .A(n6955), .ZN(n6967) );
  OAI222_X1 U8510 ( .A1(n6967), .A2(P1_U3084), .B1(n9699), .B2(n6803), .C1(
        n6802), .C2(n9704), .ZN(P1_U3349) );
  INV_X1 U8511 ( .A(n6933), .ZN(n6842) );
  OAI222_X1 U8512 ( .A1(n6842), .A2(P1_U3084), .B1(n9699), .B2(n6805), .C1(
        n6804), .C2(n9704), .ZN(P1_U3347) );
  OAI222_X1 U8513 ( .A1(n6808), .A2(P1_U3084), .B1(n9699), .B2(n6807), .C1(
        n6806), .C2(n9704), .ZN(P1_U3348) );
  OAI222_X1 U8514 ( .A1(n5079), .A2(P1_U3084), .B1(n9707), .B2(n6809), .C1(
        n4818), .C2(n9704), .ZN(P1_U3352) );
  OAI222_X1 U8515 ( .A1(n5068), .A2(P1_U3084), .B1(n9699), .B2(n6811), .C1(
        n6810), .C2(n9704), .ZN(P1_U3351) );
  INV_X1 U8516 ( .A(n6934), .ZN(n9836) );
  INV_X1 U8517 ( .A(n6812), .ZN(n6814) );
  OAI222_X1 U8518 ( .A1(n9836), .A2(P1_U3084), .B1(n9699), .B2(n6814), .C1(
        n6813), .C2(n9704), .ZN(P1_U3346) );
  OAI222_X1 U8519 ( .A1(n8661), .A2(n6815), .B1(n9212), .B2(n6814), .C1(
        P2_U3152), .C2(n7127), .ZN(P2_U3351) );
  NAND2_X1 U8520 ( .A1(n6816), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6821) );
  NAND2_X1 U8521 ( .A1(n6817), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6820) );
  NAND2_X1 U8522 ( .A1(n6818), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6819) );
  NAND3_X1 U8523 ( .A1(n6821), .A2(n6820), .A3(n6819), .ZN(n9403) );
  NAND2_X1 U8524 ( .A1(n9403), .A2(P1_U4006), .ZN(n6822) );
  OAI21_X1 U8525 ( .B1(P1_U4006), .B2(n6184), .A(n6822), .ZN(P1_U3586) );
  INV_X1 U8526 ( .A(n6823), .ZN(n6826) );
  AOI22_X1 U8527 ( .A1(n9853), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9697), .ZN(n6824) );
  OAI21_X1 U8528 ( .B1(n6826), .B2(n9699), .A(n6824), .ZN(P1_U3345) );
  OAI222_X1 U8529 ( .A1(n8661), .A2(n6827), .B1(n8665), .B2(n6826), .C1(
        P2_U3152), .C2(n6825), .ZN(P2_U3350) );
  OAI21_X1 U8530 ( .B1(n10035), .B2(n7326), .A(n5805), .ZN(n6829) );
  INV_X1 U8531 ( .A(n7952), .ZN(n7040) );
  NAND2_X1 U8532 ( .A1(n10035), .A2(n7040), .ZN(n6828) );
  NAND2_X1 U8533 ( .A1(n6829), .A2(n6828), .ZN(n9714) );
  NOR2_X1 U8534 ( .A1(n10013), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8535 ( .A(n6830), .ZN(n6869) );
  AOI22_X1 U8536 ( .A1(n9874), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9697), .ZN(n6831) );
  OAI21_X1 U8537 ( .B1(n6869), .B2(n9699), .A(n6831), .ZN(P1_U3344) );
  INV_X1 U8538 ( .A(n6832), .ZN(n6833) );
  OR2_X1 U8539 ( .A1(P1_U3083), .A2(n6833), .ZN(n9922) );
  INV_X1 U8540 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6868) );
  INV_X1 U8541 ( .A(n6948), .ZN(n6947) );
  NAND2_X1 U8542 ( .A1(n6947), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9799) );
  NOR2_X1 U8543 ( .A1(n6846), .A2(n9799), .ZN(n9395) );
  NAND2_X1 U8544 ( .A1(n9395), .A2(n5522), .ZN(n9837) );
  INV_X1 U8545 ( .A(n9837), .ZN(n9915) );
  NAND2_X1 U8546 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n9819), .ZN(n6841) );
  XNOR2_X1 U8547 ( .A(n4313), .B(n5057), .ZN(n9812) );
  INV_X1 U8548 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6834) );
  MUX2_X1 U8549 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n6834), .S(n6849), .Z(n6880)
         );
  AND2_X1 U8550 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6881) );
  NAND2_X1 U8551 ( .A1(n6880), .A2(n6881), .ZN(n6879) );
  NAND2_X1 U8552 ( .A1(n6849), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6835) );
  NAND2_X1 U8553 ( .A1(n6879), .A2(n6835), .ZN(n9813) );
  NAND2_X1 U8554 ( .A1(n9812), .A2(n9813), .ZN(n6837) );
  NAND2_X1 U8555 ( .A1(n4313), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6836) );
  NAND2_X1 U8556 ( .A1(n6837), .A2(n6836), .ZN(n6901) );
  MUX2_X1 U8557 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n5100), .S(n6909), .Z(n6900)
         );
  NAND2_X1 U8558 ( .A1(n6901), .A2(n6900), .ZN(n6899) );
  NAND2_X1 U8559 ( .A1(n6909), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6838) );
  NAND2_X1 U8560 ( .A1(n6899), .A2(n6838), .ZN(n6954) );
  INV_X1 U8561 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6839) );
  MUX2_X1 U8562 ( .A(n6839), .B(P1_REG1_REG_4__SCAN_IN), .S(n6955), .Z(n6840)
         );
  OAI21_X1 U8563 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n6955), .A(n6956), .ZN(
        n9829) );
  INV_X1 U8564 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7297) );
  MUX2_X1 U8565 ( .A(n7297), .B(P1_REG1_REG_5__SCAN_IN), .S(n9819), .Z(n9828)
         );
  INV_X1 U8566 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9985) );
  AOI22_X1 U8567 ( .A1(n6933), .A2(n9985), .B1(P1_REG1_REG_6__SCAN_IN), .B2(
        n6842), .ZN(n6843) );
  NOR2_X1 U8568 ( .A1(n6844), .A2(n6843), .ZN(n6920) );
  AOI21_X1 U8569 ( .B1(n6844), .B2(n6843), .A(n6920), .ZN(n6865) );
  NOR2_X1 U8570 ( .A1(n5522), .A2(P1_U3084), .ZN(n9798) );
  NAND2_X1 U8571 ( .A1(n9798), .A2(n6948), .ZN(n6845) );
  NAND2_X1 U8572 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3084), .ZN(n7418) );
  INV_X1 U8573 ( .A(n6846), .ZN(n9803) );
  NAND2_X1 U8574 ( .A1(n9798), .A2(n6947), .ZN(n8654) );
  INV_X1 U8575 ( .A(n8654), .ZN(n6847) );
  INV_X1 U8576 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6848) );
  XNOR2_X1 U8577 ( .A(n4313), .B(n6848), .ZN(n9811) );
  INV_X1 U8578 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7219) );
  AND2_X1 U8579 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n6950) );
  NAND2_X1 U8580 ( .A1(n6849), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6850) );
  NAND2_X1 U8581 ( .A1(n6876), .A2(n6850), .ZN(n9810) );
  NAND2_X1 U8582 ( .A1(n9811), .A2(n9810), .ZN(n9809) );
  NAND2_X1 U8583 ( .A1(n4313), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6852) );
  NAND2_X1 U8584 ( .A1(n9809), .A2(n6852), .ZN(n6904) );
  INV_X1 U8585 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6853) );
  XNOR2_X1 U8586 ( .A(n6909), .B(n6853), .ZN(n6905) );
  NAND2_X1 U8587 ( .A1(n6904), .A2(n6905), .ZN(n6903) );
  NAND2_X1 U8588 ( .A1(n6909), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6854) );
  NAND2_X1 U8589 ( .A1(n6903), .A2(n6854), .ZN(n6962) );
  MUX2_X1 U8590 ( .A(n6855), .B(P1_REG2_REG_4__SCAN_IN), .S(n6955), .Z(n6961)
         );
  OR2_X1 U8591 ( .A1(n6962), .A2(n6961), .ZN(n9821) );
  OR2_X1 U8592 ( .A1(n6955), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9822) );
  NAND2_X1 U8593 ( .A1(n9821), .A2(n9822), .ZN(n6856) );
  NOR2_X1 U8594 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n9819), .ZN(n6857) );
  AOI21_X1 U8595 ( .B1(n9819), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6857), .ZN(
        n9823) );
  NAND2_X1 U8596 ( .A1(n6856), .A2(n9823), .ZN(n9820) );
  INV_X1 U8597 ( .A(n6857), .ZN(n6858) );
  NAND2_X1 U8598 ( .A1(n9820), .A2(n6858), .ZN(n6862) );
  OR2_X1 U8599 ( .A1(n6933), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6860) );
  NAND2_X1 U8600 ( .A1(n6933), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6859) );
  NAND2_X1 U8601 ( .A1(n6860), .A2(n6859), .ZN(n6861) );
  NOR2_X1 U8602 ( .A1(n6862), .A2(n6861), .ZN(n6932) );
  AOI21_X1 U8603 ( .B1(n6862), .B2(n6861), .A(n6932), .ZN(n6863) );
  NAND2_X1 U8604 ( .A1(n9862), .A2(n6863), .ZN(n6864) );
  OAI211_X1 U8605 ( .C1(n6865), .C2(n9879), .A(n7418), .B(n6864), .ZN(n6866)
         );
  AOI21_X1 U8606 ( .B1(n6933), .B2(n9915), .A(n6866), .ZN(n6867) );
  OAI21_X1 U8607 ( .B1(n9922), .B2(n6868), .A(n6867), .ZN(P1_U3247) );
  OAI222_X1 U8608 ( .A1(n8661), .A2(n6870), .B1(n7272), .B2(P2_U3152), .C1(
        n9212), .C2(n6869), .ZN(P2_U3349) );
  NAND2_X1 U8609 ( .A1(n8913), .A2(P2_U3966), .ZN(n6871) );
  OAI21_X1 U8610 ( .B1(P2_U3966), .B2(n6185), .A(n6871), .ZN(P2_U3583) );
  INV_X1 U8611 ( .A(n6872), .ZN(n6874) );
  OAI222_X1 U8612 ( .A1(P1_U3084), .A2(n6943), .B1(n9707), .B2(n6874), .C1(
        n6873), .C2(n9704), .ZN(P1_U3343) );
  OAI222_X1 U8613 ( .A1(n8661), .A2(n6875), .B1(n8865), .B2(P2_U3152), .C1(
        n8665), .C2(n6874), .ZN(P2_U3348) );
  OAI211_X1 U8614 ( .C1(n6877), .C2(n6950), .A(n9862), .B(n6876), .ZN(n6878)
         );
  OAI21_X1 U8615 ( .B1(n9837), .B2(n5079), .A(n6878), .ZN(n6885) );
  INV_X1 U8616 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6883) );
  OAI211_X1 U8617 ( .C1(n6881), .C2(n6880), .A(n9917), .B(n6879), .ZN(n6882)
         );
  OAI21_X1 U8618 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6883), .A(n6882), .ZN(n6884) );
  AOI211_X1 U8619 ( .C1(n9854), .C2(P1_ADDR_REG_1__SCAN_IN), .A(n6885), .B(
        n6884), .ZN(n6886) );
  INV_X1 U8620 ( .A(n6886), .ZN(P1_U3242) );
  INV_X1 U8621 ( .A(n7166), .ZN(n7162) );
  INV_X1 U8622 ( .A(n5765), .ZN(n6888) );
  OAI222_X1 U8623 ( .A1(P1_U3084), .A2(n7162), .B1(n9707), .B2(n6888), .C1(
        n6887), .C2(n9704), .ZN(P1_U3342) );
  OAI222_X1 U8624 ( .A1(n8661), .A2(n6889), .B1(n7530), .B2(P2_U3152), .C1(
        n9212), .C2(n6888), .ZN(P2_U3347) );
  CLKBUF_X1 U8625 ( .A(n6890), .Z(n6893) );
  OAI21_X1 U8626 ( .B1(n6893), .B2(n6892), .A(n6891), .ZN(n6894) );
  INV_X1 U8627 ( .A(n6894), .ZN(n6949) );
  AND2_X1 U8628 ( .A1(n6896), .A2(n6895), .ZN(n7014) );
  INV_X1 U8629 ( .A(n7014), .ZN(n6996) );
  OAI22_X1 U8630 ( .A1(n9332), .A2(n6524), .B1(n7134), .B2(n9325), .ZN(n6897)
         );
  AOI21_X1 U8631 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n6996), .A(n6897), .ZN(
        n6898) );
  OAI21_X1 U8632 ( .B1(n6949), .B2(n9315), .A(n6898), .ZN(P1_U3230) );
  INV_X1 U8633 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6911) );
  OAI211_X1 U8634 ( .C1(n6901), .C2(n6900), .A(n9917), .B(n6899), .ZN(n6902)
         );
  OAI21_X1 U8635 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n5101), .A(n6902), .ZN(n6908) );
  OAI211_X1 U8636 ( .C1(n6905), .C2(n6904), .A(n9862), .B(n6903), .ZN(n6906)
         );
  INV_X1 U8637 ( .A(n6906), .ZN(n6907) );
  AOI211_X1 U8638 ( .C1(n9915), .C2(n6909), .A(n6908), .B(n6907), .ZN(n6910)
         );
  OAI21_X1 U8639 ( .B1(n9922), .B2(n6911), .A(n6910), .ZN(P1_U3244) );
  NAND2_X1 U8640 ( .A1(n6913), .A2(n6912), .ZN(n6971) );
  NOR2_X1 U8641 ( .A1(n9694), .A2(n6971), .ZN(n6914) );
  INV_X1 U8642 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6919) );
  INV_X1 U8643 ( .A(n7025), .ZN(n6917) );
  XNOR2_X1 U8644 ( .A(n6526), .B(n6519), .ZN(n8567) );
  NAND2_X1 U8645 ( .A1(n6917), .A2(n8659), .ZN(n6915) );
  OAI22_X1 U8646 ( .A1(n8567), .A2(n6915), .B1(n7134), .B2(n9550), .ZN(n9939)
         );
  INV_X1 U8647 ( .A(n9939), .ZN(n6916) );
  OAI21_X1 U8648 ( .B1(n6524), .B2(n6917), .A(n6916), .ZN(n6974) );
  NAND2_X1 U8649 ( .A1(n6974), .A2(n9983), .ZN(n6918) );
  OAI21_X1 U8650 ( .B1(n9983), .B2(n6919), .A(n6918), .ZN(P1_U3454) );
  NOR2_X1 U8651 ( .A1(n9874), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6927) );
  OR2_X1 U8652 ( .A1(n9853), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6925) );
  NOR2_X1 U8653 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6934), .ZN(n6923) );
  NOR2_X1 U8654 ( .A1(n6933), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6921) );
  INV_X1 U8655 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6922) );
  MUX2_X1 U8656 ( .A(n6922), .B(P1_REG1_REG_7__SCAN_IN), .S(n6934), .Z(n9842)
         );
  NOR2_X1 U8657 ( .A1(n9843), .A2(n9842), .ZN(n9841) );
  NOR2_X1 U8658 ( .A1(n6923), .A2(n9841), .ZN(n9857) );
  MUX2_X1 U8659 ( .A(n9988), .B(P1_REG1_REG_8__SCAN_IN), .S(n9853), .Z(n9856)
         );
  NOR2_X1 U8660 ( .A1(n9857), .A2(n9856), .ZN(n9855) );
  INV_X1 U8661 ( .A(n9855), .ZN(n6924) );
  INV_X1 U8662 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6926) );
  MUX2_X1 U8663 ( .A(n6926), .B(P1_REG1_REG_9__SCAN_IN), .S(n9874), .Z(n9877)
         );
  NOR2_X1 U8664 ( .A1(n9876), .A2(n9877), .ZN(n9875) );
  INV_X1 U8665 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7711) );
  AOI22_X1 U8666 ( .A1(n6982), .A2(n7711), .B1(P1_REG1_REG_10__SCAN_IN), .B2(
        n6943), .ZN(n6928) );
  NOR2_X1 U8667 ( .A1(n6929), .A2(n6928), .ZN(n6976) );
  AOI21_X1 U8668 ( .B1(n6929), .B2(n6928), .A(n6976), .ZN(n6946) );
  MUX2_X1 U8669 ( .A(n6455), .B(P1_REG2_REG_9__SCAN_IN), .S(n9874), .Z(n9870)
         );
  NOR2_X1 U8670 ( .A1(n9853), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6930) );
  AOI21_X1 U8671 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n9853), .A(n6930), .ZN(
        n9860) );
  AOI22_X1 U8672 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6934), .B1(n9836), .B2(
        n6931), .ZN(n9847) );
  OAI21_X1 U8673 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n9853), .A(n9859), .ZN(
        n9871) );
  NOR2_X1 U8674 ( .A1(n9870), .A2(n9871), .ZN(n9869) );
  AOI21_X1 U8675 ( .B1(n9874), .B2(P1_REG2_REG_9__SCAN_IN), .A(n9869), .ZN(
        n6939) );
  INV_X1 U8676 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6935) );
  NAND2_X1 U8677 ( .A1(n6943), .A2(n6935), .ZN(n6937) );
  NAND2_X1 U8678 ( .A1(n6982), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6936) );
  NAND2_X1 U8679 ( .A1(n6937), .A2(n6936), .ZN(n6938) );
  AOI21_X1 U8680 ( .B1(n6939), .B2(n6938), .A(n6981), .ZN(n6941) );
  NAND2_X1 U8681 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3084), .ZN(n7690) );
  INV_X1 U8682 ( .A(n7690), .ZN(n6940) );
  AOI21_X1 U8683 ( .B1(n9862), .B2(n6941), .A(n6940), .ZN(n6942) );
  OAI21_X1 U8684 ( .B1(n9837), .B2(n6943), .A(n6942), .ZN(n6944) );
  AOI21_X1 U8685 ( .B1(n9854), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n6944), .ZN(
        n6945) );
  OAI21_X1 U8686 ( .B1(n6946), .B2(n9879), .A(n6945), .ZN(P1_U3251) );
  INV_X1 U8687 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9944) );
  AOI21_X1 U8688 ( .B1(n6947), .B2(n9944), .A(n5522), .ZN(n9797) );
  MUX2_X1 U8689 ( .A(n6950), .B(n6949), .S(n6948), .Z(n6952) );
  NAND2_X1 U8690 ( .A1(n6952), .A2(n6951), .ZN(n6953) );
  OAI211_X1 U8691 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n9797), .A(n6953), .B(
        P1_U4006), .ZN(n9817) );
  INV_X1 U8692 ( .A(n6954), .ZN(n6958) );
  MUX2_X1 U8693 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6839), .S(n6955), .Z(n6957)
         );
  OAI21_X1 U8694 ( .B1(n6958), .B2(n6957), .A(n6956), .ZN(n6960) );
  NAND2_X1 U8695 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3084), .ZN(n7195) );
  INV_X1 U8696 ( .A(n7195), .ZN(n6959) );
  AOI21_X1 U8697 ( .B1(n9917), .B2(n6960), .A(n6959), .ZN(n6966) );
  NAND2_X1 U8698 ( .A1(n6962), .A2(n6961), .ZN(n6963) );
  NAND2_X1 U8699 ( .A1(n9821), .A2(n6963), .ZN(n6964) );
  NAND2_X1 U8700 ( .A1(n9862), .A2(n6964), .ZN(n6965) );
  OAI211_X1 U8701 ( .C1(n9837), .C2(n6967), .A(n6966), .B(n6965), .ZN(n6968)
         );
  AOI21_X1 U8702 ( .B1(n9854), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n6968), .ZN(
        n6969) );
  NAND2_X1 U8703 ( .A1(n9817), .A2(n6969), .ZN(P1_U3245) );
  NOR2_X1 U8704 ( .A1(n6971), .A2(n6970), .ZN(n6972) );
  INV_X1 U8705 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9804) );
  NAND2_X1 U8706 ( .A1(n6974), .A2(n9990), .ZN(n6975) );
  OAI21_X1 U8707 ( .B1(n9990), .B2(n9804), .A(n6975), .ZN(P1_U3523) );
  NOR2_X1 U8708 ( .A1(n6982), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6977) );
  NOR2_X1 U8709 ( .A1(n6977), .A2(n6976), .ZN(n6979) );
  INV_X1 U8710 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9789) );
  AOI22_X1 U8711 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n7162), .B1(n7166), .B2(
        n9789), .ZN(n6978) );
  NOR2_X1 U8712 ( .A1(n6979), .A2(n6978), .ZN(n7161) );
  AOI21_X1 U8713 ( .B1(n6979), .B2(n6978), .A(n7161), .ZN(n6990) );
  INV_X1 U8714 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6980) );
  AOI22_X1 U8715 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n7166), .B1(n7162), .B2(
        n6980), .ZN(n6984) );
  OAI21_X1 U8716 ( .B1(n6984), .B2(n6983), .A(n7165), .ZN(n6988) );
  INV_X1 U8717 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n6986) );
  NAND2_X1 U8718 ( .A1(n9915), .A2(n7166), .ZN(n6985) );
  NAND2_X1 U8719 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3084), .ZN(n7770) );
  OAI211_X1 U8720 ( .C1(n6986), .C2(n9922), .A(n6985), .B(n7770), .ZN(n6987)
         );
  AOI21_X1 U8721 ( .B1(n6988), .B2(n9862), .A(n6987), .ZN(n6989) );
  OAI21_X1 U8722 ( .B1(n6990), .B2(n9879), .A(n6989), .ZN(P1_U3252) );
  INV_X1 U8723 ( .A(n6991), .ZN(n7006) );
  AOI21_X1 U8724 ( .B1(n6993), .B2(n6992), .A(n7006), .ZN(n6998) );
  INV_X1 U8725 ( .A(n9325), .ZN(n9264) );
  AOI22_X1 U8726 ( .A1(n9264), .A2(n9357), .B1(n9308), .B2(n6526), .ZN(n6994)
         );
  OAI21_X1 U8727 ( .B1(n4393), .B2(n9332), .A(n6994), .ZN(n6995) );
  AOI21_X1 U8728 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n6996), .A(n6995), .ZN(
        n6997) );
  OAI21_X1 U8729 ( .B1(n6998), .B2(n9315), .A(n6997), .ZN(P1_U3220) );
  INV_X1 U8730 ( .A(n6999), .ZN(n7002) );
  OAI222_X1 U8731 ( .A1(n8661), .A2(n7000), .B1(n8665), .B2(n7002), .C1(
        P2_U3152), .C2(n7645), .ZN(P2_U3346) );
  INV_X1 U8732 ( .A(n7249), .ZN(n7243) );
  OAI222_X1 U8733 ( .A1(n7243), .A2(P1_U3084), .B1(n9707), .B2(n7002), .C1(
        n7001), .C2(n9704), .ZN(P1_U3341) );
  INV_X1 U8734 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7013) );
  INV_X1 U8735 ( .A(n7004), .ZN(n7005) );
  NOR3_X1 U8736 ( .A1(n7006), .A2(n7003), .A3(n7005), .ZN(n7008) );
  AND2_X1 U8737 ( .A1(n7007), .A2(n7003), .ZN(n9226) );
  OAI21_X1 U8738 ( .B1(n7008), .B2(n9226), .A(n9322), .ZN(n7012) );
  OAI22_X1 U8739 ( .A1(n9326), .A2(n7134), .B1(n7350), .B2(n9325), .ZN(n7009)
         );
  AOI21_X1 U8740 ( .B1(n7010), .B2(n9313), .A(n7009), .ZN(n7011) );
  OAI211_X1 U8741 ( .C1(n7014), .C2(n7013), .A(n7012), .B(n7011), .ZN(P1_U3235) );
  INV_X1 U8742 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7029) );
  OR2_X1 U8743 ( .A1(n8558), .A2(n7015), .ZN(n7017) );
  NAND3_X1 U8744 ( .A1(n8555), .A2(n8640), .A3(n8650), .ZN(n7016) );
  OAI21_X1 U8745 ( .B1(n7018), .B2(n7020), .A(n7019), .ZN(n7218) );
  OAI21_X1 U8746 ( .B1(n7023), .B2(n7022), .A(n7021), .ZN(n7024) );
  AOI222_X1 U8747 ( .A1(n9747), .A2(n7024), .B1(n9357), .B2(n9751), .C1(n6526), 
        .C2(n9754), .ZN(n7217) );
  OAI21_X1 U8748 ( .B1(n4393), .B2(n6524), .A(n9764), .ZN(n7026) );
  NOR2_X1 U8749 ( .A1(n7026), .A2(n7133), .ZN(n7215) );
  AOI21_X1 U8750 ( .B1(n9670), .B2(n5084), .A(n7215), .ZN(n7027) );
  OAI211_X1 U8751 ( .C1(n9672), .C2(n7218), .A(n7217), .B(n7027), .ZN(n7030)
         );
  NAND2_X1 U8752 ( .A1(n7030), .A2(n9983), .ZN(n7028) );
  OAI21_X1 U8753 ( .B1(n9983), .B2(n7029), .A(n7028), .ZN(P1_U3457) );
  INV_X2 U8754 ( .A(n9987), .ZN(n9990) );
  NAND2_X1 U8755 ( .A1(n7030), .A2(n9990), .ZN(n7031) );
  OAI21_X1 U8756 ( .B1(n9990), .B2(n6834), .A(n7031), .ZN(P1_U3524) );
  INV_X1 U8757 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7333) );
  AOI21_X1 U8758 ( .B1(n7033), .B2(P2_REG2_REG_1__SCAN_IN), .A(n9710), .ZN(
        n9728) );
  NAND2_X1 U8759 ( .A1(P2_REG2_REG_2__SCAN_IN), .A2(n9730), .ZN(n7034) );
  OAI21_X1 U8760 ( .B1(n9730), .B2(P2_REG2_REG_2__SCAN_IN), .A(n7034), .ZN(
        n9727) );
  NOR2_X1 U8761 ( .A1(n9728), .A2(n9727), .ZN(n9726) );
  AOI21_X1 U8762 ( .B1(n9730), .B2(P2_REG2_REG_2__SCAN_IN), .A(n9726), .ZN(
        n7066) );
  NAND2_X1 U8763 ( .A1(n7049), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7035) );
  OAI21_X1 U8764 ( .B1(n7049), .B2(P2_REG2_REG_3__SCAN_IN), .A(n7035), .ZN(
        n7065) );
  NOR2_X1 U8765 ( .A1(n7066), .A2(n7065), .ZN(n7064) );
  AOI21_X1 U8766 ( .B1(n7049), .B2(P2_REG2_REG_3__SCAN_IN), .A(n7064), .ZN(
        n7078) );
  NAND2_X1 U8767 ( .A1(P2_REG2_REG_4__SCAN_IN), .A2(n7047), .ZN(n7036) );
  OAI21_X1 U8768 ( .B1(n7047), .B2(P2_REG2_REG_4__SCAN_IN), .A(n7036), .ZN(
        n7077) );
  NAND2_X1 U8769 ( .A1(P2_REG2_REG_5__SCAN_IN), .A2(n7091), .ZN(n7037) );
  OAI21_X1 U8770 ( .B1(n7091), .B2(P2_REG2_REG_5__SCAN_IN), .A(n7037), .ZN(
        n7044) );
  OR2_X1 U8771 ( .A1(n7038), .A2(P2_U3152), .ZN(n7039) );
  OAI211_X1 U8772 ( .C1(n10035), .C2(n7041), .A(n7040), .B(n7039), .ZN(n7042)
         );
  NAND2_X1 U8773 ( .A1(n7042), .A2(n5805), .ZN(n7055) );
  NAND2_X1 U8774 ( .A1(n7055), .A2(n8862), .ZN(n7046) );
  NOR2_X1 U8775 ( .A1(n8663), .A2(n8687), .ZN(n7043) );
  AOI211_X1 U8776 ( .C1(n7045), .C2(n7044), .A(n7088), .B(n9725), .ZN(n7063)
         );
  NAND2_X1 U8777 ( .A1(n7046), .A2(n8663), .ZN(n10009) );
  NAND2_X1 U8778 ( .A1(P2_REG1_REG_4__SCAN_IN), .A2(n7047), .ZN(n7053) );
  MUX2_X1 U8779 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n7048), .S(n7047), .Z(n7080)
         );
  NAND2_X1 U8780 ( .A1(n7049), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7052) );
  MUX2_X1 U8781 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n7050), .S(n7049), .Z(n7068)
         );
  XNOR2_X1 U8782 ( .A(n7051), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n9734) );
  XNOR2_X1 U8783 ( .A(n9718), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n9722) );
  NAND3_X1 U8784 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .A3(n9722), .ZN(n9720) );
  OAI21_X1 U8785 ( .B1(n9718), .B2(n10108), .A(n9720), .ZN(n9733) );
  NAND2_X1 U8786 ( .A1(n9734), .A2(n9733), .ZN(n9732) );
  OAI21_X1 U8787 ( .B1(n7051), .B2(n10110), .A(n9732), .ZN(n7069) );
  NAND2_X1 U8788 ( .A1(n7068), .A2(n7069), .ZN(n7067) );
  NAND2_X1 U8789 ( .A1(n7052), .A2(n7067), .ZN(n7081) );
  NAND2_X1 U8790 ( .A1(n7080), .A2(n7081), .ZN(n7079) );
  NAND2_X1 U8791 ( .A1(n7053), .A2(n7079), .ZN(n7058) );
  MUX2_X1 U8792 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n7054), .S(n7091), .Z(n7057)
         );
  INV_X1 U8793 ( .A(n7055), .ZN(n7056) );
  NAND2_X1 U8794 ( .A1(n7056), .A2(n8687), .ZN(n10011) );
  NAND2_X1 U8795 ( .A1(n7057), .A2(n7058), .ZN(n7092) );
  OAI211_X1 U8796 ( .C1(n7058), .C2(n7057), .A(n10007), .B(n7092), .ZN(n7060)
         );
  AND2_X1 U8797 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3152), .ZN(n7392) );
  AOI21_X1 U8798 ( .B1(n10013), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n7392), .ZN(
        n7059) );
  OAI211_X1 U8799 ( .C1(n10009), .C2(n7061), .A(n7060), .B(n7059), .ZN(n7062)
         );
  OR2_X1 U8800 ( .A1(n7063), .A2(n7062), .ZN(P2_U3250) );
  AOI211_X1 U8801 ( .C1(n7066), .C2(n7065), .A(n7064), .B(n9725), .ZN(n7075)
         );
  OAI211_X1 U8802 ( .C1(n7069), .C2(n7068), .A(n10007), .B(n7067), .ZN(n7072)
         );
  NOR2_X1 U8803 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7229), .ZN(n7070) );
  AOI21_X1 U8804 ( .B1(n10013), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n7070), .ZN(
        n7071) );
  OAI211_X1 U8805 ( .C1(n10009), .C2(n7073), .A(n7072), .B(n7071), .ZN(n7074)
         );
  OR2_X1 U8806 ( .A1(n7075), .A2(n7074), .ZN(P2_U3248) );
  AOI211_X1 U8807 ( .C1(n7078), .C2(n7077), .A(n7076), .B(n9725), .ZN(n7087)
         );
  OAI211_X1 U8808 ( .C1(n7081), .C2(n7080), .A(n10007), .B(n7079), .ZN(n7084)
         );
  NAND2_X1 U8809 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n7315) );
  INV_X1 U8810 ( .A(n7315), .ZN(n7082) );
  AOI21_X1 U8811 ( .B1(n10013), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n7082), .ZN(
        n7083) );
  OAI211_X1 U8812 ( .C1(n10009), .C2(n7085), .A(n7084), .B(n7083), .ZN(n7086)
         );
  OR2_X1 U8813 ( .A1(n7087), .A2(n7086), .ZN(P2_U3249) );
  NAND2_X1 U8814 ( .A1(P2_REG2_REG_6__SCAN_IN), .A2(n7121), .ZN(n7089) );
  OAI21_X1 U8815 ( .B1(n7121), .B2(P2_REG2_REG_6__SCAN_IN), .A(n7089), .ZN(
        n7090) );
  NOR2_X1 U8816 ( .A1(n4335), .A2(n7090), .ZN(n7120) );
  AOI211_X1 U8817 ( .C1(n4335), .C2(n7090), .A(n7120), .B(n9725), .ZN(n7101)
         );
  NAND2_X1 U8818 ( .A1(P2_REG1_REG_5__SCAN_IN), .A2(n7091), .ZN(n7093) );
  NAND2_X1 U8819 ( .A1(n7093), .A2(n7092), .ZN(n7096) );
  MUX2_X1 U8820 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n7094), .S(n7121), .Z(n7095)
         );
  NAND2_X1 U8821 ( .A1(n7095), .A2(n7096), .ZN(n7114) );
  OAI211_X1 U8822 ( .C1(n7096), .C2(n7095), .A(n10007), .B(n7114), .ZN(n7098)
         );
  AND2_X1 U8823 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n7480) );
  AOI21_X1 U8824 ( .B1(n10013), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n7480), .ZN(
        n7097) );
  OAI211_X1 U8825 ( .C1(n10009), .C2(n7099), .A(n7098), .B(n7097), .ZN(n7100)
         );
  OR2_X1 U8826 ( .A1(n7101), .A2(n7100), .ZN(P2_U3251) );
  NOR2_X1 U8827 ( .A1(n7102), .A2(P2_U3152), .ZN(n7239) );
  NAND2_X1 U8828 ( .A1(n8863), .A2(n9070), .ZN(n7104) );
  NAND2_X1 U8829 ( .A1(n6115), .A2(n9068), .ZN(n7103) );
  NAND2_X1 U8830 ( .A1(n7104), .A2(n7103), .ZN(n7463) );
  AOI22_X1 U8831 ( .A1(n8834), .A2(n7546), .B1(n8734), .B2(n7463), .ZN(n7110)
         );
  OAI21_X1 U8832 ( .B1(n7107), .B2(n7106), .A(n7105), .ZN(n7108) );
  NAND2_X1 U8833 ( .A1(n7108), .A2(n10002), .ZN(n7109) );
  OAI211_X1 U8834 ( .C1(n7239), .C2(n7111), .A(n7110), .B(n7109), .ZN(P2_U3224) );
  INV_X1 U8835 ( .A(n7112), .ZN(n7129) );
  OAI222_X1 U8836 ( .A1(n8665), .A2(n7129), .B1(n7646), .B2(P2_U3152), .C1(
        n7113), .C2(n8661), .ZN(P2_U3345) );
  INV_X1 U8837 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7516) );
  NOR2_X1 U8838 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7516), .ZN(n7119) );
  NAND2_X1 U8839 ( .A1(P2_REG1_REG_6__SCAN_IN), .A2(n7121), .ZN(n7115) );
  AND2_X1 U8840 ( .A1(n7115), .A2(n7114), .ZN(n7117) );
  MUX2_X1 U8841 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n7828), .S(n7127), .Z(n7116)
         );
  NOR2_X1 U8842 ( .A1(n7117), .A2(n7116), .ZN(n7140) );
  AOI211_X1 U8843 ( .C1(n7117), .C2(n7116), .A(n7140), .B(n10011), .ZN(n7118)
         );
  AOI211_X1 U8844 ( .C1(n10013), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n7119), .B(
        n7118), .ZN(n7126) );
  XNOR2_X1 U8845 ( .A(n7148), .B(P2_REG2_REG_7__SCAN_IN), .ZN(n7122) );
  AOI211_X1 U8846 ( .C1(n7123), .C2(n7122), .A(n7147), .B(n9725), .ZN(n7124)
         );
  INV_X1 U8847 ( .A(n7124), .ZN(n7125) );
  OAI211_X1 U8848 ( .C1(n10009), .C2(n7127), .A(n7126), .B(n7125), .ZN(
        P2_U3252) );
  INV_X1 U8849 ( .A(n7611), .ZN(n7617) );
  OAI222_X1 U8850 ( .A1(P1_U3084), .A2(n7617), .B1(n9707), .B2(n7129), .C1(
        n7128), .C2(n9704), .ZN(P1_U3340) );
  INV_X1 U8851 ( .A(n7210), .ZN(n9980) );
  OAI21_X1 U8852 ( .B1(n7131), .B2(n8565), .A(n7130), .ZN(n7374) );
  INV_X1 U8853 ( .A(n7132), .ZN(n7208) );
  OAI21_X1 U8854 ( .B1(n7368), .B2(n7133), .A(n7208), .ZN(n7372) );
  OAI22_X1 U8855 ( .A1(n7372), .A2(n9975), .B1(n7368), .B2(n9973), .ZN(n7138)
         );
  XNOR2_X1 U8856 ( .A(n8565), .B(n8380), .ZN(n7137) );
  INV_X1 U8857 ( .A(n7493), .ZN(n9758) );
  OAI22_X1 U8858 ( .A1(n7134), .A2(n5531), .B1(n7350), .B2(n9550), .ZN(n7135)
         );
  AOI21_X1 U8859 ( .B1(n7374), .B2(n9758), .A(n7135), .ZN(n7136) );
  OAI21_X1 U8860 ( .B1(n9572), .B2(n7137), .A(n7136), .ZN(n7367) );
  AOI211_X1 U8861 ( .C1(n9980), .C2(n7374), .A(n7138), .B(n7367), .ZN(n9960)
         );
  NAND2_X1 U8862 ( .A1(n9987), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7139) );
  OAI21_X1 U8863 ( .B1(n9960), .B2(n9987), .A(n7139), .ZN(P1_U3525) );
  NAND2_X1 U8864 ( .A1(n7180), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7142) );
  AOI21_X1 U8865 ( .B1(n7148), .B2(P2_REG1_REG_7__SCAN_IN), .A(n7140), .ZN(
        n7175) );
  MUX2_X1 U8866 ( .A(n5716), .B(P2_REG1_REG_8__SCAN_IN), .S(n7180), .Z(n7174)
         );
  OR2_X1 U8867 ( .A1(n7175), .A2(n7174), .ZN(n7141) );
  NAND2_X1 U8868 ( .A1(n7142), .A2(n7141), .ZN(n7146) );
  INV_X1 U8869 ( .A(n7146), .ZN(n7144) );
  MUX2_X1 U8870 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n7271), .S(n7272), .Z(n7143)
         );
  AOI21_X1 U8871 ( .B1(n7144), .B2(n7143), .A(n10011), .ZN(n7153) );
  MUX2_X1 U8872 ( .A(n7271), .B(P2_REG1_REG_9__SCAN_IN), .S(n7272), .Z(n7145)
         );
  NAND2_X1 U8873 ( .A1(n7146), .A2(n7145), .ZN(n7270) );
  NAND2_X1 U8874 ( .A1(n7180), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7149) );
  OAI21_X1 U8875 ( .B1(n7180), .B2(P2_REG2_REG_8__SCAN_IN), .A(n7149), .ZN(
        n7177) );
  AOI21_X1 U8876 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n7180), .A(n7176), .ZN(
        n7151) );
  XOR2_X1 U8877 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n7272), .Z(n7150) );
  NOR2_X1 U8878 ( .A1(n7151), .A2(n7150), .ZN(n7262) );
  AOI211_X1 U8879 ( .C1(n7151), .C2(n7150), .A(n7262), .B(n9725), .ZN(n7152)
         );
  AOI21_X1 U8880 ( .B1(n7153), .B2(n7270), .A(n7152), .ZN(n7156) );
  AOI21_X1 U8881 ( .B1(n10013), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7154), .ZN(
        n7155) );
  OAI211_X1 U8882 ( .C1(n7272), .C2(n10009), .A(n7156), .B(n7155), .ZN(
        P2_U3254) );
  INV_X1 U8883 ( .A(n7157), .ZN(n7160) );
  OAI222_X1 U8884 ( .A1(n8665), .A2(n7160), .B1(n7943), .B2(P2_U3152), .C1(
        n7158), .C2(n8661), .ZN(P2_U3344) );
  INV_X1 U8885 ( .A(n7618), .ZN(n9370) );
  OAI222_X1 U8886 ( .A1(P1_U3084), .A2(n9370), .B1(n9707), .B2(n7160), .C1(
        n7159), .C2(n9704), .ZN(P1_U3339) );
  INV_X1 U8887 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9782) );
  AOI22_X1 U8888 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n7243), .B1(n7249), .B2(
        n9782), .ZN(n7163) );
  NOR2_X1 U8889 ( .A1(n7164), .A2(n7163), .ZN(n7242) );
  AOI21_X1 U8890 ( .B1(n7164), .B2(n7163), .A(n7242), .ZN(n7173) );
  NAND2_X1 U8891 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3084), .ZN(n7811) );
  OAI21_X1 U8892 ( .B1(n9837), .B2(n7243), .A(n7811), .ZN(n7171) );
  NAND2_X1 U8893 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7249), .ZN(n7167) );
  OAI21_X1 U8894 ( .B1(n7249), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7167), .ZN(
        n7168) );
  NOR2_X1 U8895 ( .A1(n7168), .A2(n7169), .ZN(n7248) );
  INV_X1 U8896 ( .A(n9862), .ZN(n9908) );
  AOI211_X1 U8897 ( .C1(n7169), .C2(n7168), .A(n7248), .B(n9908), .ZN(n7170)
         );
  AOI211_X1 U8898 ( .C1(n9854), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n7171), .B(
        n7170), .ZN(n7172) );
  OAI21_X1 U8899 ( .B1(n7173), .B2(n9879), .A(n7172), .ZN(P1_U3253) );
  XNOR2_X1 U8900 ( .A(n7175), .B(n7174), .ZN(n7184) );
  INV_X1 U8901 ( .A(n10009), .ZN(n9731) );
  AOI211_X1 U8902 ( .C1(n7178), .C2(n7177), .A(n7176), .B(n9725), .ZN(n7179)
         );
  AOI21_X1 U8903 ( .B1(n9731), .B2(n7180), .A(n7179), .ZN(n7183) );
  NAND2_X1 U8904 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n9993) );
  INV_X1 U8905 ( .A(n9993), .ZN(n7181) );
  AOI21_X1 U8906 ( .B1(n10013), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n7181), .ZN(
        n7182) );
  OAI211_X1 U8907 ( .C1(n10011), .C2(n7184), .A(n7183), .B(n7182), .ZN(
        P2_U3253) );
  NOR2_X1 U8908 ( .A1(n10000), .A2(n7467), .ZN(n7188) );
  MUX2_X1 U8909 ( .A(n7320), .B(n7467), .S(n7185), .Z(n7186) );
  AOI21_X1 U8910 ( .B1(n7461), .B2(n7186), .A(n8836), .ZN(n7187) );
  AOI211_X1 U8911 ( .C1(n8821), .C2(n8861), .A(n7188), .B(n7187), .ZN(n7189)
         );
  OAI21_X1 U8912 ( .B1(n7239), .B2(n4615), .A(n7189), .ZN(P2_U3234) );
  INV_X1 U8913 ( .A(n9329), .ZN(n9311) );
  INV_X1 U8914 ( .A(n7190), .ZN(n7361) );
  OAI21_X1 U8915 ( .B1(n7193), .B2(n7192), .A(n7191), .ZN(n7194) );
  NAND2_X1 U8916 ( .A1(n7194), .A2(n9322), .ZN(n7199) );
  NAND2_X1 U8917 ( .A1(n9356), .A2(n9308), .ZN(n7196) );
  OAI211_X1 U8918 ( .C1(n7438), .C2(n9325), .A(n7196), .B(n7195), .ZN(n7197)
         );
  AOI21_X1 U8919 ( .B1(n7357), .B2(n9313), .A(n7197), .ZN(n7198) );
  OAI211_X1 U8920 ( .C1(n9311), .C2(n7361), .A(n7199), .B(n7198), .ZN(P1_U3228) );
  OAI21_X1 U8921 ( .B1(n7201), .B2(n8564), .A(n7200), .ZN(n7457) );
  INV_X1 U8922 ( .A(n7457), .ZN(n7211) );
  OAI22_X1 U8923 ( .A1(n7287), .A2(n9550), .B1(n7202), .B2(n5531), .ZN(n7206)
         );
  XNOR2_X1 U8924 ( .A(n8564), .B(n7203), .ZN(n7204) );
  NOR2_X1 U8925 ( .A1(n7204), .A2(n9572), .ZN(n7205) );
  AOI211_X1 U8926 ( .C1(n9758), .C2(n7457), .A(n7206), .B(n7205), .ZN(n7459)
         );
  INV_X1 U8927 ( .A(n7358), .ZN(n7207) );
  AOI21_X1 U8928 ( .B1(n9230), .B2(n7208), .A(n7207), .ZN(n7452) );
  AOI22_X1 U8929 ( .A1(n7452), .A2(n9764), .B1(n9670), .B2(n9230), .ZN(n7209)
         );
  OAI211_X1 U8930 ( .C1(n7211), .C2(n7210), .A(n7459), .B(n7209), .ZN(n7213)
         );
  NAND2_X1 U8931 ( .A1(n7213), .A2(n9983), .ZN(n7212) );
  OAI21_X1 U8932 ( .B1(n9983), .B2(n5103), .A(n7212), .ZN(P1_U3463) );
  NAND2_X1 U8933 ( .A1(n7213), .A2(n9990), .ZN(n7214) );
  OAI21_X1 U8934 ( .B1(n9990), .B2(n5100), .A(n7214), .ZN(P1_U3526) );
  AOI22_X1 U8935 ( .A1(n7215), .A2(n9930), .B1(n9759), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n7216) );
  AOI21_X1 U8936 ( .B1(n7217), .B2(n7216), .A(n9578), .ZN(n7222) );
  NOR2_X1 U8937 ( .A1(n9582), .A2(n7218), .ZN(n7221) );
  OAI22_X1 U8938 ( .A1(n9568), .A2(n4393), .B1(n7219), .B2(n9945), .ZN(n7220)
         );
  OR3_X1 U8939 ( .A1(n7222), .A2(n7221), .A3(n7220), .ZN(P1_U3290) );
  NAND2_X1 U8940 ( .A1(n9358), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n7223) );
  OAI21_X1 U8941 ( .B1(n9477), .B2(n9358), .A(n7223), .ZN(P1_U3580) );
  XNOR2_X1 U8942 ( .A(n7225), .B(n7224), .ZN(n7231) );
  OAI22_X1 U8943 ( .A1(n10000), .A2(n10062), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7229), .ZN(n7228) );
  OAI22_X1 U8944 ( .A1(n9995), .A2(n7555), .B1(n7226), .B2(n8818), .ZN(n7227)
         );
  AOI211_X1 U8945 ( .C1(n8789), .C2(n7229), .A(n7228), .B(n7227), .ZN(n7230)
         );
  OAI21_X1 U8946 ( .B1(n8836), .B2(n7231), .A(n7230), .ZN(P2_U3220) );
  OAI22_X1 U8947 ( .A1(n9995), .A2(n8699), .B1(n10058), .B2(n10000), .ZN(n7232) );
  AOI21_X1 U8948 ( .B1(n9998), .B2(n8861), .A(n7232), .ZN(n7238) );
  OAI21_X1 U8949 ( .B1(n7235), .B2(n7234), .A(n7233), .ZN(n7236) );
  NAND2_X1 U8950 ( .A1(n7236), .A2(n10002), .ZN(n7237) );
  OAI211_X1 U8951 ( .C1(n7239), .C2(n8705), .A(n7238), .B(n7237), .ZN(P2_U3239) );
  INV_X1 U8952 ( .A(n7240), .ZN(n7307) );
  AOI22_X1 U8953 ( .A1(n9900), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n9697), .ZN(n7241) );
  OAI21_X1 U8954 ( .B1(n7307), .B2(n9699), .A(n7241), .ZN(P1_U3337) );
  AOI21_X1 U8955 ( .B1(n9782), .B2(n7243), .A(n7242), .ZN(n7245) );
  INV_X1 U8956 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9776) );
  AOI22_X1 U8957 ( .A1(P1_REG1_REG_13__SCAN_IN), .A2(n7617), .B1(n7611), .B2(
        n9776), .ZN(n7244) );
  NOR2_X1 U8958 ( .A1(n7245), .A2(n7244), .ZN(n7616) );
  AOI21_X1 U8959 ( .B1(n7245), .B2(n7244), .A(n7616), .ZN(n7257) );
  OR2_X1 U8960 ( .A1(n7611), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7247) );
  NAND2_X1 U8961 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n7611), .ZN(n7246) );
  NAND2_X1 U8962 ( .A1(n7247), .A2(n7246), .ZN(n7251) );
  AOI21_X1 U8963 ( .B1(n7251), .B2(n7250), .A(n7610), .ZN(n7253) );
  NAND2_X1 U8964 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7836) );
  INV_X1 U8965 ( .A(n7836), .ZN(n7252) );
  AOI21_X1 U8966 ( .B1(n9862), .B2(n7253), .A(n7252), .ZN(n7254) );
  OAI21_X1 U8967 ( .B1(n9837), .B2(n7617), .A(n7254), .ZN(n7255) );
  AOI21_X1 U8968 ( .B1(n9854), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n7255), .ZN(
        n7256) );
  OAI21_X1 U8969 ( .B1(n7257), .B2(n9879), .A(n7256), .ZN(P1_U3254) );
  INV_X1 U8970 ( .A(n7258), .ZN(n7261) );
  INV_X1 U8971 ( .A(n8183), .ZN(n8189) );
  OAI222_X1 U8972 ( .A1(n8661), .A2(n7259), .B1(n8665), .B2(n7261), .C1(
        P2_U3152), .C2(n8189), .ZN(P2_U3343) );
  INV_X1 U8973 ( .A(n9888), .ZN(n9374) );
  OAI222_X1 U8974 ( .A1(n9374), .A2(P1_U3084), .B1(n9707), .B2(n7261), .C1(
        n7260), .C2(n9704), .ZN(P1_U3338) );
  INV_X1 U8975 ( .A(n7272), .ZN(n7263) );
  AOI21_X1 U8976 ( .B1(n7263), .B2(P2_REG2_REG_9__SCAN_IN), .A(n7262), .ZN(
        n8872) );
  NAND2_X1 U8977 ( .A1(n7268), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7264) );
  OAI21_X1 U8978 ( .B1(n7268), .B2(P2_REG2_REG_10__SCAN_IN), .A(n7264), .ZN(
        n8871) );
  MUX2_X1 U8979 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n8016), .S(n7530), .Z(n7265)
         );
  INV_X1 U8980 ( .A(n7265), .ZN(n7266) );
  OAI21_X1 U8981 ( .B1(n7267), .B2(n7266), .A(n7531), .ZN(n7280) );
  MUX2_X1 U8982 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n7269), .S(n7268), .Z(n8869)
         );
  OAI21_X1 U8983 ( .B1(n7272), .B2(n7271), .A(n7270), .ZN(n8870) );
  NAND2_X1 U8984 ( .A1(n8869), .A2(n8870), .ZN(n8868) );
  OAI21_X1 U8985 ( .B1(n8865), .B2(n7269), .A(n8868), .ZN(n7275) );
  MUX2_X1 U8986 ( .A(n7273), .B(P2_REG1_REG_11__SCAN_IN), .S(n7530), .Z(n7274)
         );
  NAND2_X1 U8987 ( .A1(n7274), .A2(n7275), .ZN(n7522) );
  OAI211_X1 U8988 ( .C1(n7275), .C2(n7274), .A(n10007), .B(n7522), .ZN(n7278)
         );
  AND2_X1 U8989 ( .A1(P2_U3152), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7276) );
  AOI21_X1 U8990 ( .B1(n10013), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n7276), .ZN(
        n7277) );
  OAI211_X1 U8991 ( .C1(n10009), .C2(n7530), .A(n7278), .B(n7277), .ZN(n7279)
         );
  AOI21_X1 U8992 ( .B1(n7280), .B2(n10008), .A(n7279), .ZN(n7281) );
  INV_X1 U8993 ( .A(n7281), .ZN(P2_U3256) );
  INV_X1 U8994 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7294) );
  NAND2_X1 U8995 ( .A1(n7283), .A2(n8569), .ZN(n7284) );
  NAND2_X1 U8996 ( .A1(n7282), .A2(n7284), .ZN(n9935) );
  NAND2_X1 U8997 ( .A1(n8428), .A2(n7285), .ZN(n7286) );
  NAND2_X1 U8998 ( .A1(n7286), .A2(n8569), .ZN(n7436) );
  OAI21_X1 U8999 ( .B1(n8569), .B2(n7286), .A(n7436), .ZN(n7289) );
  OAI22_X1 U9000 ( .A1(n7287), .A2(n5531), .B1(n8431), .B2(n9550), .ZN(n7288)
         );
  AOI21_X1 U9001 ( .B1(n7289), .B2(n9747), .A(n7288), .ZN(n9933) );
  NAND2_X1 U9002 ( .A1(n7360), .A2(n9925), .ZN(n7290) );
  NAND2_X1 U9003 ( .A1(n7290), .A2(n9764), .ZN(n7291) );
  NOR2_X1 U9004 ( .A1(n7443), .A2(n7291), .ZN(n9931) );
  AOI21_X1 U9005 ( .B1(n9670), .B2(n9925), .A(n9931), .ZN(n7292) );
  OAI211_X1 U9006 ( .C1(n9935), .C2(n9672), .A(n9933), .B(n7292), .ZN(n7295)
         );
  NAND2_X1 U9007 ( .A1(n7295), .A2(n9983), .ZN(n7293) );
  OAI21_X1 U9008 ( .B1(n9983), .B2(n7294), .A(n7293), .ZN(P1_U3469) );
  NAND2_X1 U9009 ( .A1(n7295), .A2(n9990), .ZN(n7296) );
  OAI21_X1 U9010 ( .B1(n9990), .B2(n7297), .A(n7296), .ZN(P1_U3528) );
  XNOR2_X1 U9011 ( .A(n7299), .B(n7298), .ZN(n7300) );
  XNOR2_X1 U9012 ( .A(n7301), .B(n7300), .ZN(n7306) );
  NAND2_X1 U9013 ( .A1(n9353), .A2(n9308), .ZN(n7302) );
  NAND2_X1 U9014 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3084), .ZN(n9851) );
  OAI211_X1 U9015 ( .C1(n7589), .C2(n9325), .A(n7302), .B(n9851), .ZN(n7304)
         );
  NOR2_X1 U9016 ( .A1(n9332), .A2(n8436), .ZN(n7303) );
  AOI211_X1 U9017 ( .C1(n7505), .C2(n9329), .A(n7304), .B(n7303), .ZN(n7305)
         );
  OAI21_X1 U9018 ( .B1(n7306), .B2(n9315), .A(n7305), .ZN(P1_U3211) );
  OAI222_X1 U9019 ( .A1(n8661), .A2(n7309), .B1(n7308), .B2(P2_U3152), .C1(
        n8665), .C2(n7307), .ZN(P2_U3342) );
  INV_X1 U9020 ( .A(n7310), .ZN(n7311) );
  AOI21_X1 U9021 ( .B1(n7313), .B2(n7312), .A(n7311), .ZN(n7319) );
  INV_X1 U9022 ( .A(n7314), .ZN(n7755) );
  AOI22_X1 U9023 ( .A1(n9998), .A2(n8860), .B1(n8821), .B2(n8858), .ZN(n7316)
         );
  OAI211_X1 U9024 ( .C1(n10071), .C2(n10000), .A(n7316), .B(n7315), .ZN(n7317)
         );
  AOI21_X1 U9025 ( .B1(n7755), .B2(n8789), .A(n7317), .ZN(n7318) );
  OAI21_X1 U9026 ( .B1(n7319), .B2(n8836), .A(n7318), .ZN(P2_U3232) );
  NAND2_X1 U9027 ( .A1(n7461), .A2(n7320), .ZN(n10048) );
  INV_X1 U9028 ( .A(n10048), .ZN(n7339) );
  INV_X1 U9029 ( .A(n7321), .ZN(n7322) );
  NOR2_X1 U9030 ( .A1(n10035), .A2(n7322), .ZN(n7323) );
  NAND2_X1 U9031 ( .A1(n7324), .A2(n7323), .ZN(n7540) );
  INV_X1 U9032 ( .A(n7540), .ZN(n7325) );
  INV_X1 U9033 ( .A(n7544), .ZN(n7573) );
  NAND3_X1 U9034 ( .A1(n7325), .A2(n7541), .A3(n7573), .ZN(n7466) );
  NAND2_X2 U9035 ( .A1(n7466), .A2(n10025), .ZN(n9079) );
  NOR2_X1 U9036 ( .A1(n10046), .A2(n8974), .ZN(n7329) );
  MUX2_X1 U9037 ( .A(n7327), .B(n7326), .S(n7745), .Z(n7328) );
  NAND2_X1 U9038 ( .A1(n7329), .A2(n7328), .ZN(n8225) );
  NAND2_X1 U9039 ( .A1(n7330), .A2(n7745), .ZN(n7871) );
  NAND2_X1 U9040 ( .A1(n8225), .A2(n7871), .ZN(n10018) );
  AOI22_X1 U9041 ( .A1(n10048), .A2(n9084), .B1(n9068), .B2(n8861), .ZN(n10050) );
  OAI21_X1 U9042 ( .B1(n4615), .B2(n10025), .A(n10050), .ZN(n7335) );
  NOR2_X1 U9043 ( .A1(n9079), .A2(n7333), .ZN(n7334) );
  AOI21_X1 U9044 ( .B1(n7335), .B2(n9079), .A(n7334), .ZN(n7338) );
  AND2_X1 U9045 ( .A1(n10046), .A2(n6200), .ZN(n10021) );
  OR2_X1 U9046 ( .A1(n7466), .A2(n7336), .ZN(n8923) );
  INV_X1 U9047 ( .A(n8923), .ZN(n9074) );
  OAI21_X1 U9048 ( .B1(n9092), .B2(n9074), .A(n10047), .ZN(n7337) );
  OAI211_X1 U9049 ( .C1(n7339), .C2(n9094), .A(n7338), .B(n7337), .ZN(P2_U3296) );
  INV_X1 U9050 ( .A(n7340), .ZN(n7343) );
  OAI222_X1 U9051 ( .A1(n8665), .A2(n7343), .B1(n8880), .B2(P2_U3152), .C1(
        n7341), .C2(n8661), .ZN(P2_U3341) );
  INV_X1 U9052 ( .A(n9914), .ZN(n9366) );
  OAI222_X1 U9053 ( .A1(P1_U3084), .A2(n9366), .B1(n9707), .B2(n7343), .C1(
        n7342), .C2(n9704), .ZN(P1_U3336) );
  NAND2_X1 U9054 ( .A1(n7345), .A2(n7344), .ZN(n8419) );
  INV_X1 U9055 ( .A(n8566), .ZN(n7346) );
  XNOR2_X1 U9056 ( .A(n8419), .B(n7346), .ZN(n7354) );
  OR2_X1 U9057 ( .A1(n7347), .A2(n8566), .ZN(n7348) );
  NAND2_X1 U9058 ( .A1(n7349), .A2(n7348), .ZN(n9965) );
  NAND2_X1 U9059 ( .A1(n9965), .A2(n9758), .ZN(n7353) );
  OAI22_X1 U9060 ( .A1(n7438), .A2(n9550), .B1(n7350), .B2(n5531), .ZN(n7351)
         );
  INV_X1 U9061 ( .A(n7351), .ZN(n7352) );
  OAI211_X1 U9062 ( .C1(n9572), .C2(n7354), .A(n7353), .B(n7352), .ZN(n9963)
         );
  MUX2_X1 U9063 ( .A(n9963), .B(P1_REG2_REG_4__SCAN_IN), .S(n9578), .Z(n7355)
         );
  INV_X1 U9064 ( .A(n7355), .ZN(n7366) );
  AND2_X1 U9065 ( .A1(n7015), .A2(n9497), .ZN(n7356) );
  NAND2_X1 U9066 ( .A1(n7358), .A2(n7357), .ZN(n7359) );
  NAND2_X1 U9067 ( .A1(n7360), .A2(n7359), .ZN(n9962) );
  INV_X1 U9068 ( .A(n9940), .ZN(n9407) );
  OAI22_X1 U9069 ( .A1(n9568), .A2(n9961), .B1(n7361), .B2(n9949), .ZN(n7362)
         );
  INV_X1 U9070 ( .A(n7362), .ZN(n7363) );
  OAI21_X1 U9071 ( .B1(n9962), .B2(n9407), .A(n7363), .ZN(n7364) );
  AOI21_X1 U9072 ( .B1(n9965), .B2(n9768), .A(n7364), .ZN(n7365) );
  NAND2_X1 U9073 ( .A1(n7366), .A2(n7365), .ZN(P1_U3287) );
  INV_X1 U9074 ( .A(n7367), .ZN(n7376) );
  NOR2_X1 U9075 ( .A1(n9949), .A2(n7013), .ZN(n7370) );
  NOR2_X1 U9076 ( .A1(n9568), .A2(n7368), .ZN(n7369) );
  AOI211_X1 U9077 ( .C1(n9578), .C2(P1_REG2_REG_2__SCAN_IN), .A(n7370), .B(
        n7369), .ZN(n7371) );
  OAI21_X1 U9078 ( .B1(n9407), .B2(n7372), .A(n7371), .ZN(n7373) );
  AOI21_X1 U9079 ( .B1(n9768), .B2(n7374), .A(n7373), .ZN(n7375) );
  OAI21_X1 U9080 ( .B1(n7376), .B2(n9578), .A(n7375), .ZN(P1_U3289) );
  NOR2_X1 U9081 ( .A1(n4378), .A2(n7377), .ZN(n7411) );
  AOI21_X1 U9082 ( .B1(n4378), .B2(n7377), .A(n7411), .ZN(n7378) );
  NAND2_X1 U9083 ( .A1(n7378), .A2(n7379), .ZN(n7413) );
  OAI21_X1 U9084 ( .B1(n7379), .B2(n7378), .A(n7413), .ZN(n7380) );
  NAND2_X1 U9085 ( .A1(n7380), .A2(n9322), .ZN(n7385) );
  NAND2_X1 U9086 ( .A1(n9355), .A2(n9308), .ZN(n7381) );
  NAND2_X1 U9087 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3084), .ZN(n9834) );
  OAI211_X1 U9088 ( .C1(n8431), .C2(n9325), .A(n7381), .B(n9834), .ZN(n7382)
         );
  AOI21_X1 U9089 ( .B1(n7383), .B2(n9329), .A(n7382), .ZN(n7384) );
  OAI211_X1 U9090 ( .C1(n7386), .C2(n9332), .A(n7385), .B(n7384), .ZN(P1_U3225) );
  OAI21_X1 U9091 ( .B1(n7389), .B2(n7388), .A(n7387), .ZN(n7390) );
  NAND2_X1 U9092 ( .A1(n7390), .A2(n10002), .ZN(n7394) );
  INV_X1 U9093 ( .A(n8857), .ZN(n7719) );
  OAI22_X1 U9094 ( .A1(n9995), .A2(n7719), .B1(n7555), .B2(n8818), .ZN(n7391)
         );
  AOI211_X1 U9095 ( .C1(n8834), .C2(n10022), .A(n7392), .B(n7391), .ZN(n7393)
         );
  OAI211_X1 U9096 ( .C1(n10006), .C2(n10024), .A(n7394), .B(n7393), .ZN(
        P2_U3229) );
  OAI21_X1 U9097 ( .B1(n7397), .B2(n7396), .A(n7395), .ZN(n7398) );
  INV_X1 U9098 ( .A(n7398), .ZN(n7512) );
  OR2_X1 U9099 ( .A1(n7400), .A2(n8574), .ZN(n7401) );
  NAND2_X1 U9100 ( .A1(n7399), .A2(n7401), .ZN(n7403) );
  OAI22_X1 U9101 ( .A1(n8431), .A2(n5531), .B1(n7589), .B2(n9550), .ZN(n7402)
         );
  AOI21_X1 U9102 ( .B1(n7403), .B2(n9747), .A(n7402), .ZN(n7507) );
  INV_X1 U9103 ( .A(n7445), .ZN(n7405) );
  INV_X1 U9104 ( .A(n7495), .ZN(n7404) );
  AOI211_X1 U9105 ( .C1(n8441), .C2(n7405), .A(n9975), .B(n7404), .ZN(n7510)
         );
  AOI21_X1 U9106 ( .B1(n9670), .B2(n8441), .A(n7510), .ZN(n7406) );
  OAI211_X1 U9107 ( .C1(n7512), .C2(n9672), .A(n7507), .B(n7406), .ZN(n7408)
         );
  NAND2_X1 U9108 ( .A1(n7408), .A2(n9990), .ZN(n7407) );
  OAI21_X1 U9109 ( .B1(n9990), .B2(n6922), .A(n7407), .ZN(P1_U3530) );
  INV_X1 U9110 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7410) );
  NAND2_X1 U9111 ( .A1(n7408), .A2(n9983), .ZN(n7409) );
  OAI21_X1 U9112 ( .B1(n9983), .B2(n7410), .A(n7409), .ZN(P1_U3475) );
  INV_X1 U9113 ( .A(n7411), .ZN(n7412) );
  NAND2_X1 U9114 ( .A1(n7413), .A2(n7412), .ZN(n7417) );
  NAND2_X1 U9115 ( .A1(n7415), .A2(n7414), .ZN(n7416) );
  XNOR2_X1 U9116 ( .A(n7417), .B(n7416), .ZN(n7423) );
  NAND2_X1 U9117 ( .A1(n9354), .A2(n9308), .ZN(n7419) );
  OAI211_X1 U9118 ( .C1(n8438), .C2(n9325), .A(n7419), .B(n7418), .ZN(n7421)
         );
  NOR2_X1 U9119 ( .A1(n9332), .A2(n9967), .ZN(n7420) );
  AOI211_X1 U9120 ( .C1(n7446), .C2(n9329), .A(n7421), .B(n7420), .ZN(n7422)
         );
  OAI21_X1 U9121 ( .B1(n7423), .B2(n9315), .A(n7422), .ZN(P1_U3237) );
  XNOR2_X1 U9122 ( .A(n7426), .B(n7425), .ZN(n7427) );
  XNOR2_X1 U9123 ( .A(n7424), .B(n7427), .ZN(n7432) );
  INV_X1 U9124 ( .A(n8438), .ZN(n9352) );
  NAND2_X1 U9125 ( .A1(n9352), .A2(n9308), .ZN(n7428) );
  NAND2_X1 U9126 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3084), .ZN(n9866) );
  OAI211_X1 U9127 ( .C1(n7691), .C2(n9325), .A(n7428), .B(n9866), .ZN(n7430)
         );
  INV_X1 U9128 ( .A(n7498), .ZN(n9974) );
  NOR2_X1 U9129 ( .A1(n9974), .A2(n9332), .ZN(n7429) );
  AOI211_X1 U9130 ( .C1(n7497), .C2(n9329), .A(n7430), .B(n7429), .ZN(n7431)
         );
  OAI21_X1 U9131 ( .B1(n7432), .B2(n9315), .A(n7431), .ZN(P1_U3219) );
  INV_X1 U9132 ( .A(n7433), .ZN(n7434) );
  AOI21_X1 U9133 ( .B1(n8571), .B2(n7435), .A(n7434), .ZN(n7442) );
  NAND2_X1 U9134 ( .A1(n7436), .A2(n8422), .ZN(n7437) );
  XNOR2_X1 U9135 ( .A(n7437), .B(n8571), .ZN(n7440) );
  OAI22_X1 U9136 ( .A1(n8438), .A2(n9550), .B1(n7438), .B2(n5531), .ZN(n7439)
         );
  AOI21_X1 U9137 ( .B1(n7440), .B2(n9747), .A(n7439), .ZN(n7441) );
  OAI21_X1 U9138 ( .B1(n7442), .B2(n7493), .A(n7441), .ZN(n9969) );
  INV_X1 U9139 ( .A(n9969), .ZN(n7451) );
  INV_X1 U9140 ( .A(n7442), .ZN(n9971) );
  NOR2_X1 U9141 ( .A1(n7443), .A2(n9967), .ZN(n7444) );
  OR2_X1 U9142 ( .A1(n7445), .A2(n7444), .ZN(n9968) );
  AOI22_X1 U9143 ( .A1(n9578), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7446), .B2(
        n9759), .ZN(n7448) );
  NAND2_X1 U9144 ( .A1(n9941), .A2(n8434), .ZN(n7447) );
  OAI211_X1 U9145 ( .C1(n9968), .C2(n9407), .A(n7448), .B(n7447), .ZN(n7449)
         );
  AOI21_X1 U9146 ( .B1(n9971), .B2(n9768), .A(n7449), .ZN(n7450) );
  OAI21_X1 U9147 ( .B1(n7451), .B2(n9578), .A(n7450), .ZN(P1_U3285) );
  NAND2_X1 U9148 ( .A1(n7452), .A2(n9940), .ZN(n7454) );
  AOI22_X1 U9149 ( .A1(n9578), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9759), .B2(
        n5101), .ZN(n7453) );
  OAI211_X1 U9150 ( .C1(n7455), .C2(n9568), .A(n7454), .B(n7453), .ZN(n7456)
         );
  AOI21_X1 U9151 ( .B1(n7457), .B2(n9768), .A(n7456), .ZN(n7458) );
  OAI21_X1 U9152 ( .B1(n7459), .B2(n9578), .A(n7458), .ZN(P1_U3288) );
  INV_X2 U9153 ( .A(n9079), .ZN(n9017) );
  NAND2_X1 U9154 ( .A1(n6204), .A2(n7460), .ZN(n7471) );
  XNOR2_X1 U9155 ( .A(n7471), .B(n7461), .ZN(n7462) );
  NAND2_X1 U9156 ( .A1(n7462), .A2(n9084), .ZN(n7465) );
  INV_X1 U9157 ( .A(n7463), .ZN(n7464) );
  NAND2_X1 U9158 ( .A1(n7465), .A2(n7464), .ZN(n10053) );
  INV_X1 U9159 ( .A(n10053), .ZN(n7474) );
  OAI22_X1 U9160 ( .A1(n7111), .A2(n10025), .B1(n7032), .B2(n9079), .ZN(n7469)
         );
  OR2_X1 U9161 ( .A1(n7466), .A2(n8974), .ZN(n8916) );
  NAND2_X1 U9162 ( .A1(n10047), .A2(n7546), .ZN(n7545) );
  NAND2_X1 U9163 ( .A1(n7467), .A2(n10052), .ZN(n7558) );
  NAND3_X1 U9164 ( .A1(n7545), .A2(n7558), .A3(n9181), .ZN(n10051) );
  NOR2_X1 U9165 ( .A1(n8916), .A2(n10051), .ZN(n7468) );
  AOI211_X1 U9166 ( .C1(n9092), .C2(n7546), .A(n7469), .B(n7468), .ZN(n7473)
         );
  NAND2_X1 U9167 ( .A1(n8863), .A2(n10047), .ZN(n7470) );
  XNOR2_X1 U9168 ( .A(n7471), .B(n7470), .ZN(n10055) );
  NAND2_X1 U9169 ( .A1(n9006), .A2(n10055), .ZN(n7472) );
  OAI211_X1 U9170 ( .C1(n9017), .C2(n7474), .A(n7473), .B(n7472), .ZN(P2_U3295) );
  OAI21_X1 U9171 ( .B1(n7477), .B2(n7476), .A(n7475), .ZN(n7478) );
  NAND2_X1 U9172 ( .A1(n7478), .A2(n10002), .ZN(n7482) );
  OAI22_X1 U9173 ( .A1(n9995), .A2(n7720), .B1(n7634), .B2(n8818), .ZN(n7479)
         );
  AOI211_X1 U9174 ( .C1(n8834), .C2(n7640), .A(n7480), .B(n7479), .ZN(n7481)
         );
  OAI211_X1 U9175 ( .C1(n10006), .C2(n7635), .A(n7482), .B(n7481), .ZN(
        P2_U3241) );
  NAND2_X1 U9176 ( .A1(n7484), .A2(n8575), .ZN(n7485) );
  NAND2_X1 U9177 ( .A1(n7483), .A2(n7485), .ZN(n7494) );
  AOI22_X1 U9178 ( .A1(n9352), .A2(n9754), .B1(n9751), .B2(n9350), .ZN(n7492)
         );
  INV_X1 U9179 ( .A(n7399), .ZN(n7488) );
  OAI21_X1 U9180 ( .B1(n7488), .B2(n7487), .A(n7486), .ZN(n7490) );
  NAND3_X1 U9181 ( .A1(n7490), .A2(n9747), .A3(n7489), .ZN(n7491) );
  OAI211_X1 U9182 ( .C1(n7494), .C2(n7493), .A(n7492), .B(n7491), .ZN(n9977)
         );
  INV_X1 U9183 ( .A(n9977), .ZN(n7503) );
  INV_X1 U9184 ( .A(n7494), .ZN(n9979) );
  NAND2_X1 U9185 ( .A1(n7495), .A2(n7498), .ZN(n7496) );
  NAND2_X1 U9186 ( .A1(n7583), .A2(n7496), .ZN(n9976) );
  AOI22_X1 U9187 ( .A1(n9578), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7497), .B2(
        n9759), .ZN(n7500) );
  NAND2_X1 U9188 ( .A1(n9941), .A2(n7498), .ZN(n7499) );
  OAI211_X1 U9189 ( .C1(n9976), .C2(n9407), .A(n7500), .B(n7499), .ZN(n7501)
         );
  AOI21_X1 U9190 ( .B1(n9979), .B2(n9768), .A(n7501), .ZN(n7502) );
  OAI21_X1 U9191 ( .B1(n7503), .B2(n9578), .A(n7502), .ZN(P1_U3283) );
  NOR2_X1 U9192 ( .A1(n7504), .A2(n9497), .ZN(n9767) );
  OAI22_X1 U9193 ( .A1(n9568), .A2(n8436), .B1(n6931), .B2(n9945), .ZN(n7509)
         );
  NAND2_X1 U9194 ( .A1(n9759), .A2(n7505), .ZN(n7506) );
  AOI21_X1 U9195 ( .B1(n7507), .B2(n7506), .A(n9578), .ZN(n7508) );
  AOI211_X1 U9196 ( .C1(n7510), .C2(n9767), .A(n7509), .B(n7508), .ZN(n7511)
         );
  OAI21_X1 U9197 ( .B1(n7512), .B2(n9582), .A(n7511), .ZN(P1_U3284) );
  XNOR2_X1 U9198 ( .A(n7513), .B(n7514), .ZN(n7521) );
  INV_X1 U9199 ( .A(n7515), .ZN(n7798) );
  OAI22_X1 U9200 ( .A1(n7719), .A2(n8818), .B1(n10000), .B2(n7801), .ZN(n7519)
         );
  OAI22_X1 U9201 ( .A1(n9995), .A2(n7517), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7516), .ZN(n7518) );
  AOI211_X1 U9202 ( .C1(n7798), .C2(n8789), .A(n7519), .B(n7518), .ZN(n7520)
         );
  OAI21_X1 U9203 ( .B1(n7521), .B2(n8836), .A(n7520), .ZN(P2_U3215) );
  OAI21_X1 U9204 ( .B1(n7530), .B2(n7273), .A(n7522), .ZN(n7525) );
  MUX2_X1 U9205 ( .A(n7523), .B(P2_REG1_REG_12__SCAN_IN), .S(n7650), .Z(n7524)
         );
  NOR2_X1 U9206 ( .A1(n7525), .A2(n7524), .ZN(n7644) );
  AOI21_X1 U9207 ( .B1(n7525), .B2(n7524), .A(n7644), .ZN(n7529) );
  NOR2_X1 U9208 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7526), .ZN(n7527) );
  AOI21_X1 U9209 ( .B1(n10013), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n7527), .ZN(
        n7528) );
  OAI21_X1 U9210 ( .B1(n7529), .B2(n10011), .A(n7528), .ZN(n7536) );
  INV_X1 U9211 ( .A(n7530), .ZN(n7532) );
  OAI21_X1 U9212 ( .B1(n7532), .B2(P2_REG2_REG_11__SCAN_IN), .A(n7531), .ZN(
        n7534) );
  MUX2_X1 U9213 ( .A(n8081), .B(P2_REG2_REG_12__SCAN_IN), .S(n7650), .Z(n7533)
         );
  NOR2_X1 U9214 ( .A1(n7533), .A2(n7534), .ZN(n7649) );
  AOI211_X1 U9215 ( .C1(n7534), .C2(n7533), .A(n7649), .B(n9725), .ZN(n7535)
         );
  AOI211_X1 U9216 ( .C1(n9731), .C2(n7650), .A(n7536), .B(n7535), .ZN(n7537)
         );
  INV_X1 U9217 ( .A(n7537), .ZN(P2_U3257) );
  INV_X1 U9218 ( .A(n7538), .ZN(n7539) );
  NOR2_X1 U9219 ( .A1(n7540), .A2(n7539), .ZN(n7543) );
  INV_X1 U9220 ( .A(n7541), .ZN(n7542) );
  INV_X1 U9221 ( .A(n7545), .ZN(n7550) );
  NAND2_X1 U9222 ( .A1(n8861), .A2(n7546), .ZN(n7547) );
  NAND2_X1 U9223 ( .A1(n7548), .A2(n7547), .ZN(n7549) );
  OAI211_X1 U9224 ( .C1(n7550), .C2(n8861), .A(n7549), .B(n7558), .ZN(n8701)
         );
  NAND2_X1 U9225 ( .A1(n8701), .A2(n8700), .ZN(n7552) );
  NAND2_X1 U9226 ( .A1(n7226), .A2(n10058), .ZN(n7551) );
  NAND2_X1 U9227 ( .A1(n7552), .A2(n7551), .ZN(n7674) );
  NAND2_X1 U9228 ( .A1(n7674), .A2(n7675), .ZN(n7554) );
  NAND2_X1 U9229 ( .A1(n8699), .A2(n10062), .ZN(n7553) );
  NAND2_X1 U9230 ( .A1(n7554), .A2(n7553), .ZN(n7746) );
  NAND2_X1 U9231 ( .A1(n7746), .A2(n7747), .ZN(n7557) );
  NAND2_X1 U9232 ( .A1(n7555), .A2(n10071), .ZN(n7556) );
  NAND2_X1 U9233 ( .A1(n7557), .A2(n7556), .ZN(n7628) );
  XNOR2_X1 U9234 ( .A(n7628), .B(n7565), .ZN(n10019) );
  INV_X1 U9235 ( .A(n7558), .ZN(n8704) );
  NOR2_X1 U9236 ( .A1(n7753), .A2(n7756), .ZN(n7561) );
  NAND2_X1 U9237 ( .A1(n7562), .A2(n10071), .ZN(n7559) );
  INV_X1 U9238 ( .A(n7637), .ZN(n7560) );
  OAI211_X1 U9239 ( .C1(n7562), .C2(n7561), .A(n7560), .B(n9181), .ZN(n10020)
         );
  OAI21_X1 U9240 ( .B1(n7562), .B2(n10095), .A(n10020), .ZN(n7571) );
  NAND2_X1 U9241 ( .A1(n7563), .A2(n7564), .ZN(n7567) );
  INV_X1 U9242 ( .A(n7565), .ZN(n7566) );
  XNOR2_X1 U9243 ( .A(n7567), .B(n7566), .ZN(n7568) );
  NAND2_X1 U9244 ( .A1(n7568), .A2(n9084), .ZN(n7570) );
  AOI22_X1 U9245 ( .A1(n9070), .A2(n8859), .B1(n8857), .B2(n9068), .ZN(n7569)
         );
  NAND2_X1 U9246 ( .A1(n7570), .A2(n7569), .ZN(n10032) );
  AOI211_X1 U9247 ( .C1(n10101), .C2(n10019), .A(n7571), .B(n10032), .ZN(n7575) );
  OR2_X1 U9248 ( .A1(n7575), .A2(n10117), .ZN(n7572) );
  OAI21_X1 U9249 ( .B1(n10119), .B2(n7054), .A(n7572), .ZN(P2_U3525) );
  INV_X1 U9250 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7577) );
  OR2_X1 U9251 ( .A1(n7575), .A2(n10103), .ZN(n7576) );
  OAI21_X1 U9252 ( .B1(n10105), .B2(n7577), .A(n7576), .ZN(P2_U3466) );
  INV_X1 U9253 ( .A(n9389), .ZN(n9391) );
  INV_X1 U9254 ( .A(n7578), .ZN(n7580) );
  INV_X1 U9255 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7579) );
  OAI222_X1 U9256 ( .A1(n9391), .A2(P1_U3084), .B1(n9707), .B2(n7580), .C1(
        n7579), .C2(n9704), .ZN(P1_U3335) );
  OAI222_X1 U9257 ( .A1(n8661), .A2(n7581), .B1(n8665), .B2(n7580), .C1(
        P2_U3152), .C2(n8900), .ZN(P2_U3340) );
  XOR2_X1 U9258 ( .A(n7582), .B(n8576), .Z(n7702) );
  AOI21_X1 U9259 ( .B1(n7698), .B2(n7583), .A(n4533), .ZN(n7699) );
  INV_X1 U9260 ( .A(n7698), .ZN(n7585) );
  AOI22_X1 U9261 ( .A1(n9578), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7684), .B2(
        n9759), .ZN(n7584) );
  OAI21_X1 U9262 ( .B1(n7585), .B2(n9568), .A(n7584), .ZN(n7594) );
  INV_X1 U9263 ( .A(n7586), .ZN(n7588) );
  INV_X1 U9264 ( .A(n8576), .ZN(n7587) );
  AOI21_X1 U9265 ( .B1(n7588), .B2(n7587), .A(n9572), .ZN(n7592) );
  OAI22_X1 U9266 ( .A1(n7736), .A2(n9550), .B1(n7589), .B2(n5531), .ZN(n7590)
         );
  AOI21_X1 U9267 ( .B1(n7592), .B2(n7591), .A(n7590), .ZN(n7701) );
  NOR2_X1 U9268 ( .A1(n7701), .A2(n9578), .ZN(n7593) );
  AOI211_X1 U9269 ( .C1(n7699), .C2(n9940), .A(n7594), .B(n7593), .ZN(n7595)
         );
  OAI21_X1 U9270 ( .B1(n7702), .B2(n9582), .A(n7595), .ZN(P1_U3282) );
  OAI21_X1 U9271 ( .B1(n7597), .B2(n8578), .A(n7596), .ZN(n7598) );
  INV_X1 U9272 ( .A(n7598), .ZN(n7709) );
  OAI211_X1 U9273 ( .C1(n7601), .C2(n7600), .A(n7599), .B(n9747), .ZN(n7603)
         );
  AOI22_X1 U9274 ( .A1(n9751), .A2(n9753), .B1(n9350), .B2(n9754), .ZN(n7602)
         );
  NAND2_X1 U9275 ( .A1(n7603), .A2(n7602), .ZN(n7705) );
  AOI211_X1 U9276 ( .C1(n7707), .C2(n7604), .A(n9975), .B(n7737), .ZN(n7706)
         );
  NAND2_X1 U9277 ( .A1(n7706), .A2(n9767), .ZN(n7607) );
  AOI22_X1 U9278 ( .A1(n9578), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7605), .B2(
        n9759), .ZN(n7606) );
  OAI211_X1 U9279 ( .C1(n4531), .C2(n9568), .A(n7607), .B(n7606), .ZN(n7608)
         );
  AOI21_X1 U9280 ( .B1(n9945), .B2(n7705), .A(n7608), .ZN(n7609) );
  OAI21_X1 U9281 ( .B1(n7709), .B2(n9582), .A(n7609), .ZN(P1_U3281) );
  NAND2_X1 U9282 ( .A1(n7613), .A2(n7612), .ZN(n9372) );
  OAI21_X1 U9283 ( .B1(n7613), .B2(n7612), .A(n9372), .ZN(n7624) );
  INV_X1 U9284 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7615) );
  OR2_X1 U9285 ( .A1(n9837), .A2(n9370), .ZN(n7614) );
  NAND2_X1 U9286 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8095) );
  OAI211_X1 U9287 ( .C1(n9922), .C2(n7615), .A(n7614), .B(n8095), .ZN(n7623)
         );
  AOI22_X1 U9288 ( .A1(n7618), .A2(n9360), .B1(P1_REG1_REG_14__SCAN_IN), .B2(
        n9370), .ZN(n7619) );
  NOR2_X1 U9289 ( .A1(n7620), .A2(n7619), .ZN(n9359) );
  AOI21_X1 U9290 ( .B1(n7620), .B2(n7619), .A(n9359), .ZN(n7621) );
  NOR2_X1 U9291 ( .A1(n7621), .A2(n9879), .ZN(n7622) );
  AOI211_X1 U9292 ( .C1(n7624), .C2(n9862), .A(n7623), .B(n7622), .ZN(n7625)
         );
  INV_X1 U9293 ( .A(n7625), .ZN(P1_U3255) );
  NOR2_X1 U9294 ( .A1(n8858), .A2(n10022), .ZN(n7627) );
  NAND2_X1 U9295 ( .A1(n8858), .A2(n10022), .ZN(n7626) );
  OAI21_X1 U9296 ( .B1(n7628), .B2(n7627), .A(n7626), .ZN(n7717) );
  XNOR2_X1 U9297 ( .A(n7717), .B(n6122), .ZN(n10080) );
  INV_X1 U9298 ( .A(n10080), .ZN(n7643) );
  INV_X1 U9299 ( .A(n7629), .ZN(n7630) );
  AOI21_X1 U9300 ( .B1(n7632), .B2(n7631), .A(n7630), .ZN(n7633) );
  OAI222_X1 U9301 ( .A1(n9053), .A2(n7720), .B1(n9051), .B2(n7634), .C1(n9049), 
        .C2(n7633), .ZN(n10078) );
  NAND2_X1 U9302 ( .A1(n10078), .A2(n9079), .ZN(n7642) );
  OAI22_X1 U9303 ( .A1(n9079), .A2(n7636), .B1(n7635), .B2(n10025), .ZN(n7639)
         );
  OAI21_X1 U9304 ( .B1(n7637), .B2(n10076), .A(n7797), .ZN(n10077) );
  NOR2_X1 U9305 ( .A1(n10077), .A2(n8923), .ZN(n7638) );
  AOI211_X1 U9306 ( .C1(n9092), .C2(n7640), .A(n7639), .B(n7638), .ZN(n7641)
         );
  OAI211_X1 U9307 ( .C1(n7643), .C2(n9094), .A(n7642), .B(n7641), .ZN(P2_U3290) );
  AOI21_X1 U9308 ( .B1(n7645), .B2(n7523), .A(n7644), .ZN(n7648) );
  AOI22_X1 U9309 ( .A1(n7783), .A2(n5811), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n7646), .ZN(n7647) );
  NOR2_X1 U9310 ( .A1(n7648), .A2(n7647), .ZN(n7778) );
  AOI21_X1 U9311 ( .B1(n7648), .B2(n7647), .A(n7778), .ZN(n7660) );
  NOR2_X1 U9312 ( .A1(n7783), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7651) );
  AOI21_X1 U9313 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n7783), .A(n7651), .ZN(
        n7652) );
  OAI21_X1 U9314 ( .B1(n7653), .B2(n7652), .A(n7782), .ZN(n7654) );
  NAND2_X1 U9315 ( .A1(n7654), .A2(n10008), .ZN(n7659) );
  INV_X1 U9316 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7656) );
  OAI22_X1 U9317 ( .A1(n9714), .A2(n7656), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7655), .ZN(n7657) );
  AOI21_X1 U9318 ( .B1(n9731), .B2(n7783), .A(n7657), .ZN(n7658) );
  OAI211_X1 U9319 ( .C1(n7660), .C2(n10011), .A(n7659), .B(n7658), .ZN(
        P2_U3258) );
  INV_X1 U9320 ( .A(n7661), .ZN(n7664) );
  OAI222_X1 U9321 ( .A1(n8661), .A2(n7662), .B1(n8665), .B2(n7664), .C1(
        P2_U3152), .C2(n10027), .ZN(P2_U3339) );
  OAI222_X1 U9322 ( .A1(P1_U3084), .A2(n9930), .B1(n9707), .B2(n7664), .C1(
        n7663), .C2(n9704), .ZN(P1_U3334) );
  NAND3_X1 U9323 ( .A1(n7666), .A2(n7667), .A3(n7675), .ZN(n7668) );
  NAND2_X1 U9324 ( .A1(n7665), .A2(n7668), .ZN(n7669) );
  NAND2_X1 U9325 ( .A1(n7669), .A2(n9084), .ZN(n7671) );
  AOI22_X1 U9326 ( .A1(n9070), .A2(n6115), .B1(n8859), .B2(n9068), .ZN(n7670)
         );
  AND2_X1 U9327 ( .A1(n7671), .A2(n7670), .ZN(n10068) );
  OAI21_X1 U9328 ( .B1(n8702), .B2(n10062), .A(n7753), .ZN(n10063) );
  OAI22_X1 U9329 ( .A1(n10063), .A2(n8923), .B1(n10025), .B2(
        P2_REG3_REG_3__SCAN_IN), .ZN(n7673) );
  NOR2_X1 U9330 ( .A1(n9063), .A2(n10062), .ZN(n7672) );
  AOI211_X1 U9331 ( .C1(n9017), .C2(P2_REG2_REG_3__SCAN_IN), .A(n7673), .B(
        n7672), .ZN(n7677) );
  XNOR2_X1 U9332 ( .A(n7674), .B(n7675), .ZN(n10065) );
  NAND2_X1 U9333 ( .A1(n10065), .A2(n9006), .ZN(n7676) );
  OAI211_X1 U9334 ( .C1(n9017), .C2(n10068), .A(n7677), .B(n7676), .ZN(
        P2_U3293) );
  INV_X1 U9335 ( .A(n7678), .ZN(n7679) );
  AOI21_X1 U9336 ( .B1(n7681), .B2(n7680), .A(n7679), .ZN(n7687) );
  NAND2_X1 U9337 ( .A1(n9351), .A2(n9308), .ZN(n7682) );
  NAND2_X1 U9338 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3084), .ZN(n9868) );
  OAI211_X1 U9339 ( .C1(n7736), .C2(n9325), .A(n7682), .B(n9868), .ZN(n7683)
         );
  AOI21_X1 U9340 ( .B1(n7684), .B2(n9329), .A(n7683), .ZN(n7686) );
  NAND2_X1 U9341 ( .A1(n7698), .A2(n9313), .ZN(n7685) );
  OAI211_X1 U9342 ( .C1(n7687), .C2(n9315), .A(n7686), .B(n7685), .ZN(P1_U3229) );
  NAND2_X1 U9343 ( .A1(n7678), .A2(n7688), .ZN(n7763) );
  NAND2_X1 U9344 ( .A1(n7762), .A2(n7764), .ZN(n7689) );
  XNOR2_X1 U9345 ( .A(n7763), .B(n7689), .ZN(n7697) );
  OAI21_X1 U9346 ( .B1(n9326), .B2(n7691), .A(n7690), .ZN(n7692) );
  AOI21_X1 U9347 ( .B1(n9264), .B2(n9753), .A(n7692), .ZN(n7693) );
  OAI21_X1 U9348 ( .B1(n9311), .B2(n7694), .A(n7693), .ZN(n7695) );
  AOI21_X1 U9349 ( .B1(n7707), .B2(n9313), .A(n7695), .ZN(n7696) );
  OAI21_X1 U9350 ( .B1(n7697), .B2(n9315), .A(n7696), .ZN(P1_U3215) );
  INV_X1 U9351 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n7704) );
  AOI22_X1 U9352 ( .A1(n7699), .A2(n9764), .B1(n9670), .B2(n7698), .ZN(n7700)
         );
  OAI211_X1 U9353 ( .C1(n7702), .C2(n9672), .A(n7701), .B(n7700), .ZN(n7712)
         );
  NAND2_X1 U9354 ( .A1(n7712), .A2(n9983), .ZN(n7703) );
  OAI21_X1 U9355 ( .B1(n9983), .B2(n7704), .A(n7703), .ZN(P1_U3481) );
  AOI211_X1 U9356 ( .C1(n9670), .C2(n7707), .A(n7706), .B(n7705), .ZN(n7708)
         );
  OAI21_X1 U9357 ( .B1(n7709), .B2(n9672), .A(n7708), .ZN(n9692) );
  NAND2_X1 U9358 ( .A1(n9692), .A2(n9990), .ZN(n7710) );
  OAI21_X1 U9359 ( .B1(n9990), .B2(n7711), .A(n7710), .ZN(P1_U3533) );
  NAND2_X1 U9360 ( .A1(n7712), .A2(n9990), .ZN(n7713) );
  OAI21_X1 U9361 ( .B1(n9990), .B2(n6926), .A(n7713), .ZN(P1_U3532) );
  OAI21_X1 U9362 ( .B1(n7715), .B2(n6126), .A(n7714), .ZN(n7716) );
  AOI222_X1 U9363 ( .A1(n9084), .A2(n7716), .B1(n8855), .B2(n9068), .C1(n9997), 
        .C2(n9070), .ZN(n10083) );
  INV_X1 U9364 ( .A(n7717), .ZN(n7718) );
  NAND2_X1 U9365 ( .A1(n7718), .A2(n7631), .ZN(n7877) );
  NAND2_X1 U9366 ( .A1(n7719), .A2(n10076), .ZN(n7853) );
  NAND2_X1 U9367 ( .A1(n7877), .A2(n7853), .ZN(n7795) );
  NAND2_X1 U9368 ( .A1(n7795), .A2(n7855), .ZN(n7794) );
  NAND2_X1 U9369 ( .A1(n7720), .A2(n7801), .ZN(n7721) );
  AND2_X1 U9370 ( .A1(n7794), .A2(n7721), .ZN(n7723) );
  NAND2_X1 U9371 ( .A1(n7794), .A2(n7854), .ZN(n7852) );
  OAI21_X1 U9372 ( .B1(n7723), .B2(n7722), .A(n7852), .ZN(n7724) );
  INV_X1 U9373 ( .A(n7724), .ZN(n10086) );
  INV_X1 U9374 ( .A(n7725), .ZN(n7796) );
  OAI211_X1 U9375 ( .C1(n7796), .C2(n10084), .A(n9181), .B(n7866), .ZN(n10082)
         );
  INV_X1 U9376 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7726) );
  OAI22_X1 U9377 ( .A1(n9079), .A2(n7726), .B1(n10005), .B2(n10025), .ZN(n7727) );
  AOI21_X1 U9378 ( .B1(n9092), .B2(n7851), .A(n7727), .ZN(n7728) );
  OAI21_X1 U9379 ( .B1(n10082), .B2(n8916), .A(n7728), .ZN(n7729) );
  AOI21_X1 U9380 ( .B1(n10086), .B2(n9006), .A(n7729), .ZN(n7730) );
  OAI21_X1 U9381 ( .B1(n10083), .B2(n9017), .A(n7730), .ZN(P2_U3288) );
  XOR2_X1 U9382 ( .A(n7731), .B(n8579), .Z(n9788) );
  INV_X1 U9383 ( .A(n9788), .ZN(n7742) );
  OAI211_X1 U9384 ( .C1(n7733), .C2(n8579), .A(n7732), .B(n9747), .ZN(n7735)
         );
  NAND2_X1 U9385 ( .A1(n9348), .A2(n9751), .ZN(n7734) );
  OAI211_X1 U9386 ( .C1(n7736), .C2(n5531), .A(n7735), .B(n7734), .ZN(n9786)
         );
  OAI21_X1 U9387 ( .B1(n7737), .B2(n9783), .A(n9762), .ZN(n9784) );
  AOI22_X1 U9388 ( .A1(n9578), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7774), .B2(
        n9759), .ZN(n7739) );
  NAND2_X1 U9389 ( .A1(n6600), .A2(n9941), .ZN(n7738) );
  OAI211_X1 U9390 ( .C1(n9784), .C2(n9407), .A(n7739), .B(n7738), .ZN(n7740)
         );
  AOI21_X1 U9391 ( .B1(n9786), .B2(n9945), .A(n7740), .ZN(n7741) );
  OAI21_X1 U9392 ( .B1(n7742), .B2(n9582), .A(n7741), .ZN(P1_U3280) );
  INV_X1 U9393 ( .A(n7743), .ZN(n7805) );
  OAI222_X1 U9394 ( .A1(n8665), .A2(n7805), .B1(n7745), .B2(P2_U3152), .C1(
        n7744), .C2(n8661), .ZN(P2_U3338) );
  XNOR2_X1 U9395 ( .A(n7746), .B(n7747), .ZN(n10069) );
  INV_X1 U9396 ( .A(n10069), .ZN(n7761) );
  NAND3_X1 U9397 ( .A1(n7665), .A2(n7748), .A3(n7747), .ZN(n7749) );
  NAND2_X1 U9398 ( .A1(n7563), .A2(n7749), .ZN(n7750) );
  NAND2_X1 U9399 ( .A1(n7750), .A2(n9084), .ZN(n7752) );
  AOI22_X1 U9400 ( .A1(n9070), .A2(n8860), .B1(n8858), .B2(n9068), .ZN(n7751)
         );
  NAND2_X1 U9401 ( .A1(n7752), .A2(n7751), .ZN(n10074) );
  XNOR2_X1 U9402 ( .A(n7753), .B(n10071), .ZN(n7754) );
  NAND2_X1 U9403 ( .A1(n7754), .A2(n9181), .ZN(n10070) );
  INV_X1 U9404 ( .A(n10025), .ZN(n9060) );
  AOI22_X1 U9405 ( .A1(n9017), .A2(P2_REG2_REG_4__SCAN_IN), .B1(n7755), .B2(
        n9060), .ZN(n7758) );
  NAND2_X1 U9406 ( .A1(n9092), .A2(n7756), .ZN(n7757) );
  OAI211_X1 U9407 ( .C1(n10070), .C2(n8916), .A(n7758), .B(n7757), .ZN(n7759)
         );
  AOI21_X1 U9408 ( .B1(n10074), .B2(n9079), .A(n7759), .ZN(n7760) );
  OAI21_X1 U9409 ( .B1(n7761), .B2(n9094), .A(n7760), .ZN(P2_U3292) );
  NAND2_X1 U9410 ( .A1(n7763), .A2(n7762), .ZN(n7765) );
  NAND2_X1 U9411 ( .A1(n7765), .A2(n7764), .ZN(n7767) );
  AOI21_X1 U9412 ( .B1(n7767), .B2(n7766), .A(n9315), .ZN(n7769) );
  NAND2_X1 U9413 ( .A1(n7769), .A2(n7768), .ZN(n7776) );
  NAND2_X1 U9414 ( .A1(n9349), .A2(n9308), .ZN(n7771) );
  OAI211_X1 U9415 ( .C1(n7772), .C2(n9325), .A(n7771), .B(n7770), .ZN(n7773)
         );
  AOI21_X1 U9416 ( .B1(n7774), .B2(n9329), .A(n7773), .ZN(n7775) );
  OAI211_X1 U9417 ( .C1(n9783), .C2(n9332), .A(n7776), .B(n7775), .ZN(P1_U3234) );
  NOR2_X1 U9418 ( .A1(n7783), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7777) );
  NOR2_X1 U9419 ( .A1(n7778), .A2(n7777), .ZN(n7781) );
  MUX2_X1 U9420 ( .A(n7779), .B(P2_REG1_REG_14__SCAN_IN), .S(n7940), .Z(n7780)
         );
  NOR2_X1 U9421 ( .A1(n7781), .A2(n7780), .ZN(n7942) );
  AOI21_X1 U9422 ( .B1(n7781), .B2(n7780), .A(n7942), .ZN(n7791) );
  NOR2_X1 U9423 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n7940), .ZN(n7784) );
  AOI21_X1 U9424 ( .B1(n7940), .B2(P2_REG2_REG_14__SCAN_IN), .A(n7784), .ZN(
        n7785) );
  OAI21_X1 U9425 ( .B1(n7786), .B2(n7785), .A(n7939), .ZN(n7787) );
  NAND2_X1 U9426 ( .A1(n7787), .A2(n10008), .ZN(n7790) );
  AND2_X1 U9427 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8259) );
  NOR2_X1 U9428 ( .A1(n10009), .A2(n7943), .ZN(n7788) );
  AOI211_X1 U9429 ( .C1(n10013), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n8259), .B(
        n7788), .ZN(n7789) );
  OAI211_X1 U9430 ( .C1(n7791), .C2(n10011), .A(n7790), .B(n7789), .ZN(
        P2_U3259) );
  XNOR2_X1 U9431 ( .A(n7792), .B(n4619), .ZN(n7793) );
  AOI222_X1 U9432 ( .A1(n8857), .A2(n9070), .B1(n8856), .B2(n9068), .C1(n9084), 
        .C2(n7793), .ZN(n7825) );
  OAI21_X1 U9433 ( .B1(n7795), .B2(n7855), .A(n7794), .ZN(n7821) );
  AOI21_X1 U9434 ( .B1(n7822), .B2(n7797), .A(n7796), .ZN(n7823) );
  NAND2_X1 U9435 ( .A1(n7823), .A2(n9074), .ZN(n7800) );
  AOI22_X1 U9436 ( .A1(n9017), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n7798), .B2(
        n9060), .ZN(n7799) );
  OAI211_X1 U9437 ( .C1(n7801), .C2(n9063), .A(n7800), .B(n7799), .ZN(n7802)
         );
  AOI21_X1 U9438 ( .B1(n7821), .B2(n9006), .A(n7802), .ZN(n7803) );
  OAI21_X1 U9439 ( .B1(n7825), .B2(n9017), .A(n7803), .ZN(P2_U3289) );
  OAI222_X1 U9440 ( .A1(n7806), .A2(P1_U3084), .B1(n9707), .B2(n7805), .C1(
        n7804), .C2(n9704), .ZN(P1_U3333) );
  XNOR2_X1 U9441 ( .A(n7809), .B(n7808), .ZN(n7810) );
  XNOR2_X1 U9442 ( .A(n7807), .B(n7810), .ZN(n7817) );
  NAND2_X1 U9443 ( .A1(n9308), .A2(n9753), .ZN(n7812) );
  OAI211_X1 U9444 ( .C1(n9325), .C2(n7813), .A(n7812), .B(n7811), .ZN(n7815)
         );
  NOR2_X1 U9445 ( .A1(n4532), .A2(n9332), .ZN(n7814) );
  AOI211_X1 U9446 ( .C1(n9760), .C2(n9329), .A(n7815), .B(n7814), .ZN(n7816)
         );
  OAI21_X1 U9447 ( .B1(n7817), .B2(n9315), .A(n7816), .ZN(P1_U3222) );
  INV_X1 U9448 ( .A(n7818), .ZN(n7844) );
  OAI222_X1 U9449 ( .A1(n8665), .A2(n7844), .B1(n7820), .B2(P2_U3152), .C1(
        n7819), .C2(n8661), .ZN(P2_U3337) );
  INV_X1 U9450 ( .A(n7821), .ZN(n7826) );
  AOI22_X1 U9451 ( .A1(n7823), .A2(n9181), .B1(n9180), .B2(n7822), .ZN(n7824)
         );
  OAI211_X1 U9452 ( .C1(n9170), .C2(n7826), .A(n7825), .B(n7824), .ZN(n7829)
         );
  NAND2_X1 U9453 ( .A1(n7829), .A2(n10119), .ZN(n7827) );
  OAI21_X1 U9454 ( .B1(n10119), .B2(n7828), .A(n7827), .ZN(P2_U3527) );
  NAND2_X1 U9455 ( .A1(n7829), .A2(n10105), .ZN(n7830) );
  OAI21_X1 U9456 ( .B1(n10105), .B2(n5696), .A(n7830), .ZN(P2_U3472) );
  INV_X1 U9457 ( .A(n7831), .ZN(n7833) );
  NOR2_X1 U9458 ( .A1(n7833), .A2(n7832), .ZN(n7834) );
  XNOR2_X1 U9459 ( .A(n7835), .B(n7834), .ZN(n7842) );
  NAND2_X1 U9460 ( .A1(n9348), .A2(n9308), .ZN(n7837) );
  OAI211_X1 U9461 ( .C1(n7838), .C2(n9325), .A(n7837), .B(n7836), .ZN(n7840)
         );
  NOR2_X1 U9462 ( .A1(n4535), .A2(n9332), .ZN(n7839) );
  AOI211_X1 U9463 ( .C1(n7903), .C2(n9329), .A(n7840), .B(n7839), .ZN(n7841)
         );
  OAI21_X1 U9464 ( .B1(n7842), .B2(n9315), .A(n7841), .ZN(P1_U3232) );
  OAI222_X1 U9465 ( .A1(n8602), .A2(P1_U3084), .B1(n9707), .B2(n7844), .C1(
        n7843), .C2(n9704), .ZN(P1_U3332) );
  INV_X1 U9466 ( .A(n7845), .ZN(n7848) );
  OAI222_X1 U9467 ( .A1(P1_U3084), .A2(n8555), .B1(n9699), .B2(n7848), .C1(
        n7846), .C2(n9704), .ZN(P1_U3331) );
  OAI222_X1 U9468 ( .A1(n8661), .A2(n7849), .B1(n8665), .B2(n7848), .C1(
        P2_U3152), .C2(n7847), .ZN(P2_U3336) );
  INV_X1 U9469 ( .A(n7857), .ZN(n7862) );
  XNOR2_X1 U9470 ( .A(n7850), .B(n7862), .ZN(n7865) );
  NAND2_X1 U9471 ( .A1(n8856), .A2(n7851), .ZN(n7856) );
  NAND2_X1 U9472 ( .A1(n7852), .A2(n7856), .ZN(n7861) );
  AND2_X1 U9473 ( .A1(n7853), .A2(n7854), .ZN(n7875) );
  NAND2_X1 U9474 ( .A1(n7877), .A2(n7875), .ZN(n7859) );
  AND2_X1 U9475 ( .A1(n7857), .A2(n7856), .ZN(n7858) );
  AND2_X1 U9476 ( .A1(n7859), .A2(n7879), .ZN(n7860) );
  AOI21_X1 U9477 ( .B1(n7862), .B2(n7861), .A(n7860), .ZN(n7961) );
  AOI22_X1 U9478 ( .A1(n9070), .A2(n8856), .B1(n8854), .B2(n9068), .ZN(n7863)
         );
  OAI21_X1 U9479 ( .B1(n7961), .B2(n8225), .A(n7863), .ZN(n7864) );
  AOI21_X1 U9480 ( .B1(n7865), .B2(n9084), .A(n7864), .ZN(n7960) );
  AOI21_X1 U9481 ( .B1(n7957), .B2(n7866), .A(n7889), .ZN(n7958) );
  INV_X1 U9482 ( .A(n7957), .ZN(n7870) );
  INV_X1 U9483 ( .A(n7867), .ZN(n7868) );
  AOI22_X1 U9484 ( .A1(n9017), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7868), .B2(
        n9060), .ZN(n7869) );
  OAI21_X1 U9485 ( .B1(n7870), .B2(n9063), .A(n7869), .ZN(n7873) );
  NOR2_X1 U9486 ( .A1(n9017), .A2(n7871), .ZN(n8238) );
  INV_X1 U9487 ( .A(n8238), .ZN(n7895) );
  NOR2_X1 U9488 ( .A1(n7961), .A2(n7895), .ZN(n7872) );
  AOI211_X1 U9489 ( .C1(n7958), .C2(n9074), .A(n7873), .B(n7872), .ZN(n7874)
         );
  OAI21_X1 U9490 ( .B1(n9017), .B2(n7960), .A(n7874), .ZN(P2_U3287) );
  OR2_X1 U9491 ( .A1(n8855), .A2(n7957), .ZN(n7878) );
  AND2_X1 U9492 ( .A1(n7875), .A2(n7878), .ZN(n7876) );
  NAND2_X1 U9493 ( .A1(n7877), .A2(n7876), .ZN(n7880) );
  NAND2_X1 U9494 ( .A1(n7880), .A2(n4868), .ZN(n7881) );
  NAND2_X1 U9495 ( .A1(n7881), .A2(n7883), .ZN(n7988) );
  OAI21_X1 U9496 ( .B1(n7881), .B2(n7883), .A(n7988), .ZN(n10088) );
  XNOR2_X1 U9497 ( .A(n8009), .B(n7883), .ZN(n7885) );
  OAI22_X1 U9498 ( .A1(n8075), .A2(n9053), .B1(n9994), .B2(n9051), .ZN(n7884)
         );
  AOI21_X1 U9499 ( .B1(n7885), .B2(n9084), .A(n7884), .ZN(n7886) );
  OAI21_X1 U9500 ( .B1(n10088), .B2(n8225), .A(n7886), .ZN(n10091) );
  NAND2_X1 U9501 ( .A1(n10091), .A2(n9079), .ZN(n7894) );
  INV_X1 U9502 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7888) );
  OAI22_X1 U9503 ( .A1(n9079), .A2(n7888), .B1(n7887), .B2(n10025), .ZN(n7892)
         );
  INV_X1 U9504 ( .A(n7986), .ZN(n10089) );
  OR2_X1 U9505 ( .A1(n7889), .A2(n10089), .ZN(n7890) );
  NAND2_X1 U9506 ( .A1(n8018), .A2(n7890), .ZN(n10090) );
  NOR2_X1 U9507 ( .A1(n10090), .A2(n8923), .ZN(n7891) );
  AOI211_X1 U9508 ( .C1(n9092), .C2(n7986), .A(n7892), .B(n7891), .ZN(n7893)
         );
  OAI211_X1 U9509 ( .C1(n10088), .C2(n7895), .A(n7894), .B(n7893), .ZN(
        P2_U3286) );
  XNOR2_X1 U9510 ( .A(n7896), .B(n8581), .ZN(n9773) );
  OAI211_X1 U9511 ( .C1(n7898), .C2(n8581), .A(n7897), .B(n9747), .ZN(n7900)
         );
  AOI22_X1 U9512 ( .A1(n9348), .A2(n9754), .B1(n9751), .B2(n9347), .ZN(n7899)
         );
  NAND2_X1 U9513 ( .A1(n7900), .A2(n7899), .ZN(n7901) );
  AOI21_X1 U9514 ( .B1(n9773), .B2(n9758), .A(n7901), .ZN(n9775) );
  AND2_X1 U9515 ( .A1(n9763), .A2(n7904), .ZN(n7902) );
  OR2_X1 U9516 ( .A1(n7902), .A2(n7973), .ZN(n9771) );
  AOI22_X1 U9517 ( .A1(n9578), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7903), .B2(
        n9759), .ZN(n7906) );
  NAND2_X1 U9518 ( .A1(n7904), .A2(n9941), .ZN(n7905) );
  OAI211_X1 U9519 ( .C1(n9771), .C2(n9407), .A(n7906), .B(n7905), .ZN(n7907)
         );
  AOI21_X1 U9520 ( .B1(n9773), .B2(n9768), .A(n7907), .ZN(n7908) );
  OAI21_X1 U9521 ( .B1(n9775), .B2(n9578), .A(n7908), .ZN(P1_U3278) );
  INV_X1 U9522 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10156) );
  NOR2_X1 U9523 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7909) );
  AOI21_X1 U9524 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7909), .ZN(n10127) );
  NOR2_X1 U9525 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7910) );
  AOI21_X1 U9526 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7910), .ZN(n10130) );
  NOR2_X1 U9527 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7911) );
  AOI21_X1 U9528 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7911), .ZN(n10133) );
  NOR2_X1 U9529 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7912) );
  AOI21_X1 U9530 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7912), .ZN(n10136) );
  NOR2_X1 U9531 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7913) );
  AOI21_X1 U9532 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7913), .ZN(n10139) );
  NOR2_X1 U9533 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7919) );
  XNOR2_X1 U9534 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10167) );
  NAND2_X1 U9535 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7917) );
  XOR2_X1 U9536 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10165) );
  NAND2_X1 U9537 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7915) );
  XOR2_X1 U9538 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10163) );
  AOI21_X1 U9539 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10120) );
  INV_X1 U9540 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10124) );
  NAND3_X1 U9541 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10122) );
  OAI21_X1 U9542 ( .B1(n10120), .B2(n10124), .A(n10122), .ZN(n10162) );
  NAND2_X1 U9543 ( .A1(n10163), .A2(n10162), .ZN(n7914) );
  NAND2_X1 U9544 ( .A1(n7915), .A2(n7914), .ZN(n10164) );
  NAND2_X1 U9545 ( .A1(n10165), .A2(n10164), .ZN(n7916) );
  NAND2_X1 U9546 ( .A1(n7917), .A2(n7916), .ZN(n10166) );
  NOR2_X1 U9547 ( .A1(n10167), .A2(n10166), .ZN(n7918) );
  NOR2_X1 U9548 ( .A1(n7919), .A2(n7918), .ZN(n7920) );
  NOR2_X1 U9549 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7920), .ZN(n10151) );
  AND2_X1 U9550 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7920), .ZN(n10150) );
  NOR2_X1 U9551 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10150), .ZN(n7921) );
  NOR2_X1 U9552 ( .A1(n10151), .A2(n7921), .ZN(n7922) );
  NAND2_X1 U9553 ( .A1(n7922), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7924) );
  XOR2_X1 U9554 ( .A(n7922), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10153) );
  NAND2_X1 U9555 ( .A1(n10153), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7923) );
  NAND2_X1 U9556 ( .A1(n7924), .A2(n7923), .ZN(n7925) );
  NAND2_X1 U9557 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7925), .ZN(n7927) );
  XOR2_X1 U9558 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7925), .Z(n10149) );
  NAND2_X1 U9559 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10149), .ZN(n7926) );
  NAND2_X1 U9560 ( .A1(n7927), .A2(n7926), .ZN(n7928) );
  NAND2_X1 U9561 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7928), .ZN(n7930) );
  XOR2_X1 U9562 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7928), .Z(n10158) );
  NAND2_X1 U9563 ( .A1(n10158), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n7929) );
  NAND2_X1 U9564 ( .A1(n7930), .A2(n7929), .ZN(n7931) );
  AND2_X1 U9565 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7931), .ZN(n7932) );
  INV_X1 U9566 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10161) );
  XNOR2_X1 U9567 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n7931), .ZN(n10160) );
  NAND2_X1 U9568 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7933) );
  OAI21_X1 U9569 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7933), .ZN(n10147) );
  NAND2_X1 U9570 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7934) );
  OAI21_X1 U9571 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7934), .ZN(n10144) );
  AOI21_X1 U9572 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10143), .ZN(n10142) );
  NOR2_X1 U9573 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7935) );
  AOI21_X1 U9574 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7935), .ZN(n10141) );
  NAND2_X1 U9575 ( .A1(n10142), .A2(n10141), .ZN(n10140) );
  OAI21_X1 U9576 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10140), .ZN(n10138) );
  NAND2_X1 U9577 ( .A1(n10139), .A2(n10138), .ZN(n10137) );
  OAI21_X1 U9578 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10137), .ZN(n10135) );
  NAND2_X1 U9579 ( .A1(n10136), .A2(n10135), .ZN(n10134) );
  OAI21_X1 U9580 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10134), .ZN(n10132) );
  NAND2_X1 U9581 ( .A1(n10133), .A2(n10132), .ZN(n10131) );
  OAI21_X1 U9582 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10131), .ZN(n10129) );
  NAND2_X1 U9583 ( .A1(n10130), .A2(n10129), .ZN(n10128) );
  OAI21_X1 U9584 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10128), .ZN(n10126) );
  NAND2_X1 U9585 ( .A1(n10127), .A2(n10126), .ZN(n10125) );
  OAI21_X1 U9586 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10125), .ZN(n10155) );
  NOR2_X1 U9587 ( .A1(n10156), .A2(n10155), .ZN(n7936) );
  NAND2_X1 U9588 ( .A1(n10156), .A2(n10155), .ZN(n10154) );
  OAI21_X1 U9589 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7936), .A(n10154), .ZN(
        n7938) );
  XNOR2_X1 U9590 ( .A(n8910), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n7937) );
  XNOR2_X1 U9591 ( .A(n7938), .B(n7937), .ZN(ADD_1071_U4) );
  OAI21_X1 U9592 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n7940), .A(n7939), .ZN(
        n8188) );
  XNOR2_X1 U9593 ( .A(n8183), .B(n8188), .ZN(n7941) );
  NAND2_X1 U9594 ( .A1(n7941), .A2(n8164), .ZN(n8190) );
  OAI21_X1 U9595 ( .B1(n7941), .B2(n8164), .A(n8190), .ZN(n7949) );
  AOI21_X1 U9596 ( .B1(n7779), .B2(n7943), .A(n7942), .ZN(n8182) );
  XNOR2_X1 U9597 ( .A(n8189), .B(n8182), .ZN(n7944) );
  NAND2_X1 U9598 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n7944), .ZN(n8184) );
  OAI211_X1 U9599 ( .C1(P2_REG1_REG_15__SCAN_IN), .C2(n7944), .A(n10007), .B(
        n8184), .ZN(n7947) );
  NOR2_X1 U9600 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8827), .ZN(n7945) );
  AOI21_X1 U9601 ( .B1(n10013), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7945), .ZN(
        n7946) );
  OAI211_X1 U9602 ( .C1(n10009), .C2(n8189), .A(n7947), .B(n7946), .ZN(n7948)
         );
  AOI21_X1 U9603 ( .B1(n10008), .B2(n7949), .A(n7948), .ZN(n7950) );
  INV_X1 U9604 ( .A(n7950), .ZN(P2_U3260) );
  INV_X1 U9605 ( .A(n7951), .ZN(n7956) );
  AOI21_X1 U9606 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n9210), .A(n7952), .ZN(
        n7953) );
  OAI21_X1 U9607 ( .B1(n7956), .B2(n9212), .A(n7953), .ZN(P2_U3335) );
  OR2_X1 U9608 ( .A1(n7954), .A2(P1_U3084), .ZN(n8655) );
  NAND2_X1 U9609 ( .A1(n9697), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7955) );
  OAI211_X1 U9610 ( .C1(n7956), .C2(n9699), .A(n8655), .B(n7955), .ZN(P1_U3330) );
  AOI22_X1 U9611 ( .A1(n7958), .A2(n9181), .B1(n9180), .B2(n7957), .ZN(n7959)
         );
  OAI211_X1 U9612 ( .C1(n7961), .C2(n10087), .A(n7960), .B(n7959), .ZN(n7963)
         );
  NAND2_X1 U9613 ( .A1(n7963), .A2(n10119), .ZN(n7962) );
  OAI21_X1 U9614 ( .B1(n10119), .B2(n7271), .A(n7962), .ZN(P2_U3529) );
  INV_X1 U9615 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7965) );
  NAND2_X1 U9616 ( .A1(n7963), .A2(n10105), .ZN(n7964) );
  OAI21_X1 U9617 ( .B1(n10105), .B2(n7965), .A(n7964), .ZN(P2_U3478) );
  NAND2_X1 U9618 ( .A1(n7967), .A2(n7966), .ZN(n7968) );
  XOR2_X1 U9619 ( .A(n8583), .B(n7968), .Z(n9673) );
  OAI211_X1 U9620 ( .C1(n7970), .C2(n8583), .A(n7969), .B(n9747), .ZN(n7972)
         );
  AOI22_X1 U9621 ( .A1(n9754), .A2(n9752), .B1(n9346), .B2(n9751), .ZN(n7971)
         );
  NAND2_X1 U9622 ( .A1(n7972), .A2(n7971), .ZN(n9667) );
  INV_X1 U9623 ( .A(n7973), .ZN(n7975) );
  INV_X1 U9624 ( .A(n8116), .ZN(n7974) );
  AOI211_X1 U9625 ( .C1(n9669), .C2(n7975), .A(n9975), .B(n7974), .ZN(n9668)
         );
  NAND2_X1 U9626 ( .A1(n9668), .A2(n9767), .ZN(n7977) );
  AOI22_X1 U9627 ( .A1(n9578), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8098), .B2(
        n9759), .ZN(n7976) );
  OAI211_X1 U9628 ( .C1(n8101), .C2(n9568), .A(n7977), .B(n7976), .ZN(n7978)
         );
  AOI21_X1 U9629 ( .B1(n9945), .B2(n9667), .A(n7978), .ZN(n7979) );
  OAI21_X1 U9630 ( .B1(n9673), .B2(n9582), .A(n7979), .ZN(P1_U3277) );
  AND2_X1 U9631 ( .A1(n7981), .A2(n7980), .ZN(n7983) );
  AND2_X1 U9632 ( .A1(n7983), .A2(n7982), .ZN(n7984) );
  XNOR2_X1 U9633 ( .A(n7984), .B(n7991), .ZN(n7996) );
  OAI22_X1 U9634 ( .A1(n8155), .A2(n9053), .B1(n7985), .B2(n9051), .ZN(n7995)
         );
  NAND2_X1 U9635 ( .A1(n7986), .A2(n8854), .ZN(n7987) );
  NAND2_X1 U9636 ( .A1(n7988), .A2(n7987), .ZN(n8007) );
  NAND2_X1 U9637 ( .A1(n8007), .A2(n8011), .ZN(n7990) );
  NAND2_X1 U9638 ( .A1(n8040), .A2(n8853), .ZN(n7989) );
  NAND2_X1 U9639 ( .A1(n7990), .A2(n7989), .ZN(n8068) );
  NAND2_X1 U9640 ( .A1(n7992), .A2(n7991), .ZN(n7993) );
  NAND2_X1 U9641 ( .A1(n8056), .A2(n7993), .ZN(n9185) );
  NOR2_X1 U9642 ( .A1(n9185), .A2(n8225), .ZN(n7994) );
  AOI211_X1 U9643 ( .C1(n7996), .C2(n9084), .A(n7995), .B(n7994), .ZN(n9184)
         );
  INV_X1 U9644 ( .A(n9179), .ZN(n7997) );
  AOI21_X1 U9645 ( .B1(n9179), .B2(n4379), .A(n8061), .ZN(n9182) );
  NOR2_X1 U9646 ( .A1(n7997), .A2(n9063), .ZN(n8000) );
  OAI22_X1 U9647 ( .A1(n9079), .A2(n7998), .B1(n8149), .B2(n10025), .ZN(n7999)
         );
  AOI211_X1 U9648 ( .C1(n9182), .C2(n9074), .A(n8000), .B(n7999), .ZN(n8003)
         );
  INV_X1 U9649 ( .A(n9185), .ZN(n8001) );
  NAND2_X1 U9650 ( .A1(n8001), .A2(n8238), .ZN(n8002) );
  OAI211_X1 U9651 ( .C1(n9184), .C2(n9017), .A(n8003), .B(n8002), .ZN(P2_U3283) );
  INV_X1 U9652 ( .A(n8004), .ZN(n8033) );
  OAI222_X1 U9653 ( .A1(n8665), .A2(n8033), .B1(P2_U3152), .B2(n8006), .C1(
        n8005), .C2(n8661), .ZN(P2_U3334) );
  XNOR2_X1 U9654 ( .A(n8007), .B(n8011), .ZN(n8027) );
  NAND2_X1 U9655 ( .A1(n8009), .A2(n8008), .ZN(n8070) );
  NAND2_X1 U9656 ( .A1(n8070), .A2(n8010), .ZN(n8012) );
  XNOR2_X1 U9657 ( .A(n8012), .B(n8011), .ZN(n8015) );
  NAND2_X1 U9658 ( .A1(n8854), .A2(n9070), .ZN(n8014) );
  NAND2_X1 U9659 ( .A1(n8852), .A2(n9068), .ZN(n8013) );
  NAND2_X1 U9660 ( .A1(n8014), .A2(n8013), .ZN(n8039) );
  AOI21_X1 U9661 ( .B1(n8015), .B2(n9084), .A(n8039), .ZN(n8026) );
  OAI22_X1 U9662 ( .A1(n9079), .A2(n8016), .B1(n8043), .B2(n10025), .ZN(n8017)
         );
  AOI21_X1 U9663 ( .B1(n9092), .B2(n8040), .A(n8017), .ZN(n8021) );
  AOI21_X1 U9664 ( .B1(n8018), .B2(n8040), .A(n10097), .ZN(n8019) );
  AND2_X1 U9665 ( .A1(n8019), .A2(n8078), .ZN(n8024) );
  NAND2_X1 U9666 ( .A1(n8024), .A2(n9043), .ZN(n8020) );
  OAI211_X1 U9667 ( .C1(n8026), .C2(n9017), .A(n8021), .B(n8020), .ZN(n8022)
         );
  INV_X1 U9668 ( .A(n8022), .ZN(n8023) );
  OAI21_X1 U9669 ( .B1(n9094), .B2(n8027), .A(n8023), .ZN(P2_U3285) );
  AOI21_X1 U9670 ( .B1(n9180), .B2(n8040), .A(n8024), .ZN(n8025) );
  OAI211_X1 U9671 ( .C1(n8027), .C2(n9170), .A(n8026), .B(n8025), .ZN(n8030)
         );
  NAND2_X1 U9672 ( .A1(n8030), .A2(n10105), .ZN(n8028) );
  OAI21_X1 U9673 ( .B1(n10105), .B2(n8029), .A(n8028), .ZN(P2_U3484) );
  NAND2_X1 U9674 ( .A1(n8030), .A2(n10119), .ZN(n8031) );
  OAI21_X1 U9675 ( .B1(n10119), .B2(n7273), .A(n8031), .ZN(P2_U3531) );
  OAI222_X1 U9676 ( .A1(n8034), .A2(P1_U3084), .B1(n9707), .B2(n8033), .C1(
        n8032), .C2(n9704), .ZN(P1_U3329) );
  NAND2_X1 U9677 ( .A1(n8036), .A2(n8035), .ZN(n8037) );
  XOR2_X1 U9678 ( .A(n8038), .B(n8037), .Z(n8045) );
  AOI22_X1 U9679 ( .A1(n8734), .A2(n8039), .B1(P2_REG3_REG_11__SCAN_IN), .B2(
        P2_U3152), .ZN(n8042) );
  NAND2_X1 U9680 ( .A1(n8834), .A2(n8040), .ZN(n8041) );
  OAI211_X1 U9681 ( .C1(n10006), .C2(n8043), .A(n8042), .B(n8041), .ZN(n8044)
         );
  AOI21_X1 U9682 ( .B1(n8045), .B2(n10002), .A(n8044), .ZN(n8046) );
  INV_X1 U9683 ( .A(n8046), .ZN(P2_U3238) );
  XOR2_X1 U9684 ( .A(n8047), .B(n8048), .Z(n8054) );
  AOI22_X1 U9685 ( .A1(n8821), .A2(n8851), .B1(P2_REG3_REG_12__SCAN_IN), .B2(
        P2_U3152), .ZN(n8052) );
  NAND2_X1 U9686 ( .A1(n8083), .A2(n8834), .ZN(n8051) );
  OR2_X1 U9687 ( .A1(n10006), .A2(n8080), .ZN(n8050) );
  OR2_X1 U9688 ( .A1(n8818), .A2(n8075), .ZN(n8049) );
  NAND4_X1 U9689 ( .A1(n8052), .A2(n8051), .A3(n8050), .A4(n8049), .ZN(n8053)
         );
  AOI21_X1 U9690 ( .B1(n8054), .B2(n10002), .A(n8053), .ZN(n8055) );
  INV_X1 U9691 ( .A(n8055), .ZN(P2_U3226) );
  XNOR2_X1 U9692 ( .A(n8157), .B(n6135), .ZN(n9742) );
  INV_X1 U9693 ( .A(n9742), .ZN(n8067) );
  INV_X1 U9694 ( .A(n8057), .ZN(n8058) );
  AOI211_X1 U9695 ( .C1(n8156), .C2(n8059), .A(n9049), .B(n8058), .ZN(n8060)
         );
  OAI22_X1 U9696 ( .A1(n8228), .A2(n9053), .B1(n8077), .B2(n9051), .ZN(n8260)
         );
  OR2_X1 U9697 ( .A1(n8060), .A2(n8260), .ZN(n9740) );
  INV_X1 U9698 ( .A(n8264), .ZN(n9738) );
  NAND2_X1 U9699 ( .A1(n8061), .A2(n9738), .ZN(n8162) );
  OAI21_X1 U9700 ( .B1(n8061), .B2(n9738), .A(n8162), .ZN(n9739) );
  INV_X1 U9701 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8062) );
  OAI22_X1 U9702 ( .A1(n9079), .A2(n8062), .B1(n8262), .B2(n10025), .ZN(n8063)
         );
  AOI21_X1 U9703 ( .B1(n8264), .B2(n9092), .A(n8063), .ZN(n8064) );
  OAI21_X1 U9704 ( .B1(n9739), .B2(n8923), .A(n8064), .ZN(n8065) );
  AOI21_X1 U9705 ( .B1(n9740), .B2(n9079), .A(n8065), .ZN(n8066) );
  OAI21_X1 U9706 ( .B1(n9094), .B2(n8067), .A(n8066), .ZN(P2_U3282) );
  XNOR2_X1 U9707 ( .A(n8068), .B(n8074), .ZN(n10102) );
  INV_X1 U9708 ( .A(n10102), .ZN(n8087) );
  NAND2_X1 U9709 ( .A1(n8070), .A2(n8069), .ZN(n8072) );
  NAND2_X1 U9710 ( .A1(n8072), .A2(n8071), .ZN(n8073) );
  XOR2_X1 U9711 ( .A(n8074), .B(n8073), .Z(n8076) );
  OAI222_X1 U9712 ( .A1(n9053), .A2(n8077), .B1(n8076), .B2(n9049), .C1(n9051), 
        .C2(n8075), .ZN(n10099) );
  INV_X1 U9713 ( .A(n8083), .ZN(n10096) );
  INV_X1 U9714 ( .A(n8078), .ZN(n8079) );
  OAI21_X1 U9715 ( .B1(n10096), .B2(n8079), .A(n4379), .ZN(n10098) );
  OAI22_X1 U9716 ( .A1(n9079), .A2(n8081), .B1(n8080), .B2(n10025), .ZN(n8082)
         );
  AOI21_X1 U9717 ( .B1(n8083), .B2(n9092), .A(n8082), .ZN(n8084) );
  OAI21_X1 U9718 ( .B1(n10098), .B2(n8923), .A(n8084), .ZN(n8085) );
  AOI21_X1 U9719 ( .B1(n10099), .B2(n9079), .A(n8085), .ZN(n8086) );
  OAI21_X1 U9720 ( .B1(n9094), .B2(n8087), .A(n8086), .ZN(P2_U3284) );
  INV_X1 U9721 ( .A(n8090), .ZN(n8094) );
  AOI21_X1 U9722 ( .B1(n8090), .B2(n8089), .A(n8088), .ZN(n8091) );
  NOR2_X1 U9723 ( .A1(n8091), .A2(n9315), .ZN(n8092) );
  OAI21_X1 U9724 ( .B1(n8094), .B2(n8093), .A(n8092), .ZN(n8100) );
  NAND2_X1 U9725 ( .A1(n9308), .A2(n9752), .ZN(n8096) );
  OAI211_X1 U9726 ( .C1(n9325), .C2(n8175), .A(n8096), .B(n8095), .ZN(n8097)
         );
  AOI21_X1 U9727 ( .B1(n8098), .B2(n9329), .A(n8097), .ZN(n8099) );
  OAI211_X1 U9728 ( .C1(n8101), .C2(n9332), .A(n8100), .B(n8099), .ZN(P1_U3213) );
  INV_X1 U9729 ( .A(n8106), .ZN(n8103) );
  OAI21_X1 U9730 ( .B1(n8103), .B2(n8102), .A(n9322), .ZN(n8112) );
  AOI21_X1 U9731 ( .B1(n8106), .B2(n8105), .A(n8104), .ZN(n8111) );
  NAND2_X1 U9732 ( .A1(n9308), .A2(n9347), .ZN(n8107) );
  NAND2_X1 U9733 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9882) );
  OAI211_X1 U9734 ( .C1(n9325), .C2(n9570), .A(n8107), .B(n9882), .ZN(n8109)
         );
  NOR2_X1 U9735 ( .A1(n8119), .A2(n9332), .ZN(n8108) );
  AOI211_X1 U9736 ( .C1(n8117), .C2(n9329), .A(n8109), .B(n8108), .ZN(n8110)
         );
  OAI21_X1 U9737 ( .B1(n8112), .B2(n8111), .A(n8110), .ZN(P1_U3239) );
  NAND2_X1 U9738 ( .A1(n8113), .A2(n8114), .ZN(n8125) );
  INV_X1 U9739 ( .A(n8115), .ZN(n8584) );
  XNOR2_X1 U9740 ( .A(n8125), .B(n8584), .ZN(n9666) );
  AOI21_X1 U9741 ( .B1(n9662), .B2(n8116), .A(n8138), .ZN(n9663) );
  AOI22_X1 U9742 ( .A1(n9578), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n8117), .B2(
        n9759), .ZN(n8118) );
  OAI21_X1 U9743 ( .B1(n8119), .B2(n9568), .A(n8118), .ZN(n8122) );
  OAI21_X1 U9744 ( .B1(n8584), .B2(n4374), .A(n4567), .ZN(n8120) );
  AOI222_X1 U9745 ( .A1(n9747), .A2(n8120), .B1(n9347), .B2(n9754), .C1(n9345), 
        .C2(n9751), .ZN(n9665) );
  NOR2_X1 U9746 ( .A1(n9665), .A2(n9578), .ZN(n8121) );
  AOI211_X1 U9747 ( .C1(n9663), .C2(n9940), .A(n8122), .B(n8121), .ZN(n8123)
         );
  OAI21_X1 U9748 ( .B1(n9666), .B2(n9582), .A(n8123), .ZN(P1_U3276) );
  NAND2_X1 U9749 ( .A1(n8125), .A2(n8124), .ZN(n8127) );
  AND2_X1 U9750 ( .A1(n8127), .A2(n8126), .ZN(n8131) );
  AND2_X1 U9751 ( .A1(n8129), .A2(n8128), .ZN(n8130) );
  OAI21_X1 U9752 ( .B1(n8131), .B2(n8132), .A(n8130), .ZN(n9661) );
  OAI21_X1 U9753 ( .B1(n8134), .B2(n8133), .A(n8132), .ZN(n8135) );
  NAND3_X1 U9754 ( .A1(n4570), .A2(n9747), .A3(n8135), .ZN(n8137) );
  AOI22_X1 U9755 ( .A1(n9344), .A2(n9751), .B1(n9754), .B2(n9346), .ZN(n8136)
         );
  NAND2_X1 U9756 ( .A1(n8137), .A2(n8136), .ZN(n9658) );
  INV_X1 U9757 ( .A(n8138), .ZN(n8140) );
  INV_X1 U9758 ( .A(n9564), .ZN(n8139) );
  AOI211_X1 U9759 ( .C1(n5294), .C2(n8140), .A(n9975), .B(n8139), .ZN(n9659)
         );
  NAND2_X1 U9760 ( .A1(n9659), .A2(n9767), .ZN(n8142) );
  AOI22_X1 U9761 ( .A1(n9578), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n8179), .B2(
        n9759), .ZN(n8141) );
  OAI211_X1 U9762 ( .C1(n8176), .C2(n9568), .A(n8142), .B(n8141), .ZN(n8143)
         );
  AOI21_X1 U9763 ( .B1(n9658), .B2(n9945), .A(n8143), .ZN(n8144) );
  OAI21_X1 U9764 ( .B1(n9661), .B2(n9582), .A(n8144), .ZN(P1_U3275) );
  XNOR2_X1 U9765 ( .A(n8146), .B(n8145), .ZN(n8152) );
  OAI22_X1 U9766 ( .A1(n9995), .A2(n8155), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7655), .ZN(n8147) );
  AOI21_X1 U9767 ( .B1(n9998), .B2(n8852), .A(n8147), .ZN(n8148) );
  OAI21_X1 U9768 ( .B1(n8149), .B2(n10006), .A(n8148), .ZN(n8150) );
  AOI21_X1 U9769 ( .B1(n8834), .B2(n9179), .A(n8150), .ZN(n8151) );
  OAI21_X1 U9770 ( .B1(n8152), .B2(n8836), .A(n8151), .ZN(P2_U3236) );
  XOR2_X1 U9771 ( .A(n8153), .B(n8160), .Z(n8154) );
  OAI222_X1 U9772 ( .A1(n9053), .A2(n8828), .B1(n9051), .B2(n8155), .C1(n9049), 
        .C2(n8154), .ZN(n8248) );
  INV_X1 U9773 ( .A(n8248), .ZN(n8169) );
  OR2_X1 U9774 ( .A1(n8264), .A2(n8850), .ZN(n8158) );
  NAND2_X1 U9775 ( .A1(n8159), .A2(n8158), .ZN(n8161) );
  NAND2_X1 U9776 ( .A1(n8161), .A2(n8160), .ZN(n8224) );
  OAI21_X1 U9777 ( .B1(n8161), .B2(n8160), .A(n8224), .ZN(n8250) );
  INV_X1 U9778 ( .A(n8162), .ZN(n8163) );
  INV_X1 U9779 ( .A(n8833), .ZN(n8246) );
  OAI21_X1 U9780 ( .B1(n8163), .B2(n8246), .A(n8232), .ZN(n8247) );
  OAI22_X1 U9781 ( .A1(n9079), .A2(n8164), .B1(n8831), .B2(n10025), .ZN(n8165)
         );
  AOI21_X1 U9782 ( .B1(n8833), .B2(n9092), .A(n8165), .ZN(n8166) );
  OAI21_X1 U9783 ( .B1(n8247), .B2(n8923), .A(n8166), .ZN(n8167) );
  AOI21_X1 U9784 ( .B1(n8250), .B2(n9006), .A(n8167), .ZN(n8168) );
  OAI21_X1 U9785 ( .B1(n8169), .B2(n9017), .A(n8168), .ZN(P2_U3281) );
  XOR2_X1 U9786 ( .A(n8171), .B(n8170), .Z(n8172) );
  XNOR2_X1 U9787 ( .A(n8173), .B(n8172), .ZN(n8181) );
  NAND2_X1 U9788 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9894) );
  NAND2_X1 U9789 ( .A1(n9264), .A2(n9344), .ZN(n8174) );
  OAI211_X1 U9790 ( .C1(n9326), .C2(n8175), .A(n9894), .B(n8174), .ZN(n8178)
         );
  NOR2_X1 U9791 ( .A1(n8176), .A2(n9332), .ZN(n8177) );
  AOI211_X1 U9792 ( .C1(n8179), .C2(n9329), .A(n8178), .B(n8177), .ZN(n8180)
         );
  OAI21_X1 U9793 ( .B1(n8181), .B2(n9315), .A(n8180), .ZN(P1_U3224) );
  NAND2_X1 U9794 ( .A1(n8183), .A2(n8182), .ZN(n8185) );
  NAND2_X1 U9795 ( .A1(n8185), .A2(n8184), .ZN(n8187) );
  XNOR2_X1 U9796 ( .A(n8271), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8186) );
  NOR2_X1 U9797 ( .A1(n8186), .A2(n8187), .ZN(n8272) );
  AOI21_X1 U9798 ( .B1(n8187), .B2(n8186), .A(n8272), .ZN(n8200) );
  NAND2_X1 U9799 ( .A1(n8189), .A2(n8188), .ZN(n8191) );
  NAND2_X1 U9800 ( .A1(n8191), .A2(n8190), .ZN(n8194) );
  NAND2_X1 U9801 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8271), .ZN(n8192) );
  OAI21_X1 U9802 ( .B1(n8271), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8192), .ZN(
        n8193) );
  NOR2_X1 U9803 ( .A1(n8193), .A2(n8194), .ZN(n8267) );
  AOI211_X1 U9804 ( .C1(n8194), .C2(n8193), .A(n8267), .B(n9725), .ZN(n8195)
         );
  INV_X1 U9805 ( .A(n8195), .ZN(n8199) );
  INV_X1 U9806 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8196) );
  NAND2_X1 U9807 ( .A1(P2_U3152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8765) );
  OAI21_X1 U9808 ( .B1(n9714), .B2(n8196), .A(n8765), .ZN(n8197) );
  AOI21_X1 U9809 ( .B1(n9731), .B2(n8271), .A(n8197), .ZN(n8198) );
  OAI211_X1 U9810 ( .C1(n8200), .C2(n10011), .A(n8199), .B(n8198), .ZN(
        P2_U3261) );
  OAI21_X1 U9811 ( .B1(n8588), .B2(n8202), .A(n8201), .ZN(n8203) );
  AOI222_X1 U9812 ( .A1(n9747), .A2(n8203), .B1(n9344), .B2(n9754), .C1(n9343), 
        .C2(n9751), .ZN(n9652) );
  INV_X1 U9813 ( .A(n9563), .ZN(n8205) );
  INV_X1 U9814 ( .A(n9553), .ZN(n8204) );
  AOI21_X1 U9815 ( .B1(n9647), .B2(n8205), .A(n8204), .ZN(n9648) );
  NOR2_X1 U9816 ( .A1(n8206), .A2(n9568), .ZN(n8208) );
  INV_X1 U9817 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9369) );
  OAI22_X1 U9818 ( .A1(n9945), .A2(n9369), .B1(n9310), .B2(n9949), .ZN(n8207)
         );
  AOI211_X1 U9819 ( .C1(n9648), .C2(n9940), .A(n8208), .B(n8207), .ZN(n8213)
         );
  OR2_X1 U9820 ( .A1(n8210), .A2(n8209), .ZN(n9649) );
  INV_X1 U9821 ( .A(n9582), .ZN(n9427) );
  NAND3_X1 U9822 ( .A1(n9649), .A2(n8211), .A3(n9427), .ZN(n8212) );
  OAI211_X1 U9823 ( .C1(n9652), .C2(n9578), .A(n8213), .B(n8212), .ZN(P1_U3273) );
  INV_X1 U9824 ( .A(n8214), .ZN(n8218) );
  OAI222_X1 U9825 ( .A1(n8661), .A2(n8216), .B1(n8665), .B2(n8218), .C1(n8215), 
        .C2(P2_U3152), .ZN(P2_U3333) );
  OAI222_X1 U9826 ( .A1(P1_U3084), .A2(n8219), .B1(n9699), .B2(n8218), .C1(
        n8217), .C2(n9704), .ZN(P1_U3328) );
  INV_X1 U9827 ( .A(n8220), .ZN(n8241) );
  OAI222_X1 U9828 ( .A1(n9212), .A2(n8241), .B1(P2_U3152), .B2(n8222), .C1(
        n8221), .C2(n8661), .ZN(P2_U3332) );
  OR2_X1 U9829 ( .A1(n8833), .A2(n8849), .ZN(n8223) );
  XNOR2_X1 U9830 ( .A(n8289), .B(n6295), .ZN(n9171) );
  INV_X1 U9831 ( .A(n8225), .ZN(n8231) );
  NAND2_X1 U9832 ( .A1(n8226), .A2(n8288), .ZN(n8227) );
  AOI21_X1 U9833 ( .B1(n8285), .B2(n8227), .A(n9049), .ZN(n8230) );
  OAI22_X1 U9834 ( .A1(n8228), .A2(n9051), .B1(n8766), .B2(n9053), .ZN(n8229)
         );
  AOI211_X1 U9835 ( .C1(n9171), .C2(n8231), .A(n8230), .B(n8229), .ZN(n9177)
         );
  AND2_X1 U9836 ( .A1(n8232), .A2(n9172), .ZN(n8233) );
  OR2_X1 U9837 ( .A1(n8233), .A2(n8282), .ZN(n9174) );
  INV_X1 U9838 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8234) );
  OAI22_X1 U9839 ( .A1(n9079), .A2(n8234), .B1(n8769), .B2(n10025), .ZN(n8235)
         );
  AOI21_X1 U9840 ( .B1(n9172), .B2(n9092), .A(n8235), .ZN(n8236) );
  OAI21_X1 U9841 ( .B1(n9174), .B2(n8923), .A(n8236), .ZN(n8237) );
  AOI21_X1 U9842 ( .B1(n9171), .B2(n8238), .A(n8237), .ZN(n8239) );
  OAI21_X1 U9843 ( .B1(n9177), .B2(n9017), .A(n8239), .ZN(P2_U3280) );
  OAI222_X1 U9844 ( .A1(n8242), .A2(P1_U3084), .B1(n9699), .B2(n8241), .C1(
        n8240), .C2(n9704), .ZN(P1_U3327) );
  NAND2_X1 U9845 ( .A1(n8320), .A2(n8243), .ZN(n8244) );
  OAI211_X1 U9846 ( .C1(n9704), .C2(n8245), .A(n8244), .B(n9799), .ZN(P1_U3326) );
  INV_X1 U9847 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8251) );
  OAI22_X1 U9848 ( .A1(n8247), .A2(n10097), .B1(n8246), .B2(n10095), .ZN(n8249) );
  AOI211_X1 U9849 ( .C1(n10101), .C2(n8250), .A(n8249), .B(n8248), .ZN(n8253)
         );
  MUX2_X1 U9850 ( .A(n8251), .B(n8253), .S(n10105), .Z(n8252) );
  INV_X1 U9851 ( .A(n8252), .ZN(P2_U3496) );
  MUX2_X1 U9852 ( .A(n5866), .B(n8253), .S(n10119), .Z(n8254) );
  INV_X1 U9853 ( .A(n8254), .ZN(P2_U3535) );
  INV_X1 U9854 ( .A(n8255), .ZN(n8256) );
  AOI21_X1 U9855 ( .B1(n8258), .B2(n8257), .A(n8256), .ZN(n8266) );
  AOI21_X1 U9856 ( .B1(n8734), .B2(n8260), .A(n8259), .ZN(n8261) );
  OAI21_X1 U9857 ( .B1(n8262), .B2(n10006), .A(n8261), .ZN(n8263) );
  AOI21_X1 U9858 ( .B1(n8264), .B2(n8834), .A(n8263), .ZN(n8265) );
  OAI21_X1 U9859 ( .B1(n8266), .B2(n8836), .A(n8265), .ZN(P2_U3217) );
  NAND2_X1 U9860 ( .A1(n8885), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8268) );
  OAI21_X1 U9861 ( .B1(n8885), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8268), .ZN(
        n8269) );
  AOI211_X1 U9862 ( .C1(n8270), .C2(n8269), .A(n8884), .B(n9725), .ZN(n8281)
         );
  XNOR2_X1 U9863 ( .A(n8880), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8276) );
  OR2_X1 U9864 ( .A1(n8271), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8274) );
  INV_X1 U9865 ( .A(n8272), .ZN(n8273) );
  NAND2_X1 U9866 ( .A1(n8276), .A2(n8275), .ZN(n8879) );
  OAI211_X1 U9867 ( .C1(n8276), .C2(n8275), .A(n10007), .B(n8879), .ZN(n8279)
         );
  NOR2_X1 U9868 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8313), .ZN(n8277) );
  AOI21_X1 U9869 ( .B1(n10013), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8277), .ZN(
        n8278) );
  OAI211_X1 U9870 ( .C1(n10009), .C2(n8880), .A(n8279), .B(n8278), .ZN(n8280)
         );
  OR2_X1 U9871 ( .A1(n8281), .A2(n8280), .ZN(P2_U3262) );
  INV_X1 U9872 ( .A(n8282), .ZN(n8283) );
  INV_X1 U9873 ( .A(n9167), .ZN(n8292) );
  AOI211_X1 U9874 ( .C1(n9167), .C2(n8283), .A(n10097), .B(n8299), .ZN(n9166)
         );
  NAND2_X1 U9875 ( .A1(n8285), .A2(n8284), .ZN(n8286) );
  XNOR2_X1 U9876 ( .A(n8286), .B(n8290), .ZN(n8287) );
  OAI222_X1 U9877 ( .A1(n9053), .A2(n8667), .B1(n8287), .B2(n9049), .C1(n9051), 
        .C2(n8828), .ZN(n9165) );
  AOI21_X1 U9878 ( .B1(n9166), .B2(n10027), .A(n9165), .ZN(n8297) );
  OAI21_X1 U9879 ( .B1(n8291), .B2(n8290), .A(n8298), .ZN(n9164) );
  NOR2_X1 U9880 ( .A1(n8292), .A2(n9063), .ZN(n8295) );
  OAI22_X1 U9881 ( .A1(n9079), .A2(n8293), .B1(n8316), .B2(n10025), .ZN(n8294)
         );
  AOI211_X1 U9882 ( .C1(n9164), .C2(n9006), .A(n8295), .B(n8294), .ZN(n8296)
         );
  OAI21_X1 U9883 ( .B1(n8297), .B2(n9017), .A(n8296), .ZN(P2_U3279) );
  XNOR2_X1 U9884 ( .A(n8670), .B(n4327), .ZN(n9163) );
  INV_X1 U9885 ( .A(n8299), .ZN(n8301) );
  INV_X1 U9886 ( .A(n9161), .ZN(n8666) );
  INV_X1 U9887 ( .A(n9088), .ZN(n8300) );
  AOI211_X1 U9888 ( .C1(n9161), .C2(n8301), .A(n10097), .B(n8300), .ZN(n9160)
         );
  NOR2_X1 U9889 ( .A1(n8666), .A2(n9063), .ZN(n8304) );
  OAI22_X1 U9890 ( .A1(n9079), .A2(n8302), .B1(n8810), .B2(n10025), .ZN(n8303)
         );
  AOI211_X1 U9891 ( .C1(n9160), .C2(n9043), .A(n8304), .B(n8303), .ZN(n8308)
         );
  XNOR2_X1 U9892 ( .A(n8305), .B(n4327), .ZN(n8306) );
  OAI222_X1 U9893 ( .A1(n9053), .A2(n8807), .B1(n9051), .B2(n8766), .C1(n9049), 
        .C2(n8306), .ZN(n9159) );
  NAND2_X1 U9894 ( .A1(n9159), .A2(n9079), .ZN(n8307) );
  OAI211_X1 U9895 ( .C1(n9163), .C2(n9094), .A(n8308), .B(n8307), .ZN(P2_U3278) );
  INV_X1 U9896 ( .A(n8309), .ZN(n8664) );
  AOI21_X1 U9897 ( .B1(P2_DATAO_REG_28__SCAN_IN), .B2(n9697), .A(n9798), .ZN(
        n8310) );
  OAI21_X1 U9898 ( .B1(n8664), .B2(n9699), .A(n8310), .ZN(P1_U3325) );
  XNOR2_X1 U9899 ( .A(n8312), .B(n8311), .ZN(n8319) );
  OAI22_X1 U9900 ( .A1(n9995), .A2(n8667), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8313), .ZN(n8314) );
  AOI21_X1 U9901 ( .B1(n9998), .B2(n8848), .A(n8314), .ZN(n8315) );
  OAI21_X1 U9902 ( .B1(n8316), .B2(n10006), .A(n8315), .ZN(n8317) );
  AOI21_X1 U9903 ( .B1(n9167), .B2(n8834), .A(n8317), .ZN(n8318) );
  OAI21_X1 U9904 ( .B1(n8319), .B2(n8836), .A(n8318), .ZN(P2_U3230) );
  INV_X1 U9905 ( .A(n8320), .ZN(n8322) );
  OAI222_X1 U9906 ( .A1(n9212), .A2(n8322), .B1(n8687), .B2(P2_U3152), .C1(
        n8321), .C2(n8661), .ZN(P2_U3331) );
  NAND2_X1 U9907 ( .A1(n9596), .A2(n8323), .ZN(n8326) );
  NAND2_X1 U9908 ( .A1(n9335), .A2(n4388), .ZN(n8325) );
  NAND2_X1 U9909 ( .A1(n8326), .A2(n8325), .ZN(n8328) );
  XNOR2_X1 U9910 ( .A(n8328), .B(n4311), .ZN(n8331) );
  AOI22_X1 U9911 ( .A1(n9596), .A2(n8329), .B1(n6544), .B2(n9335), .ZN(n8330)
         );
  XNOR2_X1 U9912 ( .A(n8331), .B(n8330), .ZN(n8332) );
  INV_X1 U9913 ( .A(n8332), .ZN(n8336) );
  NAND3_X1 U9914 ( .A1(n8336), .A2(n9322), .A3(n8335), .ZN(n8340) );
  AOI22_X1 U9915 ( .A1(n9336), .A2(n9308), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n8334) );
  NAND2_X1 U9916 ( .A1(n9329), .A2(n9424), .ZN(n8333) );
  OAI211_X1 U9917 ( .C1(n9418), .C2(n9325), .A(n8334), .B(n8333), .ZN(n8338)
         );
  NOR3_X1 U9918 ( .A1(n8336), .A2(n8335), .A3(n9315), .ZN(n8337) );
  AOI211_X1 U9919 ( .C1(n9596), .C2(n9313), .A(n8338), .B(n8337), .ZN(n8339)
         );
  NAND2_X1 U9920 ( .A1(n9203), .A2(n5454), .ZN(n8343) );
  NAND2_X1 U9921 ( .A1(n8344), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8342) );
  INV_X1 U9922 ( .A(n9403), .ZN(n8410) );
  NAND2_X1 U9923 ( .A1(n9583), .A2(n8410), .ZN(n8600) );
  NAND2_X1 U9924 ( .A1(n9206), .A2(n5454), .ZN(n8346) );
  NAND2_X1 U9925 ( .A1(n8344), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8345) );
  OR2_X1 U9926 ( .A1(n9410), .A2(n5530), .ZN(n8599) );
  NAND2_X1 U9927 ( .A1(n8626), .A2(n8347), .ZN(n8348) );
  NAND3_X1 U9928 ( .A1(n8542), .A2(n8537), .A3(n8348), .ZN(n8631) );
  AND2_X1 U9929 ( .A1(n8349), .A2(n8528), .ZN(n8625) );
  INV_X1 U9930 ( .A(n8625), .ZN(n8402) );
  NAND2_X1 U9931 ( .A1(n8350), .A2(n9338), .ZN(n8519) );
  INV_X1 U9932 ( .A(n8351), .ZN(n8352) );
  NAND2_X1 U9933 ( .A1(n8519), .A2(n8352), .ZN(n8353) );
  NAND3_X1 U9934 ( .A1(n8530), .A2(n4560), .A3(n8353), .ZN(n8627) );
  INV_X1 U9935 ( .A(n8501), .ZN(n8354) );
  NAND2_X1 U9936 ( .A1(n8511), .A2(n8354), .ZN(n8355) );
  AND2_X1 U9937 ( .A1(n8355), .A2(n8506), .ZN(n8356) );
  AND2_X1 U9938 ( .A1(n8508), .A2(n8356), .ZN(n8512) );
  INV_X1 U9939 ( .A(n8512), .ZN(n8363) );
  AND2_X1 U9940 ( .A1(n8499), .A2(n8357), .ZN(n8476) );
  NAND2_X1 U9941 ( .A1(n8502), .A2(n8365), .ZN(n8505) );
  AND2_X1 U9942 ( .A1(n9518), .A2(n8500), .ZN(n8504) );
  OAI211_X1 U9943 ( .C1(n8476), .C2(n8505), .A(n8511), .B(n8504), .ZN(n8358)
         );
  INV_X1 U9944 ( .A(n8358), .ZN(n8359) );
  OAI211_X1 U9945 ( .C1(n8363), .C2(n8359), .A(n8412), .B(n8515), .ZN(n8360)
         );
  INV_X1 U9946 ( .A(n8360), .ZN(n8361) );
  NAND2_X1 U9947 ( .A1(n8519), .A2(n8361), .ZN(n8624) );
  OR2_X1 U9948 ( .A1(n8363), .A2(n8362), .ZN(n8622) );
  NAND2_X1 U9949 ( .A1(n8365), .A2(n8364), .ZN(n8495) );
  INV_X1 U9950 ( .A(n8480), .ZN(n8494) );
  OR2_X1 U9951 ( .A1(n8495), .A2(n8494), .ZN(n8395) );
  AND2_X1 U9952 ( .A1(n8387), .A2(n8366), .ZN(n8491) );
  INV_X1 U9953 ( .A(n8491), .ZN(n8386) );
  NAND2_X1 U9954 ( .A1(n8456), .A2(n8452), .ZN(n8460) );
  NAND2_X1 U9955 ( .A1(n8460), .A2(n8466), .ZN(n8368) );
  NAND2_X1 U9956 ( .A1(n6600), .A2(n8367), .ZN(n8485) );
  NAND3_X1 U9957 ( .A1(n8486), .A2(n8368), .A3(n8485), .ZN(n8369) );
  NOR2_X1 U9958 ( .A1(n8386), .A2(n8369), .ZN(n8385) );
  NAND4_X1 U9959 ( .A1(n8385), .A2(n8489), .A3(n8458), .A4(n8425), .ZN(n8370)
         );
  OR2_X1 U9960 ( .A1(n8395), .A2(n8370), .ZN(n8619) );
  INV_X1 U9961 ( .A(n8605), .ZN(n8371) );
  INV_X1 U9962 ( .A(n8430), .ZN(n8614) );
  AOI211_X1 U9963 ( .C1(n8373), .C2(n8371), .A(n8614), .B(n8604), .ZN(n8384)
         );
  NAND2_X1 U9964 ( .A1(n8373), .A2(n8372), .ZN(n8613) );
  INV_X1 U9965 ( .A(n8613), .ZN(n8382) );
  NAND2_X1 U9966 ( .A1(n6526), .A2(n6524), .ZN(n8375) );
  NAND2_X1 U9967 ( .A1(n6529), .A2(n4393), .ZN(n8374) );
  NAND3_X1 U9968 ( .A1(n8375), .A2(n8374), .A3(n8640), .ZN(n8376) );
  NAND2_X1 U9969 ( .A1(n8377), .A2(n8376), .ZN(n8379) );
  OAI21_X1 U9970 ( .B1(n8380), .B2(n8379), .A(n8378), .ZN(n8381) );
  NAND2_X1 U9971 ( .A1(n8382), .A2(n8381), .ZN(n8383) );
  AND2_X1 U9972 ( .A1(n8384), .A2(n8383), .ZN(n8396) );
  INV_X1 U9973 ( .A(n8385), .ZN(n8391) );
  AND2_X1 U9974 ( .A1(n8454), .A2(n8451), .ZN(n8461) );
  AND2_X1 U9975 ( .A1(n8466), .A2(n8461), .ZN(n8390) );
  OR2_X1 U9976 ( .A1(n8386), .A2(n8471), .ZN(n8389) );
  NAND2_X1 U9977 ( .A1(n8472), .A2(n8470), .ZN(n8388) );
  NAND2_X1 U9978 ( .A1(n8388), .A2(n8387), .ZN(n8477) );
  OAI211_X1 U9979 ( .C1(n8391), .C2(n8390), .A(n8389), .B(n8477), .ZN(n8392)
         );
  NAND2_X1 U9980 ( .A1(n8392), .A2(n8489), .ZN(n8393) );
  AND3_X1 U9981 ( .A1(n8393), .A2(n8481), .A3(n8478), .ZN(n8394) );
  OR2_X1 U9982 ( .A1(n8395), .A2(n8394), .ZN(n8617) );
  OAI21_X1 U9983 ( .B1(n8619), .B2(n8396), .A(n8617), .ZN(n8397) );
  INV_X1 U9984 ( .A(n8397), .ZN(n8398) );
  NOR2_X1 U9985 ( .A1(n8622), .A2(n8398), .ZN(n8399) );
  NOR2_X1 U9986 ( .A1(n8624), .A2(n8399), .ZN(n8400) );
  NOR2_X1 U9987 ( .A1(n8627), .A2(n8400), .ZN(n8401) );
  OR2_X1 U9988 ( .A1(n8402), .A2(n8401), .ZN(n8403) );
  NOR2_X1 U9989 ( .A1(n9437), .A2(n8403), .ZN(n8404) );
  NOR2_X1 U9990 ( .A1(n8631), .A2(n8404), .ZN(n8406) );
  NAND2_X1 U9991 ( .A1(n8405), .A2(n8541), .ZN(n8635) );
  OAI21_X1 U9992 ( .B1(n8406), .B2(n8635), .A(n8633), .ZN(n8407) );
  NAND2_X1 U9993 ( .A1(n8599), .A2(n8407), .ZN(n8408) );
  NAND2_X1 U9994 ( .A1(n9410), .A2(n5530), .ZN(n8597) );
  NAND2_X1 U9995 ( .A1(n8408), .A2(n8597), .ZN(n8409) );
  NAND2_X1 U9996 ( .A1(n8600), .A2(n8409), .ZN(n8411) );
  NAND2_X1 U9997 ( .A1(n8411), .A2(n8639), .ZN(n8649) );
  NAND2_X1 U9998 ( .A1(n8649), .A2(n9497), .ZN(n8648) );
  OAI211_X1 U9999 ( .C1(n8413), .C2(n8412), .A(n8528), .B(n8519), .ZN(n8414)
         );
  MUX2_X1 U10000 ( .A(n8414), .B(n8627), .S(n8536), .Z(n8415) );
  INV_X1 U10001 ( .A(n8415), .ZN(n8523) );
  INV_X1 U10002 ( .A(n9573), .ZN(n9561) );
  NAND2_X1 U10003 ( .A1(n8480), .A2(n8489), .ZN(n8416) );
  NAND2_X1 U10004 ( .A1(n8416), .A2(n8481), .ZN(n8417) );
  AOI21_X1 U10005 ( .B1(n9561), .B2(n8417), .A(n8536), .ZN(n8418) );
  NAND2_X1 U10006 ( .A1(n8418), .A2(n8476), .ZN(n8498) );
  NAND2_X1 U10007 ( .A1(n8419), .A2(n8427), .ZN(n8424) );
  INV_X1 U10008 ( .A(n8420), .ZN(n8421) );
  NAND2_X1 U10009 ( .A1(n8422), .A2(n8421), .ZN(n8423) );
  AND2_X1 U10010 ( .A1(n8423), .A2(n8429), .ZN(n8607) );
  NAND2_X1 U10011 ( .A1(n8424), .A2(n8607), .ZN(n8426) );
  NAND4_X1 U10012 ( .A1(n8426), .A2(n8536), .A3(n8610), .A4(n8425), .ZN(n8450)
         );
  NAND2_X1 U10013 ( .A1(n8428), .A2(n8427), .ZN(n8448) );
  AND4_X1 U10014 ( .A1(n8430), .A2(n8608), .A3(n8429), .A4(n8556), .ZN(n8447)
         );
  NAND2_X1 U10015 ( .A1(n8431), .A2(n8556), .ZN(n8440) );
  OAI21_X1 U10016 ( .B1(n8440), .B2(n9352), .A(n8434), .ZN(n8433) );
  OR2_X1 U10017 ( .A1(n8431), .A2(n8556), .ZN(n8435) );
  OAI21_X1 U10018 ( .B1(n8435), .B2(n8438), .A(n9967), .ZN(n8432) );
  NAND2_X1 U10019 ( .A1(n8433), .A2(n8432), .ZN(n8445) );
  OAI22_X1 U10020 ( .A1(n8435), .A2(n8434), .B1(n8438), .B2(n8556), .ZN(n8437)
         );
  NAND2_X1 U10021 ( .A1(n8437), .A2(n8436), .ZN(n8444) );
  NAND2_X1 U10022 ( .A1(n8438), .A2(n8556), .ZN(n8439) );
  OAI21_X1 U10023 ( .B1(n8440), .B2(n9967), .A(n8439), .ZN(n8442) );
  NAND2_X1 U10024 ( .A1(n8442), .A2(n8441), .ZN(n8443) );
  NAND3_X1 U10025 ( .A1(n8445), .A2(n8444), .A3(n8443), .ZN(n8446) );
  AOI21_X1 U10026 ( .B1(n8448), .B2(n8447), .A(n8446), .ZN(n8449) );
  NAND2_X1 U10027 ( .A1(n8450), .A2(n8449), .ZN(n8459) );
  NAND2_X1 U10028 ( .A1(n8459), .A2(n8451), .ZN(n8453) );
  NAND3_X1 U10029 ( .A1(n8453), .A2(n8452), .A3(n8458), .ZN(n8455) );
  NAND3_X1 U10030 ( .A1(n8455), .A2(n8466), .A3(n8454), .ZN(n8457) );
  NAND3_X1 U10031 ( .A1(n8457), .A2(n8486), .A3(n8456), .ZN(n8464) );
  NAND2_X1 U10032 ( .A1(n8459), .A2(n8458), .ZN(n8462) );
  AOI21_X1 U10033 ( .B1(n8462), .B2(n8461), .A(n8460), .ZN(n8463) );
  MUX2_X1 U10034 ( .A(n8464), .B(n8463), .S(n8536), .Z(n8465) );
  INV_X1 U10035 ( .A(n8465), .ZN(n8469) );
  OAI211_X1 U10036 ( .C1(n8466), .C2(n8556), .A(n8487), .B(n8579), .ZN(n8467)
         );
  INV_X1 U10037 ( .A(n8467), .ZN(n8468) );
  NAND2_X1 U10038 ( .A1(n8469), .A2(n8468), .ZN(n8492) );
  NAND3_X1 U10039 ( .A1(n8492), .A2(n8471), .A3(n8470), .ZN(n8474) );
  NAND3_X1 U10040 ( .A1(n8478), .A2(n8472), .A3(n8556), .ZN(n8473) );
  AOI21_X1 U10041 ( .B1(n8474), .B2(n8491), .A(n8473), .ZN(n8475) );
  NAND3_X1 U10042 ( .A1(n8476), .A2(n8475), .A3(n8481), .ZN(n8497) );
  NAND2_X1 U10043 ( .A1(n8478), .A2(n8477), .ZN(n8479) );
  NAND3_X1 U10044 ( .A1(n8480), .A2(n8489), .A3(n8479), .ZN(n8482) );
  NAND2_X1 U10045 ( .A1(n8482), .A2(n8481), .ZN(n8483) );
  NOR2_X1 U10046 ( .A1(n9573), .A2(n8483), .ZN(n8484) );
  OR3_X1 U10047 ( .A1(n8495), .A2(n8484), .A3(n8556), .ZN(n8496) );
  NAND2_X1 U10048 ( .A1(n8486), .A2(n8485), .ZN(n8488) );
  AOI21_X1 U10049 ( .B1(n8488), .B2(n8487), .A(n8556), .ZN(n8490) );
  NAND4_X1 U10050 ( .A1(n8492), .A2(n8491), .A3(n8490), .A4(n8489), .ZN(n8493)
         );
  NAND2_X1 U10051 ( .A1(n8500), .A2(n8499), .ZN(n8503) );
  INV_X1 U10052 ( .A(n8506), .ZN(n8507) );
  AOI21_X1 U10053 ( .B1(n8514), .B2(n9518), .A(n8507), .ZN(n8510) );
  NAND2_X1 U10054 ( .A1(n8515), .A2(n8511), .ZN(n8509) );
  OAI21_X1 U10055 ( .B1(n8510), .B2(n8509), .A(n8508), .ZN(n8518) );
  INV_X1 U10056 ( .A(n8511), .ZN(n8513) );
  OAI21_X1 U10057 ( .B1(n8514), .B2(n8513), .A(n8512), .ZN(n8516) );
  NAND2_X1 U10058 ( .A1(n8516), .A2(n8515), .ZN(n8517) );
  MUX2_X1 U10059 ( .A(n8518), .B(n8517), .S(n8556), .Z(n8521) );
  AND3_X1 U10060 ( .A1(n4560), .A2(n9489), .A3(n8519), .ZN(n8520) );
  NAND2_X1 U10061 ( .A1(n8521), .A2(n8520), .ZN(n8522) );
  NAND2_X1 U10062 ( .A1(n8523), .A2(n8522), .ZN(n8524) );
  NOR2_X1 U10063 ( .A1(n8530), .A2(n9337), .ZN(n8525) );
  OR2_X1 U10064 ( .A1(n9607), .A2(n8525), .ZN(n8526) );
  NAND2_X1 U10065 ( .A1(n9431), .A2(n8527), .ZN(n8535) );
  NAND2_X1 U10066 ( .A1(n9607), .A2(n8528), .ZN(n8529) );
  NAND2_X1 U10067 ( .A1(n8537), .A2(n8529), .ZN(n8533) );
  NAND2_X1 U10068 ( .A1(n8530), .A2(n9337), .ZN(n8531) );
  NAND2_X1 U10069 ( .A1(n8626), .A2(n8531), .ZN(n8532) );
  MUX2_X1 U10070 ( .A(n8533), .B(n8532), .S(n8556), .Z(n8534) );
  AND2_X1 U10071 ( .A1(n8535), .A2(n8534), .ZN(n8540) );
  MUX2_X1 U10072 ( .A(n8537), .B(n8626), .S(n8536), .Z(n8538) );
  MUX2_X1 U10073 ( .A(n8542), .B(n8541), .S(n8556), .Z(n8543) );
  NAND2_X1 U10074 ( .A1(n8544), .A2(n8543), .ZN(n8552) );
  NAND2_X1 U10075 ( .A1(n8552), .A2(n9418), .ZN(n8545) );
  INV_X1 U10076 ( .A(n9418), .ZN(n9334) );
  NAND2_X1 U10077 ( .A1(n9334), .A2(n8556), .ZN(n8548) );
  NAND2_X1 U10078 ( .A1(n9591), .A2(n8556), .ZN(n8546) );
  NOR2_X1 U10079 ( .A1(n8552), .A2(n8546), .ZN(n8547) );
  AOI21_X1 U10080 ( .B1(n8549), .B2(n8548), .A(n8547), .ZN(n8553) );
  NAND2_X1 U10081 ( .A1(n8599), .A2(n9403), .ZN(n8550) );
  AND2_X1 U10082 ( .A1(n8550), .A2(n9583), .ZN(n8554) );
  OR2_X1 U10083 ( .A1(n9418), .A2(n8556), .ZN(n8551) );
  INV_X1 U10084 ( .A(n8554), .ZN(n8638) );
  OAI21_X1 U10085 ( .B1(n8638), .B2(n8556), .A(n8555), .ZN(n8562) );
  NAND2_X1 U10086 ( .A1(n8563), .A2(n6516), .ZN(n8561) );
  NAND2_X1 U10087 ( .A1(n9403), .A2(n9333), .ZN(n8557) );
  AND2_X1 U10088 ( .A1(n9410), .A2(n8557), .ZN(n8632) );
  NAND2_X1 U10089 ( .A1(n8600), .A2(n8632), .ZN(n8559) );
  AND4_X1 U10090 ( .A1(n8559), .A2(n8640), .A3(n8558), .A4(n8639), .ZN(n8560)
         );
  OAI211_X1 U10091 ( .C1(n8563), .C2(n8562), .A(n8561), .B(n8560), .ZN(n8646)
         );
  NOR2_X1 U10092 ( .A1(n8565), .A2(n8564), .ZN(n8570) );
  NOR2_X1 U10093 ( .A1(n8566), .A2(n7018), .ZN(n8568) );
  NAND4_X1 U10094 ( .A1(n8570), .A2(n8569), .A3(n8568), .A4(n8567), .ZN(n8572)
         );
  NOR2_X1 U10095 ( .A1(n8572), .A2(n5155), .ZN(n8573) );
  NAND4_X1 U10096 ( .A1(n8576), .A2(n8575), .A3(n8574), .A4(n8573), .ZN(n8577)
         );
  NOR2_X1 U10097 ( .A1(n8578), .A2(n8577), .ZN(n8580) );
  AND4_X1 U10098 ( .A1(n8581), .A2(n9749), .A3(n8580), .A4(n8579), .ZN(n8582)
         );
  NAND4_X1 U10099 ( .A1(n8585), .A2(n8584), .A3(n8583), .A4(n8582), .ZN(n8586)
         );
  NOR2_X1 U10100 ( .A1(n8586), .A2(n9573), .ZN(n8587) );
  NAND4_X1 U10101 ( .A1(n9536), .A2(n9547), .A3(n8588), .A4(n8587), .ZN(n8589)
         );
  NOR2_X1 U10102 ( .A1(n9515), .A2(n8589), .ZN(n8590) );
  NAND3_X1 U10103 ( .A1(n9489), .A2(n9503), .A3(n8590), .ZN(n8591) );
  NOR3_X1 U10104 ( .A1(n9464), .A2(n9475), .A3(n8591), .ZN(n8592) );
  NAND2_X1 U10105 ( .A1(n8593), .A2(n8592), .ZN(n8594) );
  OR3_X1 U10106 ( .A1(n9425), .A2(n9437), .A3(n8594), .ZN(n8595) );
  NOR2_X1 U10107 ( .A1(n8596), .A2(n8595), .ZN(n8598) );
  AND3_X1 U10108 ( .A1(n8599), .A2(n8598), .A3(n8597), .ZN(n8601) );
  NAND3_X1 U10109 ( .A1(n8639), .A2(n8601), .A3(n8600), .ZN(n8603) );
  NAND2_X1 U10110 ( .A1(n8603), .A2(n8602), .ZN(n8644) );
  INV_X1 U10111 ( .A(n8604), .ZN(n8606) );
  NAND3_X1 U10112 ( .A1(n7203), .A2(n8606), .A3(n8605), .ZN(n8616) );
  INV_X1 U10113 ( .A(n8607), .ZN(n8611) );
  INV_X1 U10114 ( .A(n8608), .ZN(n8609) );
  AOI21_X1 U10115 ( .B1(n8611), .B2(n8610), .A(n8609), .ZN(n8612) );
  NAND2_X1 U10116 ( .A1(n8613), .A2(n8612), .ZN(n8615) );
  AOI21_X1 U10117 ( .B1(n8616), .B2(n8615), .A(n8614), .ZN(n8618) );
  OAI21_X1 U10118 ( .B1(n8619), .B2(n8618), .A(n8617), .ZN(n8620) );
  INV_X1 U10119 ( .A(n8620), .ZN(n8621) );
  NOR2_X1 U10120 ( .A1(n8622), .A2(n8621), .ZN(n8623) );
  NOR2_X1 U10121 ( .A1(n8624), .A2(n8623), .ZN(n8628) );
  OAI211_X1 U10122 ( .C1(n8628), .C2(n8627), .A(n8626), .B(n8625), .ZN(n8629)
         );
  INV_X1 U10123 ( .A(n8629), .ZN(n8630) );
  NOR2_X1 U10124 ( .A1(n8631), .A2(n8630), .ZN(n8636) );
  INV_X1 U10125 ( .A(n8632), .ZN(n8634) );
  OAI211_X1 U10126 ( .C1(n8636), .C2(n8635), .A(n8634), .B(n8633), .ZN(n8637)
         );
  NAND2_X1 U10127 ( .A1(n8638), .A2(n8637), .ZN(n8641) );
  NAND3_X1 U10128 ( .A1(n8641), .A2(n8640), .A3(n8639), .ZN(n8642) );
  NAND2_X1 U10129 ( .A1(n8644), .A2(n8642), .ZN(n8643) );
  MUX2_X1 U10130 ( .A(n8644), .B(n8643), .S(n9930), .Z(n8645) );
  INV_X1 U10131 ( .A(n8649), .ZN(n8651) );
  AOI21_X1 U10132 ( .B1(n8651), .B2(n8650), .A(n8655), .ZN(n8652) );
  OR2_X1 U10133 ( .A1(n8654), .A2(n8653), .ZN(n8658) );
  OAI21_X1 U10134 ( .B1(n6516), .B2(n8655), .A(P1_B_REG_SCAN_IN), .ZN(n8656)
         );
  INV_X1 U10135 ( .A(n8656), .ZN(n8657) );
  OAI21_X1 U10136 ( .B1(n8659), .B2(n8658), .A(n8657), .ZN(n8660) );
  OAI222_X1 U10137 ( .A1(n8665), .A2(n8664), .B1(n8663), .B2(P2_U3152), .C1(
        n8662), .C2(n8661), .ZN(P2_U3330) );
  NAND2_X1 U10138 ( .A1(n9161), .A2(n8846), .ZN(n8669) );
  NAND2_X1 U10139 ( .A1(n9076), .A2(n8671), .ZN(n8672) );
  OAI21_X1 U10140 ( .B1(n4468), .B2(n8807), .A(n8672), .ZN(n9057) );
  INV_X1 U10141 ( .A(n9018), .ZN(n9021) );
  AOI21_X1 U10142 ( .B1(n9135), .B2(n8997), .A(n9138), .ZN(n8981) );
  NAND2_X1 U10143 ( .A1(n8981), .A2(n8980), .ZN(n8979) );
  NAND2_X1 U10144 ( .A1(n8979), .A2(n8675), .ZN(n8963) );
  INV_X1 U10145 ( .A(n8965), .ZN(n8676) );
  AOI22_X2 U10146 ( .A1(n8963), .A2(n8676), .B1(n8758), .B2(n8954), .ZN(n8951)
         );
  INV_X1 U10148 ( .A(n9141), .ZN(n9033) );
  NAND2_X1 U10149 ( .A1(n9037), .A2(n9033), .ZN(n9026) );
  INV_X1 U10150 ( .A(n8678), .ZN(n9008) );
  NAND2_X1 U10151 ( .A1(n8983), .A2(n8758), .ZN(n8969) );
  INV_X1 U10152 ( .A(n8931), .ZN(n8679) );
  AOI21_X1 U10153 ( .B1(n9101), .B2(n8679), .A(n8918), .ZN(n9102) );
  AOI22_X1 U10154 ( .A1(n8680), .A2(n9060), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n9017), .ZN(n8681) );
  OAI21_X1 U10155 ( .B1(n8682), .B2(n9063), .A(n8681), .ZN(n8694) );
  XOR2_X1 U10156 ( .A(n8684), .B(n8683), .Z(n8692) );
  INV_X1 U10157 ( .A(n8685), .ZN(n8838) );
  NOR2_X1 U10158 ( .A1(n8687), .A2(n8686), .ZN(n8688) );
  NOR2_X1 U10159 ( .A1(n9053), .A2(n8688), .ZN(n8912) );
  NAND2_X1 U10160 ( .A1(n8838), .A2(n8912), .ZN(n8689) );
  AOI211_X1 U10161 ( .C1(n9102), .C2(n9074), .A(n8694), .B(n8693), .ZN(n8695)
         );
  OAI21_X1 U10162 ( .B1(n9106), .B2(n9094), .A(n8695), .ZN(P2_U3267) );
  INV_X1 U10163 ( .A(n7666), .ZN(n8697) );
  AOI21_X1 U10164 ( .B1(n6224), .B2(n8700), .A(n8697), .ZN(n8698) );
  OAI222_X1 U10165 ( .A1(n9053), .A2(n8699), .B1(n9051), .B2(n8696), .C1(n9049), .C2(n8698), .ZN(n10059) );
  XNOR2_X1 U10166 ( .A(n8701), .B(n8700), .ZN(n10061) );
  AOI22_X1 U10167 ( .A1(n10059), .A2(n9079), .B1(n9006), .B2(n10061), .ZN(
        n8708) );
  INV_X1 U10168 ( .A(n8702), .ZN(n8703) );
  OAI211_X1 U10169 ( .C1(n10058), .C2(n8704), .A(n8703), .B(n9181), .ZN(n10057) );
  OAI22_X1 U10170 ( .A1(n10057), .A2(n8916), .B1(n8705), .B2(n10025), .ZN(
        n8706) );
  AOI21_X1 U10171 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n9017), .A(n8706), .ZN(
        n8707) );
  OAI211_X1 U10172 ( .C1(n10058), .C2(n9063), .A(n8708), .B(n8707), .ZN(
        P2_U3294) );
  NAND2_X1 U10173 ( .A1(n8816), .A2(n8815), .ZN(n8814) );
  NAND2_X1 U10174 ( .A1(n8814), .A2(n8709), .ZN(n8712) );
  OAI211_X1 U10175 ( .C1(n8712), .C2(n8711), .A(n8710), .B(n10002), .ZN(n8718)
         );
  OAI22_X1 U10176 ( .A1(n8713), .A2(n9053), .B1(n8968), .B2(n9051), .ZN(n8946)
         );
  INV_X1 U10177 ( .A(n8946), .ZN(n8715) );
  OAI22_X1 U10178 ( .A1(n8715), .A2(n8800), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8714), .ZN(n8716) );
  AOI21_X1 U10179 ( .B1(n8941), .B2(n8789), .A(n8716), .ZN(n8717) );
  OAI211_X1 U10180 ( .C1(n8943), .C2(n10000), .A(n8718), .B(n8717), .ZN(
        P2_U3216) );
  XNOR2_X1 U10181 ( .A(n8720), .B(n8719), .ZN(n8721) );
  XNOR2_X1 U10182 ( .A(n8722), .B(n8721), .ZN(n8727) );
  AOI22_X1 U10183 ( .A1(n9998), .A2(n8844), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n8724) );
  NAND2_X1 U10184 ( .A1(n8821), .A2(n8843), .ZN(n8723) );
  OAI211_X1 U10185 ( .C1(n10006), .C2(n9009), .A(n8724), .B(n8723), .ZN(n8725)
         );
  AOI21_X1 U10186 ( .B1(n9135), .B2(n8834), .A(n8725), .ZN(n8726) );
  OAI21_X1 U10187 ( .B1(n8727), .B2(n8836), .A(n8726), .ZN(P2_U3218) );
  NAND2_X1 U10188 ( .A1(n8729), .A2(n8728), .ZN(n8731) );
  XOR2_X1 U10189 ( .A(n8731), .B(n8730), .Z(n8738) );
  NAND2_X1 U10190 ( .A1(n8846), .A2(n9070), .ZN(n8733) );
  NAND2_X1 U10191 ( .A1(n8845), .A2(n9068), .ZN(n8732) );
  NAND2_X1 U10192 ( .A1(n8733), .A2(n8732), .ZN(n9083) );
  AOI22_X1 U10193 ( .A1(n8734), .A2(n9083), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3152), .ZN(n8735) );
  OAI21_X1 U10194 ( .B1(n9077), .B2(n10006), .A(n8735), .ZN(n8736) );
  AOI21_X1 U10195 ( .B1(n9155), .B2(n8834), .A(n8736), .ZN(n8737) );
  OAI21_X1 U10196 ( .B1(n8738), .B2(n8836), .A(n8737), .ZN(P2_U3221) );
  NAND2_X1 U10197 ( .A1(n8739), .A2(n8785), .ZN(n8784) );
  NAND2_X1 U10198 ( .A1(n8784), .A2(n8740), .ZN(n8743) );
  AND2_X1 U10199 ( .A1(n8742), .A2(n8741), .ZN(n8792) );
  OAI211_X1 U10200 ( .C1(n8744), .C2(n8743), .A(n8792), .B(n10002), .ZN(n8749)
         );
  NOR2_X1 U10201 ( .A1(n10006), .A2(n9039), .ZN(n8747) );
  OAI22_X1 U10202 ( .A1(n9995), .A2(n9052), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8745), .ZN(n8746) );
  AOI211_X1 U10203 ( .C1(n9998), .C2(n8845), .A(n8747), .B(n8746), .ZN(n8748)
         );
  OAI211_X1 U10204 ( .C1(n9038), .C2(n10000), .A(n8749), .B(n8748), .ZN(
        P2_U3225) );
  NAND2_X1 U10205 ( .A1(n8751), .A2(n8750), .ZN(n8752) );
  NAND3_X1 U10206 ( .A1(n8753), .A2(n10002), .A3(n8752), .ZN(n8757) );
  AOI22_X1 U10207 ( .A1(n8842), .A2(n8821), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8754) );
  OAI21_X1 U10208 ( .B1(n9003), .B2(n8818), .A(n8754), .ZN(n8755) );
  AOI21_X1 U10209 ( .B1(n8972), .B2(n8789), .A(n8755), .ZN(n8756) );
  OAI211_X1 U10210 ( .C1(n8758), .C2(n10000), .A(n8757), .B(n8756), .ZN(
        P2_U3227) );
  NAND2_X1 U10211 ( .A1(n8760), .A2(n8759), .ZN(n8764) );
  XNOR2_X1 U10212 ( .A(n8761), .B(n8762), .ZN(n8826) );
  OAI22_X1 U10213 ( .A1(n8826), .A2(n8825), .B1(n8761), .B2(n8762), .ZN(n8763)
         );
  XOR2_X1 U10214 ( .A(n8764), .B(n8763), .Z(n8772) );
  OAI21_X1 U10215 ( .B1(n9995), .B2(n8766), .A(n8765), .ZN(n8767) );
  AOI21_X1 U10216 ( .B1(n9998), .B2(n8849), .A(n8767), .ZN(n8768) );
  OAI21_X1 U10217 ( .B1(n8769), .B2(n10006), .A(n8768), .ZN(n8770) );
  AOI21_X1 U10218 ( .B1(n9172), .B2(n8834), .A(n8770), .ZN(n8771) );
  OAI21_X1 U10219 ( .B1(n8772), .B2(n8836), .A(n8771), .ZN(P2_U3228) );
  XNOR2_X1 U10220 ( .A(n8775), .B(n8774), .ZN(n8776) );
  XNOR2_X1 U10221 ( .A(n8773), .B(n8776), .ZN(n8783) );
  OAI22_X1 U10222 ( .A1(n8818), .A2(n8778), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8777), .ZN(n8779) );
  AOI21_X1 U10223 ( .B1(n8821), .B2(n8988), .A(n8779), .ZN(n8780) );
  OAI21_X1 U10224 ( .B1(n8984), .B2(n10006), .A(n8780), .ZN(n8781) );
  AOI21_X1 U10225 ( .B1(n9127), .B2(n8834), .A(n8781), .ZN(n8782) );
  OAI21_X1 U10226 ( .B1(n8783), .B2(n8836), .A(n8782), .ZN(P2_U3231) );
  OAI211_X1 U10227 ( .C1(n8739), .C2(n8785), .A(n8784), .B(n10002), .ZN(n8791)
         );
  INV_X1 U10228 ( .A(n8786), .ZN(n9061) );
  AOI22_X1 U10229 ( .A1(n8821), .A2(n9069), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3152), .ZN(n8787) );
  OAI21_X1 U10230 ( .B1(n8807), .B2(n8818), .A(n8787), .ZN(n8788) );
  AOI21_X1 U10231 ( .B1(n9061), .B2(n8789), .A(n8788), .ZN(n8790) );
  OAI211_X1 U10232 ( .C1(n4467), .C2(n10000), .A(n8791), .B(n8790), .ZN(
        P2_U3235) );
  INV_X1 U10233 ( .A(n8792), .ZN(n8794) );
  NOR2_X1 U10234 ( .A1(n8794), .A2(n8793), .ZN(n8798) );
  XNOR2_X1 U10235 ( .A(n8796), .B(n8795), .ZN(n8797) );
  XNOR2_X1 U10236 ( .A(n8798), .B(n8797), .ZN(n8804) );
  NOR2_X1 U10237 ( .A1(n10006), .A2(n9029), .ZN(n8802) );
  AOI22_X1 U10238 ( .A1(n8997), .A2(n9068), .B1(n9070), .B2(n9069), .ZN(n9023)
         );
  OAI22_X1 U10239 ( .A1(n9023), .A2(n8800), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8799), .ZN(n8801) );
  AOI211_X1 U10240 ( .C1(n9141), .C2(n8834), .A(n8802), .B(n8801), .ZN(n8803)
         );
  OAI21_X1 U10241 ( .B1(n8804), .B2(n8836), .A(n8803), .ZN(P2_U3237) );
  XNOR2_X1 U10242 ( .A(n8805), .B(n8806), .ZN(n8813) );
  NAND2_X1 U10243 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8888) );
  OAI21_X1 U10244 ( .B1(n9995), .B2(n8807), .A(n8888), .ZN(n8808) );
  AOI21_X1 U10245 ( .B1(n9998), .B2(n8847), .A(n8808), .ZN(n8809) );
  OAI21_X1 U10246 ( .B1(n8810), .B2(n10006), .A(n8809), .ZN(n8811) );
  AOI21_X1 U10247 ( .B1(n9161), .B2(n8834), .A(n8811), .ZN(n8812) );
  OAI21_X1 U10248 ( .B1(n8813), .B2(n8836), .A(n8812), .ZN(P2_U3240) );
  INV_X1 U10249 ( .A(n9119), .ZN(n8824) );
  OAI211_X1 U10250 ( .C1(n8816), .C2(n8815), .A(n8814), .B(n10002), .ZN(n8823)
         );
  NOR2_X1 U10251 ( .A1(n8958), .A2(n10006), .ZN(n8820) );
  OAI22_X1 U10252 ( .A1(n8954), .A2(n8818), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8817), .ZN(n8819) );
  AOI211_X1 U10253 ( .C1(n8821), .C2(n8841), .A(n8820), .B(n8819), .ZN(n8822)
         );
  OAI211_X1 U10254 ( .C1(n8824), .C2(n10000), .A(n8823), .B(n8822), .ZN(
        P2_U3242) );
  XNOR2_X1 U10255 ( .A(n8826), .B(n8825), .ZN(n8837) );
  OAI22_X1 U10256 ( .A1(n9995), .A2(n8828), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8827), .ZN(n8829) );
  AOI21_X1 U10257 ( .B1(n9998), .B2(n8850), .A(n8829), .ZN(n8830) );
  OAI21_X1 U10258 ( .B1(n8831), .B2(n10006), .A(n8830), .ZN(n8832) );
  AOI21_X1 U10259 ( .B1(n8834), .B2(n8833), .A(n8832), .ZN(n8835) );
  OAI21_X1 U10260 ( .B1(n8837), .B2(n8836), .A(n8835), .ZN(P2_U3243) );
  MUX2_X1 U10261 ( .A(n8838), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8862), .Z(
        P2_U3582) );
  MUX2_X1 U10262 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8839), .S(P2_U3966), .Z(
        P2_U3581) );
  MUX2_X1 U10263 ( .A(n8840), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8862), .Z(
        P2_U3580) );
  MUX2_X1 U10264 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8841), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U10265 ( .A(n8842), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8862), .Z(
        P2_U3578) );
  MUX2_X1 U10266 ( .A(n8988), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8862), .Z(
        P2_U3577) );
  MUX2_X1 U10267 ( .A(n8843), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8862), .Z(
        P2_U3576) );
  MUX2_X1 U10268 ( .A(n8997), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8862), .Z(
        P2_U3575) );
  MUX2_X1 U10269 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8844), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U10270 ( .A(n9069), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8862), .Z(
        P2_U3573) );
  MUX2_X1 U10271 ( .A(n8845), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8862), .Z(
        P2_U3572) );
  MUX2_X1 U10272 ( .A(n9071), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8862), .Z(
        P2_U3571) );
  MUX2_X1 U10273 ( .A(n8846), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8862), .Z(
        P2_U3570) );
  MUX2_X1 U10274 ( .A(n8847), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8862), .Z(
        P2_U3569) );
  MUX2_X1 U10275 ( .A(n8848), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8862), .Z(
        P2_U3568) );
  MUX2_X1 U10276 ( .A(n8849), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8862), .Z(
        P2_U3567) );
  MUX2_X1 U10277 ( .A(n8850), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8862), .Z(
        P2_U3566) );
  MUX2_X1 U10278 ( .A(n8851), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8862), .Z(
        P2_U3565) );
  MUX2_X1 U10279 ( .A(n8852), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8862), .Z(
        P2_U3564) );
  MUX2_X1 U10280 ( .A(n8853), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8862), .Z(
        P2_U3563) );
  MUX2_X1 U10281 ( .A(n8854), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8862), .Z(
        P2_U3562) );
  MUX2_X1 U10282 ( .A(n8855), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8862), .Z(
        P2_U3561) );
  MUX2_X1 U10283 ( .A(n8856), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8862), .Z(
        P2_U3560) );
  MUX2_X1 U10284 ( .A(n9997), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8862), .Z(
        P2_U3559) );
  MUX2_X1 U10285 ( .A(n8857), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8862), .Z(
        P2_U3558) );
  MUX2_X1 U10286 ( .A(n8858), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8862), .Z(
        P2_U3557) );
  MUX2_X1 U10287 ( .A(n8859), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8862), .Z(
        P2_U3556) );
  MUX2_X1 U10288 ( .A(n8860), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8862), .Z(
        P2_U3555) );
  MUX2_X1 U10289 ( .A(n6115), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8862), .Z(
        P2_U3554) );
  MUX2_X1 U10290 ( .A(n8861), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8862), .Z(
        P2_U3553) );
  MUX2_X1 U10291 ( .A(n8863), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8862), .Z(
        P2_U3552) );
  INV_X1 U10292 ( .A(n8864), .ZN(n8867) );
  NOR2_X1 U10293 ( .A1(n10009), .A2(n8865), .ZN(n8866) );
  AOI211_X1 U10294 ( .C1(n10013), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n8867), .B(
        n8866), .ZN(n8878) );
  OAI211_X1 U10295 ( .C1(n8870), .C2(n8869), .A(n10007), .B(n8868), .ZN(n8877)
         );
  INV_X1 U10296 ( .A(n8871), .ZN(n8875) );
  INV_X1 U10297 ( .A(n8872), .ZN(n8874) );
  OAI211_X1 U10298 ( .C1(n8875), .C2(n8874), .A(n8873), .B(n10008), .ZN(n8876)
         );
  NAND3_X1 U10299 ( .A1(n8878), .A2(n8877), .A3(n8876), .ZN(P2_U3255) );
  OAI21_X1 U10300 ( .B1(n8881), .B2(n8880), .A(n8879), .ZN(n8883) );
  AOI22_X1 U10301 ( .A1(n8890), .A2(n8899), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n8900), .ZN(n8882) );
  NOR2_X1 U10302 ( .A1(n8883), .A2(n8882), .ZN(n8898) );
  AOI21_X1 U10303 ( .B1(n8883), .B2(n8882), .A(n8898), .ZN(n8893) );
  NAND2_X1 U10304 ( .A1(n8886), .A2(n8302), .ZN(n8896) );
  OAI21_X1 U10305 ( .B1(n8886), .B2(n8302), .A(n8896), .ZN(n8887) );
  NAND2_X1 U10306 ( .A1(n8887), .A2(n10008), .ZN(n8892) );
  OAI21_X1 U10307 ( .B1(n9714), .B2(n10156), .A(n8888), .ZN(n8889) );
  AOI21_X1 U10308 ( .B1(n9731), .B2(n8890), .A(n8889), .ZN(n8891) );
  OAI211_X1 U10309 ( .C1(n8893), .C2(n10011), .A(n8892), .B(n8891), .ZN(
        P2_U3263) );
  NAND2_X1 U10310 ( .A1(n8894), .A2(n8900), .ZN(n8895) );
  NAND2_X1 U10311 ( .A1(n8896), .A2(n8895), .ZN(n8897) );
  XNOR2_X1 U10312 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8897), .ZN(n8905) );
  INV_X1 U10313 ( .A(n8905), .ZN(n8903) );
  AOI21_X1 U10314 ( .B1(n8900), .B2(n8899), .A(n8898), .ZN(n8901) );
  XOR2_X1 U10315 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8901), .Z(n8904) );
  OAI21_X1 U10316 ( .B1(n8904), .B2(n10011), .A(n10009), .ZN(n8902) );
  AOI21_X1 U10317 ( .B1(n8903), .B2(n10008), .A(n8902), .ZN(n8907) );
  AOI22_X1 U10318 ( .A1(n8905), .A2(n10008), .B1(n10007), .B2(n8904), .ZN(
        n8906) );
  MUX2_X1 U10319 ( .A(n8907), .B(n8906), .S(n10027), .Z(n8909) );
  NAND2_X1 U10320 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3152), .ZN(n8908) );
  OAI211_X1 U10321 ( .C1(n8910), .C2(n9714), .A(n8909), .B(n8908), .ZN(
        P2_U3264) );
  XNOR2_X1 U10322 ( .A(n8917), .B(n9096), .ZN(n8911) );
  NAND2_X1 U10323 ( .A1(n8911), .A2(n9181), .ZN(n9095) );
  NAND2_X1 U10324 ( .A1(n8913), .A2(n8912), .ZN(n9099) );
  NOR2_X1 U10325 ( .A1(n9017), .A2(n9099), .ZN(n8921) );
  NOR2_X1 U10326 ( .A1(n9096), .A2(n9063), .ZN(n8914) );
  AOI211_X1 U10327 ( .C1(n9017), .C2(P2_REG2_REG_31__SCAN_IN), .A(n8921), .B(
        n8914), .ZN(n8915) );
  OAI21_X1 U10328 ( .B1(n9095), .B2(n8916), .A(n8915), .ZN(P2_U3265) );
  OAI21_X1 U10329 ( .B1(n8919), .B2(n8918), .A(n8917), .ZN(n9100) );
  NOR2_X1 U10330 ( .A1(n8919), .A2(n9063), .ZN(n8920) );
  AOI211_X1 U10331 ( .C1(n9017), .C2(P2_REG2_REG_30__SCAN_IN), .A(n8921), .B(
        n8920), .ZN(n8922) );
  OAI21_X1 U10332 ( .B1(n8923), .B2(n9100), .A(n8922), .ZN(P2_U3266) );
  XNOR2_X1 U10333 ( .A(n8925), .B(n8924), .ZN(n9111) );
  NAND2_X1 U10334 ( .A1(n4881), .A2(n8926), .ZN(n8928) );
  XNOR2_X1 U10335 ( .A(n8928), .B(n8927), .ZN(n8930) );
  OAI21_X1 U10336 ( .B1(n8930), .B2(n9049), .A(n8929), .ZN(n9107) );
  AOI211_X1 U10337 ( .C1(n9109), .C2(n8938), .A(n10097), .B(n8931), .ZN(n9108)
         );
  NAND2_X1 U10338 ( .A1(n9108), .A2(n9043), .ZN(n8934) );
  AOI22_X1 U10339 ( .A1(n8932), .A2(n9060), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n9017), .ZN(n8933) );
  OAI211_X1 U10340 ( .C1(n4474), .C2(n9063), .A(n8934), .B(n8933), .ZN(n8935)
         );
  AOI21_X1 U10341 ( .B1(n9107), .B2(n9079), .A(n8935), .ZN(n8936) );
  OAI21_X1 U10342 ( .B1(n9111), .B2(n9094), .A(n8936), .ZN(P2_U3268) );
  XOR2_X1 U10343 ( .A(n8944), .B(n8937), .Z(n9116) );
  INV_X1 U10344 ( .A(n8938), .ZN(n8939) );
  AOI211_X1 U10345 ( .C1(n9113), .C2(n8940), .A(n10097), .B(n8939), .ZN(n9112)
         );
  AOI22_X1 U10346 ( .A1(n8941), .A2(n9060), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n9017), .ZN(n8942) );
  OAI21_X1 U10347 ( .B1(n8943), .B2(n9063), .A(n8942), .ZN(n8949) );
  AOI21_X1 U10348 ( .B1(n8945), .B2(n8944), .A(n9049), .ZN(n8947) );
  AOI21_X1 U10349 ( .B1(n8947), .B2(n4881), .A(n8946), .ZN(n9115) );
  NOR2_X1 U10350 ( .A1(n9115), .A2(n9017), .ZN(n8948) );
  AOI211_X1 U10351 ( .C1(n9043), .C2(n9112), .A(n8949), .B(n8948), .ZN(n8950)
         );
  OAI21_X1 U10352 ( .B1(n9116), .B2(n9094), .A(n8950), .ZN(P2_U3269) );
  XOR2_X1 U10353 ( .A(n8953), .B(n8951), .Z(n9121) );
  AOI22_X1 U10354 ( .A1(n9119), .A2(n9092), .B1(n9017), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8962) );
  XOR2_X1 U10355 ( .A(n8952), .B(n8953), .Z(n8955) );
  OAI222_X1 U10356 ( .A1(n9053), .A2(n8956), .B1(n8955), .B2(n9049), .C1(n9051), .C2(n8954), .ZN(n9117) );
  AOI211_X1 U10357 ( .C1(n9119), .C2(n8969), .A(n10097), .B(n8957), .ZN(n9118)
         );
  INV_X1 U10358 ( .A(n9118), .ZN(n8959) );
  OAI22_X1 U10359 ( .A1(n8959), .A2(n8974), .B1(n10025), .B2(n8958), .ZN(n8960) );
  OAI21_X1 U10360 ( .B1(n9117), .B2(n8960), .A(n9079), .ZN(n8961) );
  OAI211_X1 U10361 ( .C1(n9121), .C2(n9094), .A(n8962), .B(n8961), .ZN(
        P2_U3270) );
  XNOR2_X1 U10362 ( .A(n8963), .B(n8965), .ZN(n9126) );
  AOI22_X1 U10363 ( .A1(n9124), .A2(n9092), .B1(n9017), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n8978) );
  NAND2_X1 U10364 ( .A1(n8989), .A2(n8964), .ZN(n8966) );
  XNOR2_X1 U10365 ( .A(n8966), .B(n8965), .ZN(n8967) );
  OAI222_X1 U10366 ( .A1(n9053), .A2(n8968), .B1(n9051), .B2(n9003), .C1(n9049), .C2(n8967), .ZN(n9122) );
  INV_X1 U10367 ( .A(n8983), .ZN(n8971) );
  INV_X1 U10368 ( .A(n8969), .ZN(n8970) );
  AOI211_X1 U10369 ( .C1(n9124), .C2(n8971), .A(n10097), .B(n8970), .ZN(n9123)
         );
  INV_X1 U10370 ( .A(n9123), .ZN(n8975) );
  INV_X1 U10371 ( .A(n8972), .ZN(n8973) );
  OAI22_X1 U10372 ( .A1(n8975), .A2(n8974), .B1(n10025), .B2(n8973), .ZN(n8976) );
  OAI21_X1 U10373 ( .B1(n9122), .B2(n8976), .A(n9079), .ZN(n8977) );
  OAI211_X1 U10374 ( .C1(n9126), .C2(n9094), .A(n8978), .B(n8977), .ZN(
        P2_U3271) );
  OAI21_X1 U10375 ( .B1(n8981), .B2(n8980), .A(n8979), .ZN(n8982) );
  INV_X1 U10376 ( .A(n8982), .ZN(n9131) );
  AOI21_X1 U10377 ( .B1(n9127), .B2(n9008), .A(n8983), .ZN(n9128) );
  INV_X1 U10378 ( .A(n9127), .ZN(n8987) );
  INV_X1 U10379 ( .A(n8984), .ZN(n8985) );
  AOI22_X1 U10380 ( .A1(n9017), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8985), .B2(
        n9060), .ZN(n8986) );
  OAI21_X1 U10381 ( .B1(n8987), .B2(n9063), .A(n8986), .ZN(n8999) );
  AND2_X1 U10382 ( .A1(n8988), .A2(n9068), .ZN(n8996) );
  INV_X1 U10383 ( .A(n8989), .ZN(n8994) );
  AOI21_X1 U10384 ( .B1(n8992), .B2(n8991), .A(n8990), .ZN(n8993) );
  NOR3_X1 U10385 ( .A1(n8994), .A2(n8993), .A3(n9049), .ZN(n8995) );
  AOI211_X1 U10386 ( .C1(n9070), .C2(n8997), .A(n8996), .B(n8995), .ZN(n9130)
         );
  NOR2_X1 U10387 ( .A1(n9130), .A2(n9017), .ZN(n8998) );
  AOI211_X1 U10388 ( .C1(n9128), .C2(n9074), .A(n8999), .B(n8998), .ZN(n9000)
         );
  OAI21_X1 U10389 ( .B1(n9131), .B2(n9094), .A(n9000), .ZN(P2_U3272) );
  XNOR2_X1 U10390 ( .A(n9001), .B(n9004), .ZN(n9002) );
  OAI222_X1 U10391 ( .A1(n9053), .A2(n9003), .B1(n9051), .B2(n9052), .C1(n9049), .C2(n9002), .ZN(n9133) );
  INV_X1 U10392 ( .A(n9133), .ZN(n9016) );
  INV_X1 U10393 ( .A(n9138), .ZN(n9007) );
  NAND2_X1 U10394 ( .A1(n9005), .A2(n9004), .ZN(n9132) );
  NAND3_X1 U10395 ( .A1(n9007), .A2(n9006), .A3(n9132), .ZN(n9015) );
  AOI211_X1 U10396 ( .C1(n9135), .C2(n9026), .A(n10097), .B(n8678), .ZN(n9134)
         );
  INV_X1 U10397 ( .A(n9135), .ZN(n9012) );
  INV_X1 U10398 ( .A(n9009), .ZN(n9010) );
  AOI22_X1 U10399 ( .A1(n9017), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n9010), .B2(
        n9060), .ZN(n9011) );
  OAI21_X1 U10400 ( .B1(n9012), .B2(n9063), .A(n9011), .ZN(n9013) );
  AOI21_X1 U10401 ( .B1(n9134), .B2(n9043), .A(n9013), .ZN(n9014) );
  OAI211_X1 U10402 ( .C1(n9017), .C2(n9016), .A(n9015), .B(n9014), .ZN(
        P2_U3273) );
  XNOR2_X1 U10403 ( .A(n9019), .B(n9018), .ZN(n9143) );
  NAND2_X1 U10404 ( .A1(n9020), .A2(n9084), .ZN(n9025) );
  AOI21_X1 U10405 ( .B1(n9044), .B2(n9022), .A(n9021), .ZN(n9024) );
  OAI21_X1 U10406 ( .B1(n9025), .B2(n9024), .A(n9023), .ZN(n9139) );
  INV_X1 U10407 ( .A(n9037), .ZN(n9028) );
  INV_X1 U10408 ( .A(n9026), .ZN(n9027) );
  AOI211_X1 U10409 ( .C1(n9141), .C2(n9028), .A(n10097), .B(n9027), .ZN(n9140)
         );
  NAND2_X1 U10410 ( .A1(n9140), .A2(n9043), .ZN(n9032) );
  INV_X1 U10411 ( .A(n9029), .ZN(n9030) );
  AOI22_X1 U10412 ( .A1(n9017), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9030), .B2(
        n9060), .ZN(n9031) );
  OAI211_X1 U10413 ( .C1(n9033), .C2(n9063), .A(n9032), .B(n9031), .ZN(n9034)
         );
  AOI21_X1 U10414 ( .B1(n9139), .B2(n9079), .A(n9034), .ZN(n9035) );
  OAI21_X1 U10415 ( .B1(n9143), .B2(n9094), .A(n9035), .ZN(P2_U3274) );
  XOR2_X1 U10416 ( .A(n9036), .B(n9047), .Z(n9148) );
  AOI211_X1 U10417 ( .C1(n9146), .C2(n9058), .A(n10097), .B(n9037), .ZN(n9145)
         );
  NOR2_X1 U10418 ( .A1(n9038), .A2(n9063), .ZN(n9042) );
  OAI22_X1 U10419 ( .A1(n9079), .A2(n9040), .B1(n9039), .B2(n10025), .ZN(n9041) );
  AOI211_X1 U10420 ( .C1(n9145), .C2(n9043), .A(n9042), .B(n9041), .ZN(n9055)
         );
  INV_X1 U10421 ( .A(n9044), .ZN(n9045) );
  AOI21_X1 U10422 ( .B1(n9047), .B2(n9046), .A(n9045), .ZN(n9048) );
  OAI222_X1 U10423 ( .A1(n9053), .A2(n9052), .B1(n9051), .B2(n9050), .C1(n9049), .C2(n9048), .ZN(n9144) );
  NAND2_X1 U10424 ( .A1(n9144), .A2(n9079), .ZN(n9054) );
  OAI211_X1 U10425 ( .C1(n9148), .C2(n9094), .A(n9055), .B(n9054), .ZN(
        P2_U3275) );
  XNOR2_X1 U10426 ( .A(n9057), .B(n9056), .ZN(n9153) );
  INV_X1 U10427 ( .A(n9058), .ZN(n9059) );
  AOI21_X1 U10428 ( .B1(n9149), .B2(n9086), .A(n9059), .ZN(n9150) );
  AOI22_X1 U10429 ( .A1(n9017), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9061), .B2(
        n9060), .ZN(n9062) );
  OAI21_X1 U10430 ( .B1(n4467), .B2(n9063), .A(n9062), .ZN(n9073) );
  NAND2_X1 U10431 ( .A1(n9080), .A2(n9064), .ZN(n9066) );
  XNOR2_X1 U10432 ( .A(n9066), .B(n9065), .ZN(n9067) );
  AOI222_X1 U10433 ( .A1(n9071), .A2(n9070), .B1(n9069), .B2(n9068), .C1(n9084), .C2(n9067), .ZN(n9152) );
  NOR2_X1 U10434 ( .A1(n9152), .A2(n9017), .ZN(n9072) );
  AOI211_X1 U10435 ( .C1(n9150), .C2(n9074), .A(n9073), .B(n9072), .ZN(n9075)
         );
  OAI21_X1 U10436 ( .B1(n9094), .B2(n9153), .A(n9075), .ZN(P2_U3276) );
  XOR2_X1 U10437 ( .A(n9076), .B(n9082), .Z(n9158) );
  OAI22_X1 U10438 ( .A1(n9079), .A2(n9078), .B1(n9077), .B2(n10025), .ZN(n9091) );
  OAI21_X1 U10439 ( .B1(n9082), .B2(n9081), .A(n9080), .ZN(n9085) );
  AOI21_X1 U10440 ( .B1(n9085), .B2(n9084), .A(n9083), .ZN(n9157) );
  INV_X1 U10441 ( .A(n9086), .ZN(n9087) );
  AOI211_X1 U10442 ( .C1(n9155), .C2(n9088), .A(n10097), .B(n9087), .ZN(n9154)
         );
  NAND2_X1 U10443 ( .A1(n9154), .A2(n10027), .ZN(n9089) );
  AOI21_X1 U10444 ( .B1(n9157), .B2(n9089), .A(n9017), .ZN(n9090) );
  AOI211_X1 U10445 ( .C1(n9092), .C2(n9155), .A(n9091), .B(n9090), .ZN(n9093)
         );
  OAI21_X1 U10446 ( .B1(n9158), .B2(n9094), .A(n9093), .ZN(P2_U3277) );
  OAI211_X1 U10447 ( .C1(n9096), .C2(n10095), .A(n9095), .B(n9099), .ZN(n9186)
         );
  MUX2_X1 U10448 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9186), .S(n10119), .Z(
        P2_U3551) );
  NAND2_X1 U10449 ( .A1(n9097), .A2(n9180), .ZN(n9098) );
  OAI211_X1 U10450 ( .C1(n9100), .C2(n10097), .A(n9099), .B(n9098), .ZN(n9187)
         );
  MUX2_X1 U10451 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9187), .S(n10119), .Z(
        P2_U3550) );
  AOI22_X1 U10452 ( .A1(n9102), .A2(n9181), .B1(n9180), .B2(n9101), .ZN(n9104)
         );
  OAI21_X1 U10453 ( .B1(n9106), .B2(n9170), .A(n9105), .ZN(n9188) );
  MUX2_X1 U10454 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n9188), .S(n10119), .Z(
        P2_U3549) );
  AOI211_X1 U10455 ( .C1(n9180), .C2(n9109), .A(n9108), .B(n9107), .ZN(n9110)
         );
  OAI21_X1 U10456 ( .B1(n9111), .B2(n9170), .A(n9110), .ZN(n9189) );
  MUX2_X1 U10457 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9189), .S(n10119), .Z(
        P2_U3548) );
  AOI21_X1 U10458 ( .B1(n9180), .B2(n9113), .A(n9112), .ZN(n9114) );
  OAI211_X1 U10459 ( .C1(n9116), .C2(n9170), .A(n9115), .B(n9114), .ZN(n9190)
         );
  MUX2_X1 U10460 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9190), .S(n10119), .Z(
        P2_U3547) );
  AOI211_X1 U10461 ( .C1(n9180), .C2(n9119), .A(n9118), .B(n9117), .ZN(n9120)
         );
  OAI21_X1 U10462 ( .B1(n9121), .B2(n9170), .A(n9120), .ZN(n9191) );
  MUX2_X1 U10463 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9191), .S(n10119), .Z(
        P2_U3546) );
  AOI211_X1 U10464 ( .C1(n9180), .C2(n9124), .A(n9123), .B(n9122), .ZN(n9125)
         );
  OAI21_X1 U10465 ( .B1(n9126), .B2(n9170), .A(n9125), .ZN(n9192) );
  MUX2_X1 U10466 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9192), .S(n10119), .Z(
        P2_U3545) );
  AOI22_X1 U10467 ( .A1(n9128), .A2(n9181), .B1(n9180), .B2(n9127), .ZN(n9129)
         );
  OAI211_X1 U10468 ( .C1(n9131), .C2(n9170), .A(n9130), .B(n9129), .ZN(n9193)
         );
  MUX2_X1 U10469 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9193), .S(n10119), .Z(
        P2_U3544) );
  NAND2_X1 U10470 ( .A1(n9132), .A2(n10101), .ZN(n9137) );
  AOI211_X1 U10471 ( .C1(n9180), .C2(n9135), .A(n9134), .B(n9133), .ZN(n9136)
         );
  OAI21_X1 U10472 ( .B1(n9138), .B2(n9137), .A(n9136), .ZN(n9194) );
  MUX2_X1 U10473 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9194), .S(n10119), .Z(
        P2_U3543) );
  AOI211_X1 U10474 ( .C1(n9180), .C2(n9141), .A(n9140), .B(n9139), .ZN(n9142)
         );
  OAI21_X1 U10475 ( .B1(n9143), .B2(n9170), .A(n9142), .ZN(n9195) );
  MUX2_X1 U10476 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9195), .S(n10119), .Z(
        P2_U3542) );
  AOI211_X1 U10477 ( .C1(n9180), .C2(n9146), .A(n9145), .B(n9144), .ZN(n9147)
         );
  OAI21_X1 U10478 ( .B1(n9148), .B2(n9170), .A(n9147), .ZN(n9196) );
  MUX2_X1 U10479 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9196), .S(n10119), .Z(
        P2_U3541) );
  AOI22_X1 U10480 ( .A1(n9150), .A2(n9181), .B1(n9180), .B2(n9149), .ZN(n9151)
         );
  OAI211_X1 U10481 ( .C1(n9153), .C2(n9170), .A(n9152), .B(n9151), .ZN(n9197)
         );
  MUX2_X1 U10482 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9197), .S(n10119), .Z(
        P2_U3540) );
  AOI21_X1 U10483 ( .B1(n9180), .B2(n9155), .A(n9154), .ZN(n9156) );
  OAI211_X1 U10484 ( .C1(n9158), .C2(n9170), .A(n9157), .B(n9156), .ZN(n9198)
         );
  MUX2_X1 U10485 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9198), .S(n10119), .Z(
        P2_U3539) );
  AOI211_X1 U10486 ( .C1(n9180), .C2(n9161), .A(n9160), .B(n9159), .ZN(n9162)
         );
  OAI21_X1 U10487 ( .B1(n9170), .B2(n9163), .A(n9162), .ZN(n9199) );
  MUX2_X1 U10488 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9199), .S(n10119), .Z(
        P2_U3538) );
  INV_X1 U10489 ( .A(n9164), .ZN(n9169) );
  AOI211_X1 U10490 ( .C1(n9180), .C2(n9167), .A(n9166), .B(n9165), .ZN(n9168)
         );
  OAI21_X1 U10491 ( .B1(n9170), .B2(n9169), .A(n9168), .ZN(n9200) );
  MUX2_X1 U10492 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9200), .S(n10119), .Z(
        P2_U3537) );
  INV_X1 U10493 ( .A(n9171), .ZN(n9178) );
  INV_X1 U10494 ( .A(n9172), .ZN(n9173) );
  OAI22_X1 U10495 ( .A1(n9174), .A2(n10097), .B1(n9173), .B2(n10095), .ZN(
        n9175) );
  INV_X1 U10496 ( .A(n9175), .ZN(n9176) );
  OAI211_X1 U10497 ( .C1(n9178), .C2(n10087), .A(n9177), .B(n9176), .ZN(n9201)
         );
  MUX2_X1 U10498 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9201), .S(n10119), .Z(
        P2_U3536) );
  AOI22_X1 U10499 ( .A1(n9182), .A2(n9181), .B1(n9180), .B2(n9179), .ZN(n9183)
         );
  OAI211_X1 U10500 ( .C1(n10087), .C2(n9185), .A(n9184), .B(n9183), .ZN(n9202)
         );
  MUX2_X1 U10501 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n9202), .S(n10119), .Z(
        P2_U3533) );
  MUX2_X1 U10502 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9186), .S(n10105), .Z(
        P2_U3519) );
  MUX2_X1 U10503 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n9187), .S(n10105), .Z(
        P2_U3518) );
  MUX2_X1 U10504 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n9188), .S(n10105), .Z(
        P2_U3517) );
  MUX2_X1 U10505 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9189), .S(n10105), .Z(
        P2_U3516) );
  MUX2_X1 U10506 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9190), .S(n10105), .Z(
        P2_U3515) );
  MUX2_X1 U10507 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9191), .S(n10105), .Z(
        P2_U3514) );
  MUX2_X1 U10508 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9192), .S(n10105), .Z(
        P2_U3513) );
  MUX2_X1 U10509 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9193), .S(n10105), .Z(
        P2_U3512) );
  MUX2_X1 U10510 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9194), .S(n10105), .Z(
        P2_U3511) );
  MUX2_X1 U10511 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9195), .S(n10105), .Z(
        P2_U3510) );
  MUX2_X1 U10512 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9196), .S(n10105), .Z(
        P2_U3509) );
  MUX2_X1 U10513 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9197), .S(n10105), .Z(
        P2_U3508) );
  MUX2_X1 U10514 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9198), .S(n10105), .Z(
        P2_U3507) );
  MUX2_X1 U10515 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9199), .S(n10105), .Z(
        P2_U3505) );
  MUX2_X1 U10516 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9200), .S(n10105), .Z(
        P2_U3502) );
  MUX2_X1 U10517 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9201), .S(n10105), .Z(
        P2_U3499) );
  MUX2_X1 U10518 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n9202), .S(n10105), .Z(
        P2_U3490) );
  INV_X1 U10519 ( .A(n9203), .ZN(n9700) );
  NOR4_X1 U10520 ( .A1(n5553), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3152), .A4(
        n5554), .ZN(n9204) );
  AOI21_X1 U10521 ( .B1(n9210), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9204), .ZN(
        n9205) );
  OAI21_X1 U10522 ( .B1(n9700), .B2(n9212), .A(n9205), .ZN(P2_U3327) );
  INV_X1 U10523 ( .A(n9206), .ZN(n9702) );
  AOI22_X1 U10524 ( .A1(n9207), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n9210), .ZN(n9208) );
  OAI21_X1 U10525 ( .B1(n9702), .B2(n9212), .A(n9208), .ZN(P2_U3328) );
  INV_X1 U10526 ( .A(n9209), .ZN(n9706) );
  AOI22_X1 U10527 ( .A1(n4613), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n9210), .ZN(n9211) );
  OAI21_X1 U10528 ( .B1(n9706), .B2(n9212), .A(n9211), .ZN(P2_U3329) );
  INV_X1 U10529 ( .A(n9213), .ZN(n9214) );
  MUX2_X1 U10530 ( .A(n9214), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  NAND2_X1 U10531 ( .A1(n4369), .A2(n9215), .ZN(n9217) );
  XNOR2_X1 U10532 ( .A(n9217), .B(n9216), .ZN(n9223) );
  OAI22_X1 U10533 ( .A1(n9325), .A2(n9491), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9218), .ZN(n9220) );
  NOR2_X1 U10534 ( .A1(n9326), .A2(n9522), .ZN(n9219) );
  AOI211_X1 U10535 ( .C1(n9495), .C2(n9329), .A(n9220), .B(n9219), .ZN(n9222)
         );
  NAND2_X1 U10536 ( .A1(n9624), .A2(n9313), .ZN(n9221) );
  OAI211_X1 U10537 ( .C1(n9223), .C2(n9315), .A(n9222), .B(n9221), .ZN(
        P1_U3214) );
  NOR3_X1 U10538 ( .A1(n9226), .A2(n4675), .A3(n9225), .ZN(n9229) );
  INV_X1 U10539 ( .A(n9227), .ZN(n9228) );
  OAI21_X1 U10540 ( .B1(n9229), .B2(n9228), .A(n9322), .ZN(n9234) );
  AOI22_X1 U10541 ( .A1(n9357), .A2(n9308), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        P1_U3084), .ZN(n9233) );
  AOI22_X1 U10542 ( .A1(n9313), .A2(n9230), .B1(n9264), .B2(n9355), .ZN(n9232)
         );
  NAND2_X1 U10543 ( .A1(n9329), .A2(n5101), .ZN(n9231) );
  NAND4_X1 U10544 ( .A1(n9234), .A2(n9233), .A3(n9232), .A4(n9231), .ZN(
        P1_U3216) );
  OAI21_X1 U10545 ( .B1(n9236), .B2(n4340), .A(n9279), .ZN(n9237) );
  NAND2_X1 U10546 ( .A1(n9237), .A2(n9322), .ZN(n9241) );
  NOR2_X1 U10547 ( .A1(n9311), .A2(n9554), .ZN(n9239) );
  NAND2_X1 U10548 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9401) );
  OAI21_X1 U10549 ( .B1(n9549), .B2(n9325), .A(n9401), .ZN(n9238) );
  AOI211_X1 U10550 ( .C1(n9308), .C2(n9577), .A(n9239), .B(n9238), .ZN(n9240)
         );
  OAI211_X1 U10551 ( .C1(n9558), .C2(n9332), .A(n9241), .B(n9240), .ZN(
        P1_U3217) );
  OAI21_X1 U10552 ( .B1(n9244), .B2(n9243), .A(n9242), .ZN(n9245) );
  NAND2_X1 U10553 ( .A1(n9245), .A2(n9322), .ZN(n9250) );
  NOR2_X1 U10554 ( .A1(n9311), .A2(n9524), .ZN(n9248) );
  OAI22_X1 U10555 ( .A1(n9549), .A2(n9326), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9246), .ZN(n9247) );
  AOI211_X1 U10556 ( .C1(n9264), .C2(n9340), .A(n9248), .B(n9247), .ZN(n9249)
         );
  OAI211_X1 U10557 ( .C1(n4525), .C2(n9332), .A(n9250), .B(n9249), .ZN(
        P1_U3221) );
  AOI21_X1 U10558 ( .B1(n9253), .B2(n9252), .A(n9320), .ZN(n9259) );
  OAI22_X1 U10559 ( .A1(n9325), .A2(n9465), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9254), .ZN(n9256) );
  NOR2_X1 U10560 ( .A1(n9326), .A2(n9491), .ZN(n9255) );
  AOI211_X1 U10561 ( .C1(n9461), .C2(n9329), .A(n9256), .B(n9255), .ZN(n9258)
         );
  NAND2_X1 U10562 ( .A1(n9612), .A2(n9313), .ZN(n9257) );
  OAI211_X1 U10563 ( .C1(n9259), .C2(n9315), .A(n9258), .B(n9257), .ZN(
        P1_U3223) );
  INV_X1 U10564 ( .A(n9261), .ZN(n9262) );
  AOI21_X1 U10565 ( .B1(n9263), .B2(n9260), .A(n9262), .ZN(n9269) );
  NOR2_X1 U10566 ( .A1(n9311), .A2(n9565), .ZN(n9267) );
  NAND2_X1 U10567 ( .A1(n9577), .A2(n9264), .ZN(n9265) );
  NAND2_X1 U10568 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9907) );
  OAI211_X1 U10569 ( .C1(n9570), .C2(n9326), .A(n9265), .B(n9907), .ZN(n9266)
         );
  AOI211_X1 U10570 ( .C1(n9654), .C2(n9313), .A(n9267), .B(n9266), .ZN(n9268)
         );
  OAI21_X1 U10571 ( .B1(n9269), .B2(n9315), .A(n9268), .ZN(P1_U3226) );
  AOI21_X1 U10572 ( .B1(n9272), .B2(n9271), .A(n9270), .ZN(n9278) );
  OAI22_X1 U10573 ( .A1(n9325), .A2(n9477), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9273), .ZN(n9275) );
  NOR2_X1 U10574 ( .A1(n9326), .A2(n9505), .ZN(n9274) );
  AOI211_X1 U10575 ( .C1(n9481), .C2(n9329), .A(n9275), .B(n9274), .ZN(n9277)
         );
  NAND2_X1 U10576 ( .A1(n9619), .A2(n9313), .ZN(n9276) );
  OAI211_X1 U10577 ( .C1(n9278), .C2(n9315), .A(n9277), .B(n9276), .ZN(
        P1_U3227) );
  INV_X1 U10578 ( .A(n9279), .ZN(n9283) );
  INV_X1 U10579 ( .A(n9280), .ZN(n9282) );
  NOR3_X1 U10580 ( .A1(n9283), .A2(n9282), .A3(n9281), .ZN(n9286) );
  INV_X1 U10581 ( .A(n9284), .ZN(n9285) );
  OAI21_X1 U10582 ( .B1(n9286), .B2(n9285), .A(n9322), .ZN(n9290) );
  AOI22_X1 U10583 ( .A1(n9343), .A2(n9308), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n9287) );
  OAI21_X1 U10584 ( .B1(n9538), .B2(n9325), .A(n9287), .ZN(n9288) );
  AOI21_X1 U10585 ( .B1(n9533), .B2(n9329), .A(n9288), .ZN(n9289) );
  OAI211_X1 U10586 ( .C1(n9535), .C2(n9332), .A(n9290), .B(n9289), .ZN(
        P1_U3231) );
  INV_X1 U10587 ( .A(n9294), .ZN(n9297) );
  AOI21_X1 U10588 ( .B1(n9294), .B2(n9293), .A(n9292), .ZN(n9295) );
  NOR2_X1 U10589 ( .A1(n9295), .A2(n9315), .ZN(n9296) );
  OAI21_X1 U10590 ( .B1(n9297), .B2(n9291), .A(n9296), .ZN(n9302) );
  OAI22_X1 U10591 ( .A1(n9325), .A2(n9505), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9298), .ZN(n9300) );
  NOR2_X1 U10592 ( .A1(n9538), .A2(n9326), .ZN(n9299) );
  AOI211_X1 U10593 ( .C1(n9509), .C2(n9329), .A(n9300), .B(n9299), .ZN(n9301)
         );
  OAI211_X1 U10594 ( .C1(n9512), .C2(n9332), .A(n9302), .B(n9301), .ZN(
        P1_U3233) );
  NAND2_X1 U10595 ( .A1(n9304), .A2(n9303), .ZN(n9305) );
  XOR2_X1 U10596 ( .A(n9306), .B(n9305), .Z(n9316) );
  NAND2_X1 U10597 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9381) );
  OAI21_X1 U10598 ( .B1(n9537), .B2(n9325), .A(n9381), .ZN(n9307) );
  AOI21_X1 U10599 ( .B1(n9308), .B2(n9344), .A(n9307), .ZN(n9309) );
  OAI21_X1 U10600 ( .B1(n9311), .B2(n9310), .A(n9309), .ZN(n9312) );
  AOI21_X1 U10601 ( .B1(n9647), .B2(n9313), .A(n9312), .ZN(n9314) );
  OAI21_X1 U10602 ( .B1(n9316), .B2(n9315), .A(n9314), .ZN(P1_U3236) );
  INV_X1 U10603 ( .A(n9317), .ZN(n9323) );
  OAI21_X1 U10604 ( .B1(n9251), .B2(n9319), .A(n9318), .ZN(n9321) );
  NAND3_X1 U10605 ( .A1(n9323), .A2(n9322), .A3(n9321), .ZN(n9331) );
  INV_X1 U10606 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9324) );
  OAI22_X1 U10607 ( .A1(n9325), .A2(n9450), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9324), .ZN(n9328) );
  NOR2_X1 U10608 ( .A1(n9326), .A2(n9477), .ZN(n9327) );
  AOI211_X1 U10609 ( .C1(n9455), .C2(n9329), .A(n9328), .B(n9327), .ZN(n9330)
         );
  OAI211_X1 U10610 ( .C1(n4848), .C2(n9332), .A(n9331), .B(n9330), .ZN(
        P1_U3238) );
  MUX2_X1 U10611 ( .A(n9333), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9358), .Z(
        P1_U3585) );
  MUX2_X1 U10612 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9334), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10613 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9335), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10614 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9336), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10615 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9337), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10616 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9338), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10617 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9339), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10618 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9340), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10619 ( .A(n9341), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9358), .Z(
        P1_U3576) );
  MUX2_X1 U10620 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9342), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10621 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9343), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10622 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9577), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10623 ( .A(n9344), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9358), .Z(
        P1_U3572) );
  MUX2_X1 U10624 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9345), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10625 ( .A(n9346), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9358), .Z(
        P1_U3570) );
  MUX2_X1 U10626 ( .A(n9347), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9358), .Z(
        P1_U3569) );
  MUX2_X1 U10627 ( .A(n9752), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9358), .Z(
        P1_U3568) );
  MUX2_X1 U10628 ( .A(n9348), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9358), .Z(
        P1_U3567) );
  MUX2_X1 U10629 ( .A(n9753), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9358), .Z(
        P1_U3566) );
  MUX2_X1 U10630 ( .A(n9349), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9358), .Z(
        P1_U3565) );
  MUX2_X1 U10631 ( .A(n9350), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9358), .Z(
        P1_U3564) );
  MUX2_X1 U10632 ( .A(n9351), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9358), .Z(
        P1_U3563) );
  MUX2_X1 U10633 ( .A(n9352), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9358), .Z(
        P1_U3562) );
  MUX2_X1 U10634 ( .A(n9353), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9358), .Z(
        P1_U3561) );
  MUX2_X1 U10635 ( .A(n9354), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9358), .Z(
        P1_U3560) );
  MUX2_X1 U10636 ( .A(n9355), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9358), .Z(
        P1_U3559) );
  MUX2_X1 U10637 ( .A(n9356), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9358), .Z(
        P1_U3558) );
  MUX2_X1 U10638 ( .A(n9357), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9358), .Z(
        P1_U3557) );
  MUX2_X1 U10639 ( .A(n6529), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9358), .Z(
        P1_U3556) );
  MUX2_X1 U10640 ( .A(n6526), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9358), .Z(
        P1_U3555) );
  INV_X1 U10641 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9392) );
  AOI22_X1 U10642 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n9391), .B1(n9389), .B2(
        n9392), .ZN(n9368) );
  INV_X1 U10643 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9365) );
  XNOR2_X1 U10644 ( .A(n9366), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9919) );
  INV_X1 U10645 ( .A(n9900), .ZN(n9364) );
  INV_X1 U10646 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9363) );
  XOR2_X1 U10647 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9900), .Z(n9902) );
  NAND2_X1 U10648 ( .A1(n9888), .A2(n9361), .ZN(n9362) );
  XNOR2_X1 U10649 ( .A(n9361), .B(n9374), .ZN(n9890) );
  NAND2_X1 U10650 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n9890), .ZN(n9889) );
  NAND2_X1 U10651 ( .A1(n9362), .A2(n9889), .ZN(n9903) );
  NAND2_X1 U10652 ( .A1(n9919), .A2(n9918), .ZN(n9916) );
  OAI21_X1 U10653 ( .B1(n9366), .B2(n9365), .A(n9916), .ZN(n9367) );
  NOR2_X1 U10654 ( .A1(n9368), .A2(n9367), .ZN(n9390) );
  AOI21_X1 U10655 ( .B1(n9368), .B2(n9367), .A(n9390), .ZN(n9387) );
  MUX2_X1 U10656 ( .A(n9369), .B(P1_REG2_REG_18__SCAN_IN), .S(n9389), .Z(n9380) );
  NAND2_X1 U10657 ( .A1(n9371), .A2(n9370), .ZN(n9373) );
  NOR2_X1 U10658 ( .A1(n9374), .A2(n9375), .ZN(n9376) );
  INV_X1 U10659 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9884) );
  NAND2_X1 U10660 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9900), .ZN(n9377) );
  OAI21_X1 U10661 ( .B1(n9900), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9377), .ZN(
        n9896) );
  NOR2_X1 U10662 ( .A1(n9897), .A2(n9896), .ZN(n9895) );
  AOI21_X1 U10663 ( .B1(n9900), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9895), .ZN(
        n9911) );
  NAND2_X1 U10664 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9914), .ZN(n9378) );
  OAI21_X1 U10665 ( .B1(n9914), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9378), .ZN(
        n9910) );
  NOR2_X1 U10666 ( .A1(n9911), .A2(n9910), .ZN(n9909) );
  AOI21_X1 U10667 ( .B1(n9380), .B2(n9379), .A(n9388), .ZN(n9383) );
  INV_X1 U10668 ( .A(n9381), .ZN(n9382) );
  AOI21_X1 U10669 ( .B1(n9862), .B2(n9383), .A(n9382), .ZN(n9384) );
  OAI21_X1 U10670 ( .B1(n9837), .B2(n9391), .A(n9384), .ZN(n9385) );
  AOI21_X1 U10671 ( .B1(n9854), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n9385), .ZN(
        n9386) );
  OAI21_X1 U10672 ( .B1(n9387), .B2(n9879), .A(n9386), .ZN(P1_U3259) );
  INV_X1 U10673 ( .A(n9398), .ZN(n9396) );
  XOR2_X1 U10674 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9393), .Z(n9397) );
  OAI21_X1 U10675 ( .B1(n9397), .B2(n9879), .A(n9837), .ZN(n9394) );
  AOI21_X1 U10676 ( .B1(n9396), .B2(n9395), .A(n9394), .ZN(n9400) );
  AOI22_X1 U10677 ( .A1(n9398), .A2(n9862), .B1(n9917), .B2(n9397), .ZN(n9399)
         );
  MUX2_X1 U10678 ( .A(n9400), .B(n9399), .S(n9930), .Z(n9402) );
  OAI211_X1 U10679 ( .C1(n4882), .C2(n9922), .A(n9402), .B(n9401), .ZN(
        P1_U3260) );
  NAND2_X1 U10680 ( .A1(n9590), .A2(n9408), .ZN(n9587) );
  XNOR2_X1 U10681 ( .A(n9587), .B(n9583), .ZN(n9585) );
  NAND2_X1 U10682 ( .A1(n9404), .A2(n9403), .ZN(n9588) );
  NOR2_X1 U10683 ( .A1(n9578), .A2(n9588), .ZN(n9411) );
  AOI21_X1 U10684 ( .B1(n9578), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9411), .ZN(
        n9406) );
  NAND2_X1 U10685 ( .A1(n9583), .A2(n9941), .ZN(n9405) );
  OAI211_X1 U10686 ( .C1(n9585), .C2(n9407), .A(n9406), .B(n9405), .ZN(
        P1_U3261) );
  INV_X1 U10687 ( .A(n9408), .ZN(n9409) );
  NAND2_X1 U10688 ( .A1(n9410), .A2(n9409), .ZN(n9586) );
  NAND3_X1 U10689 ( .A1(n9587), .A2(n9940), .A3(n9586), .ZN(n9413) );
  AOI21_X1 U10690 ( .B1(n9578), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9411), .ZN(
        n9412) );
  OAI211_X1 U10691 ( .C1(n9590), .C2(n9568), .A(n9413), .B(n9412), .ZN(
        P1_U3262) );
  OAI211_X1 U10692 ( .C1(n9415), .C2(n9433), .A(n9764), .B(n9414), .ZN(n9597)
         );
  NOR2_X1 U10693 ( .A1(n9597), .A2(n9497), .ZN(n9423) );
  INV_X1 U10694 ( .A(n9416), .ZN(n9417) );
  AOI21_X1 U10695 ( .B1(n9417), .B2(n9425), .A(n9572), .ZN(n9421) );
  OAI22_X1 U10696 ( .A1(n9450), .A2(n5531), .B1(n9418), .B2(n9550), .ZN(n9419)
         );
  AOI21_X1 U10697 ( .B1(n9421), .B2(n9420), .A(n9419), .ZN(n9599) );
  INV_X1 U10698 ( .A(n9599), .ZN(n9422) );
  AOI22_X1 U10699 ( .A1(n9596), .A2(n9941), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9578), .ZN(n9429) );
  OR2_X1 U10700 ( .A1(n9426), .A2(n9425), .ZN(n9595) );
  NAND3_X1 U10701 ( .A1(n9595), .A2(n9594), .A3(n9427), .ZN(n9428) );
  OAI211_X1 U10702 ( .C1(n9430), .C2(n9578), .A(n9429), .B(n9428), .ZN(
        P1_U3263) );
  XNOR2_X1 U10703 ( .A(n9432), .B(n9431), .ZN(n9605) );
  AOI21_X1 U10704 ( .B1(n9601), .B2(n9452), .A(n9433), .ZN(n9602) );
  AOI22_X1 U10705 ( .A1(n9578), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9434), .B2(
        n9759), .ZN(n9435) );
  OAI21_X1 U10706 ( .B1(n9436), .B2(n9568), .A(n9435), .ZN(n9443) );
  AOI21_X1 U10707 ( .B1(n4342), .B2(n9437), .A(n9572), .ZN(n9441) );
  OAI22_X1 U10708 ( .A1(n9438), .A2(n9550), .B1(n9465), .B2(n5531), .ZN(n9439)
         );
  AOI21_X1 U10709 ( .B1(n9441), .B2(n9440), .A(n9439), .ZN(n9604) );
  NOR2_X1 U10710 ( .A1(n9604), .A2(n9578), .ZN(n9442) );
  AOI211_X1 U10711 ( .C1(n9940), .C2(n9602), .A(n9443), .B(n9442), .ZN(n9444)
         );
  OAI21_X1 U10712 ( .B1(n9605), .B2(n9582), .A(n9444), .ZN(P1_U3264) );
  XNOR2_X1 U10713 ( .A(n9445), .B(n9448), .ZN(n9611) );
  AOI21_X1 U10714 ( .B1(n9448), .B2(n9447), .A(n9446), .ZN(n9449) );
  OAI222_X1 U10715 ( .A1(n9550), .A2(n9450), .B1(n5531), .B2(n9477), .C1(n9572), .C2(n9449), .ZN(n9606) );
  INV_X1 U10716 ( .A(n9451), .ZN(n9454) );
  INV_X1 U10717 ( .A(n9452), .ZN(n9453) );
  AOI21_X1 U10718 ( .B1(n9607), .B2(n9454), .A(n9453), .ZN(n9608) );
  NAND2_X1 U10719 ( .A1(n9608), .A2(n9940), .ZN(n9457) );
  AOI22_X1 U10720 ( .A1(n9578), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9455), .B2(
        n9759), .ZN(n9456) );
  OAI211_X1 U10721 ( .C1(n4848), .C2(n9568), .A(n9457), .B(n9456), .ZN(n9458)
         );
  AOI21_X1 U10722 ( .B1(n9606), .B2(n9945), .A(n9458), .ZN(n9459) );
  OAI21_X1 U10723 ( .B1(n9611), .B2(n9582), .A(n9459), .ZN(P1_U3265) );
  XNOR2_X1 U10724 ( .A(n9460), .B(n4839), .ZN(n9616) );
  XNOR2_X1 U10725 ( .A(n9463), .B(n9478), .ZN(n9613) );
  AOI22_X1 U10726 ( .A1(n9578), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9461), .B2(
        n9759), .ZN(n9462) );
  OAI21_X1 U10727 ( .B1(n9463), .B2(n9568), .A(n9462), .ZN(n9470) );
  AOI21_X1 U10728 ( .B1(n4341), .B2(n9464), .A(n9572), .ZN(n9468) );
  OAI22_X1 U10729 ( .A1(n9465), .A2(n9550), .B1(n9491), .B2(n5531), .ZN(n9466)
         );
  AOI21_X1 U10730 ( .B1(n9468), .B2(n9467), .A(n9466), .ZN(n9615) );
  NOR2_X1 U10731 ( .A1(n9615), .A2(n9578), .ZN(n9469) );
  AOI211_X1 U10732 ( .C1(n9613), .C2(n9940), .A(n9470), .B(n9469), .ZN(n9471)
         );
  OAI21_X1 U10733 ( .B1(n9616), .B2(n9582), .A(n9471), .ZN(P1_U3266) );
  XOR2_X1 U10734 ( .A(n9472), .B(n9475), .Z(n9621) );
  AOI22_X1 U10735 ( .A1(n9619), .A2(n9941), .B1(n9578), .B2(
        P1_REG2_REG_24__SCAN_IN), .ZN(n9486) );
  AOI21_X1 U10736 ( .B1(n9475), .B2(n9474), .A(n9473), .ZN(n9476) );
  OAI222_X1 U10737 ( .A1(n5531), .A2(n9505), .B1(n9550), .B2(n9477), .C1(n9572), .C2(n9476), .ZN(n9617) );
  INV_X1 U10738 ( .A(n9494), .ZN(n9480) );
  INV_X1 U10739 ( .A(n9478), .ZN(n9479) );
  AOI211_X1 U10740 ( .C1(n9619), .C2(n9480), .A(n9975), .B(n9479), .ZN(n9618)
         );
  INV_X1 U10741 ( .A(n9618), .ZN(n9483) );
  INV_X1 U10742 ( .A(n9481), .ZN(n9482) );
  OAI22_X1 U10743 ( .A1(n9483), .A2(n9497), .B1(n9949), .B2(n9482), .ZN(n9484)
         );
  OAI21_X1 U10744 ( .B1(n9617), .B2(n9484), .A(n9945), .ZN(n9485) );
  OAI211_X1 U10745 ( .C1(n9621), .C2(n9582), .A(n9486), .B(n9485), .ZN(
        P1_U3267) );
  XNOR2_X1 U10746 ( .A(n9487), .B(n9489), .ZN(n9626) );
  AOI22_X1 U10747 ( .A1(n9624), .A2(n9941), .B1(n9578), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n9501) );
  OAI211_X1 U10748 ( .C1(n9490), .C2(n9489), .A(n9488), .B(n9747), .ZN(n9493)
         );
  OR2_X1 U10749 ( .A1(n9491), .A2(n9550), .ZN(n9492) );
  OAI211_X1 U10750 ( .C1(n9522), .C2(n5531), .A(n9493), .B(n9492), .ZN(n9622)
         );
  AOI211_X1 U10751 ( .C1(n9624), .C2(n9506), .A(n9975), .B(n9494), .ZN(n9623)
         );
  INV_X1 U10752 ( .A(n9623), .ZN(n9498) );
  INV_X1 U10753 ( .A(n9495), .ZN(n9496) );
  OAI22_X1 U10754 ( .A1(n9498), .A2(n9497), .B1(n9949), .B2(n9496), .ZN(n9499)
         );
  OAI21_X1 U10755 ( .B1(n9622), .B2(n9499), .A(n9945), .ZN(n9500) );
  OAI211_X1 U10756 ( .C1(n9626), .C2(n9582), .A(n9501), .B(n9500), .ZN(
        P1_U3268) );
  XNOR2_X1 U10757 ( .A(n4333), .B(n9503), .ZN(n9631) );
  XOR2_X1 U10758 ( .A(n9503), .B(n9502), .Z(n9504) );
  OAI222_X1 U10759 ( .A1(n5531), .A2(n9538), .B1(n9550), .B2(n9505), .C1(n9504), .C2(n9572), .ZN(n9627) );
  INV_X1 U10760 ( .A(n9523), .ZN(n9508) );
  INV_X1 U10761 ( .A(n9506), .ZN(n9507) );
  AOI211_X1 U10762 ( .C1(n9629), .C2(n9508), .A(n9975), .B(n9507), .ZN(n9628)
         );
  NAND2_X1 U10763 ( .A1(n9628), .A2(n9767), .ZN(n9511) );
  AOI22_X1 U10764 ( .A1(n9578), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9509), .B2(
        n9759), .ZN(n9510) );
  OAI211_X1 U10765 ( .C1(n9512), .C2(n9568), .A(n9511), .B(n9510), .ZN(n9513)
         );
  AOI21_X1 U10766 ( .B1(n9627), .B2(n9945), .A(n9513), .ZN(n9514) );
  OAI21_X1 U10767 ( .B1(n9631), .B2(n9582), .A(n9514), .ZN(P1_U3269) );
  XNOR2_X1 U10768 ( .A(n9516), .B(n9515), .ZN(n9636) );
  INV_X1 U10769 ( .A(n9517), .ZN(n9520) );
  AOI21_X1 U10770 ( .B1(n9540), .B2(n9518), .A(n5354), .ZN(n9519) );
  NOR2_X1 U10771 ( .A1(n9520), .A2(n9519), .ZN(n9521) );
  OAI222_X1 U10772 ( .A1(n9550), .A2(n9522), .B1(n5531), .B2(n9549), .C1(n9572), .C2(n9521), .ZN(n9632) );
  AOI211_X1 U10773 ( .C1(n9634), .C2(n9531), .A(n9975), .B(n9523), .ZN(n9633)
         );
  NAND2_X1 U10774 ( .A1(n9633), .A2(n9767), .ZN(n9527) );
  INV_X1 U10775 ( .A(n9524), .ZN(n9525) );
  AOI22_X1 U10776 ( .A1(n9525), .A2(n9759), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9578), .ZN(n9526) );
  OAI211_X1 U10777 ( .C1(n4525), .C2(n9568), .A(n9527), .B(n9526), .ZN(n9528)
         );
  AOI21_X1 U10778 ( .B1(n9632), .B2(n9945), .A(n9528), .ZN(n9529) );
  OAI21_X1 U10779 ( .B1(n9636), .B2(n9582), .A(n9529), .ZN(P1_U3270) );
  XOR2_X1 U10780 ( .A(n9536), .B(n9530), .Z(n9641) );
  INV_X1 U10781 ( .A(n9531), .ZN(n9532) );
  AOI21_X1 U10782 ( .B1(n9637), .B2(n4529), .A(n9532), .ZN(n9638) );
  AOI22_X1 U10783 ( .A1(n9533), .A2(n9759), .B1(n9578), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n9534) );
  OAI21_X1 U10784 ( .B1(n9535), .B2(n9568), .A(n9534), .ZN(n9543) );
  AOI21_X1 U10785 ( .B1(n4547), .B2(n4550), .A(n9572), .ZN(n9541) );
  OAI22_X1 U10786 ( .A1(n9538), .A2(n9550), .B1(n9537), .B2(n5531), .ZN(n9539)
         );
  AOI21_X1 U10787 ( .B1(n9541), .B2(n9540), .A(n9539), .ZN(n9640) );
  NOR2_X1 U10788 ( .A1(n9640), .A2(n9578), .ZN(n9542) );
  AOI211_X1 U10789 ( .C1(n9638), .C2(n9940), .A(n9543), .B(n9542), .ZN(n9544)
         );
  OAI21_X1 U10790 ( .B1(n9641), .B2(n9582), .A(n9544), .ZN(P1_U3271) );
  XOR2_X1 U10791 ( .A(n9547), .B(n9545), .Z(n9646) );
  XOR2_X1 U10792 ( .A(n9547), .B(n9546), .Z(n9548) );
  OAI222_X1 U10793 ( .A1(n5531), .A2(n9551), .B1(n9550), .B2(n9549), .C1(n9548), .C2(n9572), .ZN(n9642) );
  AOI211_X1 U10794 ( .C1(n9644), .C2(n9553), .A(n9975), .B(n9552), .ZN(n9643)
         );
  NAND2_X1 U10795 ( .A1(n9643), .A2(n9767), .ZN(n9557) );
  INV_X1 U10796 ( .A(n9554), .ZN(n9555) );
  AOI22_X1 U10797 ( .A1(P1_REG2_REG_19__SCAN_IN), .A2(n9578), .B1(n9555), .B2(
        n9759), .ZN(n9556) );
  OAI211_X1 U10798 ( .C1(n9558), .C2(n9568), .A(n9557), .B(n9556), .ZN(n9559)
         );
  AOI21_X1 U10799 ( .B1(n9642), .B2(n9945), .A(n9559), .ZN(n9560) );
  OAI21_X1 U10800 ( .B1(n9582), .B2(n9646), .A(n9560), .ZN(P1_U3272) );
  XNOR2_X1 U10801 ( .A(n9562), .B(n9561), .ZN(n9657) );
  AOI211_X1 U10802 ( .C1(n9654), .C2(n9564), .A(n9975), .B(n9563), .ZN(n9653)
         );
  INV_X1 U10803 ( .A(n9654), .ZN(n9569) );
  INV_X1 U10804 ( .A(n9565), .ZN(n9566) );
  AOI22_X1 U10805 ( .A1(n9578), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9566), .B2(
        n9759), .ZN(n9567) );
  OAI21_X1 U10806 ( .B1(n9569), .B2(n9568), .A(n9567), .ZN(n9580) );
  NOR2_X1 U10807 ( .A1(n9570), .A2(n5531), .ZN(n9576) );
  AOI211_X1 U10808 ( .C1(n9574), .C2(n9573), .A(n9572), .B(n9571), .ZN(n9575)
         );
  AOI211_X1 U10809 ( .C1(n9751), .C2(n9577), .A(n9576), .B(n9575), .ZN(n9656)
         );
  NOR2_X1 U10810 ( .A1(n9656), .A2(n9578), .ZN(n9579) );
  AOI211_X1 U10811 ( .C1(n9653), .C2(n9767), .A(n9580), .B(n9579), .ZN(n9581)
         );
  OAI21_X1 U10812 ( .B1(n9582), .B2(n9657), .A(n9581), .ZN(P1_U3274) );
  NAND2_X1 U10813 ( .A1(n9583), .A2(n9670), .ZN(n9584) );
  OAI211_X1 U10814 ( .C1(n9585), .C2(n9975), .A(n9584), .B(n9588), .ZN(n9674)
         );
  MUX2_X1 U10815 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9674), .S(n9990), .Z(
        P1_U3554) );
  NAND3_X1 U10816 ( .A1(n9587), .A2(n9764), .A3(n9586), .ZN(n9589) );
  OAI211_X1 U10817 ( .C1(n9590), .C2(n9973), .A(n9589), .B(n9588), .ZN(n9675)
         );
  MUX2_X1 U10818 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9675), .S(n9990), .Z(
        P1_U3553) );
  MUX2_X1 U10819 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9676), .S(n9990), .Z(
        P1_U3552) );
  INV_X1 U10820 ( .A(n9672), .ZN(n9787) );
  NAND3_X1 U10821 ( .A1(n9595), .A2(n9594), .A3(n9787), .ZN(n9600) );
  NAND2_X1 U10822 ( .A1(n9596), .A2(n9670), .ZN(n9598) );
  NAND4_X1 U10823 ( .A1(n9600), .A2(n9599), .A3(n9598), .A4(n9597), .ZN(n9677)
         );
  MUX2_X1 U10824 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9677), .S(n9990), .Z(
        P1_U3551) );
  AOI22_X1 U10825 ( .A1(n9602), .A2(n9764), .B1(n9670), .B2(n9601), .ZN(n9603)
         );
  OAI211_X1 U10826 ( .C1(n9605), .C2(n9672), .A(n9604), .B(n9603), .ZN(n9678)
         );
  MUX2_X1 U10827 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9678), .S(n9990), .Z(
        P1_U3550) );
  INV_X1 U10828 ( .A(n9606), .ZN(n9610) );
  AOI22_X1 U10829 ( .A1(n9608), .A2(n9764), .B1(n9670), .B2(n9607), .ZN(n9609)
         );
  OAI211_X1 U10830 ( .C1(n9611), .C2(n9672), .A(n9610), .B(n9609), .ZN(n9679)
         );
  MUX2_X1 U10831 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9679), .S(n9990), .Z(
        P1_U3549) );
  AOI22_X1 U10832 ( .A1(n9613), .A2(n9764), .B1(n9670), .B2(n9612), .ZN(n9614)
         );
  OAI211_X1 U10833 ( .C1(n9616), .C2(n9672), .A(n9615), .B(n9614), .ZN(n9680)
         );
  MUX2_X1 U10834 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9680), .S(n9990), .Z(
        P1_U3548) );
  AOI211_X1 U10835 ( .C1(n9670), .C2(n9619), .A(n9618), .B(n9617), .ZN(n9620)
         );
  OAI21_X1 U10836 ( .B1(n9621), .B2(n9672), .A(n9620), .ZN(n9681) );
  MUX2_X1 U10837 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9681), .S(n9990), .Z(
        P1_U3547) );
  AOI211_X1 U10838 ( .C1(n9670), .C2(n9624), .A(n9623), .B(n9622), .ZN(n9625)
         );
  OAI21_X1 U10839 ( .B1(n9626), .B2(n9672), .A(n9625), .ZN(n9682) );
  MUX2_X1 U10840 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9682), .S(n9990), .Z(
        P1_U3546) );
  AOI211_X1 U10841 ( .C1(n9670), .C2(n9629), .A(n9628), .B(n9627), .ZN(n9630)
         );
  OAI21_X1 U10842 ( .B1(n9672), .B2(n9631), .A(n9630), .ZN(n9683) );
  MUX2_X1 U10843 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9683), .S(n9990), .Z(
        P1_U3545) );
  AOI211_X1 U10844 ( .C1(n9670), .C2(n9634), .A(n9633), .B(n9632), .ZN(n9635)
         );
  OAI21_X1 U10845 ( .B1(n9672), .B2(n9636), .A(n9635), .ZN(n9684) );
  MUX2_X1 U10846 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9684), .S(n9990), .Z(
        P1_U3544) );
  AOI22_X1 U10847 ( .A1(n9638), .A2(n9764), .B1(n9670), .B2(n9637), .ZN(n9639)
         );
  OAI211_X1 U10848 ( .C1(n9641), .C2(n9672), .A(n9640), .B(n9639), .ZN(n9685)
         );
  MUX2_X1 U10849 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9685), .S(n9990), .Z(
        P1_U3543) );
  AOI211_X1 U10850 ( .C1(n9670), .C2(n9644), .A(n9643), .B(n9642), .ZN(n9645)
         );
  OAI21_X1 U10851 ( .B1(n9672), .B2(n9646), .A(n9645), .ZN(n9686) );
  MUX2_X1 U10852 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9686), .S(n9990), .Z(
        P1_U3542) );
  AOI22_X1 U10853 ( .A1(n9648), .A2(n9764), .B1(n9670), .B2(n9647), .ZN(n9651)
         );
  NAND3_X1 U10854 ( .A1(n9649), .A2(n9787), .A3(n8211), .ZN(n9650) );
  NAND3_X1 U10855 ( .A1(n9652), .A2(n9651), .A3(n9650), .ZN(n9687) );
  MUX2_X1 U10856 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9687), .S(n9990), .Z(
        P1_U3541) );
  AOI21_X1 U10857 ( .B1(n9670), .B2(n9654), .A(n9653), .ZN(n9655) );
  OAI211_X1 U10858 ( .C1(n9672), .C2(n9657), .A(n9656), .B(n9655), .ZN(n9688)
         );
  MUX2_X1 U10859 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9688), .S(n9990), .Z(
        P1_U3540) );
  AOI211_X1 U10860 ( .C1(n9670), .C2(n5294), .A(n9659), .B(n9658), .ZN(n9660)
         );
  OAI21_X1 U10861 ( .B1(n9661), .B2(n9672), .A(n9660), .ZN(n9689) );
  MUX2_X1 U10862 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9689), .S(n9990), .Z(
        P1_U3539) );
  AOI22_X1 U10863 ( .A1(n9663), .A2(n9764), .B1(n9670), .B2(n9662), .ZN(n9664)
         );
  OAI211_X1 U10864 ( .C1(n9666), .C2(n9672), .A(n9665), .B(n9664), .ZN(n9690)
         );
  MUX2_X1 U10865 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9690), .S(n9990), .Z(
        P1_U3538) );
  AOI211_X1 U10866 ( .C1(n9670), .C2(n9669), .A(n9668), .B(n9667), .ZN(n9671)
         );
  OAI21_X1 U10867 ( .B1(n9673), .B2(n9672), .A(n9671), .ZN(n9691) );
  MUX2_X1 U10868 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9691), .S(n9990), .Z(
        P1_U3537) );
  MUX2_X1 U10869 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9674), .S(n9983), .Z(
        P1_U3522) );
  MUX2_X1 U10870 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9675), .S(n9983), .Z(
        P1_U3521) );
  MUX2_X1 U10871 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9677), .S(n9983), .Z(
        P1_U3519) );
  MUX2_X1 U10872 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9678), .S(n9983), .Z(
        P1_U3518) );
  MUX2_X1 U10873 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9679), .S(n9983), .Z(
        P1_U3517) );
  MUX2_X1 U10874 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9680), .S(n9983), .Z(
        P1_U3516) );
  MUX2_X1 U10875 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9681), .S(n9983), .Z(
        P1_U3515) );
  MUX2_X1 U10876 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9682), .S(n9983), .Z(
        P1_U3514) );
  MUX2_X1 U10877 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9683), .S(n9983), .Z(
        P1_U3513) );
  MUX2_X1 U10878 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9684), .S(n9983), .Z(
        P1_U3512) );
  MUX2_X1 U10879 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9685), .S(n9983), .Z(
        P1_U3511) );
  MUX2_X1 U10880 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9686), .S(n9983), .Z(
        P1_U3510) );
  MUX2_X1 U10881 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9687), .S(n9983), .Z(
        P1_U3508) );
  MUX2_X1 U10882 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9688), .S(n9983), .Z(
        P1_U3505) );
  MUX2_X1 U10883 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9689), .S(n9983), .Z(
        P1_U3502) );
  MUX2_X1 U10884 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9690), .S(n9983), .Z(
        P1_U3499) );
  MUX2_X1 U10885 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9691), .S(n9983), .Z(
        P1_U3496) );
  MUX2_X1 U10886 ( .A(P1_REG0_REG_10__SCAN_IN), .B(n9692), .S(n9983), .Z(
        P1_U3484) );
  MUX2_X1 U10887 ( .A(P1_D_REG_1__SCAN_IN), .B(n9693), .S(n9951), .Z(P1_U3441)
         );
  MUX2_X1 U10888 ( .A(P1_D_REG_0__SCAN_IN), .B(n9694), .S(n9951), .Z(P1_U3440)
         );
  NOR4_X1 U10889 ( .A1(n5018), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n9695), .ZN(n9696) );
  AOI21_X1 U10890 ( .B1(n9697), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9696), .ZN(
        n9698) );
  OAI21_X1 U10891 ( .B1(n9700), .B2(n9699), .A(n9698), .ZN(P1_U3322) );
  OAI222_X1 U10892 ( .A1(P1_U3084), .A2(n9703), .B1(n9707), .B2(n9702), .C1(
        n9701), .C2(n9704), .ZN(P1_U3323) );
  OAI222_X1 U10893 ( .A1(P1_U3084), .A2(n9708), .B1(n9707), .B2(n9706), .C1(
        n9705), .C2(n9704), .ZN(P1_U3324) );
  MUX2_X1 U10894 ( .A(n9709), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  NAND2_X1 U10895 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9711) );
  AOI21_X1 U10896 ( .B1(n9712), .B2(n9711), .A(n9710), .ZN(n9713) );
  NAND2_X1 U10897 ( .A1(n10008), .A2(n9713), .ZN(n9717) );
  OAI22_X1 U10898 ( .A1(n9714), .A2(n10124), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7111), .ZN(n9715) );
  INV_X1 U10899 ( .A(n9715), .ZN(n9716) );
  OAI211_X1 U10900 ( .C1(n10009), .C2(n9718), .A(n9717), .B(n9716), .ZN(n9719)
         );
  INV_X1 U10901 ( .A(n9719), .ZN(n9724) );
  NOR2_X1 U10902 ( .A1(n10016), .A2(n10106), .ZN(n9721) );
  OAI211_X1 U10903 ( .C1(n9722), .C2(n9721), .A(n10007), .B(n9720), .ZN(n9723)
         );
  NAND2_X1 U10904 ( .A1(n9724), .A2(n9723), .ZN(P2_U3246) );
  AOI22_X1 U10905 ( .A1(n10013), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9737) );
  AOI211_X1 U10906 ( .C1(n9728), .C2(n9727), .A(n9726), .B(n9725), .ZN(n9729)
         );
  AOI21_X1 U10907 ( .B1(n9731), .B2(n9730), .A(n9729), .ZN(n9736) );
  OAI211_X1 U10908 ( .C1(n9734), .C2(n9733), .A(n10007), .B(n9732), .ZN(n9735)
         );
  NAND3_X1 U10909 ( .A1(n9737), .A2(n9736), .A3(n9735), .ZN(P2_U3247) );
  OAI22_X1 U10910 ( .A1(n9739), .A2(n10097), .B1(n9738), .B2(n10095), .ZN(
        n9741) );
  AOI211_X1 U10911 ( .C1(n9742), .C2(n10101), .A(n9741), .B(n9740), .ZN(n9743)
         );
  AOI22_X1 U10912 ( .A1(n10119), .A2(n9743), .B1(n7779), .B2(n10117), .ZN(
        P2_U3534) );
  AOI22_X1 U10913 ( .A1(n10105), .A2(n9743), .B1(n5833), .B2(n10103), .ZN(
        P2_U3493) );
  INV_X1 U10914 ( .A(n9744), .ZN(n9745) );
  AOI21_X1 U10915 ( .B1(n9749), .B2(n9746), .A(n9745), .ZN(n9781) );
  OAI211_X1 U10916 ( .C1(n9750), .C2(n9749), .A(n9748), .B(n9747), .ZN(n9756)
         );
  AOI22_X1 U10917 ( .A1(n9754), .A2(n9753), .B1(n9752), .B2(n9751), .ZN(n9755)
         );
  NAND2_X1 U10918 ( .A1(n9756), .A2(n9755), .ZN(n9757) );
  AOI21_X1 U10919 ( .B1(n9781), .B2(n9758), .A(n9757), .ZN(n9778) );
  AOI222_X1 U10920 ( .A1(n9761), .A2(n9941), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n9578), .C1(n9760), .C2(n9759), .ZN(n9770) );
  INV_X1 U10921 ( .A(n9762), .ZN(n9765) );
  OAI211_X1 U10922 ( .C1(n9765), .C2(n4532), .A(n9764), .B(n9763), .ZN(n9777)
         );
  INV_X1 U10923 ( .A(n9777), .ZN(n9766) );
  AOI22_X1 U10924 ( .A1(n9781), .A2(n9768), .B1(n9767), .B2(n9766), .ZN(n9769)
         );
  OAI211_X1 U10925 ( .C1(n9578), .C2(n9778), .A(n9770), .B(n9769), .ZN(
        P1_U3279) );
  OAI22_X1 U10926 ( .A1(n9771), .A2(n9975), .B1(n4535), .B2(n9973), .ZN(n9772)
         );
  AOI21_X1 U10927 ( .B1(n9773), .B2(n9980), .A(n9772), .ZN(n9774) );
  AND2_X1 U10928 ( .A1(n9775), .A2(n9774), .ZN(n9791) );
  AOI22_X1 U10929 ( .A1(n9990), .A2(n9791), .B1(n9776), .B2(n9987), .ZN(
        P1_U3536) );
  OAI21_X1 U10930 ( .B1(n4532), .B2(n9973), .A(n9777), .ZN(n9780) );
  INV_X1 U10931 ( .A(n9778), .ZN(n9779) );
  AOI211_X1 U10932 ( .C1(n9980), .C2(n9781), .A(n9780), .B(n9779), .ZN(n9793)
         );
  AOI22_X1 U10933 ( .A1(n9990), .A2(n9793), .B1(n9782), .B2(n9987), .ZN(
        P1_U3535) );
  OAI22_X1 U10934 ( .A1(n9784), .A2(n9975), .B1(n9783), .B2(n9973), .ZN(n9785)
         );
  AOI211_X1 U10935 ( .C1(n9788), .C2(n9787), .A(n9786), .B(n9785), .ZN(n9795)
         );
  AOI22_X1 U10936 ( .A1(n9990), .A2(n9795), .B1(n9789), .B2(n9987), .ZN(
        P1_U3534) );
  INV_X1 U10937 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9790) );
  AOI22_X1 U10938 ( .A1(n9983), .A2(n9791), .B1(n9790), .B2(n9981), .ZN(
        P1_U3493) );
  INV_X1 U10939 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9792) );
  AOI22_X1 U10940 ( .A1(n9983), .A2(n9793), .B1(n9792), .B2(n9981), .ZN(
        P1_U3490) );
  INV_X1 U10941 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9794) );
  AOI22_X1 U10942 ( .A1(n9983), .A2(n9795), .B1(n9794), .B2(n9981), .ZN(
        P1_U3487) );
  XNOR2_X1 U10943 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XOR2_X1 U10944 ( .A(n9796), .B(P2_RD_REG_SCAN_IN), .Z(U126) );
  AOI22_X1 U10945 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n9854), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3084), .ZN(n9807) );
  XOR2_X1 U10946 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9797), .Z(n9802) );
  INV_X1 U10947 ( .A(n9798), .ZN(n9800) );
  OAI21_X1 U10948 ( .B1(n9800), .B2(n9804), .A(n9799), .ZN(n9801) );
  NAND3_X1 U10949 ( .A1(n9803), .A2(n9802), .A3(n9801), .ZN(n9806) );
  NAND3_X1 U10950 ( .A1(n9917), .A2(P1_IR_REG_0__SCAN_IN), .A3(n9804), .ZN(
        n9805) );
  NAND3_X1 U10951 ( .A1(n9807), .A2(n9806), .A3(n9805), .ZN(P1_U3241) );
  OAI22_X1 U10952 ( .A1(n9837), .A2(n5068), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7013), .ZN(n9808) );
  AOI21_X1 U10953 ( .B1(n9854), .B2(P1_ADDR_REG_2__SCAN_IN), .A(n9808), .ZN(
        n9818) );
  OAI211_X1 U10954 ( .C1(n9811), .C2(n9810), .A(n9862), .B(n9809), .ZN(n9816)
         );
  XOR2_X1 U10955 ( .A(n9813), .B(n9812), .Z(n9814) );
  NAND2_X1 U10956 ( .A1(n9917), .A2(n9814), .ZN(n9815) );
  NAND4_X1 U10957 ( .A1(n9818), .A2(n9817), .A3(n9816), .A4(n9815), .ZN(
        P1_U3243) );
  AOI22_X1 U10958 ( .A1(n9854), .A2(P1_ADDR_REG_5__SCAN_IN), .B1(n9915), .B2(
        n9819), .ZN(n9835) );
  INV_X1 U10959 ( .A(n9820), .ZN(n9827) );
  INV_X1 U10960 ( .A(n9821), .ZN(n9825) );
  INV_X1 U10961 ( .A(n9822), .ZN(n9824) );
  NOR3_X1 U10962 ( .A1(n9825), .A2(n9824), .A3(n9823), .ZN(n9826) );
  OAI21_X1 U10963 ( .B1(n9827), .B2(n9826), .A(n9862), .ZN(n9833) );
  NAND2_X1 U10964 ( .A1(n9829), .A2(n9828), .ZN(n9830) );
  NAND3_X1 U10965 ( .A1(n9917), .A2(n9831), .A3(n9830), .ZN(n9832) );
  NAND4_X1 U10966 ( .A1(n9835), .A2(n9834), .A3(n9833), .A4(n9832), .ZN(
        P1_U3246) );
  INV_X1 U10967 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9839) );
  OR2_X1 U10968 ( .A1(n9837), .A2(n9836), .ZN(n9838) );
  OAI21_X1 U10969 ( .B1(n9922), .B2(n9839), .A(n9838), .ZN(n9840) );
  INV_X1 U10970 ( .A(n9840), .ZN(n9852) );
  AOI21_X1 U10971 ( .B1(n9843), .B2(n9842), .A(n9841), .ZN(n9844) );
  OR2_X1 U10972 ( .A1(n9844), .A2(n9879), .ZN(n9850) );
  OAI21_X1 U10973 ( .B1(n9847), .B2(n9846), .A(n9845), .ZN(n9848) );
  NAND2_X1 U10974 ( .A1(n9848), .A2(n9862), .ZN(n9849) );
  NAND4_X1 U10975 ( .A1(n9852), .A2(n9851), .A3(n9850), .A4(n9849), .ZN(
        P1_U3248) );
  AOI22_X1 U10976 ( .A1(n9854), .A2(P1_ADDR_REG_8__SCAN_IN), .B1(n9915), .B2(
        n9853), .ZN(n9867) );
  AOI21_X1 U10977 ( .B1(n9857), .B2(n9856), .A(n9855), .ZN(n9858) );
  OR2_X1 U10978 ( .A1(n9858), .A2(n9879), .ZN(n9865) );
  OAI21_X1 U10979 ( .B1(n9861), .B2(n9860), .A(n9859), .ZN(n9863) );
  NAND2_X1 U10980 ( .A1(n9863), .A2(n9862), .ZN(n9864) );
  NAND4_X1 U10981 ( .A1(n9867), .A2(n9866), .A3(n9865), .A4(n9864), .ZN(
        P1_U3249) );
  INV_X1 U10982 ( .A(n9868), .ZN(n9873) );
  AOI211_X1 U10983 ( .C1(n9871), .C2(n9870), .A(n9869), .B(n9908), .ZN(n9872)
         );
  AOI211_X1 U10984 ( .C1(n9915), .C2(n9874), .A(n9873), .B(n9872), .ZN(n9881)
         );
  AOI21_X1 U10985 ( .B1(n9877), .B2(n9876), .A(n9875), .ZN(n9878) );
  OR2_X1 U10986 ( .A1(n9879), .A2(n9878), .ZN(n9880) );
  OAI211_X1 U10987 ( .C1(n10161), .C2(n9922), .A(n9881), .B(n9880), .ZN(
        P1_U3250) );
  INV_X1 U10988 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9893) );
  INV_X1 U10989 ( .A(n9882), .ZN(n9887) );
  AOI211_X1 U10990 ( .C1(n9885), .C2(n9884), .A(n9883), .B(n9908), .ZN(n9886)
         );
  AOI211_X1 U10991 ( .C1(n9915), .C2(n9888), .A(n9887), .B(n9886), .ZN(n9892)
         );
  OAI211_X1 U10992 ( .C1(n9890), .C2(P1_REG1_REG_15__SCAN_IN), .A(n9917), .B(
        n9889), .ZN(n9891) );
  OAI211_X1 U10993 ( .C1(n9893), .C2(n9922), .A(n9892), .B(n9891), .ZN(
        P1_U3256) );
  INV_X1 U10994 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9906) );
  INV_X1 U10995 ( .A(n9894), .ZN(n9899) );
  AOI211_X1 U10996 ( .C1(n9897), .C2(n9896), .A(n9895), .B(n9908), .ZN(n9898)
         );
  AOI211_X1 U10997 ( .C1(n9915), .C2(n9900), .A(n9899), .B(n9898), .ZN(n9905)
         );
  OAI211_X1 U10998 ( .C1(n9903), .C2(n9902), .A(n9917), .B(n9901), .ZN(n9904)
         );
  OAI211_X1 U10999 ( .C1(n9906), .C2(n9922), .A(n9905), .B(n9904), .ZN(
        P1_U3257) );
  INV_X1 U11000 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9923) );
  INV_X1 U11001 ( .A(n9907), .ZN(n9913) );
  AOI211_X1 U11002 ( .C1(n9911), .C2(n9910), .A(n9909), .B(n9908), .ZN(n9912)
         );
  AOI211_X1 U11003 ( .C1(n9915), .C2(n9914), .A(n9913), .B(n9912), .ZN(n9921)
         );
  OAI211_X1 U11004 ( .C1(n9919), .C2(n9918), .A(n9917), .B(n9916), .ZN(n9920)
         );
  OAI211_X1 U11005 ( .C1(n9923), .C2(n9922), .A(n9921), .B(n9920), .ZN(
        P1_U3258) );
  INV_X1 U11006 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9938) );
  INV_X1 U11007 ( .A(n9924), .ZN(n9934) );
  NAND2_X1 U11008 ( .A1(n9926), .A2(n9925), .ZN(n9927) );
  OAI21_X1 U11009 ( .B1(n9949), .B2(n9928), .A(n9927), .ZN(n9929) );
  AOI21_X1 U11010 ( .B1(n9931), .B2(n9930), .A(n9929), .ZN(n9932) );
  OAI211_X1 U11011 ( .C1(n9935), .C2(n9934), .A(n9933), .B(n9932), .ZN(n9936)
         );
  INV_X1 U11012 ( .A(n9936), .ZN(n9937) );
  AOI22_X1 U11013 ( .A1(n9578), .A2(n9938), .B1(n9937), .B2(n9945), .ZN(
        P1_U3286) );
  INV_X1 U11014 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9948) );
  NAND2_X1 U11015 ( .A1(n9939), .A2(n9945), .ZN(n9943) );
  OAI21_X1 U11016 ( .B1(n9941), .B2(n9940), .A(n6519), .ZN(n9942) );
  OAI211_X1 U11017 ( .C1(n9945), .C2(n9944), .A(n9943), .B(n9942), .ZN(n9946)
         );
  INV_X1 U11018 ( .A(n9946), .ZN(n9947) );
  OAI21_X1 U11019 ( .B1(n9949), .B2(n9948), .A(n9947), .ZN(P1_U3291) );
  AND2_X1 U11020 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9958), .ZN(P1_U3292) );
  NOR2_X1 U11021 ( .A1(n9957), .A2(n9952), .ZN(P1_U3293) );
  AND2_X1 U11022 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9958), .ZN(P1_U3294) );
  AND2_X1 U11023 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9958), .ZN(P1_U3295) );
  AND2_X1 U11024 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9958), .ZN(P1_U3296) );
  AND2_X1 U11025 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9958), .ZN(P1_U3297) );
  AND2_X1 U11026 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9958), .ZN(P1_U3298) );
  AND2_X1 U11027 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9958), .ZN(P1_U3299) );
  AND2_X1 U11028 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9958), .ZN(P1_U3300) );
  AND2_X1 U11029 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9958), .ZN(P1_U3301) );
  AND2_X1 U11030 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9958), .ZN(P1_U3302) );
  AND2_X1 U11031 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9958), .ZN(P1_U3303) );
  AND2_X1 U11032 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9958), .ZN(P1_U3304) );
  NOR2_X1 U11033 ( .A1(n9957), .A2(n9953), .ZN(P1_U3305) );
  NOR2_X1 U11034 ( .A1(n9957), .A2(n9954), .ZN(P1_U3306) );
  AND2_X1 U11035 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9958), .ZN(P1_U3307) );
  AND2_X1 U11036 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9958), .ZN(P1_U3308) );
  AND2_X1 U11037 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9958), .ZN(P1_U3309) );
  AND2_X1 U11038 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9958), .ZN(P1_U3310) );
  NOR2_X1 U11039 ( .A1(n9957), .A2(n9955), .ZN(P1_U3311) );
  AND2_X1 U11040 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9958), .ZN(P1_U3312) );
  AND2_X1 U11041 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9958), .ZN(P1_U3313) );
  AND2_X1 U11042 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9958), .ZN(P1_U3314) );
  AND2_X1 U11043 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9958), .ZN(P1_U3315) );
  AND2_X1 U11044 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9958), .ZN(P1_U3316) );
  AND2_X1 U11045 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9958), .ZN(P1_U3317) );
  NOR2_X1 U11046 ( .A1(n9957), .A2(n9956), .ZN(P1_U3318) );
  AND2_X1 U11047 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9958), .ZN(P1_U3319) );
  AND2_X1 U11048 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9958), .ZN(P1_U3320) );
  AND2_X1 U11049 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9958), .ZN(P1_U3321) );
  AOI22_X1 U11050 ( .A1(n9983), .A2(n9960), .B1(n9959), .B2(n9981), .ZN(
        P1_U3460) );
  OAI22_X1 U11051 ( .A1(n9962), .A2(n9975), .B1(n9961), .B2(n9973), .ZN(n9964)
         );
  AOI211_X1 U11052 ( .C1(n9980), .C2(n9965), .A(n9964), .B(n9963), .ZN(n9984)
         );
  INV_X1 U11053 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9966) );
  AOI22_X1 U11054 ( .A1(n9983), .A2(n9984), .B1(n9966), .B2(n9981), .ZN(
        P1_U3466) );
  OAI22_X1 U11055 ( .A1(n9968), .A2(n9975), .B1(n9967), .B2(n9973), .ZN(n9970)
         );
  AOI211_X1 U11056 ( .C1(n9980), .C2(n9971), .A(n9970), .B(n9969), .ZN(n9986)
         );
  INV_X1 U11057 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9972) );
  AOI22_X1 U11058 ( .A1(n9983), .A2(n9986), .B1(n9972), .B2(n9981), .ZN(
        P1_U3472) );
  OAI22_X1 U11059 ( .A1(n9976), .A2(n9975), .B1(n9974), .B2(n9973), .ZN(n9978)
         );
  AOI211_X1 U11060 ( .C1(n9980), .C2(n9979), .A(n9978), .B(n9977), .ZN(n9989)
         );
  INV_X1 U11061 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9982) );
  AOI22_X1 U11062 ( .A1(n9983), .A2(n9989), .B1(n9982), .B2(n9981), .ZN(
        P1_U3478) );
  AOI22_X1 U11063 ( .A1(n9990), .A2(n9984), .B1(n6839), .B2(n9987), .ZN(
        P1_U3527) );
  AOI22_X1 U11064 ( .A1(n9990), .A2(n9986), .B1(n9985), .B2(n9987), .ZN(
        P1_U3529) );
  AOI22_X1 U11065 ( .A1(n9990), .A2(n9989), .B1(n9988), .B2(n9987), .ZN(
        P1_U3531) );
  XOR2_X1 U11066 ( .A(n9992), .B(n9991), .Z(n10003) );
  OAI21_X1 U11067 ( .B1(n9995), .B2(n9994), .A(n9993), .ZN(n9996) );
  AOI21_X1 U11068 ( .B1(n9998), .B2(n9997), .A(n9996), .ZN(n9999) );
  OAI21_X1 U11069 ( .B1(n10084), .B2(n10000), .A(n9999), .ZN(n10001) );
  AOI21_X1 U11070 ( .B1(n10003), .B2(n10002), .A(n10001), .ZN(n10004) );
  OAI21_X1 U11071 ( .B1(n10006), .B2(n10005), .A(n10004), .ZN(P2_U3223) );
  AOI22_X1 U11072 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n10008), .B1(n10007), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n10017) );
  NAND2_X1 U11073 ( .A1(n10008), .A2(n7333), .ZN(n10010) );
  OAI211_X1 U11074 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n10011), .A(n10010), .B(
        n10009), .ZN(n10012) );
  INV_X1 U11075 ( .A(n10012), .ZN(n10015) );
  AOI22_X1 U11076 ( .A1(n10013), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10014) );
  OAI221_X1 U11077 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n10017), .C1(n10016), .C2(
        n10015), .A(n10014), .ZN(P2_U3245) );
  NAND2_X1 U11078 ( .A1(n10019), .A2(n10018), .ZN(n10030) );
  INV_X1 U11079 ( .A(n10020), .ZN(n10028) );
  NAND2_X1 U11080 ( .A1(n10022), .A2(n10021), .ZN(n10023) );
  OAI21_X1 U11081 ( .B1(n10025), .B2(n10024), .A(n10023), .ZN(n10026) );
  AOI21_X1 U11082 ( .B1(n10028), .B2(n10027), .A(n10026), .ZN(n10029) );
  NAND2_X1 U11083 ( .A1(n10030), .A2(n10029), .ZN(n10031) );
  NOR2_X1 U11084 ( .A1(n10032), .A2(n10031), .ZN(n10033) );
  AOI22_X1 U11085 ( .A1(n9017), .A2(n5650), .B1(n10033), .B2(n9079), .ZN(
        P2_U3291) );
  AND2_X1 U11086 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10042), .ZN(P2_U3297) );
  AND2_X1 U11087 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10042), .ZN(P2_U3298) );
  AND2_X1 U11088 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10042), .ZN(P2_U3299) );
  AND2_X1 U11089 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10042), .ZN(P2_U3300) );
  AND2_X1 U11090 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10042), .ZN(P2_U3301) );
  AND2_X1 U11091 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10042), .ZN(P2_U3302) );
  NOR2_X1 U11092 ( .A1(n10039), .A2(n10036), .ZN(P2_U3303) );
  AND2_X1 U11093 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10042), .ZN(P2_U3304) );
  AND2_X1 U11094 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10042), .ZN(P2_U3305) );
  AND2_X1 U11095 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10042), .ZN(P2_U3306) );
  AND2_X1 U11096 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10042), .ZN(P2_U3307) );
  AND2_X1 U11097 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10042), .ZN(P2_U3308) );
  AND2_X1 U11098 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10042), .ZN(P2_U3309) );
  AND2_X1 U11099 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10042), .ZN(P2_U3310) );
  AND2_X1 U11100 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10042), .ZN(P2_U3311) );
  AND2_X1 U11101 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10042), .ZN(P2_U3312) );
  AND2_X1 U11102 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10042), .ZN(P2_U3313) );
  AND2_X1 U11103 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10042), .ZN(P2_U3314) );
  AND2_X1 U11104 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10042), .ZN(P2_U3315) );
  AND2_X1 U11105 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10042), .ZN(P2_U3316) );
  AND2_X1 U11106 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10042), .ZN(P2_U3317) );
  NOR2_X1 U11107 ( .A1(n10039), .A2(n10037), .ZN(P2_U3318) );
  AND2_X1 U11108 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10042), .ZN(P2_U3319) );
  AND2_X1 U11109 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10042), .ZN(P2_U3320) );
  NOR2_X1 U11110 ( .A1(n10039), .A2(n10038), .ZN(P2_U3321) );
  AND2_X1 U11111 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10042), .ZN(P2_U3322) );
  AND2_X1 U11112 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10042), .ZN(P2_U3323) );
  AND2_X1 U11113 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10042), .ZN(P2_U3324) );
  AND2_X1 U11114 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10042), .ZN(P2_U3325) );
  AND2_X1 U11115 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10042), .ZN(P2_U3326) );
  AOI22_X1 U11116 ( .A1(n10045), .A2(n10041), .B1(n10040), .B2(n10042), .ZN(
        P2_U3437) );
  AOI22_X1 U11117 ( .A1(n10045), .A2(n10044), .B1(n10043), .B2(n10042), .ZN(
        P2_U3438) );
  AOI22_X1 U11118 ( .A1(n10048), .A2(n10101), .B1(n10047), .B2(n10046), .ZN(
        n10049) );
  AND2_X1 U11119 ( .A1(n10050), .A2(n10049), .ZN(n10107) );
  AOI22_X1 U11120 ( .A1(n10105), .A2(n10107), .B1(n5592), .B2(n10103), .ZN(
        P2_U3451) );
  OAI21_X1 U11121 ( .B1(n10052), .B2(n10095), .A(n10051), .ZN(n10054) );
  AOI211_X1 U11122 ( .C1(n10101), .C2(n10055), .A(n10054), .B(n10053), .ZN(
        n10109) );
  INV_X1 U11123 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10056) );
  AOI22_X1 U11124 ( .A1(n10105), .A2(n10109), .B1(n10056), .B2(n10103), .ZN(
        P2_U3454) );
  OAI21_X1 U11125 ( .B1(n10058), .B2(n10095), .A(n10057), .ZN(n10060) );
  AOI211_X1 U11126 ( .C1(n10101), .C2(n10061), .A(n10060), .B(n10059), .ZN(
        n10111) );
  AOI22_X1 U11127 ( .A1(n10105), .A2(n10111), .B1(n5601), .B2(n10103), .ZN(
        P2_U3457) );
  OAI22_X1 U11128 ( .A1(n10063), .A2(n10097), .B1(n10062), .B2(n10095), .ZN(
        n10064) );
  INV_X1 U11129 ( .A(n10064), .ZN(n10067) );
  NAND2_X1 U11130 ( .A1(n10065), .A2(n10101), .ZN(n10066) );
  AND3_X1 U11131 ( .A1(n10068), .A2(n10067), .A3(n10066), .ZN(n10112) );
  AOI22_X1 U11132 ( .A1(n10105), .A2(n10112), .B1(n5623), .B2(n10103), .ZN(
        P2_U3460) );
  AND2_X1 U11133 ( .A1(n10069), .A2(n10101), .ZN(n10073) );
  OAI21_X1 U11134 ( .B1(n10071), .B2(n10095), .A(n10070), .ZN(n10072) );
  NOR3_X1 U11135 ( .A1(n10074), .A2(n10073), .A3(n10072), .ZN(n10113) );
  INV_X1 U11136 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10075) );
  AOI22_X1 U11137 ( .A1(n10105), .A2(n10113), .B1(n10075), .B2(n10103), .ZN(
        P2_U3463) );
  OAI22_X1 U11138 ( .A1(n10077), .A2(n10097), .B1(n10076), .B2(n10095), .ZN(
        n10079) );
  AOI211_X1 U11139 ( .C1(n10080), .C2(n10101), .A(n10079), .B(n10078), .ZN(
        n10114) );
  INV_X1 U11140 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10081) );
  AOI22_X1 U11141 ( .A1(n10105), .A2(n10114), .B1(n10081), .B2(n10103), .ZN(
        P2_U3469) );
  OAI211_X1 U11142 ( .C1(n10084), .C2(n10095), .A(n10083), .B(n10082), .ZN(
        n10085) );
  AOI21_X1 U11143 ( .B1(n10086), .B2(n10101), .A(n10085), .ZN(n10115) );
  AOI22_X1 U11144 ( .A1(n10105), .A2(n10115), .B1(n5717), .B2(n10103), .ZN(
        P2_U3475) );
  INV_X1 U11145 ( .A(n10087), .ZN(n10094) );
  INV_X1 U11146 ( .A(n10088), .ZN(n10093) );
  OAI22_X1 U11147 ( .A1(n10090), .A2(n10097), .B1(n10089), .B2(n10095), .ZN(
        n10092) );
  AOI211_X1 U11148 ( .C1(n10094), .C2(n10093), .A(n10092), .B(n10091), .ZN(
        n10116) );
  AOI22_X1 U11149 ( .A1(n10105), .A2(n10116), .B1(n5755), .B2(n10103), .ZN(
        P2_U3481) );
  OAI22_X1 U11150 ( .A1(n10098), .A2(n10097), .B1(n10096), .B2(n10095), .ZN(
        n10100) );
  AOI211_X1 U11151 ( .C1(n10102), .C2(n10101), .A(n10100), .B(n10099), .ZN(
        n10118) );
  INV_X1 U11152 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10104) );
  AOI22_X1 U11153 ( .A1(n10105), .A2(n10118), .B1(n10104), .B2(n10103), .ZN(
        P2_U3487) );
  AOI22_X1 U11154 ( .A1(n10119), .A2(n10107), .B1(n10106), .B2(n10117), .ZN(
        P2_U3520) );
  AOI22_X1 U11155 ( .A1(n10119), .A2(n10109), .B1(n10108), .B2(n10117), .ZN(
        P2_U3521) );
  AOI22_X1 U11156 ( .A1(n10119), .A2(n10111), .B1(n10110), .B2(n10117), .ZN(
        P2_U3522) );
  AOI22_X1 U11157 ( .A1(n10119), .A2(n10112), .B1(n7050), .B2(n10117), .ZN(
        P2_U3523) );
  AOI22_X1 U11158 ( .A1(n10119), .A2(n10113), .B1(n7048), .B2(n10117), .ZN(
        P2_U3524) );
  AOI22_X1 U11159 ( .A1(n10119), .A2(n10114), .B1(n7094), .B2(n10117), .ZN(
        P2_U3526) );
  AOI22_X1 U11160 ( .A1(n10119), .A2(n10115), .B1(n5716), .B2(n10117), .ZN(
        P2_U3528) );
  AOI22_X1 U11161 ( .A1(n10119), .A2(n10116), .B1(n7269), .B2(n10117), .ZN(
        P2_U3530) );
  AOI22_X1 U11162 ( .A1(n10119), .A2(n10118), .B1(n7523), .B2(n10117), .ZN(
        P2_U3532) );
  INV_X1 U11163 ( .A(n10120), .ZN(n10121) );
  NAND2_X1 U11164 ( .A1(n10122), .A2(n10121), .ZN(n10123) );
  XOR2_X1 U11165 ( .A(n10124), .B(n10123), .Z(ADD_1071_U5) );
  XOR2_X1 U11166 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11167 ( .B1(n10127), .B2(n10126), .A(n10125), .ZN(ADD_1071_U56) );
  OAI21_X1 U11168 ( .B1(n10130), .B2(n10129), .A(n10128), .ZN(ADD_1071_U57) );
  OAI21_X1 U11169 ( .B1(n10133), .B2(n10132), .A(n10131), .ZN(ADD_1071_U58) );
  OAI21_X1 U11170 ( .B1(n10136), .B2(n10135), .A(n10134), .ZN(ADD_1071_U59) );
  OAI21_X1 U11171 ( .B1(n10139), .B2(n10138), .A(n10137), .ZN(ADD_1071_U60) );
  OAI21_X1 U11172 ( .B1(n10142), .B2(n10141), .A(n10140), .ZN(ADD_1071_U61) );
  AOI21_X1 U11173 ( .B1(n10145), .B2(n10144), .A(n10143), .ZN(ADD_1071_U62) );
  AOI21_X1 U11174 ( .B1(n10148), .B2(n10147), .A(n10146), .ZN(ADD_1071_U63) );
  XOR2_X1 U11175 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10149), .Z(ADD_1071_U49) );
  NOR2_X1 U11176 ( .A1(n10151), .A2(n10150), .ZN(n10152) );
  XOR2_X1 U11177 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10152), .Z(ADD_1071_U51) );
  XOR2_X1 U11178 ( .A(n10153), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  OAI21_X1 U11179 ( .B1(n10156), .B2(n10155), .A(n10154), .ZN(n10157) );
  XNOR2_X1 U11180 ( .A(n10157), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  XOR2_X1 U11181 ( .A(n10158), .B(P2_ADDR_REG_8__SCAN_IN), .Z(ADD_1071_U48) );
  AOI21_X1 U11182 ( .B1(n10161), .B2(n10160), .A(n10159), .ZN(ADD_1071_U47) );
  XOR2_X1 U11183 ( .A(n10163), .B(n10162), .Z(ADD_1071_U54) );
  XOR2_X1 U11184 ( .A(n10165), .B(n10164), .Z(ADD_1071_U53) );
  XNOR2_X1 U11185 ( .A(n10167), .B(n10166), .ZN(ADD_1071_U52) );
  NOR2_X1 U10147 ( .A1(n9058), .A2(n9146), .ZN(n9037) );
  INV_X1 U4818 ( .A(n6372), .ZN(n4453) );
  CLKBUF_X1 U4834 ( .A(n5684), .Z(n5917) );
  CLKBUF_X1 U4938 ( .A(n5707), .Z(n5805) );
  CLKBUF_X1 U5192 ( .A(n8324), .Z(n4388) );
  CLKBUF_X2 U5193 ( .A(n6196), .Z(n7336) );
  CLKBUF_X1 U5723 ( .A(n5559), .Z(n9207) );
  CLKBUF_X1 U6084 ( .A(n6851), .Z(n4313) );
endmodule

