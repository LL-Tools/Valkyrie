

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput63, keyinput62, keyinput61, keyinput60, keyinput59, keyinput58, 
        keyinput57, keyinput56, keyinput55, keyinput54, keyinput53, keyinput52, 
        keyinput51, keyinput50, keyinput49, keyinput48, keyinput47, keyinput46, 
        keyinput45, keyinput44, keyinput43, keyinput42, keyinput41, keyinput40, 
        keyinput39, keyinput38, keyinput37, keyinput36, keyinput35, keyinput34, 
        keyinput33, keyinput32, keyinput31, keyinput30, keyinput29, keyinput28, 
        keyinput27, keyinput26, keyinput25, keyinput24, keyinput23, keyinput22, 
        keyinput21, keyinput20, keyinput19, keyinput18, keyinput17, keyinput16, 
        keyinput15, keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, 
        keyinput9, keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, 
        keyinput3, keyinput2, keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040;

  AND4_X1 U4756 ( .A1(n4917), .A2(n4916), .A3(n4915), .A4(n4914), .ZN(n7144)
         );
  INV_X1 U4757 ( .A(n5961), .ZN(n6235) );
  CLKBUF_X2 U4758 ( .A(n6143), .Z(n4259) );
  BUF_X1 U4759 ( .A(n5960), .Z(n8646) );
  BUF_X2 U4760 ( .A(n5611), .Z(n4266) );
  AND2_X1 U4761 ( .A1(n9494), .A2(n9498), .ZN(n5657) );
  NAND2_X2 U4762 ( .A1(n6243), .A2(n6526), .ZN(n5602) );
  INV_X1 U4763 ( .A(n8561), .ZN(n4252) );
  BUF_X1 U4764 ( .A(n5648), .Z(n6133) );
  AND2_X1 U4765 ( .A1(n5523), .A2(n5522), .ZN(n5821) );
  INV_X1 U4766 ( .A(n6650), .ZN(n6655) );
  BUF_X1 U4767 ( .A(n5602), .Z(n6289) );
  INV_X1 U4768 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5818) );
  INV_X1 U4769 ( .A(n7615), .ZN(n5408) );
  INV_X1 U4770 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5169) );
  BUF_X2 U4771 ( .A(n8552), .Z(n4264) );
  AND2_X1 U4772 ( .A1(n5539), .A2(n5538), .ZN(n5635) );
  NAND2_X1 U4773 ( .A1(n9447), .A2(n8895), .ZN(n8917) );
  NAND2_X1 U4774 ( .A1(n5535), .A2(n5536), .ZN(n5538) );
  OAI22_X1 U4775 ( .A1(n7529), .A2(n7528), .B1(n7428), .B2(n8015), .ZN(n7480)
         );
  INV_X1 U4776 ( .A(n5006), .ZN(n5387) );
  NAND2_X1 U4777 ( .A1(n5700), .A2(n5699), .ZN(n8458) );
  XNOR2_X1 U4778 ( .A(n5537), .B(P1_IR_REG_30__SCAN_IN), .ZN(n9494) );
  INV_X1 U4779 ( .A(n4864), .ZN(n6274) );
  INV_X1 U4780 ( .A(n7938), .ZN(n7962) );
  INV_X1 U4781 ( .A(n8098), .ZN(n9907) );
  INV_X1 U4782 ( .A(n8646), .ZN(n9016) );
  NAND2_X1 U4784 ( .A1(n8302), .A2(n8367), .ZN(n6067) );
  NAND2_X2 U4785 ( .A1(n8282), .A2(n6130), .ZN(n6176) );
  NAND2_X2 U4786 ( .A1(n6260), .A2(n6103), .ZN(n8282) );
  XNOR2_X2 U4787 ( .A(n4861), .B(n4860), .ZN(n6396) );
  NAND4_X2 U4788 ( .A1(n4856), .A2(n4855), .A3(n4854), .A4(n4853), .ZN(n4867)
         );
  BUF_X2 U4789 ( .A(n9715), .Z(n4250) );
  XNOR2_X1 U4790 ( .A(n4882), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9715) );
  NAND2_X2 U4791 ( .A1(n6047), .A2(n8300), .ZN(n8302) );
  NOR2_X2 U4792 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5522) );
  AOI21_X2 U4793 ( .B1(n7521), .B2(n7522), .A(n7438), .ZN(n7498) );
  OAI22_X2 U4794 ( .A1(n7455), .A2(n8000), .B1(n7436), .B2(n7435), .ZN(n7521)
         );
  XNOR2_X2 U4795 ( .A(n4477), .B(n4476), .ZN(n8739) );
  NAND2_X1 U4796 ( .A1(n6067), .A2(n8365), .ZN(n8364) );
  XNOR2_X2 U4797 ( .A(n5563), .B(P1_IR_REG_21__SCAN_IN), .ZN(n8645) );
  NAND4_X2 U4798 ( .A1(n5639), .A2(n5638), .A3(n5637), .A4(n5636), .ZN(n8734)
         );
  NAND2_X2 U4799 ( .A1(n8312), .A2(n8313), .ZN(n8311) );
  AND2_X2 U4800 ( .A1(n5792), .A2(n5791), .ZN(n5793) );
  OAI211_X1 U4801 ( .C1(n8716), .C2(n6172), .A(n6191), .B(n6701), .ZN(n5589)
         );
  NAND2_X1 U4802 ( .A1(n9340), .A2(n8902), .ZN(n8922) );
  OAI21_X1 U4803 ( .B1(n5225), .B2(n4725), .A(n4722), .ZN(n5258) );
  NAND2_X1 U4804 ( .A1(n4541), .A2(n5741), .ZN(n6942) );
  INV_X2 U4805 ( .A(n9306), .ZN(n4251) );
  NAND2_X1 U4806 ( .A1(n7670), .A2(n7665), .ZN(n5413) );
  INV_X1 U4807 ( .A(n6143), .ZN(n5611) );
  CLKBUF_X2 U4808 ( .A(n6434), .Z(n4370) );
  INV_X2 U4809 ( .A(n9669), .ZN(n6774) );
  INV_X1 U4810 ( .A(n7832), .ZN(n4891) );
  INV_X2 U4811 ( .A(n4867), .ZN(n8165) );
  OAI211_X1 U4812 ( .C1(n6299), .C2(n5640), .A(n5586), .B(n5585), .ZN(n6414)
         );
  BUF_X2 U4813 ( .A(n5641), .Z(n5961) );
  BUF_X1 U4814 ( .A(n4931), .Z(n4262) );
  NOR2_X2 U4815 ( .A1(n6180), .A2(n6526), .ZN(n9224) );
  AND2_X1 U4816 ( .A1(n7394), .A2(n4852), .ZN(n4931) );
  INV_X1 U4817 ( .A(n7615), .ZN(n4849) );
  INV_X2 U4818 ( .A(n4639), .ZN(n7812) );
  NAND2_X4 U4819 ( .A1(n4737), .A2(n4738), .ZN(n4879) );
  NAND2_X1 U4820 ( .A1(n8364), .A2(n6068), .ZN(n8338) );
  MUX2_X1 U4821 ( .A(n8113), .B(n8187), .S(n9982), .Z(n8114) );
  MUX2_X1 U4822 ( .A(n8188), .B(n8187), .S(n9967), .Z(n8189) );
  AND2_X1 U4823 ( .A1(n8112), .A2(n8111), .ZN(n8187) );
  INV_X1 U4824 ( .A(n4543), .ZN(n7594) );
  NAND2_X1 U4825 ( .A1(n6012), .A2(n6011), .ZN(n9452) );
  AND2_X1 U4826 ( .A1(n5223), .A2(n7757), .ZN(n8032) );
  NAND2_X1 U4827 ( .A1(n5232), .A2(n5231), .ZN(n8231) );
  OR2_X1 U4828 ( .A1(n9851), .A2(n9850), .ZN(n4586) );
  NAND2_X1 U4829 ( .A1(n5964), .A2(n5963), .ZN(n9372) );
  NAND2_X1 U4830 ( .A1(n5214), .A2(n5213), .ZN(n8237) );
  NAND2_X1 U4831 ( .A1(n5191), .A2(n5190), .ZN(n8243) );
  AND3_X1 U4832 ( .A1(n4599), .A2(n4597), .A3(n4601), .ZN(n7905) );
  NAND2_X1 U4833 ( .A1(n7287), .A2(n7288), .ZN(n7342) );
  OR2_X1 U4834 ( .A1(n9819), .A2(n4600), .ZN(n4599) );
  NAND2_X1 U4835 ( .A1(n5920), .A2(n5919), .ZN(n9385) );
  NAND2_X1 U4836 ( .A1(n7102), .A2(n4582), .ZN(n7181) );
  NAND2_X1 U4837 ( .A1(n6664), .A2(n6663), .ZN(n6948) );
  NAND2_X1 U4838 ( .A1(n5827), .A2(n5826), .ZN(n7175) );
  NAND2_X1 U4839 ( .A1(n5076), .A2(n5075), .ZN(n9965) );
  NAND2_X1 U4840 ( .A1(n5037), .A2(n5036), .ZN(n9947) );
  NAND2_X1 U4841 ( .A1(n4502), .A2(n5063), .ZN(n9959) );
  NAND2_X1 U4842 ( .A1(n5798), .A2(n5797), .ZN(n7110) );
  OAI21_X1 U4843 ( .B1(n7085), .B2(n7084), .A(n5418), .ZN(n7090) );
  NAND2_X1 U4844 ( .A1(n5757), .A2(n5756), .ZN(n6919) );
  NAND2_X1 U4845 ( .A1(n5719), .A2(n5718), .ZN(n9676) );
  AND2_X1 U4846 ( .A1(n7129), .A2(n7695), .ZN(n7633) );
  NAND2_X1 U4847 ( .A1(n9306), .A2(n6686), .ZN(n9315) );
  NAND2_X1 U4848 ( .A1(n7667), .A2(n4872), .ZN(n6618) );
  AND2_X1 U4849 ( .A1(n7681), .A2(n7694), .ZN(n7678) );
  NAND2_X2 U4850 ( .A1(n6683), .A2(n9257), .ZN(n9306) );
  INV_X1 U4851 ( .A(n5413), .ZN(n7667) );
  AND4_X1 U4852 ( .A1(n4870), .A2(n4831), .A3(n4869), .A4(n4868), .ZN(n6721)
         );
  NAND2_X1 U4853 ( .A1(n4949), .A2(n4948), .ZN(n4962) );
  CLKBUF_X1 U4854 ( .A(n6172), .Z(n8707) );
  AND2_X1 U4855 ( .A1(n6337), .A2(n6338), .ZN(n5574) );
  BUF_X2 U4856 ( .A(n4931), .Z(n4261) );
  INV_X2 U4857 ( .A(n4908), .ZN(n5249) );
  AND2_X1 U4859 ( .A1(n4478), .A2(n4720), .ZN(n4483) );
  AND2_X2 U4860 ( .A1(n6272), .A2(n6271), .ZN(P1_U3973) );
  XNOR2_X1 U4861 ( .A(n5460), .B(n9089), .ZN(n7393) );
  INV_X2 U4862 ( .A(n5590), .ZN(n4253) );
  NAND2_X2 U4863 ( .A1(n4851), .A2(n4852), .ZN(n4913) );
  INV_X1 U4864 ( .A(n5538), .ZN(n9498) );
  INV_X1 U4865 ( .A(n4851), .ZN(n7394) );
  NAND2_X2 U4866 ( .A1(n8278), .A2(n4851), .ZN(n7615) );
  OR3_X1 U4867 ( .A1(n5851), .A2(n5850), .A3(n5849), .ZN(n5872) );
  NAND2_X1 U4868 ( .A1(n5463), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5460) );
  INV_X1 U4869 ( .A(n6338), .ZN(n8712) );
  INV_X1 U4870 ( .A(n4852), .ZN(n8278) );
  NAND2_X1 U4871 ( .A1(n5940), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5571) );
  NAND2_X1 U4872 ( .A1(n5581), .A2(n5584), .ZN(n6526) );
  NAND3_X1 U4873 ( .A1(n5560), .A2(n6150), .A3(n5551), .ZN(n6191) );
  MUX2_X1 U4874 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5534), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5535) );
  NAND2_X1 U4875 ( .A1(n5536), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5537) );
  XNOR2_X1 U4876 ( .A(n5547), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6150) );
  OR2_X1 U4877 ( .A1(n8269), .A2(n5169), .ZN(n4848) );
  NAND2_X1 U4878 ( .A1(n5568), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5938) );
  NAND2_X1 U4879 ( .A1(n4289), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4858) );
  NAND2_X1 U4880 ( .A1(n5550), .A2(n5549), .ZN(n7310) );
  NAND2_X1 U4881 ( .A1(n5549), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5547) );
  XNOR2_X1 U4882 ( .A(n6166), .B(P1_IR_REG_22__SCAN_IN), .ZN(n8716) );
  OAI21_X1 U4883 ( .B1(n5399), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5487) );
  NAND2_X1 U4884 ( .A1(n4288), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6166) );
  OR2_X1 U4885 ( .A1(n5399), .A2(n4316), .ZN(n4270) );
  OAI21_X1 U4886 ( .B1(n4288), .B2(n5555), .A(n4278), .ZN(n5559) );
  NAND2_X2 U4887 ( .A1(n6281), .A2(P1_U3086), .ZN(n9500) );
  OR2_X1 U4888 ( .A1(n5564), .A2(n5554), .ZN(n4288) );
  NAND2_X1 U4889 ( .A1(n4798), .A2(n4846), .ZN(n4797) );
  AND3_X1 U4890 ( .A1(n4393), .A2(n4840), .A3(n4838), .ZN(n4826) );
  AND2_X1 U4891 ( .A1(n4819), .A2(n4959), .ZN(n4274) );
  AND4_X1 U4892 ( .A1(n5530), .A2(n5529), .A3(n5528), .A4(n5527), .ZN(n4825)
         );
  NAND2_X1 U4893 ( .A1(n4732), .A2(n4735), .ZN(n4737) );
  AND3_X1 U4894 ( .A1(n5526), .A2(n5569), .A3(n6168), .ZN(n5530) );
  AND2_X1 U4895 ( .A1(n4942), .A2(n4919), .ZN(n4819) );
  AND3_X1 U4896 ( .A1(n5059), .A2(n4836), .A3(n4835), .ZN(n4840) );
  AND2_X1 U4897 ( .A1(n5545), .A2(n5531), .ZN(n5576) );
  INV_X1 U4898 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5397) );
  INV_X1 U4899 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5059) );
  INV_X1 U4900 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5865) );
  INV_X1 U4901 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5545) );
  INV_X1 U4902 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5569) );
  INV_X1 U4903 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4833) );
  INV_X1 U4904 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5817) );
  INV_X1 U4905 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5917) );
  INV_X1 U4906 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n9089) );
  INV_X1 U4907 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n4942) );
  INV_X1 U4908 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6168) );
  INV_X1 U4909 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5486) );
  AND2_X1 U4910 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n4732) );
  INV_X1 U4911 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4735) );
  INV_X4 U4912 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U4913 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4528) );
  AOI21_X2 U4914 ( .B1(n8033), .B2(n8032), .A(n7657), .ZN(n8021) );
  NAND2_X4 U4915 ( .A1(n7811), .A2(n4639), .ZN(n4864) );
  NOR2_X2 U4916 ( .A1(n4270), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n8269) );
  NAND2_X1 U4917 ( .A1(n6067), .A2(n4257), .ZN(n4254) );
  AND2_X2 U4918 ( .A1(n4254), .A2(n4255), .ZN(n6260) );
  OR2_X1 U4919 ( .A1(n4256), .A2(n6068), .ZN(n4255) );
  INV_X1 U4920 ( .A(n8339), .ZN(n4256) );
  AND2_X1 U4921 ( .A1(n8365), .A2(n8339), .ZN(n4257) );
  NAND2_X1 U4922 ( .A1(n8402), .A2(n5632), .ZN(n8312) );
  NAND2_X1 U4923 ( .A1(n8403), .A2(n8404), .ZN(n8402) );
  BUF_X2 U4924 ( .A(n6133), .Z(n6022) );
  AND4_X4 U4925 ( .A1(n5822), .A2(n5525), .A3(n5524), .A4(n5821), .ZN(n4258)
         );
  INV_X1 U4926 ( .A(n4258), .ZN(n5567) );
  NAND2_X1 U4927 ( .A1(n5574), .A2(n6191), .ZN(n6143) );
  OR2_X2 U4928 ( .A1(n5571), .A2(n5570), .ZN(n5573) );
  AOI211_X1 U4929 ( .C1(n6423), .C2(n6422), .A(n8424), .B(n6421), .ZN(n6426)
         );
  NAND2_X1 U4930 ( .A1(n5574), .A2(n6191), .ZN(n4260) );
  INV_X2 U4931 ( .A(n4253), .ZN(n6080) );
  XNOR2_X1 U4932 ( .A(n5669), .B(n4266), .ZN(n5671) );
  INV_X1 U4933 ( .A(n5589), .ZN(n6145) );
  NAND4_X2 U4934 ( .A1(n5707), .A2(n5706), .A3(n5705), .A4(n5704), .ZN(n8731)
         );
  NAND2_X1 U4935 ( .A1(n5771), .A2(n5770), .ZN(n7020) );
  XNOR2_X1 U4936 ( .A(n5566), .B(n5565), .ZN(n7070) );
  AND2_X2 U4937 ( .A1(n5539), .A2(n9498), .ZN(n8552) );
  AND2_X1 U4938 ( .A1(n4487), .A2(n4828), .ZN(n4486) );
  OR2_X1 U4939 ( .A1(n7654), .A2(n7655), .ZN(n7800) );
  OR2_X1 U4940 ( .A1(n9965), .A2(n7413), .ZN(n7723) );
  INV_X1 U4941 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n4841) );
  NOR2_X1 U4942 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n4842) );
  NAND2_X1 U4943 ( .A1(n4709), .A2(n4707), .ZN(n5367) );
  AOI21_X1 U4944 ( .B1(n4711), .B2(n4713), .A(n4708), .ZN(n4707) );
  NAND2_X1 U4945 ( .A1(n5331), .A2(n4711), .ZN(n4709) );
  INV_X1 U4946 ( .A(n5349), .ZN(n4708) );
  AOI21_X1 U4947 ( .B1(n4550), .B2(n7409), .A(n4326), .ZN(n4548) );
  NAND2_X1 U4949 ( .A1(n4412), .A2(n7721), .ZN(n7731) );
  NAND2_X1 U4950 ( .A1(n4414), .A2(n4413), .ZN(n4412) );
  INV_X1 U4951 ( .A(n7722), .ZN(n4413) );
  OAI21_X1 U4952 ( .B1(n8513), .B2(n8677), .A(n8680), .ZN(n8510) );
  NAND2_X1 U4953 ( .A1(n4388), .A2(n4309), .ZN(n4387) );
  NAND2_X1 U4954 ( .A1(n4390), .A2(n4389), .ZN(n4388) );
  OAI21_X1 U4955 ( .B1(n4320), .B2(n7781), .A(n4397), .ZN(n7764) );
  NAND2_X1 U4956 ( .A1(n7762), .A2(n7781), .ZN(n4397) );
  NAND2_X1 U4957 ( .A1(n4400), .A2(n4399), .ZN(n7761) );
  INV_X1 U4958 ( .A(n7767), .ZN(n4396) );
  NAND2_X1 U4959 ( .A1(n7769), .A2(n4497), .ZN(n4496) );
  NOR2_X1 U4960 ( .A1(n7801), .A2(n7626), .ZN(n4497) );
  NAND2_X1 U4961 ( .A1(n7774), .A2(n4499), .ZN(n4498) );
  AND2_X1 U4962 ( .A1(n7773), .A2(n7801), .ZN(n4499) );
  AND2_X1 U4963 ( .A1(n4727), .A2(n5240), .ZN(n4726) );
  NAND2_X1 U4964 ( .A1(n5224), .A2(n5226), .ZN(n4727) );
  NAND2_X1 U4965 ( .A1(n5011), .A2(n5010), .ZN(n4487) );
  NOR2_X1 U4966 ( .A1(n5050), .A2(n4721), .ZN(n4720) );
  INV_X1 U4967 ( .A(n5029), .ZN(n4721) );
  NOR2_X1 U4968 ( .A1(n5016), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5057) );
  AND2_X1 U4969 ( .A1(n4786), .A2(n4328), .ZN(n4784) );
  INV_X1 U4970 ( .A(n4296), .ZN(n4777) );
  NAND2_X1 U4971 ( .A1(n4772), .A2(n5414), .ZN(n8160) );
  OR2_X1 U4972 ( .A1(n7991), .A2(n7550), .ZN(n7768) );
  OR2_X1 U4973 ( .A1(n8225), .A2(n7430), .ZN(n7759) );
  OR2_X1 U4974 ( .A1(n7804), .A2(n6643), .ZN(n7652) );
  INV_X1 U4975 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5459) );
  NAND2_X1 U4976 ( .A1(n5816), .A2(n7159), .ZN(n4753) );
  NOR2_X1 U4977 ( .A1(n8954), .A2(n9427), .ZN(n8938) );
  NOR2_X1 U4978 ( .A1(n9676), .A2(n6939), .ZN(n8463) );
  AND2_X1 U4979 ( .A1(n4668), .A2(n4300), .ZN(n4667) );
  NOR2_X1 U4980 ( .A1(n4674), .A2(n8899), .ZN(n4671) );
  NAND2_X1 U4981 ( .A1(n4690), .A2(n4689), .ZN(n4688) );
  NAND2_X1 U4982 ( .A1(n5313), .A2(n5312), .ZN(n5331) );
  OAI21_X1 U4983 ( .B1(n5258), .B2(n5257), .A(n5256), .ZN(n5274) );
  NAND2_X1 U4984 ( .A1(n5164), .A2(n5163), .ZN(n5187) );
  AOI21_X1 U4985 ( .B1(n4717), .B2(n4277), .A(n4322), .ZN(n4716) );
  OR2_X1 U4986 ( .A1(n5738), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5776) );
  NAND2_X1 U4987 ( .A1(n4701), .A2(n5001), .ZN(n5012) );
  AND3_X1 U4988 ( .A1(n4885), .A2(n4884), .A3(n4883), .ZN(n8171) );
  INV_X1 U4989 ( .A(n4553), .ZN(n4551) );
  OR2_X1 U4990 ( .A1(n7806), .A2(n7805), .ZN(n4419) );
  NAND2_X1 U4991 ( .A1(n6488), .A2(n6489), .ZN(n6609) );
  XNOR2_X1 U4992 ( .A(n6840), .B(n6847), .ZN(n6839) );
  NAND2_X1 U4993 ( .A1(n4289), .A2(n4859), .ZN(n4639) );
  NAND2_X1 U4994 ( .A1(n4454), .A2(n4310), .ZN(n4859) );
  NAND2_X1 U4995 ( .A1(n5402), .A2(n4452), .ZN(n4454) );
  OR2_X1 U4996 ( .A1(n9835), .A2(n5098), .ZN(n4600) );
  NAND2_X1 U4997 ( .A1(n7902), .A2(n4598), .ZN(n4597) );
  INV_X1 U4998 ( .A(n9835), .ZN(n4598) );
  OR2_X1 U4999 ( .A1(n5339), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5359) );
  NAND2_X1 U5000 ( .A1(n7313), .A2(n5431), .ZN(n4637) );
  INV_X1 U5001 ( .A(n7627), .ZN(n5431) );
  NOR2_X1 U5002 ( .A1(n4303), .A2(n4794), .ZN(n4793) );
  XNOR2_X1 U5003 ( .A(n9959), .B(n4501), .ZN(n7627) );
  NAND2_X1 U5004 ( .A1(n6206), .A2(n5493), .ZN(n5495) );
  AND2_X1 U5005 ( .A1(n5492), .A2(n5491), .ZN(n5493) );
  AND2_X1 U5006 ( .A1(n4829), .A2(n5446), .ZN(n4811) );
  AOI21_X1 U5007 ( .B1(n4269), .B2(n4619), .A(n4610), .ZN(n4609) );
  INV_X1 U5008 ( .A(n7742), .ZN(n4610) );
  INV_X1 U5009 ( .A(n7609), .ZN(n7606) );
  INV_X1 U5010 ( .A(n8092), .ZN(n8164) );
  NAND2_X1 U5011 ( .A1(n7924), .A2(n7801), .ZN(n8080) );
  NAND2_X1 U5012 ( .A1(n7605), .A2(n5507), .ZN(n8167) );
  NAND2_X1 U5013 ( .A1(n4270), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4847) );
  CLKBUF_X1 U5014 ( .A(n5401), .Z(n5402) );
  NAND2_X1 U5015 ( .A1(n4765), .A2(n4763), .ZN(n8374) );
  NOR2_X1 U5016 ( .A1(n8377), .A2(n4764), .ZN(n4763) );
  INV_X1 U5017 ( .A(n4822), .ZN(n4764) );
  NAND2_X1 U5018 ( .A1(n5602), .A2(n6276), .ZN(n5641) );
  AND2_X1 U5019 ( .A1(n8716), .A2(n8645), .ZN(n8640) );
  INV_X1 U5020 ( .A(n6134), .ZN(n6111) );
  NOR2_X1 U5021 ( .A1(n4655), .A2(n8909), .ZN(n4654) );
  INV_X1 U5022 ( .A(n8906), .ZN(n4655) );
  NAND2_X1 U5023 ( .A1(n6029), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6051) );
  INV_X1 U5024 ( .A(n4659), .ZN(n4658) );
  OAI21_X1 U5025 ( .B1(n7115), .B2(n4662), .A(n4660), .ZN(n4659) );
  INV_X1 U5026 ( .A(n7203), .ZN(n4660) );
  NAND2_X1 U5027 ( .A1(n4529), .A2(n9301), .ZN(n4534) );
  NOR2_X1 U5028 ( .A1(n8896), .A2(n4677), .ZN(n4676) );
  INV_X1 U5029 ( .A(n8893), .ZN(n4677) );
  OR2_X1 U5030 ( .A1(n9452), .A2(n8892), .ZN(n8893) );
  INV_X1 U5031 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4770) );
  NOR2_X1 U5032 ( .A1(n6383), .A2(n6384), .ZN(n6474) );
  NAND2_X1 U5033 ( .A1(n6227), .A2(n6226), .ZN(n9417) );
  MUX2_X1 U5034 ( .A(n8471), .B(n8470), .S(n8561), .Z(n8472) );
  OAI21_X1 U5035 ( .B1(n7732), .B2(n4392), .A(n4391), .ZN(n4390) );
  AND2_X1 U5036 ( .A1(n7733), .A2(n7734), .ZN(n4392) );
  NAND2_X1 U5037 ( .A1(n7736), .A2(n7735), .ZN(n4391) );
  NOR2_X1 U5038 ( .A1(n4411), .A2(n4406), .ZN(n4405) );
  AND2_X1 U5039 ( .A1(n7752), .A2(n7751), .ZN(n4411) );
  INV_X1 U5040 ( .A(n4408), .ZN(n4406) );
  AND2_X1 U5041 ( .A1(n7752), .A2(n7801), .ZN(n4500) );
  NAND2_X1 U5042 ( .A1(n8441), .A2(n8440), .ZN(n8443) );
  NOR2_X1 U5043 ( .A1(n8439), .A2(n4252), .ZN(n8440) );
  NAND2_X1 U5044 ( .A1(n8438), .A2(n8613), .ZN(n8441) );
  NAND2_X1 U5045 ( .A1(n8608), .A2(n4252), .ZN(n8442) );
  AND3_X1 U5046 ( .A1(n4376), .A2(n4375), .A3(n9161), .ZN(n8526) );
  AND2_X1 U5047 ( .A1(n4403), .A2(n4329), .ZN(n4401) );
  NAND2_X1 U5048 ( .A1(n4387), .A2(n4385), .ZN(n7748) );
  NOR2_X1 U5049 ( .A1(n4386), .A2(n7741), .ZN(n4385) );
  NAND2_X1 U5050 ( .A1(n4394), .A2(n7983), .ZN(n7772) );
  NAND2_X1 U5051 ( .A1(n4398), .A2(n4395), .ZN(n4394) );
  OAI21_X1 U5052 ( .B1(n7764), .B2(n4315), .A(n4396), .ZN(n4395) );
  INV_X1 U5053 ( .A(n7790), .ZN(n4492) );
  OAI21_X1 U5054 ( .B1(n4295), .B2(n4364), .A(n8561), .ZN(n8546) );
  OAI21_X1 U5055 ( .B1(n4537), .B2(n4431), .A(n8921), .ZN(n4430) );
  INV_X1 U5056 ( .A(n8922), .ZN(n4428) );
  INV_X1 U5057 ( .A(n4712), .ZN(n4711) );
  OAI21_X1 U5058 ( .B1(n5330), .B2(n4713), .A(n5347), .ZN(n4712) );
  INV_X1 U5059 ( .A(n4579), .ZN(n4578) );
  AOI21_X1 U5060 ( .B1(n4579), .B2(n4577), .A(n7568), .ZN(n4576) );
  INV_X1 U5061 ( .A(n7506), .ZN(n4577) );
  NOR2_X1 U5062 ( .A1(n7650), .A2(n4741), .ZN(n4740) );
  NAND2_X1 U5063 ( .A1(n4743), .A2(n4742), .ZN(n4741) );
  NOR2_X1 U5064 ( .A1(n7941), .A2(n4744), .ZN(n4743) );
  NAND2_X1 U5065 ( .A1(n4746), .A2(n4745), .ZN(n4744) );
  NAND2_X1 U5066 ( .A1(n9748), .A2(n4372), .ZN(n7850) );
  OR2_X1 U5067 ( .A1(n9743), .A2(n4990), .ZN(n4372) );
  INV_X1 U5068 ( .A(n9804), .ZN(n4591) );
  NAND2_X1 U5069 ( .A1(n4591), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4589) );
  AOI21_X1 U5070 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n7900), .A(n9803), .ZN(
        n7901) );
  NOR2_X1 U5071 ( .A1(n9866), .A2(n4583), .ZN(n7908) );
  NOR2_X1 U5072 ( .A1(n9857), .A2(n8073), .ZN(n4583) );
  NAND2_X1 U5073 ( .A1(n4635), .A2(n7786), .ZN(n4634) );
  INV_X1 U5074 ( .A(n5346), .ZN(n4635) );
  INV_X1 U5075 ( .A(n7776), .ZN(n4631) );
  AND2_X1 U5076 ( .A1(n4787), .A2(n4792), .ZN(n4786) );
  OR2_X1 U5077 ( .A1(n7940), .A2(n7821), .ZN(n4792) );
  OR2_X1 U5078 ( .A1(n5453), .A2(n4788), .ZN(n4787) );
  NAND2_X1 U5079 ( .A1(n5452), .A2(n5451), .ZN(n4788) );
  INV_X1 U5080 ( .A(n5451), .ZN(n4789) );
  OR2_X1 U5081 ( .A1(n8250), .A2(n8081), .ZN(n7745) );
  NAND2_X1 U5082 ( .A1(n5135), .A2(n5134), .ZN(n5152) );
  INV_X1 U5083 ( .A(n5136), .ZN(n5135) );
  NAND2_X1 U5084 ( .A1(n4290), .A2(n7711), .ZN(n4626) );
  NAND2_X1 U5085 ( .A1(n6722), .A2(n4867), .ZN(n7670) );
  NAND2_X1 U5086 ( .A1(n8174), .A2(n8165), .ZN(n7665) );
  OR2_X1 U5087 ( .A1(n7949), .A2(n8201), .ZN(n7776) );
  OR2_X1 U5088 ( .A1(n8207), .A2(n7986), .ZN(n7773) );
  NAND2_X1 U5089 ( .A1(n5441), .A2(n4817), .ZN(n4814) );
  OR2_X1 U5090 ( .A1(n8231), .A2(n8041), .ZN(n7758) );
  OR2_X1 U5091 ( .A1(n8237), .A2(n7532), .ZN(n5223) );
  OR2_X1 U5092 ( .A1(n8243), .A2(n8040), .ZN(n7752) );
  AND2_X1 U5093 ( .A1(n4305), .A2(n7742), .ZN(n7740) );
  NOR2_X1 U5094 ( .A1(n9417), .A2(n9331), .ZN(n4507) );
  NOR2_X1 U5095 ( .A1(n4510), .A2(n9340), .ZN(n4508) );
  AND2_X1 U5096 ( .A1(n8979), .A2(n8918), .ZN(n4537) );
  NOR2_X1 U5097 ( .A1(n9447), .A2(n9442), .ZN(n4512) );
  INV_X1 U5098 ( .A(SI_12_), .ZN(n9025) );
  NAND2_X1 U5099 ( .A1(n9199), .A2(n8684), .ZN(n9180) );
  INV_X1 U5100 ( .A(n8623), .ZN(n4437) );
  NAND2_X1 U5101 ( .A1(n8875), .A2(n4267), .ZN(n4693) );
  OR2_X1 U5102 ( .A1(n9270), .A2(n9286), .ZN(n8675) );
  OR2_X1 U5103 ( .A1(n9311), .A2(n9284), .ZN(n8667) );
  OAI21_X1 U5104 ( .B1(n7116), .B2(n4425), .A(n7203), .ZN(n4424) );
  NAND2_X1 U5105 ( .A1(n4365), .A2(n6452), .ZN(n8465) );
  INV_X1 U5106 ( .A(n6515), .ZN(n4365) );
  OR2_X1 U5107 ( .A1(n9427), .A2(n8905), .ZN(n8923) );
  INV_X1 U5108 ( .A(n8992), .ZN(n4536) );
  OR2_X1 U5109 ( .A1(n9447), .A2(n8895), .ZN(n8567) );
  NAND2_X1 U5110 ( .A1(n4693), .A2(n4692), .ZN(n4683) );
  NAND2_X1 U5111 ( .A1(n4279), .A2(n4685), .ZN(n4684) );
  NAND2_X1 U5112 ( .A1(n4686), .A2(n4692), .ZN(n4685) );
  INV_X1 U5113 ( .A(n4688), .ZN(n4686) );
  OR2_X1 U5114 ( .A1(n5641), .A2(n4736), .ZN(n5586) );
  NAND2_X1 U5115 ( .A1(n6218), .A2(n6217), .ZN(n6231) );
  OR2_X1 U5116 ( .A1(n6216), .A2(n6215), .ZN(n6217) );
  OR2_X1 U5117 ( .A1(n6214), .A2(n6213), .ZN(n6218) );
  AND2_X1 U5118 ( .A1(n5312), .A2(n5298), .ZN(n5310) );
  AOI21_X1 U5119 ( .B1(n4726), .B2(n4724), .A(n4723), .ZN(n4722) );
  INV_X1 U5120 ( .A(n4726), .ZN(n4725) );
  INV_X1 U5121 ( .A(n5242), .ZN(n4723) );
  OR2_X1 U5122 ( .A1(n5187), .A2(n5186), .ZN(n4714) );
  NAND2_X1 U5123 ( .A1(n4702), .A2(n4704), .ZN(n5161) );
  AOI21_X1 U5124 ( .B1(n5143), .B2(n4705), .A(n4321), .ZN(n4704) );
  OR2_X1 U5125 ( .A1(n5072), .A2(n4719), .ZN(n4271) );
  INV_X1 U5126 ( .A(n5049), .ZN(n4719) );
  INV_X1 U5127 ( .A(n4718), .ZN(n4717) );
  OAI21_X1 U5128 ( .B1(n4720), .B2(n4271), .A(n5071), .ZN(n4718) );
  NAND2_X1 U5129 ( .A1(n4482), .A2(n4486), .ZN(n5030) );
  OAI21_X1 U5130 ( .B1(n6281), .B2(n4361), .A(n4360), .ZN(n4985) );
  NAND2_X1 U5131 ( .A1(n6281), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n4360) );
  XNOR2_X1 U5132 ( .A(n4876), .B(SI_1_), .ZN(n4873) );
  NOR2_X1 U5133 ( .A1(n7442), .A2(n4566), .ZN(n4565) );
  INV_X1 U5134 ( .A(n4571), .ZN(n4566) );
  INV_X1 U5135 ( .A(n8174), .ZN(n6722) );
  XNOR2_X1 U5136 ( .A(n6650), .B(n6722), .ZN(n6648) );
  NOR2_X1 U5137 ( .A1(n7515), .A2(n4580), .ZN(n4579) );
  INV_X1 U5138 ( .A(n4581), .ZN(n4580) );
  OR2_X1 U5139 ( .A1(n7422), .A2(n8081), .ZN(n4581) );
  OAI22_X1 U5140 ( .A1(n7546), .A2(n7547), .B1(n7432), .B2(n8014), .ZN(n7433)
         );
  AOI21_X1 U5141 ( .B1(n7410), .B2(n7411), .A(n4312), .ZN(n4553) );
  OAI21_X1 U5142 ( .B1(n4548), .B2(n4546), .A(n4324), .ZN(n4545) );
  INV_X1 U5143 ( .A(n7449), .ZN(n4546) );
  INV_X1 U5144 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n4857) );
  AND4_X1 U5145 ( .A1(n5184), .A2(n5183), .A3(n5182), .A4(n5181), .ZN(n7576)
         );
  NAND2_X1 U5146 ( .A1(n5485), .A2(n5484), .ZN(n6631) );
  OR2_X1 U5147 ( .A1(n6837), .A2(n6838), .ZN(n4449) );
  NAND2_X1 U5148 ( .A1(n9753), .A2(n9752), .ZN(n4596) );
  OR2_X1 U5149 ( .A1(n9787), .A2(n9788), .ZN(n4590) );
  OR2_X1 U5150 ( .A1(n5090), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5091) );
  OR2_X1 U5151 ( .A1(n9819), .A2(n5098), .ZN(n4603) );
  NAND2_X1 U5152 ( .A1(n9830), .A2(n9831), .ZN(n9829) );
  NAND2_X1 U5153 ( .A1(n9844), .A2(n7883), .ZN(n9862) );
  NAND2_X1 U5154 ( .A1(n4586), .A2(n4297), .ZN(n4585) );
  AND2_X1 U5155 ( .A1(n4585), .A2(n4584), .ZN(n9866) );
  INV_X1 U5156 ( .A(n9867), .ZN(n4584) );
  NOR2_X1 U5157 ( .A1(n5146), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n5173) );
  NAND2_X1 U5158 ( .A1(n5329), .A2(n7776), .ZN(n7950) );
  NAND2_X1 U5159 ( .A1(n5302), .A2(n5301), .ZN(n5322) );
  INV_X1 U5160 ( .A(n5303), .ZN(n5302) );
  OR2_X1 U5161 ( .A1(n5265), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5285) );
  OR2_X1 U5162 ( .A1(n5235), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5247) );
  OR2_X1 U5163 ( .A1(n5192), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5217) );
  OR2_X1 U5164 ( .A1(n5152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5179) );
  NAND2_X1 U5165 ( .A1(n5079), .A2(n5078), .ZN(n5096) );
  INV_X1 U5166 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5078) );
  INV_X1 U5167 ( .A(n5080), .ZN(n5079) );
  AND4_X1 U5168 ( .A1(n5102), .A2(n5101), .A3(n5100), .A4(n5099), .ZN(n7415)
         );
  OR2_X1 U5169 ( .A1(n5039), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5065) );
  OR2_X1 U5170 ( .A1(n7211), .A2(n7711), .ZN(n4628) );
  INV_X1 U5171 ( .A(n7827), .ZN(n7339) );
  OR2_X1 U5172 ( .A1(n4952), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n4974) );
  INV_X1 U5173 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n4910) );
  NAND2_X1 U5174 ( .A1(n4771), .A2(n5416), .ZN(n7085) );
  NAND2_X1 U5175 ( .A1(n5389), .A2(n5388), .ZN(n7654) );
  AND2_X1 U5176 ( .A1(n5345), .A2(n5344), .ZN(n7938) );
  OR2_X1 U5177 ( .A1(n7782), .A2(n7625), .ZN(n7941) );
  AND2_X1 U5178 ( .A1(n7771), .A2(n7773), .ZN(n7973) );
  OAI21_X1 U5179 ( .B1(n7995), .B2(n5270), .A(n5271), .ZN(n7982) );
  NAND2_X1 U5180 ( .A1(n4638), .A2(n7759), .ZN(n7995) );
  NAND2_X1 U5181 ( .A1(n8007), .A2(n7755), .ZN(n4638) );
  NAND2_X1 U5182 ( .A1(n8049), .A2(n5441), .ZN(n8034) );
  NAND2_X1 U5183 ( .A1(n8057), .A2(n7744), .ZN(n5440) );
  AND2_X1 U5184 ( .A1(n4800), .A2(n5435), .ZN(n4799) );
  INV_X1 U5185 ( .A(n4616), .ZN(n4615) );
  OAI21_X1 U5186 ( .B1(n8091), .B2(n4617), .A(n7737), .ZN(n4616) );
  NAND2_X1 U5187 ( .A1(n5104), .A2(n4618), .ZN(n4617) );
  INV_X1 U5188 ( .A(n5103), .ZN(n4618) );
  INV_X1 U5189 ( .A(n7740), .ZN(n8078) );
  INV_X1 U5190 ( .A(n7358), .ZN(n4613) );
  NAND2_X1 U5191 ( .A1(n7314), .A2(n7627), .ZN(n5433) );
  INV_X1 U5192 ( .A(n8080), .ZN(n8161) );
  AND2_X1 U5193 ( .A1(n5018), .A2(n5017), .ZN(n9942) );
  AND2_X1 U5194 ( .A1(n5009), .A2(n5008), .ZN(n9937) );
  INV_X1 U5195 ( .A(n9966), .ZN(n9948) );
  INV_X1 U5196 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4846) );
  INV_X1 U5197 ( .A(n4845), .ZN(n4798) );
  NAND2_X1 U5198 ( .A1(n5458), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5461) );
  NAND2_X1 U5199 ( .A1(n5461), .A2(n5459), .ZN(n5463) );
  AND2_X1 U5200 ( .A1(n5405), .A2(n5399), .ZN(n6643) );
  INV_X1 U5201 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5211) );
  OR2_X1 U5202 ( .A1(n4291), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5016) );
  NAND2_X1 U5203 ( .A1(n7020), .A2(n5775), .ZN(n5792) );
  NAND2_X1 U5204 ( .A1(n6592), .A2(n4757), .ZN(n4756) );
  AND2_X1 U5205 ( .A1(n5753), .A2(n5732), .ZN(n4755) );
  OR2_X1 U5206 ( .A1(n7019), .A2(n5768), .ZN(n5753) );
  NAND2_X1 U5207 ( .A1(n5958), .A2(n4766), .ZN(n4765) );
  INV_X1 U5208 ( .A(n4751), .ZN(n4750) );
  OAI21_X1 U5209 ( .B1(n4294), .B2(n4752), .A(n8386), .ZN(n4751) );
  NAND2_X1 U5210 ( .A1(n4754), .A2(n4294), .ZN(n7225) );
  NAND2_X1 U5211 ( .A1(n4384), .A2(n4350), .ZN(n4754) );
  INV_X1 U5212 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5849) );
  INV_X1 U5213 ( .A(n8396), .ZN(n4762) );
  INV_X1 U5214 ( .A(n7206), .ZN(n8388) );
  OR2_X1 U5215 ( .A1(n5897), .A2(n5896), .ZN(n4769) );
  OR2_X1 U5216 ( .A1(n8650), .A2(n4263), .ZN(n8705) );
  NAND2_X1 U5217 ( .A1(n8644), .A2(n8646), .ZN(n4378) );
  AND2_X1 U5218 ( .A1(n8761), .A2(n4475), .ZN(n8772) );
  NAND2_X1 U5219 ( .A1(n8760), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n4475) );
  OR2_X1 U5220 ( .A1(n8772), .A2(n8771), .ZN(n4474) );
  NOR2_X1 U5221 ( .A1(n9582), .A2(n4472), .ZN(n9540) );
  AND2_X1 U5222 ( .A1(n9587), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n4472) );
  NOR2_X1 U5223 ( .A1(n9540), .A2(n9539), .ZN(n9538) );
  OR2_X1 U5224 ( .A1(n9526), .A2(n9525), .ZN(n4467) );
  AND2_X1 U5225 ( .A1(n4467), .A2(n4466), .ZN(n9597) );
  NAND2_X1 U5226 ( .A1(n9532), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n4466) );
  OR2_X1 U5227 ( .A1(n9597), .A2(n9598), .ZN(n4465) );
  OR2_X1 U5228 ( .A1(n9608), .A2(n9609), .ZN(n4471) );
  AND2_X1 U5229 ( .A1(n4471), .A2(n4470), .ZN(n9624) );
  NAND2_X1 U5230 ( .A1(n9615), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n4470) );
  OR2_X1 U5231 ( .A1(n9624), .A2(n9623), .ZN(n4469) );
  AND2_X1 U5232 ( .A1(n4469), .A2(n4468), .ZN(n8812) );
  NAND2_X1 U5233 ( .A1(n9627), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n4468) );
  NAND2_X1 U5234 ( .A1(n8992), .A2(n4537), .ZN(n8977) );
  INV_X1 U5235 ( .A(n8917), .ZN(n4538) );
  NAND2_X1 U5236 ( .A1(n9006), .A2(n4540), .ZN(n8992) );
  AND2_X1 U5237 ( .A1(n8993), .A2(n8917), .ZN(n4540) );
  OR2_X1 U5238 ( .A1(n5945), .A2(n8418), .ZN(n5966) );
  NAND2_X1 U5239 ( .A1(n4542), .A2(n4267), .ZN(n4690) );
  NAND2_X1 U5240 ( .A1(n4267), .A2(n9284), .ZN(n4692) );
  OR2_X1 U5241 ( .A1(n9296), .A2(n4693), .ZN(n4680) );
  INV_X1 U5242 ( .A(n5889), .ZN(n5887) );
  INV_X1 U5243 ( .A(n8723), .ZN(n9286) );
  NAND2_X1 U5244 ( .A1(n4438), .A2(n4542), .ZN(n9278) );
  INV_X1 U5245 ( .A(n9280), .ZN(n4438) );
  NOR2_X1 U5246 ( .A1(n8874), .A2(n8873), .ZN(n9296) );
  NOR2_X1 U5247 ( .A1(n9408), .A2(n8725), .ZN(n8873) );
  OR2_X1 U5248 ( .A1(n9296), .A2(n9299), .ZN(n4696) );
  NOR2_X1 U5249 ( .A1(n7110), .A2(n8726), .ZN(n4662) );
  AND2_X1 U5250 ( .A1(n6973), .A2(n7115), .ZN(n7111) );
  OR2_X1 U5251 ( .A1(n8662), .A2(n8584), .ZN(n7117) );
  NOR2_X1 U5252 ( .A1(n6896), .A2(n6942), .ZN(n6915) );
  OAI211_X1 U5253 ( .C1(n8575), .C2(n4643), .A(n4640), .B(n6512), .ZN(n6565)
         );
  NOR2_X1 U5254 ( .A1(n4643), .A2(n4642), .ZN(n4641) );
  INV_X1 U5255 ( .A(n6510), .ZN(n4643) );
  NAND2_X1 U5256 ( .A1(n6453), .A2(n8575), .ZN(n6511) );
  INV_X1 U5257 ( .A(n8919), .ZN(n8979) );
  AOI21_X1 U5258 ( .B1(n4671), .B2(n4669), .A(n4318), .ZN(n4668) );
  INV_X1 U5259 ( .A(n4676), .ZN(n4669) );
  INV_X1 U5260 ( .A(n4671), .ZN(n4670) );
  NAND2_X1 U5261 ( .A1(n4676), .A2(n8894), .ZN(n4675) );
  AND2_X1 U5262 ( .A1(n8567), .A2(n8917), .ZN(n9007) );
  NOR2_X1 U5263 ( .A1(n9175), .A2(n8891), .ZN(n8894) );
  NAND2_X1 U5264 ( .A1(n8890), .A2(n8889), .ZN(n9159) );
  NAND2_X1 U5265 ( .A1(n9189), .A2(n9165), .ZN(n8889) );
  XNOR2_X1 U5266 ( .A(n6231), .B(n6230), .ZN(n7607) );
  MUX2_X1 U5267 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5583), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n5584) );
  NAND2_X1 U5268 ( .A1(n5369), .A2(n5368), .ZN(n5381) );
  XNOR2_X1 U5269 ( .A(n5331), .B(n5330), .ZN(n7308) );
  INV_X1 U5270 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5565) );
  NAND2_X1 U5271 ( .A1(n4706), .A2(n5129), .ZN(n5144) );
  NAND2_X1 U5272 ( .A1(n5127), .A2(n5126), .ZN(n4706) );
  NAND2_X1 U5273 ( .A1(n4483), .A2(n4485), .ZN(n4480) );
  AND2_X1 U5274 ( .A1(n5739), .A2(n5776), .ZN(n6549) );
  XNOR2_X1 U5275 ( .A(n5012), .B(n5011), .ZN(n6310) );
  AND2_X1 U5276 ( .A1(n5291), .A2(n5290), .ZN(n7550) );
  AND4_X1 U5277 ( .A1(n4980), .A2(n4979), .A3(n4978), .A4(n4977), .ZN(n7282)
         );
  NAND2_X1 U5278 ( .A1(n5338), .A2(n5337), .ZN(n7952) );
  NAND2_X1 U5279 ( .A1(n4418), .A2(n4311), .ZN(n4503) );
  NAND2_X1 U5280 ( .A1(n7808), .A2(n7807), .ZN(n4420) );
  XNOR2_X1 U5281 ( .A(n5400), .B(P2_IR_REG_22__SCAN_IN), .ZN(n7814) );
  NAND2_X1 U5282 ( .A1(n5399), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5400) );
  INV_X1 U5283 ( .A(n7282), .ZN(n7828) );
  INV_X1 U5284 ( .A(n7105), .ZN(n7830) );
  NAND2_X1 U5285 ( .A1(n9709), .A2(n4447), .ZN(n6383) );
  OR2_X1 U5286 ( .A1(n6382), .A2(n4250), .ZN(n4447) );
  NAND2_X1 U5287 ( .A1(n6606), .A2(n6605), .ZN(n6834) );
  OAI21_X1 U5288 ( .B1(n6839), .B2(n6610), .A(n6841), .ZN(n6842) );
  NOR2_X1 U5289 ( .A1(n5062), .A2(n5061), .ZN(n9778) );
  AND2_X1 U5290 ( .A1(n5116), .A2(n5130), .ZN(n9825) );
  XNOR2_X1 U5291 ( .A(n7912), .B(n7891), .ZN(n4607) );
  OR2_X1 U5292 ( .A1(n7915), .A2(n9732), .ZN(n4605) );
  NAND2_X1 U5293 ( .A1(n9503), .A2(n4373), .ZN(n7862) );
  OR2_X1 U5294 ( .A1(n9514), .A2(n8140), .ZN(n4373) );
  NOR3_X1 U5295 ( .A1(n7914), .A2(n4285), .A3(n4351), .ZN(n4604) );
  AOI21_X1 U5296 ( .B1(n9514), .B2(n9509), .A(n9507), .ZN(n4442) );
  OAI211_X1 U5297 ( .C1(n7946), .C2(n4779), .A(n4775), .B(n4773), .ZN(n5455)
         );
  XNOR2_X1 U5298 ( .A(n7946), .B(n4745), .ZN(n7947) );
  NAND2_X1 U5299 ( .A1(n5176), .A2(n5175), .ZN(n8143) );
  AND2_X1 U5300 ( .A1(n5086), .A2(n7726), .ZN(n4636) );
  INV_X1 U5301 ( .A(n7654), .ZN(n6208) );
  NAND2_X1 U5302 ( .A1(n5472), .A2(n5471), .ZN(n6322) );
  OR2_X1 U5303 ( .A1(n6309), .A2(n5734), .ZN(n5719) );
  AND2_X1 U5304 ( .A1(n6262), .A2(n6261), .ZN(n6103) );
  AND2_X1 U5305 ( .A1(n6260), .A2(n6261), .ZN(n6263) );
  NAND2_X1 U5306 ( .A1(n6079), .A2(n6078), .ZN(n8995) );
  OR2_X1 U5307 ( .A1(n9015), .A2(n6111), .ZN(n6037) );
  OR2_X1 U5308 ( .A1(n9171), .A2(n6111), .ZN(n6020) );
  OAI21_X1 U5309 ( .B1(n8858), .B2(n9632), .A(n4462), .ZN(n4461) );
  AOI21_X1 U5310 ( .B1(n8859), .B2(n9595), .A(n4463), .ZN(n4462) );
  NOR2_X1 U5311 ( .A1(n6238), .A2(n9308), .ZN(n8862) );
  XNOR2_X1 U5312 ( .A(n8867), .B(n8563), .ZN(n6238) );
  NAND2_X1 U5313 ( .A1(n8926), .A2(n4342), .ZN(n4652) );
  NAND2_X1 U5314 ( .A1(n4653), .A2(n4651), .ZN(n4650) );
  NOR2_X1 U5315 ( .A1(n8926), .A2(n4342), .ZN(n4651) );
  NAND2_X1 U5316 ( .A1(n8907), .A2(n4647), .ZN(n4649) );
  AND2_X1 U5317 ( .A1(n8926), .A2(n4654), .ZN(n4647) );
  NAND2_X1 U5318 ( .A1(n4534), .A2(n4530), .ZN(n4531) );
  NAND2_X1 U5319 ( .A1(n8446), .A2(n4299), .ZN(n8468) );
  AND2_X1 U5320 ( .A1(n7701), .A2(n4417), .ZN(n4416) );
  NAND2_X1 U5321 ( .A1(n7685), .A2(n7801), .ZN(n4417) );
  INV_X1 U5322 ( .A(n7743), .ZN(n4386) );
  NOR2_X1 U5323 ( .A1(n4410), .A2(n4409), .ZN(n4408) );
  NAND2_X1 U5324 ( .A1(n7754), .A2(n7781), .ZN(n4409) );
  INV_X1 U5325 ( .A(n7757), .ZN(n4410) );
  NOR2_X1 U5326 ( .A1(n4273), .A2(n4408), .ZN(n4407) );
  AND2_X1 U5327 ( .A1(n4301), .A2(n4404), .ZN(n4403) );
  AOI21_X1 U5328 ( .B1(n4273), .B2(n4308), .A(n4405), .ZN(n4404) );
  NAND2_X1 U5329 ( .A1(n8443), .A2(n8442), .ZN(n8527) );
  NAND2_X1 U5330 ( .A1(n8605), .A2(n8923), .ZN(n4364) );
  NOR2_X1 U5331 ( .A1(n7649), .A2(n7648), .ZN(n4746) );
  AOI21_X1 U5332 ( .B1(n4495), .B2(n4494), .A(n4491), .ZN(n7793) );
  INV_X1 U5333 ( .A(n7780), .ZN(n4494) );
  NAND2_X1 U5334 ( .A1(n4493), .A2(n4492), .ZN(n4491) );
  NOR2_X1 U5335 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n4839) );
  INV_X1 U5336 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n4836) );
  AND2_X1 U5337 ( .A1(n8566), .A2(n8548), .ZN(n4381) );
  NOR2_X1 U5338 ( .A1(n9205), .A2(n4516), .ZN(n4515) );
  INV_X1 U5339 ( .A(n4517), .ZN(n4516) );
  NAND2_X1 U5340 ( .A1(n5385), .A2(n5384), .ZN(n6216) );
  INV_X1 U5341 ( .A(n5332), .ZN(n4713) );
  INV_X1 U5342 ( .A(n5226), .ZN(n4724) );
  NOR2_X1 U5343 ( .A1(n5142), .A2(n5125), .ZN(n4703) );
  INV_X1 U5344 ( .A(n5129), .ZN(n4705) );
  INV_X1 U5345 ( .A(n4699), .ZN(n4698) );
  OAI21_X1 U5346 ( .B1(n4983), .B2(n4700), .A(n4997), .ZN(n4699) );
  AND2_X1 U5347 ( .A1(n4986), .A2(n4965), .ZN(n4488) );
  NOR2_X1 U5348 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P1_RD_REG_SCAN_IN), .ZN(
        n4733) );
  INV_X1 U5349 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4729) );
  NAND2_X1 U5350 ( .A1(n7242), .A2(n7241), .ZN(n7243) );
  NOR2_X1 U5351 ( .A1(n4797), .A2(n4453), .ZN(n4452) );
  NAND2_X1 U5352 ( .A1(n4843), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n4453) );
  NAND2_X1 U5353 ( .A1(n5169), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n4456) );
  NAND2_X1 U5354 ( .A1(n4457), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4458) );
  AND2_X1 U5355 ( .A1(n9879), .A2(n4451), .ZN(n7887) );
  NAND2_X1 U5356 ( .A1(n7885), .A2(n9876), .ZN(n4451) );
  NAND2_X1 U5357 ( .A1(n5454), .A2(n4790), .ZN(n4781) );
  INV_X1 U5358 ( .A(n5428), .ZN(n4794) );
  AND2_X1 U5359 ( .A1(n4304), .A2(n4803), .ZN(n4802) );
  NOR2_X1 U5360 ( .A1(n7660), .A2(n4808), .ZN(n4807) );
  INV_X1 U5361 ( .A(n5432), .ZN(n4810) );
  NOR2_X1 U5362 ( .A1(n9965), .A2(n7823), .ZN(n4808) );
  NAND2_X1 U5363 ( .A1(n6133), .A2(n8315), .ZN(n5649) );
  INV_X1 U5364 ( .A(n5841), .ZN(n4752) );
  AND2_X1 U5365 ( .A1(n7160), .A2(n4749), .ZN(n4747) );
  NOR2_X1 U5366 ( .A1(n4752), .A2(n7227), .ZN(n4749) );
  NAND2_X1 U5367 ( .A1(n5693), .A2(n5692), .ZN(n5694) );
  INV_X1 U5368 ( .A(n9494), .ZN(n5539) );
  NOR2_X1 U5369 ( .A1(n9372), .A2(n9380), .ZN(n4517) );
  AND2_X1 U5370 ( .A1(n9408), .A2(n8872), .ZN(n8620) );
  NOR2_X1 U5371 ( .A1(n9311), .A2(n9408), .ZN(n4525) );
  NAND2_X1 U5372 ( .A1(n6915), .A2(n9685), .ZN(n6803) );
  INV_X1 U5373 ( .A(n6451), .ZN(n4642) );
  NAND2_X1 U5374 ( .A1(n8406), .A2(n6437), .ZN(n6455) );
  AOI21_X1 U5375 ( .B1(n4429), .B2(n4431), .A(n4428), .ZN(n4427) );
  INV_X1 U5376 ( .A(n4430), .ZN(n4429) );
  OR2_X1 U5377 ( .A1(n9452), .A2(n8891), .ZN(n9008) );
  NAND2_X1 U5378 ( .A1(n9170), .A2(n9014), .ZN(n9013) );
  NOR2_X1 U5379 ( .A1(n9452), .A2(n9187), .ZN(n9170) );
  NAND2_X1 U5380 ( .A1(n9232), .A2(n4514), .ZN(n9187) );
  AND2_X1 U5381 ( .A1(n4515), .A2(n9459), .ZN(n4514) );
  NAND2_X1 U5382 ( .A1(n9232), .A2(n4515), .ZN(n9203) );
  OR2_X1 U5383 ( .A1(n8561), .A2(n6342), .ZN(n6433) );
  NOR2_X1 U5384 ( .A1(n6762), .A2(n6353), .ZN(n6761) );
  XNOR2_X1 U5385 ( .A(n6216), .B(n6215), .ZN(n6214) );
  AND2_X1 U5386 ( .A1(n5368), .A2(n5353), .ZN(n5366) );
  AND2_X1 U5387 ( .A1(n5349), .A2(n5336), .ZN(n5347) );
  NAND2_X1 U5388 ( .A1(n5562), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5563) );
  AND2_X1 U5389 ( .A1(n5242), .A2(n5230), .ZN(n5240) );
  INV_X1 U5390 ( .A(n4486), .ZN(n4485) );
  NAND2_X1 U5391 ( .A1(n4487), .A2(n4479), .ZN(n4478) );
  AND2_X1 U5392 ( .A1(n4828), .A2(n4484), .ZN(n4479) );
  INV_X1 U5393 ( .A(n5010), .ZN(n4484) );
  OAI21_X1 U5394 ( .B1(n6281), .B2(P1_DATAO_REG_5__SCAN_IN), .A(n4356), .ZN(
        n4963) );
  NAND2_X1 U5395 ( .A1(n6281), .A2(n6306), .ZN(n4356) );
  OAI21_X1 U5396 ( .B1(n4879), .B2(P1_DATAO_REG_2__SCAN_IN), .A(n4363), .ZN(
        n4901) );
  NAND2_X1 U5397 ( .A1(n4879), .A2(n4880), .ZN(n4363) );
  OR2_X1 U5398 ( .A1(n4563), .A2(n4821), .ZN(n4558) );
  INV_X1 U5399 ( .A(n4564), .ZN(n4563) );
  OAI21_X1 U5400 ( .B1(n4565), .B2(n4570), .A(n7470), .ZN(n4564) );
  OR2_X1 U5401 ( .A1(n4570), .A2(n4560), .ZN(n4559) );
  NAND2_X1 U5402 ( .A1(n4568), .A2(n4561), .ZN(n4560) );
  INV_X1 U5403 ( .A(n7499), .ZN(n4561) );
  OR2_X1 U5404 ( .A1(n4908), .A2(n4909), .ZN(n4916) );
  NAND2_X1 U5405 ( .A1(n5020), .A2(n5019), .ZN(n5039) );
  INV_X1 U5406 ( .A(n5021), .ZN(n5020) );
  NAND2_X1 U5407 ( .A1(n4575), .A2(n4573), .ZN(n7566) );
  AND2_X1 U5408 ( .A1(n4574), .A2(n7567), .ZN(n4573) );
  NAND2_X1 U5409 ( .A1(n4576), .A2(n4578), .ZN(n4574) );
  OR2_X1 U5410 ( .A1(n4971), .A2(n4932), .ZN(n4939) );
  NAND2_X1 U5411 ( .A1(n7440), .A2(n7949), .ZN(n4571) );
  INV_X1 U5412 ( .A(n7575), .ZN(n7596) );
  NAND2_X1 U5413 ( .A1(n4621), .A2(n7810), .ZN(n4620) );
  NAND2_X1 U5414 ( .A1(n7796), .A2(n4623), .ZN(n4622) );
  INV_X1 U5415 ( .A(n7809), .ZN(n4504) );
  NOR2_X1 U5416 ( .A1(n7651), .A2(n4739), .ZN(n7653) );
  AND4_X1 U5417 ( .A1(n5141), .A2(n5140), .A3(n5139), .A4(n5138), .ZN(n7419)
         );
  NAND2_X1 U5418 ( .A1(n4445), .A2(n4444), .ZN(n6363) );
  NAND2_X1 U5419 ( .A1(n7843), .A2(n4443), .ZN(n9711) );
  OR2_X1 U5420 ( .A1(n6380), .A2(n7842), .ZN(n4443) );
  NAND3_X1 U5421 ( .A1(n6401), .A2(n6490), .A3(P2_REG2_REG_3__SCAN_IN), .ZN(
        n6492) );
  NAND2_X1 U5422 ( .A1(n6609), .A2(n6608), .ZN(n6840) );
  AND2_X1 U5423 ( .A1(n4449), .A2(n4448), .ZN(n9738) );
  NAND2_X1 U5424 ( .A1(n7247), .A2(n7248), .ZN(n4448) );
  NAND2_X1 U5425 ( .A1(n9750), .A2(n9749), .ZN(n9748) );
  NAND2_X1 U5426 ( .A1(n7252), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4595) );
  AOI22_X1 U5427 ( .A1(n4594), .A2(n7892), .B1(n7893), .B2(
        P2_REG2_REG_9__SCAN_IN), .ZN(n9772) );
  AND2_X1 U5428 ( .A1(n5057), .A2(n5056), .ZN(n5060) );
  NAND2_X1 U5429 ( .A1(n4588), .A2(n4587), .ZN(n9803) );
  NAND2_X1 U5430 ( .A1(n4592), .A2(n4591), .ZN(n4587) );
  OR2_X1 U5431 ( .A1(n9787), .A2(n4589), .ZN(n4588) );
  XNOR2_X1 U5432 ( .A(n7856), .B(n9810), .ZN(n9812) );
  NAND2_X1 U5433 ( .A1(n9812), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n9811) );
  NAND2_X1 U5434 ( .A1(n9829), .A2(n7882), .ZN(n9845) );
  NAND2_X1 U5435 ( .A1(n9845), .A2(n9846), .ZN(n9844) );
  XNOR2_X1 U5436 ( .A(n7858), .B(n9841), .ZN(n9843) );
  NAND2_X1 U5437 ( .A1(n9843), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n9842) );
  NAND2_X1 U5438 ( .A1(n9861), .A2(n7884), .ZN(n9880) );
  NAND2_X1 U5439 ( .A1(n9880), .A2(n9881), .ZN(n9879) );
  XNOR2_X1 U5440 ( .A(n7860), .B(n9876), .ZN(n9878) );
  NAND2_X1 U5441 ( .A1(n9878), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n9877) );
  OR2_X1 U5442 ( .A1(n6631), .A2(n7222), .ZN(n6358) );
  NOR2_X1 U5443 ( .A1(n7909), .A2(n9886), .ZN(n9518) );
  NAND2_X1 U5444 ( .A1(n9504), .A2(n9505), .ZN(n9503) );
  NOR2_X1 U5445 ( .A1(n4783), .A2(n4777), .ZN(n4776) );
  NAND2_X1 U5446 ( .A1(n7650), .A2(n4790), .ZN(n4783) );
  AND2_X1 U5447 ( .A1(n4774), .A2(n4780), .ZN(n4773) );
  OAI21_X1 U5448 ( .B1(n5454), .B2(n4782), .A(n4781), .ZN(n4780) );
  NAND2_X1 U5449 ( .A1(n4778), .A2(n4777), .ZN(n4774) );
  NOR2_X1 U5450 ( .A1(n4784), .A2(n4791), .ZN(n4782) );
  NAND2_X1 U5451 ( .A1(n4629), .A2(n4633), .ZN(n7930) );
  OAI21_X1 U5452 ( .B1(n4268), .B2(n7625), .A(n7786), .ZN(n4633) );
  NOR2_X1 U5453 ( .A1(n4634), .A2(n4631), .ZN(n4630) );
  NAND2_X1 U5454 ( .A1(n5321), .A2(n5320), .ZN(n5339) );
  INV_X1 U5455 ( .A(n5322), .ZN(n5321) );
  OR2_X1 U5456 ( .A1(n5285), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5303) );
  NAND2_X1 U5457 ( .A1(n5246), .A2(n5245), .ZN(n5265) );
  INV_X1 U5458 ( .A(n5247), .ZN(n5246) );
  NAND2_X1 U5459 ( .A1(n5216), .A2(n5215), .ZN(n5235) );
  INV_X1 U5460 ( .A(n5217), .ZN(n5216) );
  NAND2_X1 U5461 ( .A1(n5178), .A2(n5177), .ZN(n5192) );
  INV_X1 U5462 ( .A(n5179), .ZN(n5178) );
  OR2_X1 U5463 ( .A1(n5119), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5136) );
  NAND2_X1 U5464 ( .A1(n5095), .A2(n5094), .ZN(n5119) );
  INV_X1 U5465 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5094) );
  INV_X1 U5466 ( .A(n5096), .ZN(n5095) );
  OR2_X1 U5467 ( .A1(n5065), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5080) );
  NAND2_X1 U5468 ( .A1(n4795), .A2(n5428), .ZN(n7272) );
  NAND2_X1 U5469 ( .A1(n4627), .A2(n4625), .ZN(n7270) );
  AND2_X1 U5470 ( .A1(n5045), .A2(n4626), .ZN(n4625) );
  AND4_X1 U5471 ( .A1(n5044), .A2(n5043), .A3(n5042), .A4(n5041), .ZN(n7555)
         );
  OR2_X1 U5472 ( .A1(n4991), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5021) );
  NAND2_X1 U5473 ( .A1(n7150), .A2(n5424), .ZN(n7212) );
  NAND2_X1 U5474 ( .A1(n4973), .A2(n4972), .ZN(n4991) );
  INV_X1 U5475 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n4972) );
  INV_X1 U5476 ( .A(n4974), .ZN(n4973) );
  AND2_X1 U5477 ( .A1(n7713), .A2(n7708), .ZN(n7701) );
  INV_X1 U5478 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n4933) );
  INV_X1 U5479 ( .A(n8159), .ZN(n8156) );
  INV_X1 U5480 ( .A(n7661), .ZN(n4872) );
  AND2_X1 U5481 ( .A1(n5506), .A2(n5488), .ZN(n6206) );
  AND2_X1 U5482 ( .A1(n5490), .A2(n7781), .ZN(n6200) );
  AND2_X1 U5483 ( .A1(n7776), .A2(n7777), .ZN(n7968) );
  AND3_X1 U5484 ( .A1(n5269), .A2(n5268), .A3(n5267), .ZN(n7987) );
  INV_X1 U5485 ( .A(n5441), .ZN(n4815) );
  AND2_X1 U5486 ( .A1(n5442), .A2(n4814), .ZN(n4813) );
  NAND2_X1 U5487 ( .A1(n5440), .A2(n4816), .ZN(n8049) );
  AOI21_X1 U5488 ( .B1(n4807), .B2(n4804), .A(n7359), .ZN(n4803) );
  INV_X1 U5489 ( .A(n4293), .ZN(n4804) );
  INV_X1 U5490 ( .A(n4807), .ZN(n4805) );
  AND4_X1 U5491 ( .A1(n5124), .A2(n5123), .A3(n5122), .A4(n5121), .ZN(n8082)
         );
  AND4_X1 U5492 ( .A1(n5085), .A2(n5084), .A3(n5083), .A4(n5082), .ZN(n7413)
         );
  NAND2_X1 U5493 ( .A1(n4809), .A2(n4806), .ZN(n7361) );
  INV_X1 U5494 ( .A(n4808), .ZN(n4806) );
  NAND2_X1 U5495 ( .A1(n5433), .A2(n4293), .ZN(n4809) );
  AND2_X1 U5496 ( .A1(n7663), .A2(n7662), .ZN(n9966) );
  AND2_X1 U5497 ( .A1(n6631), .A2(n6350), .ZN(n6637) );
  XNOR2_X1 U5498 ( .A(n5487), .B(n5486), .ZN(n6630) );
  NAND2_X1 U5499 ( .A1(n4457), .A2(n4857), .ZN(n4796) );
  OR2_X1 U5500 ( .A1(n5210), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n5396) );
  OR2_X1 U5501 ( .A1(n4881), .A2(n5169), .ZN(n4882) );
  AND2_X1 U5502 ( .A1(n8367), .A2(n6046), .ZN(n8300) );
  NAND2_X1 U5503 ( .A1(n8413), .A2(n5953), .ZN(n5958) );
  OR2_X1 U5504 ( .A1(n8415), .A2(n8414), .ZN(n5953) );
  XNOR2_X1 U5505 ( .A(n4355), .B(n5611), .ZN(n5595) );
  NAND2_X1 U5506 ( .A1(n5587), .A2(n5588), .ZN(n4355) );
  NAND2_X1 U5507 ( .A1(n6434), .A2(n5590), .ZN(n5588) );
  INV_X1 U5508 ( .A(n5709), .ZN(n5693) );
  OR2_X1 U5509 ( .A1(n5914), .A2(n5913), .ZN(n5915) );
  AND2_X1 U5510 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5681) );
  NAND2_X1 U5511 ( .A1(n8311), .A2(n4767), .ZN(n6420) );
  AND2_X1 U5512 ( .A1(n5742), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5758) );
  NAND2_X1 U5513 ( .A1(n5965), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5980) );
  INV_X1 U5514 ( .A(n5966), .ZN(n5965) );
  OR2_X1 U5515 ( .A1(n5976), .A2(n5975), .ZN(n4822) );
  NAND2_X1 U5516 ( .A1(n6013), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6030) );
  INV_X1 U5517 ( .A(n6014), .ZN(n6013) );
  INV_X1 U5518 ( .A(n6024), .ZN(n4761) );
  CLKBUF_X1 U5519 ( .A(n7160), .Z(n4374) );
  INV_X1 U5520 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5701) );
  NOR2_X1 U5521 ( .A1(n5702), .A2(n5701), .ZN(n5720) );
  NAND2_X1 U5522 ( .A1(n5681), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5702) );
  CLKBUF_X1 U5523 ( .A(n6337), .Z(n8711) );
  INV_X1 U5524 ( .A(n5722), .ZN(n8554) );
  NAND2_X1 U5525 ( .A1(n8777), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n4473) );
  NOR2_X1 U5526 ( .A1(n9538), .A2(n4343), .ZN(n9553) );
  NOR2_X1 U5527 ( .A1(n9553), .A2(n9552), .ZN(n9551) );
  AND2_X1 U5528 ( .A1(n4465), .A2(n4464), .ZN(n7011) );
  NAND2_X1 U5529 ( .A1(n7008), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n4464) );
  NOR2_X1 U5530 ( .A1(n8696), .A2(n4506), .ZN(n4505) );
  INV_X1 U5531 ( .A(n4507), .ZN(n4506) );
  INV_X1 U5532 ( .A(n8938), .ZN(n8955) );
  OR2_X1 U5533 ( .A1(n9180), .A2(n4439), .ZN(n9162) );
  INV_X1 U5534 ( .A(n8686), .ZN(n4439) );
  NAND2_X1 U5535 ( .A1(n9162), .A2(n4527), .ZN(n9164) );
  AND2_X1 U5536 ( .A1(n9161), .A2(n9163), .ZN(n4527) );
  AOI22_X1 U5537 ( .A1(n9196), .A2(n8886), .B1(n8885), .B2(n9463), .ZN(n9178)
         );
  NAND2_X1 U5538 ( .A1(n8628), .A2(n8681), .ZN(n9199) );
  NAND2_X1 U5539 ( .A1(n9232), .A2(n6228), .ZN(n9233) );
  NAND2_X1 U5540 ( .A1(n5921), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5945) );
  NAND2_X1 U5541 ( .A1(n7198), .A2(n4521), .ZN(n9268) );
  NOR2_X1 U5542 ( .A1(n9270), .A2(n4523), .ZN(n4521) );
  NAND2_X1 U5543 ( .A1(n4432), .A2(n4433), .ZN(n9253) );
  AND2_X1 U5544 ( .A1(n4434), .A2(n8675), .ZN(n4433) );
  OR2_X1 U5545 ( .A1(n4542), .A2(n4435), .ZN(n4434) );
  INV_X1 U5546 ( .A(n5872), .ZN(n5870) );
  NAND2_X1 U5547 ( .A1(n7198), .A2(n4525), .ZN(n9307) );
  NAND2_X1 U5548 ( .A1(n8488), .A2(n8494), .ZN(n4421) );
  INV_X1 U5549 ( .A(n4424), .ZN(n4423) );
  NAND2_X1 U5550 ( .A1(n7205), .A2(n8589), .ZN(n9298) );
  AND2_X1 U5551 ( .A1(n7121), .A2(n7237), .ZN(n7198) );
  NAND2_X1 U5552 ( .A1(n7198), .A2(n8871), .ZN(n9310) );
  INV_X1 U5553 ( .A(n4657), .ZN(n4656) );
  AOI21_X1 U5554 ( .B1(n4658), .B2(n4662), .A(n4313), .ZN(n4657) );
  AND2_X1 U5555 ( .A1(n8668), .A2(n9297), .ZN(n8589) );
  OR2_X1 U5556 ( .A1(n6803), .A2(n6970), .ZN(n6980) );
  NOR2_X1 U5557 ( .A1(n6980), .A2(n7110), .ZN(n7121) );
  NAND2_X1 U5558 ( .A1(n5799), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5851) );
  INV_X1 U5559 ( .A(n5801), .ZN(n5799) );
  OR2_X1 U5560 ( .A1(n8463), .A2(n6738), .ZN(n6885) );
  NAND2_X1 U5561 ( .A1(n4520), .A2(n4519), .ZN(n6896) );
  INV_X1 U5562 ( .A(n9676), .ZN(n4519) );
  OAI21_X1 U5563 ( .B1(n8446), .B2(n6561), .A(n8658), .ZN(n6795) );
  INV_X1 U5564 ( .A(n8730), .ZN(n6939) );
  NAND2_X1 U5565 ( .A1(n6500), .A2(n6451), .ZN(n6453) );
  NAND2_X1 U5566 ( .A1(n6455), .A2(n8653), .ZN(n8570) );
  NAND2_X1 U5567 ( .A1(n6435), .A2(n6756), .ZN(n6759) );
  INV_X1 U5568 ( .A(n8571), .ZN(n6435) );
  NAND2_X1 U5569 ( .A1(n4666), .A2(n4664), .ZN(n8963) );
  AND2_X1 U5570 ( .A1(n4665), .A2(n4347), .ZN(n4664) );
  NOR2_X1 U5571 ( .A1(n4536), .A2(n4535), .ZN(n8978) );
  INV_X1 U5572 ( .A(n8918), .ZN(n4535) );
  AND2_X1 U5573 ( .A1(n8568), .A2(n8626), .ZN(n9239) );
  INV_X1 U5574 ( .A(n4682), .ZN(n4681) );
  OAI21_X1 U5575 ( .B1(n4688), .B2(n4683), .A(n4345), .ZN(n4682) );
  AND2_X1 U5576 ( .A1(n6345), .A2(n8707), .ZN(n9675) );
  OAI21_X1 U5577 ( .B1(n9487), .B2(P1_D_REG_0__SCAN_IN), .A(n9489), .ZN(n6678)
         );
  INV_X1 U5578 ( .A(n6414), .ZN(n9669) );
  XNOR2_X1 U5579 ( .A(n6234), .B(n6233), .ZN(n8268) );
  OAI21_X1 U5580 ( .B1(n6231), .B2(n6230), .A(n6229), .ZN(n6234) );
  XNOR2_X1 U5581 ( .A(n6214), .B(SI_29_), .ZN(n8275) );
  XNOR2_X1 U5582 ( .A(n5580), .B(n5579), .ZN(n6243) );
  INV_X1 U5583 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5579) );
  NAND2_X1 U5584 ( .A1(n5578), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5580) );
  XNOR2_X1 U5585 ( .A(n5348), .B(n5347), .ZN(n7311) );
  NAND2_X1 U5586 ( .A1(n4710), .A2(n5332), .ZN(n5348) );
  NAND2_X1 U5587 ( .A1(n5331), .A2(n5330), .ZN(n4710) );
  OAI21_X1 U5588 ( .B1(n5274), .B2(n5273), .A(n5272), .ZN(n5281) );
  AND2_X1 U5589 ( .A1(n5293), .A2(n5279), .ZN(n5280) );
  NAND2_X1 U5590 ( .A1(n4714), .A2(n5188), .ZN(n5200) );
  OAI21_X1 U5591 ( .B1(n5030), .B2(n4271), .A(n4717), .ZN(n5089) );
  OR2_X1 U5592 ( .A1(n5776), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5777) );
  OAI21_X1 U5593 ( .B1(n5012), .B2(n5011), .A(n5010), .ZN(n5028) );
  INV_X1 U5594 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5676) );
  AND2_X1 U5595 ( .A1(n7181), .A2(n7180), .ZN(n7187) );
  AND2_X1 U5596 ( .A1(n5379), .A2(n5378), .ZN(n7937) );
  NAND2_X1 U5597 ( .A1(n4562), .A2(n4569), .ZN(n7471) );
  NAND2_X1 U5598 ( .A1(n4572), .A2(n4565), .ZN(n4562) );
  OAI21_X1 U5599 ( .B1(n7412), .B2(n4549), .A(n4548), .ZN(n7448) );
  INV_X1 U5600 ( .A(n7826), .ZN(n7378) );
  AND4_X1 U5601 ( .A1(n5197), .A2(n5196), .A3(n5195), .A4(n5194), .ZN(n8040)
         );
  OAI21_X1 U5602 ( .B1(n4558), .B2(n7472), .A(n4555), .ZN(n4554) );
  NAND2_X1 U5603 ( .A1(n4558), .A2(n4556), .ZN(n4555) );
  NAND2_X1 U5604 ( .A1(n4559), .A2(n4567), .ZN(n4556) );
  NAND2_X1 U5605 ( .A1(n5372), .A2(n5371), .ZN(n7797) );
  AND3_X1 U5606 ( .A1(n5239), .A2(n5238), .A3(n5237), .ZN(n8041) );
  AND2_X1 U5607 ( .A1(n5309), .A2(n5308), .ZN(n7986) );
  NAND2_X1 U5608 ( .A1(n7507), .A2(n7506), .ZN(n7505) );
  AND2_X1 U5609 ( .A1(n7505), .A2(n4579), .ZN(n7569) );
  NAND2_X1 U5610 ( .A1(n7505), .A2(n4581), .ZN(n7514) );
  NAND2_X1 U5611 ( .A1(n6948), .A2(n6947), .ZN(n6954) );
  NAND2_X1 U5612 ( .A1(n7342), .A2(n7341), .ZN(n7345) );
  AND4_X1 U5613 ( .A1(n5222), .A2(n5221), .A3(n5220), .A4(n5219), .ZN(n7532)
         );
  NAND2_X1 U5614 ( .A1(n4552), .A2(n4553), .ZN(n7538) );
  NAND2_X1 U5615 ( .A1(n7412), .A2(n7410), .ZN(n4552) );
  OR2_X1 U5616 ( .A1(n6670), .A2(n7924), .ZN(n7575) );
  AND2_X1 U5617 ( .A1(n7103), .A2(n7101), .ZN(n4582) );
  AND2_X1 U5618 ( .A1(n7102), .A2(n7101), .ZN(n7104) );
  AND2_X1 U5619 ( .A1(n5365), .A2(n5364), .ZN(n7948) );
  AND2_X1 U5620 ( .A1(n6662), .A2(n6661), .ZN(n7589) );
  NAND2_X1 U5621 ( .A1(n4572), .A2(n4571), .ZN(n7581) );
  NAND2_X1 U5622 ( .A1(n6666), .A2(n9896), .ZN(n7587) );
  AND4_X1 U5623 ( .A1(n5157), .A2(n5156), .A3(n5155), .A4(n5154), .ZN(n8081)
         );
  OR2_X1 U5624 ( .A1(n6670), .A2(n6669), .ZN(n7598) );
  OAI21_X1 U5625 ( .B1(n7412), .B2(n4547), .A(n4544), .ZN(n4543) );
  NAND2_X1 U5626 ( .A1(n4550), .A2(n7449), .ZN(n4547) );
  INV_X1 U5627 ( .A(n4545), .ZN(n4544) );
  INV_X1 U5628 ( .A(n7589), .ZN(n7591) );
  INV_X1 U5629 ( .A(n7558), .ZN(n7600) );
  INV_X1 U5630 ( .A(n7937), .ZN(n7820) );
  INV_X1 U5631 ( .A(n7948), .ZN(n7821) );
  INV_X1 U5632 ( .A(n7986), .ZN(n7961) );
  INV_X1 U5633 ( .A(n7987), .ZN(n8014) );
  INV_X1 U5634 ( .A(n7430), .ZN(n8026) );
  INV_X1 U5635 ( .A(n8041), .ZN(n8015) );
  INV_X1 U5636 ( .A(n7532), .ZN(n8051) );
  INV_X1 U5637 ( .A(n8040), .ZN(n8059) );
  INV_X1 U5638 ( .A(n8081), .ZN(n8058) );
  INV_X1 U5639 ( .A(n8082), .ZN(n7822) );
  INV_X1 U5640 ( .A(n7415), .ZN(n8093) );
  INV_X1 U5641 ( .A(n7413), .ZN(n7823) );
  INV_X1 U5642 ( .A(n7144), .ZN(n7831) );
  NAND2_X1 U5643 ( .A1(n4262), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4887) );
  OR2_X1 U5644 ( .A1(n6631), .A2(n6275), .ZN(n7833) );
  NAND2_X1 U5645 ( .A1(n7845), .A2(n7844), .ZN(n7843) );
  NAND2_X1 U5646 ( .A1(n6363), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n7844) );
  NOR2_X1 U5647 ( .A1(n6474), .A2(n4446), .ZN(n6478) );
  AND2_X1 U5648 ( .A1(n6475), .A2(n6476), .ZN(n4446) );
  NAND2_X1 U5649 ( .A1(n6478), .A2(n6477), .ZN(n6602) );
  NAND2_X1 U5650 ( .A1(n6834), .A2(n4450), .ZN(n6837) );
  OR2_X1 U5651 ( .A1(n6835), .A2(n6836), .ZN(n4450) );
  INV_X1 U5652 ( .A(n4449), .ZN(n7246) );
  INV_X1 U5653 ( .A(n4596), .ZN(n9755) );
  XNOR2_X1 U5654 ( .A(n5007), .B(P2_IR_REG_8__SCAN_IN), .ZN(n9743) );
  XNOR2_X1 U5655 ( .A(n4594), .B(n7261), .ZN(n7893) );
  INV_X1 U5656 ( .A(n4590), .ZN(n9786) );
  NAND2_X1 U5657 ( .A1(n4597), .A2(n4599), .ZN(n9834) );
  INV_X1 U5658 ( .A(n4586), .ZN(n9849) );
  INV_X1 U5659 ( .A(n4585), .ZN(n9868) );
  INV_X1 U5660 ( .A(n9732), .ZN(n9884) );
  INV_X1 U5661 ( .A(n7890), .ZN(n4441) );
  NOR2_X1 U5662 ( .A1(n4632), .A2(n4268), .ZN(n7942) );
  NOR2_X1 U5663 ( .A1(n7950), .A2(n5346), .ZN(n4632) );
  NAND2_X1 U5664 ( .A1(n5356), .A2(n5355), .ZN(n7940) );
  NAND2_X1 U5665 ( .A1(n5284), .A2(n5283), .ZN(n7991) );
  NAND2_X1 U5666 ( .A1(n5433), .A2(n5432), .ZN(n7324) );
  NAND2_X1 U5667 ( .A1(n6332), .A2(n5387), .ZN(n4502) );
  NAND2_X1 U5668 ( .A1(n4628), .A2(n7692), .ZN(n7297) );
  INV_X1 U5669 ( .A(n9937), .ZN(n7294) );
  AND2_X1 U5670 ( .A1(n5422), .A2(n5421), .ZN(n7131) );
  AND2_X1 U5671 ( .A1(n9904), .A2(n7062), .ZN(n8065) );
  AND2_X1 U5672 ( .A1(n7804), .A2(n7913), .ZN(n9897) );
  NAND2_X1 U5673 ( .A1(n6637), .A2(n6201), .ZN(n9896) );
  INV_X1 U5674 ( .A(n9907), .ZN(n9904) );
  OR2_X1 U5675 ( .A1(n7609), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4865) );
  INV_X1 U5676 ( .A(n9896), .ZN(n8102) );
  NAND2_X1 U5677 ( .A1(n7611), .A2(n7610), .ZN(n8183) );
  INV_X1 U5678 ( .A(n7797), .ZN(n8190) );
  XNOR2_X1 U5679 ( .A(n7967), .B(n7968), .ZN(n8204) );
  NAND2_X1 U5680 ( .A1(n5319), .A2(n5318), .ZN(n8201) );
  NAND2_X1 U5681 ( .A1(n5300), .A2(n5299), .ZN(n8207) );
  NAND2_X1 U5682 ( .A1(n4812), .A2(n5446), .ZN(n7974) );
  NAND2_X1 U5683 ( .A1(n5264), .A2(n5263), .ZN(n8219) );
  NAND2_X1 U5684 ( .A1(n5244), .A2(n5243), .ZN(n8225) );
  NAND2_X1 U5685 ( .A1(n8063), .A2(n7749), .ZN(n8048) );
  NAND2_X1 U5686 ( .A1(n5151), .A2(n5150), .ZN(n8250) );
  NAND2_X1 U5687 ( .A1(n5133), .A2(n5132), .ZN(n8256) );
  NAND2_X1 U5688 ( .A1(n4611), .A2(n4615), .ZN(n8077) );
  NAND2_X1 U5689 ( .A1(n4613), .A2(n4612), .ZN(n4611) );
  NAND2_X1 U5690 ( .A1(n5118), .A2(n5117), .ZN(n8263) );
  NAND2_X1 U5691 ( .A1(n4614), .A2(n5104), .ZN(n8089) );
  NAND2_X1 U5692 ( .A1(n7358), .A2(n5103), .ZN(n4614) );
  NAND2_X1 U5693 ( .A1(n5093), .A2(n5092), .ZN(n7659) );
  INV_X1 U5694 ( .A(n8212), .ZN(n8262) );
  NAND2_X1 U5695 ( .A1(n5402), .A2(n4455), .ZN(n5467) );
  NOR2_X1 U5696 ( .A1(n4797), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n4455) );
  INV_X1 U5697 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n9053) );
  NAND2_X1 U5698 ( .A1(n5464), .A2(n5463), .ZN(n7401) );
  INV_X1 U5699 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7224) );
  INV_X1 U5700 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n9092) );
  INV_X1 U5701 ( .A(n7814), .ZN(n7663) );
  INV_X1 U5702 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7080) );
  INV_X1 U5703 ( .A(n6643), .ZN(n7662) );
  INV_X1 U5704 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7076) );
  XNOR2_X1 U5705 ( .A(n5398), .B(n5397), .ZN(n7804) );
  OAI21_X1 U5706 ( .B1(n5396), .B2(P2_IR_REG_19__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5398) );
  INV_X1 U5707 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6934) );
  INV_X1 U5708 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6676) );
  INV_X1 U5709 ( .A(n9794), .ZN(n7900) );
  INV_X1 U5710 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6333) );
  INV_X1 U5711 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9046) );
  INV_X1 U5712 ( .A(n9761), .ZN(n7895) );
  INV_X1 U5713 ( .A(n7261), .ZN(n7892) );
  NOR2_X1 U5714 ( .A1(n4918), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n4941) );
  AND2_X1 U5715 ( .A1(n6288), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6271) );
  INV_X1 U5716 ( .A(n4756), .ZN(n6695) );
  AND2_X1 U5718 ( .A1(n6178), .A2(n9573), .ZN(n6173) );
  AND2_X1 U5719 ( .A1(n6122), .A2(n6121), .ZN(n6177) );
  NAND2_X1 U5720 ( .A1(n6132), .A2(n6131), .ZN(n9331) );
  NAND2_X1 U5721 ( .A1(n8311), .A2(n5656), .ZN(n6422) );
  OR2_X1 U5722 ( .A1(n6187), .A2(n8707), .ZN(n8419) );
  INV_X1 U5723 ( .A(n4370), .ZN(n6441) );
  CLKBUF_X1 U5724 ( .A(n8374), .Z(n8375) );
  NAND2_X1 U5725 ( .A1(n7225), .A2(n5841), .ZN(n8385) );
  AOI21_X1 U5726 ( .B1(n4374), .B2(n4384), .A(n7159), .ZN(n7228) );
  NAND2_X1 U5727 ( .A1(n6193), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9577) );
  NAND2_X1 U5728 ( .A1(n8354), .A2(n8358), .ZN(n8413) );
  NAND2_X1 U5729 ( .A1(n6179), .A2(n9257), .ZN(n8422) );
  NAND2_X1 U5730 ( .A1(n5897), .A2(n5896), .ZN(n4768) );
  AND2_X1 U5731 ( .A1(n6271), .A2(n6191), .ZN(n9486) );
  NAND2_X1 U5732 ( .A1(n8703), .A2(n4263), .ZN(n8704) );
  OR2_X1 U5733 ( .A1(n8286), .A2(n6111), .ZN(n6116) );
  INV_X1 U5734 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4476) );
  NOR2_X1 U5735 ( .A1(n9490), .A2(n8754), .ZN(n4477) );
  INV_X1 U5736 ( .A(n4474), .ZN(n8770) );
  AND2_X1 U5737 ( .A1(n9578), .A2(n6535), .ZN(n9579) );
  AND2_X1 U5738 ( .A1(n5716), .A2(n5697), .ZN(n9587) );
  INV_X1 U5739 ( .A(n4467), .ZN(n9524) );
  INV_X1 U5740 ( .A(n4465), .ZN(n9596) );
  INV_X1 U5741 ( .A(n4471), .ZN(n9607) );
  INV_X1 U5742 ( .A(n4469), .ZN(n9622) );
  OR2_X1 U5743 ( .A1(n9647), .A2(n9646), .ZN(n9656) );
  NAND2_X1 U5744 ( .A1(n4534), .A2(n4532), .ZN(n9326) );
  NAND2_X1 U5745 ( .A1(n8977), .A2(n8920), .ZN(n8965) );
  NOR2_X1 U5746 ( .A1(n4539), .A2(n4538), .ZN(n8994) );
  AND2_X1 U5747 ( .A1(n6072), .A2(n6052), .ZN(n8998) );
  NAND2_X1 U5748 ( .A1(n4687), .A2(n4690), .ZN(n9262) );
  NAND2_X1 U5749 ( .A1(n4691), .A2(n4695), .ZN(n4687) );
  NAND2_X1 U5750 ( .A1(n4680), .A2(n4692), .ZN(n4691) );
  NAND2_X1 U5751 ( .A1(n9278), .A2(n8623), .ZN(n9264) );
  NAND2_X1 U5752 ( .A1(n4694), .A2(n4695), .ZN(n9277) );
  NAND2_X1 U5753 ( .A1(n4696), .A2(n8724), .ZN(n4694) );
  NOR2_X1 U5754 ( .A1(n7111), .A2(n4662), .ZN(n7113) );
  NAND2_X1 U5755 ( .A1(n4422), .A2(n8488), .ZN(n7204) );
  NAND2_X1 U5756 ( .A1(n7117), .A2(n7116), .ZN(n4422) );
  INV_X1 U5757 ( .A(n9257), .ZN(n9312) );
  NAND2_X1 U5758 ( .A1(n6511), .A2(n6510), .ZN(n6513) );
  INV_X1 U5759 ( .A(n8982), .ZN(n9317) );
  NAND2_X1 U5760 ( .A1(n6188), .A2(n9486), .ZN(n9257) );
  OR2_X1 U5761 ( .A1(n6683), .A2(n9016), .ZN(n8982) );
  XOR2_X1 U5762 ( .A(n8932), .B(n8933), .Z(n9424) );
  NAND2_X1 U5763 ( .A1(n6106), .A2(n6105), .ZN(n9427) );
  NAND2_X1 U5764 ( .A1(n4663), .A2(n4668), .ZN(n8976) );
  OR2_X1 U5765 ( .A1(n9159), .A2(n4670), .ZN(n4663) );
  NAND2_X1 U5766 ( .A1(n4672), .A2(n4673), .ZN(n8991) );
  NAND2_X1 U5767 ( .A1(n9159), .A2(n4676), .ZN(n4672) );
  NAND2_X2 U5768 ( .A1(n6028), .A2(n6027), .ZN(n9447) );
  NAND2_X1 U5769 ( .A1(n4678), .A2(n8893), .ZN(n9004) );
  OR2_X1 U5770 ( .A1(n9159), .A2(n8894), .ZN(n4678) );
  NAND2_X1 U5771 ( .A1(n6310), .A2(n5959), .ZN(n4541) );
  INV_X1 U5772 ( .A(n8450), .ZN(n8452) );
  INV_X1 U5773 ( .A(n8315), .ZN(n7043) );
  INV_X1 U5774 ( .A(n8406), .ZN(n6994) );
  AND2_X1 U5775 ( .A1(n4276), .A2(n4645), .ZN(n4644) );
  INV_X1 U5776 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4645) );
  XNOR2_X1 U5777 ( .A(n5381), .B(n5380), .ZN(n7354) );
  CLKBUF_X1 U5778 ( .A(n6243), .Z(n8748) );
  NOR2_X1 U5779 ( .A1(n5577), .A2(n5557), .ZN(n5558) );
  NOR2_X1 U5780 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n5557) );
  INV_X1 U5781 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7079) );
  INV_X1 U5782 ( .A(n8645), .ZN(n8651) );
  INV_X1 U5783 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7069) );
  INV_X1 U5784 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n9142) );
  INV_X1 U5785 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6585) );
  AND2_X1 U5786 ( .A1(n5867), .A2(n5881), .ZN(n9627) );
  INV_X1 U5787 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6324) );
  INV_X1 U5788 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6311) );
  XNOR2_X1 U5789 ( .A(n4998), .B(n4997), .ZN(n6309) );
  XNOR2_X1 U5790 ( .A(n4503), .B(n7888), .ZN(n7818) );
  XNOR2_X1 U5791 ( .A(n4442), .B(n4441), .ZN(n4440) );
  NAND2_X1 U5792 ( .A1(n4607), .A2(n9754), .ZN(n4606) );
  AND2_X1 U5793 ( .A1(n5498), .A2(n5497), .ZN(n5499) );
  INV_X1 U5794 ( .A(n6209), .ZN(n6210) );
  OAI22_X1 U5795 ( .A1(n6208), .A2(n8126), .B1(n9982), .B2(n6207), .ZN(n6209)
         );
  INV_X1 U5796 ( .A(n4369), .ZN(n4368) );
  OAI22_X1 U5797 ( .A1(n8198), .A2(n8126), .B1(n9982), .B2(n8120), .ZN(n4369)
         );
  INV_X1 U5798 ( .A(n5517), .ZN(n5518) );
  OAI21_X1 U5799 ( .B1(n6208), .B2(n8212), .A(n5516), .ZN(n5517) );
  INV_X1 U5800 ( .A(n4367), .ZN(n4366) );
  OAI22_X1 U5801 ( .A1(n8198), .A2(n8212), .B1(n9967), .B2(n8197), .ZN(n4367)
         );
  NOR2_X1 U5802 ( .A1(n6263), .A2(n6262), .ZN(n6270) );
  OAI21_X1 U5803 ( .B1(n8860), .B2(n9016), .A(n4459), .ZN(P1_U3262) );
  AOI21_X1 U5804 ( .B1(n4461), .B2(n9016), .A(n4460), .ZN(n4459) );
  OAI21_X1 U5805 ( .B1(n9661), .B2(n4528), .A(n8861), .ZN(n4460) );
  OAI21_X1 U5806 ( .B1(n4531), .B2(n9706), .A(n4286), .ZN(n9328) );
  NAND2_X1 U5807 ( .A1(n8563), .A2(n9453), .ZN(n6258) );
  OAI21_X1 U5808 ( .B1(n4531), .B2(n9699), .A(n4284), .ZN(n9419) );
  NAND2_X1 U5809 ( .A1(n9396), .A2(n8876), .ZN(n4267) );
  AND2_X1 U5810 ( .A1(n7952), .A2(n7938), .ZN(n4268) );
  INV_X1 U5811 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9490) );
  AND2_X1 U5812 ( .A1(n4615), .A2(n4305), .ZN(n4269) );
  NAND2_X1 U5813 ( .A1(n9170), .A2(n4509), .ZN(n4272) );
  OR2_X1 U5814 ( .A1(n7175), .A2(n8388), .ZN(n8494) );
  AND2_X1 U5815 ( .A1(n8032), .A2(n4500), .ZN(n4273) );
  OR2_X1 U5816 ( .A1(n5896), .A2(n8427), .ZN(n4275) );
  AND2_X1 U5817 ( .A1(n5533), .A2(n4770), .ZN(n4276) );
  AND2_X1 U5818 ( .A1(n4271), .A2(n5087), .ZN(n4277) );
  NAND2_X1 U5819 ( .A1(n9164), .A2(n4306), .ZN(n9006) );
  INV_X1 U5820 ( .A(n9006), .ZN(n4539) );
  INV_X1 U5821 ( .A(n9340), .ZN(n8973) );
  NAND2_X1 U5822 ( .A1(n6085), .A2(n6084), .ZN(n9340) );
  AND2_X1 U5823 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n4278) );
  OR2_X1 U5824 ( .A1(n4688), .A2(n9484), .ZN(n4279) );
  AND2_X1 U5825 ( .A1(n7829), .A2(n7136), .ZN(n4280) );
  INV_X1 U5826 ( .A(n9281), .ZN(n4542) );
  AND2_X1 U5827 ( .A1(n4605), .A2(n4604), .ZN(n4281) );
  AND2_X1 U5828 ( .A1(n4652), .A2(n4648), .ZN(n4282) );
  AND2_X1 U5829 ( .A1(n7186), .A2(n7180), .ZN(n4283) );
  INV_X1 U5830 ( .A(n9270), .ZN(n9477) );
  NAND2_X1 U5831 ( .A1(n5901), .A2(n5900), .ZN(n9270) );
  OR2_X1 U5832 ( .A1(n9479), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n4284) );
  AND2_X1 U5833 ( .A1(n9875), .A2(n7913), .ZN(n4285) );
  OR2_X1 U5834 ( .A1(n9708), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n4286) );
  AND2_X1 U5835 ( .A1(n4590), .A2(n4593), .ZN(n4287) );
  INV_X1 U5836 ( .A(n5634), .ZN(n6092) );
  INV_X1 U5837 ( .A(n8716), .ZN(n6171) );
  OR3_X1 U5838 ( .A1(n5399), .A2(n4797), .A3(P2_IR_REG_27__SCAN_IN), .ZN(n4289) );
  INV_X1 U5839 ( .A(n7824), .ZN(n4501) );
  NAND2_X1 U5840 ( .A1(n6237), .A2(n6236), .ZN(n8563) );
  AND2_X1 U5841 ( .A1(n5027), .A2(n7692), .ZN(n4290) );
  INV_X1 U5842 ( .A(n7951), .ZN(n4745) );
  AOI22_X1 U5843 ( .A1(n8268), .A2(n5387), .B1(n7606), .B2(
        P1_DATAO_REG_31__SCAN_IN), .ZN(n8180) );
  INV_X1 U5844 ( .A(n8180), .ZN(n4623) );
  NAND2_X1 U5845 ( .A1(n4818), .A2(n4274), .ZN(n4291) );
  AND2_X1 U5846 ( .A1(n9170), .A2(n4512), .ZN(n4292) );
  NOR2_X1 U5847 ( .A1(n5434), .A2(n4810), .ZN(n4293) );
  NAND2_X1 U5848 ( .A1(n5880), .A2(n5879), .ZN(n4354) );
  AND2_X1 U5849 ( .A1(n7226), .A2(n4753), .ZN(n4294) );
  XNOR2_X1 U5850 ( .A(n4847), .B(P2_IR_REG_29__SCAN_IN), .ZN(n4852) );
  AND2_X1 U5851 ( .A1(n8541), .A2(n8598), .ZN(n4295) );
  INV_X1 U5852 ( .A(n8091), .ZN(n4389) );
  AND4_X1 U5853 ( .A1(n4957), .A2(n4956), .A3(n4955), .A4(n4954), .ZN(n7188)
         );
  INV_X1 U5854 ( .A(n7188), .ZN(n7829) );
  XNOR2_X1 U5855 ( .A(n7797), .B(n7937), .ZN(n7929) );
  INV_X1 U5856 ( .A(n7929), .ZN(n4742) );
  INV_X1 U5857 ( .A(n8920), .ZN(n4431) );
  INV_X1 U5858 ( .A(n7791), .ZN(n4493) );
  INV_X1 U5859 ( .A(n4570), .ZN(n4569) );
  NOR2_X1 U5860 ( .A1(n7441), .A2(n7938), .ZN(n4570) );
  NOR2_X1 U5861 ( .A1(n5453), .A2(n4789), .ZN(n4296) );
  OR2_X1 U5862 ( .A1(n9841), .A2(n7905), .ZN(n4297) );
  OR2_X1 U5863 ( .A1(n7829), .A2(n7136), .ZN(n4298) );
  NAND4_X2 U5864 ( .A1(n4890), .A2(n4889), .A3(n4888), .A4(n4887), .ZN(n7832)
         );
  AND3_X1 U5865 ( .A1(n4823), .A2(n4865), .A3(n4866), .ZN(n8174) );
  INV_X1 U5866 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6165) );
  NAND2_X1 U5867 ( .A1(n7613), .A2(n7800), .ZN(n7650) );
  AND3_X1 U5868 ( .A1(n8658), .A2(n8445), .A3(n4252), .ZN(n4299) );
  NAND2_X1 U5869 ( .A1(n4760), .A2(n8299), .ZN(n8394) );
  OR2_X1 U5870 ( .A1(n9436), .A2(n8995), .ZN(n4300) );
  OR2_X1 U5871 ( .A1(n7750), .A2(n7801), .ZN(n4301) );
  AND2_X1 U5872 ( .A1(n4474), .A2(n4473), .ZN(n4302) );
  INV_X1 U5873 ( .A(n4818), .ZN(n4918) );
  NAND2_X1 U5874 ( .A1(n4818), .A2(n4819), .ZN(n4958) );
  NAND2_X1 U5875 ( .A1(n4881), .A2(n4833), .ZN(n4897) );
  NOR2_X1 U5876 ( .A1(n9947), .A2(n7825), .ZN(n4303) );
  INV_X1 U5877 ( .A(n8696), .ZN(n9416) );
  NAND2_X1 U5878 ( .A1(n6225), .A2(n6224), .ZN(n8696) );
  NAND2_X1 U5879 ( .A1(n8263), .A2(n7822), .ZN(n4304) );
  INV_X1 U5880 ( .A(n9205), .ZN(n9463) );
  NAND2_X1 U5881 ( .A1(n5979), .A2(n5978), .ZN(n9205) );
  NAND2_X1 U5882 ( .A1(n5944), .A2(n5943), .ZN(n9380) );
  INV_X1 U5883 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5570) );
  NAND2_X1 U5884 ( .A1(n8256), .A2(n7419), .ZN(n4305) );
  AND2_X1 U5885 ( .A1(n8675), .A2(n8673), .ZN(n9263) );
  INV_X1 U5886 ( .A(n9263), .ZN(n4689) );
  AND2_X1 U5887 ( .A1(n9007), .A2(n9008), .ZN(n4306) );
  INV_X1 U5888 ( .A(n7472), .ZN(n4567) );
  OR2_X1 U5889 ( .A1(n7425), .A2(n8059), .ZN(n4307) );
  NAND2_X1 U5890 ( .A1(n7754), .A2(n7749), .ZN(n4308) );
  INV_X1 U5891 ( .A(n4619), .ZN(n4612) );
  NAND2_X1 U5892 ( .A1(n4389), .A2(n5104), .ZN(n4619) );
  AND2_X1 U5893 ( .A1(n7740), .A2(n7739), .ZN(n4309) );
  NOR2_X1 U5894 ( .A1(n7940), .A2(n7948), .ZN(n7782) );
  AND2_X1 U5895 ( .A1(n4458), .A2(n4456), .ZN(n4310) );
  AND2_X1 U5896 ( .A1(n4620), .A2(n4504), .ZN(n4311) );
  INV_X1 U5897 ( .A(n7741), .ZN(n8069) );
  INV_X1 U5898 ( .A(n4791), .ZN(n4790) );
  NOR2_X1 U5899 ( .A1(n8190), .A2(n7937), .ZN(n4791) );
  NOR2_X1 U5900 ( .A1(n7414), .A2(n7413), .ZN(n4312) );
  INV_X1 U5901 ( .A(n4817), .ZN(n4816) );
  NAND2_X1 U5902 ( .A1(n8050), .A2(n5439), .ZN(n4817) );
  AND2_X1 U5903 ( .A1(n7237), .A2(n8388), .ZN(n4313) );
  AND3_X1 U5904 ( .A1(n4383), .A2(n8457), .A3(n4382), .ZN(n4314) );
  OR2_X1 U5905 ( .A1(n7763), .A2(n7987), .ZN(n4315) );
  INV_X1 U5906 ( .A(n4510), .ZN(n4509) );
  NAND2_X1 U5907 ( .A1(n4512), .A2(n4511), .ZN(n4510) );
  INV_X1 U5908 ( .A(n4674), .ZN(n4673) );
  NAND2_X1 U5909 ( .A1(n4317), .A2(n4675), .ZN(n4674) );
  OR2_X1 U5910 ( .A1(n4797), .A2(n4796), .ZN(n4316) );
  AND2_X1 U5911 ( .A1(n8207), .A2(n7986), .ZN(n7626) );
  OR2_X1 U5912 ( .A1(n9014), .A2(n8895), .ZN(n4317) );
  INV_X1 U5913 ( .A(n8488), .ZN(n4425) );
  NOR2_X1 U5914 ( .A1(n9442), .A2(n8898), .ZN(n4318) );
  OR2_X1 U5915 ( .A1(n5399), .A2(n4845), .ZN(n4319) );
  AND2_X1 U5916 ( .A1(n7761), .A2(n7760), .ZN(n4320) );
  AND2_X1 U5917 ( .A1(n5145), .A2(SI_15_), .ZN(n4321) );
  AND2_X1 U5918 ( .A1(n5088), .A2(SI_12_), .ZN(n4322) );
  AND4_X1 U5919 ( .A1(n4842), .A2(n5211), .A3(n4841), .A4(n5397), .ZN(n4323)
         );
  INV_X1 U5920 ( .A(n8875), .ZN(n9299) );
  INV_X1 U5921 ( .A(n4550), .ZN(n4549) );
  NOR2_X1 U5922 ( .A1(n4551), .A2(n7417), .ZN(n4550) );
  NAND2_X1 U5923 ( .A1(n7418), .A2(n8082), .ZN(n4324) );
  INV_X1 U5924 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6286) );
  AND2_X1 U5925 ( .A1(n5896), .A2(n8427), .ZN(n4325) );
  NOR2_X1 U5926 ( .A1(n7416), .A2(n8093), .ZN(n4326) );
  NAND2_X1 U5927 ( .A1(n7759), .A2(n7758), .ZN(n4327) );
  INV_X1 U5928 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4457) );
  INV_X1 U5929 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4843) );
  INV_X1 U5930 ( .A(n4779), .ZN(n4778) );
  NAND2_X1 U5931 ( .A1(n5454), .A2(n4784), .ZN(n4779) );
  NAND2_X1 U5932 ( .A1(n8645), .A2(n7070), .ZN(n6338) );
  INV_X1 U5933 ( .A(n8594), .ZN(n9161) );
  OR2_X1 U5934 ( .A1(n7797), .A2(n7820), .ZN(n4328) );
  AND2_X1 U5935 ( .A1(n8006), .A2(n7757), .ZN(n4329) );
  AND2_X1 U5936 ( .A1(n8606), .A2(n8633), .ZN(n8566) );
  AND2_X1 U5937 ( .A1(n7622), .A2(n7794), .ZN(n4330) );
  NOR2_X1 U5938 ( .A1(n8603), .A2(n8646), .ZN(n4331) );
  NAND2_X1 U5939 ( .A1(n4596), .A2(n4595), .ZN(n4594) );
  AND2_X1 U5940 ( .A1(n8930), .A2(n8931), .ZN(n4332) );
  AND2_X1 U5941 ( .A1(n5198), .A2(n7749), .ZN(n4333) );
  OR2_X1 U5942 ( .A1(n5769), .A2(n6937), .ZN(n4334) );
  AND2_X1 U5943 ( .A1(n4717), .A2(n5087), .ZN(n4335) );
  AND2_X1 U5944 ( .A1(n7343), .A2(n7341), .ZN(n4336) );
  AND2_X1 U5945 ( .A1(n4298), .A2(n5421), .ZN(n4337) );
  AND2_X1 U5946 ( .A1(n7709), .A2(n4416), .ZN(n4338) );
  AND2_X1 U5947 ( .A1(n4402), .A2(n4403), .ZN(n4339) );
  INV_X1 U5948 ( .A(n4436), .ZN(n4435) );
  NOR2_X1 U5949 ( .A1(n8624), .A2(n4437), .ZN(n4436) );
  INV_X1 U5950 ( .A(n5732), .ZN(n5733) );
  NAND2_X1 U5951 ( .A1(n5731), .A2(n5730), .ZN(n5732) );
  INV_X1 U5952 ( .A(n4821), .ZN(n4568) );
  OR2_X1 U5953 ( .A1(n8183), .A2(n7612), .ZN(n7799) );
  OR2_X1 U5954 ( .A1(n4559), .A2(n4567), .ZN(n4340) );
  AND2_X1 U5955 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4341) );
  INV_X1 U5956 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n4834) );
  NAND2_X1 U5957 ( .A1(n6070), .A2(n6069), .ZN(n9436) );
  INV_X1 U5958 ( .A(n9436), .ZN(n4511) );
  NAND2_X1 U5959 ( .A1(n4628), .A2(n4290), .ZN(n7268) );
  NOR2_X1 U5960 ( .A1(n8944), .A2(n8929), .ZN(n4342) );
  AND2_X1 U5961 ( .A1(n9543), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n4343) );
  NAND2_X1 U5962 ( .A1(n4637), .A2(n4636), .ZN(n7328) );
  INV_X1 U5963 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n4361) );
  OAI21_X1 U5964 ( .B1(n5433), .B2(n4805), .A(n4803), .ZN(n8090) );
  NAND2_X1 U5965 ( .A1(n5869), .A2(n5868), .ZN(n9311) );
  NAND2_X1 U5966 ( .A1(n5848), .A2(n5847), .ZN(n9408) );
  NOR2_X1 U5967 ( .A1(n9268), .A2(n9385), .ZN(n9232) );
  NAND2_X1 U5968 ( .A1(n4765), .A2(n4822), .ZN(n8373) );
  AND2_X1 U5969 ( .A1(n5440), .A2(n5439), .ZN(n4344) );
  INV_X1 U5970 ( .A(n7949), .ZN(n7975) );
  AND2_X1 U5971 ( .A1(n5328), .A2(n5327), .ZN(n7949) );
  NAND2_X1 U5972 ( .A1(n9232), .A2(n4517), .ZN(n4518) );
  NAND2_X1 U5973 ( .A1(n7198), .A2(n4522), .ZN(n4526) );
  OR2_X1 U5974 ( .A1(n9477), .A2(n9286), .ZN(n4345) );
  INV_X1 U5975 ( .A(n4523), .ZN(n4522) );
  NAND2_X1 U5976 ( .A1(n4524), .A2(n4525), .ZN(n4523) );
  NAND2_X1 U5977 ( .A1(n5995), .A2(n5994), .ZN(n9189) );
  INV_X1 U5978 ( .A(n9189), .ZN(n9459) );
  AND2_X1 U5979 ( .A1(n5201), .A2(n5188), .ZN(n4346) );
  OR2_X1 U5980 ( .A1(n4511), .A2(n8900), .ZN(n4347) );
  INV_X1 U5981 ( .A(n4533), .ZN(n4532) );
  OAI22_X1 U5982 ( .A1(n8929), .A2(n9285), .B1(n8928), .B2(n8927), .ZN(n4533)
         );
  AND2_X1 U5983 ( .A1(n4769), .A2(n4768), .ZN(n4348) );
  AND2_X1 U5984 ( .A1(n4603), .A2(n4602), .ZN(n4349) );
  INV_X1 U5985 ( .A(n9311), .ZN(n9484) );
  INV_X1 U5986 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n4736) );
  INV_X1 U5987 ( .A(n7801), .ZN(n7781) );
  INV_X1 U5988 ( .A(n9294), .ZN(n4648) );
  OR2_X1 U5989 ( .A1(n6254), .A2(n6678), .ZN(n9706) );
  NOR2_X1 U5990 ( .A1(n6695), .A2(n5733), .ZN(n6935) );
  NAND2_X1 U5991 ( .A1(n5886), .A2(n5885), .ZN(n9396) );
  INV_X1 U5992 ( .A(n9396), .ZN(n4524) );
  NAND2_X1 U5993 ( .A1(n7090), .A2(n5419), .ZN(n7142) );
  NAND2_X1 U5994 ( .A1(n4637), .A2(n7726), .ZN(n7329) );
  AND2_X1 U5995 ( .A1(n4374), .A2(n5816), .ZN(n4350) );
  INV_X1 U5996 ( .A(n4593), .ZN(n4592) );
  NAND2_X1 U5997 ( .A1(n7897), .A2(n7898), .ZN(n4593) );
  NAND2_X1 U5998 ( .A1(n7904), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4601) );
  INV_X1 U5999 ( .A(n9654), .ZN(n4463) );
  OR3_X1 U6000 ( .A1(n6187), .A2(n8640), .A3(n9675), .ZN(n8424) );
  INV_X1 U6001 ( .A(n8424), .ZN(n9573) );
  AND2_X1 U6002 ( .A1(n6336), .A2(n6335), .ZN(n9283) );
  INV_X1 U6003 ( .A(n4520), .ZN(n6895) );
  NOR2_X1 U6004 ( .A1(n6563), .A2(n8458), .ZN(n4520) );
  XNOR2_X1 U6005 ( .A(n5212), .B(n5211), .ZN(n7888) );
  AND2_X1 U6006 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3151), .ZN(n4351) );
  INV_X1 U6007 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n4911) );
  INV_X1 U6008 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4734) );
  XNOR2_X1 U6009 ( .A(n6362), .B(n7812), .ZN(n7924) );
  NAND2_X1 U6010 ( .A1(n7812), .A2(n6394), .ZN(n4444) );
  OR2_X1 U6011 ( .A1(n7812), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n4445) );
  AND2_X1 U6012 ( .A1(n4837), .A2(n4839), .ZN(n4393) );
  NAND2_X1 U6013 ( .A1(n7946), .A2(n4296), .ZN(n4785) );
  NAND2_X1 U6014 ( .A1(n7298), .A2(n7635), .ZN(n4795) );
  NAND2_X1 U6015 ( .A1(n7984), .A2(n5445), .ZN(n4812) );
  NAND2_X1 U6016 ( .A1(n5448), .A2(n5447), .ZN(n7960) );
  NAND2_X1 U6017 ( .A1(n8329), .A2(n6010), .ZN(n6025) );
  NAND2_X1 U6018 ( .A1(n8384), .A2(n5862), .ZN(n5880) );
  NOR2_X1 U6019 ( .A1(n5794), .A2(n5793), .ZN(n9563) );
  INV_X1 U6020 ( .A(n4352), .ZN(n8348) );
  OAI21_X2 U6021 ( .B1(n5897), .B2(n4325), .A(n4275), .ZN(n4352) );
  NAND2_X2 U6022 ( .A1(n8291), .A2(n4354), .ZN(n5897) );
  OR2_X2 U6023 ( .A1(n5880), .A2(n5879), .ZN(n4353) );
  NAND2_X1 U6024 ( .A1(n4258), .A2(n4825), .ZN(n5556) );
  NAND2_X1 U6025 ( .A1(n8348), .A2(n8349), .ZN(n8347) );
  AND2_X2 U6027 ( .A1(n4354), .A2(n4353), .ZN(n8292) );
  NAND2_X2 U6028 ( .A1(n8292), .A2(n8293), .ZN(n8291) );
  NAND3_X1 U6029 ( .A1(n4760), .A2(n8299), .A3(n4762), .ZN(n8298) );
  NAND2_X1 U6030 ( .A1(n4759), .A2(n4761), .ZN(n4760) );
  NAND2_X1 U6031 ( .A1(n4756), .A2(n4755), .ZN(n5771) );
  NAND2_X1 U6032 ( .A1(n4748), .A2(n4750), .ZN(n8384) );
  NAND2_X1 U6033 ( .A1(n8374), .A2(n5993), .ZN(n8330) );
  AND2_X1 U6034 ( .A1(n5540), .A2(n5541), .ZN(n5542) );
  NAND2_X1 U6035 ( .A1(n5960), .A2(n8716), .ZN(n6337) );
  INV_X1 U6036 ( .A(n5960), .ZN(n4358) );
  MUX2_X1 U6037 ( .A(n8497), .B(n8496), .S(n4252), .Z(n8501) );
  NAND2_X1 U6038 ( .A1(n8551), .A2(n8550), .ZN(n8560) );
  AOI21_X1 U6039 ( .B1(n8531), .B2(n8922), .A(n8535), .ZN(n8532) );
  NAND2_X1 U6040 ( .A1(n8508), .A2(n8509), .ZN(n8515) );
  AOI21_X1 U6041 ( .B1(n8491), .B2(n8490), .A(n8489), .ZN(n8495) );
  NAND2_X1 U6042 ( .A1(n8465), .A2(n8460), .ZN(n8446) );
  NAND2_X1 U6043 ( .A1(n5648), .A2(n8406), .ZN(n5623) );
  NAND2_X1 U6044 ( .A1(n4380), .A2(n4331), .ZN(n4379) );
  OAI211_X1 U6045 ( .C1(n8507), .C2(n8506), .A(n9263), .B(n8505), .ZN(n8508)
         );
  NAND2_X1 U6046 ( .A1(n4697), .A2(n4986), .ZN(n4998) );
  NAND2_X1 U6047 ( .A1(n4490), .A2(n4965), .ZN(n4984) );
  XNOR2_X1 U6048 ( .A(n4259), .B(n5651), .ZN(n5653) );
  NAND2_X1 U6049 ( .A1(n4357), .A2(n5613), .ZN(n6413) );
  NAND2_X1 U6050 ( .A1(n6351), .A2(n6352), .ZN(n4357) );
  NAND2_X2 U6051 ( .A1(n4358), .A2(n8712), .ZN(n6701) );
  NAND2_X2 U6052 ( .A1(n5572), .A2(n5573), .ZN(n5960) );
  NAND2_X2 U6054 ( .A1(n6025), .A2(n6024), .ZN(n8299) );
  INV_X1 U6055 ( .A(n4986), .ZN(n4700) );
  NAND2_X1 U6056 ( .A1(n4490), .A2(n4488), .ZN(n4489) );
  INV_X1 U6057 ( .A(n5794), .ZN(n7160) );
  MUX2_X1 U6058 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9502), .S(n5602), .Z(n6782) );
  NAND2_X1 U6059 ( .A1(n4362), .A2(n4371), .ZN(n6411) );
  INV_X1 U6060 ( .A(n6413), .ZN(n4362) );
  NAND2_X1 U6061 ( .A1(n4984), .A2(n4983), .ZN(n4697) );
  NAND2_X1 U6062 ( .A1(n4379), .A2(n4378), .ZN(n8706) );
  NAND2_X1 U6063 ( .A1(n8604), .A2(n8645), .ZN(n4380) );
  OAI21_X1 U6064 ( .B1(n8521), .B2(n8522), .A(n9163), .ZN(n4377) );
  NAND2_X1 U6065 ( .A1(n4377), .A2(n4252), .ZN(n4376) );
  OAI21_X1 U6066 ( .B1(n8527), .B2(n8526), .A(n8525), .ZN(n8529) );
  AND2_X1 U6067 ( .A1(n6590), .A2(n5710), .ZN(n5711) );
  NAND3_X1 U6068 ( .A1(n4737), .A2(n4738), .A3(P1_DATAO_REG_1__SCAN_IN), .ZN(
        n4728) );
  NAND2_X1 U6069 ( .A1(n4878), .A2(n4877), .ZN(n4900) );
  NAND2_X1 U6070 ( .A1(n6760), .A2(n6440), .ZN(n6457) );
  NAND2_X1 U6071 ( .A1(n6761), .A2(n8571), .ZN(n6760) );
  INV_X1 U6072 ( .A(n8515), .ZN(n8513) );
  NAND2_X1 U6073 ( .A1(n8523), .A2(n8561), .ZN(n4375) );
  NAND2_X1 U6074 ( .A1(n4801), .A2(n4799), .ZN(n8079) );
  AOI21_X1 U6075 ( .B1(n5422), .B2(n4337), .A(n4280), .ZN(n7151) );
  OAI21_X1 U6076 ( .B1(n8196), .B2(n9969), .A(n4366), .ZN(P2_U3453) );
  OAI21_X1 U6077 ( .B1(n8196), .B2(n6211), .A(n4368), .ZN(P2_U3485) );
  NAND2_X1 U6078 ( .A1(n5559), .A2(n5558), .ZN(n7240) );
  INV_X1 U6079 ( .A(n6410), .ZN(n4371) );
  NAND2_X1 U6080 ( .A1(n5596), .A2(n5614), .ZN(n6410) );
  AOI21_X1 U6081 ( .B1(n4370), .B2(n6145), .A(n5591), .ZN(n5594) );
  OAI211_X1 U6082 ( .C1(n4440), .C2(n9508), .A(n4606), .B(n4281), .ZN(P2_U3201) );
  NAND3_X1 U6083 ( .A1(n5542), .A2(n5544), .A3(n5543), .ZN(n6434) );
  NAND2_X1 U6084 ( .A1(n8549), .A2(n4381), .ZN(n8551) );
  OAI21_X1 U6085 ( .B1(n8706), .B2(n8705), .A(n8704), .ZN(n8709) );
  OR2_X1 U6086 ( .A1(n8459), .A2(n8458), .ZN(n4382) );
  NAND2_X1 U6087 ( .A1(n8449), .A2(n8458), .ZN(n4383) );
  NAND2_X1 U6088 ( .A1(n6420), .A2(n5675), .ZN(n6572) );
  NAND2_X1 U6089 ( .A1(n8298), .A2(n8299), .ZN(n6047) );
  INV_X1 U6090 ( .A(n6423), .ZN(n5670) );
  NAND2_X2 U6091 ( .A1(n5401), .A2(n4843), .ZN(n5399) );
  AND4_X2 U6092 ( .A1(n4826), .A2(n4818), .A3(n4323), .A4(n4274), .ZN(n5401)
         );
  AND3_X2 U6093 ( .A1(n4834), .A2(n4881), .A3(n4833), .ZN(n4818) );
  OR2_X1 U6094 ( .A1(n7766), .A2(n7765), .ZN(n4398) );
  OR2_X1 U6095 ( .A1(n7753), .A2(n4407), .ZN(n4402) );
  NAND2_X1 U6096 ( .A1(n7753), .A2(n4401), .ZN(n4400) );
  AOI21_X1 U6097 ( .B1(n4401), .B2(n4407), .A(n4327), .ZN(n4399) );
  NAND3_X1 U6098 ( .A1(n7700), .A2(n4338), .A3(n4415), .ZN(n4414) );
  NAND3_X1 U6099 ( .A1(n7687), .A2(n7781), .A3(n7686), .ZN(n4415) );
  NAND4_X1 U6100 ( .A1(n4420), .A2(n7804), .A3(n7803), .A4(n4419), .ZN(n4418)
         );
  OAI22_X1 U6101 ( .A1(n7117), .A2(n4421), .B1(n7202), .B2(n4423), .ZN(n7205)
         );
  NAND2_X1 U6102 ( .A1(n8992), .A2(n4429), .ZN(n4426) );
  NAND2_X1 U6103 ( .A1(n4426), .A2(n4427), .ZN(n8949) );
  NAND2_X1 U6104 ( .A1(n9280), .A2(n4436), .ZN(n4432) );
  XNOR2_X2 U6105 ( .A(n6774), .B(n4370), .ZN(n8571) );
  NOR2_X4 U6106 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4881) );
  MUX2_X1 U6107 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n6542), .S(n8739), .Z(n8744)
         );
  NAND2_X1 U6108 ( .A1(n5012), .A2(n4483), .ZN(n4481) );
  NAND2_X1 U6109 ( .A1(n5012), .A2(n5010), .ZN(n4482) );
  NAND3_X1 U6110 ( .A1(n4481), .A2(n4480), .A3(n5049), .ZN(n5073) );
  NAND2_X1 U6111 ( .A1(n4698), .A2(n4489), .ZN(n4701) );
  NAND2_X1 U6112 ( .A1(n4962), .A2(n4961), .ZN(n4490) );
  NAND3_X1 U6113 ( .A1(n4498), .A2(n4496), .A3(n7968), .ZN(n4495) );
  NAND3_X1 U6114 ( .A1(n4737), .A2(n4738), .A3(n4341), .ZN(n4863) );
  INV_X2 U6115 ( .A(n4879), .ZN(n6276) );
  NAND3_X1 U6116 ( .A1(n4734), .A2(n4528), .A3(n4729), .ZN(n4738) );
  AND2_X1 U6117 ( .A1(n8938), .A2(n4507), .ZN(n8910) );
  NAND2_X1 U6118 ( .A1(n8938), .A2(n8944), .ZN(n8939) );
  NAND2_X1 U6119 ( .A1(n8938), .A2(n4505), .ZN(n8867) );
  NAND2_X1 U6120 ( .A1(n9170), .A2(n4508), .ZN(n8954) );
  AND2_X1 U6121 ( .A1(n4825), .A2(n5533), .ZN(n4513) );
  NAND2_X1 U6122 ( .A1(n4258), .A2(n4513), .ZN(n5582) );
  INV_X1 U6123 ( .A(n4518), .ZN(n9215) );
  INV_X1 U6124 ( .A(n4526), .ZN(n9288) );
  NOR2_X1 U6125 ( .A1(n9325), .A2(n4533), .ZN(n4530) );
  XNOR2_X1 U6126 ( .A(n8925), .B(n8566), .ZN(n4529) );
  INV_X8 U6127 ( .A(n6276), .ZN(n6281) );
  MUX2_X1 U6128 ( .A(n6304), .B(n6279), .S(n6276), .Z(n4946) );
  NAND3_X1 U6129 ( .A1(n4826), .A2(n4274), .A3(n4818), .ZN(n5146) );
  OAI211_X1 U6130 ( .C1(n7498), .C2(n4340), .A(n4557), .B(n4554), .ZN(n7478)
         );
  NAND3_X1 U6131 ( .A1(n7498), .A2(n4558), .A3(n4567), .ZN(n4557) );
  OR2_X1 U6132 ( .A1(n7498), .A2(n7499), .ZN(n4572) );
  NAND2_X1 U6133 ( .A1(n7342), .A2(n4336), .ZN(n7371) );
  NAND2_X1 U6134 ( .A1(n7507), .A2(n4576), .ZN(n4575) );
  NAND3_X1 U6135 ( .A1(n6948), .A2(n6952), .A3(n6947), .ZN(n7032) );
  OAI21_X2 U6136 ( .B1(n6642), .B2(n7652), .A(n6646), .ZN(n6650) );
  NAND2_X1 U6137 ( .A1(n7181), .A2(n4283), .ZN(n7286) );
  XNOR2_X1 U6138 ( .A(n7896), .B(n9778), .ZN(n9787) );
  INV_X1 U6139 ( .A(n4603), .ZN(n9818) );
  INV_X1 U6140 ( .A(n7902), .ZN(n4602) );
  NAND2_X1 U6141 ( .A1(n6401), .A2(n6490), .ZN(n6403) );
  NAND2_X1 U6142 ( .A1(n7358), .A2(n4269), .ZN(n4608) );
  NAND2_X1 U6143 ( .A1(n4608), .A2(n4609), .ZN(n8068) );
  NAND2_X1 U6144 ( .A1(n4624), .A2(n4622), .ZN(n4621) );
  OAI21_X1 U6145 ( .B1(n7624), .B2(n7623), .A(n4330), .ZN(n4624) );
  NAND2_X1 U6146 ( .A1(n7211), .A2(n4290), .ZN(n4627) );
  NAND2_X1 U6147 ( .A1(n5329), .A2(n4630), .ZN(n4629) );
  NAND2_X1 U6148 ( .A1(n8063), .A2(n4333), .ZN(n5199) );
  NAND2_X1 U6149 ( .A1(n8064), .A2(n5185), .ZN(n8063) );
  AND2_X1 U6150 ( .A1(n7812), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7322) );
  MUX2_X1 U6151 ( .A(P2_REG1_REG_1__SCAN_IN), .B(P2_REG2_REG_1__SCAN_IN), .S(
        n7812), .Z(n6379) );
  MUX2_X1 U6152 ( .A(P2_REG1_REG_2__SCAN_IN), .B(P2_REG2_REG_2__SCAN_IN), .S(
        n7812), .Z(n6381) );
  MUX2_X1 U6153 ( .A(P2_REG1_REG_3__SCAN_IN), .B(P2_REG2_REG_3__SCAN_IN), .S(
        n7812), .Z(n6473) );
  MUX2_X1 U6154 ( .A(P2_REG1_REG_4__SCAN_IN), .B(P2_REG2_REG_4__SCAN_IN), .S(
        n7812), .Z(n6601) );
  MUX2_X1 U6155 ( .A(P2_REG1_REG_5__SCAN_IN), .B(P2_REG2_REG_5__SCAN_IN), .S(
        n7812), .Z(n6833) );
  MUX2_X1 U6156 ( .A(P2_REG1_REG_6__SCAN_IN), .B(P2_REG2_REG_6__SCAN_IN), .S(
        n7812), .Z(n7245) );
  MUX2_X1 U6157 ( .A(P2_REG1_REG_7__SCAN_IN), .B(P2_REG2_REG_7__SCAN_IN), .S(
        n7812), .Z(n7249) );
  MUX2_X1 U6158 ( .A(P2_REG1_REG_8__SCAN_IN), .B(P2_REG2_REG_8__SCAN_IN), .S(
        n7812), .Z(n7250) );
  MUX2_X1 U6159 ( .A(P2_REG1_REG_9__SCAN_IN), .B(P2_REG2_REG_9__SCAN_IN), .S(
        n7812), .Z(n7875) );
  MUX2_X1 U6160 ( .A(P2_REG1_REG_10__SCAN_IN), .B(P2_REG2_REG_10__SCAN_IN), 
        .S(n7812), .Z(n7873) );
  MUX2_X1 U6161 ( .A(P2_REG1_REG_11__SCAN_IN), .B(P2_REG2_REG_11__SCAN_IN), 
        .S(n7812), .Z(n7872) );
  MUX2_X1 U6162 ( .A(P2_REG1_REG_12__SCAN_IN), .B(P2_REG2_REG_12__SCAN_IN), 
        .S(n7812), .Z(n7871) );
  MUX2_X1 U6163 ( .A(P2_REG1_REG_13__SCAN_IN), .B(P2_REG2_REG_13__SCAN_IN), 
        .S(n7812), .Z(n7870) );
  MUX2_X1 U6164 ( .A(P2_REG1_REG_14__SCAN_IN), .B(P2_REG2_REG_14__SCAN_IN), 
        .S(n7812), .Z(n7868) );
  MUX2_X1 U6165 ( .A(P2_REG1_REG_15__SCAN_IN), .B(P2_REG2_REG_15__SCAN_IN), 
        .S(n7812), .Z(n7867) );
  MUX2_X1 U6166 ( .A(P2_REG1_REG_16__SCAN_IN), .B(P2_REG2_REG_16__SCAN_IN), 
        .S(n7812), .Z(n7865) );
  MUX2_X1 U6167 ( .A(n7863), .B(n9887), .S(n7812), .Z(n7885) );
  MUX2_X1 U6168 ( .A(P2_REG1_REG_18__SCAN_IN), .B(P2_REG2_REG_18__SCAN_IN), 
        .S(n7812), .Z(n7886) );
  MUX2_X1 U6169 ( .A(n7889), .B(n7891), .S(n7812), .Z(n7890) );
  NAND2_X1 U6170 ( .A1(n6393), .A2(n4639), .ZN(n9732) );
  NAND2_X1 U6171 ( .A1(n6500), .A2(n4641), .ZN(n4640) );
  NAND2_X1 U6172 ( .A1(n4644), .A2(n5577), .ZN(n5536) );
  NAND2_X1 U6173 ( .A1(n5577), .A2(n4276), .ZN(n5581) );
  NAND2_X1 U6174 ( .A1(n8907), .A2(n4654), .ZN(n4653) );
  NAND2_X1 U6175 ( .A1(n4646), .A2(n4332), .ZN(P1_U3356) );
  NAND3_X1 U6176 ( .A1(n4650), .A2(n4282), .A3(n4649), .ZN(n4646) );
  NAND2_X1 U6177 ( .A1(n8907), .A2(n8906), .ZN(n8932) );
  NAND3_X1 U6178 ( .A1(n4650), .A2(n4649), .A3(n4652), .ZN(n9420) );
  AOI21_X1 U6179 ( .B1(n6973), .B2(n4658), .A(n4656), .ZN(n7197) );
  OAI21_X1 U6180 ( .B1(n6973), .B2(n4662), .A(n4658), .ZN(n4661) );
  INV_X1 U6181 ( .A(n4661), .ZN(n7196) );
  NAND2_X1 U6182 ( .A1(n9159), .A2(n4667), .ZN(n4666) );
  NAND3_X1 U6183 ( .A1(n4668), .A2(n4670), .A3(n4300), .ZN(n4665) );
  NAND2_X1 U6184 ( .A1(n9296), .A2(n4684), .ZN(n4679) );
  NAND2_X1 U6185 ( .A1(n4679), .A2(n4681), .ZN(n9247) );
  NAND2_X1 U6186 ( .A1(n9296), .A2(n9311), .ZN(n4695) );
  INV_X1 U6187 ( .A(n4696), .ZN(n9295) );
  NAND2_X1 U6188 ( .A1(n5127), .A2(n4703), .ZN(n4702) );
  NAND2_X1 U6189 ( .A1(n4714), .A2(n4346), .ZN(n5205) );
  NAND2_X1 U6190 ( .A1(n5030), .A2(n4335), .ZN(n4715) );
  NAND2_X1 U6191 ( .A1(n4715), .A2(n4716), .ZN(n5107) );
  NAND2_X1 U6192 ( .A1(n5030), .A2(n5029), .ZN(n5051) );
  OAI21_X1 U6193 ( .B1(n5225), .B2(n5224), .A(n5226), .ZN(n5241) );
  NAND3_X1 U6194 ( .A1(n4728), .A2(n4731), .A3(n4730), .ZN(n4876) );
  NAND3_X1 U6195 ( .A1(n4732), .A2(n4735), .A3(P2_DATAO_REG_1__SCAN_IN), .ZN(
        n4730) );
  NAND3_X1 U6196 ( .A1(n4733), .A2(n4734), .A3(P2_DATAO_REG_1__SCAN_IN), .ZN(
        n4731) );
  NAND3_X1 U6197 ( .A1(n7799), .A2(n4740), .A3(n7795), .ZN(n4739) );
  NAND2_X1 U6198 ( .A1(n9562), .A2(n4747), .ZN(n4748) );
  NAND2_X1 U6199 ( .A1(n6592), .A2(n5715), .ZN(n6696) );
  NOR2_X1 U6200 ( .A1(n6697), .A2(n4758), .ZN(n4757) );
  INV_X1 U6201 ( .A(n5715), .ZN(n4758) );
  INV_X1 U6202 ( .A(n6025), .ZN(n4759) );
  NAND2_X1 U6203 ( .A1(n5958), .A2(n5957), .ZN(n8320) );
  NOR2_X1 U6204 ( .A1(n5977), .A2(n5956), .ZN(n4766) );
  AND2_X1 U6205 ( .A1(n5670), .A2(n5656), .ZN(n4767) );
  NAND3_X1 U6206 ( .A1(n4769), .A2(n8427), .A3(n4768), .ZN(n8426) );
  NAND2_X1 U6207 ( .A1(n5581), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5534) );
  NAND2_X1 U6208 ( .A1(n8160), .A2(n8159), .ZN(n4771) );
  NAND2_X1 U6209 ( .A1(n7671), .A2(n7673), .ZN(n8159) );
  NAND2_X1 U6210 ( .A1(n5413), .A2(n6619), .ZN(n4772) );
  NAND2_X1 U6211 ( .A1(n7946), .A2(n4776), .ZN(n4775) );
  OAI21_X1 U6212 ( .B1(n7946), .B2(n5452), .A(n5451), .ZN(n7935) );
  NAND2_X1 U6213 ( .A1(n4785), .A2(n4786), .ZN(n7923) );
  NAND2_X1 U6214 ( .A1(n4795), .A2(n4793), .ZN(n5430) );
  NAND2_X1 U6215 ( .A1(n5433), .A2(n4802), .ZN(n4801) );
  NAND3_X1 U6216 ( .A1(n4304), .A2(n4803), .A3(n4805), .ZN(n4800) );
  NAND2_X1 U6217 ( .A1(n4812), .A2(n4811), .ZN(n5448) );
  OAI21_X2 U6218 ( .B1(n5440), .B2(n4815), .A(n4813), .ZN(n8023) );
  INV_X1 U6219 ( .A(n8566), .ZN(n8926) );
  NAND2_X1 U6220 ( .A1(n8532), .A2(n4252), .ZN(n8539) );
  NAND2_X1 U6221 ( .A1(n5367), .A2(n5366), .ZN(n5369) );
  XNOR2_X1 U6222 ( .A(n5367), .B(n5366), .ZN(n6104) );
  AOI21_X1 U6223 ( .B1(n8709), .B2(n4832), .A(n8715), .ZN(n8710) );
  NAND2_X1 U6224 ( .A1(n5294), .A2(n5293), .ZN(n5311) );
  NAND2_X1 U6225 ( .A1(n5294), .A2(n5282), .ZN(n7221) );
  NAND2_X1 U6226 ( .A1(n5470), .A2(n5469), .ZN(n6329) );
  OR2_X1 U6227 ( .A1(n7111), .A2(n6974), .ZN(n9696) );
  INV_X1 U6228 ( .A(n9159), .ZN(n9160) );
  OR2_X1 U6229 ( .A1(n6329), .A2(n5483), .ZN(n5511) );
  OR2_X1 U6230 ( .A1(n6329), .A2(P2_D_REG_1__SCAN_IN), .ZN(n5472) );
  OAI21_X1 U6231 ( .B1(n6329), .B2(P2_D_REG_0__SCAN_IN), .A(n6348), .ZN(n6642)
         );
  AOI22_X2 U6232 ( .A1(n7462), .A2(n7461), .B1(n7426), .B2(n7532), .ZN(n7529)
         );
  NOR2_X1 U6233 ( .A1(n5504), .A2(n5503), .ZN(n6212) );
  NOR2_X1 U6234 ( .A1(n5502), .A2(n5501), .ZN(n5503) );
  OR2_X1 U6235 ( .A1(n5502), .A2(n7306), .ZN(n5498) );
  NAND2_X1 U6236 ( .A1(n5415), .A2(n4891), .ZN(n7671) );
  INV_X2 U6237 ( .A(n4261), .ZN(n4971) );
  NAND2_X1 U6238 ( .A1(n4849), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4856) );
  NAND2_X1 U6239 ( .A1(n4264), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5606) );
  NAND2_X2 U6240 ( .A1(n7394), .A2(n8278), .ZN(n4908) );
  NOR2_X1 U6241 ( .A1(n5758), .A2(n5743), .ZN(n4820) );
  AND2_X1 U6242 ( .A1(n7469), .A2(n7821), .ZN(n4821) );
  OR2_X1 U6243 ( .A1(n4864), .A2(n7842), .ZN(n4823) );
  INV_X1 U6244 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5850) );
  INV_X1 U6245 ( .A(n9360), .ZN(n9406) );
  INV_X1 U6246 ( .A(n6150), .ZN(n6151) );
  NOR2_X1 U6247 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(n5552), .ZN(n4824) );
  AND2_X1 U6248 ( .A1(n6267), .A2(n6266), .ZN(n4827) );
  INV_X1 U6249 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5019) );
  AND2_X1 U6250 ( .A1(n5029), .A2(n5015), .ZN(n4828) );
  OR2_X1 U6251 ( .A1(n8207), .A2(n7961), .ZN(n4829) );
  AND2_X1 U6252 ( .A1(n6268), .A2(n4827), .ZN(n4830) );
  NAND2_X1 U6253 ( .A1(n4262), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n4831) );
  INV_X1 U6254 ( .A(n8725), .ZN(n8872) );
  INV_X1 U6255 ( .A(n7555), .ZN(n7825) );
  INV_X1 U6256 ( .A(n9408), .ZN(n8871) );
  CLKBUF_X3 U6257 ( .A(n5657), .Z(n6134) );
  OR2_X1 U6258 ( .A1(n8708), .A2(n8707), .ZN(n4832) );
  INV_X1 U6259 ( .A(n8563), .ZN(n8866) );
  INV_X2 U6260 ( .A(n9969), .ZN(n9967) );
  INV_X1 U6261 ( .A(n9982), .ZN(n6211) );
  INV_X1 U6262 ( .A(n6347), .ZN(n6331) );
  INV_X1 U6263 ( .A(n8570), .ZN(n8573) );
  NAND2_X1 U6264 ( .A1(n8537), .A2(n8561), .ZN(n8538) );
  NAND2_X1 U6265 ( .A1(n8539), .A2(n8538), .ZN(n8541) );
  INV_X1 U6266 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n4835) );
  NOR2_X1 U6267 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n4837) );
  NOR2_X1 U6268 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n4838) );
  INV_X1 U6269 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5526) );
  INV_X1 U6270 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n4844) );
  INV_X1 U6271 ( .A(n5773), .ZN(n5774) );
  INV_X1 U6272 ( .A(n6953), .ZN(n6952) );
  INV_X1 U6273 ( .A(n7701), .ZN(n5423) );
  NOR2_X1 U6274 ( .A1(n5955), .A2(n5954), .ZN(n5956) );
  NAND2_X1 U6275 ( .A1(n5772), .A2(n5774), .ZN(n5775) );
  INV_X1 U6276 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5531) );
  INV_X1 U6277 ( .A(n7635), .ZN(n5027) );
  INV_X1 U6278 ( .A(n5956), .ZN(n5957) );
  NAND2_X1 U6279 ( .A1(n5593), .A2(n5592), .ZN(n5596) );
  INV_X1 U6280 ( .A(n6030), .ZN(n6029) );
  INV_X1 U6281 ( .A(n5923), .ZN(n5921) );
  INV_X1 U6282 ( .A(n8735), .ZN(n6437) );
  NAND2_X1 U6283 ( .A1(n5381), .A2(n5380), .ZN(n5385) );
  INV_X1 U6284 ( .A(n5564), .ZN(n5561) );
  INV_X1 U6285 ( .A(SI_9_), .ZN(n9111) );
  AND2_X1 U6286 ( .A1(n7437), .A2(n7986), .ZN(n7438) );
  INV_X1 U6287 ( .A(n7409), .ZN(n7410) );
  NOR2_X1 U6288 ( .A1(n7685), .A2(n7698), .ZN(n4969) );
  INV_X1 U6289 ( .A(n7744), .ZN(n5185) );
  AND2_X1 U6290 ( .A1(n5720), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5742) );
  AND2_X1 U6291 ( .A1(n6068), .A2(n6066), .ZN(n8365) );
  NAND2_X1 U6292 ( .A1(n5960), .A2(n4263), .ZN(n6172) );
  OR2_X1 U6293 ( .A1(n6087), .A2(n6086), .ZN(n6109) );
  OR2_X1 U6294 ( .A1(n6051), .A2(n6050), .ZN(n6072) );
  OR2_X1 U6295 ( .A1(n5980), .A2(n8379), .ZN(n5996) );
  INV_X1 U6296 ( .A(n9380), .ZN(n6228) );
  INV_X1 U6297 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5842) );
  OR2_X1 U6298 ( .A1(n7420), .A2(n7419), .ZN(n7421) );
  INV_X1 U6299 ( .A(n8162), .ZN(n6955) );
  INV_X1 U6300 ( .A(n4913), .ZN(n5390) );
  OR2_X1 U6301 ( .A1(n5373), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5494) );
  NAND2_X1 U6302 ( .A1(n5358), .A2(n5357), .ZN(n5373) );
  AOI21_X1 U6303 ( .B1(n7128), .B2(n4970), .A(n4969), .ZN(n7148) );
  AND2_X2 U6304 ( .A1(n7814), .A2(n6643), .ZN(n7801) );
  AND2_X1 U6305 ( .A1(n9897), .A2(n9966), .ZN(n6201) );
  OR2_X1 U6306 ( .A1(n6642), .A2(n6322), .ZN(n5506) );
  XOR2_X1 U6307 ( .A(n7624), .B(n7650), .Z(n5502) );
  INV_X1 U6308 ( .A(n8167), .ZN(n8037) );
  NOR2_X1 U6309 ( .A1(n6639), .A2(n6321), .ZN(n6668) );
  NAND2_X1 U6310 ( .A1(n5870), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5889) );
  INV_X1 U6311 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5782) );
  OR2_X1 U6312 ( .A1(n5996), .A2(n8334), .ZN(n6014) );
  OR2_X1 U6313 ( .A1(n5903), .A2(n5902), .ZN(n5923) );
  NAND2_X1 U6314 ( .A1(n5758), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5783) );
  INV_X1 U6315 ( .A(n9165), .ZN(n8887) );
  OR2_X1 U6316 ( .A1(n5641), .A2(n4880), .ZN(n5622) );
  NAND2_X1 U6317 ( .A1(n5887), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5903) );
  AND2_X1 U6318 ( .A1(n6109), .A2(n6088), .ZN(n8970) );
  INV_X1 U6319 ( .A(n9648), .ZN(n9632) );
  OR2_X1 U6320 ( .A1(n6540), .A2(n8749), .ZN(n9654) );
  INV_X1 U6321 ( .A(n9232), .ZN(n9248) );
  INV_X1 U6322 ( .A(n8724), .ZN(n9284) );
  INV_X1 U6323 ( .A(n8620), .ZN(n9297) );
  NOR2_X1 U6324 ( .A1(n9308), .A2(n8646), .ZN(n6188) );
  AND2_X1 U6325 ( .A1(n6247), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6679) );
  AND2_X1 U6326 ( .A1(n6526), .A2(n8640), .ZN(n9222) );
  OR2_X1 U6327 ( .A1(n6788), .A2(n8485), .ZN(n6913) );
  INV_X1 U6328 ( .A(n9224), .ZN(n9285) );
  NAND2_X1 U6329 ( .A1(n6438), .A2(n8570), .ZN(n6449) );
  AND2_X1 U6330 ( .A1(n5332), .A2(n5317), .ZN(n5330) );
  INV_X1 U6331 ( .A(n7598), .ZN(n7573) );
  INV_X1 U6332 ( .A(n7888), .ZN(n7913) );
  AND3_X1 U6333 ( .A1(n5252), .A2(n5251), .A3(n5250), .ZN(n7430) );
  OR2_X1 U6334 ( .A1(n4913), .A2(n4886), .ZN(n4889) );
  OR2_X1 U6335 ( .A1(n6360), .A2(n6359), .ZN(n9875) );
  INV_X1 U6336 ( .A(n9720), .ZN(n9874) );
  OR2_X1 U6337 ( .A1(n9897), .A2(n9948), .ZN(n8096) );
  AND2_X1 U6338 ( .A1(n7768), .A2(n7770), .ZN(n7983) );
  AND2_X1 U6339 ( .A1(n6669), .A2(n7801), .ZN(n8092) );
  INV_X1 U6340 ( .A(n7955), .ZN(n8086) );
  INV_X1 U6341 ( .A(n8126), .ZN(n8152) );
  AND2_X1 U6342 ( .A1(n6204), .A2(n6203), .ZN(n6205) );
  AND2_X1 U6343 ( .A1(n7917), .A2(n7916), .ZN(n8181) );
  AND2_X1 U6344 ( .A1(n9897), .A2(n7663), .ZN(n9953) );
  NAND2_X1 U6345 ( .A1(n5501), .A2(n7155), .ZN(n9962) );
  OR2_X1 U6346 ( .A1(n6665), .A2(n5510), .ZN(n5514) );
  OR2_X1 U6347 ( .A1(n5783), .A2(n5782), .ZN(n5801) );
  OR2_X1 U6348 ( .A1(n8983), .A2(n6111), .ZN(n6079) );
  INV_X1 U6349 ( .A(n4265), .ZN(n6137) );
  INV_X1 U6350 ( .A(n9645), .ZN(n9595) );
  AND2_X1 U6351 ( .A1(n6552), .A2(n8748), .ZN(n9648) );
  AND2_X1 U6352 ( .A1(n8494), .A2(n8493), .ZN(n7203) );
  INV_X1 U6353 ( .A(n9283), .ZN(n9301) );
  INV_X1 U6354 ( .A(n9315), .ZN(n9005) );
  AND2_X1 U6355 ( .A1(n9708), .A2(n9675), .ZN(n9360) );
  AND2_X1 U6356 ( .A1(n6171), .A2(n8651), .ZN(n6345) );
  AND2_X1 U6357 ( .A1(n9701), .A2(n9675), .ZN(n9453) );
  AND2_X1 U6358 ( .A1(n6255), .A2(n6678), .ZN(n9479) );
  AND2_X1 U6359 ( .A1(n5779), .A2(n5795), .ZN(n9532) );
  INV_X1 U6360 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5819) );
  AND2_X1 U6361 ( .A1(n6641), .A2(n6640), .ZN(n7558) );
  AND2_X1 U6362 ( .A1(n7621), .A2(n5395), .ZN(n7655) );
  INV_X1 U6363 ( .A(n7550), .ZN(n8000) );
  INV_X1 U6364 ( .A(n7419), .ZN(n8094) );
  OR2_X1 U6365 ( .A1(P2_U3150), .A2(n6356), .ZN(n9720) );
  OR2_X1 U6366 ( .A1(n5495), .A2(n8096), .ZN(n7955) );
  INV_X1 U6367 ( .A(n8065), .ZN(n8105) );
  NAND2_X1 U6368 ( .A1(n5495), .A2(n9896), .ZN(n8098) );
  NAND2_X1 U6369 ( .A1(n9982), .A2(n9962), .ZN(n8155) );
  AND2_X2 U6370 ( .A1(n6206), .A2(n6205), .ZN(n9982) );
  NAND2_X1 U6371 ( .A1(n9967), .A2(n9966), .ZN(n8212) );
  NAND2_X1 U6372 ( .A1(n9967), .A2(n9962), .ZN(n8266) );
  AND2_X1 U6373 ( .A1(n5514), .A2(n5513), .ZN(n9969) );
  AND2_X1 U6374 ( .A1(n6637), .A2(n6329), .ZN(n6347) );
  AND2_X1 U6375 ( .A1(n6630), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6350) );
  INV_X1 U6376 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6586) );
  INV_X1 U6377 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6327) );
  INV_X1 U6378 ( .A(n9447), .ZN(n9014) );
  INV_X1 U6379 ( .A(n7175), .ZN(n7237) );
  NAND2_X1 U6380 ( .A1(n6116), .A2(n6115), .ZN(n8721) );
  NAND2_X1 U6381 ( .A1(n6037), .A2(n6036), .ZN(n9166) );
  OR2_X1 U6382 ( .A1(n6540), .A2(n6527), .ZN(n9645) );
  NAND2_X1 U6383 ( .A1(n9306), .A2(n6702), .ZN(n9294) );
  NAND2_X1 U6384 ( .A1(n8563), .A2(n9360), .ZN(n6252) );
  INV_X1 U6385 ( .A(n9706), .ZN(n9403) );
  INV_X1 U6386 ( .A(n9706), .ZN(n9708) );
  INV_X1 U6387 ( .A(n9453), .ZN(n9483) );
  INV_X1 U6388 ( .A(n9479), .ZN(n9699) );
  INV_X1 U6389 ( .A(n9699), .ZN(n9701) );
  NAND2_X1 U6390 ( .A1(n9487), .A2(n9486), .ZN(n9667) );
  INV_X1 U6391 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6712) );
  INV_X1 U6392 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9022) );
  INV_X1 U6393 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6306) );
  INV_X1 U6394 ( .A(n7833), .ZN(P2_U3893) );
  NAND4_X1 U6395 ( .A1(n4844), .A2(n9089), .A3(n5459), .A4(n5486), .ZN(n4845)
         );
  XNOR2_X2 U6396 ( .A(n4848), .B(P2_IR_REG_30__SCAN_IN), .ZN(n4851) );
  INV_X1 U6397 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n4850) );
  OR2_X1 U6398 ( .A1(n4908), .A2(n4850), .ZN(n4855) );
  INV_X1 U6399 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6723) );
  OR2_X1 U6400 ( .A1(n4913), .A2(n6723), .ZN(n4854) );
  NAND2_X1 U6401 ( .A1(n4931), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4853) );
  XNOR2_X2 U6402 ( .A(n4858), .B(n4857), .ZN(n7811) );
  INV_X1 U6403 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4861) );
  NAND2_X1 U6404 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4860) );
  INV_X1 U6405 ( .A(n6396), .ZN(n7842) );
  NAND2_X2 U6406 ( .A1(n4864), .A2(n6276), .ZN(n5006) );
  AND2_X1 U6407 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4862) );
  NAND2_X1 U6408 ( .A1(n4879), .A2(n4862), .ZN(n5600) );
  NAND2_X1 U6409 ( .A1(n5600), .A2(n4863), .ZN(n4874) );
  XNOR2_X1 U6410 ( .A(n4873), .B(n4874), .ZN(n5575) );
  OR2_X1 U6411 ( .A1(n5006), .A2(n5575), .ZN(n4866) );
  NAND2_X4 U6412 ( .A1(n4864), .A2(n6281), .ZN(n7609) );
  NAND2_X1 U6413 ( .A1(n5249), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n4870) );
  INV_X1 U6414 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6716) );
  OR2_X1 U6415 ( .A1(n4913), .A2(n6716), .ZN(n4869) );
  INV_X1 U6416 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6394) );
  OR2_X1 U6417 ( .A1(n7615), .A2(n6394), .ZN(n4868) );
  NAND2_X1 U6418 ( .A1(n6276), .A2(SI_0_), .ZN(n4871) );
  XNOR2_X1 U6419 ( .A(n4871), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8279) );
  MUX2_X1 U6420 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8279), .S(n4864), .Z(n6470) );
  NAND2_X1 U6421 ( .A1(n6721), .A2(n6470), .ZN(n7661) );
  NAND2_X1 U6422 ( .A1(n6618), .A2(n7665), .ZN(n8157) );
  INV_X1 U6423 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6277) );
  OR2_X1 U6424 ( .A1(n7609), .A2(n6277), .ZN(n4885) );
  INV_X1 U6425 ( .A(n4873), .ZN(n4875) );
  NAND2_X1 U6426 ( .A1(n4875), .A2(n4874), .ZN(n4878) );
  NAND2_X1 U6427 ( .A1(n4876), .A2(SI_1_), .ZN(n4877) );
  INV_X1 U6428 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n4880) );
  XNOR2_X1 U6429 ( .A(n4901), .B(SI_2_), .ZN(n4899) );
  XNOR2_X1 U6430 ( .A(n4900), .B(n4899), .ZN(n6285) );
  OR2_X1 U6431 ( .A1(n5006), .A2(n6285), .ZN(n4884) );
  NAND2_X1 U6432 ( .A1(n6274), .A2(n4250), .ZN(n4883) );
  NAND2_X1 U6433 ( .A1(n5249), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n4890) );
  INV_X1 U6434 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n4886) );
  NAND2_X1 U6435 ( .A1(n4849), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4888) );
  NAND2_X1 U6436 ( .A1(n7832), .A2(n8171), .ZN(n7673) );
  NAND2_X1 U6437 ( .A1(n8157), .A2(n8156), .ZN(n4892) );
  NAND2_X1 U6438 ( .A1(n4892), .A2(n7671), .ZN(n7059) );
  NAND2_X1 U6439 ( .A1(n4261), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4896) );
  NAND2_X1 U6440 ( .A1(n5408), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4895) );
  NAND2_X1 U6441 ( .A1(n5249), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n4894) );
  OR2_X1 U6442 ( .A1(n4913), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n4893) );
  NAND4_X1 U6443 ( .A1(n4896), .A2(n4895), .A3(n4894), .A4(n4893), .ZN(n8162)
         );
  NAND2_X1 U6444 ( .A1(n4897), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4898) );
  XNOR2_X1 U6445 ( .A(n4898), .B(n4834), .ZN(n6481) );
  INV_X1 U6446 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6278) );
  OR2_X1 U6447 ( .A1(n7609), .A2(n6278), .ZN(n4907) );
  NAND2_X1 U6448 ( .A1(n4900), .A2(n4899), .ZN(n4904) );
  INV_X1 U6449 ( .A(n4901), .ZN(n4902) );
  NAND2_X1 U6450 ( .A1(n4902), .A2(SI_2_), .ZN(n4903) );
  NAND2_X1 U6451 ( .A1(n4904), .A2(n4903), .ZN(n4922) );
  INV_X1 U6452 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n4905) );
  MUX2_X1 U6453 ( .A(n6278), .B(n4905), .S(n4879), .Z(n4923) );
  XNOR2_X1 U6454 ( .A(n4923), .B(SI_3_), .ZN(n4921) );
  XNOR2_X1 U6455 ( .A(n4922), .B(n4921), .ZN(n6283) );
  OR2_X1 U6456 ( .A1(n5006), .A2(n6283), .ZN(n4906) );
  OAI211_X1 U6457 ( .C1(n4864), .C2(n6481), .A(n4907), .B(n4906), .ZN(n7063)
         );
  XNOR2_X1 U6458 ( .A(n8162), .B(n7063), .ZN(n7060) );
  NAND2_X1 U6459 ( .A1(n7059), .A2(n7060), .ZN(n7082) );
  NAND2_X1 U6460 ( .A1(n6955), .A2(n7063), .ZN(n7693) );
  NAND2_X1 U6461 ( .A1(n4261), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4917) );
  INV_X1 U6462 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n4909) );
  NAND2_X1 U6463 ( .A1(n4911), .A2(n4910), .ZN(n4935) );
  NAND2_X1 U6464 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n4912) );
  AND2_X1 U6465 ( .A1(n4935), .A2(n4912), .ZN(n6958) );
  OR2_X1 U6466 ( .A1(n4913), .A2(n6958), .ZN(n4915) );
  INV_X1 U6467 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7094) );
  OR2_X1 U6468 ( .A1(n7615), .A2(n7094), .ZN(n4914) );
  NAND2_X1 U6469 ( .A1(n4918), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4920) );
  INV_X1 U6470 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4919) );
  XNOR2_X1 U6471 ( .A(n4920), .B(n4919), .ZN(n6607) );
  INV_X1 U6472 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6279) );
  OR2_X1 U6473 ( .A1(n7609), .A2(n6279), .ZN(n4928) );
  NAND2_X1 U6474 ( .A1(n4922), .A2(n4921), .ZN(n4926) );
  INV_X1 U6475 ( .A(n4923), .ZN(n4924) );
  NAND2_X1 U6476 ( .A1(n4924), .A2(SI_3_), .ZN(n4925) );
  NAND2_X1 U6477 ( .A1(n4926), .A2(n4925), .ZN(n4945) );
  INV_X1 U6478 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6304) );
  XNOR2_X1 U6479 ( .A(n4946), .B(SI_4_), .ZN(n4944) );
  XNOR2_X1 U6480 ( .A(n4945), .B(n4944), .ZN(n6303) );
  OR2_X1 U6481 ( .A1(n5006), .A2(n6303), .ZN(n4927) );
  OAI211_X1 U6482 ( .C1(n4864), .C2(n6607), .A(n4928), .B(n4927), .ZN(n7096)
         );
  NAND2_X1 U6483 ( .A1(n7144), .A2(n7096), .ZN(n7681) );
  AND2_X1 U6484 ( .A1(n7693), .A2(n7681), .ZN(n4929) );
  NAND2_X1 U6485 ( .A1(n7082), .A2(n4929), .ZN(n7128) );
  INV_X1 U6486 ( .A(n7681), .ZN(n4930) );
  INV_X1 U6487 ( .A(n7096), .ZN(n9918) );
  NAND2_X1 U6488 ( .A1(n7831), .A2(n9918), .ZN(n7694) );
  OR2_X1 U6489 ( .A1(n4930), .A2(n7678), .ZN(n7127) );
  NAND2_X1 U6490 ( .A1(n5249), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n4940) );
  INV_X1 U6491 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n4932) );
  INV_X1 U6492 ( .A(n4935), .ZN(n4934) );
  NAND2_X1 U6493 ( .A1(n4934), .A2(n4933), .ZN(n4952) );
  NAND2_X1 U6494 ( .A1(n4935), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n4936) );
  AND2_X1 U6495 ( .A1(n4952), .A2(n4936), .ZN(n7141) );
  OR2_X1 U6496 ( .A1(n4913), .A2(n7141), .ZN(n4938) );
  INV_X1 U6497 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6610) );
  OR2_X1 U6498 ( .A1(n7615), .A2(n6610), .ZN(n4937) );
  AND4_X2 U6499 ( .A1(n4940), .A2(n4939), .A3(n4938), .A4(n4937), .ZN(n7105)
         );
  OR2_X1 U6500 ( .A1(n4941), .A2(n5169), .ZN(n4943) );
  XNOR2_X1 U6501 ( .A(n4943), .B(n4942), .ZN(n6847) );
  NAND2_X1 U6502 ( .A1(n4945), .A2(n4944), .ZN(n4949) );
  INV_X1 U6503 ( .A(n4946), .ZN(n4947) );
  NAND2_X1 U6504 ( .A1(n4947), .A2(SI_4_), .ZN(n4948) );
  XNOR2_X1 U6505 ( .A(n4963), .B(SI_5_), .ZN(n4961) );
  XNOR2_X1 U6506 ( .A(n4962), .B(n4961), .ZN(n6305) );
  OR2_X1 U6507 ( .A1(n5006), .A2(n6305), .ZN(n4951) );
  OR2_X1 U6508 ( .A1(n7609), .A2(n6286), .ZN(n4950) );
  OAI211_X1 U6509 ( .C1(n4864), .C2(n6847), .A(n4951), .B(n4950), .ZN(n7039)
         );
  NAND2_X1 U6510 ( .A1(n7105), .A2(n7039), .ZN(n7129) );
  INV_X1 U6511 ( .A(n7039), .ZN(n9921) );
  NAND2_X1 U6512 ( .A1(n7830), .A2(n9921), .ZN(n7695) );
  NAND2_X1 U6513 ( .A1(n5249), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n4957) );
  OR2_X1 U6514 ( .A1(n4971), .A2(n9974), .ZN(n4956) );
  NAND2_X1 U6515 ( .A1(n4952), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n4953) );
  AND2_X1 U6516 ( .A1(n4974), .A2(n4953), .ZN(n7134) );
  OR2_X1 U6517 ( .A1(n4913), .A2(n7134), .ZN(n4955) );
  INV_X1 U6518 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7133) );
  OR2_X1 U6519 ( .A1(n7615), .A2(n7133), .ZN(n4954) );
  NAND2_X1 U6520 ( .A1(n4958), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4960) );
  INV_X1 U6521 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n4959) );
  XNOR2_X1 U6522 ( .A(n4960), .B(n4959), .ZN(n7253) );
  INV_X1 U6523 ( .A(n4963), .ZN(n4964) );
  NAND2_X1 U6524 ( .A1(n4964), .A2(SI_5_), .ZN(n4965) );
  INV_X1 U6525 ( .A(SI_6_), .ZN(n9076) );
  XNOR2_X1 U6526 ( .A(n4985), .B(n9076), .ZN(n4983) );
  XNOR2_X1 U6527 ( .A(n4984), .B(n4983), .ZN(n6301) );
  OR2_X1 U6528 ( .A1(n5006), .A2(n6301), .ZN(n4967) );
  OR2_X1 U6529 ( .A1(n7609), .A2(n4361), .ZN(n4966) );
  OAI211_X1 U6530 ( .C1(n4864), .C2(n7253), .A(n4967), .B(n4966), .ZN(n7136)
         );
  INV_X1 U6531 ( .A(n7136), .ZN(n9927) );
  NAND2_X1 U6532 ( .A1(n7829), .A2(n9927), .ZN(n7688) );
  AND2_X1 U6533 ( .A1(n7633), .A2(n7688), .ZN(n4968) );
  AND2_X1 U6534 ( .A1(n7127), .A2(n4968), .ZN(n4970) );
  INV_X1 U6535 ( .A(n7688), .ZN(n7685) );
  NAND2_X1 U6536 ( .A1(n7188), .A2(n7136), .ZN(n7683) );
  AND2_X1 U6537 ( .A1(n7129), .A2(n7683), .ZN(n7698) );
  NAND2_X1 U6538 ( .A1(n5249), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n4980) );
  INV_X1 U6539 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7259) );
  OR2_X1 U6540 ( .A1(n4971), .A2(n7259), .ZN(n4979) );
  NAND2_X1 U6541 ( .A1(n4974), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n4975) );
  AND2_X1 U6542 ( .A1(n4991), .A2(n4975), .ZN(n7191) );
  OR2_X1 U6543 ( .A1(n4913), .A2(n7191), .ZN(n4978) );
  INV_X1 U6544 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n4976) );
  OR2_X1 U6545 ( .A1(n7615), .A2(n4976), .ZN(n4977) );
  NAND2_X1 U6546 ( .A1(n4291), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4981) );
  MUX2_X1 U6547 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4981), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n4982) );
  NAND2_X1 U6548 ( .A1(n4982), .A2(n5016), .ZN(n7256) );
  NAND2_X1 U6549 ( .A1(n4985), .A2(SI_6_), .ZN(n4986) );
  INV_X1 U6550 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6308) );
  INV_X1 U6551 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n4987) );
  MUX2_X1 U6552 ( .A(n6308), .B(n4987), .S(n6281), .Z(n4999) );
  XNOR2_X1 U6553 ( .A(n4999), .B(SI_7_), .ZN(n4997) );
  OR2_X1 U6554 ( .A1(n6309), .A2(n5006), .ZN(n4989) );
  OR2_X1 U6555 ( .A1(n7609), .A2(n6308), .ZN(n4988) );
  OAI211_X1 U6556 ( .C1(n4864), .C2(n7256), .A(n4989), .B(n4988), .ZN(n7182)
         );
  NAND2_X1 U6557 ( .A1(n7282), .A2(n7182), .ZN(n7713) );
  INV_X1 U6558 ( .A(n7182), .ZN(n9932) );
  NAND2_X1 U6559 ( .A1(n7828), .A2(n9932), .ZN(n7708) );
  NAND2_X1 U6560 ( .A1(n7148), .A2(n7701), .ZN(n7149) );
  NAND2_X1 U6561 ( .A1(n7149), .A2(n7708), .ZN(n7211) );
  NAND2_X1 U6562 ( .A1(n5249), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n4996) );
  INV_X1 U6563 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n4990) );
  OR2_X1 U6564 ( .A1(n4971), .A2(n4990), .ZN(n4995) );
  NAND2_X1 U6565 ( .A1(n5408), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4994) );
  NAND2_X1 U6566 ( .A1(n4991), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n4992) );
  AND2_X1 U6567 ( .A1(n5021), .A2(n4992), .ZN(n7285) );
  OR2_X1 U6568 ( .A1(n4913), .A2(n7285), .ZN(n4993) );
  NAND4_X1 U6569 ( .A1(n4996), .A2(n4995), .A3(n4994), .A4(n4993), .ZN(n7827)
         );
  INV_X1 U6570 ( .A(n4999), .ZN(n5000) );
  NAND2_X1 U6571 ( .A1(n5000), .A2(SI_7_), .ZN(n5001) );
  INV_X1 U6572 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6312) );
  MUX2_X1 U6573 ( .A(n6312), .B(n6311), .S(n6281), .Z(n5003) );
  INV_X1 U6574 ( .A(SI_8_), .ZN(n5002) );
  NAND2_X1 U6575 ( .A1(n5003), .A2(n5002), .ZN(n5010) );
  INV_X1 U6576 ( .A(n5003), .ZN(n5004) );
  NAND2_X1 U6577 ( .A1(n5004), .A2(SI_8_), .ZN(n5005) );
  NAND2_X1 U6578 ( .A1(n5010), .A2(n5005), .ZN(n5011) );
  NAND2_X1 U6579 ( .A1(n6310), .A2(n5387), .ZN(n5009) );
  NAND2_X1 U6580 ( .A1(n5016), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5007) );
  AOI22_X1 U6581 ( .A1(n7606), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6274), .B2(
        n9743), .ZN(n5008) );
  AND2_X1 U6582 ( .A1(n7827), .A2(n9937), .ZN(n7711) );
  NAND2_X1 U6583 ( .A1(n7339), .A2(n7294), .ZN(n7692) );
  MUX2_X1 U6584 ( .A(n6327), .B(n6324), .S(n6281), .Z(n5013) );
  NAND2_X1 U6585 ( .A1(n5013), .A2(n9111), .ZN(n5029) );
  INV_X1 U6586 ( .A(n5013), .ZN(n5014) );
  NAND2_X1 U6587 ( .A1(n5014), .A2(SI_9_), .ZN(n5015) );
  XNOR2_X1 U6588 ( .A(n5028), .B(n4828), .ZN(n6323) );
  NAND2_X1 U6589 ( .A1(n6323), .A2(n5387), .ZN(n5018) );
  OR2_X1 U6590 ( .A1(n5057), .A2(n5169), .ZN(n5033) );
  XNOR2_X1 U6591 ( .A(n5033), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7261) );
  AOI22_X1 U6592 ( .A1(n7606), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6274), .B2(
        n7261), .ZN(n5017) );
  NAND2_X1 U6593 ( .A1(n5249), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5026) );
  NAND2_X1 U6594 ( .A1(n4262), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5025) );
  NAND2_X1 U6595 ( .A1(n5408), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5024) );
  NAND2_X1 U6596 ( .A1(n5021), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5022) );
  AND2_X1 U6597 ( .A1(n5039), .A2(n5022), .ZN(n7337) );
  OR2_X1 U6598 ( .A1(n4913), .A2(n7337), .ZN(n5023) );
  NAND4_X1 U6599 ( .A1(n5026), .A2(n5025), .A3(n5024), .A4(n5023), .ZN(n7826)
         );
  NAND2_X1 U6600 ( .A1(n9942), .A2(n7826), .ZN(n7690) );
  INV_X1 U6601 ( .A(n9942), .ZN(n7349) );
  NAND2_X1 U6602 ( .A1(n7349), .A2(n7378), .ZN(n7702) );
  NAND2_X1 U6603 ( .A1(n7690), .A2(n7702), .ZN(n7635) );
  INV_X1 U6604 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5031) );
  MUX2_X1 U6605 ( .A(n9046), .B(n5031), .S(n6281), .Z(n5047) );
  XNOR2_X1 U6606 ( .A(n5047), .B(SI_10_), .ZN(n5046) );
  XNOR2_X1 U6607 ( .A(n5051), .B(n5046), .ZN(n6325) );
  NAND2_X1 U6608 ( .A1(n6325), .A2(n5387), .ZN(n5037) );
  INV_X1 U6609 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5032) );
  NAND2_X1 U6610 ( .A1(n5033), .A2(n5032), .ZN(n5034) );
  NAND2_X1 U6611 ( .A1(n5034), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5035) );
  XNOR2_X1 U6612 ( .A(n5035), .B(P2_IR_REG_10__SCAN_IN), .ZN(n9761) );
  AOI22_X1 U6613 ( .A1(n7606), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6274), .B2(
        n9761), .ZN(n5036) );
  NAND2_X1 U6614 ( .A1(n5249), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5044) );
  INV_X1 U6615 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n5038) );
  OR2_X1 U6616 ( .A1(n4971), .A2(n5038), .ZN(n5043) );
  NAND2_X1 U6617 ( .A1(n5039), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5040) );
  AND2_X1 U6618 ( .A1(n5065), .A2(n5040), .ZN(n7375) );
  OR2_X1 U6619 ( .A1(n4913), .A2(n7375), .ZN(n5042) );
  INV_X1 U6620 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7276) );
  OR2_X1 U6621 ( .A1(n7615), .A2(n7276), .ZN(n5041) );
  OR2_X1 U6622 ( .A1(n9947), .A2(n7555), .ZN(n7719) );
  NAND2_X1 U6623 ( .A1(n9947), .A2(n7555), .ZN(n7720) );
  NAND2_X1 U6624 ( .A1(n7719), .A2(n7720), .ZN(n7636) );
  INV_X1 U6625 ( .A(n7690), .ZN(n7704) );
  NOR2_X1 U6626 ( .A1(n7636), .A2(n7704), .ZN(n5045) );
  NAND2_X1 U6627 ( .A1(n7270), .A2(n7720), .ZN(n7313) );
  INV_X1 U6628 ( .A(n5046), .ZN(n5050) );
  INV_X1 U6629 ( .A(n5047), .ZN(n5048) );
  NAND2_X1 U6630 ( .A1(n5048), .A2(SI_10_), .ZN(n5049) );
  MUX2_X1 U6631 ( .A(n6333), .B(n9022), .S(n6281), .Z(n5053) );
  INV_X1 U6632 ( .A(SI_11_), .ZN(n5052) );
  NAND2_X1 U6633 ( .A1(n5053), .A2(n5052), .ZN(n5071) );
  INV_X1 U6634 ( .A(n5053), .ZN(n5054) );
  NAND2_X1 U6635 ( .A1(n5054), .A2(SI_11_), .ZN(n5055) );
  NAND2_X1 U6636 ( .A1(n5071), .A2(n5055), .ZN(n5072) );
  XNOR2_X1 U6637 ( .A(n5073), .B(n5072), .ZN(n6332) );
  NOR2_X1 U6638 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5056) );
  NOR2_X1 U6639 ( .A1(n5060), .A2(n5169), .ZN(n5058) );
  MUX2_X1 U6640 ( .A(n5169), .B(n5058), .S(P2_IR_REG_11__SCAN_IN), .Z(n5062)
         );
  NAND2_X1 U6641 ( .A1(n5060), .A2(n5059), .ZN(n5090) );
  INV_X1 U6642 ( .A(n5090), .ZN(n5061) );
  AOI22_X1 U6643 ( .A1(n7606), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6274), .B2(
        n9778), .ZN(n5063) );
  INV_X1 U6644 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n5064) );
  OR2_X1 U6645 ( .A1(n4971), .A2(n5064), .ZN(n5070) );
  NAND2_X1 U6646 ( .A1(n5408), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5069) );
  NAND2_X1 U6647 ( .A1(n5249), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5068) );
  NAND2_X1 U6648 ( .A1(n5065), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5066) );
  AND2_X1 U6649 ( .A1(n5080), .A2(n5066), .ZN(n7559) );
  OR2_X1 U6650 ( .A1(n4913), .A2(n7559), .ZN(n5067) );
  NAND4_X1 U6651 ( .A1(n5070), .A2(n5069), .A3(n5068), .A4(n5067), .ZN(n7824)
         );
  NAND2_X1 U6652 ( .A1(n9959), .A2(n4501), .ZN(n7726) );
  MUX2_X1 U6653 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n6281), .Z(n5088) );
  XNOR2_X1 U6654 ( .A(n5088), .B(n9025), .ZN(n5087) );
  XNOR2_X1 U6655 ( .A(n5089), .B(n5087), .ZN(n6369) );
  NAND2_X1 U6656 ( .A1(n6369), .A2(n5387), .ZN(n5076) );
  NAND2_X1 U6657 ( .A1(n5090), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5074) );
  XNOR2_X1 U6658 ( .A(n5074), .B(P2_IR_REG_12__SCAN_IN), .ZN(n9794) );
  AOI22_X1 U6659 ( .A1(n7606), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6274), .B2(
        n9794), .ZN(n5075) );
  NAND2_X1 U6660 ( .A1(n5249), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5085) );
  INV_X1 U6661 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n5077) );
  OR2_X1 U6662 ( .A1(n4971), .A2(n5077), .ZN(n5084) );
  INV_X1 U6663 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7326) );
  OR2_X1 U6664 ( .A1(n7615), .A2(n7326), .ZN(n5083) );
  NAND2_X1 U6665 ( .A1(n5080), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5081) );
  AND2_X1 U6666 ( .A1(n5096), .A2(n5081), .ZN(n7494) );
  OR2_X1 U6667 ( .A1(n4913), .A2(n7494), .ZN(n5082) );
  NAND2_X1 U6668 ( .A1(n9965), .A2(n7413), .ZN(n7725) );
  NAND2_X1 U6669 ( .A1(n7723), .A2(n7725), .ZN(n7628) );
  INV_X1 U6670 ( .A(n7628), .ZN(n5086) );
  NAND2_X1 U6671 ( .A1(n7328), .A2(n7723), .ZN(n7358) );
  MUX2_X1 U6672 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6281), .Z(n5108) );
  XNOR2_X1 U6673 ( .A(n5108), .B(SI_13_), .ZN(n5105) );
  XNOR2_X1 U6674 ( .A(n5107), .B(n5105), .ZN(n6373) );
  NAND2_X1 U6675 ( .A1(n6373), .A2(n5387), .ZN(n5093) );
  NAND2_X1 U6676 ( .A1(n5091), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5112) );
  XNOR2_X1 U6677 ( .A(n5112), .B(P2_IR_REG_13__SCAN_IN), .ZN(n9810) );
  AOI22_X1 U6678 ( .A1(n7606), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6274), .B2(
        n9810), .ZN(n5092) );
  NAND2_X1 U6679 ( .A1(n5249), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5102) );
  INV_X1 U6680 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7386) );
  OR2_X1 U6681 ( .A1(n4971), .A2(n7386), .ZN(n5101) );
  NAND2_X1 U6682 ( .A1(n5096), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5097) );
  AND2_X1 U6683 ( .A1(n5119), .A2(n5097), .ZN(n7542) );
  OR2_X1 U6684 ( .A1(n4913), .A2(n7542), .ZN(n5100) );
  INV_X1 U6685 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n5098) );
  OR2_X1 U6686 ( .A1(n7615), .A2(n5098), .ZN(n5099) );
  NAND2_X1 U6687 ( .A1(n7659), .A2(n7415), .ZN(n5103) );
  OR2_X1 U6688 ( .A1(n7659), .A2(n7415), .ZN(n5104) );
  INV_X1 U6689 ( .A(n5105), .ZN(n5106) );
  NAND2_X1 U6690 ( .A1(n5107), .A2(n5106), .ZN(n5110) );
  NAND2_X1 U6691 ( .A1(n5108), .A2(SI_13_), .ZN(n5109) );
  NAND2_X1 U6692 ( .A1(n5110), .A2(n5109), .ZN(n5127) );
  MUX2_X1 U6693 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6281), .Z(n5128) );
  XNOR2_X1 U6694 ( .A(n5128), .B(SI_14_), .ZN(n5125) );
  XNOR2_X1 U6695 ( .A(n5127), .B(n5125), .ZN(n6377) );
  NAND2_X1 U6696 ( .A1(n6377), .A2(n5387), .ZN(n5118) );
  INV_X1 U6697 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5111) );
  NAND2_X1 U6698 ( .A1(n5112), .A2(n5111), .ZN(n5113) );
  NAND2_X1 U6699 ( .A1(n5113), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5115) );
  INV_X1 U6700 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5114) );
  OR2_X1 U6701 ( .A1(n5115), .A2(n5114), .ZN(n5116) );
  NAND2_X1 U6702 ( .A1(n5115), .A2(n5114), .ZN(n5130) );
  AOI22_X1 U6703 ( .A1(n7606), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6274), .B2(
        n9825), .ZN(n5117) );
  NAND2_X1 U6704 ( .A1(n5249), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5124) );
  INV_X1 U6705 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8151) );
  OR2_X1 U6706 ( .A1(n4971), .A2(n8151), .ZN(n5123) );
  NAND2_X1 U6707 ( .A1(n5119), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5120) );
  AND2_X1 U6708 ( .A1(n5136), .A2(n5120), .ZN(n8100) );
  OR2_X1 U6709 ( .A1(n4913), .A2(n8100), .ZN(n5122) );
  INV_X1 U6710 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7903) );
  OR2_X1 U6711 ( .A1(n7615), .A2(n7903), .ZN(n5121) );
  OR2_X1 U6712 ( .A1(n8263), .A2(n8082), .ZN(n7738) );
  NAND2_X1 U6713 ( .A1(n8263), .A2(n8082), .ZN(n7737) );
  NAND2_X1 U6714 ( .A1(n7738), .A2(n7737), .ZN(n8091) );
  INV_X1 U6715 ( .A(n5125), .ZN(n5126) );
  NAND2_X1 U6716 ( .A1(n5128), .A2(SI_14_), .ZN(n5129) );
  MUX2_X1 U6717 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6281), .Z(n5145) );
  XNOR2_X1 U6718 ( .A(n5145), .B(SI_15_), .ZN(n5142) );
  XNOR2_X1 U6719 ( .A(n5144), .B(n5142), .ZN(n6427) );
  NAND2_X1 U6720 ( .A1(n6427), .A2(n5387), .ZN(n5133) );
  NAND2_X1 U6721 ( .A1(n5130), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5131) );
  XNOR2_X1 U6722 ( .A(n5131), .B(P2_IR_REG_15__SCAN_IN), .ZN(n9841) );
  AOI22_X1 U6723 ( .A1(n7606), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n9841), .B2(
        n6274), .ZN(n5132) );
  NAND2_X1 U6724 ( .A1(n5249), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5141) );
  INV_X1 U6725 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9040) );
  OR2_X1 U6726 ( .A1(n4971), .A2(n9040), .ZN(n5140) );
  INV_X1 U6727 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5134) );
  NAND2_X1 U6728 ( .A1(n5136), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5137) );
  AND2_X1 U6729 ( .A1(n5152), .A2(n5137), .ZN(n7595) );
  OR2_X1 U6730 ( .A1(n4913), .A2(n7595), .ZN(n5139) );
  INV_X1 U6731 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n9850) );
  OR2_X1 U6732 ( .A1(n7615), .A2(n9850), .ZN(n5138) );
  OR2_X1 U6733 ( .A1(n8256), .A2(n7419), .ZN(n7742) );
  INV_X1 U6734 ( .A(n5142), .ZN(n5143) );
  MUX2_X1 U6735 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n6281), .Z(n5162) );
  XNOR2_X1 U6736 ( .A(n5162), .B(SI_16_), .ZN(n5159) );
  XNOR2_X1 U6737 ( .A(n5161), .B(n5159), .ZN(n6522) );
  NAND2_X1 U6738 ( .A1(n6522), .A2(n5387), .ZN(n5151) );
  NAND2_X1 U6739 ( .A1(n5146), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5147) );
  MUX2_X1 U6740 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5147), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n5148) );
  INV_X1 U6741 ( .A(n5148), .ZN(n5149) );
  NOR2_X1 U6742 ( .A1(n5149), .A2(n5173), .ZN(n9857) );
  AOI22_X1 U6743 ( .A1(n7606), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6274), .B2(
        n9857), .ZN(n5150) );
  NAND2_X1 U6744 ( .A1(n5249), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5157) );
  INV_X1 U6745 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9050) );
  OR2_X1 U6746 ( .A1(n4971), .A2(n9050), .ZN(n5156) );
  NAND2_X1 U6747 ( .A1(n5152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5153) );
  AND2_X1 U6748 ( .A1(n5179), .A2(n5153), .ZN(n7508) );
  OR2_X1 U6749 ( .A1(n4913), .A2(n7508), .ZN(n5155) );
  INV_X1 U6750 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8073) );
  OR2_X1 U6751 ( .A1(n7615), .A2(n8073), .ZN(n5154) );
  NAND2_X1 U6752 ( .A1(n8250), .A2(n8081), .ZN(n7746) );
  INV_X1 U6753 ( .A(n7745), .ZN(n5158) );
  AOI21_X1 U6754 ( .B1(n8068), .B2(n7746), .A(n5158), .ZN(n8064) );
  INV_X1 U6755 ( .A(n5159), .ZN(n5160) );
  NAND2_X1 U6756 ( .A1(n5161), .A2(n5160), .ZN(n5164) );
  NAND2_X1 U6757 ( .A1(n5162), .A2(SI_16_), .ZN(n5163) );
  MUX2_X1 U6758 ( .A(n6586), .B(n6585), .S(n6281), .Z(n5166) );
  INV_X1 U6759 ( .A(SI_17_), .ZN(n5165) );
  NAND2_X1 U6760 ( .A1(n5166), .A2(n5165), .ZN(n5188) );
  INV_X1 U6761 ( .A(n5166), .ZN(n5167) );
  NAND2_X1 U6762 ( .A1(n5167), .A2(SI_17_), .ZN(n5168) );
  NAND2_X1 U6763 ( .A1(n5188), .A2(n5168), .ZN(n5186) );
  XNOR2_X1 U6764 ( .A(n5187), .B(n5186), .ZN(n6584) );
  NAND2_X1 U6765 ( .A1(n6584), .A2(n5387), .ZN(n5176) );
  NOR2_X1 U6766 ( .A1(n5173), .A2(n5169), .ZN(n5170) );
  MUX2_X1 U6767 ( .A(n5169), .B(n5170), .S(P2_IR_REG_17__SCAN_IN), .Z(n5171)
         );
  INV_X1 U6768 ( .A(n5171), .ZN(n5174) );
  INV_X1 U6769 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5172) );
  NAND2_X1 U6770 ( .A1(n5173), .A2(n5172), .ZN(n5210) );
  AND2_X1 U6771 ( .A1(n5174), .A2(n5210), .ZN(n9876) );
  AOI22_X1 U6772 ( .A1(n7606), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6274), .B2(
        n9876), .ZN(n5175) );
  NAND2_X1 U6773 ( .A1(n5249), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5184) );
  INV_X1 U6774 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n7863) );
  OR2_X1 U6775 ( .A1(n4971), .A2(n7863), .ZN(n5183) );
  INV_X1 U6776 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5177) );
  NAND2_X1 U6777 ( .A1(n5179), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5180) );
  AND2_X1 U6778 ( .A1(n5192), .A2(n5180), .ZN(n8061) );
  OR2_X1 U6779 ( .A1(n4913), .A2(n8061), .ZN(n5182) );
  INV_X1 U6780 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9887) );
  OR2_X1 U6781 ( .A1(n7615), .A2(n9887), .ZN(n5181) );
  OR2_X1 U6782 ( .A1(n8143), .A2(n7576), .ZN(n7751) );
  NAND2_X1 U6783 ( .A1(n8143), .A2(n7576), .ZN(n7749) );
  NAND2_X1 U6784 ( .A1(n7751), .A2(n7749), .ZN(n7744) );
  MUX2_X1 U6785 ( .A(n6676), .B(n6712), .S(n6281), .Z(n5202) );
  XNOR2_X1 U6786 ( .A(n5202), .B(SI_18_), .ZN(n5201) );
  XNOR2_X1 U6787 ( .A(n5200), .B(n5201), .ZN(n6675) );
  NAND2_X1 U6788 ( .A1(n6675), .A2(n5387), .ZN(n5191) );
  NAND2_X1 U6789 ( .A1(n5210), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5189) );
  XNOR2_X1 U6790 ( .A(n5189), .B(P2_IR_REG_18__SCAN_IN), .ZN(n9514) );
  AOI22_X1 U6791 ( .A1(n7606), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6274), .B2(
        n9514), .ZN(n5190) );
  NAND2_X1 U6792 ( .A1(n5249), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5197) );
  INV_X1 U6793 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8140) );
  OR2_X1 U6794 ( .A1(n4971), .A2(n8140), .ZN(n5196) );
  NAND2_X1 U6795 ( .A1(n5192), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5193) );
  AND2_X1 U6796 ( .A1(n5217), .A2(n5193), .ZN(n7572) );
  OR2_X1 U6797 ( .A1(n7572), .A2(n4913), .ZN(n5195) );
  INV_X1 U6798 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8053) );
  OR2_X1 U6799 ( .A1(n7615), .A2(n8053), .ZN(n5194) );
  NAND2_X1 U6800 ( .A1(n8243), .A2(n8040), .ZN(n7754) );
  NAND2_X1 U6801 ( .A1(n7752), .A2(n7754), .ZN(n8050) );
  INV_X1 U6802 ( .A(n8050), .ZN(n5198) );
  NAND2_X1 U6803 ( .A1(n5199), .A2(n7752), .ZN(n8033) );
  INV_X1 U6804 ( .A(n5202), .ZN(n5203) );
  NAND2_X1 U6805 ( .A1(n5203), .A2(SI_18_), .ZN(n5204) );
  NAND2_X1 U6806 ( .A1(n5205), .A2(n5204), .ZN(n5225) );
  MUX2_X1 U6807 ( .A(n6934), .B(n9142), .S(n6281), .Z(n5207) );
  INV_X1 U6808 ( .A(SI_19_), .ZN(n5206) );
  NAND2_X1 U6809 ( .A1(n5207), .A2(n5206), .ZN(n5226) );
  INV_X1 U6810 ( .A(n5207), .ZN(n5208) );
  NAND2_X1 U6811 ( .A1(n5208), .A2(SI_19_), .ZN(n5209) );
  NAND2_X1 U6812 ( .A1(n5226), .A2(n5209), .ZN(n5224) );
  XNOR2_X1 U6813 ( .A(n5225), .B(n5224), .ZN(n6933) );
  NAND2_X1 U6814 ( .A1(n6933), .A2(n5387), .ZN(n5214) );
  NAND2_X1 U6815 ( .A1(n5396), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5212) );
  AOI22_X1 U6816 ( .A1(n7606), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7913), .B2(
        n6274), .ZN(n5213) );
  INV_X1 U6817 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5215) );
  NAND2_X1 U6818 ( .A1(n5217), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5218) );
  NAND2_X1 U6819 ( .A1(n5235), .A2(n5218), .ZN(n8045) );
  NAND2_X1 U6820 ( .A1(n5390), .A2(n8045), .ZN(n5222) );
  INV_X1 U6821 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8236) );
  OR2_X1 U6822 ( .A1(n4908), .A2(n8236), .ZN(n5221) );
  INV_X1 U6823 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8137) );
  OR2_X1 U6824 ( .A1(n4971), .A2(n8137), .ZN(n5220) );
  INV_X1 U6825 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8044) );
  OR2_X1 U6826 ( .A1(n7615), .A2(n8044), .ZN(n5219) );
  NAND2_X1 U6827 ( .A1(n8237), .A2(n7532), .ZN(n7757) );
  INV_X1 U6828 ( .A(n5223), .ZN(n7657) );
  MUX2_X1 U6829 ( .A(n7076), .B(n7069), .S(n6281), .Z(n5228) );
  INV_X1 U6830 ( .A(SI_20_), .ZN(n5227) );
  NAND2_X1 U6831 ( .A1(n5228), .A2(n5227), .ZN(n5242) );
  INV_X1 U6832 ( .A(n5228), .ZN(n5229) );
  NAND2_X1 U6833 ( .A1(n5229), .A2(SI_20_), .ZN(n5230) );
  XNOR2_X1 U6834 ( .A(n5241), .B(n5240), .ZN(n7068) );
  NAND2_X1 U6835 ( .A1(n7068), .A2(n5387), .ZN(n5232) );
  OR2_X1 U6836 ( .A1(n7609), .A2(n7076), .ZN(n5231) );
  NAND2_X1 U6837 ( .A1(n4261), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5234) );
  NAND2_X1 U6838 ( .A1(n5249), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5233) );
  AND2_X1 U6839 ( .A1(n5234), .A2(n5233), .ZN(n5239) );
  NAND2_X1 U6840 ( .A1(n5235), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5236) );
  NAND2_X1 U6841 ( .A1(n5247), .A2(n5236), .ZN(n8029) );
  NAND2_X1 U6842 ( .A1(n8029), .A2(n5390), .ZN(n5238) );
  NAND2_X1 U6843 ( .A1(n5408), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5237) );
  NAND2_X1 U6844 ( .A1(n8021), .A2(n7758), .ZN(n8007) );
  MUX2_X1 U6845 ( .A(n7080), .B(n7079), .S(n6281), .Z(n5254) );
  XNOR2_X1 U6846 ( .A(n5254), .B(SI_21_), .ZN(n5253) );
  XNOR2_X1 U6847 ( .A(n5258), .B(n5253), .ZN(n7078) );
  NAND2_X1 U6848 ( .A1(n7078), .A2(n5387), .ZN(n5244) );
  OR2_X1 U6849 ( .A1(n7609), .A2(n7080), .ZN(n5243) );
  INV_X1 U6850 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5245) );
  NAND2_X1 U6851 ( .A1(n5247), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5248) );
  NAND2_X1 U6852 ( .A1(n5265), .A2(n5248), .ZN(n8018) );
  NAND2_X1 U6853 ( .A1(n8018), .A2(n5390), .ZN(n5252) );
  AOI22_X1 U6854 ( .A1(n5249), .A2(P2_REG0_REG_21__SCAN_IN), .B1(n4262), .B2(
        P2_REG1_REG_21__SCAN_IN), .ZN(n5251) );
  NAND2_X1 U6855 ( .A1(n5408), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5250) );
  NAND2_X1 U6856 ( .A1(n8225), .A2(n7430), .ZN(n7760) );
  NAND2_X1 U6857 ( .A1(n8231), .A2(n8041), .ZN(n8006) );
  AND2_X1 U6858 ( .A1(n7760), .A2(n8006), .ZN(n7755) );
  INV_X1 U6859 ( .A(n5253), .ZN(n5257) );
  INV_X1 U6860 ( .A(n5254), .ZN(n5255) );
  NAND2_X1 U6861 ( .A1(n5255), .A2(SI_21_), .ZN(n5256) );
  INV_X1 U6862 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7391) );
  MUX2_X1 U6863 ( .A(n9092), .B(n7391), .S(n6281), .Z(n5260) );
  INV_X1 U6864 ( .A(SI_22_), .ZN(n5259) );
  NAND2_X1 U6865 ( .A1(n5260), .A2(n5259), .ZN(n5272) );
  INV_X1 U6866 ( .A(n5260), .ZN(n5261) );
  NAND2_X1 U6867 ( .A1(n5261), .A2(SI_22_), .ZN(n5262) );
  NAND2_X1 U6868 ( .A1(n5272), .A2(n5262), .ZN(n5273) );
  XNOR2_X1 U6869 ( .A(n5274), .B(n5273), .ZN(n7178) );
  NAND2_X1 U6870 ( .A1(n7178), .A2(n5387), .ZN(n5264) );
  OR2_X1 U6871 ( .A1(n7609), .A2(n9092), .ZN(n5263) );
  NAND2_X1 U6872 ( .A1(n5265), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5266) );
  NAND2_X1 U6873 ( .A1(n5285), .A2(n5266), .ZN(n7996) );
  NAND2_X1 U6874 ( .A1(n7996), .A2(n5390), .ZN(n5269) );
  AOI22_X1 U6875 ( .A1(n5249), .A2(P2_REG0_REG_22__SCAN_IN), .B1(n4261), .B2(
        P2_REG1_REG_22__SCAN_IN), .ZN(n5268) );
  NAND2_X1 U6876 ( .A1(n5408), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5267) );
  NOR2_X1 U6877 ( .A1(n8219), .A2(n7987), .ZN(n5270) );
  NAND2_X1 U6878 ( .A1(n8219), .A2(n7987), .ZN(n5271) );
  INV_X1 U6879 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5275) );
  MUX2_X1 U6880 ( .A(n7224), .B(n5275), .S(n6281), .Z(n5277) );
  INV_X1 U6881 ( .A(SI_23_), .ZN(n5276) );
  NAND2_X1 U6882 ( .A1(n5277), .A2(n5276), .ZN(n5293) );
  INV_X1 U6883 ( .A(n5277), .ZN(n5278) );
  NAND2_X1 U6884 ( .A1(n5278), .A2(SI_23_), .ZN(n5279) );
  NAND2_X1 U6885 ( .A1(n5281), .A2(n5280), .ZN(n5294) );
  OR2_X1 U6886 ( .A1(n5281), .A2(n5280), .ZN(n5282) );
  NAND2_X1 U6887 ( .A1(n7221), .A2(n5387), .ZN(n5284) );
  OR2_X1 U6888 ( .A1(n7609), .A2(n7224), .ZN(n5283) );
  NAND2_X1 U6889 ( .A1(n5285), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5286) );
  NAND2_X1 U6890 ( .A1(n5303), .A2(n5286), .ZN(n7990) );
  NAND2_X1 U6891 ( .A1(n7990), .A2(n5390), .ZN(n5291) );
  INV_X1 U6892 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n7989) );
  NAND2_X1 U6893 ( .A1(n5249), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5288) );
  NAND2_X1 U6894 ( .A1(n4262), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5287) );
  OAI211_X1 U6895 ( .C1(n7989), .C2(n7615), .A(n5288), .B(n5287), .ZN(n5289)
         );
  INV_X1 U6896 ( .A(n5289), .ZN(n5290) );
  NAND2_X1 U6897 ( .A1(n7982), .A2(n7768), .ZN(n5292) );
  NAND2_X1 U6898 ( .A1(n7991), .A2(n7550), .ZN(n7770) );
  NAND2_X1 U6899 ( .A1(n5292), .A2(n7770), .ZN(n7972) );
  INV_X1 U6900 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7399) );
  INV_X1 U6901 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7239) );
  MUX2_X1 U6902 ( .A(n7399), .B(n7239), .S(n6281), .Z(n5296) );
  INV_X1 U6903 ( .A(SI_24_), .ZN(n5295) );
  NAND2_X1 U6904 ( .A1(n5296), .A2(n5295), .ZN(n5312) );
  INV_X1 U6905 ( .A(n5296), .ZN(n5297) );
  NAND2_X1 U6906 ( .A1(n5297), .A2(SI_24_), .ZN(n5298) );
  XNOR2_X1 U6907 ( .A(n5311), .B(n5310), .ZN(n7238) );
  NAND2_X1 U6908 ( .A1(n7238), .A2(n5387), .ZN(n5300) );
  OR2_X1 U6909 ( .A1(n7609), .A2(n7399), .ZN(n5299) );
  INV_X1 U6910 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5301) );
  NAND2_X1 U6911 ( .A1(n5303), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5304) );
  NAND2_X1 U6912 ( .A1(n5322), .A2(n5304), .ZN(n7979) );
  NAND2_X1 U6913 ( .A1(n7979), .A2(n5390), .ZN(n5309) );
  INV_X1 U6914 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8206) );
  NAND2_X1 U6915 ( .A1(n5408), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5306) );
  NAND2_X1 U6916 ( .A1(n4261), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5305) );
  OAI211_X1 U6917 ( .C1(n4908), .C2(n8206), .A(n5306), .B(n5305), .ZN(n5307)
         );
  INV_X1 U6918 ( .A(n5307), .ZN(n5308) );
  OAI21_X2 U6919 ( .B1(n7972), .B2(n7626), .A(n7773), .ZN(n7967) );
  NAND2_X1 U6920 ( .A1(n5311), .A2(n5310), .ZN(n5313) );
  INV_X1 U6921 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7309) );
  MUX2_X1 U6922 ( .A(n9053), .B(n7309), .S(n6281), .Z(n5315) );
  INV_X1 U6923 ( .A(SI_25_), .ZN(n5314) );
  NAND2_X1 U6924 ( .A1(n5315), .A2(n5314), .ZN(n5332) );
  INV_X1 U6925 ( .A(n5315), .ZN(n5316) );
  NAND2_X1 U6926 ( .A1(n5316), .A2(SI_25_), .ZN(n5317) );
  NAND2_X1 U6927 ( .A1(n7308), .A2(n5387), .ZN(n5319) );
  OR2_X1 U6928 ( .A1(n7609), .A2(n9053), .ZN(n5318) );
  INV_X1 U6929 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5320) );
  NAND2_X1 U6930 ( .A1(n5322), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5323) );
  NAND2_X1 U6931 ( .A1(n5339), .A2(n5323), .ZN(n7966) );
  NAND2_X1 U6932 ( .A1(n7966), .A2(n5390), .ZN(n5328) );
  INV_X1 U6933 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9039) );
  NAND2_X1 U6934 ( .A1(n5249), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5325) );
  NAND2_X1 U6935 ( .A1(n5408), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5324) );
  OAI211_X1 U6936 ( .C1(n4971), .C2(n9039), .A(n5325), .B(n5324), .ZN(n5326)
         );
  INV_X1 U6937 ( .A(n5326), .ZN(n5327) );
  NAND2_X1 U6938 ( .A1(n8201), .A2(n7949), .ZN(n7777) );
  NAND2_X1 U6939 ( .A1(n7967), .A2(n7777), .ZN(n5329) );
  INV_X1 U6940 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7319) );
  INV_X1 U6941 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7312) );
  MUX2_X1 U6942 ( .A(n7319), .B(n7312), .S(n6281), .Z(n5334) );
  INV_X1 U6943 ( .A(SI_26_), .ZN(n5333) );
  NAND2_X1 U6944 ( .A1(n5334), .A2(n5333), .ZN(n5349) );
  INV_X1 U6945 ( .A(n5334), .ZN(n5335) );
  NAND2_X1 U6946 ( .A1(n5335), .A2(SI_26_), .ZN(n5336) );
  NAND2_X1 U6947 ( .A1(n7311), .A2(n5387), .ZN(n5338) );
  OR2_X1 U6948 ( .A1(n7609), .A2(n7319), .ZN(n5337) );
  NAND2_X1 U6949 ( .A1(n5339), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5340) );
  NAND2_X1 U6950 ( .A1(n5359), .A2(n5340), .ZN(n7953) );
  NAND2_X1 U6951 ( .A1(n7953), .A2(n5390), .ZN(n5345) );
  INV_X1 U6952 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8197) );
  NAND2_X1 U6953 ( .A1(n4262), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5342) );
  NAND2_X1 U6954 ( .A1(n5408), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5341) );
  OAI211_X1 U6955 ( .C1(n8197), .C2(n4908), .A(n5342), .B(n5341), .ZN(n5343)
         );
  INV_X1 U6956 ( .A(n5343), .ZN(n5344) );
  NOR2_X1 U6957 ( .A1(n7952), .A2(n7938), .ZN(n5346) );
  INV_X1 U6958 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5354) );
  INV_X1 U6959 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7395) );
  MUX2_X1 U6960 ( .A(n5354), .B(n7395), .S(n6281), .Z(n5351) );
  INV_X1 U6961 ( .A(SI_27_), .ZN(n5350) );
  NAND2_X1 U6962 ( .A1(n5351), .A2(n5350), .ZN(n5368) );
  INV_X1 U6963 ( .A(n5351), .ZN(n5352) );
  NAND2_X1 U6964 ( .A1(n5352), .A2(SI_27_), .ZN(n5353) );
  NAND2_X1 U6965 ( .A1(n6104), .A2(n5387), .ZN(n5356) );
  OR2_X1 U6966 ( .A1(n7609), .A2(n5354), .ZN(n5355) );
  INV_X1 U6967 ( .A(n5359), .ZN(n5358) );
  INV_X1 U6968 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5357) );
  NAND2_X1 U6969 ( .A1(n5359), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5360) );
  NAND2_X1 U6970 ( .A1(n5373), .A2(n5360), .ZN(n7939) );
  NAND2_X1 U6971 ( .A1(n7939), .A2(n5390), .ZN(n5365) );
  INV_X1 U6972 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9048) );
  NAND2_X1 U6973 ( .A1(n5408), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5362) );
  NAND2_X1 U6974 ( .A1(n4261), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5361) );
  OAI211_X1 U6975 ( .C1(n4908), .C2(n9048), .A(n5362), .B(n5361), .ZN(n5363)
         );
  INV_X1 U6976 ( .A(n5363), .ZN(n5364) );
  NAND2_X1 U6977 ( .A1(n7940), .A2(n7948), .ZN(n7784) );
  INV_X1 U6978 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7357) );
  INV_X1 U6979 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n5370) );
  MUX2_X1 U6980 ( .A(n7357), .B(n5370), .S(n6281), .Z(n5383) );
  XNOR2_X1 U6981 ( .A(n5383), .B(SI_28_), .ZN(n5380) );
  NAND2_X1 U6982 ( .A1(n7354), .A2(n5387), .ZN(n5372) );
  OR2_X1 U6983 ( .A1(n7609), .A2(n7357), .ZN(n5371) );
  NAND2_X1 U6984 ( .A1(n5373), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5374) );
  NAND2_X1 U6985 ( .A1(n5494), .A2(n5374), .ZN(n7931) );
  NAND2_X1 U6986 ( .A1(n7931), .A2(n5390), .ZN(n5379) );
  INV_X1 U6987 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8188) );
  NAND2_X1 U6988 ( .A1(n4261), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5376) );
  NAND2_X1 U6989 ( .A1(n5408), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5375) );
  OAI211_X1 U6990 ( .C1(n4908), .C2(n8188), .A(n5376), .B(n5375), .ZN(n5377)
         );
  INV_X1 U6991 ( .A(n5377), .ZN(n5378) );
  OAI22_X1 U6992 ( .A1(n7930), .A2(n7929), .B1(n7937), .B2(n7797), .ZN(n7624)
         );
  INV_X1 U6993 ( .A(SI_28_), .ZN(n5382) );
  NAND2_X1 U6994 ( .A1(n5383), .A2(n5382), .ZN(n5384) );
  INV_X1 U6995 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9077) );
  INV_X1 U6996 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n5386) );
  MUX2_X1 U6997 ( .A(n9077), .B(n5386), .S(n6281), .Z(n6215) );
  NAND2_X1 U6998 ( .A1(n8275), .A2(n5387), .ZN(n5389) );
  OR2_X1 U6999 ( .A1(n7609), .A2(n9077), .ZN(n5388) );
  INV_X1 U7000 ( .A(n5494), .ZN(n5391) );
  NAND2_X1 U7001 ( .A1(n5391), .A2(n5390), .ZN(n7621) );
  INV_X1 U7002 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n5515) );
  NAND2_X1 U7003 ( .A1(n4262), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5393) );
  NAND2_X1 U7004 ( .A1(n5408), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5392) );
  OAI211_X1 U7005 ( .C1(n4908), .C2(n5515), .A(n5393), .B(n5392), .ZN(n5394)
         );
  INV_X1 U7006 ( .A(n5394), .ZN(n5395) );
  NAND2_X1 U7007 ( .A1(n7654), .A2(n7655), .ZN(n7613) );
  NAND2_X1 U7008 ( .A1(n7804), .A2(n7888), .ZN(n6645) );
  INV_X1 U7009 ( .A(n5402), .ZN(n5403) );
  NAND2_X1 U7010 ( .A1(n5403), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5404) );
  MUX2_X1 U7011 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5404), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n5405) );
  OR2_X1 U7012 ( .A1(n6645), .A2(n7781), .ZN(n6466) );
  INV_X1 U7013 ( .A(n7804), .ZN(n5489) );
  NAND2_X1 U7014 ( .A1(n7888), .A2(n9948), .ZN(n5406) );
  AOI21_X1 U7015 ( .B1(n5489), .B2(n7663), .A(n5406), .ZN(n5407) );
  NAND2_X1 U7016 ( .A1(n6466), .A2(n5407), .ZN(n7155) );
  INV_X1 U7017 ( .A(n7811), .ZN(n6362) );
  INV_X1 U7018 ( .A(n7924), .ZN(n6669) );
  INV_X1 U7019 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8186) );
  NAND2_X1 U7020 ( .A1(n5408), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5410) );
  NAND2_X1 U7021 ( .A1(n4262), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5409) );
  OAI211_X1 U7022 ( .C1(n4908), .C2(n8186), .A(n5410), .B(n5409), .ZN(n5411)
         );
  INV_X1 U7023 ( .A(n5411), .ZN(n5412) );
  NAND2_X1 U7024 ( .A1(n7621), .A2(n5412), .ZN(n7819) );
  AOI21_X1 U7025 ( .B1(P2_B_REG_SCAN_IN), .B2(n4864), .A(n8080), .ZN(n7916) );
  AOI22_X1 U7026 ( .A1(n8092), .A2(n7820), .B1(n7819), .B2(n7916), .ZN(n5457)
         );
  INV_X1 U7027 ( .A(n6721), .ZN(n7834) );
  NAND2_X1 U7028 ( .A1(n7834), .A2(n6470), .ZN(n6619) );
  NAND2_X1 U7029 ( .A1(n8165), .A2(n6722), .ZN(n5414) );
  INV_X1 U7030 ( .A(n8171), .ZN(n5415) );
  OR2_X1 U7031 ( .A1(n7832), .A2(n5415), .ZN(n5416) );
  NOR2_X1 U7032 ( .A1(n8162), .A2(n7063), .ZN(n7084) );
  INV_X1 U7033 ( .A(n7678), .ZN(n5417) );
  NAND2_X1 U7034 ( .A1(n8162), .A2(n7063), .ZN(n7086) );
  AND2_X1 U7035 ( .A1(n5417), .A2(n7086), .ZN(n5418) );
  NAND2_X1 U7036 ( .A1(n7144), .A2(n9918), .ZN(n5419) );
  NAND2_X1 U7037 ( .A1(n7830), .A2(n7039), .ZN(n5420) );
  NAND2_X1 U7038 ( .A1(n7142), .A2(n5420), .ZN(n5422) );
  NAND2_X1 U7039 ( .A1(n7105), .A2(n9921), .ZN(n5421) );
  NAND2_X1 U7040 ( .A1(n7151), .A2(n5423), .ZN(n7150) );
  NAND2_X1 U7041 ( .A1(n7282), .A2(n9932), .ZN(n5424) );
  NAND2_X1 U7042 ( .A1(n7827), .A2(n7294), .ZN(n5425) );
  NAND2_X1 U7043 ( .A1(n7212), .A2(n5425), .ZN(n5427) );
  NAND2_X1 U7044 ( .A1(n7339), .A2(n9937), .ZN(n5426) );
  NAND2_X1 U7045 ( .A1(n5427), .A2(n5426), .ZN(n7298) );
  NAND2_X1 U7046 ( .A1(n9942), .A2(n7378), .ZN(n5428) );
  NAND2_X1 U7047 ( .A1(n9947), .A2(n7825), .ZN(n5429) );
  NAND2_X1 U7048 ( .A1(n5430), .A2(n5429), .ZN(n7314) );
  NAND2_X1 U7049 ( .A1(n9959), .A2(n7824), .ZN(n5432) );
  AND2_X1 U7050 ( .A1(n9965), .A2(n7823), .ZN(n5434) );
  NOR2_X1 U7051 ( .A1(n7659), .A2(n8093), .ZN(n7660) );
  NAND2_X1 U7052 ( .A1(n7659), .A2(n8093), .ZN(n7734) );
  OR2_X1 U7053 ( .A1(n8263), .A2(n7822), .ZN(n5435) );
  NOR2_X1 U7054 ( .A1(n8256), .A2(n8094), .ZN(n5436) );
  INV_X1 U7055 ( .A(n8256), .ZN(n7604) );
  OAI22_X1 U7056 ( .A1(n8079), .A2(n5436), .B1(n7419), .B2(n7604), .ZN(n8070)
         );
  NAND2_X1 U7057 ( .A1(n7745), .A2(n7746), .ZN(n7741) );
  NAND2_X1 U7058 ( .A1(n8070), .A2(n7741), .ZN(n5438) );
  NAND2_X1 U7059 ( .A1(n8250), .A2(n8058), .ZN(n5437) );
  NAND2_X1 U7060 ( .A1(n5438), .A2(n5437), .ZN(n8057) );
  INV_X1 U7061 ( .A(n7576), .ZN(n8071) );
  NAND2_X1 U7062 ( .A1(n8143), .A2(n8071), .ZN(n5439) );
  INV_X1 U7063 ( .A(n8032), .ZN(n8035) );
  OR2_X1 U7064 ( .A1(n8243), .A2(n8059), .ZN(n8036) );
  AND2_X1 U7065 ( .A1(n8035), .A2(n8036), .ZN(n5441) );
  NAND2_X1 U7066 ( .A1(n7758), .A2(n8006), .ZN(n8024) );
  NAND2_X1 U7067 ( .A1(n8237), .A2(n8051), .ZN(n8022) );
  AND2_X1 U7068 ( .A1(n8024), .A2(n8022), .ZN(n5442) );
  OR2_X1 U7069 ( .A1(n8231), .A2(n8015), .ZN(n8010) );
  NAND2_X1 U7070 ( .A1(n8023), .A2(n8010), .ZN(n5443) );
  NAND2_X1 U7071 ( .A1(n7759), .A2(n7760), .ZN(n8009) );
  NAND2_X1 U7072 ( .A1(n5443), .A2(n8009), .ZN(n8013) );
  OR2_X1 U7073 ( .A1(n8225), .A2(n8026), .ZN(n5444) );
  NAND2_X1 U7074 ( .A1(n8013), .A2(n5444), .ZN(n7998) );
  XNOR2_X1 U7075 ( .A(n8219), .B(n7987), .ZN(n7999) );
  NAND2_X1 U7076 ( .A1(n7998), .A2(n7999), .ZN(n7997) );
  OR2_X1 U7077 ( .A1(n8219), .A2(n8014), .ZN(n7765) );
  NAND2_X1 U7078 ( .A1(n7997), .A2(n7765), .ZN(n7984) );
  NAND2_X1 U7079 ( .A1(n7991), .A2(n8000), .ZN(n5445) );
  INV_X1 U7080 ( .A(n7991), .ZN(n8213) );
  NAND2_X1 U7081 ( .A1(n8213), .A2(n7550), .ZN(n5446) );
  NAND2_X1 U7082 ( .A1(n8207), .A2(n7961), .ZN(n5447) );
  AND2_X1 U7083 ( .A1(n8201), .A2(n7975), .ZN(n5450) );
  OR2_X1 U7084 ( .A1(n8201), .A2(n7975), .ZN(n5449) );
  OAI21_X2 U7085 ( .B1(n7960), .B2(n5450), .A(n5449), .ZN(n7946) );
  NOR2_X1 U7086 ( .A1(n7952), .A2(n7962), .ZN(n5452) );
  NAND2_X1 U7087 ( .A1(n7952), .A2(n7962), .ZN(n5451) );
  AND2_X1 U7088 ( .A1(n7940), .A2(n7821), .ZN(n5453) );
  INV_X1 U7089 ( .A(n7650), .ZN(n5454) );
  NAND2_X1 U7090 ( .A1(n5489), .A2(n6643), .ZN(n7605) );
  NAND2_X1 U7091 ( .A1(n7913), .A2(n7814), .ZN(n5507) );
  NAND2_X1 U7092 ( .A1(n5455), .A2(n8167), .ZN(n5456) );
  OAI211_X1 U7093 ( .C1(n5502), .C2(n7155), .A(n5457), .B(n5456), .ZN(n5504)
         );
  NAND2_X1 U7094 ( .A1(n5487), .A2(n5486), .ZN(n5458) );
  INV_X1 U7095 ( .A(n5461), .ZN(n5462) );
  NAND2_X1 U7096 ( .A1(n5462), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n5464) );
  XNOR2_X1 U7097 ( .A(n7401), .B(P2_B_REG_SCAN_IN), .ZN(n5465) );
  NAND2_X1 U7098 ( .A1(n7393), .A2(n5465), .ZN(n5470) );
  NAND2_X1 U7099 ( .A1(n4319), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5466) );
  MUX2_X1 U7100 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5466), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5468) );
  NAND2_X1 U7101 ( .A1(n5468), .A2(n5467), .ZN(n7321) );
  INV_X1 U7102 ( .A(n7321), .ZN(n5469) );
  NAND2_X1 U7103 ( .A1(n7401), .A2(n7321), .ZN(n6348) );
  NAND2_X1 U7104 ( .A1(n7393), .A2(n7321), .ZN(n5471) );
  NOR2_X1 U7105 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .ZN(
        n5476) );
  NOR4_X1 U7106 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n5475) );
  NOR4_X1 U7107 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n5474) );
  NOR4_X1 U7108 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_31__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n5473) );
  NAND4_X1 U7109 ( .A1(n5476), .A2(n5475), .A3(n5474), .A4(n5473), .ZN(n5482)
         );
  NOR4_X1 U7110 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n5480) );
  NOR4_X1 U7111 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n5479) );
  NOR4_X1 U7112 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5478) );
  NOR4_X1 U7113 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n5477) );
  NAND4_X1 U7114 ( .A1(n5480), .A2(n5479), .A3(n5478), .A4(n5477), .ZN(n5481)
         );
  NOR2_X1 U7115 ( .A1(n5482), .A2(n5481), .ZN(n5483) );
  INV_X1 U7116 ( .A(n7393), .ZN(n5485) );
  NOR2_X1 U7117 ( .A1(n7401), .A2(n7321), .ZN(n5484) );
  NAND2_X1 U7118 ( .A1(n6645), .A2(n7801), .ZN(n6629) );
  AND3_X1 U7119 ( .A1(n5511), .A2(n6637), .A3(n6629), .ZN(n5488) );
  NAND3_X1 U7120 ( .A1(n5489), .A2(n7814), .A3(n7888), .ZN(n5490) );
  INV_X1 U7121 ( .A(n6200), .ZN(n6202) );
  NAND2_X1 U7122 ( .A1(n6642), .A2(n6202), .ZN(n5492) );
  NAND2_X1 U7123 ( .A1(n6322), .A2(n6200), .ZN(n5491) );
  NAND2_X1 U7124 ( .A1(n5504), .A2(n8098), .ZN(n5500) );
  AND2_X1 U7125 ( .A1(n9897), .A2(n6643), .ZN(n9903) );
  NAND2_X1 U7126 ( .A1(n8098), .A2(n9903), .ZN(n7306) );
  NOR2_X1 U7127 ( .A1(n5494), .A2(n9896), .ZN(n7918) );
  NOR2_X1 U7128 ( .A1(n6208), .A2(n7955), .ZN(n5496) );
  AOI211_X1 U7129 ( .C1(n9907), .C2(P2_REG2_REG_29__SCAN_IN), .A(n7918), .B(
        n5496), .ZN(n5497) );
  NAND2_X1 U7130 ( .A1(n5500), .A2(n5499), .ZN(P2_U3204) );
  INV_X1 U7131 ( .A(n9953), .ZN(n5501) );
  INV_X1 U7132 ( .A(n5511), .ZN(n5505) );
  NOR2_X1 U7133 ( .A1(n5506), .A2(n5505), .ZN(n6635) );
  NAND2_X1 U7134 ( .A1(n6635), .A2(n6637), .ZN(n6665) );
  INV_X1 U7135 ( .A(n7652), .ZN(n5509) );
  INV_X1 U7136 ( .A(n5507), .ZN(n5508) );
  NAND2_X1 U7137 ( .A1(n5509), .A2(n5508), .ZN(n6628) );
  AND2_X1 U7138 ( .A1(n6628), .A2(n6466), .ZN(n5510) );
  NAND3_X1 U7139 ( .A1(n6642), .A2(n6322), .A3(n5511), .ZN(n6639) );
  INV_X1 U7140 ( .A(n6637), .ZN(n6321) );
  NOR2_X1 U7141 ( .A1(n7801), .A2(n9966), .ZN(n5512) );
  NAND2_X1 U7142 ( .A1(n6628), .A2(n5512), .ZN(n6659) );
  NAND2_X1 U7143 ( .A1(n6659), .A2(n8096), .ZN(n6627) );
  NAND2_X1 U7144 ( .A1(n6668), .A2(n6627), .ZN(n5513) );
  OR2_X1 U7145 ( .A1(n9967), .A2(n5515), .ZN(n5516) );
  OAI21_X1 U7146 ( .B1(n6212), .B2(n9969), .A(n5518), .ZN(P2_U3456) );
  INV_X2 U7147 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X2 U7148 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5620) );
  NOR2_X1 U7149 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5519) );
  AND2_X2 U7150 ( .A1(n5620), .A2(n5519), .ZN(n5822) );
  NOR2_X2 U7151 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5521) );
  INV_X1 U7152 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5520) );
  AND4_X2 U7153 ( .A1(n5521), .A2(n5842), .A3(n5865), .A4(n5520), .ZN(n5525)
         );
  AND3_X2 U7154 ( .A1(n5819), .A2(n5818), .A3(n5817), .ZN(n5524) );
  NOR2_X1 U7155 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5523) );
  NOR2_X1 U7156 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5529) );
  NOR2_X1 U7157 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5528) );
  NOR2_X1 U7158 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5527) );
  INV_X1 U7159 ( .A(n5576), .ZN(n5532) );
  NOR2_X1 U7160 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(n5532), .ZN(n5533) );
  NAND2_X1 U7161 ( .A1(n8552), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5544) );
  NAND2_X1 U7162 ( .A1(n5657), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5543) );
  AND2_X2 U7163 ( .A1(n9494), .A2(n5538), .ZN(n5634) );
  NAND2_X1 U7164 ( .A1(n5634), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5541) );
  NAND2_X1 U7165 ( .A1(n5635), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5540) );
  NAND2_X1 U7166 ( .A1(n5577), .A2(n5545), .ZN(n5549) );
  NAND2_X1 U7167 ( .A1(n5556), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5548) );
  MUX2_X1 U7168 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5548), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n5550) );
  INV_X1 U7169 ( .A(n7310), .ZN(n5551) );
  NAND3_X1 U7170 ( .A1(n5917), .A2(n5569), .A3(n5570), .ZN(n5552) );
  NAND2_X1 U7171 ( .A1(n4258), .A2(n4824), .ZN(n5564) );
  INV_X1 U7172 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5553) );
  NAND2_X1 U7173 ( .A1(n5565), .A2(n5553), .ZN(n5554) );
  NAND2_X1 U7174 ( .A1(n6165), .A2(n6168), .ZN(n5555) );
  INV_X2 U7175 ( .A(n5556), .ZN(n5577) );
  INV_X1 U7176 ( .A(n7240), .ZN(n5560) );
  NAND2_X1 U7177 ( .A1(n5561), .A2(n5565), .ZN(n5562) );
  NAND2_X1 U7178 ( .A1(n5564), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5566) );
  AND2_X2 U7179 ( .A1(n6191), .A2(n8712), .ZN(n5590) );
  OAI21_X2 U7180 ( .B1(n5567), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5916) );
  NAND2_X1 U7181 ( .A1(n5916), .A2(n5917), .ZN(n5568) );
  NAND2_X1 U7182 ( .A1(n5938), .A2(n5569), .ZN(n5940) );
  NAND2_X1 U7183 ( .A1(n5571), .A2(n5570), .ZN(n5572) );
  INV_X1 U7184 ( .A(n4263), .ZN(n6342) );
  NAND2_X1 U7185 ( .A1(n5589), .A2(n4260), .ZN(n5597) );
  INV_X1 U7186 ( .A(n5575), .ZN(n6299) );
  NAND2_X1 U7187 ( .A1(n5577), .A2(n5576), .ZN(n5578) );
  NAND2_X1 U7188 ( .A1(n5582), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5583) );
  NAND2_X1 U7189 ( .A1(n5602), .A2(n6281), .ZN(n5640) );
  INV_X2 U7190 ( .A(n5602), .ZN(n5619) );
  NAND2_X1 U7191 ( .A1(n5619), .A2(n8739), .ZN(n5585) );
  NAND2_X1 U7192 ( .A1(n5597), .A2(n6414), .ZN(n5587) );
  INV_X1 U7193 ( .A(n5595), .ZN(n5593) );
  INV_X2 U7194 ( .A(n4253), .ZN(n6021) );
  AND2_X1 U7195 ( .A1(n6414), .A2(n5590), .ZN(n5591) );
  INV_X1 U7196 ( .A(n5594), .ZN(n5592) );
  NAND2_X1 U7197 ( .A1(n5595), .A2(n5594), .ZN(n5614) );
  INV_X1 U7199 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n8754) );
  NAND2_X1 U7200 ( .A1(n6281), .A2(SI_0_), .ZN(n5599) );
  INV_X1 U7201 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5598) );
  NAND2_X1 U7202 ( .A1(n5599), .A2(n5598), .ZN(n5601) );
  AND2_X1 U7203 ( .A1(n5601), .A2(n5600), .ZN(n9502) );
  NAND2_X1 U7204 ( .A1(n5634), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5605) );
  NAND2_X1 U7205 ( .A1(n5635), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5604) );
  NAND2_X1 U7206 ( .A1(n5657), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5603) );
  AND3_X1 U7207 ( .A1(n5605), .A2(n5604), .A3(n5603), .ZN(n5607) );
  NAND2_X2 U7208 ( .A1(n5607), .A2(n5606), .ZN(n6762) );
  AOI22_X2 U7209 ( .A1(n5648), .A2(n6782), .B1(n6762), .B2(n5590), .ZN(n5612)
         );
  INV_X1 U7210 ( .A(n6191), .ZN(n6272) );
  NAND2_X1 U7211 ( .A1(n6272), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5608) );
  NAND2_X1 U7212 ( .A1(n5612), .A2(n5608), .ZN(n6351) );
  NAND2_X1 U7213 ( .A1(n6762), .A2(n6145), .ZN(n5610) );
  AOI22_X1 U7214 ( .A1(n6782), .A2(n5590), .B1(n6272), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n5609) );
  NAND2_X1 U7215 ( .A1(n5610), .A2(n5609), .ZN(n6352) );
  NAND2_X1 U7216 ( .A1(n5612), .A2(n4266), .ZN(n5613) );
  NAND2_X1 U7217 ( .A1(n6411), .A2(n5614), .ZN(n8403) );
  NAND2_X1 U7218 ( .A1(n4265), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5618) );
  NAND2_X1 U7219 ( .A1(n5657), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5617) );
  NAND2_X1 U7220 ( .A1(n5634), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5616) );
  NAND2_X1 U7221 ( .A1(n5635), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5615) );
  NAND4_X2 U7222 ( .A1(n5618), .A2(n5615), .A3(n5616), .A4(n5617), .ZN(n8735)
         );
  NAND2_X1 U7223 ( .A1(n8735), .A2(n5590), .ZN(n5624) );
  OR2_X1 U7224 ( .A1(n5620), .A2(n9490), .ZN(n5643) );
  XNOR2_X1 U7225 ( .A(n5643), .B(P1_IR_REG_2__SCAN_IN), .ZN(n8760) );
  NAND2_X1 U7226 ( .A1(n5619), .A2(n8760), .ZN(n5621) );
  OAI211_X1 U7227 ( .C1(n6285), .C2(n5640), .A(n5622), .B(n5621), .ZN(n8406)
         );
  NAND2_X1 U7228 ( .A1(n5624), .A2(n5623), .ZN(n5625) );
  XNOR2_X1 U7229 ( .A(n5625), .B(n5611), .ZN(n5630) );
  INV_X1 U7230 ( .A(n5630), .ZN(n5628) );
  AND2_X1 U7231 ( .A1(n8406), .A2(n5590), .ZN(n5626) );
  AOI21_X1 U7232 ( .B1(n8735), .B2(n6145), .A(n5626), .ZN(n5629) );
  INV_X1 U7233 ( .A(n5629), .ZN(n5627) );
  NAND2_X1 U7234 ( .A1(n5628), .A2(n5627), .ZN(n5631) );
  NAND2_X1 U7235 ( .A1(n5630), .A2(n5629), .ZN(n5632) );
  AND2_X1 U7236 ( .A1(n5631), .A2(n5632), .ZN(n8404) );
  NAND2_X1 U7237 ( .A1(n4265), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5639) );
  INV_X1 U7238 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5633) );
  NAND2_X1 U7239 ( .A1(n6134), .A2(n5633), .ZN(n5638) );
  NAND2_X1 U7240 ( .A1(n5634), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5637) );
  INV_X2 U7241 ( .A(n5635), .ZN(n5722) );
  NAND2_X1 U7242 ( .A1(n6239), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5636) );
  NAND2_X1 U7243 ( .A1(n8734), .A2(n6021), .ZN(n5650) );
  OR2_X1 U7244 ( .A1(n5961), .A2(n4905), .ZN(n5647) );
  INV_X1 U7245 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5642) );
  NAND2_X1 U7246 ( .A1(n5643), .A2(n5642), .ZN(n5644) );
  NAND2_X1 U7247 ( .A1(n5644), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5645) );
  XNOR2_X1 U7248 ( .A(n5645), .B(P1_IR_REG_3__SCAN_IN), .ZN(n8777) );
  NAND2_X1 U7249 ( .A1(n5619), .A2(n8777), .ZN(n5646) );
  OAI211_X1 U7250 ( .C1(n6283), .C2(n5734), .A(n5647), .B(n5646), .ZN(n8315)
         );
  NAND2_X1 U7251 ( .A1(n5650), .A2(n5649), .ZN(n5651) );
  AND2_X1 U7252 ( .A1(n8315), .A2(n6080), .ZN(n5652) );
  AOI21_X1 U7253 ( .B1(n8734), .B2(n6145), .A(n5652), .ZN(n5654) );
  XNOR2_X1 U7254 ( .A(n5653), .B(n5654), .ZN(n8313) );
  INV_X1 U7255 ( .A(n5653), .ZN(n5655) );
  NAND2_X1 U7256 ( .A1(n5655), .A2(n5654), .ZN(n5656) );
  NOR2_X1 U7257 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5658) );
  NOR2_X1 U7258 ( .A1(n5681), .A2(n5658), .ZN(n6867) );
  NAND2_X1 U7259 ( .A1(n6134), .A2(n6867), .ZN(n5662) );
  NAND2_X1 U7260 ( .A1(n4265), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U7261 ( .A1(n6239), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5660) );
  NAND2_X1 U7262 ( .A1(n5634), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5659) );
  NAND4_X1 U7263 ( .A1(n5662), .A2(n5661), .A3(n5660), .A4(n5659), .ZN(n8733)
         );
  NAND2_X1 U7264 ( .A1(n8733), .A2(n6021), .ZN(n5668) );
  OR2_X1 U7265 ( .A1(n5734), .A2(n6303), .ZN(n5666) );
  OR2_X1 U7266 ( .A1(n5822), .A2(n9490), .ZN(n5663) );
  XNOR2_X1 U7267 ( .A(n5663), .B(n5676), .ZN(n6543) );
  OAI22_X1 U7268 ( .A1(n5961), .A2(n6304), .B1(n6289), .B2(n6543), .ZN(n5664)
         );
  INV_X1 U7269 ( .A(n5664), .ZN(n5665) );
  NAND2_X1 U7270 ( .A1(n5666), .A2(n5665), .ZN(n6454) );
  NAND2_X1 U7271 ( .A1(n6454), .A2(n6133), .ZN(n5667) );
  NAND2_X1 U7272 ( .A1(n5668), .A2(n5667), .ZN(n5669) );
  AOI22_X1 U7273 ( .A1(n8733), .A2(n6145), .B1(n6021), .B2(n6454), .ZN(n5672)
         );
  XNOR2_X1 U7274 ( .A(n5671), .B(n5672), .ZN(n6423) );
  INV_X1 U7275 ( .A(n5671), .ZN(n5674) );
  INV_X1 U7276 ( .A(n5672), .ZN(n5673) );
  NAND2_X1 U7277 ( .A1(n5674), .A2(n5673), .ZN(n5675) );
  OR2_X1 U7278 ( .A1(n6305), .A2(n5734), .ZN(n5680) );
  NAND2_X1 U7279 ( .A1(n5822), .A2(n5676), .ZN(n5695) );
  NAND2_X1 U7280 ( .A1(n5695), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5677) );
  XNOR2_X1 U7281 ( .A(n5677), .B(n5819), .ZN(n6544) );
  OAI22_X1 U7282 ( .A1(n5961), .A2(n6306), .B1(n6289), .B2(n6544), .ZN(n5678)
         );
  INV_X1 U7283 ( .A(n5678), .ZN(n5679) );
  NAND2_X1 U7284 ( .A1(n5680), .A2(n5679), .ZN(n8450) );
  NAND2_X1 U7285 ( .A1(n8450), .A2(n6022), .ZN(n5688) );
  OAI21_X1 U7286 ( .B1(n5681), .B2(P1_REG3_REG_5__SCAN_IN), .A(n5702), .ZN(
        n6705) );
  INV_X1 U7287 ( .A(n6705), .ZN(n5682) );
  NAND2_X1 U7288 ( .A1(n6134), .A2(n5682), .ZN(n5686) );
  NAND2_X1 U7289 ( .A1(n4265), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5685) );
  INV_X2 U7290 ( .A(n6092), .ZN(n8553) );
  NAND2_X1 U7291 ( .A1(n8553), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5684) );
  NAND2_X1 U7292 ( .A1(n8554), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5683) );
  NAND4_X1 U7293 ( .A1(n5686), .A2(n5685), .A3(n5684), .A4(n5683), .ZN(n8732)
         );
  NAND2_X1 U7294 ( .A1(n8732), .A2(n6021), .ZN(n5687) );
  NAND2_X1 U7295 ( .A1(n5688), .A2(n5687), .ZN(n5689) );
  XNOR2_X1 U7296 ( .A(n5689), .B(n4259), .ZN(n5709) );
  NAND2_X1 U7297 ( .A1(n8450), .A2(n6021), .ZN(n5691) );
  NAND2_X1 U7298 ( .A1(n8732), .A2(n4359), .ZN(n5690) );
  NAND2_X1 U7299 ( .A1(n5691), .A2(n5690), .ZN(n6575) );
  INV_X1 U7300 ( .A(n6575), .ZN(n5692) );
  NAND2_X1 U7301 ( .A1(n6572), .A2(n5694), .ZN(n5712) );
  OR2_X1 U7302 ( .A1(n6301), .A2(n5734), .ZN(n5700) );
  INV_X1 U7303 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6302) );
  NOR2_X1 U7304 ( .A1(n5695), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5736) );
  OR2_X1 U7305 ( .A1(n5736), .A2(n9490), .ZN(n5696) );
  NAND2_X1 U7306 ( .A1(n5696), .A2(n5818), .ZN(n5716) );
  OR2_X1 U7307 ( .A1(n5696), .A2(n5818), .ZN(n5697) );
  INV_X1 U7308 ( .A(n9587), .ZN(n6300) );
  OAI22_X1 U7309 ( .A1(n5961), .A2(n6302), .B1(n6289), .B2(n6300), .ZN(n5698)
         );
  INV_X1 U7310 ( .A(n5698), .ZN(n5699) );
  NAND2_X1 U7311 ( .A1(n4264), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5707) );
  AND2_X1 U7312 ( .A1(n5702), .A2(n5701), .ZN(n5703) );
  NOR2_X1 U7313 ( .A1(n5720), .A2(n5703), .ZN(n6875) );
  NAND2_X1 U7314 ( .A1(n5657), .A2(n6875), .ZN(n5706) );
  NAND2_X1 U7315 ( .A1(n8553), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5705) );
  NAND2_X1 U7316 ( .A1(n6239), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5704) );
  AOI22_X1 U7317 ( .A1(n8458), .A2(n6080), .B1(n4359), .B2(n8731), .ZN(n5713)
         );
  AOI22_X1 U7318 ( .A1(n8458), .A2(n6133), .B1(n6021), .B2(n8731), .ZN(n5708)
         );
  XNOR2_X1 U7319 ( .A(n5708), .B(n4259), .ZN(n5714) );
  XOR2_X1 U7320 ( .A(n5713), .B(n5714), .Z(n6590) );
  NAND2_X1 U7321 ( .A1(n5709), .A2(n6575), .ZN(n5710) );
  NAND2_X1 U7322 ( .A1(n5712), .A2(n5711), .ZN(n6592) );
  NAND2_X1 U7323 ( .A1(n5714), .A2(n5713), .ZN(n5715) );
  NAND2_X1 U7324 ( .A1(n5716), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5717) );
  XNOR2_X1 U7325 ( .A(n5717), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9543) );
  AOI22_X1 U7326 ( .A1(n6235), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5619), .B2(
        n9543), .ZN(n5718) );
  NOR2_X1 U7327 ( .A1(n5720), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5721) );
  OR2_X1 U7328 ( .A1(n5742), .A2(n5721), .ZN(n6694) );
  INV_X1 U7329 ( .A(n6694), .ZN(n6898) );
  NAND2_X1 U7330 ( .A1(n6134), .A2(n6898), .ZN(n5726) );
  NAND2_X1 U7331 ( .A1(n4264), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5725) );
  NAND2_X1 U7332 ( .A1(n8553), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5724) );
  INV_X2 U7333 ( .A(n5722), .ZN(n6239) );
  NAND2_X1 U7334 ( .A1(n6239), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5723) );
  NAND4_X1 U7335 ( .A1(n5726), .A2(n5725), .A3(n5724), .A4(n5723), .ZN(n8730)
         );
  AOI22_X1 U7336 ( .A1(n9676), .A2(n6022), .B1(n6080), .B2(n8730), .ZN(n5727)
         );
  XNOR2_X1 U7337 ( .A(n5727), .B(n4259), .ZN(n5728) );
  AOI22_X1 U7338 ( .A1(n9676), .A2(n6080), .B1(n4359), .B2(n8730), .ZN(n5729)
         );
  XNOR2_X1 U7339 ( .A(n5728), .B(n5729), .ZN(n6697) );
  INV_X1 U7340 ( .A(n5728), .ZN(n5731) );
  INV_X1 U7341 ( .A(n5729), .ZN(n5730) );
  INV_X2 U7342 ( .A(n5734), .ZN(n5959) );
  NOR2_X1 U7343 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5735) );
  NAND2_X1 U7344 ( .A1(n5736), .A2(n5735), .ZN(n5738) );
  NAND2_X1 U7345 ( .A1(n5738), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5737) );
  MUX2_X1 U7346 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5737), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n5739) );
  INV_X1 U7347 ( .A(n6549), .ZN(n9557) );
  OAI22_X1 U7348 ( .A1(n5961), .A2(n6311), .B1(n6289), .B2(n9557), .ZN(n5740)
         );
  INV_X1 U7349 ( .A(n5740), .ZN(n5741) );
  NAND2_X1 U7350 ( .A1(n6942), .A2(n6022), .ZN(n5749) );
  NOR2_X1 U7351 ( .A1(n5742), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5743) );
  NAND2_X1 U7352 ( .A1(n6134), .A2(n4820), .ZN(n5747) );
  NAND2_X1 U7353 ( .A1(n4264), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5746) );
  NAND2_X1 U7354 ( .A1(n6239), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5745) );
  NAND2_X1 U7355 ( .A1(n8553), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5744) );
  NAND4_X1 U7356 ( .A1(n5747), .A2(n5746), .A3(n5745), .A4(n5744), .ZN(n8729)
         );
  NAND2_X1 U7357 ( .A1(n8729), .A2(n6021), .ZN(n5748) );
  NAND2_X1 U7358 ( .A1(n5749), .A2(n5748), .ZN(n5750) );
  XNOR2_X1 U7359 ( .A(n5750), .B(n4266), .ZN(n7019) );
  NAND2_X1 U7360 ( .A1(n6942), .A2(n6080), .ZN(n5752) );
  NAND2_X1 U7361 ( .A1(n8729), .A2(n4359), .ZN(n5751) );
  AND2_X1 U7362 ( .A1(n5752), .A2(n5751), .ZN(n5768) );
  NAND2_X1 U7363 ( .A1(n6323), .A2(n5959), .ZN(n5757) );
  NAND2_X1 U7364 ( .A1(n5776), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5754) );
  XNOR2_X1 U7365 ( .A(n5754), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7006) );
  INV_X1 U7366 ( .A(n7006), .ZN(n6557) );
  OAI22_X1 U7367 ( .A1(n5961), .A2(n6324), .B1(n6289), .B2(n6557), .ZN(n5755)
         );
  INV_X1 U7368 ( .A(n5755), .ZN(n5756) );
  NAND2_X1 U7369 ( .A1(n6919), .A2(n6022), .ZN(n5765) );
  OR2_X1 U7370 ( .A1(n5758), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5759) );
  AND2_X1 U7371 ( .A1(n5783), .A2(n5759), .ZN(n7026) );
  NAND2_X1 U7372 ( .A1(n6134), .A2(n7026), .ZN(n5763) );
  NAND2_X1 U7373 ( .A1(n4264), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5762) );
  NAND2_X1 U7374 ( .A1(n8553), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5761) );
  NAND2_X1 U7375 ( .A1(n6239), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5760) );
  NAND4_X1 U7376 ( .A1(n5763), .A2(n5762), .A3(n5761), .A4(n5760), .ZN(n8728)
         );
  NAND2_X1 U7377 ( .A1(n8728), .A2(n6080), .ZN(n5764) );
  NAND2_X1 U7378 ( .A1(n5765), .A2(n5764), .ZN(n5766) );
  XNOR2_X1 U7379 ( .A(n5766), .B(n4259), .ZN(n5772) );
  AND2_X1 U7380 ( .A1(n8728), .A2(n4359), .ZN(n5767) );
  AOI21_X1 U7381 ( .B1(n6919), .B2(n6021), .A(n5767), .ZN(n5773) );
  XNOR2_X1 U7382 ( .A(n5772), .B(n5773), .ZN(n7021) );
  INV_X1 U7383 ( .A(n7019), .ZN(n5769) );
  INV_X1 U7384 ( .A(n5768), .ZN(n6937) );
  AND2_X1 U7385 ( .A1(n7021), .A2(n4334), .ZN(n5770) );
  NAND2_X1 U7386 ( .A1(n6325), .A2(n5959), .ZN(n5781) );
  NAND2_X1 U7387 ( .A1(n5777), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5778) );
  OR2_X1 U7388 ( .A1(n5778), .A2(n5817), .ZN(n5779) );
  NAND2_X1 U7389 ( .A1(n5778), .A2(n5817), .ZN(n5795) );
  AOI22_X1 U7390 ( .A1(n6235), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5619), .B2(
        n9532), .ZN(n5780) );
  NAND2_X1 U7391 ( .A1(n5781), .A2(n5780), .ZN(n6970) );
  NAND2_X1 U7392 ( .A1(n5783), .A2(n5782), .ZN(n5784) );
  NAND2_X1 U7393 ( .A1(n5801), .A2(n5784), .ZN(n9576) );
  INV_X1 U7394 ( .A(n9576), .ZN(n5785) );
  NAND2_X1 U7395 ( .A1(n6134), .A2(n5785), .ZN(n5789) );
  NAND2_X1 U7396 ( .A1(n4265), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5788) );
  NAND2_X1 U7397 ( .A1(n8553), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5787) );
  NAND2_X1 U7398 ( .A1(n6239), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5786) );
  NAND4_X1 U7399 ( .A1(n5789), .A2(n5788), .A3(n5787), .A4(n5786), .ZN(n8727)
         );
  AOI22_X1 U7400 ( .A1(n6970), .A2(n6022), .B1(n6021), .B2(n8727), .ZN(n5790)
         );
  XOR2_X1 U7401 ( .A(n4259), .B(n5790), .Z(n5791) );
  NOR2_X2 U7402 ( .A1(n5792), .A2(n5791), .ZN(n5794) );
  AOI22_X1 U7403 ( .A1(n6970), .A2(n6080), .B1(n4359), .B2(n8727), .ZN(n9564)
         );
  NAND2_X1 U7404 ( .A1(n9563), .A2(n9564), .ZN(n9562) );
  NAND2_X1 U7405 ( .A1(n6332), .A2(n5959), .ZN(n5798) );
  NAND2_X1 U7406 ( .A1(n5795), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5796) );
  XNOR2_X1 U7407 ( .A(n5796), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7008) );
  AOI22_X1 U7408 ( .A1(n6235), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5619), .B2(
        n7008), .ZN(n5797) );
  NAND2_X1 U7409 ( .A1(n7110), .A2(n6022), .ZN(n5808) );
  INV_X1 U7410 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5800) );
  NAND2_X1 U7411 ( .A1(n5801), .A2(n5800), .ZN(n5802) );
  AND2_X1 U7412 ( .A1(n5851), .A2(n5802), .ZN(n7165) );
  NAND2_X1 U7413 ( .A1(n6134), .A2(n7165), .ZN(n5806) );
  NAND2_X1 U7414 ( .A1(n4265), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5805) );
  NAND2_X1 U7415 ( .A1(n8553), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5804) );
  NAND2_X1 U7416 ( .A1(n6239), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5803) );
  NAND4_X1 U7417 ( .A1(n5806), .A2(n5805), .A3(n5804), .A4(n5803), .ZN(n8726)
         );
  NAND2_X1 U7418 ( .A1(n8726), .A2(n6080), .ZN(n5807) );
  NAND2_X1 U7419 ( .A1(n5808), .A2(n5807), .ZN(n5809) );
  XNOR2_X1 U7420 ( .A(n5809), .B(n4266), .ZN(n5811) );
  AND2_X1 U7421 ( .A1(n8726), .A2(n4359), .ZN(n5810) );
  AOI21_X1 U7422 ( .B1(n7110), .B2(n6080), .A(n5810), .ZN(n5812) );
  NAND2_X1 U7423 ( .A1(n5811), .A2(n5812), .ZN(n5816) );
  INV_X1 U7424 ( .A(n5811), .ZN(n5814) );
  INV_X1 U7425 ( .A(n5812), .ZN(n5813) );
  NAND2_X1 U7426 ( .A1(n5814), .A2(n5813), .ZN(n5815) );
  NAND2_X1 U7427 ( .A1(n5816), .A2(n5815), .ZN(n7159) );
  INV_X1 U7428 ( .A(n5816), .ZN(n7227) );
  NAND2_X1 U7429 ( .A1(n6369), .A2(n5959), .ZN(n5827) );
  INV_X1 U7430 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6370) );
  NAND3_X1 U7431 ( .A1(n5819), .A2(n5818), .A3(n5817), .ZN(n5820) );
  NOR2_X1 U7432 ( .A1(n5820), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5823) );
  AND3_X1 U7433 ( .A1(n5823), .A2(n5822), .A3(n5821), .ZN(n5843) );
  OR2_X1 U7434 ( .A1(n5843), .A2(n9490), .ZN(n5824) );
  XNOR2_X1 U7435 ( .A(n5824), .B(P1_IR_REG_12__SCAN_IN), .ZN(n8819) );
  INV_X1 U7436 ( .A(n8819), .ZN(n7013) );
  OAI22_X1 U7437 ( .A1(n5961), .A2(n6370), .B1(n6289), .B2(n7013), .ZN(n5825)
         );
  INV_X1 U7438 ( .A(n5825), .ZN(n5826) );
  NAND2_X1 U7439 ( .A1(n7175), .A2(n6022), .ZN(n5833) );
  NAND2_X1 U7440 ( .A1(n4264), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5831) );
  XNOR2_X1 U7441 ( .A(n5851), .B(P1_REG3_REG_12__SCAN_IN), .ZN(n7234) );
  NAND2_X1 U7442 ( .A1(n6134), .A2(n7234), .ZN(n5830) );
  NAND2_X1 U7443 ( .A1(n8553), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5829) );
  NAND2_X1 U7444 ( .A1(n6239), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5828) );
  NAND4_X1 U7445 ( .A1(n5831), .A2(n5830), .A3(n5829), .A4(n5828), .ZN(n7206)
         );
  NAND2_X1 U7446 ( .A1(n7206), .A2(n6021), .ZN(n5832) );
  NAND2_X1 U7447 ( .A1(n5833), .A2(n5832), .ZN(n5834) );
  XNOR2_X1 U7448 ( .A(n5834), .B(n4266), .ZN(n5836) );
  AND2_X1 U7449 ( .A1(n7206), .A2(n4359), .ZN(n5835) );
  AOI21_X1 U7450 ( .B1(n7175), .B2(n6080), .A(n5835), .ZN(n5837) );
  NAND2_X1 U7451 ( .A1(n5836), .A2(n5837), .ZN(n5841) );
  INV_X1 U7452 ( .A(n5836), .ZN(n5839) );
  INV_X1 U7453 ( .A(n5837), .ZN(n5838) );
  NAND2_X1 U7454 ( .A1(n5839), .A2(n5838), .ZN(n5840) );
  AND2_X1 U7455 ( .A1(n5841), .A2(n5840), .ZN(n7226) );
  NAND2_X1 U7456 ( .A1(n6373), .A2(n5959), .ZN(n5848) );
  INV_X1 U7457 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6376) );
  NAND2_X1 U7458 ( .A1(n5843), .A2(n5842), .ZN(n5863) );
  NAND2_X1 U7459 ( .A1(n5863), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5845) );
  INV_X1 U7460 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5844) );
  XNOR2_X1 U7461 ( .A(n5845), .B(n5844), .ZN(n8821) );
  OAI22_X1 U7462 ( .A1(n5961), .A2(n6376), .B1(n6289), .B2(n8821), .ZN(n5846)
         );
  INV_X1 U7463 ( .A(n5846), .ZN(n5847) );
  NAND2_X1 U7464 ( .A1(n4264), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5856) );
  OAI21_X1 U7465 ( .B1(n5851), .B2(n5849), .A(n5850), .ZN(n5852) );
  AND2_X1 U7466 ( .A1(n5852), .A2(n5872), .ZN(n8391) );
  NAND2_X1 U7467 ( .A1(n6134), .A2(n8391), .ZN(n5855) );
  NAND2_X1 U7468 ( .A1(n8553), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5854) );
  NAND2_X1 U7469 ( .A1(n8554), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5853) );
  NAND4_X1 U7470 ( .A1(n5856), .A2(n5855), .A3(n5854), .A4(n5853), .ZN(n8725)
         );
  INV_X1 U7471 ( .A(n4359), .ZN(n6026) );
  OAI22_X1 U7472 ( .A1(n8871), .A2(n4253), .B1(n8872), .B2(n6026), .ZN(n5860)
         );
  NAND2_X1 U7473 ( .A1(n9408), .A2(n6022), .ZN(n5858) );
  NAND2_X1 U7474 ( .A1(n8725), .A2(n6080), .ZN(n5857) );
  NAND2_X1 U7475 ( .A1(n5858), .A2(n5857), .ZN(n5859) );
  XNOR2_X1 U7476 ( .A(n5859), .B(n4259), .ZN(n5861) );
  XOR2_X1 U7477 ( .A(n5860), .B(n5861), .Z(n8386) );
  OR2_X1 U7478 ( .A1(n5861), .A2(n5860), .ZN(n5862) );
  NAND2_X1 U7479 ( .A1(n6377), .A2(n5959), .ZN(n5869) );
  OR2_X1 U7480 ( .A1(n5863), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n5864) );
  NAND2_X1 U7481 ( .A1(n5864), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5866) );
  OR2_X1 U7482 ( .A1(n5866), .A2(n5865), .ZN(n5867) );
  NAND2_X1 U7483 ( .A1(n5866), .A2(n5865), .ZN(n5881) );
  AOI22_X1 U7484 ( .A1(n6235), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5619), .B2(
        n9627), .ZN(n5868) );
  NAND2_X1 U7485 ( .A1(n4265), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5877) );
  INV_X1 U7486 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5871) );
  NAND2_X1 U7487 ( .A1(n5872), .A2(n5871), .ZN(n5873) );
  AND2_X1 U7488 ( .A1(n5889), .A2(n5873), .ZN(n9313) );
  NAND2_X1 U7489 ( .A1(n6134), .A2(n9313), .ZN(n5876) );
  NAND2_X1 U7490 ( .A1(n8553), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5875) );
  NAND2_X1 U7491 ( .A1(n6239), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5874) );
  NAND4_X1 U7492 ( .A1(n5877), .A2(n5876), .A3(n5875), .A4(n5874), .ZN(n8724)
         );
  AOI22_X1 U7493 ( .A1(n9311), .A2(n6022), .B1(n6021), .B2(n8724), .ZN(n5878)
         );
  XNOR2_X1 U7494 ( .A(n5878), .B(n4259), .ZN(n5879) );
  AOI22_X1 U7495 ( .A1(n9311), .A2(n6021), .B1(n4359), .B2(n8724), .ZN(n8293)
         );
  NAND2_X1 U7496 ( .A1(n6427), .A2(n5959), .ZN(n5886) );
  INV_X1 U7497 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6429) );
  NAND2_X1 U7498 ( .A1(n5881), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5883) );
  INV_X1 U7499 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5882) );
  XNOR2_X1 U7500 ( .A(n5883), .B(n5882), .ZN(n9631) );
  OAI22_X1 U7501 ( .A1(n5961), .A2(n6429), .B1(n6289), .B2(n9631), .ZN(n5884)
         );
  INV_X1 U7502 ( .A(n5884), .ZN(n5885) );
  INV_X1 U7503 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5888) );
  NAND2_X1 U7504 ( .A1(n5889), .A2(n5888), .ZN(n5890) );
  AND2_X1 U7505 ( .A1(n5903), .A2(n5890), .ZN(n9289) );
  NAND2_X1 U7506 ( .A1(n6134), .A2(n9289), .ZN(n5894) );
  NAND2_X1 U7507 ( .A1(n4265), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5893) );
  NAND2_X1 U7508 ( .A1(n8553), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5892) );
  NAND2_X1 U7509 ( .A1(n8554), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5891) );
  NAND4_X1 U7510 ( .A1(n5894), .A2(n5893), .A3(n5892), .A4(n5891), .ZN(n8876)
         );
  AOI22_X1 U7511 ( .A1(n9396), .A2(n6022), .B1(n6080), .B2(n8876), .ZN(n5895)
         );
  XNOR2_X1 U7512 ( .A(n5895), .B(n4259), .ZN(n5896) );
  AOI22_X1 U7513 ( .A1(n9396), .A2(n6021), .B1(n4359), .B2(n8876), .ZN(n8427)
         );
  NAND2_X1 U7514 ( .A1(n6522), .A2(n5959), .ZN(n5901) );
  INV_X1 U7515 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6523) );
  NAND2_X1 U7516 ( .A1(n5567), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5898) );
  XNOR2_X1 U7517 ( .A(n5898), .B(P1_IR_REG_16__SCAN_IN), .ZN(n8834) );
  INV_X1 U7518 ( .A(n8834), .ZN(n8825) );
  OAI22_X1 U7519 ( .A1(n5961), .A2(n6523), .B1(n6289), .B2(n8825), .ZN(n5899)
         );
  INV_X1 U7520 ( .A(n5899), .ZN(n5900) );
  NAND2_X1 U7521 ( .A1(n9270), .A2(n6022), .ZN(n5910) );
  NAND2_X1 U7522 ( .A1(n4264), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5908) );
  INV_X1 U7523 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5902) );
  NAND2_X1 U7524 ( .A1(n5903), .A2(n5902), .ZN(n5904) );
  AND2_X1 U7525 ( .A1(n5923), .A2(n5904), .ZN(n9271) );
  NAND2_X1 U7526 ( .A1(n9271), .A2(n6134), .ZN(n5907) );
  NAND2_X1 U7527 ( .A1(n8553), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5906) );
  NAND2_X1 U7528 ( .A1(n6239), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5905) );
  NAND4_X1 U7529 ( .A1(n5908), .A2(n5907), .A3(n5906), .A4(n5905), .ZN(n8723)
         );
  NAND2_X1 U7530 ( .A1(n8723), .A2(n6080), .ZN(n5909) );
  NAND2_X1 U7531 ( .A1(n5910), .A2(n5909), .ZN(n5911) );
  XNOR2_X1 U7532 ( .A(n5911), .B(n4259), .ZN(n5914) );
  AOI22_X1 U7533 ( .A1(n9270), .A2(n6021), .B1(n4359), .B2(n8723), .ZN(n5912)
         );
  XNOR2_X1 U7534 ( .A(n5914), .B(n5912), .ZN(n8349) );
  INV_X1 U7535 ( .A(n5912), .ZN(n5913) );
  NAND2_X1 U7536 ( .A1(n8347), .A2(n5915), .ZN(n8355) );
  NAND2_X1 U7537 ( .A1(n6584), .A2(n5959), .ZN(n5920) );
  XNOR2_X1 U7538 ( .A(n5916), .B(n5917), .ZN(n8850) );
  OAI22_X1 U7539 ( .A1(n5961), .A2(n6585), .B1(n6289), .B2(n8850), .ZN(n5918)
         );
  INV_X1 U7540 ( .A(n5918), .ZN(n5919) );
  NAND2_X1 U7541 ( .A1(n9385), .A2(n6022), .ZN(n5930) );
  INV_X1 U7542 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9470) );
  INV_X1 U7543 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5922) );
  NAND2_X1 U7544 ( .A1(n5923), .A2(n5922), .ZN(n5924) );
  NAND2_X1 U7545 ( .A1(n5945), .A2(n5924), .ZN(n9258) );
  OR2_X1 U7546 ( .A1(n9258), .A2(n6111), .ZN(n5928) );
  NAND2_X1 U7547 ( .A1(n8553), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5926) );
  NAND2_X1 U7548 ( .A1(n4264), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5925) );
  AND2_X1 U7549 ( .A1(n5926), .A2(n5925), .ZN(n5927) );
  OAI211_X1 U7550 ( .C1(n5722), .C2(n9470), .A(n5928), .B(n5927), .ZN(n8878)
         );
  NAND2_X1 U7551 ( .A1(n8878), .A2(n6080), .ZN(n5929) );
  NAND2_X1 U7552 ( .A1(n5930), .A2(n5929), .ZN(n5931) );
  XNOR2_X1 U7553 ( .A(n5931), .B(n4259), .ZN(n5934) );
  NAND2_X1 U7554 ( .A1(n9385), .A2(n6080), .ZN(n5933) );
  NAND2_X1 U7555 ( .A1(n8878), .A2(n4359), .ZN(n5932) );
  NAND2_X1 U7556 ( .A1(n5933), .A2(n5932), .ZN(n5935) );
  NAND2_X1 U7557 ( .A1(n5934), .A2(n5935), .ZN(n8356) );
  NAND2_X1 U7558 ( .A1(n8355), .A2(n8356), .ZN(n8354) );
  INV_X1 U7559 ( .A(n5934), .ZN(n5937) );
  INV_X1 U7560 ( .A(n5935), .ZN(n5936) );
  NAND2_X1 U7561 ( .A1(n5937), .A2(n5936), .ZN(n8358) );
  NAND2_X1 U7562 ( .A1(n6675), .A2(n5959), .ZN(n5944) );
  INV_X1 U7563 ( .A(n5938), .ZN(n5939) );
  NAND2_X1 U7564 ( .A1(n5939), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n5941) );
  NAND2_X1 U7565 ( .A1(n5941), .A2(n5940), .ZN(n9653) );
  OAI22_X1 U7566 ( .A1(n5961), .A2(n6712), .B1(n6289), .B2(n9653), .ZN(n5942)
         );
  INV_X1 U7567 ( .A(n5942), .ZN(n5943) );
  NAND2_X1 U7568 ( .A1(n9380), .A2(n6022), .ZN(n5950) );
  INV_X1 U7569 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8418) );
  NAND2_X1 U7570 ( .A1(n5945), .A2(n8418), .ZN(n5946) );
  NAND2_X1 U7571 ( .A1(n5966), .A2(n5946), .ZN(n9243) );
  AOI22_X1 U7572 ( .A1(n8553), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n6239), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n5948) );
  NAND2_X1 U7573 ( .A1(n4264), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5947) );
  OAI211_X1 U7574 ( .C1(n9243), .C2(n6111), .A(n5948), .B(n5947), .ZN(n9225)
         );
  NAND2_X1 U7575 ( .A1(n9225), .A2(n6080), .ZN(n5949) );
  NAND2_X1 U7576 ( .A1(n5950), .A2(n5949), .ZN(n5951) );
  XNOR2_X1 U7577 ( .A(n5951), .B(n4266), .ZN(n8415) );
  AND2_X1 U7578 ( .A1(n9225), .A2(n4359), .ZN(n5952) );
  AOI21_X1 U7579 ( .B1(n9380), .B2(n6080), .A(n5952), .ZN(n8414) );
  INV_X1 U7580 ( .A(n8415), .ZN(n5955) );
  INV_X1 U7581 ( .A(n8414), .ZN(n5954) );
  NAND2_X1 U7582 ( .A1(n6933), .A2(n5959), .ZN(n5964) );
  OAI22_X1 U7583 ( .A1(n5961), .A2(n9142), .B1(n8646), .B2(n6289), .ZN(n5962)
         );
  INV_X1 U7584 ( .A(n5962), .ZN(n5963) );
  NAND2_X1 U7585 ( .A1(n9372), .A2(n6022), .ZN(n5971) );
  INV_X1 U7586 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n8855) );
  INV_X1 U7587 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8324) );
  NAND2_X1 U7588 ( .A1(n5966), .A2(n8324), .ZN(n5967) );
  NAND2_X1 U7589 ( .A1(n5980), .A2(n5967), .ZN(n9216) );
  OR2_X1 U7590 ( .A1(n9216), .A2(n6111), .ZN(n5969) );
  AOI22_X1 U7591 ( .A1(n8553), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n8554), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n5968) );
  OAI211_X1 U7592 ( .C1(n6137), .C2(n8855), .A(n5969), .B(n5968), .ZN(n8883)
         );
  NAND2_X1 U7593 ( .A1(n8883), .A2(n6021), .ZN(n5970) );
  NAND2_X1 U7594 ( .A1(n5971), .A2(n5970), .ZN(n5972) );
  XNOR2_X1 U7595 ( .A(n5972), .B(n4259), .ZN(n8322) );
  NAND2_X1 U7596 ( .A1(n9372), .A2(n6080), .ZN(n5974) );
  NAND2_X1 U7597 ( .A1(n8883), .A2(n4359), .ZN(n5973) );
  NAND2_X1 U7598 ( .A1(n5974), .A2(n5973), .ZN(n8321) );
  NOR2_X1 U7599 ( .A1(n8322), .A2(n8321), .ZN(n5977) );
  INV_X1 U7600 ( .A(n8322), .ZN(n5976) );
  INV_X1 U7601 ( .A(n8321), .ZN(n5975) );
  NAND2_X1 U7602 ( .A1(n7068), .A2(n5959), .ZN(n5979) );
  NAND2_X1 U7603 ( .A1(n6235), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5978) );
  NAND2_X1 U7604 ( .A1(n9205), .A2(n6022), .ZN(n5988) );
  INV_X1 U7605 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8379) );
  NAND2_X1 U7606 ( .A1(n5980), .A2(n8379), .ZN(n5981) );
  NAND2_X1 U7607 ( .A1(n5996), .A2(n5981), .ZN(n9206) );
  OR2_X1 U7608 ( .A1(n9206), .A2(n6111), .ZN(n5986) );
  INV_X1 U7609 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9461) );
  NAND2_X1 U7610 ( .A1(n8553), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5983) );
  NAND2_X1 U7611 ( .A1(n4265), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5982) );
  OAI211_X1 U7612 ( .C1(n9461), .C2(n5722), .A(n5983), .B(n5982), .ZN(n5984)
         );
  INV_X1 U7613 ( .A(n5984), .ZN(n5985) );
  NAND2_X1 U7614 ( .A1(n5986), .A2(n5985), .ZN(n9223) );
  NAND2_X1 U7615 ( .A1(n9223), .A2(n6080), .ZN(n5987) );
  NAND2_X1 U7616 ( .A1(n5988), .A2(n5987), .ZN(n5989) );
  XNOR2_X1 U7617 ( .A(n5989), .B(n4266), .ZN(n5992) );
  AND2_X1 U7618 ( .A1(n9223), .A2(n4359), .ZN(n5990) );
  AOI21_X1 U7619 ( .B1(n9205), .B2(n6080), .A(n5990), .ZN(n5991) );
  NAND2_X1 U7620 ( .A1(n5992), .A2(n5991), .ZN(n5993) );
  OAI21_X1 U7621 ( .B1(n5992), .B2(n5991), .A(n5993), .ZN(n8377) );
  NAND2_X1 U7622 ( .A1(n7078), .A2(n5959), .ZN(n5995) );
  NAND2_X1 U7623 ( .A1(n6235), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5994) );
  INV_X1 U7624 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8334) );
  NAND2_X1 U7625 ( .A1(n5996), .A2(n8334), .ZN(n5997) );
  AND2_X1 U7626 ( .A1(n6014), .A2(n5997), .ZN(n9190) );
  NAND2_X1 U7627 ( .A1(n9190), .A2(n6134), .ZN(n6002) );
  INV_X1 U7628 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9365) );
  NAND2_X1 U7629 ( .A1(n5634), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5999) );
  NAND2_X1 U7630 ( .A1(n8554), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5998) );
  OAI211_X1 U7631 ( .C1(n6137), .C2(n9365), .A(n5999), .B(n5998), .ZN(n6000)
         );
  INV_X1 U7632 ( .A(n6000), .ZN(n6001) );
  NAND2_X1 U7633 ( .A1(n6002), .A2(n6001), .ZN(n9165) );
  OAI22_X1 U7634 ( .A1(n9459), .A2(n4253), .B1(n8887), .B2(n6026), .ZN(n6007)
         );
  NAND2_X1 U7635 ( .A1(n9189), .A2(n6022), .ZN(n6004) );
  NAND2_X1 U7636 ( .A1(n9165), .A2(n6021), .ZN(n6003) );
  NAND2_X1 U7637 ( .A1(n6004), .A2(n6003), .ZN(n6005) );
  XNOR2_X1 U7638 ( .A(n6005), .B(n4259), .ZN(n6006) );
  XOR2_X1 U7639 ( .A(n6007), .B(n6006), .Z(n8331) );
  NAND2_X1 U7640 ( .A1(n8330), .A2(n8331), .ZN(n8329) );
  INV_X1 U7641 ( .A(n6006), .ZN(n6009) );
  INV_X1 U7642 ( .A(n6007), .ZN(n6008) );
  NAND2_X1 U7643 ( .A1(n6009), .A2(n6008), .ZN(n6010) );
  NAND2_X1 U7644 ( .A1(n7178), .A2(n5959), .ZN(n6012) );
  NAND2_X1 U7645 ( .A1(n6235), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6011) );
  INV_X1 U7646 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8397) );
  NAND2_X1 U7647 ( .A1(n6014), .A2(n8397), .ZN(n6015) );
  NAND2_X1 U7648 ( .A1(n6030), .A2(n6015), .ZN(n9171) );
  INV_X1 U7649 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9061) );
  NAND2_X1 U7650 ( .A1(n6239), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6017) );
  NAND2_X1 U7651 ( .A1(n8553), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6016) );
  OAI211_X1 U7652 ( .C1(n9061), .C2(n6137), .A(n6017), .B(n6016), .ZN(n6018)
         );
  INV_X1 U7653 ( .A(n6018), .ZN(n6019) );
  NAND2_X1 U7654 ( .A1(n6020), .A2(n6019), .ZN(n8892) );
  AOI22_X1 U7655 ( .A1(n9452), .A2(n6022), .B1(n6080), .B2(n8892), .ZN(n6023)
         );
  XNOR2_X1 U7656 ( .A(n6023), .B(n4259), .ZN(n6024) );
  INV_X1 U7657 ( .A(n9452), .ZN(n9175) );
  INV_X1 U7658 ( .A(n8892), .ZN(n8891) );
  OAI22_X1 U7659 ( .A1(n9175), .A2(n4253), .B1(n8891), .B2(n6026), .ZN(n8396)
         );
  NAND2_X1 U7660 ( .A1(n7221), .A2(n5959), .ZN(n6028) );
  NAND2_X1 U7661 ( .A1(n6235), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6027) );
  NAND2_X1 U7662 ( .A1(n9447), .A2(n6022), .ZN(n6039) );
  INV_X1 U7663 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8307) );
  NAND2_X1 U7664 ( .A1(n6030), .A2(n8307), .ZN(n6031) );
  NAND2_X1 U7665 ( .A1(n6051), .A2(n6031), .ZN(n9015) );
  INV_X1 U7666 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n6034) );
  NAND2_X1 U7667 ( .A1(n8553), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6033) );
  NAND2_X1 U7668 ( .A1(n8554), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6032) );
  OAI211_X1 U7669 ( .C1(n6034), .C2(n6137), .A(n6033), .B(n6032), .ZN(n6035)
         );
  INV_X1 U7670 ( .A(n6035), .ZN(n6036) );
  NAND2_X1 U7671 ( .A1(n9166), .A2(n6080), .ZN(n6038) );
  NAND2_X1 U7672 ( .A1(n6039), .A2(n6038), .ZN(n6040) );
  XNOR2_X1 U7673 ( .A(n6040), .B(n4266), .ZN(n6042) );
  AND2_X1 U7674 ( .A1(n9166), .A2(n4359), .ZN(n6041) );
  AOI21_X1 U7675 ( .B1(n9447), .B2(n6080), .A(n6041), .ZN(n6043) );
  NAND2_X1 U7676 ( .A1(n6042), .A2(n6043), .ZN(n8367) );
  INV_X1 U7677 ( .A(n6042), .ZN(n6045) );
  INV_X1 U7678 ( .A(n6043), .ZN(n6044) );
  NAND2_X1 U7679 ( .A1(n6045), .A2(n6044), .ZN(n6046) );
  NAND2_X1 U7680 ( .A1(n7238), .A2(n5959), .ZN(n6049) );
  NAND2_X1 U7681 ( .A1(n6235), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6048) );
  NAND2_X2 U7682 ( .A1(n6049), .A2(n6048), .ZN(n9442) );
  NAND2_X1 U7683 ( .A1(n9442), .A2(n6022), .ZN(n6059) );
  INV_X1 U7684 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6050) );
  NAND2_X1 U7685 ( .A1(n6051), .A2(n6050), .ZN(n6052) );
  NAND2_X1 U7686 ( .A1(n8998), .A2(n6134), .ZN(n6057) );
  INV_X1 U7687 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9349) );
  NAND2_X1 U7688 ( .A1(n8553), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6054) );
  NAND2_X1 U7689 ( .A1(n6239), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6053) );
  OAI211_X1 U7690 ( .C1(n9349), .C2(n6137), .A(n6054), .B(n6053), .ZN(n6055)
         );
  INV_X1 U7691 ( .A(n6055), .ZN(n6056) );
  NAND2_X1 U7692 ( .A1(n6057), .A2(n6056), .ZN(n8898) );
  NAND2_X1 U7693 ( .A1(n8898), .A2(n6080), .ZN(n6058) );
  NAND2_X1 U7694 ( .A1(n6059), .A2(n6058), .ZN(n6060) );
  XNOR2_X1 U7695 ( .A(n6060), .B(n4266), .ZN(n6062) );
  AND2_X1 U7696 ( .A1(n8898), .A2(n4359), .ZN(n6061) );
  AOI21_X1 U7697 ( .B1(n9442), .B2(n6080), .A(n6061), .ZN(n6063) );
  NAND2_X1 U7698 ( .A1(n6062), .A2(n6063), .ZN(n6068) );
  INV_X1 U7699 ( .A(n6062), .ZN(n6065) );
  INV_X1 U7700 ( .A(n6063), .ZN(n6064) );
  NAND2_X1 U7701 ( .A1(n6065), .A2(n6064), .ZN(n6066) );
  NAND2_X1 U7702 ( .A1(n7308), .A2(n5959), .ZN(n6070) );
  NAND2_X1 U7703 ( .A1(n6235), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6069) );
  NAND2_X1 U7704 ( .A1(n9436), .A2(n6022), .ZN(n6082) );
  INV_X1 U7705 ( .A(n6072), .ZN(n6071) );
  NAND2_X1 U7706 ( .A1(n6071), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6087) );
  INV_X1 U7707 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8343) );
  NAND2_X1 U7708 ( .A1(n6072), .A2(n8343), .ZN(n6073) );
  NAND2_X1 U7709 ( .A1(n6087), .A2(n6073), .ZN(n8983) );
  INV_X1 U7710 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U7711 ( .A1(n8553), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6075) );
  NAND2_X1 U7712 ( .A1(n8554), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6074) );
  OAI211_X1 U7713 ( .C1(n6137), .C2(n6076), .A(n6075), .B(n6074), .ZN(n6077)
         );
  INV_X1 U7714 ( .A(n6077), .ZN(n6078) );
  NAND2_X1 U7715 ( .A1(n8995), .A2(n6021), .ZN(n6081) );
  NAND2_X1 U7716 ( .A1(n6082), .A2(n6081), .ZN(n6083) );
  XNOR2_X1 U7717 ( .A(n6083), .B(n4259), .ZN(n6100) );
  AOI22_X1 U7718 ( .A1(n9436), .A2(n6080), .B1(n4359), .B2(n8995), .ZN(n6101)
         );
  XNOR2_X1 U7719 ( .A(n6100), .B(n6101), .ZN(n8339) );
  NAND2_X1 U7720 ( .A1(n7311), .A2(n5959), .ZN(n6085) );
  NAND2_X1 U7721 ( .A1(n6235), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6084) );
  NAND2_X1 U7722 ( .A1(n9340), .A2(n6022), .ZN(n6097) );
  INV_X1 U7723 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U7724 ( .A1(n6087), .A2(n6086), .ZN(n6088) );
  NAND2_X1 U7725 ( .A1(n8970), .A2(n5657), .ZN(n6095) );
  INV_X1 U7726 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n6091) );
  NAND2_X1 U7727 ( .A1(n4264), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6090) );
  NAND2_X1 U7728 ( .A1(n6239), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6089) );
  OAI211_X1 U7729 ( .C1(n6092), .C2(n6091), .A(n6090), .B(n6089), .ZN(n6093)
         );
  INV_X1 U7730 ( .A(n6093), .ZN(n6094) );
  NAND2_X1 U7731 ( .A1(n6095), .A2(n6094), .ZN(n8722) );
  NAND2_X1 U7732 ( .A1(n8722), .A2(n6080), .ZN(n6096) );
  NAND2_X1 U7733 ( .A1(n6097), .A2(n6096), .ZN(n6098) );
  XNOR2_X1 U7734 ( .A(n6098), .B(n4259), .ZN(n6127) );
  AND2_X1 U7735 ( .A1(n8722), .A2(n4359), .ZN(n6099) );
  AOI21_X1 U7736 ( .B1(n9340), .B2(n5590), .A(n6099), .ZN(n6125) );
  XNOR2_X1 U7737 ( .A(n6127), .B(n6125), .ZN(n6262) );
  INV_X1 U7738 ( .A(n6100), .ZN(n6102) );
  NAND2_X1 U7739 ( .A1(n6102), .A2(n6101), .ZN(n6261) );
  NAND2_X1 U7740 ( .A1(n6104), .A2(n5959), .ZN(n6106) );
  NAND2_X1 U7741 ( .A1(n6235), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6105) );
  NAND2_X1 U7742 ( .A1(n9427), .A2(n6022), .ZN(n6118) );
  INV_X1 U7743 ( .A(n6109), .ZN(n6107) );
  NAND2_X1 U7744 ( .A1(n6107), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n8911) );
  INV_X1 U7745 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6108) );
  NAND2_X1 U7746 ( .A1(n6109), .A2(n6108), .ZN(n6110) );
  NAND2_X1 U7747 ( .A1(n8911), .A2(n6110), .ZN(n8286) );
  INV_X1 U7748 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9121) );
  NAND2_X1 U7749 ( .A1(n8553), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6113) );
  NAND2_X1 U7750 ( .A1(n4265), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6112) );
  OAI211_X1 U7751 ( .C1(n5722), .C2(n9121), .A(n6113), .B(n6112), .ZN(n6114)
         );
  INV_X1 U7752 ( .A(n6114), .ZN(n6115) );
  NAND2_X1 U7753 ( .A1(n8721), .A2(n6021), .ZN(n6117) );
  NAND2_X1 U7754 ( .A1(n6118), .A2(n6117), .ZN(n6119) );
  XNOR2_X1 U7755 ( .A(n6119), .B(n4266), .ZN(n6122) );
  INV_X1 U7756 ( .A(n6122), .ZN(n6124) );
  AND2_X1 U7757 ( .A1(n8721), .A2(n4359), .ZN(n6120) );
  AOI21_X1 U7758 ( .B1(n9427), .B2(n5590), .A(n6120), .ZN(n6121) );
  INV_X1 U7759 ( .A(n6121), .ZN(n6123) );
  AOI21_X1 U7760 ( .B1(n6124), .B2(n6123), .A(n6177), .ZN(n8280) );
  INV_X1 U7761 ( .A(n8280), .ZN(n6129) );
  INV_X1 U7762 ( .A(n6125), .ZN(n6126) );
  NAND2_X1 U7763 ( .A1(n6127), .A2(n6126), .ZN(n8281) );
  INV_X1 U7764 ( .A(n8281), .ZN(n6128) );
  NOR2_X1 U7765 ( .A1(n6129), .A2(n6128), .ZN(n6130) );
  INV_X1 U7766 ( .A(n6176), .ZN(n8284) );
  NAND2_X1 U7767 ( .A1(n7354), .A2(n5959), .ZN(n6132) );
  NAND2_X1 U7768 ( .A1(n6235), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6131) );
  NAND2_X1 U7769 ( .A1(n9331), .A2(n6022), .ZN(n6142) );
  XNOR2_X1 U7770 ( .A(n8911), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n8941) );
  NAND2_X1 U7771 ( .A1(n8941), .A2(n6134), .ZN(n6140) );
  INV_X1 U7772 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9332) );
  NAND2_X1 U7773 ( .A1(n8553), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6136) );
  NAND2_X1 U7774 ( .A1(n8554), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6135) );
  OAI211_X1 U7775 ( .C1(n6137), .C2(n9332), .A(n6136), .B(n6135), .ZN(n6138)
         );
  INV_X1 U7776 ( .A(n6138), .ZN(n6139) );
  NAND2_X1 U7777 ( .A1(n6140), .A2(n6139), .ZN(n8908) );
  NAND2_X1 U7778 ( .A1(n8908), .A2(n5590), .ZN(n6141) );
  NAND2_X1 U7779 ( .A1(n6142), .A2(n6141), .ZN(n6144) );
  XNOR2_X1 U7780 ( .A(n6144), .B(n4259), .ZN(n6147) );
  AOI22_X1 U7781 ( .A1(n9331), .A2(n5590), .B1(n4359), .B2(n8908), .ZN(n6146)
         );
  XNOR2_X1 U7782 ( .A(n6147), .B(n6146), .ZN(n6178) );
  NAND2_X1 U7783 ( .A1(n7310), .A2(P1_B_REG_SCAN_IN), .ZN(n6148) );
  MUX2_X1 U7784 ( .A(P1_B_REG_SCAN_IN), .B(n6148), .S(n7240), .Z(n6149) );
  NAND2_X1 U7785 ( .A1(n6150), .A2(n6149), .ZN(n9487) );
  NAND2_X1 U7786 ( .A1(n7240), .A2(n6151), .ZN(n9489) );
  INV_X1 U7787 ( .A(n6678), .ZN(n6164) );
  NOR4_X1 U7788 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6155) );
  NOR4_X1 U7789 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n6154) );
  NOR4_X1 U7790 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6153) );
  NOR4_X1 U7791 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6152) );
  AND4_X1 U7792 ( .A1(n6155), .A2(n6154), .A3(n6153), .A4(n6152), .ZN(n6161)
         );
  NOR2_X1 U7793 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .ZN(
        n6159) );
  NOR4_X1 U7794 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n6158) );
  NOR4_X1 U7795 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n6157) );
  NOR4_X1 U7796 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n6156) );
  AND4_X1 U7797 ( .A1(n6159), .A2(n6158), .A3(n6157), .A4(n6156), .ZN(n6160)
         );
  NAND2_X1 U7798 ( .A1(n6161), .A2(n6160), .ZN(n6245) );
  INV_X1 U7799 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9141) );
  NOR2_X1 U7800 ( .A1(n6245), .A2(n9141), .ZN(n6162) );
  NAND2_X1 U7801 ( .A1(n6151), .A2(n7310), .ZN(n9488) );
  OAI21_X1 U7802 ( .B1(n9487), .B2(n6162), .A(n9488), .ZN(n6163) );
  INV_X1 U7803 ( .A(n6163), .ZN(n6680) );
  NAND2_X1 U7804 ( .A1(n6164), .A2(n6680), .ZN(n6189) );
  INV_X1 U7805 ( .A(n6189), .ZN(n6170) );
  NAND2_X1 U7806 ( .A1(n6166), .A2(n6165), .ZN(n6167) );
  NAND2_X1 U7807 ( .A1(n6167), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6169) );
  XNOR2_X1 U7808 ( .A(n6169), .B(n6168), .ZN(n6288) );
  NAND2_X1 U7809 ( .A1(n6170), .A2(n9486), .ZN(n6187) );
  NAND2_X1 U7810 ( .A1(n8284), .A2(n6173), .ZN(n6199) );
  INV_X1 U7811 ( .A(n6177), .ZN(n6175) );
  INV_X1 U7812 ( .A(n6178), .ZN(n6174) );
  NAND4_X1 U7813 ( .A1(n6176), .A2(n6175), .A3(n6174), .A4(n9573), .ZN(n6198)
         );
  NAND3_X1 U7814 ( .A1(n6178), .A2(n9573), .A3(n6177), .ZN(n6197) );
  NAND2_X1 U7815 ( .A1(n6345), .A2(n6342), .ZN(n6685) );
  OR2_X1 U7816 ( .A1(n6187), .A2(n6685), .ZN(n6179) );
  NAND2_X2 U7817 ( .A1(n6345), .A2(n4263), .ZN(n9308) );
  INV_X1 U7818 ( .A(n8640), .ZN(n6180) );
  NAND2_X1 U7819 ( .A1(n6134), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n6181) );
  OR2_X1 U7820 ( .A1(n8911), .A2(n6181), .ZN(n6186) );
  NAND2_X1 U7821 ( .A1(n8554), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6184) );
  NAND2_X1 U7822 ( .A1(n8553), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6183) );
  NAND2_X1 U7823 ( .A1(n4264), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6182) );
  AND3_X1 U7824 ( .A1(n6184), .A2(n6183), .A3(n6182), .ZN(n6185) );
  NAND2_X1 U7825 ( .A1(n6186), .A2(n6185), .ZN(n8720) );
  AOI22_X1 U7826 ( .A1(n8721), .A2(n9224), .B1(n9222), .B2(n8720), .ZN(n8936)
         );
  INV_X1 U7827 ( .A(n6188), .ZN(n6248) );
  NAND2_X1 U7828 ( .A1(n6189), .A2(n6248), .ZN(n6192) );
  NAND2_X1 U7829 ( .A1(n8640), .A2(n8707), .ZN(n6190) );
  AND3_X1 U7830 ( .A1(n6191), .A2(n6288), .A3(n6190), .ZN(n6247) );
  NAND2_X1 U7831 ( .A1(n6192), .A2(n6247), .ZN(n6193) );
  INV_X1 U7832 ( .A(n9577), .ZN(n8433) );
  AOI22_X1 U7833 ( .A1(n8941), .A2(n8433), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n6194) );
  OAI21_X1 U7834 ( .B1(n8936), .B2(n8419), .A(n6194), .ZN(n6195) );
  AOI21_X1 U7835 ( .B1(n9331), .B2(n8422), .A(n6195), .ZN(n6196) );
  NAND4_X1 U7836 ( .A1(n6199), .A2(n6198), .A3(n6197), .A4(n6196), .ZN(
        P1_U3220) );
  OAI21_X1 U7837 ( .B1(n6642), .B2(n6201), .A(n6200), .ZN(n6204) );
  NAND2_X1 U7838 ( .A1(n6322), .A2(n6202), .ZN(n6203) );
  NAND2_X1 U7839 ( .A1(n9982), .A2(n9966), .ZN(n8126) );
  INV_X1 U7840 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6207) );
  OAI21_X1 U7841 ( .B1(n6212), .B2(n6211), .A(n6210), .ZN(P2_U3488) );
  INV_X1 U7842 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6251) );
  INV_X1 U7843 ( .A(SI_29_), .ZN(n6213) );
  INV_X1 U7844 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7608) );
  INV_X1 U7845 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n6219) );
  MUX2_X1 U7846 ( .A(n7608), .B(n6219), .S(n6281), .Z(n6221) );
  INV_X1 U7847 ( .A(SI_30_), .ZN(n6220) );
  NAND2_X1 U7848 ( .A1(n6221), .A2(n6220), .ZN(n6229) );
  INV_X1 U7849 ( .A(n6221), .ZN(n6222) );
  NAND2_X1 U7850 ( .A1(n6222), .A2(SI_30_), .ZN(n6223) );
  NAND2_X1 U7851 ( .A1(n6229), .A2(n6223), .ZN(n6230) );
  NAND2_X1 U7852 ( .A1(n7607), .A2(n5959), .ZN(n6225) );
  NAND2_X1 U7853 ( .A1(n6235), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n6224) );
  NAND2_X1 U7854 ( .A1(n8275), .A2(n5959), .ZN(n6227) );
  NAND2_X1 U7855 ( .A1(n6235), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6226) );
  NOR2_X1 U7856 ( .A1(n6414), .A2(n6782), .ZN(n6439) );
  AND2_X1 U7857 ( .A1(n6439), .A2(n6994), .ZN(n6505) );
  NAND2_X1 U7858 ( .A1(n6505), .A2(n7043), .ZN(n6504) );
  NOR2_X1 U7859 ( .A1(n6504), .A2(n6454), .ZN(n6518) );
  NAND2_X1 U7860 ( .A1(n6518), .A2(n8452), .ZN(n6563) );
  INV_X1 U7861 ( .A(n6919), .ZN(n9685) );
  MUX2_X1 U7862 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n6281), .Z(n6232) );
  INV_X1 U7863 ( .A(SI_31_), .ZN(n9091) );
  XNOR2_X1 U7864 ( .A(n6232), .B(n9091), .ZN(n6233) );
  NAND2_X1 U7865 ( .A1(n8268), .A2(n5959), .ZN(n6237) );
  NAND2_X1 U7866 ( .A1(n6235), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U7867 ( .A1(n4264), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6242) );
  NAND2_X1 U7868 ( .A1(n5634), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6241) );
  NAND2_X1 U7869 ( .A1(n6239), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6240) );
  AND3_X1 U7870 ( .A1(n6242), .A2(n6241), .A3(n6240), .ZN(n8637) );
  INV_X1 U7871 ( .A(P1_B_REG_SCAN_IN), .ZN(n9148) );
  OR2_X1 U7872 ( .A1(n8748), .A2(n9148), .ZN(n6244) );
  NAND2_X1 U7873 ( .A1(n9222), .A2(n6244), .ZN(n8928) );
  NOR2_X1 U7874 ( .A1(n8637), .A2(n8928), .ZN(n8863) );
  NOR2_X1 U7875 ( .A1(n8862), .A2(n8863), .ZN(n6256) );
  INV_X1 U7876 ( .A(n9487), .ZN(n6246) );
  NAND2_X1 U7877 ( .A1(n6246), .A2(n6245), .ZN(n6250) );
  OAI21_X1 U7878 ( .B1(n9487), .B2(P1_D_REG_1__SCAN_IN), .A(n9488), .ZN(n6249)
         );
  NAND4_X1 U7879 ( .A1(n6250), .A2(n6679), .A3(n6249), .A4(n6248), .ZN(n6254)
         );
  MUX2_X1 U7880 ( .A(n6251), .B(n6256), .S(n9708), .Z(n6253) );
  NAND2_X1 U7881 ( .A1(n6253), .A2(n6252), .ZN(P1_U3553) );
  INV_X1 U7882 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6257) );
  INV_X1 U7883 ( .A(n6254), .ZN(n6255) );
  MUX2_X1 U7884 ( .A(n6257), .B(n6256), .S(n9701), .Z(n6259) );
  NAND2_X1 U7885 ( .A1(n6259), .A2(n6258), .ZN(P1_U3521) );
  NAND2_X1 U7886 ( .A1(n8282), .A2(n9573), .ZN(n6269) );
  NAND2_X1 U7887 ( .A1(n9340), .A2(n8422), .ZN(n6268) );
  NAND2_X1 U7888 ( .A1(n8721), .A2(n9222), .ZN(n6265) );
  NAND2_X1 U7889 ( .A1(n8995), .A2(n9224), .ZN(n6264) );
  NAND2_X1 U7890 ( .A1(n6265), .A2(n6264), .ZN(n8966) );
  INV_X1 U7891 ( .A(n8419), .ZN(n9568) );
  NAND2_X1 U7892 ( .A1(n8966), .A2(n9568), .ZN(n6267) );
  AOI22_X1 U7893 ( .A1(n8970), .A2(n8433), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n6266) );
  OAI21_X1 U7894 ( .B1(n6270), .B2(n6269), .A(n4830), .ZN(P1_U3240) );
  INV_X1 U7895 ( .A(n6630), .ZN(n7222) );
  NAND2_X1 U7896 ( .A1(n7801), .A2(n6630), .ZN(n6273) );
  NAND2_X1 U7897 ( .A1(n6358), .A2(n6273), .ZN(n6361) );
  OAI21_X1 U7898 ( .B1(n6361), .B2(n6274), .A(P2_STATE_REG_SCAN_IN), .ZN(
        P2_U3150) );
  INV_X1 U7899 ( .A(n6350), .ZN(n6275) );
  AND2_X1 U7900 ( .A1(n6281), .A2(P2_U3151), .ZN(n8273) );
  INV_X2 U7901 ( .A(n8273), .ZN(n8276) );
  AND2_X1 U7902 ( .A1(n6276), .A2(P2_U3151), .ZN(n7353) );
  INV_X2 U7903 ( .A(n7353), .ZN(n8277) );
  INV_X1 U7904 ( .A(n4250), .ZN(n6398) );
  OAI222_X1 U7905 ( .A1(n8276), .A2(n6277), .B1(n8277), .B2(n6285), .C1(n6398), 
        .C2(P2_U3151), .ZN(P2_U3293) );
  OAI222_X1 U7906 ( .A1(n8276), .A2(n6278), .B1(n8277), .B2(n6283), .C1(n6481), 
        .C2(P2_U3151), .ZN(P2_U3292) );
  OAI222_X1 U7907 ( .A1(n8276), .A2(n6279), .B1(n8277), .B2(n6303), .C1(n6607), 
        .C2(P2_U3151), .ZN(P2_U3291) );
  INV_X1 U7908 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6280) );
  OAI222_X1 U7909 ( .A1(P2_U3151), .A2(n6396), .B1(n8277), .B2(n6299), .C1(
        n6280), .C2(n8276), .ZN(P2_U3294) );
  NOR2_X1 U7910 ( .A1(n6281), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9497) );
  AOI22_X1 U7911 ( .A1(n8777), .A2(P1_STATE_REG_SCAN_IN), .B1(n9497), .B2(
        P2_DATAO_REG_3__SCAN_IN), .ZN(n6282) );
  OAI21_X1 U7912 ( .B1(n6283), .B2(n9500), .A(n6282), .ZN(P1_U3352) );
  AOI22_X1 U7913 ( .A1(n9497), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n8760), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6284) );
  OAI21_X1 U7914 ( .B1(n6285), .B2(n9500), .A(n6284), .ZN(P1_U3353) );
  OAI222_X1 U7915 ( .A1(n6847), .A2(P2_U3151), .B1(n8277), .B2(n6305), .C1(
        n6286), .C2(n8276), .ZN(P2_U3290) );
  OAI222_X1 U7916 ( .A1(n7253), .A2(P2_U3151), .B1(n8277), .B2(n6301), .C1(
        n4361), .C2(n8276), .ZN(P2_U3289) );
  INV_X1 U7917 ( .A(n9486), .ZN(n6287) );
  OR2_X1 U7918 ( .A1(n6288), .A2(P1_U3086), .ZN(n8715) );
  NAND2_X1 U7919 ( .A1(n6287), .A2(n8715), .ZN(n6293) );
  NAND2_X1 U7920 ( .A1(n8640), .A2(n6288), .ZN(n6290) );
  AND2_X1 U7921 ( .A1(n6290), .A2(n6289), .ZN(n6292) );
  INV_X1 U7922 ( .A(n6292), .ZN(n6291) );
  NAND2_X1 U7923 ( .A1(n6293), .A2(n6291), .ZN(n9661) );
  INV_X1 U7924 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6298) );
  NAND2_X1 U7925 ( .A1(n6293), .A2(n6292), .ZN(n6540) );
  INV_X1 U7926 ( .A(n6540), .ZN(n6552) );
  INV_X1 U7927 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6294) );
  INV_X1 U7928 ( .A(n6526), .ZN(n8749) );
  OAI21_X1 U7929 ( .B1(n8748), .B2(P1_REG2_REG_0__SCAN_IN), .A(n8749), .ZN(
        n8753) );
  AOI21_X1 U7930 ( .B1(n8748), .B2(n6294), .A(n8753), .ZN(n6295) );
  XNOR2_X1 U7931 ( .A(n6295), .B(n8754), .ZN(n6296) );
  AOI22_X1 U7932 ( .A1(n6552), .A2(n6296), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n6297) );
  OAI21_X1 U7933 ( .B1(n9661), .B2(n6298), .A(n6297), .ZN(P1_U3243) );
  INV_X1 U7934 ( .A(n9497), .ZN(n7398) );
  INV_X1 U7935 ( .A(n8739), .ZN(n6541) );
  OAI222_X1 U7936 ( .A1(n7398), .A2(n4736), .B1(n9500), .B2(n6299), .C1(
        P1_U3086), .C2(n6541), .ZN(P1_U3354) );
  OAI222_X1 U7937 ( .A1(n7398), .A2(n6302), .B1(n9500), .B2(n6301), .C1(
        P1_U3086), .C2(n6300), .ZN(P1_U3349) );
  OAI222_X1 U7938 ( .A1(n7398), .A2(n6304), .B1(n9500), .B2(n6303), .C1(
        P1_U3086), .C2(n6543), .ZN(P1_U3351) );
  OAI222_X1 U7939 ( .A1(n7398), .A2(n6306), .B1(n9500), .B2(n6305), .C1(
        P1_U3086), .C2(n6544), .ZN(P1_U3350) );
  AOI22_X1 U7940 ( .A1(n9543), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n9497), .ZN(n6307) );
  OAI21_X1 U7941 ( .B1(n6309), .B2(n9500), .A(n6307), .ZN(P1_U3348) );
  OAI222_X1 U7942 ( .A1(n7256), .A2(P2_U3151), .B1(n8277), .B2(n6309), .C1(
        n6308), .C2(n8276), .ZN(P2_U3288) );
  INV_X1 U7943 ( .A(n9661), .ZN(n8835) );
  NOR2_X1 U7944 ( .A1(n8835), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U7945 ( .A(n6310), .ZN(n6313) );
  OAI222_X1 U7946 ( .A1(n7398), .A2(n6311), .B1(n9500), .B2(n6313), .C1(
        P1_U3086), .C2(n9557), .ZN(P1_U3347) );
  INV_X1 U7947 ( .A(n9743), .ZN(n7252) );
  OAI222_X1 U7948 ( .A1(n7252), .A2(P2_U3151), .B1(n8277), .B2(n6313), .C1(
        n6312), .C2(n8276), .ZN(P2_U3287) );
  INV_X1 U7949 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6315) );
  NAND2_X1 U7950 ( .A1(n6762), .A2(P1_U3973), .ZN(n6314) );
  OAI21_X1 U7951 ( .B1(P1_U3973), .B2(n6315), .A(n6314), .ZN(P1_U3554) );
  INV_X1 U7952 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6317) );
  INV_X1 U7953 ( .A(n8637), .ZN(n8558) );
  NAND2_X1 U7954 ( .A1(n8558), .A2(P1_U3973), .ZN(n6316) );
  OAI21_X1 U7955 ( .B1(P1_U3973), .B2(n6317), .A(n6316), .ZN(P1_U3585) );
  INV_X1 U7956 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n9138) );
  NAND2_X1 U7957 ( .A1(n8876), .A2(P1_U3973), .ZN(n6318) );
  OAI21_X1 U7958 ( .B1(n9138), .B2(P1_U3973), .A(n6318), .ZN(P1_U3569) );
  INV_X1 U7959 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6372) );
  NAND2_X1 U7960 ( .A1(n7206), .A2(P1_U3973), .ZN(n6319) );
  OAI21_X1 U7961 ( .B1(n6372), .B2(P1_U3973), .A(n6319), .ZN(P1_U3566) );
  NAND2_X1 U7962 ( .A1(n6321), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6320) );
  OAI21_X1 U7963 ( .B1(n6322), .B2(n6321), .A(n6320), .ZN(P2_U3377) );
  INV_X1 U7964 ( .A(n6323), .ZN(n6328) );
  OAI222_X1 U7965 ( .A1(n9500), .A2(n6328), .B1(n6557), .B2(P1_U3086), .C1(
        n6324), .C2(n7398), .ZN(P1_U3346) );
  INV_X1 U7966 ( .A(n6325), .ZN(n6330) );
  AOI22_X1 U7967 ( .A1(n9532), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9497), .ZN(n6326) );
  OAI21_X1 U7968 ( .B1(n6330), .B2(n9500), .A(n6326), .ZN(P1_U3345) );
  OAI222_X1 U7969 ( .A1(P2_U3151), .A2(n7892), .B1(n8277), .B2(n6328), .C1(
        n6327), .C2(n8276), .ZN(P2_U3286) );
  INV_X1 U7970 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n9085) );
  NOR2_X1 U7971 ( .A1(n6347), .A2(n9085), .ZN(P2_U3255) );
  INV_X1 U7972 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n9110) );
  NOR2_X1 U7973 ( .A1(n6347), .A2(n9110), .ZN(P2_U3239) );
  INV_X1 U7974 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n9074) );
  NOR2_X1 U7975 ( .A1(n6347), .A2(n9074), .ZN(P2_U3258) );
  INV_X1 U7976 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n9117) );
  NOR2_X1 U7977 ( .A1(n6347), .A2(n9117), .ZN(P2_U3235) );
  OAI222_X1 U7978 ( .A1(n8276), .A2(n9046), .B1(n8277), .B2(n6330), .C1(
        P2_U3151), .C2(n7895), .ZN(P2_U3285) );
  AND2_X1 U7979 ( .A1(n6331), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U7980 ( .A1(n6331), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U7981 ( .A1(n6331), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U7982 ( .A1(n6331), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U7983 ( .A1(n6331), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U7984 ( .A1(n6331), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U7985 ( .A1(n6331), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U7986 ( .A1(n6331), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U7987 ( .A1(n6331), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  INV_X1 U7988 ( .A(n9778), .ZN(n7898) );
  INV_X1 U7989 ( .A(n6332), .ZN(n6334) );
  OAI222_X1 U7990 ( .A1(n7898), .A2(P2_U3151), .B1(n8277), .B2(n6334), .C1(
        n6333), .C2(n8276), .ZN(P2_U3284) );
  INV_X1 U7991 ( .A(n7008), .ZN(n9602) );
  OAI222_X1 U7992 ( .A1(n7398), .A2(n9022), .B1(n9500), .B2(n6334), .C1(
        P1_U3086), .C2(n9602), .ZN(P1_U3344) );
  INV_X1 U7993 ( .A(n9222), .ZN(n9287) );
  NOR2_X1 U7994 ( .A1(n6441), .A2(n9287), .ZN(n6778) );
  NAND2_X1 U7995 ( .A1(n8716), .A2(n9016), .ZN(n6336) );
  OR2_X1 U7996 ( .A1(n8651), .A2(n4263), .ZN(n6335) );
  OR2_X1 U7997 ( .A1(n8711), .A2(n6338), .ZN(n6340) );
  INV_X1 U7998 ( .A(n6345), .ZN(n6339) );
  AND2_X1 U7999 ( .A1(n6340), .A2(n6339), .ZN(n6777) );
  NAND2_X1 U8000 ( .A1(n8711), .A2(n8707), .ZN(n6341) );
  NAND2_X1 U8001 ( .A1(n6777), .A2(n6341), .ZN(n9305) );
  NAND2_X1 U8002 ( .A1(n9016), .A2(n6171), .ZN(n8561) );
  NAND2_X1 U8003 ( .A1(n9305), .A2(n6433), .ZN(n9689) );
  INV_X1 U8004 ( .A(n9689), .ZN(n9411) );
  INV_X1 U8005 ( .A(n6782), .ZN(n6353) );
  INV_X1 U8006 ( .A(n6761), .ZN(n6343) );
  NAND2_X1 U8007 ( .A1(n6762), .A2(n6353), .ZN(n8652) );
  AND2_X1 U8008 ( .A1(n6343), .A2(n8652), .ZN(n8572) );
  AOI21_X1 U8009 ( .B1(n9283), .B2(n9411), .A(n8572), .ZN(n6344) );
  AOI211_X1 U8010 ( .C1(n6345), .C2(n6782), .A(n6778), .B(n6344), .ZN(n6581)
         );
  NAND2_X1 U8011 ( .A1(n9706), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6346) );
  OAI21_X1 U8012 ( .B1(n6581), .B2(n9706), .A(n6346), .ZN(P1_U3522) );
  AND2_X1 U8013 ( .A1(n6331), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8014 ( .A1(n6331), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8015 ( .A1(n6331), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8016 ( .A1(n6331), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8017 ( .A1(n6331), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8018 ( .A1(n6331), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8019 ( .A1(n6331), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8020 ( .A1(n6331), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8021 ( .A1(n6331), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8022 ( .A1(n6331), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8023 ( .A1(n6331), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8024 ( .A1(n6331), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8025 ( .A1(n6331), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8026 ( .A1(n6331), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8027 ( .A1(n6331), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8028 ( .A1(n6331), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8029 ( .A1(n6331), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  INV_X1 U8030 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9021) );
  INV_X1 U8031 ( .A(n6348), .ZN(n6349) );
  AOI22_X1 U8032 ( .A1(n6331), .A2(n9021), .B1(n6350), .B2(n6349), .ZN(
        P2_U3376) );
  XNOR2_X1 U8033 ( .A(n6352), .B(n6351), .ZN(n8750) );
  NAND2_X1 U8034 ( .A1(n9577), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8408) );
  INV_X1 U8035 ( .A(n8422), .ZN(n9570) );
  OR2_X1 U8036 ( .A1(n8419), .A2(n9287), .ZN(n8429) );
  OAI22_X1 U8037 ( .A1(n9570), .A2(n6353), .B1(n8429), .B2(n6441), .ZN(n6354)
         );
  AOI21_X1 U8038 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n8408), .A(n6354), .ZN(
        n6355) );
  OAI21_X1 U8039 ( .B1(n8424), .B2(n8750), .A(n6355), .ZN(P1_U3232) );
  INV_X1 U8040 ( .A(n6358), .ZN(n6356) );
  INV_X1 U8041 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6368) );
  NAND2_X1 U8042 ( .A1(n7322), .A2(n7811), .ZN(n6357) );
  NOR2_X1 U8043 ( .A1(n6361), .A2(n6357), .ZN(n6360) );
  OR2_X1 U8044 ( .A1(n7811), .A2(P2_U3151), .ZN(n7355) );
  NOR2_X1 U8045 ( .A1(n6358), .A2(n7355), .ZN(n6359) );
  NOR2_X1 U8046 ( .A1(n6361), .A2(n7355), .ZN(n6393) );
  NOR2_X2 U8047 ( .A1(n7833), .A2(n6362), .ZN(n9883) );
  INV_X1 U8048 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9107) );
  OAI21_X1 U8049 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n6363), .A(n7844), .ZN(n6364) );
  OAI21_X1 U8050 ( .B1(n6393), .B2(n9883), .A(n6364), .ZN(n6365) );
  OAI21_X1 U8051 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n6716), .A(n6365), .ZN(n6366) );
  AOI21_X1 U8052 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n9875), .A(n6366), .ZN(n6367) );
  OAI21_X1 U8053 ( .B1(n9720), .B2(n6368), .A(n6367), .ZN(P2_U3182) );
  INV_X1 U8054 ( .A(n6369), .ZN(n6371) );
  OAI222_X1 U8055 ( .A1(n9500), .A2(n6371), .B1(n7013), .B2(P1_U3086), .C1(
        n6370), .C2(n7398), .ZN(P1_U3343) );
  OAI222_X1 U8056 ( .A1(n7900), .A2(P2_U3151), .B1(n8276), .B2(n6372), .C1(
        n6371), .C2(n8277), .ZN(P2_U3283) );
  INV_X1 U8057 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6374) );
  INV_X1 U8058 ( .A(n6373), .ZN(n6375) );
  INV_X1 U8059 ( .A(n9810), .ZN(n7869) );
  OAI222_X1 U8060 ( .A1(n8276), .A2(n6374), .B1(n8277), .B2(n6375), .C1(n7869), 
        .C2(P2_U3151), .ZN(P2_U3282) );
  OAI222_X1 U8061 ( .A1(n7398), .A2(n6376), .B1(n9500), .B2(n6375), .C1(
        P1_U3086), .C2(n8821), .ZN(P1_U3342) );
  INV_X1 U8062 ( .A(n6377), .ZN(n6419) );
  AOI22_X1 U8063 ( .A1(n9627), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n9497), .ZN(n6378) );
  OAI21_X1 U8064 ( .B1(n6419), .B2(n9500), .A(n6378), .ZN(P1_U3341) );
  XNOR2_X1 U8065 ( .A(n6473), .B(n6481), .ZN(n6384) );
  INV_X1 U8066 ( .A(n6381), .ZN(n6382) );
  INV_X1 U8067 ( .A(n6379), .ZN(n6380) );
  XOR2_X1 U8068 ( .A(n6396), .B(n6379), .Z(n7845) );
  XNOR2_X1 U8069 ( .A(n6381), .B(n4250), .ZN(n9710) );
  NAND2_X1 U8070 ( .A1(n9711), .A2(n9710), .ZN(n9709) );
  AOI21_X1 U8071 ( .B1(n6384), .B2(n6383), .A(n6474), .ZN(n6409) );
  INV_X1 U8072 ( .A(n9883), .ZN(n9508) );
  INV_X1 U8073 ( .A(n6481), .ZN(n6476) );
  NOR2_X1 U8074 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n4911), .ZN(n6672) );
  XNOR2_X1 U8075 ( .A(n4250), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n9723) );
  NAND2_X1 U8076 ( .A1(n4881), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6389) );
  NAND2_X1 U8077 ( .A1(n6396), .A2(n6389), .ZN(n6388) );
  INV_X1 U8078 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6385) );
  NAND2_X1 U8079 ( .A1(n6385), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6386) );
  OR2_X1 U8080 ( .A1(n6386), .A2(n4881), .ZN(n6387) );
  NAND2_X1 U8081 ( .A1(n6388), .A2(n6387), .ZN(n7839) );
  NAND2_X1 U8082 ( .A1(n7839), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6390) );
  NAND2_X1 U8083 ( .A1(n6390), .A2(n6389), .ZN(n9722) );
  NAND2_X1 U8084 ( .A1(n9723), .A2(n9722), .ZN(n6392) );
  NAND2_X1 U8085 ( .A1(n6398), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6391) );
  NAND2_X1 U8086 ( .A1(n6392), .A2(n6391), .ZN(n6482) );
  XNOR2_X1 U8087 ( .A(n6482), .B(n6476), .ZN(n6480) );
  XOR2_X1 U8088 ( .A(n6480), .B(P2_REG1_REG_3__SCAN_IN), .Z(n6405) );
  NAND2_X1 U8089 ( .A1(n6393), .A2(n7812), .ZN(n9890) );
  INV_X1 U8090 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7065) );
  NOR2_X1 U8091 ( .A1(n6394), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6395) );
  NAND2_X1 U8092 ( .A1(n4881), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6397) );
  OAI21_X1 U8093 ( .B1(n6396), .B2(n6395), .A(n6397), .ZN(n7836) );
  INV_X1 U8094 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7835) );
  OR2_X1 U8095 ( .A1(n7836), .A2(n7835), .ZN(n7838) );
  NAND2_X1 U8096 ( .A1(n7838), .A2(n6397), .ZN(n9713) );
  XNOR2_X1 U8097 ( .A(n9715), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n9714) );
  NAND2_X1 U8098 ( .A1(n9713), .A2(n9714), .ZN(n9712) );
  NAND2_X1 U8099 ( .A1(n6398), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6399) );
  NAND2_X1 U8100 ( .A1(n9712), .A2(n6399), .ZN(n6400) );
  NAND2_X1 U8101 ( .A1(n6400), .A2(n6481), .ZN(n6490) );
  OR2_X1 U8102 ( .A1(n6400), .A2(n6481), .ZN(n6401) );
  INV_X1 U8103 ( .A(n6492), .ZN(n6402) );
  AOI21_X1 U8104 ( .B1(n7065), .B2(n6403), .A(n6402), .ZN(n6404) );
  OAI22_X1 U8105 ( .A1(n6405), .A2(n9732), .B1(n9890), .B2(n6404), .ZN(n6406)
         );
  AOI211_X1 U8106 ( .C1(n6476), .C2(n9875), .A(n6672), .B(n6406), .ZN(n6408)
         );
  NAND2_X1 U8107 ( .A1(n9874), .A2(P2_ADDR_REG_3__SCAN_IN), .ZN(n6407) );
  OAI211_X1 U8108 ( .C1(n6409), .C2(n9508), .A(n6408), .B(n6407), .ZN(P2_U3185) );
  INV_X1 U8109 ( .A(n6411), .ZN(n6412) );
  AOI21_X1 U8110 ( .B1(n6413), .B2(n6410), .A(n6412), .ZN(n6417) );
  INV_X1 U8111 ( .A(n8429), .ZN(n8407) );
  AOI22_X1 U8112 ( .A1(n8407), .A2(n8735), .B1(n6774), .B2(n8422), .ZN(n6416)
         );
  NOR2_X1 U8113 ( .A1(n8419), .A2(n9285), .ZN(n8409) );
  AOI22_X1 U8114 ( .A1(n8409), .A2(n6762), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n8408), .ZN(n6415) );
  OAI211_X1 U8115 ( .C1(n6417), .C2(n8424), .A(n6416), .B(n6415), .ZN(P1_U3222) );
  INV_X1 U8116 ( .A(n9825), .ZN(n7904) );
  INV_X1 U8117 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6418) );
  OAI222_X1 U8118 ( .A1(n7904), .A2(P2_U3151), .B1(n8277), .B2(n6419), .C1(
        n6418), .C2(n8276), .ZN(P2_U3281) );
  INV_X1 U8119 ( .A(n6420), .ZN(n6421) );
  AOI22_X1 U8120 ( .A1(n9224), .A2(n8734), .B1(n8732), .B2(n9222), .ZN(n6460)
         );
  AOI22_X1 U8121 ( .A1(n8433), .A2(n6867), .B1(n8422), .B2(n6454), .ZN(n6424)
         );
  NAND2_X1 U8122 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n8784) );
  OAI211_X1 U8123 ( .C1(n6460), .C2(n8419), .A(n6424), .B(n8784), .ZN(n6425)
         );
  OR2_X1 U8124 ( .A1(n6426), .A2(n6425), .ZN(P1_U3230) );
  INV_X1 U8125 ( .A(n9841), .ZN(n7866) );
  INV_X1 U8126 ( .A(n6427), .ZN(n6428) );
  OAI222_X1 U8127 ( .A1(n7866), .A2(P2_U3151), .B1(n8277), .B2(n6428), .C1(
        n8276), .C2(n9138), .ZN(P2_U3280) );
  OAI222_X1 U8128 ( .A1(n7398), .A2(n6429), .B1(n9500), .B2(n6428), .C1(
        P1_U3086), .C2(n9631), .ZN(P1_U3340) );
  INV_X1 U8129 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6432) );
  INV_X1 U8130 ( .A(n6470), .ZN(n6713) );
  NOR2_X1 U8131 ( .A1(n6721), .A2(n6470), .ZN(n7664) );
  INV_X1 U8132 ( .A(n7664), .ZN(n7666) );
  NAND2_X1 U8133 ( .A1(n7666), .A2(n7661), .ZN(n6465) );
  OAI21_X1 U8134 ( .B1(n8167), .B2(n9962), .A(n6465), .ZN(n6430) );
  OR2_X1 U8135 ( .A1(n8165), .A2(n8080), .ZN(n6467) );
  OAI211_X1 U8136 ( .C1(n6713), .C2(n9948), .A(n6430), .B(n6467), .ZN(n8179)
         );
  NAND2_X1 U8137 ( .A1(n8179), .A2(n9967), .ZN(n6431) );
  OAI21_X1 U8138 ( .B1(n6432), .B2(n9967), .A(n6431), .ZN(P2_U3390) );
  INV_X1 U8139 ( .A(n6433), .ZN(n9695) );
  NAND2_X1 U8140 ( .A1(n6762), .A2(n6782), .ZN(n6756) );
  NAND2_X1 U8141 ( .A1(n6441), .A2(n9669), .ZN(n6436) );
  NAND2_X1 U8142 ( .A1(n6759), .A2(n6436), .ZN(n6438) );
  NAND2_X1 U8143 ( .A1(n8735), .A2(n6994), .ZN(n8653) );
  OAI21_X1 U8144 ( .B1(n6438), .B2(n8570), .A(n6449), .ZN(n6677) );
  INV_X1 U8145 ( .A(n6439), .ZN(n6771) );
  AOI211_X1 U8146 ( .C1(n8406), .C2(n6771), .A(n9308), .B(n6505), .ZN(n6689)
         );
  NAND2_X1 U8147 ( .A1(n6441), .A2(n6774), .ZN(n6440) );
  XNOR2_X1 U8148 ( .A(n6457), .B(n8570), .ZN(n6444) );
  INV_X1 U8149 ( .A(n9305), .ZN(n6979) );
  INV_X1 U8150 ( .A(n8734), .ZN(n6450) );
  OAI22_X1 U8151 ( .A1(n6441), .A2(n9285), .B1(n6450), .B2(n9287), .ZN(n6442)
         );
  AOI21_X1 U8152 ( .B1(n6677), .B2(n6979), .A(n6442), .ZN(n6443) );
  OAI21_X1 U8153 ( .B1(n9283), .B2(n6444), .A(n6443), .ZN(n6682) );
  AOI211_X1 U8154 ( .C1(n9695), .C2(n6677), .A(n6689), .B(n6682), .ZN(n6997)
         );
  INV_X1 U8155 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6445) );
  OAI22_X1 U8156 ( .A1(n9406), .A2(n6994), .B1(n9403), .B2(n6445), .ZN(n6446)
         );
  INV_X1 U8157 ( .A(n6446), .ZN(n6447) );
  OAI21_X1 U8158 ( .B1(n6997), .B2(n9706), .A(n6447), .ZN(P1_U3524) );
  NAND2_X1 U8159 ( .A1(n6437), .A2(n6994), .ZN(n6448) );
  NAND2_X1 U8160 ( .A1(n6449), .A2(n6448), .ZN(n6501) );
  NAND2_X1 U8161 ( .A1(n6450), .A2(n8315), .ZN(n6458) );
  NAND2_X1 U8162 ( .A1(n8734), .A2(n7043), .ZN(n8654) );
  NAND2_X1 U8163 ( .A1(n6458), .A2(n8654), .ZN(n8574) );
  NAND2_X1 U8164 ( .A1(n6501), .A2(n8574), .ZN(n6500) );
  NAND2_X1 U8165 ( .A1(n6450), .A2(n7043), .ZN(n6451) );
  INV_X1 U8166 ( .A(n8733), .ZN(n6516) );
  NAND2_X1 U8167 ( .A1(n6516), .A2(n6454), .ZN(n8460) );
  INV_X1 U8168 ( .A(n6454), .ZN(n6989) );
  AND2_X1 U8169 ( .A1(n8733), .A2(n6989), .ZN(n8656) );
  INV_X1 U8170 ( .A(n8656), .ZN(n6452) );
  NAND2_X1 U8171 ( .A1(n8460), .A2(n6452), .ZN(n8575) );
  OAI21_X1 U8172 ( .B1(n6453), .B2(n8575), .A(n6511), .ZN(n6871) );
  AOI211_X1 U8173 ( .C1(n6454), .C2(n6504), .A(n9308), .B(n6518), .ZN(n6866)
         );
  INV_X1 U8174 ( .A(n6455), .ZN(n6456) );
  OAI21_X1 U8175 ( .B1(n6457), .B2(n6456), .A(n8653), .ZN(n6502) );
  NAND2_X1 U8176 ( .A1(n6502), .A2(n6458), .ZN(n6459) );
  NAND2_X1 U8177 ( .A1(n6459), .A2(n8654), .ZN(n6515) );
  XOR2_X1 U8178 ( .A(n6515), .B(n8575), .Z(n6461) );
  OAI21_X1 U8179 ( .B1(n6461), .B2(n9283), .A(n6460), .ZN(n6865) );
  AOI211_X1 U8180 ( .C1(n9689), .C2(n6871), .A(n6866), .B(n6865), .ZN(n6992)
         );
  INV_X1 U8181 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6462) );
  OAI22_X1 U8182 ( .A1(n9406), .A2(n6989), .B1(n9403), .B2(n6462), .ZN(n6463)
         );
  INV_X1 U8183 ( .A(n6463), .ZN(n6464) );
  OAI21_X1 U8184 ( .B1(n6992), .B2(n9706), .A(n6464), .ZN(P1_U3526) );
  INV_X1 U8185 ( .A(n6465), .ZN(n7629) );
  INV_X1 U8186 ( .A(n6466), .ZN(n6667) );
  NOR3_X1 U8187 ( .A1(n7629), .A2(n9966), .A3(n6667), .ZN(n6469) );
  INV_X1 U8188 ( .A(n6467), .ZN(n6468) );
  OAI21_X1 U8189 ( .B1(n6469), .B2(n6468), .A(n8098), .ZN(n6472) );
  AOI22_X1 U8190 ( .A1(n8086), .A2(n6470), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n8102), .ZN(n6471) );
  OAI211_X1 U8191 ( .C1(n6394), .C2(n8098), .A(n6472), .B(n6471), .ZN(P2_U3233) );
  INV_X1 U8192 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6499) );
  INV_X1 U8193 ( .A(n6473), .ZN(n6475) );
  XOR2_X1 U8194 ( .A(n6607), .B(n6601), .Z(n6477) );
  OAI211_X1 U8195 ( .C1(n6478), .C2(n6477), .A(n6602), .B(n9883), .ZN(n6498)
         );
  INV_X1 U8196 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6479) );
  MUX2_X1 U8197 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6479), .S(n6607), .Z(n6486)
         );
  NAND2_X1 U8198 ( .A1(n6480), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6484) );
  NAND2_X1 U8199 ( .A1(n6482), .A2(n6481), .ZN(n6483) );
  NAND2_X1 U8200 ( .A1(n6484), .A2(n6483), .ZN(n6485) );
  NAND2_X1 U8201 ( .A1(n6485), .A2(n6486), .ZN(n6600) );
  OAI21_X1 U8202 ( .B1(n6486), .B2(n6485), .A(n6600), .ZN(n6496) );
  INV_X1 U8203 ( .A(n9875), .ZN(n9511) );
  AND2_X1 U8204 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n6957) );
  INV_X1 U8205 ( .A(n6957), .ZN(n6487) );
  OAI21_X1 U8206 ( .B1(n9511), .B2(n6607), .A(n6487), .ZN(n6495) );
  NAND2_X1 U8207 ( .A1(n6492), .A2(n6490), .ZN(n6488) );
  XNOR2_X1 U8208 ( .A(n6607), .B(n7094), .ZN(n6489) );
  INV_X1 U8209 ( .A(n6489), .ZN(n6491) );
  NAND3_X1 U8210 ( .A1(n6492), .A2(n6491), .A3(n6490), .ZN(n6493) );
  AOI21_X1 U8211 ( .B1(n6609), .B2(n6493), .A(n9890), .ZN(n6494) );
  AOI211_X1 U8212 ( .C1(n9884), .C2(n6496), .A(n6495), .B(n6494), .ZN(n6497)
         );
  OAI211_X1 U8213 ( .C1(n6499), .C2(n9720), .A(n6498), .B(n6497), .ZN(P2_U3186) );
  OAI21_X1 U8214 ( .B1(n6501), .B2(n8574), .A(n6500), .ZN(n6930) );
  INV_X1 U8215 ( .A(n6930), .ZN(n6506) );
  XNOR2_X1 U8216 ( .A(n6502), .B(n8574), .ZN(n6503) );
  OAI22_X1 U8217 ( .A1(n6437), .A2(n9285), .B1(n6516), .B2(n9287), .ZN(n8316)
         );
  AOI21_X1 U8218 ( .B1(n6503), .B2(n9301), .A(n8316), .ZN(n6932) );
  INV_X1 U8219 ( .A(n9308), .ZN(n9373) );
  OAI211_X1 U8220 ( .C1(n6505), .C2(n7043), .A(n9373), .B(n6504), .ZN(n6928)
         );
  OAI211_X1 U8221 ( .C1(n6506), .C2(n9411), .A(n6932), .B(n6928), .ZN(n7045)
         );
  INV_X1 U8222 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6507) );
  OAI22_X1 U8223 ( .A1(n9406), .A2(n7043), .B1(n9403), .B2(n6507), .ZN(n6508)
         );
  AOI21_X1 U8224 ( .B1(n7045), .B2(n9403), .A(n6508), .ZN(n6509) );
  INV_X1 U8225 ( .A(n6509), .ZN(P1_U3525) );
  NAND2_X1 U8226 ( .A1(n6516), .A2(n6989), .ZN(n6510) );
  NAND2_X1 U8227 ( .A1(n8452), .A2(n8732), .ZN(n8658) );
  INV_X1 U8228 ( .A(n8732), .ZN(n8448) );
  NAND2_X1 U8229 ( .A1(n8448), .A2(n8450), .ZN(n8461) );
  AND2_X1 U8230 ( .A1(n8658), .A2(n8461), .ZN(n8578) );
  INV_X1 U8231 ( .A(n8578), .ZN(n6512) );
  OAI21_X1 U8232 ( .B1(n6513), .B2(n6512), .A(n6565), .ZN(n6514) );
  INV_X1 U8233 ( .A(n6514), .ZN(n6710) );
  XNOR2_X1 U8234 ( .A(n8446), .B(n8578), .ZN(n6517) );
  INV_X1 U8235 ( .A(n8731), .ZN(n8454) );
  OAI22_X1 U8236 ( .A1(n8454), .A2(n9287), .B1(n6516), .B2(n9285), .ZN(n6576)
         );
  AOI21_X1 U8237 ( .B1(n6517), .B2(n9301), .A(n6576), .ZN(n6703) );
  OAI211_X1 U8238 ( .C1(n6518), .C2(n8452), .A(n9373), .B(n6563), .ZN(n6704)
         );
  OAI211_X1 U8239 ( .C1(n6710), .C2(n9411), .A(n6703), .B(n6704), .ZN(n7056)
         );
  INV_X1 U8240 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6519) );
  OAI22_X1 U8241 ( .A1(n9406), .A2(n8452), .B1(n9403), .B2(n6519), .ZN(n6520)
         );
  AOI21_X1 U8242 ( .B1(n7056), .B2(n9403), .A(n6520), .ZN(n6521) );
  INV_X1 U8243 ( .A(n6521), .ZN(P1_U3527) );
  INV_X1 U8244 ( .A(n6522), .ZN(n6525) );
  OAI222_X1 U8245 ( .A1(n7398), .A2(n6523), .B1(n9500), .B2(n6525), .C1(
        P1_U3086), .C2(n8825), .ZN(P1_U3339) );
  INV_X1 U8246 ( .A(n9857), .ZN(n7907) );
  INV_X1 U8247 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6524) );
  OAI222_X1 U8248 ( .A1(n7907), .A2(P2_U3151), .B1(n8277), .B2(n6525), .C1(
        n6524), .C2(n8276), .ZN(P2_U3279) );
  NOR2_X1 U8249 ( .A1(n6526), .A2(n8748), .ZN(n8752) );
  INV_X1 U8250 ( .A(n8752), .ZN(n6527) );
  NOR2_X1 U8251 ( .A1(n7006), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6528) );
  AOI21_X1 U8252 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n7006), .A(n6528), .ZN(
        n6539) );
  INV_X1 U8253 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6769) );
  MUX2_X1 U8254 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n6769), .S(n8739), .Z(n8741)
         );
  AND2_X1 U8255 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n8751) );
  NAND2_X1 U8256 ( .A1(n8741), .A2(n8751), .ZN(n8740) );
  NAND2_X1 U8257 ( .A1(n8739), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6529) );
  NAND2_X1 U8258 ( .A1(n8740), .A2(n6529), .ZN(n8765) );
  INV_X1 U8259 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6684) );
  XNOR2_X1 U8260 ( .A(n8760), .B(n6684), .ZN(n8766) );
  NAND2_X1 U8261 ( .A1(n8765), .A2(n8766), .ZN(n8764) );
  NAND2_X1 U8262 ( .A1(n8760), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6530) );
  NAND2_X1 U8263 ( .A1(n8764), .A2(n6530), .ZN(n8779) );
  INV_X1 U8264 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6925) );
  XNOR2_X1 U8265 ( .A(n8777), .B(n6925), .ZN(n8780) );
  NAND2_X1 U8266 ( .A1(n8779), .A2(n8780), .ZN(n8778) );
  NAND2_X1 U8267 ( .A1(n8777), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6531) );
  NAND2_X1 U8268 ( .A1(n8778), .A2(n6531), .ZN(n8791) );
  XNOR2_X1 U8269 ( .A(n6543), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n8792) );
  NAND2_X1 U8270 ( .A1(n8791), .A2(n8792), .ZN(n8790) );
  INV_X1 U8271 ( .A(n6543), .ZN(n8789) );
  NAND2_X1 U8272 ( .A1(n8789), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6532) );
  NAND2_X1 U8273 ( .A1(n8790), .A2(n6532), .ZN(n8806) );
  INV_X1 U8274 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9051) );
  MUX2_X1 U8275 ( .A(n9051), .B(P1_REG2_REG_5__SCAN_IN), .S(n6544), .Z(n8807)
         );
  NAND2_X1 U8276 ( .A1(n8806), .A2(n8807), .ZN(n8805) );
  OR2_X1 U8277 ( .A1(n6544), .A2(n9051), .ZN(n6533) );
  NAND2_X1 U8278 ( .A1(n8805), .A2(n6533), .ZN(n9578) );
  NAND2_X1 U8279 ( .A1(n9587), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6534) );
  OAI21_X1 U8280 ( .B1(n9587), .B2(P1_REG2_REG_6__SCAN_IN), .A(n6534), .ZN(
        n9580) );
  INV_X1 U8281 ( .A(n9580), .ZN(n6535) );
  AOI21_X1 U8282 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n9587), .A(n9579), .ZN(
        n9537) );
  NAND2_X1 U8283 ( .A1(n9543), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6536) );
  OAI21_X1 U8284 ( .B1(n9543), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6536), .ZN(
        n9536) );
  NOR2_X1 U8285 ( .A1(n9537), .A2(n9536), .ZN(n9535) );
  AOI21_X1 U8286 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n9543), .A(n9535), .ZN(
        n9548) );
  NAND2_X1 U8287 ( .A1(n6549), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6537) );
  OAI21_X1 U8288 ( .B1(n6549), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6537), .ZN(
        n9549) );
  NOR2_X1 U8289 ( .A1(n9548), .A2(n9549), .ZN(n9547) );
  AOI21_X1 U8290 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n6549), .A(n9547), .ZN(
        n6538) );
  NAND2_X1 U8291 ( .A1(n6539), .A2(n6538), .ZN(n7000) );
  OAI21_X1 U8292 ( .B1(n6539), .B2(n6538), .A(n7000), .ZN(n6559) );
  INV_X1 U8293 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9704) );
  AOI22_X1 U8294 ( .A1(n7006), .A2(P1_REG1_REG_9__SCAN_IN), .B1(n9704), .B2(
        n6557), .ZN(n6551) );
  INV_X1 U8295 ( .A(n6544), .ZN(n8804) );
  XOR2_X1 U8296 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n8760), .Z(n8763) );
  INV_X1 U8297 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6542) );
  NAND3_X1 U8298 ( .A1(n8744), .A2(P1_IR_REG_0__SCAN_IN), .A3(
        P1_REG1_REG_0__SCAN_IN), .ZN(n8742) );
  OAI21_X1 U8299 ( .B1(n6542), .B2(n6541), .A(n8742), .ZN(n8762) );
  NAND2_X1 U8300 ( .A1(n8763), .A2(n8762), .ZN(n8761) );
  XNOR2_X1 U8301 ( .A(n8777), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n8771) );
  XOR2_X1 U8302 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6543), .Z(n8786) );
  NOR2_X1 U8303 ( .A1(n4302), .A2(n8786), .ZN(n8785) );
  AOI21_X1 U8304 ( .B1(n8789), .B2(P1_REG1_REG_4__SCAN_IN), .A(n8785), .ZN(
        n8799) );
  XOR2_X1 U8305 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6544), .Z(n8798) );
  NOR2_X1 U8306 ( .A1(n8799), .A2(n8798), .ZN(n8797) );
  AOI21_X1 U8307 ( .B1(n8804), .B2(P1_REG1_REG_5__SCAN_IN), .A(n8797), .ZN(
        n9584) );
  NAND2_X1 U8308 ( .A1(n9587), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6545) );
  OAI21_X1 U8309 ( .B1(n9587), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6545), .ZN(
        n9583) );
  NOR2_X1 U8310 ( .A1(n9584), .A2(n9583), .ZN(n9582) );
  INV_X1 U8311 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6546) );
  MUX2_X1 U8312 ( .A(n6546), .B(P1_REG1_REG_7__SCAN_IN), .S(n9543), .Z(n9539)
         );
  OR2_X1 U8313 ( .A1(n6549), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6548) );
  NAND2_X1 U8314 ( .A1(n6549), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6547) );
  NAND2_X1 U8315 ( .A1(n6548), .A2(n6547), .ZN(n9552) );
  AOI21_X1 U8316 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n6549), .A(n9551), .ZN(
        n6550) );
  NAND2_X1 U8317 ( .A1(n6551), .A2(n6550), .ZN(n7005) );
  OAI21_X1 U8318 ( .B1(n6551), .B2(n6550), .A(n7005), .ZN(n6553) );
  NAND2_X1 U8319 ( .A1(n6553), .A2(n9648), .ZN(n6556) );
  INV_X1 U8320 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6554) );
  NOR2_X1 U8321 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6554), .ZN(n7025) );
  AOI21_X1 U8322 ( .B1(n8835), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n7025), .ZN(
        n6555) );
  OAI211_X1 U8323 ( .C1(n9654), .C2(n6557), .A(n6556), .B(n6555), .ZN(n6558)
         );
  AOI21_X1 U8324 ( .B1(n9595), .B2(n6559), .A(n6558), .ZN(n6560) );
  INV_X1 U8325 ( .A(n6560), .ZN(P1_U3252) );
  INV_X1 U8326 ( .A(n8461), .ZN(n6561) );
  OR2_X1 U8327 ( .A1(n8454), .A2(n8458), .ZN(n8445) );
  NAND2_X1 U8328 ( .A1(n8458), .A2(n8454), .ZN(n8462) );
  AND2_X1 U8329 ( .A1(n8445), .A2(n8462), .ZN(n8579) );
  XNOR2_X1 U8330 ( .A(n6795), .B(n8579), .ZN(n6562) );
  OAI222_X1 U8331 ( .A1(n9287), .A2(n6939), .B1(n9285), .B2(n8448), .C1(n9283), 
        .C2(n6562), .ZN(n6874) );
  AOI211_X1 U8332 ( .C1(n8458), .C2(n6563), .A(n9308), .B(n4520), .ZN(n6878)
         );
  NOR2_X1 U8333 ( .A1(n6874), .A2(n6878), .ZN(n7053) );
  NAND2_X1 U8334 ( .A1(n8452), .A2(n8448), .ZN(n6564) );
  NAND2_X1 U8335 ( .A1(n6565), .A2(n6564), .ZN(n6567) );
  INV_X1 U8336 ( .A(n8579), .ZN(n6566) );
  NAND2_X1 U8337 ( .A1(n6567), .A2(n6566), .ZN(n6737) );
  OAI21_X1 U8338 ( .B1(n6567), .B2(n6566), .A(n6737), .ZN(n7051) );
  NAND2_X1 U8339 ( .A1(n9403), .A2(n9689), .ZN(n9388) );
  INV_X1 U8340 ( .A(n9388), .ZN(n6570) );
  INV_X1 U8341 ( .A(n8458), .ZN(n7048) );
  INV_X1 U8342 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6568) );
  OAI22_X1 U8343 ( .A1(n9406), .A2(n7048), .B1(n9403), .B2(n6568), .ZN(n6569)
         );
  AOI21_X1 U8344 ( .B1(n7051), .B2(n6570), .A(n6569), .ZN(n6571) );
  OAI21_X1 U8345 ( .B1(n7053), .B2(n9706), .A(n6571), .ZN(P1_U3528) );
  INV_X1 U8346 ( .A(n6572), .ZN(n6573) );
  NAND2_X1 U8347 ( .A1(n6573), .A2(n5693), .ZN(n6588) );
  OAI21_X1 U8348 ( .B1(n6573), .B2(n5693), .A(n6588), .ZN(n6574) );
  NOR2_X1 U8349 ( .A1(n6574), .A2(n6575), .ZN(n6591) );
  AOI21_X1 U8350 ( .B1(n6575), .B2(n6574), .A(n6591), .ZN(n6580) );
  NAND2_X1 U8351 ( .A1(n9568), .A2(n6576), .ZN(n6577) );
  NAND2_X1 U8352 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n8801) );
  OAI211_X1 U8353 ( .C1(n9577), .C2(n6705), .A(n6577), .B(n8801), .ZN(n6578)
         );
  AOI21_X1 U8354 ( .B1(n8450), .B2(n8422), .A(n6578), .ZN(n6579) );
  OAI21_X1 U8355 ( .B1(n6580), .B2(n8424), .A(n6579), .ZN(P1_U3227) );
  INV_X1 U8356 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6583) );
  OR2_X1 U8357 ( .A1(n6581), .A2(n9699), .ZN(n6582) );
  OAI21_X1 U8358 ( .B1(n9701), .B2(n6583), .A(n6582), .ZN(P1_U3453) );
  INV_X1 U8359 ( .A(n6584), .ZN(n6587) );
  OAI222_X1 U8360 ( .A1(n7398), .A2(n6585), .B1(n9500), .B2(n6587), .C1(
        P1_U3086), .C2(n8850), .ZN(P1_U3338) );
  INV_X1 U8361 ( .A(n9876), .ZN(n7864) );
  OAI222_X1 U8362 ( .A1(n7864), .A2(P2_U3151), .B1(n8277), .B2(n6587), .C1(
        n6586), .C2(n8276), .ZN(P2_U3278) );
  INV_X1 U8363 ( .A(n6588), .ZN(n6589) );
  NOR3_X1 U8364 ( .A1(n6591), .A2(n6590), .A3(n6589), .ZN(n6594) );
  INV_X1 U8365 ( .A(n6592), .ZN(n6593) );
  OAI21_X1 U8366 ( .B1(n6594), .B2(n6593), .A(n9573), .ZN(n6598) );
  NAND2_X1 U8367 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9588) );
  INV_X1 U8368 ( .A(n9588), .ZN(n6596) );
  INV_X1 U8369 ( .A(n8409), .ZN(n8430) );
  OAI22_X1 U8370 ( .A1(n8430), .A2(n8448), .B1(n6939), .B2(n8429), .ZN(n6595)
         );
  AOI211_X1 U8371 ( .C1(n8433), .C2(n6875), .A(n6596), .B(n6595), .ZN(n6597)
         );
  OAI211_X1 U8372 ( .C1(n7048), .C2(n9570), .A(n6598), .B(n6597), .ZN(P1_U3239) );
  NAND2_X1 U8373 ( .A1(n6607), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6599) );
  NAND2_X1 U8374 ( .A1(n6600), .A2(n6599), .ZN(n6848) );
  INV_X1 U8375 ( .A(n6847), .ZN(n6836) );
  XNOR2_X1 U8376 ( .A(n6848), .B(n6836), .ZN(n6850) );
  XOR2_X1 U8377 ( .A(n6850), .B(P2_REG1_REG_5__SCAN_IN), .Z(n6616) );
  INV_X1 U8378 ( .A(n6607), .ZN(n6604) );
  INV_X1 U8379 ( .A(n6601), .ZN(n6603) );
  OAI21_X1 U8380 ( .B1(n6604), .B2(n6603), .A(n6602), .ZN(n6606) );
  XOR2_X1 U8381 ( .A(n6847), .B(n6833), .Z(n6605) );
  OAI211_X1 U8382 ( .C1(n6606), .C2(n6605), .A(n6834), .B(n9883), .ZN(n6615)
         );
  INV_X1 U8383 ( .A(n9890), .ZN(n9754) );
  NAND2_X1 U8384 ( .A1(n6607), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6608) );
  XNOR2_X1 U8385 ( .A(n6839), .B(n6610), .ZN(n6613) );
  INV_X1 U8386 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n9093) );
  AND2_X1 U8387 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7038) );
  AOI21_X1 U8388 ( .B1(n9875), .B2(n6836), .A(n7038), .ZN(n6611) );
  OAI21_X1 U8389 ( .B1(n9720), .B2(n9093), .A(n6611), .ZN(n6612) );
  AOI21_X1 U8390 ( .B1(n9754), .B2(n6613), .A(n6612), .ZN(n6614) );
  OAI211_X1 U8391 ( .C1(n6616), .C2(n9732), .A(n6615), .B(n6614), .ZN(P2_U3187) );
  NAND2_X1 U8392 ( .A1(n5413), .A2(n7661), .ZN(n6617) );
  NAND2_X1 U8393 ( .A1(n6618), .A2(n6617), .ZN(n8175) );
  INV_X1 U8394 ( .A(n8175), .ZN(n6626) );
  INV_X1 U8395 ( .A(n7155), .ZN(n8158) );
  NAND2_X1 U8396 ( .A1(n8175), .A2(n8158), .ZN(n6623) );
  AOI22_X1 U8397 ( .A1(n7834), .A2(n8092), .B1(n8161), .B2(n7832), .ZN(n6622)
         );
  XNOR2_X1 U8398 ( .A(n5413), .B(n6619), .ZN(n6620) );
  NAND2_X1 U8399 ( .A1(n6620), .A2(n8167), .ZN(n6621) );
  AND3_X1 U8400 ( .A1(n6623), .A2(n6622), .A3(n6621), .ZN(n8177) );
  MUX2_X1 U8401 ( .A(n8177), .B(n7835), .S(n9907), .Z(n6625) );
  AOI22_X1 U8402 ( .A1(n8086), .A2(n8174), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8102), .ZN(n6624) );
  OAI211_X1 U8403 ( .C1(n6626), .C2(n7306), .A(n6625), .B(n6624), .ZN(P2_U3232) );
  INV_X1 U8404 ( .A(n6627), .ZN(n6634) );
  INV_X1 U8405 ( .A(n6628), .ZN(n6660) );
  NAND3_X1 U8406 ( .A1(n6631), .A2(n6630), .A3(n6629), .ZN(n6632) );
  AOI21_X1 U8407 ( .B1(n6639), .B2(n6660), .A(n6632), .ZN(n6633) );
  OAI21_X1 U8408 ( .B1(n6635), .B2(n6634), .A(n6633), .ZN(n6636) );
  NAND2_X1 U8409 ( .A1(n6636), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6641) );
  NAND2_X1 U8410 ( .A1(n6637), .A2(n6667), .ZN(n7813) );
  INV_X1 U8411 ( .A(n7813), .ZN(n6638) );
  NAND2_X1 U8412 ( .A1(n6639), .A2(n6638), .ZN(n6640) );
  NAND2_X1 U8413 ( .A1(n7804), .A2(n6643), .ZN(n6644) );
  AND2_X1 U8414 ( .A1(n6645), .A2(n6644), .ZN(n6646) );
  INV_X1 U8415 ( .A(n6648), .ZN(n6647) );
  NAND2_X1 U8416 ( .A1(n6647), .A2(n8165), .ZN(n6654) );
  NAND2_X1 U8417 ( .A1(n6648), .A2(n4867), .ZN(n6649) );
  NAND2_X1 U8418 ( .A1(n6654), .A2(n6649), .ZN(n6719) );
  INV_X1 U8419 ( .A(n6719), .ZN(n6653) );
  NAND2_X1 U8420 ( .A1(n6655), .A2(n6713), .ZN(n6651) );
  AND2_X1 U8421 ( .A1(n7661), .A2(n6651), .ZN(n6720) );
  INV_X1 U8422 ( .A(n6720), .ZN(n6652) );
  NAND2_X1 U8423 ( .A1(n6653), .A2(n6652), .ZN(n6717) );
  NAND2_X1 U8424 ( .A1(n6717), .A2(n6654), .ZN(n6729) );
  XNOR2_X1 U8425 ( .A(n6650), .B(n8171), .ZN(n6656) );
  XNOR2_X1 U8426 ( .A(n6656), .B(n4891), .ZN(n6730) );
  NAND2_X1 U8427 ( .A1(n6729), .A2(n6730), .ZN(n6728) );
  INV_X1 U8428 ( .A(n6656), .ZN(n6657) );
  NAND2_X1 U8429 ( .A1(n6657), .A2(n4891), .ZN(n6658) );
  AND2_X1 U8430 ( .A1(n6728), .A2(n6658), .ZN(n6664) );
  INV_X1 U8431 ( .A(n7063), .ZN(n9912) );
  XNOR2_X1 U8432 ( .A(n7439), .B(n9912), .ZN(n6946) );
  XNOR2_X1 U8433 ( .A(n6946), .B(n6955), .ZN(n6663) );
  OR2_X1 U8434 ( .A1(n6665), .A2(n6659), .ZN(n6662) );
  NAND2_X1 U8435 ( .A1(n6668), .A2(n6660), .ZN(n6661) );
  OAI211_X1 U8436 ( .C1(n6664), .C2(n6663), .A(n6948), .B(n7591), .ZN(n6674)
         );
  OR2_X1 U8437 ( .A1(n6665), .A2(n9948), .ZN(n6666) );
  NAND2_X1 U8438 ( .A1(n6668), .A2(n6667), .ZN(n6670) );
  OAI22_X1 U8439 ( .A1(n4891), .A2(n7575), .B1(n7598), .B2(n7144), .ZN(n6671)
         );
  AOI211_X1 U8440 ( .C1(n7063), .C2(n7587), .A(n6672), .B(n6671), .ZN(n6673)
         );
  OAI211_X1 U8441 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n7558), .A(n6674), .B(
        n6673), .ZN(P2_U3158) );
  INV_X1 U8442 ( .A(n9514), .ZN(n7911) );
  INV_X1 U8443 ( .A(n6675), .ZN(n6711) );
  OAI222_X1 U8444 ( .A1(P2_U3151), .A2(n7911), .B1(n8277), .B2(n6711), .C1(
        n6676), .C2(n8276), .ZN(P2_U3277) );
  INV_X1 U8445 ( .A(n6677), .ZN(n6692) );
  NAND3_X1 U8446 ( .A1(n6680), .A2(n6679), .A3(n6678), .ZN(n6683) );
  INV_X1 U8447 ( .A(n6701), .ZN(n6681) );
  NAND2_X1 U8448 ( .A1(n9306), .A2(n6681), .ZN(n9320) );
  NAND2_X1 U8449 ( .A1(n6682), .A2(n9306), .ZN(n6691) );
  INV_X1 U8450 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n8757) );
  OAI22_X1 U8451 ( .A1(n9306), .A2(n6684), .B1(n8757), .B2(n9257), .ZN(n6688)
         );
  INV_X1 U8452 ( .A(n6685), .ZN(n6686) );
  NOR2_X1 U8453 ( .A1(n9315), .A2(n6994), .ZN(n6687) );
  AOI211_X1 U8454 ( .C1(n6689), .C2(n9317), .A(n6688), .B(n6687), .ZN(n6690)
         );
  OAI211_X1 U8455 ( .C1(n6692), .C2(n9320), .A(n6691), .B(n6690), .ZN(P1_U3291) );
  AOI22_X1 U8456 ( .A1(n8409), .A2(n8731), .B1(n8407), .B2(n8729), .ZN(n6693)
         );
  NAND2_X1 U8457 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n9544) );
  OAI211_X1 U8458 ( .C1(n6694), .C2(n9577), .A(n6693), .B(n9544), .ZN(n6699)
         );
  AOI211_X1 U8459 ( .C1(n6697), .C2(n6696), .A(n8424), .B(n6695), .ZN(n6698)
         );
  AOI211_X1 U8460 ( .C1(n9676), .C2(n8422), .A(n6699), .B(n6698), .ZN(n6700)
         );
  INV_X1 U8461 ( .A(n6700), .ZN(P1_U3213) );
  NAND2_X1 U8462 ( .A1(n9305), .A2(n6701), .ZN(n6702) );
  MUX2_X1 U8463 ( .A(n9051), .B(n6703), .S(n9306), .Z(n6709) );
  INV_X1 U8464 ( .A(n6704), .ZN(n6707) );
  OAI22_X1 U8465 ( .A1(n9315), .A2(n8452), .B1(n6705), .B2(n9257), .ZN(n6706)
         );
  AOI21_X1 U8466 ( .B1(n6707), .B2(n9317), .A(n6706), .ZN(n6708) );
  OAI211_X1 U8467 ( .C1(n6710), .C2(n9294), .A(n6709), .B(n6708), .ZN(P1_U3288) );
  OAI222_X1 U8468 ( .A1(n7398), .A2(n6712), .B1(n9653), .B2(P1_U3086), .C1(
        n9500), .C2(n6711), .ZN(P1_U3337) );
  NOR2_X1 U8469 ( .A1(n7600), .A2(P2_U3151), .ZN(n6735) );
  INV_X1 U8470 ( .A(n7587), .ZN(n7603) );
  OAI22_X1 U8471 ( .A1(n7603), .A2(n6713), .B1(n7589), .B2(n7629), .ZN(n6714)
         );
  AOI21_X1 U8472 ( .B1(n7573), .B2(n4867), .A(n6714), .ZN(n6715) );
  OAI21_X1 U8473 ( .B1(n6735), .B2(n6716), .A(n6715), .ZN(P2_U3172) );
  INV_X1 U8474 ( .A(n6717), .ZN(n6718) );
  AOI21_X1 U8475 ( .B1(n6720), .B2(n6719), .A(n6718), .ZN(n6727) );
  OAI22_X1 U8476 ( .A1(n7603), .A2(n6722), .B1(n6721), .B2(n7575), .ZN(n6725)
         );
  NOR2_X1 U8477 ( .A1(n6735), .A2(n6723), .ZN(n6724) );
  AOI211_X1 U8478 ( .C1(n7573), .C2(n7832), .A(n6725), .B(n6724), .ZN(n6726)
         );
  OAI21_X1 U8479 ( .B1(n7589), .B2(n6727), .A(n6726), .ZN(P2_U3162) );
  OAI21_X1 U8480 ( .B1(n6730), .B2(n6729), .A(n6728), .ZN(n6731) );
  NAND2_X1 U8481 ( .A1(n6731), .A2(n7591), .ZN(n6734) );
  OAI22_X1 U8482 ( .A1(n7603), .A2(n8171), .B1(n8165), .B2(n7575), .ZN(n6732)
         );
  AOI21_X1 U8483 ( .B1(n7573), .B2(n8162), .A(n6732), .ZN(n6733) );
  OAI211_X1 U8484 ( .C1(n6735), .C2(n4886), .A(n6734), .B(n6733), .ZN(P2_U3177) );
  OR2_X1 U8485 ( .A1(n8458), .A2(n8731), .ZN(n6736) );
  NAND2_X1 U8486 ( .A1(n6737), .A2(n6736), .ZN(n6882) );
  NAND2_X1 U8487 ( .A1(n9676), .A2(n6939), .ZN(n8466) );
  INV_X1 U8488 ( .A(n8466), .ZN(n6738) );
  NAND2_X1 U8489 ( .A1(n6882), .A2(n6885), .ZN(n6884) );
  OR2_X1 U8490 ( .A1(n9676), .A2(n8730), .ZN(n6739) );
  NAND2_X1 U8491 ( .A1(n6884), .A2(n6739), .ZN(n6740) );
  INV_X1 U8492 ( .A(n8729), .ZN(n7023) );
  OR2_X1 U8493 ( .A1(n6942), .A2(n7023), .ZN(n8469) );
  NAND2_X1 U8494 ( .A1(n6942), .A2(n7023), .ZN(n8475) );
  NAND2_X1 U8495 ( .A1(n8469), .A2(n8475), .ZN(n6741) );
  NAND2_X1 U8496 ( .A1(n6740), .A2(n6741), .ZN(n6787) );
  OAI21_X1 U8497 ( .B1(n6740), .B2(n6741), .A(n6787), .ZN(n6829) );
  INV_X1 U8498 ( .A(n6829), .ZN(n6755) );
  INV_X1 U8499 ( .A(n6741), .ZN(n6746) );
  INV_X1 U8500 ( .A(n8445), .ZN(n6742) );
  OR2_X1 U8501 ( .A1(n6795), .A2(n6742), .ZN(n6886) );
  NAND2_X1 U8502 ( .A1(n6886), .A2(n8462), .ZN(n6744) );
  INV_X1 U8503 ( .A(n6885), .ZN(n6743) );
  NAND2_X1 U8504 ( .A1(n6744), .A2(n6743), .ZN(n6888) );
  NAND2_X1 U8505 ( .A1(n6888), .A2(n8466), .ZN(n6745) );
  NAND2_X1 U8506 ( .A1(n6745), .A2(n6746), .ZN(n6906) );
  OAI21_X1 U8507 ( .B1(n6746), .B2(n6745), .A(n6906), .ZN(n6748) );
  INV_X1 U8508 ( .A(n8728), .ZN(n6938) );
  OAI22_X1 U8509 ( .A1(n6939), .A2(n9285), .B1(n6938), .B2(n9287), .ZN(n6747)
         );
  AOI21_X1 U8510 ( .B1(n6748), .B2(n9301), .A(n6747), .ZN(n6749) );
  OAI21_X1 U8511 ( .B1(n6755), .B2(n9305), .A(n6749), .ZN(n6827) );
  NAND2_X1 U8512 ( .A1(n6827), .A2(n9306), .ZN(n6754) );
  AOI211_X1 U8513 ( .C1(n6942), .C2(n6896), .A(n9308), .B(n6915), .ZN(n6828)
         );
  INV_X1 U8514 ( .A(n6942), .ZN(n6751) );
  AOI22_X1 U8515 ( .A1(n4251), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n4820), .B2(
        n9312), .ZN(n6750) );
  OAI21_X1 U8516 ( .B1(n6751), .B2(n9315), .A(n6750), .ZN(n6752) );
  AOI21_X1 U8517 ( .B1(n6828), .B2(n9317), .A(n6752), .ZN(n6753) );
  OAI211_X1 U8518 ( .C1(n6755), .C2(n9320), .A(n6754), .B(n6753), .ZN(P1_U3285) );
  INV_X1 U8519 ( .A(n6756), .ZN(n6757) );
  NAND2_X1 U8520 ( .A1(n8571), .A2(n6757), .ZN(n6758) );
  NAND2_X1 U8521 ( .A1(n6759), .A2(n6758), .ZN(n9671) );
  NAND2_X1 U8522 ( .A1(n9671), .A2(n6979), .ZN(n6768) );
  OAI21_X1 U8523 ( .B1(n6761), .B2(n8571), .A(n6760), .ZN(n6766) );
  NAND2_X1 U8524 ( .A1(n6762), .A2(n9224), .ZN(n6764) );
  NAND2_X1 U8525 ( .A1(n8735), .A2(n9222), .ZN(n6763) );
  NAND2_X1 U8526 ( .A1(n6764), .A2(n6763), .ZN(n6765) );
  AOI21_X1 U8527 ( .B1(n6766), .B2(n9301), .A(n6765), .ZN(n6767) );
  AND2_X1 U8528 ( .A1(n6768), .A2(n6767), .ZN(n9673) );
  NOR2_X1 U8529 ( .A1(n9306), .A2(n6769), .ZN(n6773) );
  AOI21_X1 U8530 ( .B1(n6774), .B2(n6782), .A(n9308), .ZN(n6770) );
  NAND2_X1 U8531 ( .A1(n6771), .A2(n6770), .ZN(n9668) );
  INV_X1 U8532 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n8736) );
  OAI22_X1 U8533 ( .A1(n8982), .A2(n9668), .B1(n8736), .B2(n9257), .ZN(n6772)
         );
  AOI211_X1 U8534 ( .C1(n9005), .C2(n6774), .A(n6773), .B(n6772), .ZN(n6776)
         );
  INV_X1 U8535 ( .A(n9320), .ZN(n6986) );
  NAND2_X1 U8536 ( .A1(n9671), .A2(n6986), .ZN(n6775) );
  OAI211_X1 U8537 ( .C1(n4251), .C2(n9673), .A(n6776), .B(n6775), .ZN(P1_U3292) );
  INV_X1 U8538 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6785) );
  INV_X1 U8539 ( .A(n6777), .ZN(n6780) );
  AOI21_X1 U8540 ( .B1(n9312), .B2(P1_REG3_REG_0__SCAN_IN), .A(n6778), .ZN(
        n6779) );
  OAI21_X1 U8541 ( .B1(n8572), .B2(n6780), .A(n6779), .ZN(n6781) );
  NAND2_X1 U8542 ( .A1(n6781), .A2(n9306), .ZN(n6784) );
  NOR2_X1 U8543 ( .A1(n8982), .A2(n9308), .ZN(n9229) );
  OAI21_X1 U8544 ( .B1(n9229), .B2(n9005), .A(n6782), .ZN(n6783) );
  OAI211_X1 U8545 ( .C1(n6785), .C2(n9306), .A(n6784), .B(n6783), .ZN(P1_U3293) );
  OR2_X1 U8546 ( .A1(n6942), .A2(n8729), .ZN(n6786) );
  NAND2_X1 U8547 ( .A1(n6787), .A2(n6786), .ZN(n6914) );
  OR2_X1 U8548 ( .A1(n6919), .A2(n6938), .ZN(n8484) );
  INV_X1 U8549 ( .A(n8484), .ZN(n6788) );
  AND2_X1 U8550 ( .A1(n6919), .A2(n6938), .ZN(n8485) );
  NAND2_X1 U8551 ( .A1(n6914), .A2(n6913), .ZN(n6912) );
  OR2_X1 U8552 ( .A1(n6919), .A2(n8728), .ZN(n6789) );
  NAND2_X1 U8553 ( .A1(n6912), .A2(n6789), .ZN(n6790) );
  INV_X1 U8554 ( .A(n8727), .ZN(n7162) );
  OR2_X1 U8555 ( .A1(n6970), .A2(n7162), .ZN(n8487) );
  NAND2_X1 U8556 ( .A1(n6970), .A2(n7162), .ZN(n8490) );
  NAND2_X1 U8557 ( .A1(n8487), .A2(n8490), .ZN(n8584) );
  NAND2_X1 U8558 ( .A1(n6790), .A2(n8584), .ZN(n6972) );
  OAI21_X1 U8559 ( .B1(n6790), .B2(n8584), .A(n6972), .ZN(n6962) );
  INV_X1 U8560 ( .A(n6962), .ZN(n7075) );
  AND2_X1 U8561 ( .A1(n8475), .A2(n8466), .ZN(n8470) );
  INV_X1 U8562 ( .A(n8470), .ZN(n6791) );
  AND2_X1 U8563 ( .A1(n6791), .A2(n8469), .ZN(n6904) );
  NAND2_X1 U8564 ( .A1(n6904), .A2(n8484), .ZN(n6793) );
  INV_X1 U8565 ( .A(n8485), .ZN(n6792) );
  NAND2_X1 U8566 ( .A1(n6793), .A2(n6792), .ZN(n8583) );
  INV_X1 U8567 ( .A(n8583), .ZN(n6794) );
  NAND3_X1 U8568 ( .A1(n6795), .A2(n6794), .A3(n8462), .ZN(n6798) );
  AND2_X1 U8569 ( .A1(n8484), .A2(n8469), .ZN(n8474) );
  INV_X1 U8570 ( .A(n8474), .ZN(n8582) );
  INV_X1 U8571 ( .A(n8463), .ZN(n8577) );
  NAND2_X1 U8572 ( .A1(n8577), .A2(n8445), .ZN(n6796) );
  NOR2_X1 U8573 ( .A1(n8582), .A2(n6796), .ZN(n6797) );
  OR2_X1 U8574 ( .A1(n6797), .A2(n8583), .ZN(n8660) );
  NAND2_X1 U8575 ( .A1(n6798), .A2(n8660), .ZN(n8662) );
  NAND2_X1 U8576 ( .A1(n8662), .A2(n8584), .ZN(n6799) );
  NAND2_X1 U8577 ( .A1(n7117), .A2(n6799), .ZN(n6802) );
  NAND2_X1 U8578 ( .A1(n8728), .A2(n9224), .ZN(n6801) );
  NAND2_X1 U8579 ( .A1(n8726), .A2(n9222), .ZN(n6800) );
  NAND2_X1 U8580 ( .A1(n6801), .A2(n6800), .ZN(n9567) );
  AOI21_X1 U8581 ( .B1(n6802), .B2(n9301), .A(n9567), .ZN(n6969) );
  INV_X1 U8582 ( .A(n6803), .ZN(n6916) );
  INV_X1 U8583 ( .A(n6970), .ZN(n9571) );
  OAI211_X1 U8584 ( .C1(n6916), .C2(n9571), .A(n9373), .B(n6980), .ZN(n6964)
         );
  NAND2_X1 U8585 ( .A1(n6969), .A2(n6964), .ZN(n7073) );
  INV_X1 U8586 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6804) );
  OAI22_X1 U8587 ( .A1(n9571), .A2(n9406), .B1(n9403), .B2(n6804), .ZN(n6805)
         );
  AOI21_X1 U8588 ( .B1(n7073), .B2(n9403), .A(n6805), .ZN(n6806) );
  OAI21_X1 U8589 ( .B1(n7075), .B2(n9388), .A(n6806), .ZN(P1_U3532) );
  INV_X1 U8590 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n9992) );
  INV_X1 U8591 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9660) );
  NOR2_X1 U8592 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n6807) );
  AOI21_X1 U8593 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n6807), .ZN(n9995) );
  NOR2_X1 U8594 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n6808) );
  AOI21_X1 U8595 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n6808), .ZN(n9998) );
  NOR2_X1 U8596 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n6809) );
  AOI21_X1 U8597 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n6809), .ZN(n10001) );
  NOR2_X1 U8598 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n6810) );
  AOI21_X1 U8599 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n6810), .ZN(n10004) );
  NOR2_X1 U8600 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(P2_ADDR_REG_13__SCAN_IN), 
        .ZN(n6811) );
  AOI21_X1 U8601 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n6811), .ZN(n10007) );
  NOR2_X1 U8602 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(P2_ADDR_REG_12__SCAN_IN), 
        .ZN(n6812) );
  AOI21_X1 U8603 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n6812), .ZN(n10010) );
  NOR2_X1 U8604 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n6813) );
  AOI21_X1 U8605 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n6813), .ZN(n10013) );
  NOR2_X1 U8606 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n6814) );
  AOI21_X1 U8607 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n6814), .ZN(n10016) );
  NOR2_X1 U8608 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n6815) );
  AOI21_X1 U8609 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n6815), .ZN(n10025) );
  NOR2_X1 U8610 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n6816) );
  AOI21_X1 U8611 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n6816), .ZN(n10031) );
  NOR2_X1 U8612 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n6817) );
  AOI21_X1 U8613 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n6817), .ZN(n10028) );
  NOR2_X1 U8614 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(P2_ADDR_REG_6__SCAN_IN), 
        .ZN(n6818) );
  AOI21_X1 U8615 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n6818), .ZN(n10019) );
  NOR2_X1 U8616 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n6819) );
  AOI21_X1 U8617 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n6819), .ZN(n10022) );
  AND2_X1 U8618 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n6820) );
  NOR2_X1 U8619 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n6820), .ZN(n9984) );
  INV_X1 U8620 ( .A(n9984), .ZN(n9985) );
  INV_X1 U8621 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9987) );
  NAND3_X1 U8622 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n9986) );
  NAND2_X1 U8623 ( .A1(n9987), .A2(n9986), .ZN(n9983) );
  NAND2_X1 U8624 ( .A1(n9985), .A2(n9983), .ZN(n10034) );
  NAND2_X1 U8625 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n6821) );
  OAI21_X1 U8626 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n6821), .ZN(n10033) );
  NOR2_X1 U8627 ( .A1(n10034), .A2(n10033), .ZN(n10032) );
  AOI21_X1 U8628 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n10032), .ZN(n10037) );
  NAND2_X1 U8629 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n6822) );
  OAI21_X1 U8630 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n6822), .ZN(n10036) );
  NOR2_X1 U8631 ( .A1(n10037), .A2(n10036), .ZN(n10035) );
  AOI21_X1 U8632 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n10035), .ZN(n10040) );
  NOR2_X1 U8633 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n6823) );
  AOI21_X1 U8634 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n6823), .ZN(n10039) );
  NAND2_X1 U8635 ( .A1(n10040), .A2(n10039), .ZN(n10038) );
  OAI21_X1 U8636 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10038), .ZN(n10021) );
  NAND2_X1 U8637 ( .A1(n10022), .A2(n10021), .ZN(n10020) );
  OAI21_X1 U8638 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10020), .ZN(n10018) );
  NAND2_X1 U8639 ( .A1(n10019), .A2(n10018), .ZN(n10017) );
  OAI21_X1 U8640 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n10017), .ZN(n10027) );
  NAND2_X1 U8641 ( .A1(n10028), .A2(n10027), .ZN(n10026) );
  OAI21_X1 U8642 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10026), .ZN(n10030) );
  NAND2_X1 U8643 ( .A1(n10031), .A2(n10030), .ZN(n10029) );
  OAI21_X1 U8644 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10029), .ZN(n10024) );
  NAND2_X1 U8645 ( .A1(n10025), .A2(n10024), .ZN(n10023) );
  OAI21_X1 U8646 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10023), .ZN(n10015) );
  NAND2_X1 U8647 ( .A1(n10016), .A2(n10015), .ZN(n10014) );
  OAI21_X1 U8648 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10014), .ZN(n10012) );
  NAND2_X1 U8649 ( .A1(n10013), .A2(n10012), .ZN(n10011) );
  OAI21_X1 U8650 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10011), .ZN(n10009) );
  NAND2_X1 U8651 ( .A1(n10010), .A2(n10009), .ZN(n10008) );
  OAI21_X1 U8652 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n10008), .ZN(n10006) );
  NAND2_X1 U8653 ( .A1(n10007), .A2(n10006), .ZN(n10005) );
  OAI21_X1 U8654 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n10005), .ZN(n10003) );
  NAND2_X1 U8655 ( .A1(n10004), .A2(n10003), .ZN(n10002) );
  OAI21_X1 U8656 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10002), .ZN(n10000) );
  NAND2_X1 U8657 ( .A1(n10001), .A2(n10000), .ZN(n9999) );
  OAI21_X1 U8658 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9999), .ZN(n9997) );
  NAND2_X1 U8659 ( .A1(n9998), .A2(n9997), .ZN(n9996) );
  OAI21_X1 U8660 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9996), .ZN(n9994) );
  NAND2_X1 U8661 ( .A1(n9995), .A2(n9994), .ZN(n9993) );
  OAI21_X1 U8662 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9993), .ZN(n6824) );
  OR2_X1 U8663 ( .A1(n9660), .A2(n6824), .ZN(n9991) );
  NAND2_X1 U8664 ( .A1(n9992), .A2(n9991), .ZN(n9988) );
  NAND2_X1 U8665 ( .A1(n9660), .A2(n6824), .ZN(n9990) );
  NAND2_X1 U8666 ( .A1(n9988), .A2(n9990), .ZN(n6826) );
  XNOR2_X1 U8667 ( .A(n4528), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n6825) );
  XNOR2_X1 U8668 ( .A(n6826), .B(n6825), .ZN(ADD_1068_U4) );
  AOI211_X1 U8669 ( .C1(n9695), .C2(n6829), .A(n6828), .B(n6827), .ZN(n6864)
         );
  INV_X1 U8670 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6830) );
  NOR2_X1 U8671 ( .A1(n9403), .A2(n6830), .ZN(n6831) );
  AOI21_X1 U8672 ( .B1(n9360), .B2(n6942), .A(n6831), .ZN(n6832) );
  OAI21_X1 U8673 ( .B1(n6864), .B2(n9706), .A(n6832), .ZN(P1_U3530) );
  XNOR2_X1 U8674 ( .A(n7245), .B(n7253), .ZN(n6838) );
  INV_X1 U8675 ( .A(n6833), .ZN(n6835) );
  AOI21_X1 U8676 ( .B1(n6838), .B2(n6837), .A(n7246), .ZN(n6860) );
  MUX2_X1 U8677 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n7133), .S(n7253), .Z(n6843)
         );
  NAND2_X1 U8678 ( .A1(n6840), .A2(n6847), .ZN(n6841) );
  NAND2_X1 U8679 ( .A1(n6842), .A2(n6843), .ZN(n7242) );
  OAI21_X1 U8680 ( .B1(n6843), .B2(n6842), .A(n7242), .ZN(n6858) );
  INV_X1 U8681 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n6846) );
  INV_X1 U8682 ( .A(n7253), .ZN(n7248) );
  INV_X1 U8683 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6844) );
  NOR2_X1 U8684 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6844), .ZN(n7107) );
  AOI21_X1 U8685 ( .B1(n9875), .B2(n7248), .A(n7107), .ZN(n6845) );
  OAI21_X1 U8686 ( .B1(n9720), .B2(n6846), .A(n6845), .ZN(n6857) );
  AND2_X1 U8687 ( .A1(n6848), .A2(n6847), .ZN(n6849) );
  AOI21_X1 U8688 ( .B1(n6850), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6849), .ZN(
        n6854) );
  INV_X1 U8689 ( .A(n6854), .ZN(n6852) );
  INV_X1 U8690 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9974) );
  MUX2_X1 U8691 ( .A(n9974), .B(P2_REG1_REG_6__SCAN_IN), .S(n7253), .Z(n6853)
         );
  INV_X1 U8692 ( .A(n6853), .ZN(n6851) );
  NAND2_X1 U8693 ( .A1(n6852), .A2(n6851), .ZN(n7255) );
  NAND2_X1 U8694 ( .A1(n6854), .A2(n6853), .ZN(n6855) );
  AOI21_X1 U8695 ( .B1(n7255), .B2(n6855), .A(n9732), .ZN(n6856) );
  AOI211_X1 U8696 ( .C1(n9754), .C2(n6858), .A(n6857), .B(n6856), .ZN(n6859)
         );
  OAI21_X1 U8697 ( .B1(n6860), .B2(n9508), .A(n6859), .ZN(P2_U3188) );
  INV_X1 U8698 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n6861) );
  NOR2_X1 U8699 ( .A1(n9479), .A2(n6861), .ZN(n6862) );
  AOI21_X1 U8700 ( .B1(n9453), .B2(n6942), .A(n6862), .ZN(n6863) );
  OAI21_X1 U8701 ( .B1(n6864), .B2(n9699), .A(n6863), .ZN(P1_U3477) );
  INV_X1 U8702 ( .A(n6865), .ZN(n6873) );
  NAND2_X1 U8703 ( .A1(n6866), .A2(n9317), .ZN(n6869) );
  AOI22_X1 U8704 ( .A1(n4251), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n6867), .B2(
        n9312), .ZN(n6868) );
  OAI211_X1 U8705 ( .C1(n6989), .C2(n9315), .A(n6869), .B(n6868), .ZN(n6870)
         );
  AOI21_X1 U8706 ( .B1(n4648), .B2(n6871), .A(n6870), .ZN(n6872) );
  OAI21_X1 U8707 ( .B1(n6873), .B2(n4251), .A(n6872), .ZN(P1_U3289) );
  INV_X1 U8708 ( .A(n7051), .ZN(n6881) );
  NAND2_X1 U8709 ( .A1(n6874), .A2(n9306), .ZN(n6880) );
  AOI22_X1 U8710 ( .A1(n4251), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n6875), .B2(
        n9312), .ZN(n6876) );
  OAI21_X1 U8711 ( .B1(n7048), .B2(n9315), .A(n6876), .ZN(n6877) );
  AOI21_X1 U8712 ( .B1(n6878), .B2(n9317), .A(n6877), .ZN(n6879) );
  OAI211_X1 U8713 ( .C1(n6881), .C2(n9294), .A(n6880), .B(n6879), .ZN(P1_U3287) );
  OR2_X1 U8714 ( .A1(n6882), .A2(n6885), .ZN(n6883) );
  NAND2_X1 U8715 ( .A1(n6884), .A2(n6883), .ZN(n9680) );
  NAND2_X1 U8716 ( .A1(n9680), .A2(n6979), .ZN(n6894) );
  NAND3_X1 U8717 ( .A1(n6886), .A2(n8462), .A3(n6885), .ZN(n6887) );
  NAND2_X1 U8718 ( .A1(n6888), .A2(n6887), .ZN(n6892) );
  NAND2_X1 U8719 ( .A1(n8731), .A2(n9224), .ZN(n6890) );
  NAND2_X1 U8720 ( .A1(n8729), .A2(n9222), .ZN(n6889) );
  NAND2_X1 U8721 ( .A1(n6890), .A2(n6889), .ZN(n6891) );
  AOI21_X1 U8722 ( .B1(n6892), .B2(n9301), .A(n6891), .ZN(n6893) );
  AND2_X1 U8723 ( .A1(n6894), .A2(n6893), .ZN(n9682) );
  AOI21_X1 U8724 ( .B1(n6895), .B2(n9676), .A(n9308), .ZN(n6897) );
  NAND2_X1 U8725 ( .A1(n6897), .A2(n6896), .ZN(n9678) );
  AOI22_X1 U8726 ( .A1(n4251), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n6898), .B2(
        n9312), .ZN(n6900) );
  NAND2_X1 U8727 ( .A1(n9005), .A2(n9676), .ZN(n6899) );
  OAI211_X1 U8728 ( .C1(n9678), .C2(n8982), .A(n6900), .B(n6899), .ZN(n6901)
         );
  AOI21_X1 U8729 ( .B1(n9680), .B2(n6986), .A(n6901), .ZN(n6902) );
  OAI21_X1 U8730 ( .B1(n9682), .B2(n4251), .A(n6902), .ZN(P1_U3286) );
  NAND2_X1 U8731 ( .A1(n7833), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6903) );
  OAI21_X1 U8732 ( .B1(n7655), .B2(n7833), .A(n6903), .ZN(P2_U3520) );
  INV_X1 U8733 ( .A(n6904), .ZN(n6905) );
  NAND2_X1 U8734 ( .A1(n6906), .A2(n6905), .ZN(n6908) );
  INV_X1 U8735 ( .A(n6913), .ZN(n6907) );
  XNOR2_X1 U8736 ( .A(n6908), .B(n6907), .ZN(n6909) );
  NAND2_X1 U8737 ( .A1(n6909), .A2(n9301), .ZN(n6911) );
  NAND2_X1 U8738 ( .A1(n8729), .A2(n9224), .ZN(n6910) );
  NAND2_X1 U8739 ( .A1(n6911), .A2(n6910), .ZN(n9686) );
  INV_X1 U8740 ( .A(n9686), .ZN(n6924) );
  OAI21_X1 U8741 ( .B1(n6914), .B2(n6913), .A(n6912), .ZN(n9688) );
  INV_X1 U8742 ( .A(n6915), .ZN(n6917) );
  AOI211_X1 U8743 ( .C1(n6919), .C2(n6917), .A(n9308), .B(n6916), .ZN(n6918)
         );
  AOI21_X1 U8744 ( .B1(n9222), .B2(n8727), .A(n6918), .ZN(n9684) );
  AOI22_X1 U8745 ( .A1(n4251), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7026), .B2(
        n9312), .ZN(n6921) );
  NAND2_X1 U8746 ( .A1(n6919), .A2(n9005), .ZN(n6920) );
  OAI211_X1 U8747 ( .C1(n9684), .C2(n8982), .A(n6921), .B(n6920), .ZN(n6922)
         );
  AOI21_X1 U8748 ( .B1(n4648), .B2(n9688), .A(n6922), .ZN(n6923) );
  OAI21_X1 U8749 ( .B1(n4251), .B2(n6924), .A(n6923), .ZN(P1_U3284) );
  OAI22_X1 U8750 ( .A1(n9306), .A2(n6925), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9257), .ZN(n6926) );
  AOI21_X1 U8751 ( .B1(n9005), .B2(n8315), .A(n6926), .ZN(n6927) );
  OAI21_X1 U8752 ( .B1(n8982), .B2(n6928), .A(n6927), .ZN(n6929) );
  AOI21_X1 U8753 ( .B1(n6930), .B2(n4648), .A(n6929), .ZN(n6931) );
  OAI21_X1 U8754 ( .B1(n6932), .B2(n4251), .A(n6931), .ZN(P1_U3290) );
  INV_X1 U8755 ( .A(n6933), .ZN(n7397) );
  OAI222_X1 U8756 ( .A1(P2_U3151), .A2(n7888), .B1(n8277), .B2(n7397), .C1(
        n6934), .C2(n8276), .ZN(P2_U3276) );
  XNOR2_X1 U8757 ( .A(n6935), .B(n7019), .ZN(n6936) );
  NOR2_X1 U8758 ( .A1(n6936), .A2(n6937), .ZN(n7018) );
  AOI21_X1 U8759 ( .B1(n6937), .B2(n6936), .A(n7018), .ZN(n6945) );
  NAND2_X1 U8760 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9559) );
  INV_X1 U8761 ( .A(n9559), .ZN(n6941) );
  OAI22_X1 U8762 ( .A1(n8430), .A2(n6939), .B1(n6938), .B2(n8429), .ZN(n6940)
         );
  AOI211_X1 U8763 ( .C1(n8433), .C2(n4820), .A(n6941), .B(n6940), .ZN(n6944)
         );
  NAND2_X1 U8764 ( .A1(n6942), .A2(n8422), .ZN(n6943) );
  OAI211_X1 U8765 ( .C1(n6945), .C2(n8424), .A(n6944), .B(n6943), .ZN(P1_U3221) );
  NAND2_X1 U8766 ( .A1(n6946), .A2(n8162), .ZN(n6947) );
  XNOR2_X1 U8767 ( .A(n7439), .B(n7096), .ZN(n6949) );
  NAND2_X1 U8768 ( .A1(n6949), .A2(n7144), .ZN(n7031) );
  INV_X1 U8769 ( .A(n6949), .ZN(n6950) );
  NAND2_X1 U8770 ( .A1(n7831), .A2(n6950), .ZN(n6951) );
  NAND2_X1 U8771 ( .A1(n7031), .A2(n6951), .ZN(n6953) );
  INV_X1 U8772 ( .A(n7032), .ZN(n7030) );
  AOI21_X1 U8773 ( .B1(n6954), .B2(n6953), .A(n7030), .ZN(n6961) );
  OAI22_X1 U8774 ( .A1(n6955), .A2(n7575), .B1(n7598), .B2(n7105), .ZN(n6956)
         );
  AOI211_X1 U8775 ( .C1(n7096), .C2(n7587), .A(n6957), .B(n6956), .ZN(n6960)
         );
  INV_X1 U8776 ( .A(n6958), .ZN(n7095) );
  NAND2_X1 U8777 ( .A1(n7600), .A2(n7095), .ZN(n6959) );
  OAI211_X1 U8778 ( .C1(n6961), .C2(n7589), .A(n6960), .B(n6959), .ZN(P2_U3170) );
  NAND2_X1 U8779 ( .A1(n6962), .A2(n4648), .ZN(n6968) );
  INV_X1 U8780 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6963) );
  OAI22_X1 U8781 ( .A1(n9306), .A2(n6963), .B1(n9576), .B2(n9257), .ZN(n6966)
         );
  NOR2_X1 U8782 ( .A1(n6964), .A2(n8982), .ZN(n6965) );
  AOI211_X1 U8783 ( .C1(n9005), .C2(n6970), .A(n6966), .B(n6965), .ZN(n6967)
         );
  OAI211_X1 U8784 ( .C1(n4251), .C2(n6969), .A(n6968), .B(n6967), .ZN(P1_U3283) );
  OR2_X1 U8785 ( .A1(n6970), .A2(n8727), .ZN(n6971) );
  NAND2_X1 U8786 ( .A1(n6972), .A2(n6971), .ZN(n6973) );
  INV_X1 U8787 ( .A(n8726), .ZN(n7112) );
  OR2_X1 U8788 ( .A1(n7110), .A2(n7112), .ZN(n8488) );
  NAND2_X1 U8789 ( .A1(n7110), .A2(n7112), .ZN(n8492) );
  NAND2_X1 U8790 ( .A1(n8488), .A2(n8492), .ZN(n7115) );
  NOR2_X1 U8791 ( .A1(n6973), .A2(n7115), .ZN(n6974) );
  NAND2_X1 U8792 ( .A1(n7117), .A2(n8490), .ZN(n6975) );
  XNOR2_X1 U8793 ( .A(n6975), .B(n7115), .ZN(n6977) );
  AOI22_X1 U8794 ( .A1(n9224), .A2(n8727), .B1(n7206), .B2(n9222), .ZN(n6976)
         );
  OAI21_X1 U8795 ( .B1(n6977), .B2(n9283), .A(n6976), .ZN(n6978) );
  AOI21_X1 U8796 ( .B1(n9696), .B2(n6979), .A(n6978), .ZN(n9698) );
  NAND2_X1 U8797 ( .A1(n6980), .A2(n7110), .ZN(n6981) );
  NAND2_X1 U8798 ( .A1(n6981), .A2(n9373), .ZN(n6982) );
  OR2_X1 U8799 ( .A1(n6982), .A2(n7121), .ZN(n9691) );
  AOI22_X1 U8800 ( .A1(n4251), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7165), .B2(
        n9312), .ZN(n6984) );
  NAND2_X1 U8801 ( .A1(n7110), .A2(n9005), .ZN(n6983) );
  OAI211_X1 U8802 ( .C1(n9691), .C2(n8982), .A(n6984), .B(n6983), .ZN(n6985)
         );
  AOI21_X1 U8803 ( .B1(n9696), .B2(n6986), .A(n6985), .ZN(n6987) );
  OAI21_X1 U8804 ( .B1(n9698), .B2(n4251), .A(n6987), .ZN(P1_U3282) );
  INV_X1 U8805 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6988) );
  OAI22_X1 U8806 ( .A1(n9483), .A2(n6989), .B1(n9701), .B2(n6988), .ZN(n6990)
         );
  INV_X1 U8807 ( .A(n6990), .ZN(n6991) );
  OAI21_X1 U8808 ( .B1(n6992), .B2(n9699), .A(n6991), .ZN(P1_U3465) );
  INV_X1 U8809 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6993) );
  OAI22_X1 U8810 ( .A1(n9483), .A2(n6994), .B1(n9701), .B2(n6993), .ZN(n6995)
         );
  INV_X1 U8811 ( .A(n6995), .ZN(n6996) );
  OAI21_X1 U8812 ( .B1(n6997), .B2(n9699), .A(n6996), .ZN(P1_U3459) );
  NOR2_X1 U8813 ( .A1(n8819), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6998) );
  AOI21_X1 U8814 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n8819), .A(n6998), .ZN(
        n7003) );
  NAND2_X1 U8815 ( .A1(n9532), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6999) );
  OAI21_X1 U8816 ( .B1(n9532), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6999), .ZN(
        n9528) );
  OAI21_X1 U8817 ( .B1(n7006), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7000), .ZN(
        n9529) );
  NOR2_X1 U8818 ( .A1(n9528), .A2(n9529), .ZN(n9527) );
  AOI21_X1 U8819 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n9532), .A(n9527), .ZN(
        n9592) );
  NAND2_X1 U8820 ( .A1(n7008), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7001) );
  OAI21_X1 U8821 ( .B1(n7008), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7001), .ZN(
        n9593) );
  NOR2_X1 U8822 ( .A1(n9592), .A2(n9593), .ZN(n9591) );
  AOI21_X1 U8823 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n7008), .A(n9591), .ZN(
        n7002) );
  NAND2_X1 U8824 ( .A1(n7003), .A2(n7002), .ZN(n8818) );
  OAI21_X1 U8825 ( .B1(n7003), .B2(n7002), .A(n8818), .ZN(n7004) );
  NAND2_X1 U8826 ( .A1(n7004), .A2(n9595), .ZN(n7017) );
  MUX2_X1 U8827 ( .A(n6804), .B(P1_REG1_REG_10__SCAN_IN), .S(n9532), .Z(n9525)
         );
  OAI21_X1 U8828 ( .B1(n7006), .B2(P1_REG1_REG_9__SCAN_IN), .A(n7005), .ZN(
        n9526) );
  INV_X1 U8829 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7007) );
  MUX2_X1 U8830 ( .A(n7007), .B(P1_REG1_REG_11__SCAN_IN), .S(n7008), .Z(n9598)
         );
  INV_X1 U8831 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7009) );
  AOI22_X1 U8832 ( .A1(n8819), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n7009), .B2(
        n7013), .ZN(n7010) );
  NAND2_X1 U8833 ( .A1(n7011), .A2(n7010), .ZN(n8811) );
  OAI21_X1 U8834 ( .B1(n7011), .B2(n7010), .A(n8811), .ZN(n7015) );
  NAND2_X1 U8835 ( .A1(n8835), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n7012) );
  NAND2_X1 U8836 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7231) );
  OAI211_X1 U8837 ( .C1(n9654), .C2(n7013), .A(n7012), .B(n7231), .ZN(n7014)
         );
  AOI21_X1 U8838 ( .B1(n7015), .B2(n9648), .A(n7014), .ZN(n7016) );
  NAND2_X1 U8839 ( .A1(n7017), .A2(n7016), .ZN(P1_U3255) );
  AOI21_X1 U8840 ( .B1(n6935), .B2(n7019), .A(n7018), .ZN(n7022) );
  OAI211_X1 U8841 ( .C1(n7022), .C2(n7021), .A(n9573), .B(n7020), .ZN(n7028)
         );
  OAI22_X1 U8842 ( .A1(n8430), .A2(n7023), .B1(n7162), .B2(n8429), .ZN(n7024)
         );
  AOI211_X1 U8843 ( .C1(n8433), .C2(n7026), .A(n7025), .B(n7024), .ZN(n7027)
         );
  OAI211_X1 U8844 ( .C1(n9685), .C2(n9570), .A(n7028), .B(n7027), .ZN(P1_U3231) );
  INV_X1 U8845 ( .A(n7031), .ZN(n7029) );
  INV_X4 U8846 ( .A(n6655), .ZN(n7439) );
  XNOR2_X1 U8847 ( .A(n7439), .B(n9921), .ZN(n7099) );
  XNOR2_X1 U8848 ( .A(n7099), .B(n7105), .ZN(n7033) );
  NOR3_X1 U8849 ( .A1(n7030), .A2(n7029), .A3(n7033), .ZN(n7036) );
  NAND2_X1 U8850 ( .A1(n7032), .A2(n7031), .ZN(n7034) );
  NAND2_X1 U8851 ( .A1(n7034), .A2(n7033), .ZN(n7102) );
  INV_X1 U8852 ( .A(n7102), .ZN(n7035) );
  OAI21_X1 U8853 ( .B1(n7036), .B2(n7035), .A(n7591), .ZN(n7041) );
  OAI22_X1 U8854 ( .A1(n7144), .A2(n7575), .B1(n7598), .B2(n7188), .ZN(n7037)
         );
  AOI211_X1 U8855 ( .C1(n7039), .C2(n7587), .A(n7038), .B(n7037), .ZN(n7040)
         );
  OAI211_X1 U8856 ( .C1(n7141), .C2(n7558), .A(n7041), .B(n7040), .ZN(P2_U3167) );
  INV_X1 U8857 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n7042) );
  OAI22_X1 U8858 ( .A1(n9483), .A2(n7043), .B1(n9701), .B2(n7042), .ZN(n7044)
         );
  AOI21_X1 U8859 ( .B1(n7045), .B2(n9701), .A(n7044), .ZN(n7046) );
  INV_X1 U8860 ( .A(n7046), .ZN(P1_U3462) );
  NAND2_X1 U8861 ( .A1(n9479), .A2(n9689), .ZN(n9472) );
  INV_X1 U8862 ( .A(n9472), .ZN(n7050) );
  INV_X1 U8863 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7047) );
  OAI22_X1 U8864 ( .A1(n9483), .A2(n7048), .B1(n9479), .B2(n7047), .ZN(n7049)
         );
  AOI21_X1 U8865 ( .B1(n7051), .B2(n7050), .A(n7049), .ZN(n7052) );
  OAI21_X1 U8866 ( .B1(n7053), .B2(n9699), .A(n7052), .ZN(P1_U3471) );
  INV_X1 U8867 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7054) );
  OAI22_X1 U8868 ( .A1(n9483), .A2(n8452), .B1(n9479), .B2(n7054), .ZN(n7055)
         );
  AOI21_X1 U8869 ( .B1(n7056), .B2(n9701), .A(n7055), .ZN(n7057) );
  INV_X1 U8870 ( .A(n7057), .ZN(P1_U3468) );
  INV_X1 U8871 ( .A(n7060), .ZN(n7630) );
  XNOR2_X1 U8872 ( .A(n7085), .B(n7630), .ZN(n7058) );
  AOI222_X1 U8873 ( .A1(n8167), .A2(n7058), .B1(n7831), .B2(n8161), .C1(n7832), 
        .C2(n8092), .ZN(n9911) );
  XNOR2_X1 U8874 ( .A(n7059), .B(n7060), .ZN(n9914) );
  INV_X1 U8875 ( .A(n9903), .ZN(n7061) );
  NAND2_X1 U8876 ( .A1(n7061), .A2(n7155), .ZN(n7062) );
  AOI22_X1 U8877 ( .A1(n8086), .A2(n7063), .B1(n4911), .B2(n8102), .ZN(n7064)
         );
  OAI21_X1 U8878 ( .B1(n7065), .B2(n8098), .A(n7064), .ZN(n7066) );
  AOI21_X1 U8879 ( .B1(n9914), .B2(n8065), .A(n7066), .ZN(n7067) );
  OAI21_X1 U8880 ( .B1(n9911), .B2(n9907), .A(n7067), .ZN(P2_U3230) );
  INV_X1 U8881 ( .A(n7068), .ZN(n7077) );
  OAI222_X1 U8882 ( .A1(n9500), .A2(n7077), .B1(n4263), .B2(P1_U3086), .C1(
        n7069), .C2(n7398), .ZN(P1_U3335) );
  INV_X1 U8883 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7071) );
  OAI22_X1 U8884 ( .A1(n9571), .A2(n9483), .B1(n9479), .B2(n7071), .ZN(n7072)
         );
  AOI21_X1 U8885 ( .B1(n7073), .B2(n9701), .A(n7072), .ZN(n7074) );
  OAI21_X1 U8886 ( .B1(n7075), .B2(n9472), .A(n7074), .ZN(P1_U3483) );
  OAI222_X1 U8887 ( .A1(n7804), .A2(P2_U3151), .B1(n8277), .B2(n7077), .C1(
        n7076), .C2(n8276), .ZN(P2_U3275) );
  INV_X1 U8888 ( .A(n7078), .ZN(n7081) );
  OAI222_X1 U8889 ( .A1(n9500), .A2(n7081), .B1(n8651), .B2(P1_U3086), .C1(
        n7079), .C2(n7398), .ZN(P1_U3334) );
  OAI222_X1 U8890 ( .A1(n7662), .A2(P2_U3151), .B1(n8277), .B2(n7081), .C1(
        n7080), .C2(n8276), .ZN(P2_U3274) );
  NAND2_X1 U8891 ( .A1(n7082), .A2(n7693), .ZN(n7083) );
  XOR2_X1 U8892 ( .A(n7678), .B(n7083), .Z(n9916) );
  OR2_X1 U8893 ( .A1(n7085), .A2(n7084), .ZN(n7087) );
  NAND2_X1 U8894 ( .A1(n7087), .A2(n7086), .ZN(n7088) );
  NAND2_X1 U8895 ( .A1(n7088), .A2(n7678), .ZN(n7089) );
  NAND2_X1 U8896 ( .A1(n7090), .A2(n7089), .ZN(n7093) );
  NAND2_X1 U8897 ( .A1(n8162), .A2(n8092), .ZN(n7091) );
  OAI21_X1 U8898 ( .B1(n7105), .B2(n8080), .A(n7091), .ZN(n7092) );
  AOI21_X1 U8899 ( .B1(n7093), .B2(n8167), .A(n7092), .ZN(n9917) );
  MUX2_X1 U8900 ( .A(n9917), .B(n7094), .S(n9907), .Z(n7098) );
  AOI22_X1 U8901 ( .A1(n8086), .A2(n7096), .B1(n8102), .B2(n7095), .ZN(n7097)
         );
  OAI211_X1 U8902 ( .C1(n8105), .C2(n9916), .A(n7098), .B(n7097), .ZN(P2_U3229) );
  INV_X1 U8903 ( .A(n7099), .ZN(n7100) );
  NAND2_X1 U8904 ( .A1(n7100), .A2(n7105), .ZN(n7101) );
  XNOR2_X1 U8905 ( .A(n7439), .B(n9927), .ZN(n7179) );
  XNOR2_X1 U8906 ( .A(n7179), .B(n7188), .ZN(n7103) );
  OAI211_X1 U8907 ( .C1(n7104), .C2(n7103), .A(n7181), .B(n7591), .ZN(n7109)
         );
  OAI22_X1 U8908 ( .A1(n7105), .A2(n7575), .B1(n7598), .B2(n7282), .ZN(n7106)
         );
  AOI211_X1 U8909 ( .C1(n7136), .C2(n7587), .A(n7107), .B(n7106), .ZN(n7108)
         );
  OAI211_X1 U8910 ( .C1(n7134), .C2(n7558), .A(n7109), .B(n7108), .ZN(P2_U3179) );
  INV_X1 U8911 ( .A(n7110), .ZN(n9693) );
  NAND2_X1 U8912 ( .A1(n7175), .A2(n8388), .ZN(n8493) );
  AOI21_X1 U8913 ( .B1(n7113), .B2(n7203), .A(n7196), .ZN(n7168) );
  INV_X1 U8914 ( .A(n8490), .ZN(n7114) );
  NOR2_X1 U8915 ( .A1(n7115), .A2(n7114), .ZN(n7116) );
  XNOR2_X1 U8916 ( .A(n7204), .B(n7203), .ZN(n7120) );
  NAND2_X1 U8917 ( .A1(n8725), .A2(n9222), .ZN(n7119) );
  NAND2_X1 U8918 ( .A1(n8726), .A2(n9224), .ZN(n7118) );
  AND2_X1 U8919 ( .A1(n7119), .A2(n7118), .ZN(n7232) );
  OAI21_X1 U8920 ( .B1(n7120), .B2(n9283), .A(n7232), .ZN(n7169) );
  INV_X1 U8921 ( .A(n7121), .ZN(n7122) );
  AOI211_X1 U8922 ( .C1(n7175), .C2(n7122), .A(n9308), .B(n7198), .ZN(n7170)
         );
  NAND2_X1 U8923 ( .A1(n7170), .A2(n9317), .ZN(n7124) );
  AOI22_X1 U8924 ( .A1(n4251), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7234), .B2(
        n9312), .ZN(n7123) );
  OAI211_X1 U8925 ( .C1(n7237), .C2(n9315), .A(n7124), .B(n7123), .ZN(n7125)
         );
  AOI21_X1 U8926 ( .B1(n9306), .B2(n7169), .A(n7125), .ZN(n7126) );
  OAI21_X1 U8927 ( .B1(n7168), .B2(n9294), .A(n7126), .ZN(P1_U3281) );
  XNOR2_X1 U8928 ( .A(n7188), .B(n9927), .ZN(n7632) );
  AND2_X1 U8929 ( .A1(n7128), .A2(n7127), .ZN(n7140) );
  NAND2_X1 U8930 ( .A1(n7140), .A2(n7633), .ZN(n7139) );
  NAND2_X1 U8931 ( .A1(n7139), .A2(n7129), .ZN(n7130) );
  XOR2_X1 U8932 ( .A(n7632), .B(n7130), .Z(n9928) );
  XNOR2_X1 U8933 ( .A(n7131), .B(n7632), .ZN(n7132) );
  AOI222_X1 U8934 ( .A1(n8167), .A2(n7132), .B1(n7828), .B2(n8161), .C1(n7830), 
        .C2(n8092), .ZN(n9926) );
  MUX2_X1 U8935 ( .A(n7133), .B(n9926), .S(n9904), .Z(n7138) );
  INV_X1 U8936 ( .A(n7134), .ZN(n7135) );
  AOI22_X1 U8937 ( .A1(n8086), .A2(n7136), .B1(n8102), .B2(n7135), .ZN(n7137)
         );
  OAI211_X1 U8938 ( .C1(n9928), .C2(n8105), .A(n7138), .B(n7137), .ZN(P2_U3227) );
  OAI21_X1 U8939 ( .B1(n7140), .B2(n7633), .A(n7139), .ZN(n9924) );
  OAI22_X1 U8940 ( .A1(n7955), .A2(n9921), .B1(n7141), .B2(n9896), .ZN(n7146)
         );
  XNOR2_X1 U8941 ( .A(n7142), .B(n7633), .ZN(n7143) );
  OAI222_X1 U8942 ( .A1(n8080), .A2(n7188), .B1(n8164), .B2(n7144), .C1(n8037), 
        .C2(n7143), .ZN(n9922) );
  MUX2_X1 U8943 ( .A(n9922), .B(P2_REG2_REG_5__SCAN_IN), .S(n9907), .Z(n7145)
         );
  AOI211_X1 U8944 ( .C1(n9924), .C2(n8065), .A(n7146), .B(n7145), .ZN(n7147)
         );
  INV_X1 U8945 ( .A(n7147), .ZN(P2_U3228) );
  OAI21_X1 U8946 ( .B1(n7148), .B2(n7701), .A(n7149), .ZN(n9933) );
  OAI21_X1 U8947 ( .B1(n7151), .B2(n5423), .A(n7150), .ZN(n7152) );
  NAND2_X1 U8948 ( .A1(n7152), .A2(n8167), .ZN(n7154) );
  AOI22_X1 U8949 ( .A1(n7829), .A2(n8092), .B1(n8161), .B2(n7827), .ZN(n7153)
         );
  OAI211_X1 U8950 ( .C1(n7155), .C2(n9933), .A(n7154), .B(n7153), .ZN(n9935)
         );
  NAND2_X1 U8951 ( .A1(n9935), .A2(n8098), .ZN(n7158) );
  OAI22_X1 U8952 ( .A1(n9904), .A2(n4976), .B1(n7191), .B2(n9896), .ZN(n7156)
         );
  AOI21_X1 U8953 ( .B1(n8086), .B2(n7182), .A(n7156), .ZN(n7157) );
  OAI211_X1 U8954 ( .C1(n9933), .C2(n7306), .A(n7158), .B(n7157), .ZN(P2_U3226) );
  AND3_X1 U8955 ( .A1(n4384), .A2(n4374), .A3(n7159), .ZN(n7161) );
  OAI21_X1 U8956 ( .B1(n7228), .B2(n7161), .A(n9573), .ZN(n7167) );
  NAND2_X1 U8957 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9604) );
  INV_X1 U8958 ( .A(n9604), .ZN(n7164) );
  OAI22_X1 U8959 ( .A1(n8430), .A2(n7162), .B1(n8388), .B2(n8429), .ZN(n7163)
         );
  AOI211_X1 U8960 ( .C1(n7165), .C2(n8433), .A(n7164), .B(n7163), .ZN(n7166)
         );
  OAI211_X1 U8961 ( .C1(n9693), .C2(n9570), .A(n7167), .B(n7166), .ZN(P1_U3236) );
  INV_X1 U8962 ( .A(n7168), .ZN(n7171) );
  AOI211_X1 U8963 ( .C1(n7171), .C2(n9689), .A(n7170), .B(n7169), .ZN(n7177)
         );
  INV_X1 U8964 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7172) );
  OAI22_X1 U8965 ( .A1(n7237), .A2(n9483), .B1(n9479), .B2(n7172), .ZN(n7173)
         );
  INV_X1 U8966 ( .A(n7173), .ZN(n7174) );
  OAI21_X1 U8967 ( .B1(n7177), .B2(n9699), .A(n7174), .ZN(P1_U3489) );
  AOI22_X1 U8968 ( .A1(n7175), .A2(n9360), .B1(n9706), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n7176) );
  OAI21_X1 U8969 ( .B1(n7177), .B2(n9706), .A(n7176), .ZN(P1_U3534) );
  INV_X1 U8970 ( .A(n7178), .ZN(n7390) );
  OAI222_X1 U8971 ( .A1(P2_U3151), .A2(n7663), .B1(n8277), .B2(n7390), .C1(
        n9092), .C2(n8276), .ZN(P2_U3273) );
  NAND2_X1 U8972 ( .A1(n7829), .A2(n7179), .ZN(n7180) );
  XNOR2_X1 U8973 ( .A(n7439), .B(n7182), .ZN(n7183) );
  NAND2_X1 U8974 ( .A1(n7183), .A2(n7282), .ZN(n7289) );
  INV_X1 U8975 ( .A(n7183), .ZN(n7184) );
  NAND2_X1 U8976 ( .A1(n7828), .A2(n7184), .ZN(n7185) );
  AND2_X1 U8977 ( .A1(n7289), .A2(n7185), .ZN(n7186) );
  OAI21_X1 U8978 ( .B1(n7187), .B2(n7186), .A(n7286), .ZN(n7194) );
  NOR2_X1 U8979 ( .A1(n7603), .A2(n9932), .ZN(n7193) );
  AND2_X1 U8980 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n9728) );
  AOI21_X1 U8981 ( .B1(n7573), .B2(n7827), .A(n9728), .ZN(n7190) );
  OR2_X1 U8982 ( .A1(n7575), .A2(n7188), .ZN(n7189) );
  OAI211_X1 U8983 ( .C1(n7191), .C2(n7558), .A(n7190), .B(n7189), .ZN(n7192)
         );
  AOI211_X1 U8984 ( .C1(n7194), .C2(n7591), .A(n7193), .B(n7192), .ZN(n7195)
         );
  INV_X1 U8985 ( .A(n7195), .ZN(P2_U3153) );
  NOR2_X1 U8986 ( .A1(n9408), .A2(n8872), .ZN(n8498) );
  INV_X1 U8987 ( .A(n8498), .ZN(n8668) );
  NOR2_X1 U8988 ( .A1(n7197), .A2(n8589), .ZN(n8874) );
  AOI21_X1 U8989 ( .B1(n7197), .B2(n8589), .A(n8874), .ZN(n9412) );
  INV_X1 U8990 ( .A(n7198), .ZN(n7200) );
  INV_X1 U8991 ( .A(n9310), .ZN(n7199) );
  AOI211_X1 U8992 ( .C1(n9408), .C2(n7200), .A(n9308), .B(n7199), .ZN(n9407)
         );
  AOI22_X1 U8993 ( .A1(n4251), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n8391), .B2(
        n9312), .ZN(n7201) );
  OAI21_X1 U8994 ( .B1(n8871), .B2(n9315), .A(n7201), .ZN(n7209) );
  INV_X1 U8995 ( .A(n8494), .ZN(n7202) );
  OAI21_X1 U8996 ( .B1(n8589), .B2(n7205), .A(n9298), .ZN(n7207) );
  AOI222_X1 U8997 ( .A1(n9301), .A2(n7207), .B1(n7206), .B2(n9224), .C1(n8724), 
        .C2(n9222), .ZN(n9410) );
  NOR2_X1 U8998 ( .A1(n9410), .A2(n4251), .ZN(n7208) );
  AOI211_X1 U8999 ( .C1(n9407), .C2(n9317), .A(n7209), .B(n7208), .ZN(n7210)
         );
  OAI21_X1 U9000 ( .B1(n9412), .B2(n9294), .A(n7210), .ZN(P1_U3280) );
  XNOR2_X1 U9001 ( .A(n7827), .B(n9937), .ZN(n7637) );
  XOR2_X1 U9002 ( .A(n7211), .B(n7637), .Z(n9938) );
  XOR2_X1 U9003 ( .A(n7212), .B(n7637), .Z(n7213) );
  OAI222_X1 U9004 ( .A1(n8080), .A2(n7378), .B1(n8164), .B2(n7282), .C1(n7213), 
        .C2(n8037), .ZN(n9940) );
  NAND2_X1 U9005 ( .A1(n9940), .A2(n8098), .ZN(n7217) );
  INV_X1 U9006 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7214) );
  OAI22_X1 U9007 ( .A1(n9904), .A2(n7214), .B1(n7285), .B2(n9896), .ZN(n7215)
         );
  AOI21_X1 U9008 ( .B1(n8086), .B2(n7294), .A(n7215), .ZN(n7216) );
  OAI211_X1 U9009 ( .C1(n8105), .C2(n9938), .A(n7217), .B(n7216), .ZN(P2_U3225) );
  INV_X1 U9010 ( .A(n7221), .ZN(n7220) );
  INV_X1 U9011 ( .A(n8715), .ZN(n7218) );
  AOI21_X1 U9012 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n9497), .A(n7218), .ZN(
        n7219) );
  OAI21_X1 U9013 ( .B1(n7220), .B2(n9500), .A(n7219), .ZN(P1_U3332) );
  NAND2_X1 U9014 ( .A1(n7221), .A2(n7353), .ZN(n7223) );
  NAND2_X1 U9015 ( .A1(n7222), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7817) );
  OAI211_X1 U9016 ( .C1(n7224), .C2(n8276), .A(n7223), .B(n7817), .ZN(P2_U3272) );
  INV_X1 U9017 ( .A(n7225), .ZN(n7230) );
  NOR3_X1 U9018 ( .A1(n7228), .A2(n7227), .A3(n7226), .ZN(n7229) );
  OAI21_X1 U9019 ( .B1(n7230), .B2(n7229), .A(n9573), .ZN(n7236) );
  OAI21_X1 U9020 ( .B1(n8419), .B2(n7232), .A(n7231), .ZN(n7233) );
  AOI21_X1 U9021 ( .B1(n7234), .B2(n8433), .A(n7233), .ZN(n7235) );
  OAI211_X1 U9022 ( .C1(n7237), .C2(n9570), .A(n7236), .B(n7235), .ZN(P1_U3224) );
  INV_X1 U9023 ( .A(n7238), .ZN(n7400) );
  OAI222_X1 U9024 ( .A1(n9500), .A2(n7400), .B1(P1_U3086), .B2(n7240), .C1(
        n7239), .C2(n7398), .ZN(P1_U3331) );
  NAND2_X1 U9025 ( .A1(n7253), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7241) );
  XNOR2_X1 U9026 ( .A(n7243), .B(n7256), .ZN(n9727) );
  INV_X1 U9027 ( .A(n7256), .ZN(n9729) );
  INV_X1 U9028 ( .A(n7243), .ZN(n7244) );
  OAI22_X1 U9029 ( .A1(n9727), .A2(n4976), .B1(n9729), .B2(n7244), .ZN(n9753)
         );
  MUX2_X1 U9030 ( .A(n7214), .B(P2_REG2_REG_8__SCAN_IN), .S(n9743), .Z(n9752)
         );
  INV_X1 U9031 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7302) );
  XNOR2_X1 U9032 ( .A(n7893), .B(n7302), .ZN(n7267) );
  XNOR2_X1 U9033 ( .A(n7875), .B(n7892), .ZN(n7876) );
  XNOR2_X1 U9034 ( .A(n7250), .B(n9743), .ZN(n9745) );
  INV_X1 U9035 ( .A(n7245), .ZN(n7247) );
  XNOR2_X1 U9036 ( .A(n7249), .B(n7256), .ZN(n9737) );
  OAI22_X1 U9037 ( .A1(n9738), .A2(n9737), .B1(n7249), .B2(n7256), .ZN(n9746)
         );
  NAND2_X1 U9038 ( .A1(n9745), .A2(n9746), .ZN(n9744) );
  OAI21_X1 U9039 ( .B1(n7250), .B2(n7252), .A(n9744), .ZN(n7874) );
  XNOR2_X1 U9040 ( .A(n7876), .B(n7874), .ZN(n7251) );
  NOR2_X1 U9041 ( .A1(n7251), .A2(n9508), .ZN(n7265) );
  AOI22_X1 U9042 ( .A1(n9743), .A2(n4990), .B1(P2_REG1_REG_8__SCAN_IN), .B2(
        n7252), .ZN(n9749) );
  NAND2_X1 U9043 ( .A1(n7253), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7254) );
  NAND2_X1 U9044 ( .A1(n7255), .A2(n7254), .ZN(n7257) );
  XNOR2_X1 U9045 ( .A(n7257), .B(n7256), .ZN(n9730) );
  INV_X1 U9046 ( .A(n7257), .ZN(n7258) );
  OAI22_X1 U9047 ( .A1(n9730), .A2(n7259), .B1(n9729), .B2(n7258), .ZN(n9750)
         );
  XNOR2_X1 U9048 ( .A(n7850), .B(n7261), .ZN(n7851) );
  INV_X1 U9049 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7260) );
  XNOR2_X1 U9050 ( .A(n7851), .B(n7260), .ZN(n7263) );
  NAND2_X1 U9051 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7333) );
  NAND2_X1 U9052 ( .A1(n9875), .A2(n7261), .ZN(n7262) );
  OAI211_X1 U9053 ( .C1(n9732), .C2(n7263), .A(n7333), .B(n7262), .ZN(n7264)
         );
  AOI211_X1 U9054 ( .C1(n9874), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n7265), .B(
        n7264), .ZN(n7266) );
  OAI21_X1 U9055 ( .B1(n7267), .B2(n9890), .A(n7266), .ZN(P2_U3191) );
  NAND2_X1 U9056 ( .A1(n7268), .A2(n7690), .ZN(n7269) );
  NAND2_X1 U9057 ( .A1(n7269), .A2(n7636), .ZN(n7271) );
  NAND2_X1 U9058 ( .A1(n7271), .A2(n7270), .ZN(n9952) );
  INV_X1 U9059 ( .A(n9952), .ZN(n7280) );
  XOR2_X1 U9060 ( .A(n7272), .B(n7636), .Z(n7275) );
  OAI22_X1 U9061 ( .A1(n4501), .A2(n8080), .B1(n7378), .B2(n8164), .ZN(n7273)
         );
  AOI21_X1 U9062 ( .B1(n9952), .B2(n8158), .A(n7273), .ZN(n7274) );
  OAI21_X1 U9063 ( .B1(n7275), .B2(n8037), .A(n7274), .ZN(n9950) );
  NAND2_X1 U9064 ( .A1(n9950), .A2(n8098), .ZN(n7279) );
  OAI22_X1 U9065 ( .A1(n9904), .A2(n7276), .B1(n7375), .B2(n9896), .ZN(n7277)
         );
  AOI21_X1 U9066 ( .B1(n8086), .B2(n9947), .A(n7277), .ZN(n7278) );
  OAI211_X1 U9067 ( .C1(n7280), .C2(n7306), .A(n7279), .B(n7278), .ZN(P2_U3223) );
  INV_X1 U9068 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7281) );
  NOR2_X1 U9069 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7281), .ZN(n9742) );
  NOR2_X1 U9070 ( .A1(n7575), .A2(n7282), .ZN(n7283) );
  AOI211_X1 U9071 ( .C1(n7573), .C2(n7826), .A(n9742), .B(n7283), .ZN(n7284)
         );
  OAI21_X1 U9072 ( .B1(n7285), .B2(n7558), .A(n7284), .ZN(n7293) );
  NAND2_X1 U9073 ( .A1(n7286), .A2(n7289), .ZN(n7287) );
  XNOR2_X1 U9074 ( .A(n9937), .B(n7439), .ZN(n7338) );
  XNOR2_X1 U9075 ( .A(n7338), .B(n7339), .ZN(n7288) );
  INV_X1 U9076 ( .A(n7288), .ZN(n7290) );
  NAND3_X1 U9077 ( .A1(n7286), .A2(n7290), .A3(n7289), .ZN(n7291) );
  AOI21_X1 U9078 ( .B1(n7342), .B2(n7291), .A(n7589), .ZN(n7292) );
  AOI211_X1 U9079 ( .C1(n7294), .C2(n7587), .A(n7293), .B(n7292), .ZN(n7295)
         );
  INV_X1 U9080 ( .A(n7295), .ZN(P2_U3161) );
  INV_X1 U9081 ( .A(n7268), .ZN(n7296) );
  AOI21_X1 U9082 ( .B1(n7297), .B2(n7635), .A(n7296), .ZN(n9945) );
  INV_X1 U9083 ( .A(n9945), .ZN(n7307) );
  XOR2_X1 U9084 ( .A(n7298), .B(n7635), .Z(n7301) );
  OAI22_X1 U9085 ( .A1(n7339), .A2(n8164), .B1(n7555), .B2(n8080), .ZN(n7299)
         );
  AOI21_X1 U9086 ( .B1(n9945), .B2(n8158), .A(n7299), .ZN(n7300) );
  OAI21_X1 U9087 ( .B1(n8037), .B2(n7301), .A(n7300), .ZN(n9943) );
  NAND2_X1 U9088 ( .A1(n9943), .A2(n8098), .ZN(n7305) );
  OAI22_X1 U9089 ( .A1(n9904), .A2(n7302), .B1(n7337), .B2(n9896), .ZN(n7303)
         );
  AOI21_X1 U9090 ( .B1(n8086), .B2(n7349), .A(n7303), .ZN(n7304) );
  OAI211_X1 U9091 ( .C1(n7307), .C2(n7306), .A(n7305), .B(n7304), .ZN(P2_U3224) );
  INV_X1 U9092 ( .A(n7308), .ZN(n7392) );
  OAI222_X1 U9093 ( .A1(n9500), .A2(n7392), .B1(P1_U3086), .B2(n7310), .C1(
        n7309), .C2(n7398), .ZN(P1_U3330) );
  INV_X1 U9094 ( .A(n7311), .ZN(n7320) );
  OAI222_X1 U9095 ( .A1(n9500), .A2(n7320), .B1(P1_U3086), .B2(n6151), .C1(
        n7312), .C2(n7398), .ZN(P1_U3329) );
  XNOR2_X1 U9096 ( .A(n7313), .B(n7627), .ZN(n9956) );
  XNOR2_X1 U9097 ( .A(n7314), .B(n7627), .ZN(n7315) );
  OAI222_X1 U9098 ( .A1(n8164), .A2(n7555), .B1(n8080), .B2(n7413), .C1(n8037), 
        .C2(n7315), .ZN(n9957) );
  NAND2_X1 U9099 ( .A1(n9957), .A2(n8098), .ZN(n7318) );
  INV_X1 U9100 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n9788) );
  OAI22_X1 U9101 ( .A1(n9904), .A2(n9788), .B1(n7559), .B2(n9896), .ZN(n7316)
         );
  AOI21_X1 U9102 ( .B1(n9959), .B2(n8086), .A(n7316), .ZN(n7317) );
  OAI211_X1 U9103 ( .C1(n9956), .C2(n8105), .A(n7318), .B(n7317), .ZN(P2_U3222) );
  OAI222_X1 U9104 ( .A1(n7321), .A2(P2_U3151), .B1(n8277), .B2(n7320), .C1(
        n7319), .C2(n8276), .ZN(P2_U3269) );
  INV_X1 U9105 ( .A(n6104), .ZN(n7396) );
  AOI21_X1 U9106 ( .B1(n8273), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n7322), .ZN(
        n7323) );
  OAI21_X1 U9107 ( .B1(n7396), .B2(n8277), .A(n7323), .ZN(P2_U3268) );
  XNOR2_X1 U9108 ( .A(n7324), .B(n7628), .ZN(n7325) );
  OAI222_X1 U9109 ( .A1(n8080), .A2(n7415), .B1(n8164), .B2(n4501), .C1(n7325), 
        .C2(n8037), .ZN(n9963) );
  INV_X1 U9110 ( .A(n9963), .ZN(n7332) );
  OAI22_X1 U9111 ( .A1(n9904), .A2(n7326), .B1(n7494), .B2(n9896), .ZN(n7327)
         );
  AOI21_X1 U9112 ( .B1(n9965), .B2(n8086), .A(n7327), .ZN(n7331) );
  NAND2_X1 U9113 ( .A1(n7329), .A2(n7628), .ZN(n9961) );
  NAND3_X1 U9114 ( .A1(n7328), .A2(n9961), .A3(n8065), .ZN(n7330) );
  OAI211_X1 U9115 ( .C1(n7332), .C2(n9907), .A(n7331), .B(n7330), .ZN(P2_U3221) );
  INV_X1 U9116 ( .A(n7333), .ZN(n7334) );
  AOI21_X1 U9117 ( .B1(n7573), .B2(n7825), .A(n7334), .ZN(n7336) );
  OR2_X1 U9118 ( .A1(n7575), .A2(n7339), .ZN(n7335) );
  OAI211_X1 U9119 ( .C1(n7337), .C2(n7558), .A(n7336), .B(n7335), .ZN(n7348)
         );
  XNOR2_X1 U9120 ( .A(n9942), .B(n7439), .ZN(n7369) );
  XNOR2_X1 U9121 ( .A(n7369), .B(n7826), .ZN(n7346) );
  INV_X1 U9122 ( .A(n7338), .ZN(n7340) );
  NAND2_X1 U9123 ( .A1(n7340), .A2(n7339), .ZN(n7341) );
  INV_X1 U9124 ( .A(n7346), .ZN(n7343) );
  INV_X1 U9125 ( .A(n7371), .ZN(n7344) );
  AOI211_X1 U9126 ( .C1(n7346), .C2(n7345), .A(n7589), .B(n7344), .ZN(n7347)
         );
  AOI211_X1 U9127 ( .C1(n7349), .C2(n7587), .A(n7348), .B(n7347), .ZN(n7350)
         );
  INV_X1 U9128 ( .A(n7350), .ZN(P2_U3171) );
  INV_X1 U9129 ( .A(n7354), .ZN(n7352) );
  AOI22_X1 U9130 ( .A1(n8749), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n9497), .ZN(n7351) );
  OAI21_X1 U9131 ( .B1(n7352), .B2(n9500), .A(n7351), .ZN(P1_U3327) );
  NAND2_X1 U9132 ( .A1(n7354), .A2(n7353), .ZN(n7356) );
  OAI211_X1 U9133 ( .C1(n8276), .C2(n7357), .A(n7356), .B(n7355), .ZN(P2_U3267) );
  INV_X1 U9134 ( .A(n7734), .ZN(n7359) );
  OR2_X1 U9135 ( .A1(n7660), .A2(n7359), .ZN(n7640) );
  XNOR2_X1 U9136 ( .A(n7358), .B(n7640), .ZN(n7389) );
  INV_X1 U9137 ( .A(n7640), .ZN(n7360) );
  XNOR2_X1 U9138 ( .A(n7361), .B(n7360), .ZN(n7363) );
  OAI22_X1 U9139 ( .A1(n8082), .A2(n8080), .B1(n7413), .B2(n8164), .ZN(n7362)
         );
  AOI21_X1 U9140 ( .B1(n7363), .B2(n8167), .A(n7362), .ZN(n7385) );
  INV_X1 U9141 ( .A(n7385), .ZN(n7366) );
  INV_X1 U9142 ( .A(n7659), .ZN(n7364) );
  OAI22_X1 U9143 ( .A1(n7364), .A2(n8096), .B1(n7542), .B2(n9896), .ZN(n7365)
         );
  OAI21_X1 U9144 ( .B1(n7366), .B2(n7365), .A(n8098), .ZN(n7368) );
  NAND2_X1 U9145 ( .A1(n9907), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7367) );
  OAI211_X1 U9146 ( .C1(n7389), .C2(n8105), .A(n7368), .B(n7367), .ZN(P2_U3220) );
  NAND2_X1 U9147 ( .A1(n7369), .A2(n7826), .ZN(n7370) );
  NAND2_X1 U9148 ( .A1(n7371), .A2(n7370), .ZN(n7412) );
  XNOR2_X1 U9149 ( .A(n7412), .B(n7555), .ZN(n7372) );
  XNOR2_X1 U9150 ( .A(n9947), .B(n6655), .ZN(n7402) );
  INV_X1 U9151 ( .A(n7402), .ZN(n7405) );
  NAND2_X1 U9152 ( .A1(n7372), .A2(n7405), .ZN(n7486) );
  OAI21_X1 U9153 ( .B1(n7372), .B2(n7405), .A(n7486), .ZN(n7373) );
  NAND2_X1 U9154 ( .A1(n7373), .A2(n7591), .ZN(n7381) );
  NAND2_X1 U9155 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n9775) );
  INV_X1 U9156 ( .A(n9775), .ZN(n7374) );
  AOI21_X1 U9157 ( .B1(n7573), .B2(n7824), .A(n7374), .ZN(n7377) );
  OR2_X1 U9158 ( .A1(n7558), .A2(n7375), .ZN(n7376) );
  OAI211_X1 U9159 ( .C1(n7378), .C2(n7575), .A(n7377), .B(n7376), .ZN(n7379)
         );
  AOI21_X1 U9160 ( .B1(n9947), .B2(n7587), .A(n7379), .ZN(n7380) );
  NAND2_X1 U9161 ( .A1(n7381), .A2(n7380), .ZN(P2_U3157) );
  INV_X1 U9162 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7382) );
  MUX2_X1 U9163 ( .A(n7382), .B(n7385), .S(n9967), .Z(n7384) );
  NAND2_X1 U9164 ( .A1(n7659), .A2(n8262), .ZN(n7383) );
  OAI211_X1 U9165 ( .C1(n7389), .C2(n8266), .A(n7384), .B(n7383), .ZN(P2_U3429) );
  MUX2_X1 U9166 ( .A(n7386), .B(n7385), .S(n9982), .Z(n7388) );
  NAND2_X1 U9167 ( .A1(n7659), .A2(n8152), .ZN(n7387) );
  OAI211_X1 U9168 ( .C1(n8155), .C2(n7389), .A(n7388), .B(n7387), .ZN(P2_U3472) );
  OAI222_X1 U9169 ( .A1(n7398), .A2(n7391), .B1(n9500), .B2(n7390), .C1(
        P1_U3086), .C2(n6171), .ZN(P1_U3333) );
  OAI222_X1 U9170 ( .A1(n7393), .A2(P2_U3151), .B1(n8277), .B2(n7392), .C1(
        n9053), .C2(n8276), .ZN(P2_U3270) );
  INV_X1 U9171 ( .A(n7607), .ZN(n9496) );
  OAI222_X1 U9172 ( .A1(n7394), .A2(P2_U3151), .B1(n8277), .B2(n9496), .C1(
        n7608), .C2(n8276), .ZN(P2_U3265) );
  OAI222_X1 U9173 ( .A1(n9500), .A2(n7396), .B1(n8748), .B2(P1_U3086), .C1(
        n7395), .C2(n7398), .ZN(P1_U3328) );
  OAI222_X1 U9174 ( .A1(n7398), .A2(n9142), .B1(n9500), .B2(n7397), .C1(
        P1_U3086), .C2(n8646), .ZN(P1_U3336) );
  OAI222_X1 U9175 ( .A1(n7401), .A2(P2_U3151), .B1(n8277), .B2(n7400), .C1(
        n7399), .C2(n8276), .ZN(P2_U3271) );
  XNOR2_X1 U9176 ( .A(n8250), .B(n7439), .ZN(n7422) );
  XNOR2_X1 U9177 ( .A(n9959), .B(n7439), .ZN(n7487) );
  NOR2_X1 U9178 ( .A1(n7487), .A2(n4501), .ZN(n7488) );
  INV_X1 U9179 ( .A(n7488), .ZN(n7404) );
  NAND2_X1 U9180 ( .A1(n7402), .A2(n7825), .ZN(n7403) );
  NAND2_X1 U9181 ( .A1(n7404), .A2(n7403), .ZN(n7411) );
  AND2_X1 U9182 ( .A1(n7405), .A2(n7555), .ZN(n7406) );
  INV_X1 U9183 ( .A(n7406), .ZN(n7408) );
  XNOR2_X1 U9184 ( .A(n9965), .B(n7439), .ZN(n7414) );
  XNOR2_X1 U9185 ( .A(n7414), .B(n7823), .ZN(n7490) );
  OAI21_X1 U9186 ( .B1(n7406), .B2(n4501), .A(n7487), .ZN(n7407) );
  OAI211_X1 U9187 ( .C1(n7824), .C2(n7408), .A(n7490), .B(n7407), .ZN(n7409)
         );
  XNOR2_X1 U9188 ( .A(n7659), .B(n7439), .ZN(n7536) );
  NOR2_X1 U9189 ( .A1(n7536), .A2(n7415), .ZN(n7417) );
  INV_X1 U9190 ( .A(n7536), .ZN(n7416) );
  XNOR2_X1 U9191 ( .A(n8263), .B(n7439), .ZN(n7418) );
  XNOR2_X1 U9192 ( .A(n7418), .B(n7822), .ZN(n7449) );
  XNOR2_X1 U9193 ( .A(n8256), .B(n7439), .ZN(n7420) );
  XNOR2_X1 U9194 ( .A(n7420), .B(n8094), .ZN(n7593) );
  NAND2_X1 U9195 ( .A1(n7594), .A2(n7593), .ZN(n7592) );
  NAND2_X1 U9196 ( .A1(n7592), .A2(n7421), .ZN(n7507) );
  XNOR2_X1 U9197 ( .A(n7422), .B(n8058), .ZN(n7506) );
  XNOR2_X1 U9198 ( .A(n8143), .B(n7439), .ZN(n7423) );
  XNOR2_X1 U9199 ( .A(n7423), .B(n7576), .ZN(n7515) );
  AND2_X1 U9200 ( .A1(n7423), .A2(n7576), .ZN(n7568) );
  XNOR2_X1 U9201 ( .A(n8243), .B(n7439), .ZN(n7424) );
  XNOR2_X1 U9202 ( .A(n7424), .B(n8059), .ZN(n7567) );
  INV_X1 U9203 ( .A(n7424), .ZN(n7425) );
  NAND2_X1 U9204 ( .A1(n7566), .A2(n4307), .ZN(n7462) );
  XNOR2_X1 U9205 ( .A(n8237), .B(n7439), .ZN(n7426) );
  XNOR2_X1 U9206 ( .A(n7426), .B(n8051), .ZN(n7461) );
  XNOR2_X1 U9207 ( .A(n8231), .B(n7439), .ZN(n7427) );
  XNOR2_X1 U9208 ( .A(n7427), .B(n8041), .ZN(n7528) );
  INV_X1 U9209 ( .A(n7427), .ZN(n7428) );
  XNOR2_X1 U9210 ( .A(n8225), .B(n7439), .ZN(n7429) );
  XNOR2_X1 U9211 ( .A(n7429), .B(n8026), .ZN(n7479) );
  AOI22_X2 U9212 ( .A1(n7480), .A2(n7479), .B1(n7430), .B2(n7429), .ZN(n7546)
         );
  XNOR2_X1 U9213 ( .A(n8219), .B(n7439), .ZN(n7431) );
  XNOR2_X1 U9214 ( .A(n7431), .B(n7987), .ZN(n7547) );
  INV_X1 U9215 ( .A(n7431), .ZN(n7432) );
  XNOR2_X1 U9216 ( .A(n7991), .B(n7439), .ZN(n7434) );
  XNOR2_X1 U9217 ( .A(n7433), .B(n7434), .ZN(n7455) );
  INV_X1 U9218 ( .A(n7433), .ZN(n7436) );
  INV_X1 U9219 ( .A(n7434), .ZN(n7435) );
  XNOR2_X1 U9220 ( .A(n8207), .B(n6650), .ZN(n7437) );
  XNOR2_X1 U9221 ( .A(n7437), .B(n7961), .ZN(n7522) );
  XNOR2_X1 U9222 ( .A(n8201), .B(n7439), .ZN(n7440) );
  XNOR2_X1 U9223 ( .A(n7440), .B(n7949), .ZN(n7499) );
  XNOR2_X1 U9224 ( .A(n7952), .B(n6655), .ZN(n7582) );
  NOR2_X1 U9225 ( .A1(n7582), .A2(n7962), .ZN(n7442) );
  INV_X1 U9226 ( .A(n7582), .ZN(n7441) );
  XNOR2_X1 U9227 ( .A(n7940), .B(n7439), .ZN(n7468) );
  XNOR2_X1 U9228 ( .A(n7468), .B(n7821), .ZN(n7470) );
  XNOR2_X1 U9229 ( .A(n7471), .B(n7470), .ZN(n7447) );
  AOI22_X1 U9230 ( .A1(n7962), .A2(n7596), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n7444) );
  NAND2_X1 U9231 ( .A1(n7939), .A2(n7600), .ZN(n7443) );
  OAI211_X1 U9232 ( .C1(n7937), .C2(n7598), .A(n7444), .B(n7443), .ZN(n7445)
         );
  AOI21_X1 U9233 ( .B1(n7940), .B2(n7587), .A(n7445), .ZN(n7446) );
  OAI21_X1 U9234 ( .B1(n7447), .B2(n7589), .A(n7446), .ZN(P2_U3154) );
  XOR2_X1 U9235 ( .A(n7449), .B(n7448), .Z(n7454) );
  AOI22_X1 U9236 ( .A1(n7573), .A2(n8094), .B1(P2_REG3_REG_14__SCAN_IN), .B2(
        P2_U3151), .ZN(n7451) );
  NAND2_X1 U9237 ( .A1(n7596), .A2(n8093), .ZN(n7450) );
  OAI211_X1 U9238 ( .C1(n8100), .C2(n7558), .A(n7451), .B(n7450), .ZN(n7452)
         );
  AOI21_X1 U9239 ( .B1(n8263), .B2(n7587), .A(n7452), .ZN(n7453) );
  OAI21_X1 U9240 ( .B1(n7454), .B2(n7589), .A(n7453), .ZN(P2_U3155) );
  XNOR2_X1 U9241 ( .A(n7455), .B(n7550), .ZN(n7460) );
  AOI22_X1 U9242 ( .A1(n8014), .A2(n7596), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n7457) );
  NAND2_X1 U9243 ( .A1(n7600), .A2(n7990), .ZN(n7456) );
  OAI211_X1 U9244 ( .C1(n7986), .C2(n7598), .A(n7457), .B(n7456), .ZN(n7458)
         );
  AOI21_X1 U9245 ( .B1(n7991), .B2(n7587), .A(n7458), .ZN(n7459) );
  OAI21_X1 U9246 ( .B1(n7460), .B2(n7589), .A(n7459), .ZN(P2_U3156) );
  XOR2_X1 U9247 ( .A(n7462), .B(n7461), .Z(n7467) );
  NAND2_X1 U9248 ( .A1(n7600), .A2(n8045), .ZN(n7464) );
  AOI22_X1 U9249 ( .A1(n7573), .A2(n8015), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3151), .ZN(n7463) );
  OAI211_X1 U9250 ( .C1(n8040), .C2(n7575), .A(n7464), .B(n7463), .ZN(n7465)
         );
  AOI21_X1 U9251 ( .B1(n8237), .B2(n7587), .A(n7465), .ZN(n7466) );
  OAI21_X1 U9252 ( .B1(n7467), .B2(n7589), .A(n7466), .ZN(P2_U3159) );
  INV_X1 U9253 ( .A(n7468), .ZN(n7469) );
  XNOR2_X1 U9254 ( .A(n7929), .B(n7439), .ZN(n7472) );
  INV_X1 U9255 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n7473) );
  OAI22_X1 U9256 ( .A1(n7948), .A2(n7575), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7473), .ZN(n7476) );
  INV_X1 U9257 ( .A(n7931), .ZN(n7474) );
  OAI22_X1 U9258 ( .A1(n7655), .A2(n7598), .B1(n7474), .B2(n7558), .ZN(n7475)
         );
  AOI211_X1 U9259 ( .C1(n7797), .C2(n7587), .A(n7476), .B(n7475), .ZN(n7477)
         );
  OAI21_X1 U9260 ( .B1(n7478), .B2(n7589), .A(n7477), .ZN(P2_U3160) );
  XOR2_X1 U9261 ( .A(n7480), .B(n7479), .Z(n7485) );
  AOI22_X1 U9262 ( .A1(n8014), .A2(n7573), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n7482) );
  NAND2_X1 U9263 ( .A1(n7600), .A2(n8018), .ZN(n7481) );
  OAI211_X1 U9264 ( .C1(n8041), .C2(n7575), .A(n7482), .B(n7481), .ZN(n7483)
         );
  AOI21_X1 U9265 ( .B1(n8225), .B2(n7587), .A(n7483), .ZN(n7484) );
  OAI21_X1 U9266 ( .B1(n7485), .B2(n7589), .A(n7484), .ZN(P2_U3163) );
  OAI21_X1 U9267 ( .B1(n7825), .B2(n7412), .A(n7486), .ZN(n7561) );
  XNOR2_X1 U9268 ( .A(n7487), .B(n4501), .ZN(n7562) );
  NOR2_X1 U9269 ( .A1(n7561), .A2(n7562), .ZN(n7560) );
  NOR2_X1 U9270 ( .A1(n7560), .A2(n7488), .ZN(n7489) );
  XOR2_X1 U9271 ( .A(n7490), .B(n7489), .Z(n7497) );
  NAND2_X1 U9272 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n9807) );
  INV_X1 U9273 ( .A(n9807), .ZN(n7492) );
  NOR2_X1 U9274 ( .A1(n7575), .A2(n4501), .ZN(n7491) );
  AOI211_X1 U9275 ( .C1(n7573), .C2(n8093), .A(n7492), .B(n7491), .ZN(n7493)
         );
  OAI21_X1 U9276 ( .B1(n7494), .B2(n7558), .A(n7493), .ZN(n7495) );
  AOI21_X1 U9277 ( .B1(n9965), .B2(n7587), .A(n7495), .ZN(n7496) );
  OAI21_X1 U9278 ( .B1(n7497), .B2(n7589), .A(n7496), .ZN(P2_U3164) );
  XOR2_X1 U9279 ( .A(n7499), .B(n7498), .Z(n7504) );
  AOI22_X1 U9280 ( .A1(n7962), .A2(n7573), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n7501) );
  NAND2_X1 U9281 ( .A1(n7600), .A2(n7966), .ZN(n7500) );
  OAI211_X1 U9282 ( .C1(n7986), .C2(n7575), .A(n7501), .B(n7500), .ZN(n7502)
         );
  AOI21_X1 U9283 ( .B1(n8201), .B2(n7587), .A(n7502), .ZN(n7503) );
  OAI21_X1 U9284 ( .B1(n7504), .B2(n7589), .A(n7503), .ZN(P2_U3165) );
  INV_X1 U9285 ( .A(n8250), .ZN(n7513) );
  OAI211_X1 U9286 ( .C1(n7507), .C2(n7506), .A(n7505), .B(n7591), .ZN(n7512)
         );
  INV_X1 U9287 ( .A(n7508), .ZN(n8074) );
  NAND2_X1 U9288 ( .A1(n7596), .A2(n8094), .ZN(n7509) );
  NAND2_X1 U9289 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n9871) );
  OAI211_X1 U9290 ( .C1(n7576), .C2(n7598), .A(n7509), .B(n9871), .ZN(n7510)
         );
  AOI21_X1 U9291 ( .B1(n8074), .B2(n7600), .A(n7510), .ZN(n7511) );
  OAI211_X1 U9292 ( .C1(n7513), .C2(n7603), .A(n7512), .B(n7511), .ZN(P2_U3166) );
  AOI21_X1 U9293 ( .B1(n7515), .B2(n7514), .A(n7569), .ZN(n7520) );
  AOI22_X1 U9294 ( .A1(n7573), .A2(n8059), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3151), .ZN(n7517) );
  NAND2_X1 U9295 ( .A1(n7596), .A2(n8058), .ZN(n7516) );
  OAI211_X1 U9296 ( .C1(n8061), .C2(n7558), .A(n7517), .B(n7516), .ZN(n7518)
         );
  AOI21_X1 U9297 ( .B1(n8143), .B2(n7587), .A(n7518), .ZN(n7519) );
  OAI21_X1 U9298 ( .B1(n7520), .B2(n7589), .A(n7519), .ZN(P2_U3168) );
  XOR2_X1 U9299 ( .A(n7522), .B(n7521), .Z(n7527) );
  AOI22_X1 U9300 ( .A1(n7975), .A2(n7573), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n7524) );
  NAND2_X1 U9301 ( .A1(n7600), .A2(n7979), .ZN(n7523) );
  OAI211_X1 U9302 ( .C1(n7550), .C2(n7575), .A(n7524), .B(n7523), .ZN(n7525)
         );
  AOI21_X1 U9303 ( .B1(n8207), .B2(n7587), .A(n7525), .ZN(n7526) );
  OAI21_X1 U9304 ( .B1(n7527), .B2(n7589), .A(n7526), .ZN(P2_U3169) );
  XOR2_X1 U9305 ( .A(n7529), .B(n7528), .Z(n7535) );
  NAND2_X1 U9306 ( .A1(n7600), .A2(n8029), .ZN(n7531) );
  AOI22_X1 U9307 ( .A1(n7573), .A2(n8026), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n7530) );
  OAI211_X1 U9308 ( .C1(n7532), .C2(n7575), .A(n7531), .B(n7530), .ZN(n7533)
         );
  AOI21_X1 U9309 ( .B1(n8231), .B2(n7587), .A(n7533), .ZN(n7534) );
  OAI21_X1 U9310 ( .B1(n7535), .B2(n7589), .A(n7534), .ZN(P2_U3173) );
  XNOR2_X1 U9311 ( .A(n7536), .B(n8093), .ZN(n7537) );
  XNOR2_X1 U9312 ( .A(n7538), .B(n7537), .ZN(n7545) );
  NAND2_X1 U9313 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n9822) );
  INV_X1 U9314 ( .A(n9822), .ZN(n7540) );
  NOR2_X1 U9315 ( .A1(n7598), .A2(n8082), .ZN(n7539) );
  AOI211_X1 U9316 ( .C1(n7596), .C2(n7823), .A(n7540), .B(n7539), .ZN(n7541)
         );
  OAI21_X1 U9317 ( .B1(n7542), .B2(n7558), .A(n7541), .ZN(n7543) );
  AOI21_X1 U9318 ( .B1(n7659), .B2(n7587), .A(n7543), .ZN(n7544) );
  OAI21_X1 U9319 ( .B1(n7545), .B2(n7589), .A(n7544), .ZN(P2_U3174) );
  XOR2_X1 U9320 ( .A(n7547), .B(n7546), .Z(n7553) );
  NAND2_X1 U9321 ( .A1(n7600), .A2(n7996), .ZN(n7549) );
  AOI22_X1 U9322 ( .A1(n7596), .A2(n8026), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n7548) );
  OAI211_X1 U9323 ( .C1(n7550), .C2(n7598), .A(n7549), .B(n7548), .ZN(n7551)
         );
  AOI21_X1 U9324 ( .B1(n8219), .B2(n7587), .A(n7551), .ZN(n7552) );
  OAI21_X1 U9325 ( .B1(n7553), .B2(n7589), .A(n7552), .ZN(P2_U3175) );
  NAND2_X1 U9326 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n9791) );
  INV_X1 U9327 ( .A(n9791), .ZN(n7554) );
  AOI21_X1 U9328 ( .B1(n7573), .B2(n7823), .A(n7554), .ZN(n7557) );
  OR2_X1 U9329 ( .A1(n7575), .A2(n7555), .ZN(n7556) );
  OAI211_X1 U9330 ( .C1(n7559), .C2(n7558), .A(n7557), .B(n7556), .ZN(n7564)
         );
  AOI211_X1 U9331 ( .C1(n7562), .C2(n7561), .A(n7589), .B(n7560), .ZN(n7563)
         );
  AOI211_X1 U9332 ( .C1(n9959), .C2(n7587), .A(n7564), .B(n7563), .ZN(n7565)
         );
  INV_X1 U9333 ( .A(n7565), .ZN(P2_U3176) );
  INV_X1 U9334 ( .A(n8243), .ZN(n7580) );
  INV_X1 U9335 ( .A(n7566), .ZN(n7571) );
  NOR3_X1 U9336 ( .A1(n7569), .A2(n7568), .A3(n7567), .ZN(n7570) );
  OAI21_X1 U9337 ( .B1(n7571), .B2(n7570), .A(n7591), .ZN(n7579) );
  INV_X1 U9338 ( .A(n7572), .ZN(n8054) );
  AOI22_X1 U9339 ( .A1(n7573), .A2(n8051), .B1(P2_REG3_REG_18__SCAN_IN), .B2(
        P2_U3151), .ZN(n7574) );
  OAI21_X1 U9340 ( .B1(n7576), .B2(n7575), .A(n7574), .ZN(n7577) );
  AOI21_X1 U9341 ( .B1(n8054), .B2(n7600), .A(n7577), .ZN(n7578) );
  OAI211_X1 U9342 ( .C1(n7580), .C2(n7603), .A(n7579), .B(n7578), .ZN(P2_U3178) );
  XNOR2_X1 U9343 ( .A(n7582), .B(n7962), .ZN(n7583) );
  XNOR2_X1 U9344 ( .A(n7581), .B(n7583), .ZN(n7590) );
  AOI22_X1 U9345 ( .A1(n7975), .A2(n7596), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n7585) );
  NAND2_X1 U9346 ( .A1(n7953), .A2(n7600), .ZN(n7584) );
  OAI211_X1 U9347 ( .C1(n7948), .C2(n7598), .A(n7585), .B(n7584), .ZN(n7586)
         );
  AOI21_X1 U9348 ( .B1(n7952), .B2(n7587), .A(n7586), .ZN(n7588) );
  OAI21_X1 U9349 ( .B1(n7590), .B2(n7589), .A(n7588), .ZN(P2_U3180) );
  OAI211_X1 U9350 ( .C1(n7594), .C2(n7593), .A(n7592), .B(n7591), .ZN(n7602)
         );
  INV_X1 U9351 ( .A(n7595), .ZN(n8085) );
  NAND2_X1 U9352 ( .A1(n7596), .A2(n7822), .ZN(n7597) );
  NAND2_X1 U9353 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9854) );
  OAI211_X1 U9354 ( .C1(n8081), .C2(n7598), .A(n7597), .B(n9854), .ZN(n7599)
         );
  AOI21_X1 U9355 ( .B1(n8085), .B2(n7600), .A(n7599), .ZN(n7601) );
  OAI211_X1 U9356 ( .C1(n7604), .C2(n7603), .A(n7602), .B(n7601), .ZN(P2_U3181) );
  INV_X1 U9357 ( .A(n7605), .ZN(n7810) );
  NAND2_X1 U9358 ( .A1(n7607), .A2(n5387), .ZN(n7611) );
  OR2_X1 U9359 ( .A1(n7609), .A2(n7608), .ZN(n7610) );
  INV_X1 U9360 ( .A(n7819), .ZN(n7612) );
  INV_X1 U9361 ( .A(n7800), .ZN(n7623) );
  NAND2_X1 U9362 ( .A1(n8183), .A2(n7612), .ZN(n7795) );
  AND2_X1 U9363 ( .A1(n7795), .A2(n7613), .ZN(n7794) );
  INV_X1 U9364 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n7618) );
  NAND2_X1 U9365 ( .A1(n4261), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n7617) );
  INV_X1 U9366 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n7614) );
  OR2_X1 U9367 ( .A1(n7615), .A2(n7614), .ZN(n7616) );
  OAI211_X1 U9368 ( .C1(n4908), .C2(n7618), .A(n7617), .B(n7616), .ZN(n7619)
         );
  INV_X1 U9369 ( .A(n7619), .ZN(n7620) );
  NAND2_X1 U9370 ( .A1(n7621), .A2(n7620), .ZN(n7917) );
  OAI21_X1 U9371 ( .B1(n8183), .B2(n7917), .A(n8180), .ZN(n7622) );
  NAND2_X1 U9372 ( .A1(n8180), .A2(n7917), .ZN(n7803) );
  INV_X1 U9373 ( .A(n7803), .ZN(n7651) );
  INV_X1 U9374 ( .A(n7799), .ZN(n7796) );
  INV_X1 U9375 ( .A(n7784), .ZN(n7625) );
  XNOR2_X1 U9376 ( .A(n7952), .B(n7938), .ZN(n7951) );
  INV_X1 U9377 ( .A(n7968), .ZN(n7649) );
  INV_X1 U9378 ( .A(n7626), .ZN(n7771) );
  INV_X1 U9379 ( .A(n8024), .ZN(n7645) );
  NOR2_X1 U9380 ( .A1(n7628), .A2(n7627), .ZN(n7730) );
  NAND4_X1 U9381 ( .A1(n7629), .A2(n7667), .A3(n8156), .A4(n7678), .ZN(n7631)
         );
  NOR2_X1 U9382 ( .A1(n7631), .A2(n7630), .ZN(n7634) );
  NAND4_X1 U9383 ( .A1(n7634), .A2(n7701), .A3(n7633), .A4(n7632), .ZN(n7638)
         );
  NOR4_X1 U9384 ( .A1(n7638), .A2(n7637), .A3(n7636), .A4(n7635), .ZN(n7639)
         );
  NAND3_X1 U9385 ( .A1(n7640), .A2(n7730), .A3(n7639), .ZN(n7641) );
  OR2_X1 U9386 ( .A1(n7641), .A2(n8091), .ZN(n7642) );
  OR4_X1 U9387 ( .A1(n8078), .A2(n7744), .A3(n7642), .A4(n7741), .ZN(n7643) );
  NOR2_X1 U9388 ( .A1(n8050), .A2(n7643), .ZN(n7644) );
  NAND3_X1 U9389 ( .A1(n7645), .A2(n8032), .A3(n7644), .ZN(n7646) );
  NOR2_X1 U9390 ( .A1(n7646), .A2(n8009), .ZN(n7647) );
  INV_X1 U9391 ( .A(n7999), .ZN(n7994) );
  NAND4_X1 U9392 ( .A1(n7973), .A2(n7983), .A3(n7647), .A4(n7994), .ZN(n7648)
         );
  OAI22_X1 U9393 ( .A1(n7653), .A2(n7652), .B1(n8180), .B2(n7917), .ZN(n7809)
         );
  NAND2_X1 U9394 ( .A1(n7654), .A2(n7801), .ZN(n7656) );
  NOR2_X1 U9395 ( .A1(n7655), .A2(n7781), .ZN(n7925) );
  AOI21_X1 U9396 ( .B1(n7800), .B2(n7656), .A(n7925), .ZN(n7791) );
  MUX2_X1 U9397 ( .A(n7820), .B(n7797), .S(n7781), .Z(n7792) );
  INV_X1 U9398 ( .A(n7758), .ZN(n7658) );
  NOR2_X1 U9399 ( .A1(n7658), .A2(n7657), .ZN(n7750) );
  MUX2_X1 U9400 ( .A(n8093), .B(n7659), .S(n7801), .Z(n7733) );
  INV_X1 U9401 ( .A(n7733), .ZN(n7736) );
  INV_X1 U9402 ( .A(n7660), .ZN(n7735) );
  AOI22_X1 U9403 ( .A1(n7664), .A2(n7663), .B1(n7662), .B2(n7661), .ZN(n7669)
         );
  INV_X1 U9404 ( .A(n7665), .ZN(n7674) );
  NAND3_X1 U9405 ( .A1(n7667), .A2(n7801), .A3(n7666), .ZN(n7668) );
  OAI211_X1 U9406 ( .C1(n7669), .C2(n7674), .A(n8156), .B(n7668), .ZN(n7675)
         );
  INV_X1 U9407 ( .A(n7670), .ZN(n7672) );
  OAI211_X1 U9408 ( .C1(n7675), .C2(n7672), .A(n7671), .B(n7693), .ZN(n7677)
         );
  NAND2_X1 U9409 ( .A1(n8162), .A2(n9912), .ZN(n7680) );
  OAI211_X1 U9410 ( .C1(n7675), .C2(n7674), .A(n7680), .B(n7673), .ZN(n7676)
         );
  MUX2_X1 U9411 ( .A(n7677), .B(n7676), .S(n7801), .Z(n7679) );
  NAND2_X1 U9412 ( .A1(n7679), .A2(n7678), .ZN(n7697) );
  INV_X1 U9413 ( .A(n7680), .ZN(n7682) );
  OAI211_X1 U9414 ( .C1(n7697), .C2(n7682), .A(n7698), .B(n7681), .ZN(n7687)
         );
  INV_X1 U9415 ( .A(n7695), .ZN(n7684) );
  OAI21_X1 U9416 ( .B1(n7685), .B2(n7684), .A(n7683), .ZN(n7686) );
  INV_X1 U9417 ( .A(n7711), .ZN(n7689) );
  NAND2_X1 U9418 ( .A1(n7690), .A2(n7689), .ZN(n7691) );
  NAND2_X1 U9419 ( .A1(n7691), .A2(n7801), .ZN(n7707) );
  AND2_X1 U9420 ( .A1(n7702), .A2(n7692), .ZN(n7712) );
  AND2_X1 U9421 ( .A1(n7707), .A2(n7712), .ZN(n7709) );
  INV_X1 U9422 ( .A(n7693), .ZN(n7696) );
  OAI211_X1 U9423 ( .C1(n7697), .C2(n7696), .A(n7695), .B(n7694), .ZN(n7699)
         );
  NAND3_X1 U9424 ( .A1(n7699), .A2(n7698), .A3(n7801), .ZN(n7700) );
  INV_X1 U9425 ( .A(n7702), .ZN(n7706) );
  INV_X1 U9426 ( .A(n7720), .ZN(n7705) );
  INV_X1 U9427 ( .A(n7719), .ZN(n7703) );
  OAI33_X1 U9428 ( .A1(n7707), .A2(n7706), .A3(n7705), .B1(n7801), .B2(n7704), 
        .B3(n7703), .ZN(n7718) );
  INV_X1 U9429 ( .A(n7708), .ZN(n7710) );
  OAI21_X1 U9430 ( .B1(n7711), .B2(n7710), .A(n7709), .ZN(n7717) );
  INV_X1 U9431 ( .A(n7712), .ZN(n7715) );
  NAND2_X1 U9432 ( .A1(n7713), .A2(n7801), .ZN(n7714) );
  NOR2_X1 U9433 ( .A1(n7715), .A2(n7714), .ZN(n7716) );
  AOI22_X1 U9434 ( .A1(n7718), .A2(n7717), .B1(n7716), .B2(n7720), .ZN(n7722)
         );
  MUX2_X1 U9435 ( .A(n7720), .B(n7719), .S(n7801), .Z(n7721) );
  INV_X1 U9436 ( .A(n7723), .ZN(n7724) );
  AOI21_X1 U9437 ( .B1(n7726), .B2(n7725), .A(n7724), .ZN(n7728) );
  NOR2_X1 U9438 ( .A1(n7728), .A2(n7730), .ZN(n7727) );
  MUX2_X1 U9439 ( .A(n7728), .B(n7727), .S(n7801), .Z(n7729) );
  AOI21_X1 U9440 ( .B1(n7731), .B2(n7730), .A(n7729), .ZN(n7732) );
  MUX2_X1 U9441 ( .A(n7738), .B(n7737), .S(n7781), .Z(n7739) );
  MUX2_X1 U9442 ( .A(n7742), .B(n4305), .S(n7801), .Z(n7743) );
  MUX2_X1 U9443 ( .A(n7746), .B(n7745), .S(n7801), .Z(n7747) );
  NAND3_X1 U9444 ( .A1(n7748), .A2(n5185), .A3(n7747), .ZN(n7753) );
  INV_X1 U9445 ( .A(n7755), .ZN(n7756) );
  OAI21_X1 U9446 ( .B1(n4339), .B2(n7756), .A(n7759), .ZN(n7762) );
  INV_X1 U9447 ( .A(n8219), .ZN(n7763) );
  MUX2_X1 U9448 ( .A(n7763), .B(n7987), .S(n7781), .Z(n7767) );
  INV_X1 U9449 ( .A(n7764), .ZN(n7766) );
  NAND3_X1 U9450 ( .A1(n7772), .A2(n7773), .A3(n7768), .ZN(n7769) );
  NAND3_X1 U9451 ( .A1(n7772), .A2(n7771), .A3(n7770), .ZN(n7774) );
  NOR2_X1 U9452 ( .A1(n7938), .A2(n7781), .ZN(n7775) );
  AOI21_X1 U9453 ( .B1(n7952), .B2(n7781), .A(n7775), .ZN(n7785) );
  MUX2_X1 U9454 ( .A(n7962), .B(n7952), .S(n7801), .Z(n7783) );
  INV_X1 U9455 ( .A(n7941), .ZN(n7779) );
  MUX2_X1 U9456 ( .A(n7777), .B(n7776), .S(n7801), .Z(n7778) );
  OAI211_X1 U9457 ( .C1(n7785), .C2(n7783), .A(n7779), .B(n7778), .ZN(n7780)
         );
  INV_X1 U9458 ( .A(n7940), .ZN(n8192) );
  AOI21_X1 U9459 ( .B1(n7948), .B2(n7801), .A(n8192), .ZN(n7789) );
  AOI21_X1 U9460 ( .B1(n7781), .B2(n7821), .A(n7940), .ZN(n7788) );
  INV_X1 U9461 ( .A(n7782), .ZN(n7786) );
  NAND4_X1 U9462 ( .A1(n7786), .A2(n7785), .A3(n7784), .A4(n7783), .ZN(n7787)
         );
  OAI21_X1 U9463 ( .B1(n7789), .B2(n7788), .A(n7787), .ZN(n7790) );
  AOI21_X1 U9464 ( .B1(n4493), .B2(n7792), .A(n7793), .ZN(n7798) );
  NAND2_X1 U9465 ( .A1(n7793), .A2(n7792), .ZN(n7802) );
  OAI211_X1 U9466 ( .C1(n7798), .C2(n7820), .A(n7794), .B(n7802), .ZN(n7808)
         );
  OAI21_X1 U9467 ( .B1(n7796), .B2(n7801), .A(n7795), .ZN(n7807) );
  NOR2_X1 U9468 ( .A1(n7798), .A2(n7797), .ZN(n7806) );
  NAND4_X1 U9469 ( .A1(n7802), .A2(n7801), .A3(n7800), .A4(n7799), .ZN(n7805)
         );
  NOR3_X1 U9470 ( .A1(n7813), .A2(n7812), .A3(n7811), .ZN(n7816) );
  OAI21_X1 U9471 ( .B1(n7817), .B2(n7814), .A(P2_B_REG_SCAN_IN), .ZN(n7815) );
  OAI22_X1 U9472 ( .A1(n7818), .A2(n7817), .B1(n7816), .B2(n7815), .ZN(
        P2_U3296) );
  MUX2_X1 U9473 ( .A(n7917), .B(P2_DATAO_REG_31__SCAN_IN), .S(n7833), .Z(
        P2_U3522) );
  MUX2_X1 U9474 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n7819), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U9475 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n7820), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9476 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n7821), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9477 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n7962), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U9478 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n7975), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9479 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n7961), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9480 ( .A(n8000), .B(P2_DATAO_REG_23__SCAN_IN), .S(n7833), .Z(
        P2_U3514) );
  MUX2_X1 U9481 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8014), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9482 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8026), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9483 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8015), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9484 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8051), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9485 ( .A(n8059), .B(P2_DATAO_REG_18__SCAN_IN), .S(n7833), .Z(
        P2_U3509) );
  MUX2_X1 U9486 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8071), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9487 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8058), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9488 ( .A(n8094), .B(P2_DATAO_REG_15__SCAN_IN), .S(n7833), .Z(
        P2_U3506) );
  MUX2_X1 U9489 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n7822), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U9490 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8093), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U9491 ( .A(n7823), .B(P2_DATAO_REG_12__SCAN_IN), .S(n7833), .Z(
        P2_U3503) );
  MUX2_X1 U9492 ( .A(n7824), .B(P2_DATAO_REG_11__SCAN_IN), .S(n7833), .Z(
        P2_U3502) );
  MUX2_X1 U9493 ( .A(n7825), .B(P2_DATAO_REG_10__SCAN_IN), .S(n7833), .Z(
        P2_U3501) );
  MUX2_X1 U9494 ( .A(n7826), .B(P2_DATAO_REG_9__SCAN_IN), .S(n7833), .Z(
        P2_U3500) );
  MUX2_X1 U9495 ( .A(n7827), .B(P2_DATAO_REG_8__SCAN_IN), .S(n7833), .Z(
        P2_U3499) );
  MUX2_X1 U9496 ( .A(n7828), .B(P2_DATAO_REG_7__SCAN_IN), .S(n7833), .Z(
        P2_U3498) );
  MUX2_X1 U9497 ( .A(n7829), .B(P2_DATAO_REG_6__SCAN_IN), .S(n7833), .Z(
        P2_U3497) );
  MUX2_X1 U9498 ( .A(n7830), .B(P2_DATAO_REG_5__SCAN_IN), .S(n7833), .Z(
        P2_U3496) );
  MUX2_X1 U9499 ( .A(n7831), .B(P2_DATAO_REG_4__SCAN_IN), .S(n7833), .Z(
        P2_U3495) );
  MUX2_X1 U9500 ( .A(n8162), .B(P2_DATAO_REG_3__SCAN_IN), .S(n7833), .Z(
        P2_U3494) );
  MUX2_X1 U9501 ( .A(n7832), .B(P2_DATAO_REG_2__SCAN_IN), .S(n7833), .Z(
        P2_U3493) );
  MUX2_X1 U9502 ( .A(n4867), .B(P2_DATAO_REG_1__SCAN_IN), .S(n7833), .Z(
        P2_U3492) );
  MUX2_X1 U9503 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n7834), .S(P2_U3893), .Z(
        P2_U3491) );
  NAND2_X1 U9504 ( .A1(n7836), .A2(n7835), .ZN(n7837) );
  NAND2_X1 U9505 ( .A1(n7838), .A2(n7837), .ZN(n7841) );
  XNOR2_X1 U9506 ( .A(n7839), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n7840) );
  AOI22_X1 U9507 ( .A1(n9754), .A2(n7841), .B1(n9884), .B2(n7840), .ZN(n7849)
         );
  AOI22_X1 U9508 ( .A1(n9875), .A2(n7842), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        P2_U3151), .ZN(n7848) );
  OAI211_X1 U9509 ( .C1(n7845), .C2(n7844), .A(n7843), .B(n9883), .ZN(n7847)
         );
  NAND2_X1 U9510 ( .A1(n9874), .A2(P2_ADDR_REG_1__SCAN_IN), .ZN(n7846) );
  NAND4_X1 U9511 ( .A1(n7849), .A2(n7848), .A3(n7847), .A4(n7846), .ZN(
        P2_U3183) );
  AOI22_X1 U9512 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n7911), .B1(n9514), .B2(
        n8140), .ZN(n9505) );
  AOI22_X1 U9513 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n7907), .B1(n9857), .B2(
        n9050), .ZN(n9860) );
  AOI22_X1 U9514 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n7904), .B1(n9825), .B2(
        n8151), .ZN(n9828) );
  AOI22_X1 U9515 ( .A1(n9794), .A2(n5077), .B1(P2_REG1_REG_12__SCAN_IN), .B2(
        n7900), .ZN(n9797) );
  NAND2_X1 U9516 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n7895), .ZN(n7853) );
  AOI22_X1 U9517 ( .A1(n9761), .A2(n5038), .B1(P2_REG1_REG_10__SCAN_IN), .B2(
        n7895), .ZN(n9767) );
  AOI22_X1 U9518 ( .A1(n7851), .A2(P2_REG1_REG_9__SCAN_IN), .B1(n7892), .B2(
        n7850), .ZN(n7852) );
  INV_X1 U9519 ( .A(n7852), .ZN(n9766) );
  NAND2_X1 U9520 ( .A1(n9767), .A2(n9766), .ZN(n9765) );
  NAND2_X1 U9521 ( .A1(n7853), .A2(n9765), .ZN(n7854) );
  NAND2_X1 U9522 ( .A1(n7854), .A2(n7898), .ZN(n7855) );
  XNOR2_X1 U9523 ( .A(n7854), .B(n9778), .ZN(n9780) );
  NAND2_X1 U9524 ( .A1(P2_REG1_REG_11__SCAN_IN), .A2(n9780), .ZN(n9779) );
  NAND2_X1 U9525 ( .A1(n7855), .A2(n9779), .ZN(n9796) );
  NAND2_X1 U9526 ( .A1(n9797), .A2(n9796), .ZN(n9795) );
  OAI21_X1 U9527 ( .B1(n9794), .B2(n5077), .A(n9795), .ZN(n7856) );
  NAND2_X1 U9528 ( .A1(n7869), .A2(n7856), .ZN(n7857) );
  NAND2_X1 U9529 ( .A1(n7857), .A2(n9811), .ZN(n9827) );
  NAND2_X1 U9530 ( .A1(n9828), .A2(n9827), .ZN(n9826) );
  OAI21_X1 U9531 ( .B1(n9825), .B2(n8151), .A(n9826), .ZN(n7858) );
  NAND2_X1 U9532 ( .A1(n7866), .A2(n7858), .ZN(n7859) );
  NAND2_X1 U9533 ( .A1(n7859), .A2(n9842), .ZN(n9859) );
  NAND2_X1 U9534 ( .A1(n9860), .A2(n9859), .ZN(n9858) );
  OAI21_X1 U9535 ( .B1(n9857), .B2(n9050), .A(n9858), .ZN(n7860) );
  NAND2_X1 U9536 ( .A1(n7864), .A2(n7860), .ZN(n7861) );
  NAND2_X1 U9537 ( .A1(n7861), .A2(n9877), .ZN(n9504) );
  XNOR2_X1 U9538 ( .A(n7888), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n7889) );
  XNOR2_X1 U9539 ( .A(n7862), .B(n7889), .ZN(n7915) );
  XNOR2_X1 U9540 ( .A(n7885), .B(n7864), .ZN(n9881) );
  OR2_X1 U9541 ( .A1(n7865), .A2(n7907), .ZN(n7884) );
  XNOR2_X1 U9542 ( .A(n7865), .B(n9857), .ZN(n9863) );
  OR2_X1 U9543 ( .A1(n7867), .A2(n7866), .ZN(n7883) );
  XNOR2_X1 U9544 ( .A(n7867), .B(n9841), .ZN(n9846) );
  OR2_X1 U9545 ( .A1(n7868), .A2(n7904), .ZN(n7882) );
  XNOR2_X1 U9546 ( .A(n7868), .B(n9825), .ZN(n9831) );
  OR2_X1 U9547 ( .A1(n7870), .A2(n7869), .ZN(n7881) );
  XNOR2_X1 U9548 ( .A(n7870), .B(n9810), .ZN(n9815) );
  OR2_X1 U9549 ( .A1(n7871), .A2(n7900), .ZN(n7880) );
  XNOR2_X1 U9550 ( .A(n7871), .B(n9794), .ZN(n9800) );
  OR2_X1 U9551 ( .A1(n7872), .A2(n7898), .ZN(n7879) );
  XNOR2_X1 U9552 ( .A(n7872), .B(n9778), .ZN(n9783) );
  OR2_X1 U9553 ( .A1(n7873), .A2(n7895), .ZN(n7878) );
  XNOR2_X1 U9554 ( .A(n7873), .B(n9761), .ZN(n9763) );
  INV_X1 U9555 ( .A(n7874), .ZN(n7877) );
  OAI22_X1 U9556 ( .A1(n7877), .A2(n7876), .B1(n7875), .B2(n7892), .ZN(n9764)
         );
  NAND2_X1 U9557 ( .A1(n9763), .A2(n9764), .ZN(n9762) );
  NAND2_X1 U9558 ( .A1(n7878), .A2(n9762), .ZN(n9782) );
  NAND2_X1 U9559 ( .A1(n9783), .A2(n9782), .ZN(n9781) );
  NAND2_X1 U9560 ( .A1(n7879), .A2(n9781), .ZN(n9799) );
  NAND2_X1 U9561 ( .A1(n9800), .A2(n9799), .ZN(n9798) );
  NAND2_X1 U9562 ( .A1(n7880), .A2(n9798), .ZN(n9814) );
  NAND2_X1 U9563 ( .A1(n9815), .A2(n9814), .ZN(n9813) );
  NAND2_X1 U9564 ( .A1(n7881), .A2(n9813), .ZN(n9830) );
  NAND2_X1 U9565 ( .A1(n9863), .A2(n9862), .ZN(n9861) );
  NAND2_X1 U9566 ( .A1(n7887), .A2(n7886), .ZN(n9509) );
  NOR2_X1 U9567 ( .A1(n7887), .A2(n7886), .ZN(n9507) );
  XNOR2_X1 U9568 ( .A(n7888), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n7891) );
  NOR2_X1 U9569 ( .A1(n9720), .A2(n4734), .ZN(n7914) );
  NAND2_X1 U9570 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n7895), .ZN(n7894) );
  OAI21_X1 U9571 ( .B1(n7895), .B2(P2_REG2_REG_10__SCAN_IN), .A(n7894), .ZN(
        n9771) );
  NOR2_X1 U9572 ( .A1(n9772), .A2(n9771), .ZN(n9770) );
  AOI21_X1 U9573 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n7895), .A(n9770), .ZN(
        n7896) );
  INV_X1 U9574 ( .A(n7896), .ZN(n7897) );
  NAND2_X1 U9575 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n7900), .ZN(n7899) );
  OAI21_X1 U9576 ( .B1(n7900), .B2(P2_REG2_REG_12__SCAN_IN), .A(n7899), .ZN(
        n9804) );
  NOR2_X1 U9577 ( .A1(n9810), .A2(n7901), .ZN(n7902) );
  XNOR2_X1 U9578 ( .A(n9810), .B(n7901), .ZN(n9819) );
  XNOR2_X1 U9579 ( .A(n9825), .B(n7903), .ZN(n9835) );
  XNOR2_X1 U9580 ( .A(n9841), .B(n7905), .ZN(n9851) );
  NOR2_X1 U9581 ( .A1(n7907), .A2(n8073), .ZN(n7906) );
  AOI21_X1 U9582 ( .B1(n8073), .B2(n7907), .A(n7906), .ZN(n9867) );
  NOR2_X1 U9583 ( .A1(n9876), .A2(n7908), .ZN(n7909) );
  XNOR2_X1 U9584 ( .A(n9876), .B(n7908), .ZN(n9888) );
  NOR2_X1 U9585 ( .A1(n9887), .A2(n9888), .ZN(n9886) );
  NOR2_X1 U9586 ( .A1(n7911), .A2(n8053), .ZN(n7910) );
  AOI21_X1 U9587 ( .B1(n8053), .B2(n7911), .A(n7910), .ZN(n9517) );
  NOR2_X1 U9588 ( .A1(n9518), .A2(n9517), .ZN(n9516) );
  AOI21_X1 U9589 ( .B1(n7911), .B2(P2_REG2_REG_18__SCAN_IN), .A(n9516), .ZN(
        n7912) );
  AOI21_X1 U9590 ( .B1(n8181), .B2(n8098), .A(n7918), .ZN(n7921) );
  NAND2_X1 U9591 ( .A1(n9907), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n7919) );
  OAI211_X1 U9592 ( .C1(n8180), .C2(n7955), .A(n7921), .B(n7919), .ZN(P2_U3202) );
  INV_X1 U9593 ( .A(n8183), .ZN(n7922) );
  NAND2_X1 U9594 ( .A1(n9907), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n7920) );
  OAI211_X1 U9595 ( .C1(n7922), .C2(n7955), .A(n7921), .B(n7920), .ZN(P2_U3203) );
  XNOR2_X1 U9596 ( .A(n7923), .B(n7929), .ZN(n7928) );
  NAND2_X1 U9597 ( .A1(n7925), .A2(n7924), .ZN(n7926) );
  OAI21_X1 U9598 ( .B1(n7948), .B2(n8164), .A(n7926), .ZN(n7927) );
  AOI21_X1 U9599 ( .B1(n7928), .B2(n8167), .A(n7927), .ZN(n8112) );
  XNOR2_X1 U9600 ( .A(n7930), .B(n4742), .ZN(n8110) );
  AOI22_X1 U9601 ( .A1(n7931), .A2(n8102), .B1(n9907), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n7932) );
  OAI21_X1 U9602 ( .B1(n8190), .B2(n7955), .A(n7932), .ZN(n7933) );
  AOI21_X1 U9603 ( .B1(n8110), .B2(n8065), .A(n7933), .ZN(n7934) );
  OAI21_X1 U9604 ( .B1(n8112), .B2(n9907), .A(n7934), .ZN(P2_U3205) );
  XNOR2_X1 U9605 ( .A(n7935), .B(n7941), .ZN(n7936) );
  OAI222_X1 U9606 ( .A1(n8164), .A2(n7938), .B1(n8080), .B2(n7937), .C1(n7936), 
        .C2(n8037), .ZN(n8191) );
  AOI21_X1 U9607 ( .B1(n8102), .B2(n7939), .A(n8191), .ZN(n7945) );
  AOI22_X1 U9608 ( .A1(n7940), .A2(n8086), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n9907), .ZN(n7944) );
  XNOR2_X1 U9609 ( .A(n7942), .B(n7941), .ZN(n8115) );
  NAND2_X1 U9610 ( .A1(n8115), .A2(n8065), .ZN(n7943) );
  OAI211_X1 U9611 ( .C1(n7945), .C2(n9907), .A(n7944), .B(n7943), .ZN(P2_U3206) );
  OAI222_X1 U9612 ( .A1(n8164), .A2(n7949), .B1(n8080), .B2(n7948), .C1(n7947), 
        .C2(n8037), .ZN(n8118) );
  INV_X1 U9613 ( .A(n8118), .ZN(n7958) );
  XNOR2_X1 U9614 ( .A(n7950), .B(n7951), .ZN(n8119) );
  INV_X1 U9615 ( .A(n7952), .ZN(n8198) );
  AOI22_X1 U9616 ( .A1(n7953), .A2(n8102), .B1(n9907), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n7954) );
  OAI21_X1 U9617 ( .B1(n8198), .B2(n7955), .A(n7954), .ZN(n7956) );
  AOI21_X1 U9618 ( .B1(n8119), .B2(n8065), .A(n7956), .ZN(n7957) );
  OAI21_X1 U9619 ( .B1(n7958), .B2(n9907), .A(n7957), .ZN(P2_U3207) );
  INV_X1 U9620 ( .A(n8201), .ZN(n7959) );
  NOR2_X1 U9621 ( .A1(n7959), .A2(n8096), .ZN(n7965) );
  XNOR2_X1 U9622 ( .A(n7960), .B(n7968), .ZN(n7963) );
  AOI222_X1 U9623 ( .A1(n8167), .A2(n7963), .B1(n7962), .B2(n8161), .C1(n7961), 
        .C2(n8092), .ZN(n8199) );
  INV_X1 U9624 ( .A(n8199), .ZN(n7964) );
  AOI211_X1 U9625 ( .C1(n8102), .C2(n7966), .A(n7965), .B(n7964), .ZN(n7971)
         );
  INV_X1 U9626 ( .A(n8204), .ZN(n7969) );
  AOI22_X1 U9627 ( .A1(n7969), .A2(n8065), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n9907), .ZN(n7970) );
  OAI21_X1 U9628 ( .B1(n7971), .B2(n9907), .A(n7970), .ZN(P2_U3208) );
  XOR2_X1 U9629 ( .A(n7973), .B(n7972), .Z(n8210) );
  INV_X1 U9630 ( .A(n8207), .ZN(n7977) );
  XOR2_X1 U9631 ( .A(n7974), .B(n7973), .Z(n7976) );
  AOI222_X1 U9632 ( .A1(n8167), .A2(n7976), .B1(n8000), .B2(n8092), .C1(n7975), 
        .C2(n8161), .ZN(n8205) );
  OAI21_X1 U9633 ( .B1(n7977), .B2(n8096), .A(n8205), .ZN(n7978) );
  NAND2_X1 U9634 ( .A1(n7978), .A2(n8098), .ZN(n7981) );
  AOI22_X1 U9635 ( .A1(n7979), .A2(n8102), .B1(n9907), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n7980) );
  OAI211_X1 U9636 ( .C1(n8210), .C2(n8105), .A(n7981), .B(n7980), .ZN(P2_U3209) );
  XOR2_X1 U9637 ( .A(n7983), .B(n7982), .Z(n8214) );
  XNOR2_X1 U9638 ( .A(n7984), .B(n7983), .ZN(n7985) );
  OAI222_X1 U9639 ( .A1(n8164), .A2(n7987), .B1(n8080), .B2(n7986), .C1(n8037), 
        .C2(n7985), .ZN(n8211) );
  INV_X1 U9640 ( .A(n8211), .ZN(n7988) );
  MUX2_X1 U9641 ( .A(n7989), .B(n7988), .S(n9904), .Z(n7993) );
  AOI22_X1 U9642 ( .A1(n7991), .A2(n8086), .B1(n8102), .B2(n7990), .ZN(n7992)
         );
  OAI211_X1 U9643 ( .C1(n8214), .C2(n8105), .A(n7993), .B(n7992), .ZN(P2_U3210) );
  XNOR2_X1 U9644 ( .A(n7995), .B(n7994), .ZN(n8222) );
  INV_X1 U9645 ( .A(n7996), .ZN(n8002) );
  OAI21_X1 U9646 ( .B1(n7999), .B2(n7998), .A(n7997), .ZN(n8001) );
  AOI222_X1 U9647 ( .A1(n8167), .A2(n8001), .B1(n8000), .B2(n8161), .C1(n8026), 
        .C2(n8092), .ZN(n8217) );
  OAI21_X1 U9648 ( .B1(n8002), .B2(n9896), .A(n8217), .ZN(n8003) );
  NAND2_X1 U9649 ( .A1(n8003), .A2(n8098), .ZN(n8005) );
  AOI22_X1 U9650 ( .A1(n8219), .A2(n8086), .B1(P2_REG2_REG_22__SCAN_IN), .B2(
        n9907), .ZN(n8004) );
  OAI211_X1 U9651 ( .C1(n8222), .C2(n8105), .A(n8005), .B(n8004), .ZN(P2_U3211) );
  NAND2_X1 U9652 ( .A1(n8007), .A2(n8006), .ZN(n8008) );
  XNOR2_X1 U9653 ( .A(n8008), .B(n8009), .ZN(n8228) );
  INV_X1 U9654 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8017) );
  INV_X1 U9655 ( .A(n8009), .ZN(n8011) );
  NAND3_X1 U9656 ( .A1(n8023), .A2(n8011), .A3(n8010), .ZN(n8012) );
  NAND2_X1 U9657 ( .A1(n8013), .A2(n8012), .ZN(n8016) );
  AOI222_X1 U9658 ( .A1(n8167), .A2(n8016), .B1(n8015), .B2(n8092), .C1(n8014), 
        .C2(n8161), .ZN(n8223) );
  MUX2_X1 U9659 ( .A(n8017), .B(n8223), .S(n9904), .Z(n8020) );
  AOI22_X1 U9660 ( .A1(n8225), .A2(n8086), .B1(n8102), .B2(n8018), .ZN(n8019)
         );
  OAI211_X1 U9661 ( .C1(n8228), .C2(n8105), .A(n8020), .B(n8019), .ZN(P2_U3212) );
  XNOR2_X1 U9662 ( .A(n8021), .B(n8024), .ZN(n8234) );
  INV_X1 U9663 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8028) );
  AND2_X1 U9664 ( .A1(n8034), .A2(n8022), .ZN(n8025) );
  OAI21_X1 U9665 ( .B1(n8025), .B2(n8024), .A(n8023), .ZN(n8027) );
  AOI222_X1 U9666 ( .A1(n8167), .A2(n8027), .B1(n8051), .B2(n8092), .C1(n8026), 
        .C2(n8161), .ZN(n8229) );
  MUX2_X1 U9667 ( .A(n8028), .B(n8229), .S(n9904), .Z(n8031) );
  AOI22_X1 U9668 ( .A1(n8231), .A2(n8086), .B1(n8102), .B2(n8029), .ZN(n8030)
         );
  OAI211_X1 U9669 ( .C1(n8234), .C2(n8105), .A(n8031), .B(n8030), .ZN(P2_U3213) );
  XNOR2_X1 U9670 ( .A(n8033), .B(n8032), .ZN(n8240) );
  INV_X1 U9671 ( .A(n8034), .ZN(n8039) );
  AOI21_X1 U9672 ( .B1(n8049), .B2(n8036), .A(n8035), .ZN(n8038) );
  NOR3_X1 U9673 ( .A1(n8039), .A2(n8038), .A3(n8037), .ZN(n8043) );
  OAI22_X1 U9674 ( .A1(n8041), .A2(n8080), .B1(n8040), .B2(n8164), .ZN(n8042)
         );
  NOR2_X1 U9675 ( .A1(n8043), .A2(n8042), .ZN(n8235) );
  MUX2_X1 U9676 ( .A(n8044), .B(n8235), .S(n9904), .Z(n8047) );
  AOI22_X1 U9677 ( .A1(n8237), .A2(n8086), .B1(n8102), .B2(n8045), .ZN(n8046)
         );
  OAI211_X1 U9678 ( .C1(n8240), .C2(n8105), .A(n8047), .B(n8046), .ZN(P2_U3214) );
  XNOR2_X1 U9679 ( .A(n8048), .B(n8050), .ZN(n8246) );
  OAI21_X1 U9680 ( .B1(n4344), .B2(n8050), .A(n8049), .ZN(n8052) );
  AOI222_X1 U9681 ( .A1(n8167), .A2(n8052), .B1(n8071), .B2(n8092), .C1(n8051), 
        .C2(n8161), .ZN(n8241) );
  MUX2_X1 U9682 ( .A(n8053), .B(n8241), .S(n9904), .Z(n8056) );
  AOI22_X1 U9683 ( .A1(n8243), .A2(n8086), .B1(n8102), .B2(n8054), .ZN(n8055)
         );
  OAI211_X1 U9684 ( .C1(n8246), .C2(n8105), .A(n8056), .B(n8055), .ZN(P2_U3215) );
  XNOR2_X1 U9685 ( .A(n8057), .B(n5185), .ZN(n8060) );
  AOI222_X1 U9686 ( .A1(n8167), .A2(n8060), .B1(n8059), .B2(n8161), .C1(n8058), 
        .C2(n8092), .ZN(n8146) );
  OAI22_X1 U9687 ( .A1(n8098), .A2(n9887), .B1(n8061), .B2(n9896), .ZN(n8062)
         );
  AOI21_X1 U9688 ( .B1(n8143), .B2(n8086), .A(n8062), .ZN(n8067) );
  OAI21_X1 U9689 ( .B1(n8064), .B2(n5185), .A(n8063), .ZN(n8144) );
  NAND2_X1 U9690 ( .A1(n8144), .A2(n8065), .ZN(n8066) );
  OAI211_X1 U9691 ( .C1(n8146), .C2(n9907), .A(n8067), .B(n8066), .ZN(P2_U3216) );
  XNOR2_X1 U9692 ( .A(n8068), .B(n8069), .ZN(n8253) );
  XNOR2_X1 U9693 ( .A(n8070), .B(n8069), .ZN(n8072) );
  AOI222_X1 U9694 ( .A1(n8167), .A2(n8072), .B1(n8071), .B2(n8161), .C1(n8094), 
        .C2(n8092), .ZN(n8248) );
  MUX2_X1 U9695 ( .A(n8073), .B(n8248), .S(n9904), .Z(n8076) );
  AOI22_X1 U9696 ( .A1(n8250), .A2(n8086), .B1(n8102), .B2(n8074), .ZN(n8075)
         );
  OAI211_X1 U9697 ( .C1(n8253), .C2(n8105), .A(n8076), .B(n8075), .ZN(P2_U3217) );
  XNOR2_X1 U9698 ( .A(n8077), .B(n8078), .ZN(n8259) );
  XNOR2_X1 U9699 ( .A(n8079), .B(n8078), .ZN(n8084) );
  OAI22_X1 U9700 ( .A1(n8082), .A2(n8164), .B1(n8081), .B2(n8080), .ZN(n8083)
         );
  AOI21_X1 U9701 ( .B1(n8084), .B2(n8167), .A(n8083), .ZN(n8255) );
  MUX2_X1 U9702 ( .A(n8255), .B(n9850), .S(n9907), .Z(n8088) );
  AOI22_X1 U9703 ( .A1(n8256), .A2(n8086), .B1(n8102), .B2(n8085), .ZN(n8087)
         );
  OAI211_X1 U9704 ( .C1(n8259), .C2(n8105), .A(n8088), .B(n8087), .ZN(P2_U3218) );
  XOR2_X1 U9705 ( .A(n8089), .B(n8091), .Z(n8267) );
  INV_X1 U9706 ( .A(n8263), .ZN(n8097) );
  XOR2_X1 U9707 ( .A(n8090), .B(n8091), .Z(n8095) );
  AOI222_X1 U9708 ( .A1(n8167), .A2(n8095), .B1(n8094), .B2(n8161), .C1(n8093), 
        .C2(n8092), .ZN(n8260) );
  OAI21_X1 U9709 ( .B1(n8097), .B2(n8096), .A(n8260), .ZN(n8099) );
  NAND2_X1 U9710 ( .A1(n8099), .A2(n8098), .ZN(n8104) );
  INV_X1 U9711 ( .A(n8100), .ZN(n8101) );
  AOI22_X1 U9712 ( .A1(n9907), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8102), .B2(
        n8101), .ZN(n8103) );
  OAI211_X1 U9713 ( .C1(n8267), .C2(n8105), .A(n8104), .B(n8103), .ZN(P2_U3219) );
  NAND2_X1 U9714 ( .A1(n6211), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8106) );
  NAND2_X1 U9715 ( .A1(n8181), .A2(n9982), .ZN(n8107) );
  OAI211_X1 U9716 ( .C1(n8180), .C2(n8126), .A(n8106), .B(n8107), .ZN(P2_U3490) );
  INV_X1 U9717 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8109) );
  NAND2_X1 U9718 ( .A1(n8183), .A2(n8152), .ZN(n8108) );
  OAI211_X1 U9719 ( .C1(n9982), .C2(n8109), .A(n8108), .B(n8107), .ZN(P2_U3489) );
  INV_X1 U9720 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8113) );
  NAND2_X1 U9721 ( .A1(n8110), .A2(n9962), .ZN(n8111) );
  OAI21_X1 U9722 ( .B1(n8190), .B2(n8126), .A(n8114), .ZN(P2_U3487) );
  MUX2_X1 U9723 ( .A(n8191), .B(P2_REG1_REG_27__SCAN_IN), .S(n6211), .Z(n8117)
         );
  INV_X1 U9724 ( .A(n8115), .ZN(n8193) );
  OAI22_X1 U9725 ( .A1(n8193), .A2(n8155), .B1(n8192), .B2(n8126), .ZN(n8116)
         );
  OR2_X1 U9726 ( .A1(n8117), .A2(n8116), .ZN(P2_U3486) );
  INV_X1 U9727 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8120) );
  AOI21_X1 U9728 ( .B1(n8119), .B2(n9962), .A(n8118), .ZN(n8196) );
  MUX2_X1 U9729 ( .A(n9039), .B(n8199), .S(n9982), .Z(n8122) );
  NAND2_X1 U9730 ( .A1(n8201), .A2(n8152), .ZN(n8121) );
  OAI211_X1 U9731 ( .C1(n8204), .C2(n8155), .A(n8122), .B(n8121), .ZN(P2_U3484) );
  INV_X1 U9732 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8123) );
  MUX2_X1 U9733 ( .A(n8123), .B(n8205), .S(n9982), .Z(n8125) );
  NAND2_X1 U9734 ( .A1(n8207), .A2(n8152), .ZN(n8124) );
  OAI211_X1 U9735 ( .C1(n8155), .C2(n8210), .A(n8125), .B(n8124), .ZN(P2_U3483) );
  MUX2_X1 U9736 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8211), .S(n9982), .Z(n8128)
         );
  OAI22_X1 U9737 ( .A1(n8214), .A2(n8155), .B1(n8213), .B2(n8126), .ZN(n8127)
         );
  OR2_X1 U9738 ( .A1(n8128), .A2(n8127), .ZN(P2_U3482) );
  INV_X1 U9739 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9054) );
  MUX2_X1 U9740 ( .A(n9054), .B(n8217), .S(n9982), .Z(n8130) );
  NAND2_X1 U9741 ( .A1(n8219), .A2(n8152), .ZN(n8129) );
  OAI211_X1 U9742 ( .C1(n8155), .C2(n8222), .A(n8130), .B(n8129), .ZN(P2_U3481) );
  INV_X1 U9743 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8131) );
  MUX2_X1 U9744 ( .A(n8131), .B(n8223), .S(n9982), .Z(n8133) );
  NAND2_X1 U9745 ( .A1(n8225), .A2(n8152), .ZN(n8132) );
  OAI211_X1 U9746 ( .C1(n8155), .C2(n8228), .A(n8133), .B(n8132), .ZN(P2_U3480) );
  INV_X1 U9747 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8134) );
  MUX2_X1 U9748 ( .A(n8134), .B(n8229), .S(n9982), .Z(n8136) );
  NAND2_X1 U9749 ( .A1(n8231), .A2(n8152), .ZN(n8135) );
  OAI211_X1 U9750 ( .C1(n8234), .C2(n8155), .A(n8136), .B(n8135), .ZN(P2_U3479) );
  MUX2_X1 U9751 ( .A(n8137), .B(n8235), .S(n9982), .Z(n8139) );
  NAND2_X1 U9752 ( .A1(n8237), .A2(n8152), .ZN(n8138) );
  OAI211_X1 U9753 ( .C1(n8240), .C2(n8155), .A(n8139), .B(n8138), .ZN(P2_U3478) );
  MUX2_X1 U9754 ( .A(n8140), .B(n8241), .S(n9982), .Z(n8142) );
  NAND2_X1 U9755 ( .A1(n8243), .A2(n8152), .ZN(n8141) );
  OAI211_X1 U9756 ( .C1(n8155), .C2(n8246), .A(n8142), .B(n8141), .ZN(P2_U3477) );
  AOI22_X1 U9757 ( .A1(n8144), .A2(n9962), .B1(n9966), .B2(n8143), .ZN(n8145)
         );
  NAND2_X1 U9758 ( .A1(n8146), .A2(n8145), .ZN(n8247) );
  MUX2_X1 U9759 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8247), .S(n9982), .Z(
        P2_U3476) );
  MUX2_X1 U9760 ( .A(n9050), .B(n8248), .S(n9982), .Z(n8148) );
  NAND2_X1 U9761 ( .A1(n8250), .A2(n8152), .ZN(n8147) );
  OAI211_X1 U9762 ( .C1(n8253), .C2(n8155), .A(n8148), .B(n8147), .ZN(P2_U3475) );
  MUX2_X1 U9763 ( .A(n9040), .B(n8255), .S(n9982), .Z(n8150) );
  NAND2_X1 U9764 ( .A1(n8256), .A2(n8152), .ZN(n8149) );
  OAI211_X1 U9765 ( .C1(n8155), .C2(n8259), .A(n8150), .B(n8149), .ZN(P2_U3474) );
  MUX2_X1 U9766 ( .A(n8151), .B(n8260), .S(n9982), .Z(n8154) );
  NAND2_X1 U9767 ( .A1(n8263), .A2(n8152), .ZN(n8153) );
  OAI211_X1 U9768 ( .C1(n8267), .C2(n8155), .A(n8154), .B(n8153), .ZN(P2_U3473) );
  XNOR2_X1 U9769 ( .A(n8157), .B(n8156), .ZN(n9902) );
  NAND2_X1 U9770 ( .A1(n9902), .A2(n8158), .ZN(n8170) );
  XNOR2_X1 U9771 ( .A(n8160), .B(n8159), .ZN(n8168) );
  NAND2_X1 U9772 ( .A1(n8162), .A2(n8161), .ZN(n8163) );
  OAI21_X1 U9773 ( .B1(n8165), .B2(n8164), .A(n8163), .ZN(n8166) );
  AOI21_X1 U9774 ( .B1(n8168), .B2(n8167), .A(n8166), .ZN(n8169) );
  AND2_X1 U9775 ( .A1(n8170), .A2(n8169), .ZN(n9899) );
  NOR2_X1 U9776 ( .A1(n8171), .A2(n9948), .ZN(n9895) );
  AOI21_X1 U9777 ( .B1(n9902), .B2(n9953), .A(n9895), .ZN(n8172) );
  AND2_X1 U9778 ( .A1(n9899), .A2(n8172), .ZN(n9909) );
  INV_X1 U9779 ( .A(n9909), .ZN(n8173) );
  MUX2_X1 U9780 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n8173), .S(n9982), .Z(
        P2_U3461) );
  AOI22_X1 U9781 ( .A1(n8175), .A2(n9953), .B1(n9966), .B2(n8174), .ZN(n8176)
         );
  AND2_X1 U9782 ( .A1(n8177), .A2(n8176), .ZN(n9908) );
  INV_X1 U9783 ( .A(n9908), .ZN(n8178) );
  MUX2_X1 U9784 ( .A(n8178), .B(P2_REG1_REG_1__SCAN_IN), .S(n6211), .Z(
        P2_U3460) );
  MUX2_X1 U9785 ( .A(n8179), .B(P2_REG1_REG_0__SCAN_IN), .S(n6211), .Z(
        P2_U3459) );
  NAND2_X1 U9786 ( .A1(n4623), .A2(n8262), .ZN(n8182) );
  NAND2_X1 U9787 ( .A1(n8181), .A2(n9967), .ZN(n8184) );
  OAI211_X1 U9788 ( .C1(n7618), .C2(n9967), .A(n8182), .B(n8184), .ZN(P2_U3458) );
  NAND2_X1 U9789 ( .A1(n8183), .A2(n8262), .ZN(n8185) );
  OAI211_X1 U9790 ( .C1(n9967), .C2(n8186), .A(n8185), .B(n8184), .ZN(P2_U3457) );
  OAI21_X1 U9791 ( .B1(n8190), .B2(n8212), .A(n8189), .ZN(P2_U3455) );
  MUX2_X1 U9792 ( .A(n8191), .B(P2_REG0_REG_27__SCAN_IN), .S(n9969), .Z(n8195)
         );
  OAI22_X1 U9793 ( .A1(n8193), .A2(n8266), .B1(n8192), .B2(n8212), .ZN(n8194)
         );
  OR2_X1 U9794 ( .A1(n8195), .A2(n8194), .ZN(P2_U3454) );
  INV_X1 U9795 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8200) );
  MUX2_X1 U9796 ( .A(n8200), .B(n8199), .S(n9967), .Z(n8203) );
  NAND2_X1 U9797 ( .A1(n8201), .A2(n8262), .ZN(n8202) );
  OAI211_X1 U9798 ( .C1(n8204), .C2(n8266), .A(n8203), .B(n8202), .ZN(P2_U3452) );
  MUX2_X1 U9799 ( .A(n8206), .B(n8205), .S(n9967), .Z(n8209) );
  NAND2_X1 U9800 ( .A1(n8207), .A2(n8262), .ZN(n8208) );
  OAI211_X1 U9801 ( .C1(n8210), .C2(n8266), .A(n8209), .B(n8208), .ZN(P2_U3451) );
  MUX2_X1 U9802 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8211), .S(n9967), .Z(n8216)
         );
  OAI22_X1 U9803 ( .A1(n8214), .A2(n8266), .B1(n8213), .B2(n8212), .ZN(n8215)
         );
  OR2_X1 U9804 ( .A1(n8216), .A2(n8215), .ZN(P2_U3450) );
  INV_X1 U9805 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8218) );
  MUX2_X1 U9806 ( .A(n8218), .B(n8217), .S(n9967), .Z(n8221) );
  NAND2_X1 U9807 ( .A1(n8219), .A2(n8262), .ZN(n8220) );
  OAI211_X1 U9808 ( .C1(n8222), .C2(n8266), .A(n8221), .B(n8220), .ZN(P2_U3449) );
  INV_X1 U9809 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8224) );
  MUX2_X1 U9810 ( .A(n8224), .B(n8223), .S(n9967), .Z(n8227) );
  NAND2_X1 U9811 ( .A1(n8225), .A2(n8262), .ZN(n8226) );
  OAI211_X1 U9812 ( .C1(n8228), .C2(n8266), .A(n8227), .B(n8226), .ZN(P2_U3448) );
  INV_X1 U9813 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8230) );
  MUX2_X1 U9814 ( .A(n8230), .B(n8229), .S(n9967), .Z(n8233) );
  NAND2_X1 U9815 ( .A1(n8231), .A2(n8262), .ZN(n8232) );
  OAI211_X1 U9816 ( .C1(n8234), .C2(n8266), .A(n8233), .B(n8232), .ZN(P2_U3447) );
  MUX2_X1 U9817 ( .A(n8236), .B(n8235), .S(n9967), .Z(n8239) );
  NAND2_X1 U9818 ( .A1(n8237), .A2(n8262), .ZN(n8238) );
  OAI211_X1 U9819 ( .C1(n8240), .C2(n8266), .A(n8239), .B(n8238), .ZN(P2_U3446) );
  INV_X1 U9820 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8242) );
  MUX2_X1 U9821 ( .A(n8242), .B(n8241), .S(n9967), .Z(n8245) );
  NAND2_X1 U9822 ( .A1(n8243), .A2(n8262), .ZN(n8244) );
  OAI211_X1 U9823 ( .C1(n8246), .C2(n8266), .A(n8245), .B(n8244), .ZN(P2_U3444) );
  MUX2_X1 U9824 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8247), .S(n9967), .Z(
        P2_U3441) );
  INV_X1 U9825 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8249) );
  MUX2_X1 U9826 ( .A(n8249), .B(n8248), .S(n9967), .Z(n8252) );
  NAND2_X1 U9827 ( .A1(n8250), .A2(n8262), .ZN(n8251) );
  OAI211_X1 U9828 ( .C1(n8253), .C2(n8266), .A(n8252), .B(n8251), .ZN(P2_U3438) );
  INV_X1 U9829 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8254) );
  MUX2_X1 U9830 ( .A(n8255), .B(n8254), .S(n9969), .Z(n8258) );
  NAND2_X1 U9831 ( .A1(n8256), .A2(n8262), .ZN(n8257) );
  OAI211_X1 U9832 ( .C1(n8259), .C2(n8266), .A(n8258), .B(n8257), .ZN(P2_U3435) );
  INV_X1 U9833 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8261) );
  MUX2_X1 U9834 ( .A(n8261), .B(n8260), .S(n9967), .Z(n8265) );
  NAND2_X1 U9835 ( .A1(n8263), .A2(n8262), .ZN(n8264) );
  OAI211_X1 U9836 ( .C1(n8267), .C2(n8266), .A(n8265), .B(n8264), .ZN(P2_U3432) );
  INV_X1 U9837 ( .A(n8268), .ZN(n9493) );
  INV_X1 U9838 ( .A(n8269), .ZN(n8271) );
  NOR4_X1 U9839 ( .A1(n8271), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n5169), .ZN(n8272) );
  AOI21_X1 U9840 ( .B1(n8273), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8272), .ZN(
        n8274) );
  OAI21_X1 U9841 ( .B1(n9493), .B2(n8277), .A(n8274), .ZN(P2_U3264) );
  INV_X1 U9842 ( .A(n8275), .ZN(n9501) );
  OAI222_X1 U9843 ( .A1(P2_U3151), .A2(n8278), .B1(n8277), .B2(n9501), .C1(
        n9077), .C2(n8276), .ZN(P2_U3266) );
  MUX2_X1 U9844 ( .A(n8279), .B(P2_IR_REG_0__SCAN_IN), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  AOI21_X1 U9845 ( .B1(n8282), .B2(n8281), .A(n8280), .ZN(n8283) );
  OAI21_X1 U9846 ( .B1(n8284), .B2(n8283), .A(n9573), .ZN(n8290) );
  AND2_X1 U9847 ( .A1(n8722), .A2(n9224), .ZN(n8285) );
  AOI21_X1 U9848 ( .B1(n8908), .B2(n9222), .A(n8285), .ZN(n8952) );
  INV_X1 U9849 ( .A(n8286), .ZN(n8956) );
  AOI22_X1 U9850 ( .A1(n8956), .A2(n8433), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n8287) );
  OAI21_X1 U9851 ( .B1(n8952), .B2(n8419), .A(n8287), .ZN(n8288) );
  AOI21_X1 U9852 ( .B1(n9427), .B2(n8422), .A(n8288), .ZN(n8289) );
  NAND2_X1 U9853 ( .A1(n8290), .A2(n8289), .ZN(P1_U3214) );
  OAI21_X1 U9854 ( .B1(n8293), .B2(n8292), .A(n8291), .ZN(n8294) );
  NAND2_X1 U9855 ( .A1(n8294), .A2(n9573), .ZN(n8297) );
  AOI22_X1 U9856 ( .A1(n9224), .A2(n8725), .B1(n8876), .B2(n9222), .ZN(n9304)
         );
  NAND2_X1 U9857 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9628) );
  OAI21_X1 U9858 ( .B1(n8419), .B2(n9304), .A(n9628), .ZN(n8295) );
  AOI21_X1 U9859 ( .B1(n9313), .B2(n8433), .A(n8295), .ZN(n8296) );
  OAI211_X1 U9860 ( .C1(n9484), .C2(n9570), .A(n8297), .B(n8296), .ZN(P1_U3215) );
  INV_X1 U9861 ( .A(n8298), .ZN(n8395) );
  INV_X1 U9862 ( .A(n8299), .ZN(n8301) );
  NOR3_X1 U9863 ( .A1(n8395), .A2(n8301), .A3(n8300), .ZN(n8304) );
  INV_X1 U9864 ( .A(n8302), .ZN(n8303) );
  OAI21_X1 U9865 ( .B1(n8304), .B2(n8303), .A(n9573), .ZN(n8310) );
  NAND2_X1 U9866 ( .A1(n8898), .A2(n9222), .ZN(n8306) );
  NAND2_X1 U9867 ( .A1(n8892), .A2(n9224), .ZN(n8305) );
  NAND2_X1 U9868 ( .A1(n8306), .A2(n8305), .ZN(n9010) );
  OAI22_X1 U9869 ( .A1(n9015), .A2(n9577), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8307), .ZN(n8308) );
  AOI21_X1 U9870 ( .B1(n9010), .B2(n9568), .A(n8308), .ZN(n8309) );
  OAI211_X1 U9871 ( .C1(n9014), .C2(n9570), .A(n8310), .B(n8309), .ZN(P1_U3216) );
  OAI21_X1 U9872 ( .B1(n8313), .B2(n8312), .A(n8311), .ZN(n8314) );
  NAND2_X1 U9873 ( .A1(n8314), .A2(n9573), .ZN(n8319) );
  AOI22_X1 U9874 ( .A1(n9568), .A2(n8316), .B1(n8422), .B2(n8315), .ZN(n8318)
         );
  MUX2_X1 U9875 ( .A(n9577), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n8317) );
  NAND3_X1 U9876 ( .A1(n8319), .A2(n8318), .A3(n8317), .ZN(P1_U3218) );
  XNOR2_X1 U9877 ( .A(n8322), .B(n8321), .ZN(n8323) );
  XNOR2_X1 U9878 ( .A(n8320), .B(n8323), .ZN(n8328) );
  OAI22_X1 U9879 ( .A1(n9577), .A2(n9216), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8324), .ZN(n8326) );
  INV_X1 U9880 ( .A(n9225), .ZN(n8880) );
  INV_X1 U9881 ( .A(n9223), .ZN(n8885) );
  OAI22_X1 U9882 ( .A1(n8430), .A2(n8880), .B1(n8885), .B2(n8429), .ZN(n8325)
         );
  AOI211_X1 U9883 ( .C1(n9372), .C2(n8422), .A(n8326), .B(n8325), .ZN(n8327)
         );
  OAI21_X1 U9884 ( .B1(n8328), .B2(n8424), .A(n8327), .ZN(P1_U3219) );
  OAI21_X1 U9885 ( .B1(n8331), .B2(n8330), .A(n8329), .ZN(n8332) );
  NAND2_X1 U9886 ( .A1(n8332), .A2(n9573), .ZN(n8337) );
  AND2_X1 U9887 ( .A1(n9223), .A2(n9224), .ZN(n8333) );
  AOI21_X1 U9888 ( .B1(n8892), .B2(n9222), .A(n8333), .ZN(n9185) );
  OAI22_X1 U9889 ( .A1(n9185), .A2(n8419), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8334), .ZN(n8335) );
  AOI21_X1 U9890 ( .B1(n9190), .B2(n8433), .A(n8335), .ZN(n8336) );
  OAI211_X1 U9891 ( .C1(n9459), .C2(n9570), .A(n8337), .B(n8336), .ZN(P1_U3223) );
  OAI21_X1 U9892 ( .B1(n8339), .B2(n8338), .A(n6260), .ZN(n8340) );
  NAND2_X1 U9893 ( .A1(n8340), .A2(n9573), .ZN(n8346) );
  NAND2_X1 U9894 ( .A1(n8722), .A2(n9222), .ZN(n8342) );
  NAND2_X1 U9895 ( .A1(n8898), .A2(n9224), .ZN(n8341) );
  NAND2_X1 U9896 ( .A1(n8342), .A2(n8341), .ZN(n8980) );
  OAI22_X1 U9897 ( .A1(n8983), .A2(n9577), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8343), .ZN(n8344) );
  AOI21_X1 U9898 ( .B1(n8980), .B2(n9568), .A(n8344), .ZN(n8345) );
  OAI211_X1 U9899 ( .C1(n4511), .C2(n9570), .A(n8346), .B(n8345), .ZN(P1_U3225) );
  OAI21_X1 U9900 ( .B1(n8349), .B2(n8348), .A(n8347), .ZN(n8350) );
  NAND2_X1 U9901 ( .A1(n8350), .A2(n9573), .ZN(n8353) );
  AOI22_X1 U9902 ( .A1(n8878), .A2(n9222), .B1(n8876), .B2(n9224), .ZN(n9266)
         );
  NAND2_X1 U9903 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8817) );
  OAI21_X1 U9904 ( .B1(n8419), .B2(n9266), .A(n8817), .ZN(n8351) );
  AOI21_X1 U9905 ( .B1(n9271), .B2(n8433), .A(n8351), .ZN(n8352) );
  OAI211_X1 U9906 ( .C1(n9477), .C2(n9570), .A(n8353), .B(n8352), .ZN(P1_U3226) );
  INV_X1 U9907 ( .A(n8354), .ZN(n8359) );
  AOI21_X1 U9908 ( .B1(n8356), .B2(n8358), .A(n8355), .ZN(n8357) );
  AOI21_X1 U9909 ( .B1(n8359), .B2(n8358), .A(n8357), .ZN(n8363) );
  OAI22_X1 U9910 ( .A1(n8880), .A2(n9287), .B1(n9286), .B2(n9285), .ZN(n9254)
         );
  NAND2_X1 U9911 ( .A1(n9254), .A2(n9568), .ZN(n8360) );
  NAND2_X1 U9912 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8836) );
  OAI211_X1 U9913 ( .C1(n9577), .C2(n9258), .A(n8360), .B(n8836), .ZN(n8361)
         );
  AOI21_X1 U9914 ( .B1(n9385), .B2(n8422), .A(n8361), .ZN(n8362) );
  OAI21_X1 U9915 ( .B1(n8363), .B2(n8424), .A(n8362), .ZN(P1_U3228) );
  INV_X1 U9916 ( .A(n8365), .ZN(n8366) );
  NAND3_X1 U9917 ( .A1(n8302), .A2(n8367), .A3(n8366), .ZN(n8368) );
  AOI21_X1 U9918 ( .B1(n8364), .B2(n8368), .A(n8424), .ZN(n8372) );
  INV_X1 U9919 ( .A(n9442), .ZN(n9001) );
  AOI22_X1 U9920 ( .A1(n8998), .A2(n8433), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n8370) );
  AOI22_X1 U9921 ( .A1(n8995), .A2(n8407), .B1(n8409), .B2(n9166), .ZN(n8369)
         );
  OAI211_X1 U9922 ( .C1(n9001), .C2(n9570), .A(n8370), .B(n8369), .ZN(n8371)
         );
  OR2_X1 U9923 ( .A1(n8372), .A2(n8371), .ZN(P1_U3229) );
  INV_X1 U9924 ( .A(n8375), .ZN(n8376) );
  AOI21_X1 U9925 ( .B1(n8373), .B2(n8377), .A(n8376), .ZN(n8383) );
  NOR2_X1 U9926 ( .A1(n9577), .A2(n9206), .ZN(n8381) );
  AND2_X1 U9927 ( .A1(n8883), .A2(n9224), .ZN(n8378) );
  AOI21_X1 U9928 ( .B1(n9165), .B2(n9222), .A(n8378), .ZN(n9201) );
  OAI22_X1 U9929 ( .A1(n9201), .A2(n8419), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8379), .ZN(n8380) );
  AOI211_X1 U9930 ( .C1(n9205), .C2(n8422), .A(n8381), .B(n8380), .ZN(n8382)
         );
  OAI21_X1 U9931 ( .B1(n8383), .B2(n8424), .A(n8382), .ZN(P1_U3233) );
  OAI21_X1 U9932 ( .B1(n8386), .B2(n8385), .A(n8384), .ZN(n8387) );
  NAND2_X1 U9933 ( .A1(n8387), .A2(n9573), .ZN(n8393) );
  NAND2_X1 U9934 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9616) );
  INV_X1 U9935 ( .A(n9616), .ZN(n8390) );
  OAI22_X1 U9936 ( .A1(n8430), .A2(n8388), .B1(n9284), .B2(n8429), .ZN(n8389)
         );
  AOI211_X1 U9937 ( .C1(n8433), .C2(n8391), .A(n8390), .B(n8389), .ZN(n8392)
         );
  OAI211_X1 U9938 ( .C1(n8871), .C2(n9570), .A(n8393), .B(n8392), .ZN(P1_U3234) );
  AOI21_X1 U9939 ( .B1(n8396), .B2(n8394), .A(n8395), .ZN(n8401) );
  OAI22_X1 U9940 ( .A1(n9171), .A2(n9577), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8397), .ZN(n8399) );
  INV_X1 U9941 ( .A(n9166), .ZN(n8895) );
  OAI22_X1 U9942 ( .A1(n8895), .A2(n8429), .B1(n8887), .B2(n8430), .ZN(n8398)
         );
  AOI211_X1 U9943 ( .C1(n9452), .C2(n8422), .A(n8399), .B(n8398), .ZN(n8400)
         );
  OAI21_X1 U9944 ( .B1(n8401), .B2(n8424), .A(n8400), .ZN(P1_U3235) );
  OAI21_X1 U9945 ( .B1(n8404), .B2(n8403), .A(n8402), .ZN(n8405) );
  NAND2_X1 U9946 ( .A1(n8405), .A2(n9573), .ZN(n8412) );
  AOI22_X1 U9947 ( .A1(n8407), .A2(n8734), .B1(n8406), .B2(n8422), .ZN(n8411)
         );
  AOI22_X1 U9948 ( .A1(n8409), .A2(n4370), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n8408), .ZN(n8410) );
  NAND3_X1 U9949 ( .A1(n8412), .A2(n8411), .A3(n8410), .ZN(P1_U3237) );
  XNOR2_X1 U9950 ( .A(n8415), .B(n8414), .ZN(n8416) );
  XNOR2_X1 U9951 ( .A(n8413), .B(n8416), .ZN(n8425) );
  NOR2_X1 U9952 ( .A1(n9577), .A2(n9243), .ZN(n8421) );
  AND2_X1 U9953 ( .A1(n8878), .A2(n9224), .ZN(n8417) );
  AOI21_X1 U9954 ( .B1(n8883), .B2(n9222), .A(n8417), .ZN(n9241) );
  OAI22_X1 U9955 ( .A1(n9241), .A2(n8419), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8418), .ZN(n8420) );
  AOI211_X1 U9956 ( .C1(n9380), .C2(n8422), .A(n8421), .B(n8420), .ZN(n8423)
         );
  OAI21_X1 U9957 ( .B1(n8425), .B2(n8424), .A(n8423), .ZN(P1_U3238) );
  OAI21_X1 U9958 ( .B1(n4348), .B2(n8427), .A(n8426), .ZN(n8428) );
  NAND2_X1 U9959 ( .A1(n8428), .A2(n9573), .ZN(n8435) );
  NAND2_X1 U9960 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9642) );
  INV_X1 U9961 ( .A(n9642), .ZN(n8432) );
  OAI22_X1 U9962 ( .A1(n8430), .A2(n9284), .B1(n9286), .B2(n8429), .ZN(n8431)
         );
  AOI211_X1 U9963 ( .C1(n8433), .C2(n9289), .A(n8432), .B(n8431), .ZN(n8434)
         );
  OAI211_X1 U9964 ( .C1(n4524), .C2(n9570), .A(n8435), .B(n8434), .ZN(P1_U3241) );
  NAND2_X1 U9965 ( .A1(n9452), .A2(n8891), .ZN(n8437) );
  NAND2_X1 U9966 ( .A1(n9008), .A2(n8437), .ZN(n8594) );
  NAND2_X1 U9967 ( .A1(n9189), .A2(n8887), .ZN(n8519) );
  INV_X1 U9968 ( .A(n8519), .ZN(n8436) );
  NAND2_X1 U9969 ( .A1(n9161), .A2(n8436), .ZN(n8438) );
  AND2_X1 U9970 ( .A1(n8917), .A2(n8437), .ZN(n8613) );
  INV_X1 U9971 ( .A(n8567), .ZN(n8439) );
  NAND2_X1 U9972 ( .A1(n8567), .A2(n9008), .ZN(n8608) );
  OR2_X1 U9973 ( .A1(n9189), .A2(n8887), .ZN(n8686) );
  OR2_X1 U9974 ( .A1(n9205), .A2(n8885), .ZN(n8684) );
  AND2_X1 U9975 ( .A1(n8686), .A2(n8684), .ZN(n8512) );
  NAND2_X1 U9976 ( .A1(n9270), .A2(n9286), .ZN(n8673) );
  INV_X1 U9977 ( .A(n8878), .ZN(n8877) );
  OR2_X1 U9978 ( .A1(n9385), .A2(n8877), .ZN(n9237) );
  AND2_X1 U9979 ( .A1(n9237), .A2(n8675), .ZN(n8444) );
  MUX2_X1 U9980 ( .A(n8673), .B(n8444), .S(n8561), .Z(n8509) );
  NAND2_X1 U9981 ( .A1(n8732), .A2(n8561), .ZN(n8453) );
  INV_X1 U9982 ( .A(n8453), .ZN(n8447) );
  AOI22_X1 U9983 ( .A1(n8447), .A2(n8452), .B1(n8731), .B2(n8561), .ZN(n8459)
         );
  NAND2_X1 U9984 ( .A1(n8448), .A2(n4252), .ZN(n8451) );
  OAI22_X1 U9985 ( .A1(n8451), .A2(n8452), .B1(n8561), .B2(n8731), .ZN(n8449)
         );
  OAI21_X1 U9986 ( .B1(n8451), .B2(n8731), .A(n8450), .ZN(n8456) );
  OAI21_X1 U9987 ( .B1(n8454), .B2(n8453), .A(n8452), .ZN(n8455) );
  NAND2_X1 U9988 ( .A1(n8456), .A2(n8455), .ZN(n8457) );
  AND4_X1 U9989 ( .A1(n8462), .A2(n8461), .A3(n8460), .A4(n8561), .ZN(n8464)
         );
  AOI21_X1 U9990 ( .B1(n8465), .B2(n8464), .A(n8463), .ZN(n8467) );
  NAND4_X1 U9991 ( .A1(n8468), .A2(n4314), .A3(n8467), .A4(n8466), .ZN(n8473)
         );
  AND2_X1 U9992 ( .A1(n8469), .A2(n8577), .ZN(n8471) );
  NAND2_X1 U9993 ( .A1(n8473), .A2(n8472), .ZN(n8477) );
  MUX2_X1 U9994 ( .A(n8475), .B(n8474), .S(n8561), .Z(n8476) );
  NAND2_X1 U9995 ( .A1(n8477), .A2(n8476), .ZN(n8486) );
  INV_X1 U9996 ( .A(n8486), .ZN(n8479) );
  NAND2_X1 U9997 ( .A1(n8494), .A2(n8488), .ZN(n8480) );
  INV_X1 U9998 ( .A(n8487), .ZN(n8478) );
  NOR2_X1 U9999 ( .A1(n8480), .A2(n8478), .ZN(n8664) );
  OAI21_X1 U10000 ( .B1(n8485), .B2(n8479), .A(n8664), .ZN(n8483) );
  INV_X1 U10001 ( .A(n8480), .ZN(n8588) );
  NAND2_X1 U10002 ( .A1(n8492), .A2(n8490), .ZN(n8482) );
  INV_X1 U10003 ( .A(n8493), .ZN(n8481) );
  AOI21_X1 U10004 ( .B1(n8588), .B2(n8482), .A(n8481), .ZN(n8665) );
  NAND2_X1 U10005 ( .A1(n8483), .A2(n8665), .ZN(n8497) );
  OAI21_X1 U10006 ( .B1(n8486), .B2(n8485), .A(n8484), .ZN(n8491) );
  NAND2_X1 U10007 ( .A1(n8488), .A2(n8487), .ZN(n8489) );
  NAND2_X1 U10008 ( .A1(n8493), .A2(n8492), .ZN(n8569) );
  OAI21_X1 U10009 ( .B1(n8495), .B2(n8569), .A(n8494), .ZN(n8496) );
  NAND2_X1 U10010 ( .A1(n9311), .A2(n9284), .ZN(n8503) );
  NAND2_X1 U10011 ( .A1(n8667), .A2(n8503), .ZN(n8875) );
  MUX2_X1 U10012 ( .A(n8620), .B(n8498), .S(n4252), .Z(n8499) );
  OR2_X1 U10013 ( .A1(n8875), .A2(n8499), .ZN(n8500) );
  AOI21_X1 U10014 ( .B1(n8501), .B2(n8589), .A(n8500), .ZN(n8507) );
  INV_X1 U10015 ( .A(n8876), .ZN(n8502) );
  OR2_X1 U10016 ( .A1(n9396), .A2(n8502), .ZN(n8670) );
  NAND2_X1 U10017 ( .A1(n8670), .A2(n8667), .ZN(n8504) );
  NAND2_X1 U10018 ( .A1(n9396), .A2(n8502), .ZN(n8623) );
  NAND2_X1 U10019 ( .A1(n8623), .A2(n8503), .ZN(n8672) );
  MUX2_X1 U10020 ( .A(n8504), .B(n8672), .S(n4252), .Z(n8506) );
  MUX2_X1 U10021 ( .A(n8623), .B(n8670), .S(n4252), .Z(n8505) );
  NAND2_X1 U10022 ( .A1(n9380), .A2(n8880), .ZN(n8626) );
  NAND2_X1 U10023 ( .A1(n9385), .A2(n8877), .ZN(n8625) );
  NAND2_X1 U10024 ( .A1(n8626), .A2(n8625), .ZN(n8677) );
  INV_X1 U10025 ( .A(n8883), .ZN(n8882) );
  OR2_X1 U10026 ( .A1(n9372), .A2(n8882), .ZN(n8517) );
  OR2_X1 U10027 ( .A1(n9380), .A2(n8880), .ZN(n8568) );
  AND2_X1 U10028 ( .A1(n8517), .A2(n8568), .ZN(n8680) );
  NAND2_X1 U10029 ( .A1(n9372), .A2(n8882), .ZN(n8681) );
  NAND2_X1 U10030 ( .A1(n9205), .A2(n8885), .ZN(n9179) );
  NAND3_X1 U10031 ( .A1(n8510), .A2(n8681), .A3(n9179), .ZN(n8511) );
  NAND3_X1 U10032 ( .A1(n8567), .A2(n8512), .A3(n8511), .ZN(n8523) );
  INV_X1 U10033 ( .A(n8512), .ZN(n8522) );
  INV_X1 U10034 ( .A(n8625), .ZN(n8514) );
  AND2_X1 U10035 ( .A1(n8568), .A2(n9237), .ZN(n8679) );
  OAI21_X1 U10036 ( .B1(n8515), .B2(n8514), .A(n8679), .ZN(n8516) );
  NAND3_X1 U10037 ( .A1(n8516), .A2(n8681), .A3(n8626), .ZN(n8518) );
  NAND2_X1 U10038 ( .A1(n8518), .A2(n8517), .ZN(n8521) );
  NAND2_X1 U10039 ( .A1(n8519), .A2(n9179), .ZN(n8520) );
  NAND2_X1 U10040 ( .A1(n8520), .A2(n8686), .ZN(n9163) );
  INV_X1 U10041 ( .A(n8898), .ZN(n8897) );
  OR2_X1 U10042 ( .A1(n9442), .A2(n8897), .ZN(n8918) );
  NAND2_X1 U10043 ( .A1(n9442), .A2(n8897), .ZN(n8614) );
  NAND2_X1 U10044 ( .A1(n8918), .A2(n8614), .ZN(n8990) );
  NOR2_X1 U10045 ( .A1(n8917), .A2(n8561), .ZN(n8524) );
  NOR2_X1 U10046 ( .A1(n8990), .A2(n8524), .ZN(n8525) );
  MUX2_X1 U10047 ( .A(n8614), .B(n8918), .S(n4252), .Z(n8528) );
  NAND2_X1 U10048 ( .A1(n8529), .A2(n8528), .ZN(n8533) );
  INV_X1 U10049 ( .A(n8995), .ZN(n8900) );
  NAND2_X1 U10050 ( .A1(n9436), .A2(n8900), .ZN(n8920) );
  NAND2_X1 U10051 ( .A1(n8533), .A2(n8920), .ZN(n8530) );
  OR2_X1 U10052 ( .A1(n9436), .A2(n8900), .ZN(n8612) );
  NAND2_X1 U10053 ( .A1(n8530), .A2(n8612), .ZN(n8531) );
  INV_X1 U10054 ( .A(n8722), .ZN(n8902) );
  NOR2_X1 U10055 ( .A1(n9340), .A2(n8902), .ZN(n8535) );
  NAND2_X1 U10056 ( .A1(n8533), .A2(n8612), .ZN(n8534) );
  NAND3_X1 U10057 ( .A1(n8534), .A2(n8922), .A3(n8920), .ZN(n8536) );
  INV_X1 U10058 ( .A(n8535), .ZN(n8607) );
  NAND2_X1 U10059 ( .A1(n8536), .A2(n8607), .ZN(n8537) );
  INV_X1 U10060 ( .A(n8721), .ZN(n8905) );
  NAND2_X1 U10061 ( .A1(n9427), .A2(n8905), .ZN(n8598) );
  INV_X1 U10062 ( .A(n8908), .ZN(n8929) );
  OR2_X1 U10063 ( .A1(n8929), .A2(n9331), .ZN(n8605) );
  MUX2_X1 U10064 ( .A(n4252), .B(n9427), .S(n8721), .Z(n8540) );
  NAND2_X1 U10065 ( .A1(n8541), .A2(n8540), .ZN(n8543) );
  NAND2_X1 U10066 ( .A1(n9331), .A2(n8929), .ZN(n8924) );
  NAND2_X1 U10067 ( .A1(n8924), .A2(n8598), .ZN(n8618) );
  NAND2_X1 U10068 ( .A1(n8618), .A2(n4252), .ZN(n8542) );
  NAND2_X1 U10069 ( .A1(n8543), .A2(n8542), .ZN(n8544) );
  NAND2_X1 U10070 ( .A1(n8544), .A2(n8605), .ZN(n8545) );
  NAND2_X1 U10071 ( .A1(n8546), .A2(n8545), .ZN(n8549) );
  INV_X1 U10072 ( .A(n8720), .ZN(n8547) );
  OR2_X1 U10073 ( .A1(n9417), .A2(n8547), .ZN(n8606) );
  NAND2_X1 U10074 ( .A1(n9417), .A2(n8547), .ZN(n8633) );
  OR2_X1 U10075 ( .A1(n8924), .A2(n4252), .ZN(n8548) );
  MUX2_X1 U10076 ( .A(n8633), .B(n8606), .S(n8561), .Z(n8550) );
  MUX2_X1 U10077 ( .A(n8560), .B(n4252), .S(n8696), .Z(n8559) );
  OR2_X1 U10078 ( .A1(n8563), .A2(n8637), .ZN(n8699) );
  NAND2_X1 U10079 ( .A1(n4265), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8557) );
  NAND2_X1 U10080 ( .A1(n8553), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8556) );
  NAND2_X1 U10081 ( .A1(n8554), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8555) );
  NAND3_X1 U10082 ( .A1(n8557), .A2(n8556), .A3(n8555), .ZN(n8719) );
  NAND2_X1 U10083 ( .A1(n8558), .A2(n8719), .ZN(n8635) );
  NAND3_X1 U10084 ( .A1(n8559), .A2(n8699), .A3(n8635), .ZN(n8565) );
  MUX2_X1 U10085 ( .A(n8561), .B(n8560), .S(n8696), .Z(n8562) );
  NAND3_X1 U10086 ( .A1(n8562), .A2(n8563), .A3(n8719), .ZN(n8564) );
  NAND2_X1 U10087 ( .A1(n8563), .A2(n8637), .ZN(n8701) );
  NAND3_X1 U10088 ( .A1(n8565), .A2(n8564), .A3(n8701), .ZN(n8649) );
  NAND2_X1 U10089 ( .A1(n8649), .A2(n8716), .ZN(n8604) );
  NAND2_X1 U10090 ( .A1(n8612), .A2(n8920), .ZN(n8919) );
  INV_X1 U10091 ( .A(n8990), .ZN(n8993) );
  NAND2_X1 U10092 ( .A1(n8684), .A2(n9179), .ZN(n9197) );
  XNOR2_X1 U10093 ( .A(n9372), .B(n8882), .ZN(n9213) );
  NAND2_X1 U10094 ( .A1(n8670), .A2(n8623), .ZN(n9281) );
  INV_X1 U10095 ( .A(n8569), .ZN(n8587) );
  NAND4_X1 U10096 ( .A1(n8573), .A2(n8572), .A3(n8651), .A4(n8571), .ZN(n8576)
         );
  NOR3_X1 U10097 ( .A1(n8576), .A2(n8575), .A3(n8574), .ZN(n8580) );
  NAND4_X1 U10098 ( .A1(n8580), .A2(n8579), .A3(n8578), .A4(n8577), .ZN(n8581)
         );
  OR3_X1 U10099 ( .A1(n8583), .A2(n8582), .A3(n8581), .ZN(n8585) );
  NOR2_X1 U10100 ( .A1(n8585), .A2(n8584), .ZN(n8586) );
  NAND4_X1 U10101 ( .A1(n8589), .A2(n8588), .A3(n8587), .A4(n8586), .ZN(n8590)
         );
  OR3_X1 U10102 ( .A1(n9281), .A2(n8590), .A3(n8875), .ZN(n8591) );
  NOR2_X1 U10103 ( .A1(n4689), .A2(n8591), .ZN(n8592) );
  XNOR2_X1 U10104 ( .A(n9385), .B(n8878), .ZN(n9252) );
  NAND3_X1 U10105 ( .A1(n9239), .A2(n8592), .A3(n9252), .ZN(n8593) );
  NOR3_X1 U10106 ( .A1(n9197), .A2(n9213), .A3(n8593), .ZN(n8596) );
  XNOR2_X1 U10107 ( .A(n9189), .B(n8887), .ZN(n9181) );
  NOR2_X1 U10108 ( .A1(n8594), .A2(n9181), .ZN(n8595) );
  NAND4_X1 U10109 ( .A1(n8993), .A2(n9007), .A3(n8596), .A4(n8595), .ZN(n8597)
         );
  OR2_X1 U10110 ( .A1(n8919), .A2(n8597), .ZN(n8599) );
  NAND2_X1 U10111 ( .A1(n8605), .A2(n8924), .ZN(n8933) );
  NAND2_X1 U10112 ( .A1(n8923), .A2(n8598), .ZN(n8948) );
  NAND2_X1 U10113 ( .A1(n8607), .A2(n8922), .ZN(n8964) );
  OR4_X1 U10114 ( .A1(n8599), .A2(n8933), .A3(n8948), .A4(n8964), .ZN(n8600)
         );
  NOR2_X1 U10115 ( .A1(n8926), .A2(n8600), .ZN(n8602) );
  XNOR2_X1 U10116 ( .A(n8696), .B(n8719), .ZN(n8601) );
  NAND4_X1 U10117 ( .A1(n8699), .A2(n8701), .A3(n8602), .A4(n8601), .ZN(n8642)
         );
  INV_X1 U10118 ( .A(n8642), .ZN(n8603) );
  NAND2_X1 U10119 ( .A1(n8606), .A2(n8605), .ZN(n8695) );
  NAND2_X1 U10120 ( .A1(n8923), .A2(n8607), .ZN(n8691) );
  NAND2_X1 U10121 ( .A1(n8608), .A2(n8917), .ZN(n8609) );
  NAND2_X1 U10122 ( .A1(n8918), .A2(n8609), .ZN(n8610) );
  NAND2_X1 U10123 ( .A1(n8610), .A2(n8614), .ZN(n8611) );
  AND2_X1 U10124 ( .A1(n8612), .A2(n8611), .ZN(n8619) );
  NAND3_X1 U10125 ( .A1(n8614), .A2(n8613), .A3(n9163), .ZN(n8615) );
  AOI21_X1 U10126 ( .B1(n8619), .B2(n8615), .A(n4431), .ZN(n8616) );
  NOR2_X1 U10127 ( .A1(n8691), .A2(n8616), .ZN(n8617) );
  OR2_X1 U10128 ( .A1(n8618), .A2(n8617), .ZN(n8693) );
  INV_X1 U10129 ( .A(n8619), .ZN(n8688) );
  NOR2_X1 U10130 ( .A1(n8875), .A2(n8620), .ZN(n8621) );
  NAND2_X1 U10131 ( .A1(n9298), .A2(n8621), .ZN(n8622) );
  NAND2_X1 U10132 ( .A1(n8622), .A2(n8667), .ZN(n9280) );
  INV_X1 U10133 ( .A(n8673), .ZN(n8624) );
  NAND2_X1 U10134 ( .A1(n9253), .A2(n8625), .ZN(n9238) );
  NAND2_X1 U10135 ( .A1(n9238), .A2(n8679), .ZN(n8627) );
  NAND2_X1 U10136 ( .A1(n8627), .A2(n8626), .ZN(n9221) );
  INV_X1 U10137 ( .A(n9213), .ZN(n9220) );
  NAND2_X1 U10138 ( .A1(n9221), .A2(n9220), .ZN(n8628) );
  OAI21_X1 U10139 ( .B1(n8688), .B2(n9162), .A(n8922), .ZN(n8629) );
  INV_X1 U10140 ( .A(n8629), .ZN(n8630) );
  NOR2_X1 U10141 ( .A1(n8691), .A2(n8630), .ZN(n8631) );
  NOR2_X1 U10142 ( .A1(n8693), .A2(n8631), .ZN(n8632) );
  NOR2_X1 U10143 ( .A1(n8695), .A2(n8632), .ZN(n8636) );
  INV_X1 U10144 ( .A(n8719), .ZN(n8927) );
  NAND2_X1 U10145 ( .A1(n8696), .A2(n8927), .ZN(n8634) );
  NAND2_X1 U10146 ( .A1(n8634), .A2(n8633), .ZN(n8697) );
  OAI22_X1 U10147 ( .A1(n8636), .A2(n8697), .B1(n8696), .B2(n8635), .ZN(n8639)
         );
  NAND2_X1 U10148 ( .A1(n8696), .A2(n8637), .ZN(n8638) );
  NAND3_X1 U10149 ( .A1(n8639), .A2(n8699), .A3(n8638), .ZN(n8641) );
  NAND3_X1 U10150 ( .A1(n8641), .A2(n8640), .A3(n8701), .ZN(n8643) );
  NAND2_X1 U10151 ( .A1(n8643), .A2(n8642), .ZN(n8644) );
  OR2_X1 U10152 ( .A1(n8701), .A2(n8646), .ZN(n8648) );
  OAI211_X1 U10153 ( .C1(n8699), .C2(n8646), .A(n8645), .B(n6171), .ZN(n8647)
         );
  AOI21_X1 U10154 ( .B1(n8649), .B2(n8648), .A(n8647), .ZN(n8650) );
  AOI21_X1 U10155 ( .B1(n4370), .B2(n9669), .A(n8651), .ZN(n8655) );
  NAND4_X1 U10156 ( .A1(n8655), .A2(n8654), .A3(n8653), .A4(n8652), .ZN(n8657)
         );
  NOR2_X1 U10157 ( .A1(n8657), .A2(n8656), .ZN(n8659) );
  NAND3_X1 U10158 ( .A1(n8660), .A2(n8659), .A3(n8658), .ZN(n8661) );
  NAND2_X1 U10159 ( .A1(n8662), .A2(n8661), .ZN(n8663) );
  NAND2_X1 U10160 ( .A1(n8664), .A2(n8663), .ZN(n8666) );
  NAND3_X1 U10161 ( .A1(n8666), .A2(n8665), .A3(n9297), .ZN(n8669) );
  AND3_X1 U10162 ( .A1(n8669), .A2(n8668), .A3(n8667), .ZN(n8671) );
  OAI21_X1 U10163 ( .B1(n8672), .B2(n8671), .A(n8670), .ZN(n8674) );
  NAND2_X1 U10164 ( .A1(n8674), .A2(n8673), .ZN(n8676) );
  AND2_X1 U10165 ( .A1(n8676), .A2(n8675), .ZN(n8678) );
  AOI21_X1 U10166 ( .B1(n8679), .B2(n8678), .A(n8677), .ZN(n8683) );
  INV_X1 U10167 ( .A(n8680), .ZN(n8682) );
  OAI21_X1 U10168 ( .B1(n8683), .B2(n8682), .A(n8681), .ZN(n8685) );
  NAND3_X1 U10169 ( .A1(n8686), .A2(n8685), .A3(n8684), .ZN(n8687) );
  OAI21_X1 U10170 ( .B1(n8688), .B2(n8687), .A(n8922), .ZN(n8689) );
  INV_X1 U10171 ( .A(n8689), .ZN(n8690) );
  NOR2_X1 U10172 ( .A1(n8691), .A2(n8690), .ZN(n8692) );
  NOR2_X1 U10173 ( .A1(n8693), .A2(n8692), .ZN(n8694) );
  NOR2_X1 U10174 ( .A1(n8695), .A2(n8694), .ZN(n8698) );
  OAI22_X1 U10175 ( .A1(n8698), .A2(n8697), .B1(n8927), .B2(n8696), .ZN(n8700)
         );
  NAND2_X1 U10176 ( .A1(n8700), .A2(n8699), .ZN(n8702) );
  NAND2_X1 U10177 ( .A1(n8702), .A2(n8701), .ZN(n8708) );
  NAND2_X1 U10178 ( .A1(n8708), .A2(n9016), .ZN(n8703) );
  INV_X1 U10179 ( .A(n8710), .ZN(n8718) );
  INV_X1 U10180 ( .A(n8711), .ZN(n8713) );
  NAND4_X1 U10181 ( .A1(n8712), .A2(n8713), .A3(n9486), .A4(n8752), .ZN(n8714)
         );
  OAI211_X1 U10182 ( .C1(n8716), .C2(n8715), .A(n8714), .B(P1_B_REG_SCAN_IN), 
        .ZN(n8717) );
  NAND2_X1 U10183 ( .A1(n8718), .A2(n8717), .ZN(P1_U3242) );
  MUX2_X1 U10184 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n8719), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10185 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n8720), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10186 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n8908), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10187 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n8721), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10188 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n8722), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10189 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n8995), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10190 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n8898), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10191 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9166), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10192 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n8892), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10193 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9165), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10194 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9223), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10195 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n8883), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10196 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9225), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10197 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n8878), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10198 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n8723), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10199 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n8724), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10200 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n8725), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10201 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n8726), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10202 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n8727), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10203 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n8728), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10204 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n8729), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10205 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n8730), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10206 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n8731), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10207 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n8732), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10208 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n8733), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10209 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n8734), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10210 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n8735), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10211 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n4370), .S(P1_U3973), .Z(
        P1_U3555) );
  INV_X1 U10212 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n8737) );
  OAI22_X1 U10213 ( .A1(n9661), .A2(n8737), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8736), .ZN(n8738) );
  AOI21_X1 U10214 ( .B1(n8739), .B2(n4463), .A(n8738), .ZN(n8747) );
  OAI211_X1 U10215 ( .C1(n8751), .C2(n8741), .A(n9595), .B(n8740), .ZN(n8746)
         );
  AND2_X1 U10216 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n8743) );
  OAI211_X1 U10217 ( .C1(n8744), .C2(n8743), .A(n9648), .B(n8742), .ZN(n8745)
         );
  NAND3_X1 U10218 ( .A1(n8747), .A2(n8746), .A3(n8745), .ZN(P1_U3244) );
  NAND3_X1 U10219 ( .A1(n8750), .A2(n8749), .A3(n8748), .ZN(n8756) );
  AOI22_X1 U10220 ( .A1(n8754), .A2(n8753), .B1(n8752), .B2(n8751), .ZN(n8755)
         );
  NAND3_X1 U10221 ( .A1(n8756), .A2(P1_U3973), .A3(n8755), .ZN(n8795) );
  INV_X1 U10222 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n8758) );
  OAI22_X1 U10223 ( .A1(n9661), .A2(n8758), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8757), .ZN(n8759) );
  AOI21_X1 U10224 ( .B1(n8760), .B2(n4463), .A(n8759), .ZN(n8769) );
  OAI211_X1 U10225 ( .C1(n8763), .C2(n8762), .A(n9648), .B(n8761), .ZN(n8768)
         );
  OAI211_X1 U10226 ( .C1(n8766), .C2(n8765), .A(n9595), .B(n8764), .ZN(n8767)
         );
  NAND4_X1 U10227 ( .A1(n8795), .A2(n8769), .A3(n8768), .A4(n8767), .ZN(
        P1_U3245) );
  AOI211_X1 U10228 ( .C1(n8772), .C2(n8771), .A(n8770), .B(n9632), .ZN(n8773)
         );
  INV_X1 U10229 ( .A(n8773), .ZN(n8783) );
  INV_X1 U10230 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n8775) );
  NAND2_X1 U10231 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n8774) );
  OAI21_X1 U10232 ( .B1(n9661), .B2(n8775), .A(n8774), .ZN(n8776) );
  AOI21_X1 U10233 ( .B1(n8777), .B2(n4463), .A(n8776), .ZN(n8782) );
  OAI211_X1 U10234 ( .C1(n8780), .C2(n8779), .A(n9595), .B(n8778), .ZN(n8781)
         );
  NAND3_X1 U10235 ( .A1(n8783), .A2(n8782), .A3(n8781), .ZN(P1_U3246) );
  INV_X1 U10236 ( .A(n8784), .ZN(n8788) );
  AOI211_X1 U10237 ( .C1(n4302), .C2(n8786), .A(n8785), .B(n9632), .ZN(n8787)
         );
  AOI211_X1 U10238 ( .C1(n8835), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n8788), .B(
        n8787), .ZN(n8796) );
  NAND2_X1 U10239 ( .A1(n4463), .A2(n8789), .ZN(n8794) );
  OAI211_X1 U10240 ( .C1(n8792), .C2(n8791), .A(n9595), .B(n8790), .ZN(n8793)
         );
  NAND4_X1 U10241 ( .A1(n8796), .A2(n8795), .A3(n8794), .A4(n8793), .ZN(
        P1_U3247) );
  AOI211_X1 U10242 ( .C1(n8799), .C2(n8798), .A(n9632), .B(n8797), .ZN(n8800)
         );
  INV_X1 U10243 ( .A(n8800), .ZN(n8810) );
  INV_X1 U10244 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n8802) );
  OAI21_X1 U10245 ( .B1(n9661), .B2(n8802), .A(n8801), .ZN(n8803) );
  AOI21_X1 U10246 ( .B1(n8804), .B2(n4463), .A(n8803), .ZN(n8809) );
  OAI211_X1 U10247 ( .C1(n8807), .C2(n8806), .A(n9595), .B(n8805), .ZN(n8808)
         );
  NAND3_X1 U10248 ( .A1(n8810), .A2(n8809), .A3(n8808), .ZN(P1_U3248) );
  INV_X1 U10249 ( .A(n8821), .ZN(n9615) );
  OAI21_X1 U10250 ( .B1(n8819), .B2(P1_REG1_REG_12__SCAN_IN), .A(n8811), .ZN(
        n9608) );
  XNOR2_X1 U10251 ( .A(n9615), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n9609) );
  XNOR2_X1 U10252 ( .A(n9627), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n9623) );
  NOR2_X1 U10253 ( .A1(n8812), .A2(n9631), .ZN(n8813) );
  INV_X1 U10254 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9634) );
  XNOR2_X1 U10255 ( .A(n9631), .B(n8812), .ZN(n9635) );
  NOR2_X1 U10256 ( .A1(n9634), .A2(n9635), .ZN(n9633) );
  NOR2_X1 U10257 ( .A1(n8813), .A2(n9633), .ZN(n8815) );
  INV_X1 U10258 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9392) );
  AOI22_X1 U10259 ( .A1(n8834), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n9392), .B2(
        n8825), .ZN(n8814) );
  NAND2_X1 U10260 ( .A1(n8814), .A2(n8815), .ZN(n8833) );
  OAI21_X1 U10261 ( .B1(n8815), .B2(n8814), .A(n8833), .ZN(n8830) );
  NAND2_X1 U10262 ( .A1(n8835), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n8816) );
  OAI211_X1 U10263 ( .C1(n9654), .C2(n8825), .A(n8817), .B(n8816), .ZN(n8829)
         );
  OAI21_X1 U10264 ( .B1(n8819), .B2(P1_REG2_REG_12__SCAN_IN), .A(n8818), .ZN(
        n9612) );
  INV_X1 U10265 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n8820) );
  XNOR2_X1 U10266 ( .A(n8821), .B(n8820), .ZN(n9611) );
  NOR2_X1 U10267 ( .A1(n9612), .A2(n9611), .ZN(n9610) );
  AOI21_X1 U10268 ( .B1(n9615), .B2(P1_REG2_REG_13__SCAN_IN), .A(n9610), .ZN(
        n9621) );
  NAND2_X1 U10269 ( .A1(n9627), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n8822) );
  OAI21_X1 U10270 ( .B1(n9627), .B2(P1_REG2_REG_14__SCAN_IN), .A(n8822), .ZN(
        n9620) );
  NOR2_X1 U10271 ( .A1(n9621), .A2(n9620), .ZN(n9619) );
  AOI21_X1 U10272 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n9627), .A(n9619), .ZN(
        n8823) );
  NOR2_X1 U10273 ( .A1(n8823), .A2(n9631), .ZN(n8824) );
  INV_X1 U10274 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9637) );
  XNOR2_X1 U10275 ( .A(n9631), .B(n8823), .ZN(n9638) );
  NOR2_X1 U10276 ( .A1(n9637), .A2(n9638), .ZN(n9636) );
  NOR2_X1 U10277 ( .A1(n8824), .A2(n9636), .ZN(n8827) );
  INV_X1 U10278 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9034) );
  AOI22_X1 U10279 ( .A1(n8834), .A2(n9034), .B1(P1_REG2_REG_16__SCAN_IN), .B2(
        n8825), .ZN(n8826) );
  NOR2_X1 U10280 ( .A1(n8827), .A2(n8826), .ZN(n8832) );
  AOI211_X1 U10281 ( .C1(n8827), .C2(n8826), .A(n8832), .B(n9645), .ZN(n8828)
         );
  AOI211_X1 U10282 ( .C1(n9648), .C2(n8830), .A(n8829), .B(n8828), .ZN(n8831)
         );
  INV_X1 U10283 ( .A(n8831), .ZN(P1_U3259) );
  XNOR2_X1 U10284 ( .A(n8850), .B(P1_REG2_REG_17__SCAN_IN), .ZN(n8842) );
  AOI21_X1 U10285 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n8834), .A(n8832), .ZN(
        n8843) );
  XOR2_X1 U10286 ( .A(n8842), .B(n8843), .Z(n8841) );
  OAI21_X1 U10287 ( .B1(n8834), .B2(P1_REG1_REG_16__SCAN_IN), .A(n8833), .ZN(
        n8852) );
  XNOR2_X1 U10288 ( .A(n8850), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n8851) );
  XNOR2_X1 U10289 ( .A(n8852), .B(n8851), .ZN(n8839) );
  NAND2_X1 U10290 ( .A1(n8835), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n8837) );
  OAI211_X1 U10291 ( .C1(n9654), .C2(n8850), .A(n8837), .B(n8836), .ZN(n8838)
         );
  AOI21_X1 U10292 ( .B1(n8839), .B2(n9648), .A(n8838), .ZN(n8840) );
  OAI21_X1 U10293 ( .B1(n8841), .B2(n9645), .A(n8840), .ZN(P1_U3260) );
  NAND2_X1 U10294 ( .A1(n8843), .A2(n8842), .ZN(n8845) );
  INV_X1 U10295 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9249) );
  NAND2_X1 U10296 ( .A1(n8850), .A2(n9249), .ZN(n8844) );
  NAND2_X1 U10297 ( .A1(n8845), .A2(n8844), .ZN(n9647) );
  INV_X1 U10298 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9235) );
  OR2_X1 U10299 ( .A1(n9653), .A2(n9235), .ZN(n8847) );
  NAND2_X1 U10300 ( .A1(n9653), .A2(n9235), .ZN(n8846) );
  NAND2_X1 U10301 ( .A1(n8847), .A2(n8846), .ZN(n9646) );
  NAND2_X1 U10302 ( .A1(n9656), .A2(n8847), .ZN(n8849) );
  INV_X1 U10303 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n8848) );
  XNOR2_X1 U10304 ( .A(n8849), .B(n8848), .ZN(n8857) );
  INV_X1 U10305 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9386) );
  AOI22_X1 U10306 ( .A1(n8852), .A2(n8851), .B1(n9386), .B2(n8850), .ZN(n9651)
         );
  INV_X1 U10307 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9381) );
  NOR2_X1 U10308 ( .A1(n9653), .A2(n9381), .ZN(n8853) );
  AOI21_X1 U10309 ( .B1(n9381), .B2(n9653), .A(n8853), .ZN(n9650) );
  NAND2_X1 U10310 ( .A1(n9651), .A2(n9650), .ZN(n9649) );
  INV_X1 U10311 ( .A(n8853), .ZN(n8854) );
  NAND2_X1 U10312 ( .A1(n9649), .A2(n8854), .ZN(n8856) );
  XNOR2_X1 U10313 ( .A(n8856), .B(n8855), .ZN(n8858) );
  AOI22_X1 U10314 ( .A1(n8857), .A2(n9595), .B1(n9648), .B2(n8858), .ZN(n8860)
         );
  INV_X1 U10315 ( .A(n8857), .ZN(n8859) );
  NAND2_X1 U10316 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n8861) );
  NAND2_X1 U10317 ( .A1(n8862), .A2(n9317), .ZN(n8865) );
  INV_X1 U10318 ( .A(n8863), .ZN(n9321) );
  NOR2_X1 U10319 ( .A1(n4251), .A2(n9321), .ZN(n8869) );
  AOI21_X1 U10320 ( .B1(n4251), .B2(P1_REG2_REG_31__SCAN_IN), .A(n8869), .ZN(
        n8864) );
  OAI211_X1 U10321 ( .C1(n8866), .C2(n9315), .A(n8865), .B(n8864), .ZN(
        P1_U3263) );
  OAI211_X1 U10322 ( .C1(n9416), .C2(n8910), .A(n9373), .B(n8867), .ZN(n9322)
         );
  NOR2_X1 U10323 ( .A1(n9416), .A2(n9315), .ZN(n8868) );
  AOI211_X1 U10324 ( .C1(n4251), .C2(P1_REG2_REG_30__SCAN_IN), .A(n8869), .B(
        n8868), .ZN(n8870) );
  OAI21_X1 U10325 ( .B1(n9322), .B2(n8982), .A(n8870), .ZN(P1_U3264) );
  INV_X1 U10326 ( .A(n9385), .ZN(n9250) );
  NOR2_X1 U10327 ( .A1(n9250), .A2(n8877), .ZN(n8879) );
  OAI22_X1 U10328 ( .A1(n9247), .A2(n8879), .B1(n8878), .B2(n9385), .ZN(n9231)
         );
  INV_X1 U10329 ( .A(n9239), .ZN(n8881) );
  AOI22_X1 U10330 ( .A1(n9231), .A2(n8881), .B1(n8880), .B2(n6228), .ZN(n9214)
         );
  INV_X1 U10331 ( .A(n9372), .ZN(n9219) );
  NAND2_X1 U10332 ( .A1(n9219), .A2(n8882), .ZN(n8884) );
  AOI22_X1 U10333 ( .A1(n9214), .A2(n8884), .B1(n8883), .B2(n9372), .ZN(n9196)
         );
  NAND2_X1 U10334 ( .A1(n9205), .A2(n9223), .ZN(n8886) );
  NAND2_X1 U10335 ( .A1(n9459), .A2(n8887), .ZN(n8888) );
  NAND2_X1 U10336 ( .A1(n9178), .A2(n8888), .ZN(n8890) );
  NOR2_X1 U10337 ( .A1(n9447), .A2(n9166), .ZN(n8896) );
  NOR2_X1 U10338 ( .A1(n9001), .A2(n8897), .ZN(n8899) );
  NOR2_X1 U10339 ( .A1(n8973), .A2(n8902), .ZN(n8901) );
  OR2_X1 U10340 ( .A1(n8963), .A2(n8901), .ZN(n8904) );
  NAND2_X1 U10341 ( .A1(n8973), .A2(n8902), .ZN(n8903) );
  NAND2_X1 U10342 ( .A1(n8904), .A2(n8903), .ZN(n8947) );
  NAND2_X1 U10343 ( .A1(n8947), .A2(n8948), .ZN(n8907) );
  INV_X1 U10344 ( .A(n9427), .ZN(n8958) );
  NAND2_X1 U10345 ( .A1(n8958), .A2(n8905), .ZN(n8906) );
  NOR2_X1 U10346 ( .A1(n9331), .A2(n8908), .ZN(n8909) );
  INV_X1 U10347 ( .A(n9331), .ZN(n8944) );
  AOI211_X1 U10348 ( .C1(n9417), .C2(n8939), .A(n9308), .B(n8910), .ZN(n9325)
         );
  INV_X1 U10349 ( .A(n9417), .ZN(n8915) );
  INV_X1 U10350 ( .A(n8911), .ZN(n8912) );
  NAND3_X1 U10351 ( .A1(n8912), .A2(P1_REG3_REG_28__SCAN_IN), .A3(n9312), .ZN(
        n8914) );
  NAND2_X1 U10352 ( .A1(n4251), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8913) );
  OAI211_X1 U10353 ( .C1(n8915), .C2(n9315), .A(n8914), .B(n8913), .ZN(n8916)
         );
  AOI21_X1 U10354 ( .B1(n9325), .B2(n9317), .A(n8916), .ZN(n8931) );
  INV_X1 U10355 ( .A(n8964), .ZN(n8921) );
  OR2_X1 U10356 ( .A1(n8949), .A2(n8948), .ZN(n8951) );
  NAND2_X1 U10357 ( .A1(n8951), .A2(n8923), .ZN(n8934) );
  OAI21_X1 U10358 ( .B1(n8934), .B2(n8933), .A(n8924), .ZN(n8925) );
  NAND2_X1 U10359 ( .A1(n9326), .A2(n9306), .ZN(n8930) );
  XNOR2_X1 U10360 ( .A(n8934), .B(n8933), .ZN(n8935) );
  NAND2_X1 U10361 ( .A1(n8935), .A2(n9301), .ZN(n8937) );
  NAND2_X1 U10362 ( .A1(n8937), .A2(n8936), .ZN(n9329) );
  INV_X1 U10363 ( .A(n8939), .ZN(n8940) );
  AOI211_X1 U10364 ( .C1(n9331), .C2(n8955), .A(n9308), .B(n8940), .ZN(n9330)
         );
  NAND2_X1 U10365 ( .A1(n9330), .A2(n9317), .ZN(n8943) );
  AOI22_X1 U10366 ( .A1(n8941), .A2(n9312), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n4251), .ZN(n8942) );
  OAI211_X1 U10367 ( .C1(n8944), .C2(n9315), .A(n8943), .B(n8942), .ZN(n8945)
         );
  AOI21_X1 U10368 ( .B1(n9306), .B2(n9329), .A(n8945), .ZN(n8946) );
  OAI21_X1 U10369 ( .B1(n9424), .B2(n9294), .A(n8946), .ZN(P1_U3265) );
  XOR2_X1 U10370 ( .A(n8947), .B(n8948), .Z(n9429) );
  NAND2_X1 U10371 ( .A1(n8949), .A2(n8948), .ZN(n8950) );
  NAND3_X1 U10372 ( .A1(n8951), .A2(n9301), .A3(n8950), .ZN(n8953) );
  AND2_X1 U10373 ( .A1(n8953), .A2(n8952), .ZN(n9335) );
  INV_X1 U10374 ( .A(n9335), .ZN(n8961) );
  INV_X1 U10375 ( .A(n8954), .ZN(n8969) );
  OAI211_X1 U10376 ( .C1(n8969), .C2(n8958), .A(n9373), .B(n8955), .ZN(n9334)
         );
  NOR2_X1 U10377 ( .A1(n9334), .A2(n8982), .ZN(n8960) );
  AOI22_X1 U10378 ( .A1(n8956), .A2(n9312), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n4251), .ZN(n8957) );
  OAI21_X1 U10379 ( .B1(n8958), .B2(n9315), .A(n8957), .ZN(n8959) );
  AOI211_X1 U10380 ( .C1(n8961), .C2(n9306), .A(n8960), .B(n8959), .ZN(n8962)
         );
  OAI21_X1 U10381 ( .B1(n9429), .B2(n9294), .A(n8962), .ZN(P1_U3266) );
  XNOR2_X1 U10382 ( .A(n8963), .B(n8964), .ZN(n9433) );
  XNOR2_X1 U10383 ( .A(n8965), .B(n8964), .ZN(n8968) );
  INV_X1 U10384 ( .A(n8966), .ZN(n8967) );
  OAI21_X1 U10385 ( .B1(n8968), .B2(n9283), .A(n8967), .ZN(n9338) );
  AOI211_X1 U10386 ( .C1(n9340), .C2(n4272), .A(n9308), .B(n8969), .ZN(n9339)
         );
  NAND2_X1 U10387 ( .A1(n9339), .A2(n9317), .ZN(n8972) );
  AOI22_X1 U10388 ( .A1(n8970), .A2(n9312), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n4251), .ZN(n8971) );
  OAI211_X1 U10389 ( .C1(n8973), .C2(n9315), .A(n8972), .B(n8971), .ZN(n8974)
         );
  AOI21_X1 U10390 ( .B1(n9306), .B2(n9338), .A(n8974), .ZN(n8975) );
  OAI21_X1 U10391 ( .B1(n9433), .B2(n9294), .A(n8975), .ZN(P1_U3267) );
  XNOR2_X1 U10392 ( .A(n8976), .B(n8979), .ZN(n9438) );
  OAI21_X1 U10393 ( .B1(n8979), .B2(n8978), .A(n8977), .ZN(n8981) );
  AOI21_X1 U10394 ( .B1(n8981), .B2(n9301), .A(n8980), .ZN(n9344) );
  INV_X1 U10395 ( .A(n9344), .ZN(n8988) );
  OAI211_X1 U10396 ( .C1(n4511), .C2(n4292), .A(n4272), .B(n9373), .ZN(n9343)
         );
  NOR2_X1 U10397 ( .A1(n9343), .A2(n8982), .ZN(n8987) );
  INV_X1 U10398 ( .A(n8983), .ZN(n8984) );
  AOI22_X1 U10399 ( .A1(n8984), .A2(n9312), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n4251), .ZN(n8985) );
  OAI21_X1 U10400 ( .B1(n4511), .B2(n9315), .A(n8985), .ZN(n8986) );
  AOI211_X1 U10401 ( .C1(n8988), .C2(n9306), .A(n8987), .B(n8986), .ZN(n8989)
         );
  OAI21_X1 U10402 ( .B1(n9438), .B2(n9294), .A(n8989), .ZN(P1_U3268) );
  XNOR2_X1 U10403 ( .A(n8991), .B(n8990), .ZN(n9444) );
  OAI211_X1 U10404 ( .C1(n8994), .C2(n8993), .A(n8992), .B(n9301), .ZN(n8997)
         );
  AOI22_X1 U10405 ( .A1(n8995), .A2(n9222), .B1(n9224), .B2(n9166), .ZN(n8996)
         );
  NAND2_X1 U10406 ( .A1(n8997), .A2(n8996), .ZN(n9347) );
  AOI211_X1 U10407 ( .C1(n9442), .C2(n9013), .A(n9308), .B(n4292), .ZN(n9348)
         );
  NAND2_X1 U10408 ( .A1(n9348), .A2(n9317), .ZN(n9000) );
  AOI22_X1 U10409 ( .A1(n8998), .A2(n9312), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n4251), .ZN(n8999) );
  OAI211_X1 U10410 ( .C1(n9001), .C2(n9315), .A(n9000), .B(n8999), .ZN(n9002)
         );
  AOI21_X1 U10411 ( .B1(n9306), .B2(n9347), .A(n9002), .ZN(n9003) );
  OAI21_X1 U10412 ( .B1(n9444), .B2(n9294), .A(n9003), .ZN(P1_U3269) );
  XNOR2_X1 U10413 ( .A(n9004), .B(n9007), .ZN(n9449) );
  AOI22_X1 U10414 ( .A1(n9447), .A2(n9005), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n4251), .ZN(n9019) );
  AOI21_X1 U10415 ( .B1(n9008), .B2(n9164), .A(n9007), .ZN(n9009) );
  OAI21_X1 U10416 ( .B1(n4539), .B2(n9009), .A(n9301), .ZN(n9012) );
  INV_X1 U10417 ( .A(n9010), .ZN(n9011) );
  NAND2_X1 U10418 ( .A1(n9012), .A2(n9011), .ZN(n9352) );
  OAI211_X1 U10419 ( .C1(n9014), .C2(n9170), .A(n9373), .B(n9013), .ZN(n9353)
         );
  OAI22_X1 U10420 ( .A1(n9353), .A2(n9016), .B1(n9257), .B2(n9015), .ZN(n9017)
         );
  OAI21_X1 U10421 ( .B1(n9352), .B2(n9017), .A(n9306), .ZN(n9018) );
  OAI211_X1 U10422 ( .C1(n9449), .C2(n9294), .A(n9019), .B(n9018), .ZN(n9158)
         );
  AOI22_X1 U10423 ( .A1(n9022), .A2(keyinput6), .B1(keyinput57), .B2(n9021), 
        .ZN(n9020) );
  OAI221_X1 U10424 ( .B1(n9022), .B2(keyinput6), .C1(n9021), .C2(keyinput57), 
        .A(n9020), .ZN(n9032) );
  INV_X1 U10425 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n9024) );
  AOI22_X1 U10426 ( .A1(n9025), .A2(keyinput34), .B1(keyinput45), .B2(n9024), 
        .ZN(n9023) );
  OAI221_X1 U10427 ( .B1(n9025), .B2(keyinput34), .C1(n9024), .C2(keyinput45), 
        .A(n9023), .ZN(n9031) );
  INV_X1 U10428 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9481) );
  AOI22_X1 U10429 ( .A1(n9142), .A2(keyinput62), .B1(keyinput19), .B2(n9481), 
        .ZN(n9026) );
  OAI221_X1 U10430 ( .B1(n9142), .B2(keyinput62), .C1(n9481), .C2(keyinput19), 
        .A(n9026), .ZN(n9030) );
  INV_X1 U10431 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9028) );
  AOI22_X1 U10432 ( .A1(n9028), .A2(keyinput37), .B1(n6546), .B2(keyinput63), 
        .ZN(n9027) );
  OAI221_X1 U10433 ( .B1(n9028), .B2(keyinput37), .C1(n6546), .C2(keyinput63), 
        .A(n9027), .ZN(n9029) );
  NOR4_X1 U10434 ( .A1(n9032), .A2(n9031), .A3(n9030), .A4(n9029), .ZN(n9104)
         );
  AOI22_X1 U10435 ( .A1(n9034), .A2(keyinput31), .B1(n9461), .B2(keyinput20), 
        .ZN(n9033) );
  OAI221_X1 U10436 ( .B1(n9034), .B2(keyinput31), .C1(n9461), .C2(keyinput20), 
        .A(n9033), .ZN(n9044) );
  INV_X1 U10437 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n9665) );
  AOI22_X1 U10438 ( .A1(n7989), .A2(keyinput0), .B1(n9665), .B2(keyinput46), 
        .ZN(n9035) );
  OAI221_X1 U10439 ( .B1(n7989), .B2(keyinput0), .C1(n9665), .C2(keyinput46), 
        .A(n9035), .ZN(n9043) );
  INV_X1 U10440 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9037) );
  AOI22_X1 U10441 ( .A1(n5850), .A2(keyinput61), .B1(keyinput38), .B2(n9037), 
        .ZN(n9036) );
  OAI221_X1 U10442 ( .B1(n5850), .B2(keyinput61), .C1(n9037), .C2(keyinput38), 
        .A(n9036), .ZN(n9042) );
  AOI22_X1 U10443 ( .A1(n9040), .A2(keyinput2), .B1(n9039), .B2(keyinput48), 
        .ZN(n9038) );
  OAI221_X1 U10444 ( .B1(n9040), .B2(keyinput2), .C1(n9039), .C2(keyinput48), 
        .A(n9038), .ZN(n9041) );
  NOR4_X1 U10445 ( .A1(n9044), .A2(n9043), .A3(n9042), .A4(n9041), .ZN(n9103)
         );
  AOI22_X1 U10446 ( .A1(n7614), .A2(keyinput59), .B1(n9046), .B2(keyinput49), 
        .ZN(n9045) );
  OAI221_X1 U10447 ( .B1(n7614), .B2(keyinput59), .C1(n9046), .C2(keyinput49), 
        .A(n9045), .ZN(n9058) );
  INV_X1 U10448 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9960) );
  AOI22_X1 U10449 ( .A1(n9048), .A2(keyinput56), .B1(keyinput1), .B2(n9960), 
        .ZN(n9047) );
  OAI221_X1 U10450 ( .B1(n9048), .B2(keyinput56), .C1(n9960), .C2(keyinput1), 
        .A(n9047), .ZN(n9057) );
  AOI22_X1 U10451 ( .A1(n9051), .A2(keyinput40), .B1(keyinput53), .B2(n9050), 
        .ZN(n9049) );
  OAI221_X1 U10452 ( .B1(n9051), .B2(keyinput40), .C1(n9050), .C2(keyinput53), 
        .A(n9049), .ZN(n9056) );
  AOI22_X1 U10453 ( .A1(n9054), .A2(keyinput10), .B1(n9053), .B2(keyinput18), 
        .ZN(n9052) );
  OAI221_X1 U10454 ( .B1(n9054), .B2(keyinput10), .C1(n9053), .C2(keyinput18), 
        .A(n9052), .ZN(n9055) );
  NOR4_X1 U10455 ( .A1(n9058), .A2(n9057), .A3(n9056), .A4(n9055), .ZN(n9102)
         );
  INV_X1 U10456 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n9663) );
  AOI22_X1 U10457 ( .A1(n9148), .A2(keyinput33), .B1(n9663), .B2(keyinput47), 
        .ZN(n9059) );
  OAI221_X1 U10458 ( .B1(n9148), .B2(keyinput33), .C1(n9663), .C2(keyinput47), 
        .A(n9059), .ZN(n9063) );
  INV_X1 U10459 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n9137) );
  AOI22_X1 U10460 ( .A1(n9137), .A2(keyinput50), .B1(n9061), .B2(keyinput36), 
        .ZN(n9060) );
  OAI221_X1 U10461 ( .B1(n9137), .B2(keyinput50), .C1(n9061), .C2(keyinput36), 
        .A(n9060), .ZN(n9062) );
  NOR2_X1 U10462 ( .A1(n9063), .A2(n9062), .ZN(n9072) );
  AOI22_X1 U10463 ( .A1(n7259), .A2(keyinput54), .B1(n9850), .B2(keyinput22), 
        .ZN(n9064) );
  OAI221_X1 U10464 ( .B1(n7259), .B2(keyinput54), .C1(n9850), .C2(keyinput22), 
        .A(n9064), .ZN(n9070) );
  XNOR2_X1 U10465 ( .A(SI_17_), .B(keyinput51), .ZN(n9068) );
  XNOR2_X1 U10466 ( .A(P2_IR_REG_11__SCAN_IN), .B(keyinput32), .ZN(n9067) );
  XNOR2_X1 U10467 ( .A(P1_REG0_REG_16__SCAN_IN), .B(keyinput3), .ZN(n9066) );
  XNOR2_X1 U10468 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput16), .ZN(n9065) );
  NAND4_X1 U10469 ( .A1(n9068), .A2(n9067), .A3(n9066), .A4(n9065), .ZN(n9069)
         );
  NOR2_X1 U10470 ( .A1(n9070), .A2(n9069), .ZN(n9071) );
  AND2_X1 U10471 ( .A1(n9072), .A2(n9071), .ZN(n9100) );
  AOI22_X1 U10472 ( .A1(n5077), .A2(keyinput43), .B1(n9074), .B2(keyinput30), 
        .ZN(n9073) );
  OAI221_X1 U10473 ( .B1(n5077), .B2(keyinput43), .C1(n9074), .C2(keyinput30), 
        .A(n9073), .ZN(n9082) );
  AOI22_X1 U10474 ( .A1(n9077), .A2(keyinput42), .B1(n9076), .B2(keyinput52), 
        .ZN(n9075) );
  OAI221_X1 U10475 ( .B1(n9077), .B2(keyinput42), .C1(n9076), .C2(keyinput52), 
        .A(n9075), .ZN(n9081) );
  XNOR2_X1 U10476 ( .A(P1_REG2_REG_2__SCAN_IN), .B(keyinput21), .ZN(n9079) );
  XNOR2_X1 U10477 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput12), .ZN(n9078) );
  NAND2_X1 U10478 ( .A1(n9079), .A2(n9078), .ZN(n9080) );
  NOR3_X1 U10479 ( .A1(n9082), .A2(n9081), .A3(n9080), .ZN(n9099) );
  INV_X1 U10480 ( .A(SI_15_), .ZN(n9084) );
  AOI22_X1 U10481 ( .A1(n9084), .A2(keyinput4), .B1(n9138), .B2(keyinput25), 
        .ZN(n9083) );
  OAI221_X1 U10482 ( .B1(n9084), .B2(keyinput4), .C1(n9138), .C2(keyinput25), 
        .A(n9083), .ZN(n9087) );
  XNOR2_X1 U10483 ( .A(n9085), .B(keyinput39), .ZN(n9086) );
  NOR2_X1 U10484 ( .A1(n9087), .A2(n9086), .ZN(n9098) );
  INV_X1 U10485 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9590) );
  AOI22_X1 U10486 ( .A1(n9590), .A2(keyinput60), .B1(n9089), .B2(keyinput55), 
        .ZN(n9088) );
  OAI221_X1 U10487 ( .B1(n9590), .B2(keyinput60), .C1(n9089), .C2(keyinput55), 
        .A(n9088), .ZN(n9096) );
  AOI22_X1 U10488 ( .A1(n9092), .A2(keyinput24), .B1(keyinput17), .B2(n9091), 
        .ZN(n9090) );
  OAI221_X1 U10489 ( .B1(n9092), .B2(keyinput24), .C1(n9091), .C2(keyinput17), 
        .A(n9090), .ZN(n9095) );
  XNOR2_X1 U10490 ( .A(n9093), .B(keyinput58), .ZN(n9094) );
  NOR3_X1 U10491 ( .A1(n9096), .A2(n9095), .A3(n9094), .ZN(n9097) );
  AND4_X1 U10492 ( .A1(n9100), .A2(n9099), .A3(n9098), .A4(n9097), .ZN(n9101)
         );
  AND4_X1 U10493 ( .A1(n9104), .A2(n9103), .A3(n9102), .A4(n9101), .ZN(n9128)
         );
  INV_X1 U10494 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9690) );
  AOI22_X1 U10495 ( .A1(n7473), .A2(keyinput13), .B1(n9690), .B2(keyinput41), 
        .ZN(n9105) );
  OAI221_X1 U10496 ( .B1(n7473), .B2(keyinput13), .C1(n9690), .C2(keyinput41), 
        .A(n9105), .ZN(n9115) );
  INV_X1 U10497 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n9664) );
  AOI22_X1 U10498 ( .A1(n9107), .A2(keyinput27), .B1(n9664), .B2(keyinput5), 
        .ZN(n9106) );
  OAI221_X1 U10499 ( .B1(n9107), .B2(keyinput27), .C1(n9664), .C2(keyinput5), 
        .A(n9106), .ZN(n9114) );
  AOI22_X1 U10500 ( .A1(n9386), .A2(keyinput14), .B1(n6091), .B2(keyinput9), 
        .ZN(n9108) );
  OAI221_X1 U10501 ( .B1(n9386), .B2(keyinput14), .C1(n6091), .C2(keyinput9), 
        .A(n9108), .ZN(n9113) );
  AOI22_X1 U10502 ( .A1(n9111), .A2(keyinput35), .B1(keyinput44), .B2(n9110), 
        .ZN(n9109) );
  OAI221_X1 U10503 ( .B1(n9111), .B2(keyinput35), .C1(n9110), .C2(keyinput44), 
        .A(n9109), .ZN(n9112) );
  NOR4_X1 U10504 ( .A1(n9115), .A2(n9114), .A3(n9113), .A4(n9112), .ZN(n9127)
         );
  AOI22_X1 U10505 ( .A1(n9117), .A2(keyinput29), .B1(n9249), .B2(keyinput7), 
        .ZN(n9116) );
  OAI221_X1 U10506 ( .B1(n9117), .B2(keyinput29), .C1(n9249), .C2(keyinput7), 
        .A(n9116), .ZN(n9125) );
  AOI22_X1 U10507 ( .A1(n5019), .A2(keyinput11), .B1(n9141), .B2(keyinput15), 
        .ZN(n9118) );
  OAI221_X1 U10508 ( .B1(n5019), .B2(keyinput11), .C1(n9141), .C2(keyinput15), 
        .A(n9118), .ZN(n9124) );
  INV_X1 U10509 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n9662) );
  AOI22_X1 U10510 ( .A1(n9992), .A2(keyinput26), .B1(n9662), .B2(keyinput8), 
        .ZN(n9119) );
  OAI221_X1 U10511 ( .B1(n9992), .B2(keyinput26), .C1(n9662), .C2(keyinput8), 
        .A(n9119), .ZN(n9123) );
  INV_X1 U10512 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9618) );
  AOI22_X1 U10513 ( .A1(n9121), .A2(keyinput23), .B1(keyinput28), .B2(n9618), 
        .ZN(n9120) );
  OAI221_X1 U10514 ( .B1(n9121), .B2(keyinput23), .C1(n9618), .C2(keyinput28), 
        .A(n9120), .ZN(n9122) );
  NOR4_X1 U10515 ( .A1(n9125), .A2(n9124), .A3(n9123), .A4(n9122), .ZN(n9126)
         );
  NAND3_X1 U10516 ( .A1(n9128), .A2(n9127), .A3(n9126), .ZN(n9156) );
  NAND4_X1 U10517 ( .A1(P2_D_REG_0__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .A3(P1_DATAO_REG_29__SCAN_IN), .A4(P2_ADDR_REG_10__SCAN_IN), .ZN(n9132) );
  NAND4_X1 U10518 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_REG1_REG_25__SCAN_IN), 
        .A3(P2_REG2_REG_23__SCAN_IN), .A4(P2_REG1_REG_31__SCAN_IN), .ZN(n9131)
         );
  NAND4_X1 U10519 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), 
        .A3(P2_D_REG_10__SCAN_IN), .A4(P2_REG1_REG_12__SCAN_IN), .ZN(n9130) );
  NAND4_X1 U10520 ( .A1(P1_REG0_REG_27__SCAN_IN), .A2(P2_REG1_REG_16__SCAN_IN), 
        .A3(P2_REG2_REG_15__SCAN_IN), .A4(SI_31_), .ZN(n9129) );
  NOR4_X1 U10521 ( .A1(n9132), .A2(n9131), .A3(n9130), .A4(n9129), .ZN(n9136)
         );
  NOR4_X1 U10522 ( .A1(P2_REG2_REG_31__SCAN_IN), .A2(P2_REG1_REG_15__SCAN_IN), 
        .A3(P2_ADDR_REG_18__SCAN_IN), .A4(n5019), .ZN(n9135) );
  NOR4_X1 U10523 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_REG0_REG_9__SCAN_IN), 
        .A3(P1_REG2_REG_5__SCAN_IN), .A4(P1_REG2_REG_2__SCAN_IN), .ZN(n9134)
         );
  NOR4_X1 U10524 ( .A1(P1_REG2_REG_26__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_13__SCAN_IN), .A4(P1_ADDR_REG_12__SCAN_IN), .ZN(n9133)
         );
  AND4_X1 U10525 ( .A1(n9136), .A2(n9135), .A3(n9134), .A4(n9133), .ZN(n9154)
         );
  NOR4_X1 U10526 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .A3(P2_ADDR_REG_5__SCAN_IN), .A4(n9137), .ZN(n9153) );
  NOR4_X1 U10527 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_REG1_REG_22__SCAN_IN), 
        .A3(P2_REG0_REG_11__SCAN_IN), .A4(P2_REG1_REG_7__SCAN_IN), .ZN(n9152)
         );
  NAND4_X1 U10528 ( .A1(SI_17_), .A2(SI_15_), .A3(SI_12_), .A4(n9138), .ZN(
        n9140) );
  NAND3_X1 U10529 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(
        P1_DATAO_REG_10__SCAN_IN), .A3(SI_9_), .ZN(n9139) );
  NOR3_X1 U10530 ( .A1(SI_6_), .A2(n9140), .A3(n9139), .ZN(n9150) );
  INV_X1 U10531 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9475) );
  NOR3_X1 U10532 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(P1_REG0_REG_14__SCAN_IN), 
        .A3(P1_REG1_REG_7__SCAN_IN), .ZN(n9146) );
  NOR4_X1 U10533 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(P1_REG0_REG_20__SCAN_IN), 
        .A3(P1_REG1_REG_17__SCAN_IN), .A4(n9249), .ZN(n9145) );
  NOR4_X1 U10534 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P1_DATAO_REG_25__SCAN_IN), 
        .A3(P2_REG0_REG_27__SCAN_IN), .A4(n9141), .ZN(n9144) );
  NOR4_X1 U10535 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_REG3_REG_13__SCAN_IN), 
        .A3(P1_REG1_REG_22__SCAN_IN), .A4(n9142), .ZN(n9143) );
  NAND4_X1 U10536 ( .A1(n9146), .A2(n9145), .A3(n9144), .A4(n9143), .ZN(n9147)
         );
  NOR4_X1 U10537 ( .A1(n9148), .A2(n9662), .A3(n9475), .A4(n9147), .ZN(n9149)
         );
  AND4_X1 U10538 ( .A1(n9150), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(n9149), .ZN(n9151) );
  NAND4_X1 U10539 ( .A1(n9154), .A2(n9153), .A3(n9152), .A4(n9151), .ZN(n9155)
         );
  XNOR2_X1 U10540 ( .A(n9156), .B(n9155), .ZN(n9157) );
  XNOR2_X1 U10541 ( .A(n9158), .B(n9157), .ZN(P1_U3270) );
  XNOR2_X1 U10542 ( .A(n9160), .B(n9161), .ZN(n9455) );
  AOI21_X1 U10543 ( .B1(n9163), .B2(n9162), .A(n9161), .ZN(n9169) );
  NAND2_X1 U10544 ( .A1(n9164), .A2(n9301), .ZN(n9168) );
  AOI22_X1 U10545 ( .A1(n9166), .A2(n9222), .B1(n9224), .B2(n9165), .ZN(n9167)
         );
  OAI21_X1 U10546 ( .B1(n9169), .B2(n9168), .A(n9167), .ZN(n9358) );
  AOI211_X1 U10547 ( .C1(n9452), .C2(n9187), .A(n9308), .B(n9170), .ZN(n9357)
         );
  NAND2_X1 U10548 ( .A1(n9357), .A2(n9317), .ZN(n9174) );
  INV_X1 U10549 ( .A(n9171), .ZN(n9172) );
  AOI22_X1 U10550 ( .A1(n9172), .A2(n9312), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n4251), .ZN(n9173) );
  OAI211_X1 U10551 ( .C1(n9175), .C2(n9315), .A(n9174), .B(n9173), .ZN(n9176)
         );
  AOI21_X1 U10552 ( .B1(n9306), .B2(n9358), .A(n9176), .ZN(n9177) );
  OAI21_X1 U10553 ( .B1(n9455), .B2(n9294), .A(n9177), .ZN(P1_U3271) );
  XOR2_X1 U10554 ( .A(n9181), .B(n9178), .Z(n9364) );
  INV_X1 U10555 ( .A(n9364), .ZN(n9195) );
  NAND2_X1 U10556 ( .A1(n9180), .A2(n9179), .ZN(n9183) );
  INV_X1 U10557 ( .A(n9181), .ZN(n9182) );
  XNOR2_X1 U10558 ( .A(n9183), .B(n9182), .ZN(n9184) );
  NAND2_X1 U10559 ( .A1(n9184), .A2(n9301), .ZN(n9186) );
  NAND2_X1 U10560 ( .A1(n9186), .A2(n9185), .ZN(n9362) );
  INV_X1 U10561 ( .A(n9187), .ZN(n9188) );
  AOI211_X1 U10562 ( .C1(n9189), .C2(n9203), .A(n9308), .B(n9188), .ZN(n9363)
         );
  NAND2_X1 U10563 ( .A1(n9363), .A2(n9317), .ZN(n9192) );
  AOI22_X1 U10564 ( .A1(n9190), .A2(n9312), .B1(n4251), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n9191) );
  OAI211_X1 U10565 ( .C1(n9459), .C2(n9315), .A(n9192), .B(n9191), .ZN(n9193)
         );
  AOI21_X1 U10566 ( .B1(n9306), .B2(n9362), .A(n9193), .ZN(n9194) );
  OAI21_X1 U10567 ( .B1(n9195), .B2(n9294), .A(n9194), .ZN(P1_U3272) );
  XNOR2_X1 U10568 ( .A(n9196), .B(n9197), .ZN(n9369) );
  INV_X1 U10569 ( .A(n9369), .ZN(n9212) );
  INV_X1 U10570 ( .A(n9197), .ZN(n9198) );
  XNOR2_X1 U10571 ( .A(n9199), .B(n9198), .ZN(n9200) );
  NAND2_X1 U10572 ( .A1(n9200), .A2(n9301), .ZN(n9202) );
  NAND2_X1 U10573 ( .A1(n9202), .A2(n9201), .ZN(n9367) );
  INV_X1 U10574 ( .A(n9203), .ZN(n9204) );
  AOI211_X1 U10575 ( .C1(n9205), .C2(n4518), .A(n9308), .B(n9204), .ZN(n9368)
         );
  NAND2_X1 U10576 ( .A1(n9368), .A2(n9317), .ZN(n9209) );
  INV_X1 U10577 ( .A(n9206), .ZN(n9207) );
  AOI22_X1 U10578 ( .A1(n4251), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9207), .B2(
        n9312), .ZN(n9208) );
  OAI211_X1 U10579 ( .C1(n9463), .C2(n9315), .A(n9209), .B(n9208), .ZN(n9210)
         );
  AOI21_X1 U10580 ( .B1(n9306), .B2(n9367), .A(n9210), .ZN(n9211) );
  OAI21_X1 U10581 ( .B1(n9212), .B2(n9294), .A(n9211), .ZN(P1_U3273) );
  XNOR2_X1 U10582 ( .A(n9214), .B(n9213), .ZN(n9377) );
  AOI21_X1 U10583 ( .B1(n9372), .B2(n9233), .A(n9215), .ZN(n9374) );
  INV_X1 U10584 ( .A(n9216), .ZN(n9217) );
  AOI22_X1 U10585 ( .A1(n4251), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9217), .B2(
        n9312), .ZN(n9218) );
  OAI21_X1 U10586 ( .B1(n9219), .B2(n9315), .A(n9218), .ZN(n9228) );
  XNOR2_X1 U10587 ( .A(n9221), .B(n9220), .ZN(n9226) );
  AOI222_X1 U10588 ( .A1(n9301), .A2(n9226), .B1(n9225), .B2(n9224), .C1(n9223), .C2(n9222), .ZN(n9376) );
  NOR2_X1 U10589 ( .A1(n9376), .A2(n4251), .ZN(n9227) );
  AOI211_X1 U10590 ( .C1(n9374), .C2(n9229), .A(n9228), .B(n9227), .ZN(n9230)
         );
  OAI21_X1 U10591 ( .B1(n9377), .B2(n9294), .A(n9230), .ZN(P1_U3274) );
  XNOR2_X1 U10592 ( .A(n9231), .B(n9239), .ZN(n9468) );
  INV_X1 U10593 ( .A(n9233), .ZN(n9234) );
  AOI211_X1 U10594 ( .C1(n9380), .C2(n9248), .A(n9308), .B(n9234), .ZN(n9379)
         );
  OAI22_X1 U10595 ( .A1(n6228), .A2(n9315), .B1(n9235), .B2(n9306), .ZN(n9236)
         );
  AOI21_X1 U10596 ( .B1(n9379), .B2(n9317), .A(n9236), .ZN(n9246) );
  NAND2_X1 U10597 ( .A1(n9238), .A2(n9237), .ZN(n9240) );
  XNOR2_X1 U10598 ( .A(n9240), .B(n9239), .ZN(n9242) );
  OAI21_X1 U10599 ( .B1(n9242), .B2(n9283), .A(n9241), .ZN(n9378) );
  NOR2_X1 U10600 ( .A1(n9243), .A2(n9257), .ZN(n9244) );
  OAI21_X1 U10601 ( .B1(n9378), .B2(n9244), .A(n9306), .ZN(n9245) );
  OAI211_X1 U10602 ( .C1(n9468), .C2(n9294), .A(n9246), .B(n9245), .ZN(
        P1_U3275) );
  XOR2_X1 U10603 ( .A(n9252), .B(n9247), .Z(n9473) );
  AOI211_X1 U10604 ( .C1(n9385), .C2(n9268), .A(n9308), .B(n9232), .ZN(n9384)
         );
  OAI22_X1 U10605 ( .A1(n9250), .A2(n9315), .B1(n9249), .B2(n9306), .ZN(n9251)
         );
  AOI21_X1 U10606 ( .B1(n9384), .B2(n9317), .A(n9251), .ZN(n9261) );
  XNOR2_X1 U10607 ( .A(n9253), .B(n9252), .ZN(n9256) );
  INV_X1 U10608 ( .A(n9254), .ZN(n9255) );
  OAI21_X1 U10609 ( .B1(n9256), .B2(n9283), .A(n9255), .ZN(n9383) );
  NOR2_X1 U10610 ( .A1(n9258), .A2(n9257), .ZN(n9259) );
  OAI21_X1 U10611 ( .B1(n9383), .B2(n9259), .A(n9306), .ZN(n9260) );
  OAI211_X1 U10612 ( .C1(n9473), .C2(n9294), .A(n9261), .B(n9260), .ZN(
        P1_U3276) );
  XNOR2_X1 U10613 ( .A(n9262), .B(n4689), .ZN(n9391) );
  INV_X1 U10614 ( .A(n9391), .ZN(n9276) );
  XNOR2_X1 U10615 ( .A(n9264), .B(n9263), .ZN(n9265) );
  NAND2_X1 U10616 ( .A1(n9265), .A2(n9301), .ZN(n9267) );
  NAND2_X1 U10617 ( .A1(n9267), .A2(n9266), .ZN(n9389) );
  INV_X1 U10618 ( .A(n9268), .ZN(n9269) );
  AOI211_X1 U10619 ( .C1(n9270), .C2(n4526), .A(n9308), .B(n9269), .ZN(n9390)
         );
  NAND2_X1 U10620 ( .A1(n9390), .A2(n9317), .ZN(n9273) );
  AOI22_X1 U10621 ( .A1(n4251), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9271), .B2(
        n9312), .ZN(n9272) );
  OAI211_X1 U10622 ( .C1(n9477), .C2(n9315), .A(n9273), .B(n9272), .ZN(n9274)
         );
  AOI21_X1 U10623 ( .B1(n9306), .B2(n9389), .A(n9274), .ZN(n9275) );
  OAI21_X1 U10624 ( .B1(n9276), .B2(n9294), .A(n9275), .ZN(P1_U3277) );
  XNOR2_X1 U10625 ( .A(n9277), .B(n9281), .ZN(n9398) );
  INV_X1 U10626 ( .A(n9278), .ZN(n9279) );
  AOI21_X1 U10627 ( .B1(n9281), .B2(n9280), .A(n9279), .ZN(n9282) );
  OAI222_X1 U10628 ( .A1(n9287), .A2(n9286), .B1(n9285), .B2(n9284), .C1(n9283), .C2(n9282), .ZN(n9394) );
  AOI211_X1 U10629 ( .C1(n9396), .C2(n9307), .A(n9308), .B(n9288), .ZN(n9395)
         );
  NAND2_X1 U10630 ( .A1(n9395), .A2(n9317), .ZN(n9291) );
  AOI22_X1 U10631 ( .A1(n4251), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9289), .B2(
        n9312), .ZN(n9290) );
  OAI211_X1 U10632 ( .C1(n4524), .C2(n9315), .A(n9291), .B(n9290), .ZN(n9292)
         );
  AOI21_X1 U10633 ( .B1(n9394), .B2(n9306), .A(n9292), .ZN(n9293) );
  OAI21_X1 U10634 ( .B1(n9398), .B2(n9294), .A(n9293), .ZN(P1_U3278) );
  AOI21_X1 U10635 ( .B1(n9296), .B2(n9299), .A(n9295), .ZN(n9399) );
  NAND2_X1 U10636 ( .A1(n9298), .A2(n9297), .ZN(n9300) );
  XNOR2_X1 U10637 ( .A(n9300), .B(n9299), .ZN(n9302) );
  NAND2_X1 U10638 ( .A1(n9302), .A2(n9301), .ZN(n9303) );
  OAI211_X1 U10639 ( .C1(n9399), .C2(n9305), .A(n9304), .B(n9303), .ZN(n9400)
         );
  NAND2_X1 U10640 ( .A1(n9400), .A2(n9306), .ZN(n9319) );
  INV_X1 U10641 ( .A(n9307), .ZN(n9309) );
  AOI211_X1 U10642 ( .C1(n9311), .C2(n9310), .A(n9309), .B(n9308), .ZN(n9401)
         );
  AOI22_X1 U10643 ( .A1(n4251), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9313), .B2(
        n9312), .ZN(n9314) );
  OAI21_X1 U10644 ( .B1(n9484), .B2(n9315), .A(n9314), .ZN(n9316) );
  AOI21_X1 U10645 ( .B1(n9401), .B2(n9317), .A(n9316), .ZN(n9318) );
  OAI211_X1 U10646 ( .C1(n9399), .C2(n9320), .A(n9319), .B(n9318), .ZN(
        P1_U3279) );
  INV_X1 U10647 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9323) );
  AND2_X1 U10648 ( .A1(n9322), .A2(n9321), .ZN(n9413) );
  MUX2_X1 U10649 ( .A(n9323), .B(n9413), .S(n9708), .Z(n9324) );
  OAI21_X1 U10650 ( .B1(n9416), .B2(n9406), .A(n9324), .ZN(P1_U3552) );
  NAND2_X1 U10651 ( .A1(n9417), .A2(n9360), .ZN(n9327) );
  OAI211_X1 U10652 ( .C1(n9420), .C2(n9388), .A(n9328), .B(n9327), .ZN(
        P1_U3551) );
  AOI211_X1 U10653 ( .C1(n9675), .C2(n9331), .A(n9330), .B(n9329), .ZN(n9421)
         );
  MUX2_X1 U10654 ( .A(n9332), .B(n9421), .S(n9708), .Z(n9333) );
  OAI21_X1 U10655 ( .B1(n9424), .B2(n9388), .A(n9333), .ZN(P1_U3550) );
  NAND2_X1 U10656 ( .A1(n9335), .A2(n9334), .ZN(n9425) );
  MUX2_X1 U10657 ( .A(n9425), .B(P1_REG1_REG_27__SCAN_IN), .S(n9706), .Z(n9336) );
  AOI21_X1 U10658 ( .B1(n9360), .B2(n9427), .A(n9336), .ZN(n9337) );
  OAI21_X1 U10659 ( .B1(n9429), .B2(n9388), .A(n9337), .ZN(P1_U3549) );
  INV_X1 U10660 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9341) );
  AOI211_X1 U10661 ( .C1(n9675), .C2(n9340), .A(n9339), .B(n9338), .ZN(n9430)
         );
  MUX2_X1 U10662 ( .A(n9341), .B(n9430), .S(n9708), .Z(n9342) );
  OAI21_X1 U10663 ( .B1(n9433), .B2(n9388), .A(n9342), .ZN(P1_U3548) );
  NAND2_X1 U10664 ( .A1(n9344), .A2(n9343), .ZN(n9434) );
  MUX2_X1 U10665 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9434), .S(n9708), .Z(n9345) );
  AOI21_X1 U10666 ( .B1(n9360), .B2(n9436), .A(n9345), .ZN(n9346) );
  OAI21_X1 U10667 ( .B1(n9438), .B2(n9388), .A(n9346), .ZN(P1_U3547) );
  NOR2_X1 U10668 ( .A1(n9348), .A2(n9347), .ZN(n9439) );
  MUX2_X1 U10669 ( .A(n9349), .B(n9439), .S(n9403), .Z(n9351) );
  NAND2_X1 U10670 ( .A1(n9442), .A2(n9360), .ZN(n9350) );
  OAI211_X1 U10671 ( .C1(n9444), .C2(n9388), .A(n9351), .B(n9350), .ZN(
        P1_U3546) );
  INV_X1 U10672 ( .A(n9352), .ZN(n9354) );
  NAND2_X1 U10673 ( .A1(n9354), .A2(n9353), .ZN(n9445) );
  MUX2_X1 U10674 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9445), .S(n9708), .Z(n9355) );
  AOI21_X1 U10675 ( .B1(n9360), .B2(n9447), .A(n9355), .ZN(n9356) );
  OAI21_X1 U10676 ( .B1(n9449), .B2(n9388), .A(n9356), .ZN(P1_U3545) );
  OR2_X1 U10677 ( .A1(n9358), .A2(n9357), .ZN(n9450) );
  MUX2_X1 U10678 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9450), .S(n9403), .Z(n9359) );
  AOI21_X1 U10679 ( .B1(n9360), .B2(n9452), .A(n9359), .ZN(n9361) );
  OAI21_X1 U10680 ( .B1(n9455), .B2(n9388), .A(n9361), .ZN(P1_U3544) );
  AOI211_X1 U10681 ( .C1(n9364), .C2(n9689), .A(n9363), .B(n9362), .ZN(n9456)
         );
  MUX2_X1 U10682 ( .A(n9365), .B(n9456), .S(n9403), .Z(n9366) );
  OAI21_X1 U10683 ( .B1(n9459), .B2(n9406), .A(n9366), .ZN(P1_U3543) );
  INV_X1 U10684 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9370) );
  AOI211_X1 U10685 ( .C1(n9369), .C2(n9689), .A(n9368), .B(n9367), .ZN(n9460)
         );
  MUX2_X1 U10686 ( .A(n9370), .B(n9460), .S(n9403), .Z(n9371) );
  OAI21_X1 U10687 ( .B1(n9463), .B2(n9406), .A(n9371), .ZN(P1_U3542) );
  AOI22_X1 U10688 ( .A1(n9374), .A2(n9373), .B1(n9675), .B2(n9372), .ZN(n9375)
         );
  OAI211_X1 U10689 ( .C1(n9377), .C2(n9411), .A(n9376), .B(n9375), .ZN(n9464)
         );
  MUX2_X1 U10690 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9464), .S(n9403), .Z(
        P1_U3541) );
  AOI211_X1 U10691 ( .C1(n9675), .C2(n9380), .A(n9379), .B(n9378), .ZN(n9465)
         );
  MUX2_X1 U10692 ( .A(n9381), .B(n9465), .S(n9403), .Z(n9382) );
  OAI21_X1 U10693 ( .B1(n9468), .B2(n9388), .A(n9382), .ZN(P1_U3540) );
  AOI211_X1 U10694 ( .C1(n9675), .C2(n9385), .A(n9384), .B(n9383), .ZN(n9469)
         );
  MUX2_X1 U10695 ( .A(n9386), .B(n9469), .S(n9403), .Z(n9387) );
  OAI21_X1 U10696 ( .B1(n9473), .B2(n9388), .A(n9387), .ZN(P1_U3539) );
  AOI211_X1 U10697 ( .C1(n9391), .C2(n9689), .A(n9390), .B(n9389), .ZN(n9474)
         );
  MUX2_X1 U10698 ( .A(n9392), .B(n9474), .S(n9403), .Z(n9393) );
  OAI21_X1 U10699 ( .B1(n9477), .B2(n9406), .A(n9393), .ZN(P1_U3538) );
  AOI211_X1 U10700 ( .C1(n9675), .C2(n9396), .A(n9395), .B(n9394), .ZN(n9397)
         );
  OAI21_X1 U10701 ( .B1(n9398), .B2(n9411), .A(n9397), .ZN(n9478) );
  MUX2_X1 U10702 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9478), .S(n9403), .Z(
        P1_U3537) );
  INV_X1 U10703 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9404) );
  INV_X1 U10704 ( .A(n9399), .ZN(n9402) );
  AOI211_X1 U10705 ( .C1(n9695), .C2(n9402), .A(n9401), .B(n9400), .ZN(n9480)
         );
  MUX2_X1 U10706 ( .A(n9404), .B(n9480), .S(n9403), .Z(n9405) );
  OAI21_X1 U10707 ( .B1(n9484), .B2(n9406), .A(n9405), .ZN(P1_U3536) );
  AOI21_X1 U10708 ( .B1(n9675), .B2(n9408), .A(n9407), .ZN(n9409) );
  OAI211_X1 U10709 ( .C1(n9412), .C2(n9411), .A(n9410), .B(n9409), .ZN(n9485)
         );
  MUX2_X1 U10710 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9485), .S(n9708), .Z(
        P1_U3535) );
  INV_X1 U10711 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9414) );
  MUX2_X1 U10712 ( .A(n9414), .B(n9413), .S(n9479), .Z(n9415) );
  OAI21_X1 U10713 ( .B1(n9416), .B2(n9483), .A(n9415), .ZN(P1_U3520) );
  NAND2_X1 U10714 ( .A1(n9417), .A2(n9453), .ZN(n9418) );
  OAI211_X1 U10715 ( .C1(n9420), .C2(n9472), .A(n9419), .B(n9418), .ZN(
        P1_U3519) );
  INV_X1 U10716 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9422) );
  MUX2_X1 U10717 ( .A(n9422), .B(n9421), .S(n9479), .Z(n9423) );
  OAI21_X1 U10718 ( .B1(n9424), .B2(n9472), .A(n9423), .ZN(P1_U3518) );
  MUX2_X1 U10719 ( .A(n9425), .B(P1_REG0_REG_27__SCAN_IN), .S(n9699), .Z(n9426) );
  AOI21_X1 U10720 ( .B1(n9453), .B2(n9427), .A(n9426), .ZN(n9428) );
  OAI21_X1 U10721 ( .B1(n9429), .B2(n9472), .A(n9428), .ZN(P1_U3517) );
  INV_X1 U10722 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9431) );
  MUX2_X1 U10723 ( .A(n9431), .B(n9430), .S(n9479), .Z(n9432) );
  OAI21_X1 U10724 ( .B1(n9433), .B2(n9472), .A(n9432), .ZN(P1_U3516) );
  MUX2_X1 U10725 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9434), .S(n9479), .Z(n9435) );
  AOI21_X1 U10726 ( .B1(n9453), .B2(n9436), .A(n9435), .ZN(n9437) );
  OAI21_X1 U10727 ( .B1(n9438), .B2(n9472), .A(n9437), .ZN(P1_U3515) );
  INV_X1 U10728 ( .A(n9439), .ZN(n9440) );
  MUX2_X1 U10729 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9440), .S(n9479), .Z(n9441) );
  AOI21_X1 U10730 ( .B1(n9453), .B2(n9442), .A(n9441), .ZN(n9443) );
  OAI21_X1 U10731 ( .B1(n9444), .B2(n9472), .A(n9443), .ZN(P1_U3514) );
  MUX2_X1 U10732 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9445), .S(n9479), .Z(n9446) );
  AOI21_X1 U10733 ( .B1(n9453), .B2(n9447), .A(n9446), .ZN(n9448) );
  OAI21_X1 U10734 ( .B1(n9449), .B2(n9472), .A(n9448), .ZN(P1_U3513) );
  MUX2_X1 U10735 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9450), .S(n9479), .Z(n9451) );
  AOI21_X1 U10736 ( .B1(n9453), .B2(n9452), .A(n9451), .ZN(n9454) );
  OAI21_X1 U10737 ( .B1(n9455), .B2(n9472), .A(n9454), .ZN(P1_U3512) );
  INV_X1 U10738 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9457) );
  MUX2_X1 U10739 ( .A(n9457), .B(n9456), .S(n9479), .Z(n9458) );
  OAI21_X1 U10740 ( .B1(n9459), .B2(n9483), .A(n9458), .ZN(P1_U3511) );
  MUX2_X1 U10741 ( .A(n9461), .B(n9460), .S(n9479), .Z(n9462) );
  OAI21_X1 U10742 ( .B1(n9463), .B2(n9483), .A(n9462), .ZN(P1_U3510) );
  MUX2_X1 U10743 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9464), .S(n9701), .Z(
        P1_U3509) );
  INV_X1 U10744 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9466) );
  MUX2_X1 U10745 ( .A(n9466), .B(n9465), .S(n9479), .Z(n9467) );
  OAI21_X1 U10746 ( .B1(n9468), .B2(n9472), .A(n9467), .ZN(P1_U3507) );
  MUX2_X1 U10747 ( .A(n9470), .B(n9469), .S(n9479), .Z(n9471) );
  OAI21_X1 U10748 ( .B1(n9473), .B2(n9472), .A(n9471), .ZN(P1_U3504) );
  MUX2_X1 U10749 ( .A(n9475), .B(n9474), .S(n9479), .Z(n9476) );
  OAI21_X1 U10750 ( .B1(n9477), .B2(n9483), .A(n9476), .ZN(P1_U3501) );
  MUX2_X1 U10751 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9478), .S(n9701), .Z(
        P1_U3498) );
  MUX2_X1 U10752 ( .A(n9481), .B(n9480), .S(n9479), .Z(n9482) );
  OAI21_X1 U10753 ( .B1(n9484), .B2(n9483), .A(n9482), .ZN(P1_U3495) );
  MUX2_X1 U10754 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9485), .S(n9701), .Z(
        P1_U3492) );
  MUX2_X1 U10755 ( .A(n9488), .B(P1_D_REG_1__SCAN_IN), .S(n9667), .Z(P1_U3440)
         );
  MUX2_X1 U10756 ( .A(n9489), .B(P1_D_REG_0__SCAN_IN), .S(n9667), .Z(P1_U3439)
         );
  NOR4_X1 U10757 ( .A1(n5536), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), .A4(
        n9490), .ZN(n9491) );
  AOI21_X1 U10758 ( .B1(n9497), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9491), .ZN(
        n9492) );
  OAI21_X1 U10759 ( .B1(n9493), .B2(n9500), .A(n9492), .ZN(P1_U3324) );
  AOI22_X1 U10760 ( .A1(n9494), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n9497), .ZN(n9495) );
  OAI21_X1 U10761 ( .B1(n9496), .B2(n9500), .A(n9495), .ZN(P1_U3325) );
  AOI22_X1 U10762 ( .A1(n9498), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n9497), .ZN(n9499) );
  OAI21_X1 U10763 ( .B1(n9501), .B2(n9500), .A(n9499), .ZN(P1_U3326) );
  MUX2_X1 U10764 ( .A(n9502), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  OAI21_X1 U10765 ( .B1(n9505), .B2(n9504), .A(n9503), .ZN(n9506) );
  AOI22_X1 U10766 ( .A1(n9506), .A2(n9884), .B1(n9874), .B2(
        P2_ADDR_REG_18__SCAN_IN), .ZN(n9523) );
  INV_X1 U10767 ( .A(n9507), .ZN(n9510) );
  AOI21_X1 U10768 ( .B1(n9510), .B2(n9509), .A(n9508), .ZN(n9515) );
  NAND3_X1 U10769 ( .A1(n9510), .A2(P2_U3893), .A3(n9509), .ZN(n9512) );
  NAND3_X1 U10770 ( .A1(n9512), .A2(n9511), .A3(n9514), .ZN(n9513) );
  OAI21_X1 U10771 ( .B1(n9515), .B2(n9514), .A(n9513), .ZN(n9522) );
  NAND2_X1 U10772 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_U3151), .ZN(n9521) );
  AOI21_X1 U10773 ( .B1(n9518), .B2(n9517), .A(n9516), .ZN(n9519) );
  OR2_X1 U10774 ( .A1(n9519), .A2(n9890), .ZN(n9520) );
  NAND4_X1 U10775 ( .A1(n9523), .A2(n9522), .A3(n9521), .A4(n9520), .ZN(
        P2_U3200) );
  INV_X1 U10776 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9534) );
  AOI211_X1 U10777 ( .C1(n9526), .C2(n9525), .A(n9524), .B(n9632), .ZN(n9531)
         );
  AOI211_X1 U10778 ( .C1(n9529), .C2(n9528), .A(n9527), .B(n9645), .ZN(n9530)
         );
  AOI211_X1 U10779 ( .C1(n4463), .C2(n9532), .A(n9531), .B(n9530), .ZN(n9533)
         );
  NAND2_X1 U10780 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9565) );
  OAI211_X1 U10781 ( .C1(n9661), .C2(n9534), .A(n9533), .B(n9565), .ZN(
        P1_U3253) );
  INV_X1 U10782 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9546) );
  AOI211_X1 U10783 ( .C1(n9537), .C2(n9536), .A(n9535), .B(n9645), .ZN(n9542)
         );
  AOI211_X1 U10784 ( .C1(n9540), .C2(n9539), .A(n9538), .B(n9632), .ZN(n9541)
         );
  AOI211_X1 U10785 ( .C1(n4463), .C2(n9543), .A(n9542), .B(n9541), .ZN(n9545)
         );
  OAI211_X1 U10786 ( .C1(n9661), .C2(n9546), .A(n9545), .B(n9544), .ZN(
        P1_U3250) );
  INV_X1 U10787 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9561) );
  AOI21_X1 U10788 ( .B1(n9549), .B2(n9548), .A(n9547), .ZN(n9550) );
  NAND2_X1 U10789 ( .A1(n9595), .A2(n9550), .ZN(n9556) );
  AOI21_X1 U10790 ( .B1(n9553), .B2(n9552), .A(n9551), .ZN(n9554) );
  NAND2_X1 U10791 ( .A1(n9648), .A2(n9554), .ZN(n9555) );
  OAI211_X1 U10792 ( .C1(n9654), .C2(n9557), .A(n9556), .B(n9555), .ZN(n9558)
         );
  INV_X1 U10793 ( .A(n9558), .ZN(n9560) );
  OAI211_X1 U10794 ( .C1(n9661), .C2(n9561), .A(n9560), .B(n9559), .ZN(
        P1_U3251) );
  OAI21_X1 U10795 ( .B1(n9564), .B2(n9563), .A(n4384), .ZN(n9574) );
  INV_X1 U10796 ( .A(n9565), .ZN(n9566) );
  AOI21_X1 U10797 ( .B1(n9568), .B2(n9567), .A(n9566), .ZN(n9569) );
  OAI21_X1 U10798 ( .B1(n9571), .B2(n9570), .A(n9569), .ZN(n9572) );
  AOI21_X1 U10799 ( .B1(n9574), .B2(n9573), .A(n9572), .ZN(n9575) );
  OAI21_X1 U10800 ( .B1(n9577), .B2(n9576), .A(n9575), .ZN(P1_U3217) );
  XNOR2_X1 U10801 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10802 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10803 ( .A(n9578), .ZN(n9581) );
  AOI211_X1 U10804 ( .C1(n9581), .C2(n9580), .A(n9579), .B(n9645), .ZN(n9586)
         );
  AOI211_X1 U10805 ( .C1(n9584), .C2(n9583), .A(n9632), .B(n9582), .ZN(n9585)
         );
  AOI211_X1 U10806 ( .C1(n4463), .C2(n9587), .A(n9586), .B(n9585), .ZN(n9589)
         );
  OAI211_X1 U10807 ( .C1(n9661), .C2(n9590), .A(n9589), .B(n9588), .ZN(
        P1_U3249) );
  INV_X1 U10808 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9606) );
  AOI21_X1 U10809 ( .B1(n9593), .B2(n9592), .A(n9591), .ZN(n9594) );
  NAND2_X1 U10810 ( .A1(n9595), .A2(n9594), .ZN(n9601) );
  AOI21_X1 U10811 ( .B1(n9598), .B2(n9597), .A(n9596), .ZN(n9599) );
  NAND2_X1 U10812 ( .A1(n9648), .A2(n9599), .ZN(n9600) );
  OAI211_X1 U10813 ( .C1(n9654), .C2(n9602), .A(n9601), .B(n9600), .ZN(n9603)
         );
  INV_X1 U10814 ( .A(n9603), .ZN(n9605) );
  OAI211_X1 U10815 ( .C1(n9661), .C2(n9606), .A(n9605), .B(n9604), .ZN(
        P1_U3254) );
  AOI211_X1 U10816 ( .C1(n9609), .C2(n9608), .A(n9632), .B(n9607), .ZN(n9614)
         );
  AOI211_X1 U10817 ( .C1(n9612), .C2(n9611), .A(n9645), .B(n9610), .ZN(n9613)
         );
  AOI211_X1 U10818 ( .C1(n4463), .C2(n9615), .A(n9614), .B(n9613), .ZN(n9617)
         );
  OAI211_X1 U10819 ( .C1(n9618), .C2(n9661), .A(n9617), .B(n9616), .ZN(
        P1_U3256) );
  INV_X1 U10820 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9630) );
  AOI211_X1 U10821 ( .C1(n9621), .C2(n9620), .A(n9619), .B(n9645), .ZN(n9626)
         );
  AOI211_X1 U10822 ( .C1(n9624), .C2(n9623), .A(n9632), .B(n9622), .ZN(n9625)
         );
  AOI211_X1 U10823 ( .C1(n4463), .C2(n9627), .A(n9626), .B(n9625), .ZN(n9629)
         );
  OAI211_X1 U10824 ( .C1(n9661), .C2(n9630), .A(n9629), .B(n9628), .ZN(
        P1_U3257) );
  INV_X1 U10825 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9644) );
  INV_X1 U10826 ( .A(n9631), .ZN(n9641) );
  AOI211_X1 U10827 ( .C1(n9635), .C2(n9634), .A(n9633), .B(n9632), .ZN(n9640)
         );
  AOI211_X1 U10828 ( .C1(n9638), .C2(n9637), .A(n9636), .B(n9645), .ZN(n9639)
         );
  AOI211_X1 U10829 ( .C1(n4463), .C2(n9641), .A(n9640), .B(n9639), .ZN(n9643)
         );
  OAI211_X1 U10830 ( .C1(n9661), .C2(n9644), .A(n9643), .B(n9642), .ZN(
        P1_U3258) );
  AOI21_X1 U10831 ( .B1(n9647), .B2(n9646), .A(n9645), .ZN(n9657) );
  OAI211_X1 U10832 ( .C1(n9651), .C2(n9650), .A(n9649), .B(n9648), .ZN(n9652)
         );
  OAI21_X1 U10833 ( .B1(n9654), .B2(n9653), .A(n9652), .ZN(n9655) );
  AOI21_X1 U10834 ( .B1(n9657), .B2(n9656), .A(n9655), .ZN(n9659) );
  NAND2_X1 U10835 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3086), .ZN(n9658) );
  OAI211_X1 U10836 ( .C1(n9661), .C2(n9660), .A(n9659), .B(n9658), .ZN(
        P1_U3261) );
  AND2_X1 U10837 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9667), .ZN(P1_U3294) );
  AND2_X1 U10838 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9667), .ZN(P1_U3295) );
  AND2_X1 U10839 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9667), .ZN(P1_U3296) );
  AND2_X1 U10840 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9667), .ZN(P1_U3297) );
  AND2_X1 U10841 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9667), .ZN(P1_U3298) );
  AND2_X1 U10842 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9667), .ZN(P1_U3299) );
  AND2_X1 U10843 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9667), .ZN(P1_U3300) );
  AND2_X1 U10844 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9667), .ZN(P1_U3301) );
  AND2_X1 U10845 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9667), .ZN(P1_U3302) );
  AND2_X1 U10846 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9667), .ZN(P1_U3303) );
  INV_X1 U10847 ( .A(n9667), .ZN(n9666) );
  NOR2_X1 U10848 ( .A1(n9666), .A2(n9662), .ZN(P1_U3304) );
  AND2_X1 U10849 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9667), .ZN(P1_U3305) );
  NOR2_X1 U10850 ( .A1(n9666), .A2(n9663), .ZN(P1_U3306) );
  AND2_X1 U10851 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9667), .ZN(P1_U3307) );
  AND2_X1 U10852 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9667), .ZN(P1_U3308) );
  AND2_X1 U10853 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9667), .ZN(P1_U3309) );
  AND2_X1 U10854 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9667), .ZN(P1_U3310) );
  AND2_X1 U10855 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9667), .ZN(P1_U3311) );
  AND2_X1 U10856 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9667), .ZN(P1_U3312) );
  NOR2_X1 U10857 ( .A1(n9666), .A2(n9664), .ZN(P1_U3313) );
  AND2_X1 U10858 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9667), .ZN(P1_U3314) );
  AND2_X1 U10859 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9667), .ZN(P1_U3315) );
  AND2_X1 U10860 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9667), .ZN(P1_U3316) );
  AND2_X1 U10861 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9667), .ZN(P1_U3317) );
  AND2_X1 U10862 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9667), .ZN(P1_U3318) );
  AND2_X1 U10863 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9667), .ZN(P1_U3319) );
  AND2_X1 U10864 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9667), .ZN(P1_U3320) );
  AND2_X1 U10865 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9667), .ZN(P1_U3321) );
  NOR2_X1 U10866 ( .A1(n9666), .A2(n9665), .ZN(P1_U3322) );
  AND2_X1 U10867 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9667), .ZN(P1_U3323) );
  INV_X1 U10868 ( .A(n9675), .ZN(n9692) );
  OAI21_X1 U10869 ( .B1(n9669), .B2(n9692), .A(n9668), .ZN(n9670) );
  AOI21_X1 U10870 ( .B1(n9671), .B2(n9695), .A(n9670), .ZN(n9672) );
  AND2_X1 U10871 ( .A1(n9673), .A2(n9672), .ZN(n9702) );
  INV_X1 U10872 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9674) );
  AOI22_X1 U10873 ( .A1(n9701), .A2(n9702), .B1(n9674), .B2(n9699), .ZN(
        P1_U3456) );
  NAND2_X1 U10874 ( .A1(n9676), .A2(n9675), .ZN(n9677) );
  NAND2_X1 U10875 ( .A1(n9678), .A2(n9677), .ZN(n9679) );
  AOI21_X1 U10876 ( .B1(n9680), .B2(n9695), .A(n9679), .ZN(n9681) );
  AND2_X1 U10877 ( .A1(n9682), .A2(n9681), .ZN(n9703) );
  INV_X1 U10878 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9683) );
  AOI22_X1 U10879 ( .A1(n9701), .A2(n9703), .B1(n9683), .B2(n9699), .ZN(
        P1_U3474) );
  OAI21_X1 U10880 ( .B1(n9685), .B2(n9692), .A(n9684), .ZN(n9687) );
  AOI211_X1 U10881 ( .C1(n9689), .C2(n9688), .A(n9687), .B(n9686), .ZN(n9705)
         );
  AOI22_X1 U10882 ( .A1(n9701), .A2(n9705), .B1(n9690), .B2(n9699), .ZN(
        P1_U3480) );
  OAI21_X1 U10883 ( .B1(n9693), .B2(n9692), .A(n9691), .ZN(n9694) );
  AOI21_X1 U10884 ( .B1(n9696), .B2(n9695), .A(n9694), .ZN(n9697) );
  AND2_X1 U10885 ( .A1(n9698), .A2(n9697), .ZN(n9707) );
  INV_X1 U10886 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9700) );
  AOI22_X1 U10887 ( .A1(n9701), .A2(n9707), .B1(n9700), .B2(n9699), .ZN(
        P1_U3486) );
  AOI22_X1 U10888 ( .A1(n9708), .A2(n9702), .B1(n6542), .B2(n9706), .ZN(
        P1_U3523) );
  AOI22_X1 U10889 ( .A1(n9708), .A2(n9703), .B1(n6546), .B2(n9706), .ZN(
        P1_U3529) );
  AOI22_X1 U10890 ( .A1(n9708), .A2(n9705), .B1(n9704), .B2(n9706), .ZN(
        P1_U3531) );
  AOI22_X1 U10891 ( .A1(n9708), .A2(n9707), .B1(n7007), .B2(n9706), .ZN(
        P1_U3533) );
  INV_X1 U10892 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n9719) );
  OAI211_X1 U10893 ( .C1(n9711), .C2(n9710), .A(n9709), .B(n9883), .ZN(n9718)
         );
  OAI21_X1 U10894 ( .B1(n9714), .B2(n9713), .A(n9712), .ZN(n9716) );
  AOI22_X1 U10895 ( .A1(n9754), .A2(n9716), .B1(n4250), .B2(n9875), .ZN(n9717)
         );
  OAI211_X1 U10896 ( .C1(n9720), .C2(n9719), .A(n9718), .B(n9717), .ZN(n9721)
         );
  INV_X1 U10897 ( .A(n9721), .ZN(n9726) );
  XNOR2_X1 U10898 ( .A(n9723), .B(n9722), .ZN(n9724) );
  NAND2_X1 U10899 ( .A1(n9884), .A2(n9724), .ZN(n9725) );
  OAI211_X1 U10900 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n4886), .A(n9726), .B(
        n9725), .ZN(P2_U3184) );
  XNOR2_X1 U10901 ( .A(n9727), .B(P2_REG2_REG_7__SCAN_IN), .ZN(n9735) );
  AOI21_X1 U10902 ( .B1(n9875), .B2(n9729), .A(n9728), .ZN(n9734) );
  XNOR2_X1 U10903 ( .A(n9730), .B(P2_REG1_REG_7__SCAN_IN), .ZN(n9731) );
  OR2_X1 U10904 ( .A1(n9732), .A2(n9731), .ZN(n9733) );
  OAI211_X1 U10905 ( .C1(n9890), .C2(n9735), .A(n9734), .B(n9733), .ZN(n9736)
         );
  INV_X1 U10906 ( .A(n9736), .ZN(n9741) );
  XNOR2_X1 U10907 ( .A(n9738), .B(n9737), .ZN(n9739) );
  AOI22_X1 U10908 ( .A1(n9739), .A2(n9883), .B1(n9874), .B2(
        P2_ADDR_REG_7__SCAN_IN), .ZN(n9740) );
  NAND2_X1 U10909 ( .A1(n9741), .A2(n9740), .ZN(P2_U3189) );
  AOI21_X1 U10910 ( .B1(n9743), .B2(n9875), .A(n9742), .ZN(n9760) );
  OAI21_X1 U10911 ( .B1(n9746), .B2(n9745), .A(n9744), .ZN(n9747) );
  AOI22_X1 U10912 ( .A1(n9747), .A2(n9883), .B1(n9874), .B2(
        P2_ADDR_REG_8__SCAN_IN), .ZN(n9759) );
  OAI21_X1 U10913 ( .B1(n9750), .B2(n9749), .A(n9748), .ZN(n9751) );
  NAND2_X1 U10914 ( .A1(n9751), .A2(n9884), .ZN(n9758) );
  NOR2_X1 U10915 ( .A1(n9753), .A2(n9752), .ZN(n9756) );
  OAI21_X1 U10916 ( .B1(n9756), .B2(n9755), .A(n9754), .ZN(n9757) );
  NAND4_X1 U10917 ( .A1(n9760), .A2(n9759), .A3(n9758), .A4(n9757), .ZN(
        P2_U3190) );
  AOI22_X1 U10918 ( .A1(n9761), .A2(n9875), .B1(P2_ADDR_REG_10__SCAN_IN), .B2(
        n9874), .ZN(n9777) );
  OAI21_X1 U10919 ( .B1(n9764), .B2(n9763), .A(n9762), .ZN(n9769) );
  OAI21_X1 U10920 ( .B1(n9767), .B2(n9766), .A(n9765), .ZN(n9768) );
  AOI22_X1 U10921 ( .A1(n9769), .A2(n9883), .B1(n9884), .B2(n9768), .ZN(n9776)
         );
  AOI21_X1 U10922 ( .B1(n9772), .B2(n9771), .A(n9770), .ZN(n9773) );
  OR2_X1 U10923 ( .A1(n9773), .A2(n9890), .ZN(n9774) );
  NAND4_X1 U10924 ( .A1(n9777), .A2(n9776), .A3(n9775), .A4(n9774), .ZN(
        P2_U3192) );
  AOI22_X1 U10925 ( .A1(n9874), .A2(P2_ADDR_REG_11__SCAN_IN), .B1(n9778), .B2(
        n9875), .ZN(n9793) );
  OAI21_X1 U10926 ( .B1(n9780), .B2(P2_REG1_REG_11__SCAN_IN), .A(n9779), .ZN(
        n9785) );
  OAI21_X1 U10927 ( .B1(n9783), .B2(n9782), .A(n9781), .ZN(n9784) );
  AOI22_X1 U10928 ( .A1(n9785), .A2(n9884), .B1(n9883), .B2(n9784), .ZN(n9792)
         );
  AOI21_X1 U10929 ( .B1(n9788), .B2(n9787), .A(n9786), .ZN(n9789) );
  OR2_X1 U10930 ( .A1(n9789), .A2(n9890), .ZN(n9790) );
  NAND4_X1 U10931 ( .A1(n9793), .A2(n9792), .A3(n9791), .A4(n9790), .ZN(
        P2_U3193) );
  AOI22_X1 U10932 ( .A1(n9794), .A2(n9875), .B1(n9874), .B2(
        P2_ADDR_REG_12__SCAN_IN), .ZN(n9809) );
  OAI21_X1 U10933 ( .B1(n9797), .B2(n9796), .A(n9795), .ZN(n9802) );
  OAI21_X1 U10934 ( .B1(n9800), .B2(n9799), .A(n9798), .ZN(n9801) );
  AOI22_X1 U10935 ( .A1(n9802), .A2(n9884), .B1(n9883), .B2(n9801), .ZN(n9808)
         );
  AOI21_X1 U10936 ( .B1(n4287), .B2(n9804), .A(n9803), .ZN(n9805) );
  OR2_X1 U10937 ( .A1(n9805), .A2(n9890), .ZN(n9806) );
  NAND4_X1 U10938 ( .A1(n9809), .A2(n9808), .A3(n9807), .A4(n9806), .ZN(
        P2_U3194) );
  AOI22_X1 U10939 ( .A1(n9810), .A2(n9875), .B1(n9874), .B2(
        P2_ADDR_REG_13__SCAN_IN), .ZN(n9824) );
  OAI21_X1 U10940 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n9812), .A(n9811), .ZN(
        n9817) );
  OAI21_X1 U10941 ( .B1(n9815), .B2(n9814), .A(n9813), .ZN(n9816) );
  AOI22_X1 U10942 ( .A1(n9817), .A2(n9884), .B1(n9883), .B2(n9816), .ZN(n9823)
         );
  AOI21_X1 U10943 ( .B1(n9819), .B2(n5098), .A(n9818), .ZN(n9820) );
  OR2_X1 U10944 ( .A1(n9890), .A2(n9820), .ZN(n9821) );
  NAND4_X1 U10945 ( .A1(n9824), .A2(n9823), .A3(n9822), .A4(n9821), .ZN(
        P2_U3195) );
  AOI22_X1 U10946 ( .A1(n9825), .A2(n9875), .B1(n9874), .B2(
        P2_ADDR_REG_14__SCAN_IN), .ZN(n9840) );
  OAI21_X1 U10947 ( .B1(n9828), .B2(n9827), .A(n9826), .ZN(n9833) );
  OAI21_X1 U10948 ( .B1(n9831), .B2(n9830), .A(n9829), .ZN(n9832) );
  AOI22_X1 U10949 ( .A1(n9833), .A2(n9884), .B1(n9883), .B2(n9832), .ZN(n9839)
         );
  NAND2_X1 U10950 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3151), .ZN(n9838) );
  AOI21_X1 U10951 ( .B1(n4349), .B2(n9835), .A(n9834), .ZN(n9836) );
  OR2_X1 U10952 ( .A1(n9836), .A2(n9890), .ZN(n9837) );
  NAND4_X1 U10953 ( .A1(n9840), .A2(n9839), .A3(n9838), .A4(n9837), .ZN(
        P2_U3196) );
  AOI22_X1 U10954 ( .A1(n9841), .A2(n9875), .B1(n9874), .B2(
        P2_ADDR_REG_15__SCAN_IN), .ZN(n9856) );
  OAI21_X1 U10955 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n9843), .A(n9842), .ZN(
        n9848) );
  OAI21_X1 U10956 ( .B1(n9846), .B2(n9845), .A(n9844), .ZN(n9847) );
  AOI22_X1 U10957 ( .A1(n9848), .A2(n9884), .B1(n9883), .B2(n9847), .ZN(n9855)
         );
  AOI21_X1 U10958 ( .B1(n9851), .B2(n9850), .A(n9849), .ZN(n9852) );
  OR2_X1 U10959 ( .A1(n9890), .A2(n9852), .ZN(n9853) );
  NAND4_X1 U10960 ( .A1(n9856), .A2(n9855), .A3(n9854), .A4(n9853), .ZN(
        P2_U3197) );
  AOI22_X1 U10961 ( .A1(n9857), .A2(n9875), .B1(n9874), .B2(
        P2_ADDR_REG_16__SCAN_IN), .ZN(n9873) );
  OAI21_X1 U10962 ( .B1(n9860), .B2(n9859), .A(n9858), .ZN(n9865) );
  OAI21_X1 U10963 ( .B1(n9863), .B2(n9862), .A(n9861), .ZN(n9864) );
  AOI22_X1 U10964 ( .A1(n9865), .A2(n9884), .B1(n9883), .B2(n9864), .ZN(n9872)
         );
  AOI21_X1 U10965 ( .B1(n9868), .B2(n9867), .A(n9866), .ZN(n9869) );
  OR2_X1 U10966 ( .A1(n9869), .A2(n9890), .ZN(n9870) );
  NAND4_X1 U10967 ( .A1(n9873), .A2(n9872), .A3(n9871), .A4(n9870), .ZN(
        P2_U3198) );
  AOI22_X1 U10968 ( .A1(n9876), .A2(n9875), .B1(n9874), .B2(
        P2_ADDR_REG_17__SCAN_IN), .ZN(n9894) );
  OAI21_X1 U10969 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n9878), .A(n9877), .ZN(
        n9885) );
  OAI21_X1 U10970 ( .B1(n9881), .B2(n9880), .A(n9879), .ZN(n9882) );
  AOI22_X1 U10971 ( .A1(n9885), .A2(n9884), .B1(n9883), .B2(n9882), .ZN(n9893)
         );
  NAND2_X1 U10972 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3151), .ZN(n9892) );
  AOI21_X1 U10973 ( .B1(n9888), .B2(n9887), .A(n9886), .ZN(n9889) );
  OR2_X1 U10974 ( .A1(n9890), .A2(n9889), .ZN(n9891) );
  NAND4_X1 U10975 ( .A1(n9894), .A2(n9893), .A3(n9892), .A4(n9891), .ZN(
        P2_U3199) );
  INV_X1 U10976 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9906) );
  INV_X1 U10977 ( .A(n9895), .ZN(n9898) );
  OAI22_X1 U10978 ( .A1(n9898), .A2(n9897), .B1(n4886), .B2(n9896), .ZN(n9901)
         );
  INV_X1 U10979 ( .A(n9899), .ZN(n9900) );
  AOI211_X1 U10980 ( .C1(n9903), .C2(n9902), .A(n9901), .B(n9900), .ZN(n9905)
         );
  AOI22_X1 U10981 ( .A1(n9907), .A2(n9906), .B1(n9905), .B2(n9904), .ZN(
        P2_U3231) );
  AOI22_X1 U10982 ( .A1(n9969), .A2(n4850), .B1(n9908), .B2(n9967), .ZN(
        P2_U3393) );
  INV_X1 U10983 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9910) );
  AOI22_X1 U10984 ( .A1(n9969), .A2(n9910), .B1(n9909), .B2(n9967), .ZN(
        P2_U3396) );
  INV_X1 U10985 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9915) );
  OAI21_X1 U10986 ( .B1(n9912), .B2(n9948), .A(n9911), .ZN(n9913) );
  AOI21_X1 U10987 ( .B1(n9962), .B2(n9914), .A(n9913), .ZN(n9971) );
  AOI22_X1 U10988 ( .A1(n9969), .A2(n9915), .B1(n9971), .B2(n9967), .ZN(
        P2_U3399) );
  INV_X1 U10989 ( .A(n9916), .ZN(n9920) );
  OAI21_X1 U10990 ( .B1(n9918), .B2(n9948), .A(n9917), .ZN(n9919) );
  AOI21_X1 U10991 ( .B1(n9920), .B2(n9962), .A(n9919), .ZN(n9972) );
  AOI22_X1 U10992 ( .A1(n9969), .A2(n4909), .B1(n9972), .B2(n9967), .ZN(
        P2_U3402) );
  INV_X1 U10993 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9925) );
  NOR2_X1 U10994 ( .A1(n9921), .A2(n9948), .ZN(n9923) );
  AOI211_X1 U10995 ( .C1(n9962), .C2(n9924), .A(n9923), .B(n9922), .ZN(n9973)
         );
  AOI22_X1 U10996 ( .A1(n9969), .A2(n9925), .B1(n9973), .B2(n9967), .ZN(
        P2_U3405) );
  INV_X1 U10997 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9931) );
  INV_X1 U10998 ( .A(n9926), .ZN(n9930) );
  INV_X1 U10999 ( .A(n9962), .ZN(n9955) );
  OAI22_X1 U11000 ( .A1(n9928), .A2(n9955), .B1(n9927), .B2(n9948), .ZN(n9929)
         );
  NOR2_X1 U11001 ( .A1(n9930), .A2(n9929), .ZN(n9975) );
  AOI22_X1 U11002 ( .A1(n9969), .A2(n9931), .B1(n9975), .B2(n9967), .ZN(
        P2_U3408) );
  INV_X1 U11003 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9936) );
  OAI22_X1 U11004 ( .A1(n9933), .A2(n5501), .B1(n9932), .B2(n9948), .ZN(n9934)
         );
  NOR2_X1 U11005 ( .A1(n9935), .A2(n9934), .ZN(n9976) );
  AOI22_X1 U11006 ( .A1(n9969), .A2(n9936), .B1(n9976), .B2(n9967), .ZN(
        P2_U3411) );
  INV_X1 U11007 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9941) );
  OAI22_X1 U11008 ( .A1(n9938), .A2(n9955), .B1(n9937), .B2(n9948), .ZN(n9939)
         );
  NOR2_X1 U11009 ( .A1(n9940), .A2(n9939), .ZN(n9977) );
  AOI22_X1 U11010 ( .A1(n9969), .A2(n9941), .B1(n9977), .B2(n9967), .ZN(
        P2_U3414) );
  INV_X1 U11011 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9946) );
  NOR2_X1 U11012 ( .A1(n9942), .A2(n9948), .ZN(n9944) );
  AOI211_X1 U11013 ( .C1(n9945), .C2(n9953), .A(n9944), .B(n9943), .ZN(n9978)
         );
  AOI22_X1 U11014 ( .A1(n9969), .A2(n9946), .B1(n9978), .B2(n9967), .ZN(
        P2_U3417) );
  INV_X1 U11015 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9954) );
  INV_X1 U11016 ( .A(n9947), .ZN(n9949) );
  NOR2_X1 U11017 ( .A1(n9949), .A2(n9948), .ZN(n9951) );
  AOI211_X1 U11018 ( .C1(n9953), .C2(n9952), .A(n9951), .B(n9950), .ZN(n9979)
         );
  AOI22_X1 U11019 ( .A1(n9969), .A2(n9954), .B1(n9979), .B2(n9967), .ZN(
        P2_U3420) );
  NOR2_X1 U11020 ( .A1(n9956), .A2(n9955), .ZN(n9958) );
  AOI211_X1 U11021 ( .C1(n9966), .C2(n9959), .A(n9958), .B(n9957), .ZN(n9980)
         );
  AOI22_X1 U11022 ( .A1(n9969), .A2(n9960), .B1(n9980), .B2(n9967), .ZN(
        P2_U3423) );
  INV_X1 U11023 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9968) );
  AND3_X1 U11024 ( .A1(n7328), .A2(n9962), .A3(n9961), .ZN(n9964) );
  AOI211_X1 U11025 ( .C1(n9966), .C2(n9965), .A(n9964), .B(n9963), .ZN(n9981)
         );
  AOI22_X1 U11026 ( .A1(n9969), .A2(n9968), .B1(n9981), .B2(n9967), .ZN(
        P2_U3426) );
  INV_X1 U11027 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9970) );
  AOI22_X1 U11028 ( .A1(n9982), .A2(n9971), .B1(n9970), .B2(n6211), .ZN(
        P2_U3462) );
  AOI22_X1 U11029 ( .A1(n9982), .A2(n9972), .B1(n6479), .B2(n6211), .ZN(
        P2_U3463) );
  AOI22_X1 U11030 ( .A1(n9982), .A2(n9973), .B1(n4932), .B2(n6211), .ZN(
        P2_U3464) );
  AOI22_X1 U11031 ( .A1(n9982), .A2(n9975), .B1(n9974), .B2(n6211), .ZN(
        P2_U3465) );
  AOI22_X1 U11032 ( .A1(n9982), .A2(n9976), .B1(n7259), .B2(n6211), .ZN(
        P2_U3466) );
  AOI22_X1 U11033 ( .A1(n9982), .A2(n9977), .B1(n4990), .B2(n6211), .ZN(
        P2_U3467) );
  AOI22_X1 U11034 ( .A1(n9982), .A2(n9978), .B1(n7260), .B2(n6211), .ZN(
        P2_U3468) );
  AOI22_X1 U11035 ( .A1(n9982), .A2(n9979), .B1(n5038), .B2(n6211), .ZN(
        P2_U3469) );
  AOI22_X1 U11036 ( .A1(n9982), .A2(n9980), .B1(n5064), .B2(n6211), .ZN(
        P2_U3470) );
  AOI22_X1 U11037 ( .A1(n9982), .A2(n9981), .B1(n5077), .B2(n6211), .ZN(
        P2_U3471) );
  OAI222_X1 U11038 ( .A1(n9987), .A2(n9986), .B1(n9987), .B2(n9985), .C1(n9984), .C2(n9983), .ZN(ADD_1068_U5) );
  XOR2_X1 U11039 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  INV_X1 U11040 ( .A(n9990), .ZN(n9989) );
  OAI222_X1 U11041 ( .A1(n9992), .A2(n9991), .B1(n9992), .B2(n9990), .C1(n9989), .C2(n9988), .ZN(ADD_1068_U55) );
  OAI21_X1 U11042 ( .B1(n9995), .B2(n9994), .A(n9993), .ZN(ADD_1068_U56) );
  OAI21_X1 U11043 ( .B1(n9998), .B2(n9997), .A(n9996), .ZN(ADD_1068_U57) );
  OAI21_X1 U11044 ( .B1(n10001), .B2(n10000), .A(n9999), .ZN(ADD_1068_U58) );
  OAI21_X1 U11045 ( .B1(n10004), .B2(n10003), .A(n10002), .ZN(ADD_1068_U59) );
  OAI21_X1 U11046 ( .B1(n10007), .B2(n10006), .A(n10005), .ZN(ADD_1068_U60) );
  OAI21_X1 U11047 ( .B1(n10010), .B2(n10009), .A(n10008), .ZN(ADD_1068_U61) );
  OAI21_X1 U11048 ( .B1(n10013), .B2(n10012), .A(n10011), .ZN(ADD_1068_U62) );
  OAI21_X1 U11049 ( .B1(n10016), .B2(n10015), .A(n10014), .ZN(ADD_1068_U63) );
  OAI21_X1 U11050 ( .B1(n10019), .B2(n10018), .A(n10017), .ZN(ADD_1068_U50) );
  OAI21_X1 U11051 ( .B1(n10022), .B2(n10021), .A(n10020), .ZN(ADD_1068_U51) );
  OAI21_X1 U11052 ( .B1(n10025), .B2(n10024), .A(n10023), .ZN(ADD_1068_U47) );
  OAI21_X1 U11053 ( .B1(n10028), .B2(n10027), .A(n10026), .ZN(ADD_1068_U49) );
  OAI21_X1 U11054 ( .B1(n10031), .B2(n10030), .A(n10029), .ZN(ADD_1068_U48) );
  AOI21_X1 U11055 ( .B1(n10034), .B2(n10033), .A(n10032), .ZN(ADD_1068_U54) );
  AOI21_X1 U11056 ( .B1(n10037), .B2(n10036), .A(n10035), .ZN(ADD_1068_U53) );
  OAI21_X1 U11057 ( .B1(n10040), .B2(n10039), .A(n10038), .ZN(ADD_1068_U52) );
  CLKBUF_X2 U4783 ( .A(n5597), .Z(n5648) );
  CLKBUF_X1 U4858 ( .A(n6145), .Z(n4359) );
  CLKBUF_X1 U4948 ( .A(n5640), .Z(n5734) );
  CLKBUF_X1 U5717 ( .A(n9562), .Z(n4384) );
  CLKBUF_X2 U6026 ( .A(n8552), .Z(n4265) );
  CLKBUF_X1 U6053 ( .A(n7070), .Z(n4263) );
endmodule

