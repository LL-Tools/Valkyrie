

module b20_C_gen_AntiSAT_k_128_8 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, 
        ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, 
        ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, 
        ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, 
        ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, 
        P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, 
        P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, 
        P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, 
        P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, 
        P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, 
        P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, 
        P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, 
        P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, 
        P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, 
        P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, 
        P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, 
        P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, 
        P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, 
        P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, 
        P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, 
        P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, 
        P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, 
        P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, 
        P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, 
        P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, 
        P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, 
        P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, 
        P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, 
        P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, 
        P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, 
        P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, 
        P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, 
        P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, 
        P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, 
        P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, 
        P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10152;

  MUX2_X1 U4854 ( .A(n8798), .B(n8749), .S(n8755), .Z(n8750) );
  MUX2_X1 U4855 ( .A(n8799), .B(n8798), .S(n10088), .Z(n8800) );
  INV_X1 U4856 ( .A(n7033), .ZN(n4848) );
  INV_X1 U4857 ( .A(n5096), .ZN(n5471) );
  NAND2_X1 U4858 ( .A1(n6400), .A2(n6399), .ZN(n6423) );
  INV_X1 U4859 ( .A(n5683), .ZN(n5897) );
  INV_X2 U4860 ( .A(n5491), .ZN(n5356) );
  INV_X1 U4861 ( .A(n5216), .ZN(n5081) );
  INV_X1 U4863 ( .A(n10152), .ZN(n4349) );
  NOR2_X1 U4864 ( .A1(n4472), .A2(n4471), .ZN(n4469) );
  INV_X1 U4865 ( .A(n6686), .ZN(n5903) );
  OR2_X1 U4866 ( .A1(n6384), .A2(n6383), .ZN(n6385) );
  INV_X1 U4867 ( .A(n5048), .ZN(n5057) );
  INV_X1 U4868 ( .A(n5514), .ZN(n5405) );
  XNOR2_X1 U4869 ( .A(n8210), .B(n8589), .ZN(n8580) );
  OR2_X1 U4870 ( .A1(n5392), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5403) );
  INV_X1 U4871 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5210) );
  OAI211_X2 U4872 ( .C1(n9261), .C2(n6021), .A(n7917), .B(n6647), .ZN(n6507)
         );
  INV_X1 U4873 ( .A(n6941), .ZN(n7099) );
  CLKBUF_X2 U4874 ( .A(n5509), .Z(n8529) );
  NAND2_X1 U4875 ( .A1(n6321), .A2(n6180), .ZN(n6369) );
  NOR2_X1 U4877 ( .A1(n9393), .A2(n9392), .ZN(n9396) );
  AND2_X1 U4878 ( .A1(n6168), .A2(n5495), .ZN(n8563) );
  INV_X1 U4879 ( .A(n7614), .ZN(n8369) );
  INV_X1 U4880 ( .A(n8786), .ZN(n8755) );
  INV_X1 U4881 ( .A(n6096), .ZN(n9381) );
  NOR2_X2 U4882 ( .A1(n9490), .A2(n9483), .ZN(n4572) );
  NAND2_X2 U4883 ( .A1(n7756), .A2(n7757), .ZN(n7755) );
  OAI21_X2 U4884 ( .B1(n6956), .B2(n6962), .A(n6997), .ZN(n6963) );
  INV_X2 U4885 ( .A(n4928), .ZN(n6663) );
  XNOR2_X2 U4886 ( .A(n6878), .B(n5523), .ZN(n7044) );
  AOI21_X2 U4887 ( .B1(n4848), .B2(n4843), .A(n4840), .ZN(n7756) );
  OAI21_X2 U4888 ( .B1(n8301), .B2(n8169), .A(n4816), .ZN(n8308) );
  NAND2_X2 U4889 ( .A1(n5092), .A2(n5109), .ZN(n10022) );
  OAI21_X2 U4890 ( .B1(n5091), .B2(n5090), .A(n5089), .ZN(n5092) );
  OR4_X2 U4891 ( .A1(n6639), .A2(n6615), .A3(n8974), .A4(n6614), .ZN(n6636) );
  XNOR2_X2 U4892 ( .A(n5021), .B(n5044), .ZN(n6968) );
  AOI21_X1 U4893 ( .B1(n6059), .B2(n6058), .A(n6057), .ZN(n9400) );
  AOI21_X1 U4894 ( .B1(P2_REG1_REG_16__SCAN_IN), .B2(n8481), .A(n8471), .ZN(
        n8492) );
  INV_X1 U4895 ( .A(n9662), .ZN(n9570) );
  OR2_X1 U4896 ( .A1(n7861), .A2(n4791), .ZN(n4787) );
  OAI21_X1 U4897 ( .B1(n7735), .B2(n5530), .A(n6233), .ZN(n7781) );
  INV_X4 U4898 ( .A(n7358), .ZN(n8173) );
  INV_X4 U4899 ( .A(n6434), .ZN(n6601) );
  INV_X1 U4900 ( .A(n5099), .ZN(n10062) );
  INV_X1 U4901 ( .A(n7924), .ZN(n7699) );
  INV_X1 U4902 ( .A(n8368), .ZN(n7642) );
  INV_X1 U4903 ( .A(n8896), .ZN(n9956) );
  INV_X1 U4904 ( .A(n5101), .ZN(n5100) );
  NAND4_X1 U4905 ( .A1(n5071), .A2(n5070), .A3(n5069), .A4(n5068), .ZN(n6878)
         );
  INV_X2 U4906 ( .A(n6835), .ZN(n6060) );
  NAND4_X1 U4907 ( .A1(n5680), .A2(n5679), .A3(n5678), .A4(n5677), .ZN(n9284)
         );
  CLKBUF_X3 U4908 ( .A(n5081), .Z(n6161) );
  NAND2_X2 U4909 ( .A1(n5509), .A2(n6968), .ZN(n5088) );
  INV_X8 U4910 ( .A(n6663), .ZN(n4350) );
  INV_X2 U4911 ( .A(n5111), .ZN(n4786) );
  OR2_X1 U4912 ( .A1(n9396), .A2(n9395), .ZN(n9607) );
  OR2_X1 U4913 ( .A1(n8579), .A2(n8580), .ZN(n4593) );
  AOI21_X1 U4914 ( .B1(n9412), .B2(n9411), .A(n5995), .ZN(n6006) );
  NAND2_X1 U4915 ( .A1(n8184), .A2(n8183), .ZN(n8250) );
  OAI21_X1 U4916 ( .B1(n8946), .B2(n4831), .A(n4828), .ZN(n8989) );
  NOR2_X1 U4917 ( .A1(n4462), .A2(n4461), .ZN(n4468) );
  INV_X1 U4918 ( .A(n4668), .ZN(n9427) );
  NAND2_X1 U4919 ( .A1(n6552), .A2(n6553), .ZN(n8964) );
  NAND2_X1 U4920 ( .A1(n5489), .A2(n5488), .ZN(n8558) );
  NAND2_X1 U4921 ( .A1(n4483), .A2(n4482), .ZN(n6552) );
  OR2_X1 U4922 ( .A1(n9431), .A2(n6643), .ZN(n4908) );
  NAND2_X1 U4923 ( .A1(n5446), .A2(n5445), .ZN(n8210) );
  XNOR2_X1 U4924 ( .A(n6154), .B(n6153), .ZN(n6156) );
  OR2_X1 U4925 ( .A1(n8234), .A2(n8230), .ZN(n8168) );
  XNOR2_X1 U4926 ( .A(n8492), .B(n8505), .ZN(n8472) );
  NAND2_X1 U4927 ( .A1(n5415), .A2(n5414), .ZN(n8818) );
  NAND2_X1 U4928 ( .A1(n5945), .A2(n5944), .ZN(n9483) );
  INV_X1 U4929 ( .A(n8604), .ZN(n8578) );
  NAND2_X1 U4930 ( .A1(n5439), .A2(n5438), .ZN(n8604) );
  NAND2_X1 U4931 ( .A1(n5535), .A2(n6251), .ZN(n8005) );
  NAND2_X1 U4932 ( .A1(n5423), .A2(n5422), .ZN(n8628) );
  NAND2_X1 U4933 ( .A1(n5915), .A2(n5914), .ZN(n9647) );
  NAND2_X1 U4934 ( .A1(n4787), .A2(n4388), .ZN(n8291) );
  NAND2_X1 U4935 ( .A1(n5893), .A2(n5892), .ZN(n9657) );
  OR2_X1 U4936 ( .A1(n7706), .A2(n4634), .ZN(n4631) );
  NAND2_X1 U4937 ( .A1(n7559), .A2(n9081), .ZN(n9908) );
  NAND2_X1 U4938 ( .A1(n5041), .A2(n5040), .ZN(n5418) );
  OR2_X1 U4939 ( .A1(n7558), .A2(n9032), .ZN(n7559) );
  INV_X1 U4940 ( .A(n5416), .ZN(n5041) );
  NAND2_X1 U4941 ( .A1(n4695), .A2(n4566), .ZN(n7384) );
  AND2_X1 U4942 ( .A1(n9941), .A2(n4417), .ZN(n9917) );
  NAND2_X1 U4943 ( .A1(n5649), .A2(n5648), .ZN(n9672) );
  AND2_X1 U4944 ( .A1(n4805), .A2(n4802), .ZN(n7637) );
  NAND2_X1 U4945 ( .A1(n7473), .A2(n5757), .ZN(n9924) );
  NAND2_X1 U4946 ( .A1(n5848), .A2(n5847), .ZN(n9679) );
  OAI21_X1 U4947 ( .B1(n6829), .B2(n6823), .A(n6822), .ZN(n6821) );
  NAND2_X1 U4948 ( .A1(n4744), .A2(n4380), .ZN(n4747) );
  OAI21_X1 U4949 ( .B1(n9047), .B2(n9019), .A(n9217), .ZN(n7105) );
  OR2_X1 U4951 ( .A1(n6411), .A2(n6601), .ZN(n4916) );
  AND2_X1 U4952 ( .A1(n4624), .A2(n7403), .ZN(n7009) );
  INV_X2 U4953 ( .A(n6906), .ZN(n7358) );
  AND2_X1 U4954 ( .A1(n7067), .A2(n9970), .ZN(n6896) );
  NOR2_X1 U4955 ( .A1(n6866), .A2(n6648), .ZN(P2_U3893) );
  NOR2_X1 U4956 ( .A1(n7006), .A2(n7005), .ZN(n7430) );
  NAND4_X2 U4957 ( .A1(n5108), .A2(n5107), .A3(n5106), .A4(n5105), .ZN(n8370)
         );
  AND2_X1 U4958 ( .A1(n5561), .A2(n5560), .ZN(n5563) );
  NAND2_X1 U4959 ( .A1(n5674), .A2(n4644), .ZN(n7089) );
  OAI211_X1 U4960 ( .C1(n6686), .C2(n6756), .A(n5696), .B(n5695), .ZN(n8896)
         );
  XNOR2_X1 U4961 ( .A(n5552), .B(n5556), .ZN(n8129) );
  NAND4_X1 U4962 ( .A1(n5087), .A2(n5086), .A3(n5085), .A4(n5084), .ZN(n5101)
         );
  NAND3_X1 U4963 ( .A1(n5654), .A2(n4496), .A3(n5655), .ZN(n6417) );
  NAND2_X1 U4964 ( .A1(n5550), .A2(n5551), .ZN(n8202) );
  INV_X1 U4965 ( .A(n5673), .ZN(n5904) );
  CLKBUF_X1 U4966 ( .A(n5675), .Z(n6686) );
  AND2_X2 U4967 ( .A1(n5057), .A2(n5049), .ZN(n5491) );
  AND2_X1 U4968 ( .A1(n5048), .A2(n5056), .ZN(n5082) );
  XNOR2_X1 U4969 ( .A(n6020), .B(n6019), .ZN(n9204) );
  AND2_X2 U4970 ( .A1(n5624), .A2(n5623), .ZN(n5685) );
  NAND2_X1 U4971 ( .A1(n5048), .A2(n5049), .ZN(n5216) );
  AND2_X2 U4972 ( .A1(n5501), .A2(n5502), .ZN(n5555) );
  AND2_X1 U4973 ( .A1(n5498), .A2(n5497), .ZN(n5501) );
  CLKBUF_X1 U4974 ( .A(n6048), .Z(n4351) );
  OR2_X1 U4975 ( .A1(n5020), .A2(n5210), .ZN(n5021) );
  AND2_X1 U4976 ( .A1(n8873), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5047) );
  OAI21_X1 U4977 ( .B1(n5622), .B2(n4913), .A(n9724), .ZN(n8130) );
  NAND2_X2 U4978 ( .A1(n6669), .A2(P1_U3086), .ZN(n9729) );
  NOR2_X1 U4979 ( .A1(n5619), .A2(n5618), .ZN(n5622) );
  XNOR2_X1 U4980 ( .A(n5619), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5626) );
  NOR2_X1 U4981 ( .A1(n5016), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n4898) );
  XNOR2_X1 U4982 ( .A(n4667), .B(n5636), .ZN(n8108) );
  AND2_X1 U4983 ( .A1(n4892), .A2(n4605), .ZN(n4604) );
  OAI211_X1 U4984 ( .C1(n5074), .C2(n4537), .A(n5075), .B(n4536), .ZN(n6956)
         );
  AND2_X1 U4985 ( .A1(n5001), .A2(n5002), .ZN(n4605) );
  AND3_X1 U4986 ( .A1(n5003), .A2(n5305), .A3(n5348), .ZN(n5007) );
  AND4_X1 U4987 ( .A1(n5608), .A2(n5607), .A3(n5606), .A4(n5605), .ZN(n5609)
         );
  INV_X4 U4988 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U4989 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5025) );
  INV_X4 U4990 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U4991 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9386) );
  INV_X1 U4992 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4717) );
  INV_X1 U4993 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5142) );
  INV_X1 U4994 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5348) );
  NOR2_X1 U4995 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n5611) );
  INV_X1 U4996 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6010) );
  INV_X1 U4997 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6067) );
  INV_X1 U4998 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5002) );
  INV_X1 U4999 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5305) );
  INV_X1 U5000 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6016) );
  NAND2_X2 U5001 ( .A1(n8076), .A2(n8075), .ZN(n8145) );
  AOI22_X2 U5002 ( .A1(n9511), .A2(n5932), .B1(n9533), .B2(n9513), .ZN(n9489)
         );
  NOR2_X1 U5003 ( .A1(n6320), .A2(n4909), .ZN(n6330) );
  NOR2_X1 U5004 ( .A1(n5258), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5308) );
  OR2_X1 U5005 ( .A1(n9626), .A2(n6041), .ZN(n9172) );
  NAND2_X1 U5006 ( .A1(n9555), .A2(n9102), .ZN(n4662) );
  NOR2_X1 U5007 ( .A1(n9088), .A2(n4700), .ZN(n4699) );
  INV_X1 U5008 ( .A(n9230), .ZN(n4700) );
  OAI21_X2 U5009 ( .B1(n5209), .B2(n4768), .A(n4765), .ZN(n5257) );
  AOI21_X1 U5010 ( .B1(n4769), .B2(n4767), .A(n4766), .ZN(n4765) );
  INV_X1 U5011 ( .A(n4769), .ZN(n4768) );
  INV_X1 U5012 ( .A(n4961), .ZN(n4766) );
  NAND2_X1 U5013 ( .A1(n6647), .A2(n6396), .ZN(n6551) );
  NOR2_X1 U5014 ( .A1(n9095), .A2(n9094), .ZN(n4526) );
  NAND2_X1 U5015 ( .A1(n9120), .A2(n4516), .ZN(n4514) );
  NAND2_X1 U5016 ( .A1(n4504), .A2(n4514), .ZN(n4503) );
  INV_X1 U5017 ( .A(n9121), .ZN(n4504) );
  MUX2_X1 U5018 ( .A(n9176), .B(n9182), .S(n9155), .Z(n9121) );
  AOI21_X1 U5019 ( .B1(n4421), .B2(n4727), .A(n4723), .ZN(n4722) );
  INV_X1 U5020 ( .A(n5482), .ZN(n4723) );
  INV_X1 U5021 ( .A(n8910), .ZN(n4484) );
  OR2_X1 U5022 ( .A1(n9054), .A2(n9052), .ZN(n6033) );
  INV_X1 U5023 ( .A(n7862), .ZN(n4792) );
  OAI21_X1 U5024 ( .B1(n6326), .B2(n6325), .A(n4390), .ZN(n6327) );
  NOR2_X1 U5025 ( .A1(n6323), .A2(n6322), .ZN(n6324) );
  XOR2_X1 U5026 ( .A(n5047), .B(P2_IR_REG_29__SCAN_IN), .Z(n5049) );
  NAND2_X1 U5027 ( .A1(n7456), .A2(n7455), .ZN(n4640) );
  AND2_X1 U5028 ( .A1(n4898), .A2(n5211), .ZN(n5020) );
  AND3_X1 U5029 ( .A1(n4548), .A2(n4445), .A3(n4547), .ZN(n8402) );
  AND3_X1 U5030 ( .A1(n4534), .A2(n4532), .A3(n4444), .ZN(n8457) );
  NOR2_X1 U5031 ( .A1(n8818), .A2(n8253), .ZN(n6337) );
  NAND2_X1 U5032 ( .A1(n4860), .A2(n4862), .ZN(n4856) );
  NOR2_X1 U5033 ( .A1(n5345), .A2(n4859), .ZN(n4858) );
  INV_X1 U5034 ( .A(n4860), .ZN(n4859) );
  OR2_X1 U5035 ( .A1(n8860), .A2(n8712), .ZN(n6274) );
  OR2_X1 U5036 ( .A1(n8149), .A2(n8150), .ZN(n6258) );
  OR2_X1 U5037 ( .A1(n8041), .A2(n8097), .ZN(n6251) );
  NAND2_X1 U5038 ( .A1(n5142), .A2(n5127), .ZN(n4893) );
  NOR2_X1 U5039 ( .A1(n4385), .A2(n4833), .ZN(n4832) );
  INV_X1 U5040 ( .A(n6544), .ZN(n4833) );
  INV_X1 U5041 ( .A(n6552), .ZN(n6555) );
  INV_X1 U5042 ( .A(n6647), .ZN(n6607) );
  INV_X1 U5043 ( .A(n8130), .ZN(n5623) );
  NAND2_X1 U5044 ( .A1(n6045), .A2(n4704), .ZN(n4703) );
  INV_X1 U5045 ( .A(n9189), .ZN(n4704) );
  NOR2_X1 U5046 ( .A1(n6062), .A2(n9402), .ZN(n4581) );
  NAND2_X1 U5047 ( .A1(n9418), .A2(n6061), .ZN(n6062) );
  NAND2_X1 U5048 ( .A1(n9466), .A2(n6042), .ZN(n4702) );
  OAI21_X1 U5049 ( .B1(n6156), .B2(n7305), .A(n6155), .ZN(n6171) );
  OR2_X1 U5050 ( .A1(n6154), .A2(n6153), .ZN(n6155) );
  OAI21_X1 U5051 ( .B1(n4979), .B2(n4763), .A(n4759), .ZN(n5378) );
  AOI21_X1 U5052 ( .B1(n4982), .B2(n5364), .A(n4366), .ZN(n4763) );
  INV_X1 U5053 ( .A(n4760), .ZN(n4759) );
  OAI21_X1 U5054 ( .B1(n4764), .B2(n4762), .A(n4761), .ZN(n4760) );
  NAND2_X1 U5055 ( .A1(n4755), .A2(n4422), .ZN(n4754) );
  INV_X1 U5056 ( .A(n4757), .ZN(n4755) );
  AOI21_X1 U5057 ( .B1(n4971), .B2(n4970), .A(n4758), .ZN(n4757) );
  INV_X1 U5058 ( .A(n5320), .ZN(n4758) );
  XNOR2_X1 U5059 ( .A(n4972), .B(n7292), .ZN(n5320) );
  NOR2_X1 U5060 ( .A1(n4746), .A2(n4966), .ZN(n4745) );
  NAND2_X1 U5061 ( .A1(n4956), .A2(n4955), .ZN(n5209) );
  AOI21_X1 U5062 ( .B1(n4737), .B2(n4740), .A(n4736), .ZN(n4735) );
  NAND2_X1 U5063 ( .A1(n7536), .A2(n4808), .ZN(n4806) );
  NOR2_X1 U5064 ( .A1(n7456), .A2(n7455), .ZN(n7650) );
  XNOR2_X1 U5065 ( .A(n8402), .B(n8403), .ZN(n8390) );
  NAND2_X1 U5066 ( .A1(n4593), .A2(n4586), .ZN(n4585) );
  NOR2_X1 U5067 ( .A1(n4592), .A2(n4587), .ZN(n4586) );
  INV_X1 U5068 ( .A(n4590), .ZN(n4587) );
  NOR2_X1 U5069 ( .A1(n8028), .A2(n4603), .ZN(n4602) );
  INV_X1 U5070 ( .A(n6230), .ZN(n4603) );
  NAND2_X1 U5071 ( .A1(n7610), .A2(n5148), .ZN(n5150) );
  NAND2_X1 U5072 ( .A1(n4596), .A2(n7626), .ZN(n4595) );
  AND2_X1 U5073 ( .A1(n6213), .A2(n6199), .ZN(n4596) );
  INV_X1 U5074 ( .A(n8612), .ZN(n8588) );
  AND2_X1 U5075 ( .A1(n5508), .A2(n6187), .ZN(n8666) );
  NAND2_X1 U5076 ( .A1(n5323), .A2(n4423), .ZN(n4797) );
  NAND2_X1 U5077 ( .A1(n5323), .A2(n5322), .ZN(n5336) );
  AND2_X1 U5078 ( .A1(n6585), .A2(n4829), .ZN(n4828) );
  NAND2_X1 U5079 ( .A1(n8917), .A2(n4830), .ZN(n4829) );
  AND2_X1 U5080 ( .A1(n8990), .A2(n8987), .ZN(n6585) );
  INV_X1 U5081 ( .A(n6574), .ZN(n4830) );
  NAND2_X1 U5082 ( .A1(n5599), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5948) );
  INV_X1 U5083 ( .A(n5925), .ZN(n5599) );
  OR2_X1 U5084 ( .A1(n5973), .A2(n8919), .ZN(n5975) );
  NAND2_X1 U5085 ( .A1(n4466), .A2(n4465), .ZN(n8946) );
  OAI21_X1 U5086 ( .B1(n6555), .B2(n4461), .A(n4460), .ZN(n4466) );
  AOI21_X1 U5087 ( .B1(n8964), .B2(n4463), .A(n4459), .ZN(n4465) );
  AOI21_X1 U5088 ( .B1(n8885), .B2(n6553), .A(n4467), .ZN(n4460) );
  AOI21_X1 U5089 ( .B1(n6417), .B2(n6407), .A(n6416), .ZN(n6418) );
  NAND2_X1 U5090 ( .A1(n4675), .A2(n4356), .ZN(n4674) );
  INV_X1 U5091 ( .A(n4678), .ZN(n4675) );
  AOI21_X1 U5092 ( .B1(n4680), .B2(n4679), .A(n4392), .ZN(n4678) );
  NAND2_X1 U5093 ( .A1(n4680), .A2(n4356), .ZN(n4676) );
  INV_X1 U5094 ( .A(n9440), .ZN(n6043) );
  INV_X1 U5095 ( .A(n4647), .ZN(n9511) );
  OAI21_X1 U5096 ( .B1(n9565), .B2(n4651), .A(n4648), .ZN(n4647) );
  NAND2_X1 U5097 ( .A1(n4652), .A2(n5921), .ZN(n4651) );
  INV_X1 U5098 ( .A(n4649), .ZN(n4648) );
  NAND2_X1 U5099 ( .A1(n4407), .A2(n4662), .ZN(n4659) );
  NAND2_X1 U5100 ( .A1(n9583), .A2(n9584), .ZN(n4694) );
  AOI21_X1 U5101 ( .B1(n4697), .B2(n4699), .A(n6036), .ZN(n4696) );
  INV_X1 U5102 ( .A(n6035), .ZN(n4697) );
  NOR2_X1 U5103 ( .A1(n4698), .A2(n9915), .ZN(n4568) );
  INV_X1 U5104 ( .A(n4699), .ZN(n4698) );
  NAND2_X1 U5105 ( .A1(n6841), .A2(n5671), .ZN(n7082) );
  OR2_X1 U5106 ( .A1(n6417), .A2(n6835), .ZN(n5671) );
  NAND2_X1 U5107 ( .A1(n5675), .A2(n4364), .ZN(n4835) );
  INV_X1 U5109 ( .A(n8357), .ZN(n8577) );
  AND2_X1 U5110 ( .A1(n9233), .A2(n9229), .ZN(n4524) );
  NAND2_X1 U5111 ( .A1(n4528), .A2(n4527), .ZN(n9095) );
  NAND2_X1 U5112 ( .A1(n9087), .A2(n4516), .ZN(n4527) );
  NAND2_X1 U5113 ( .A1(n4513), .A2(n4511), .ZN(n4502) );
  INV_X1 U5114 ( .A(n4514), .ZN(n4512) );
  OAI21_X1 U5115 ( .B1(n4508), .B2(n9128), .A(n4505), .ZN(n9133) );
  INV_X1 U5116 ( .A(n4506), .ZN(n4505) );
  OAI21_X1 U5117 ( .B1(n4507), .B2(n9128), .A(n9127), .ZN(n4506) );
  AOI21_X1 U5118 ( .B1(n9393), .B2(n4729), .A(n4728), .ZN(n4730) );
  NAND2_X1 U5119 ( .A1(n9389), .A2(n9275), .ZN(n4729) );
  INV_X1 U5120 ( .A(n9144), .ZN(n4728) );
  AND2_X1 U5121 ( .A1(n6033), .A2(n6031), .ZN(n9218) );
  NAND2_X1 U5122 ( .A1(n5487), .A2(n5486), .ZN(n6154) );
  NAND2_X1 U5123 ( .A1(n4724), .A2(n4722), .ZN(n5487) );
  INV_X1 U5124 ( .A(n5429), .ZN(n4726) );
  NOR2_X1 U5125 ( .A1(n5186), .A2(n4742), .ZN(n4741) );
  INV_X1 U5126 ( .A(n4945), .ZN(n4742) );
  INV_X1 U5127 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4720) );
  NOR2_X1 U5128 ( .A1(n5012), .A2(n4800), .ZN(n5013) );
  INV_X1 U5129 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5012) );
  AND2_X1 U5130 ( .A1(n8741), .A2(n8549), .ZN(n6374) );
  NAND2_X1 U5131 ( .A1(n10027), .A2(n7017), .ZN(n4531) );
  NOR2_X1 U5132 ( .A1(n7004), .A2(n7441), .ZN(n7006) );
  NAND2_X1 U5133 ( .A1(n4620), .A2(n4622), .ZN(n4624) );
  NOR2_X1 U5134 ( .A1(n4623), .A2(n4400), .ZN(n4620) );
  INV_X1 U5135 ( .A(n7419), .ZN(n4626) );
  NAND3_X1 U5136 ( .A1(n4632), .A2(n4438), .A3(n4631), .ZN(n8396) );
  INV_X1 U5137 ( .A(n8399), .ZN(n4629) );
  NOR2_X1 U5138 ( .A1(n5542), .A2(n8604), .ZN(n4869) );
  INV_X1 U5139 ( .A(n6348), .ZN(n4884) );
  NAND2_X1 U5140 ( .A1(n5564), .A2(n6783), .ZN(n7369) );
  INV_X1 U5141 ( .A(n7846), .ZN(n6144) );
  NAND2_X1 U5142 ( .A1(n8812), .A2(n8588), .ZN(n4879) );
  NAND2_X1 U5143 ( .A1(n4878), .A2(n4372), .ZN(n4877) );
  OR2_X1 U5144 ( .A1(n8256), .A2(n8588), .ZN(n6305) );
  INV_X1 U5145 ( .A(n6299), .ZN(n4609) );
  OR2_X1 U5146 ( .A1(n8836), .A2(n8667), .ZN(n6290) );
  OR2_X1 U5147 ( .A1(n8773), .A2(n8246), .ZN(n6289) );
  OR2_X1 U5148 ( .A1(n8867), .A2(n8346), .ZN(n6266) );
  AND2_X1 U5149 ( .A1(n7975), .A2(n5238), .ZN(n4897) );
  INV_X1 U5150 ( .A(n5254), .ZN(n4896) );
  INV_X1 U5151 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5579) );
  AND2_X1 U5152 ( .A1(n5308), .A2(n5307), .ZN(n5323) );
  OAI21_X1 U5153 ( .B1(n7755), .B2(n4822), .A(n4821), .ZN(n6505) );
  AOI21_X1 U5154 ( .B1(n7849), .B2(n6496), .A(n4403), .ZN(n4821) );
  INV_X1 U5155 ( .A(n7849), .ZN(n4822) );
  INV_X1 U5156 ( .A(n6516), .ZN(n4471) );
  INV_X1 U5157 ( .A(n4826), .ZN(n4825) );
  OAI21_X1 U5158 ( .B1(n8927), .B2(n4827), .A(n8936), .ZN(n4826) );
  INV_X1 U5159 ( .A(n8935), .ZN(n4824) );
  INV_X1 U5160 ( .A(n6521), .ZN(n4827) );
  NAND2_X1 U5161 ( .A1(n4480), .A2(n6488), .ZN(n4841) );
  INV_X1 U5162 ( .A(n8945), .ZN(n4459) );
  INV_X1 U5163 ( .A(n7132), .ZN(n4846) );
  AND2_X1 U5164 ( .A1(n6516), .A2(n8996), .ZN(n4472) );
  OAI21_X1 U5165 ( .B1(n4674), .B2(n4671), .A(n4404), .ZN(n4670) );
  INV_X1 U5166 ( .A(n5981), .ZN(n4671) );
  INV_X1 U5167 ( .A(n4676), .ZN(n4673) );
  NOR2_X1 U5168 ( .A1(n9530), .A2(n4559), .ZN(n4558) );
  INV_X1 U5169 ( .A(n9248), .ZN(n4559) );
  OR2_X1 U5170 ( .A1(n9679), .A2(n9002), .ZN(n9229) );
  OR2_X1 U5171 ( .A1(n9914), .A2(n7852), .ZN(n9085) );
  OR2_X1 U5172 ( .A1(n7882), .A2(n5812), .ZN(n9081) );
  NOR2_X1 U5173 ( .A1(n7512), .A2(n7391), .ZN(n4571) );
  NAND2_X1 U5174 ( .A1(n9218), .A2(n7105), .ZN(n4695) );
  AND2_X1 U5175 ( .A1(n4419), .A2(n4915), .ZN(n4851) );
  NAND2_X1 U5176 ( .A1(n4751), .A2(n4749), .ZN(n5347) );
  NOR2_X1 U5177 ( .A1(n4753), .A2(n4750), .ZN(n4749) );
  INV_X1 U5178 ( .A(n4978), .ZN(n4750) );
  INV_X1 U5179 ( .A(n5741), .ZN(n4853) );
  OAI21_X1 U5180 ( .B1(n5257), .B2(SI_13_), .A(n5255), .ZN(n4963) );
  NAND2_X1 U5181 ( .A1(n4960), .A2(SI_12_), .ZN(n4961) );
  AND2_X1 U5182 ( .A1(n4410), .A2(n4958), .ZN(n4774) );
  INV_X1 U5183 ( .A(n4379), .ZN(n4775) );
  AOI21_X1 U5184 ( .B1(n4741), .B2(n4739), .A(n4738), .ZN(n4737) );
  INV_X1 U5185 ( .A(n4949), .ZN(n4738) );
  INV_X1 U5186 ( .A(n5173), .ZN(n4739) );
  INV_X1 U5187 ( .A(n4741), .ZN(n4740) );
  NAND2_X1 U5188 ( .A1(n4928), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4922) );
  AND2_X1 U5189 ( .A1(n4783), .A2(n8332), .ZN(n4782) );
  NAND2_X1 U5190 ( .A1(n8331), .A2(n4784), .ZN(n4783) );
  INV_X1 U5191 ( .A(n8186), .ZN(n4784) );
  INV_X1 U5192 ( .A(n8331), .ZN(n4785) );
  NAND2_X1 U5193 ( .A1(n4782), .A2(n4785), .ZN(n4779) );
  NOR2_X1 U5194 ( .A1(n8205), .A2(n4781), .ZN(n4780) );
  INV_X1 U5195 ( .A(n4782), .ZN(n4781) );
  NAND2_X1 U5196 ( .A1(n7952), .A2(n7960), .ZN(n4794) );
  NAND2_X1 U5197 ( .A1(n4793), .A2(n4792), .ZN(n7953) );
  INV_X1 U5198 ( .A(n7861), .ZN(n4793) );
  NAND2_X1 U5199 ( .A1(n7533), .A2(n8370), .ZN(n4808) );
  OR2_X1 U5200 ( .A1(n7362), .A2(n7363), .ZN(n4809) );
  NAND2_X1 U5201 ( .A1(n4807), .A2(n4809), .ZN(n7581) );
  INV_X1 U5202 ( .A(n4806), .ZN(n4807) );
  NAND2_X1 U5203 ( .A1(n4792), .A2(n8019), .ZN(n4791) );
  AOI21_X1 U5204 ( .B1(n4813), .B2(n4811), .A(n4425), .ZN(n4810) );
  INV_X1 U5205 ( .A(n4813), .ZN(n4812) );
  NAND2_X1 U5206 ( .A1(n6866), .A2(n6788), .ZN(n6390) );
  AND2_X1 U5207 ( .A1(n6334), .A2(n6333), .ZN(n6382) );
  NOR3_X1 U5208 ( .A1(n6382), .A2(n6374), .A3(n6903), .ZN(n6381) );
  NAND2_X1 U5209 ( .A1(n4588), .A2(n4393), .ZN(n6189) );
  OAI21_X1 U5210 ( .B1(n4585), .B2(n6323), .A(n4582), .ZN(n4588) );
  AND2_X1 U5211 ( .A1(n4589), .A2(n4583), .ZN(n4582) );
  OAI21_X1 U5212 ( .B1(n6956), .B2(n6955), .A(n7015), .ZN(n6958) );
  AND2_X1 U5213 ( .A1(n4546), .A2(n7415), .ZN(n7434) );
  NAND2_X1 U5214 ( .A1(n7492), .A2(n4545), .ZN(n4546) );
  NOR2_X1 U5215 ( .A1(n7020), .A2(n4355), .ZN(n4545) );
  AOI22_X1 U5216 ( .A1(n7442), .A2(n7443), .B1(n6986), .B2(n7020), .ZN(n7425)
         );
  OAI21_X1 U5217 ( .B1(n7019), .B2(n4355), .A(n4543), .ZN(n7415) );
  INV_X1 U5218 ( .A(n4544), .ZN(n4543) );
  OAI21_X1 U5219 ( .B1(n4355), .B2(n7488), .A(n7020), .ZN(n4544) );
  NOR2_X1 U5220 ( .A1(n7411), .A2(n7412), .ZN(n4623) );
  NAND2_X1 U5221 ( .A1(n4640), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4639) );
  OAI21_X1 U5222 ( .B1(n4712), .B2(P2_REG2_REG_9__SCAN_IN), .A(n4711), .ZN(
        n4542) );
  INV_X1 U5223 ( .A(n7668), .ZN(n4711) );
  AOI21_X1 U5224 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n7708), .A(n7705), .ZN(
        n7806) );
  OR2_X1 U5225 ( .A1(n7707), .A2(n4441), .ZN(n4547) );
  NAND2_X1 U5226 ( .A1(n7812), .A2(n4549), .ZN(n4548) );
  INV_X1 U5227 ( .A(n7814), .ZN(n4549) );
  OR2_X1 U5228 ( .A1(n7707), .A2(n7935), .ZN(n4551) );
  XNOR2_X1 U5229 ( .A(n8396), .B(n8389), .ZN(n8384) );
  OR2_X1 U5230 ( .A1(n8390), .A2(n4367), .ZN(n4534) );
  INV_X1 U5231 ( .A(n8406), .ZN(n4533) );
  NAND2_X1 U5232 ( .A1(n4535), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4714) );
  INV_X1 U5233 ( .A(n8390), .ZN(n4535) );
  NOR2_X1 U5234 ( .A1(n8428), .A2(n8431), .ZN(n8459) );
  INV_X1 U5235 ( .A(n5490), .ZN(n8547) );
  OAI21_X1 U5236 ( .B1(n4878), .B2(n4871), .A(n4868), .ZN(n8575) );
  NAND2_X1 U5237 ( .A1(n4873), .A2(n4872), .ZN(n4871) );
  AOI21_X1 U5238 ( .B1(n4873), .B2(n4870), .A(n4869), .ZN(n4868) );
  INV_X1 U5239 ( .A(n5440), .ZN(n4872) );
  OAI21_X1 U5240 ( .B1(n8592), .B2(n6310), .A(n6308), .ZN(n8579) );
  NAND2_X1 U5241 ( .A1(n4600), .A2(n4395), .ZN(n5536) );
  NAND2_X1 U5242 ( .A1(n5239), .A2(n4897), .ZN(n7974) );
  INV_X1 U5243 ( .A(n8361), .ZN(n8097) );
  INV_X1 U5244 ( .A(n4887), .ZN(n4886) );
  OAI21_X1 U5245 ( .B1(n4889), .B2(n4888), .A(n8030), .ZN(n4887) );
  NAND2_X1 U5246 ( .A1(n4406), .A2(n5208), .ZN(n4888) );
  INV_X1 U5247 ( .A(n7781), .ZN(n5531) );
  AND2_X1 U5248 ( .A1(n5533), .A2(n7931), .ZN(n7888) );
  AND4_X1 U5249 ( .A1(n5236), .A2(n5235), .A3(n5234), .A4(n5233), .ZN(n8052)
         );
  NAND2_X1 U5250 ( .A1(n4864), .A2(n5133), .ZN(n4866) );
  AND2_X1 U5251 ( .A1(n7691), .A2(n4597), .ZN(n4594) );
  AND2_X1 U5252 ( .A1(n6214), .A2(n6208), .ZN(n7691) );
  NAND2_X1 U5253 ( .A1(n5100), .A2(n5099), .ZN(n6199) );
  INV_X1 U5254 ( .A(n6197), .ZN(n5527) );
  NAND2_X1 U5255 ( .A1(n7046), .A2(n7375), .ZN(n7045) );
  NAND2_X1 U5256 ( .A1(n7376), .A2(n5544), .ZN(n7892) );
  NOR2_X1 U5257 ( .A1(n7899), .A2(n6144), .ZN(n6880) );
  OR2_X1 U5258 ( .A1(n8549), .A2(n8548), .ZN(n8744) );
  OR2_X1 U5259 ( .A1(n6310), .A2(n6311), .ZN(n8591) );
  NAND2_X1 U5260 ( .A1(n4874), .A2(n4879), .ZN(n4873) );
  INV_X1 U5261 ( .A(n4875), .ZN(n4874) );
  OR2_X1 U5262 ( .A1(n6337), .A2(n6336), .ZN(n8619) );
  OR2_X1 U5263 ( .A1(n8830), .A2(n5396), .ZN(n6292) );
  NAND2_X1 U5264 ( .A1(n8634), .A2(n8637), .ZN(n4611) );
  NAND2_X1 U5265 ( .A1(n5361), .A2(n4919), .ZN(n4891) );
  NAND2_X1 U5266 ( .A1(n6911), .A2(n6659), .ZN(n8669) );
  INV_X1 U5267 ( .A(n5543), .ZN(n8539) );
  AOI21_X1 U5268 ( .B1(n6340), .B2(n4861), .A(n4397), .ZN(n4860) );
  INV_X1 U5269 ( .A(n5318), .ZN(n4861) );
  OAI22_X1 U5270 ( .A1(n8724), .A2(n5300), .B1(n8217), .B2(n8355), .ZN(n8708)
         );
  INV_X1 U5271 ( .A(n8728), .ZN(n8711) );
  INV_X1 U5272 ( .A(n8666), .ZN(n8731) );
  NOR2_X1 U5273 ( .A1(n8077), .A2(n8144), .ZN(n4601) );
  OR2_X1 U5274 ( .A1(n6383), .A2(n6392), .ZN(n7899) );
  INV_X1 U5275 ( .A(n8793), .ZN(n8745) );
  INV_X1 U5276 ( .A(n6876), .ZN(n6885) );
  INV_X1 U5277 ( .A(n6390), .ZN(n6879) );
  NAND2_X1 U5278 ( .A1(n4455), .A2(n4454), .ZN(n5016) );
  NOR2_X1 U5279 ( .A1(n5014), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n4454) );
  INV_X1 U5280 ( .A(n5015), .ZN(n4455) );
  AND2_X1 U5281 ( .A1(n4619), .A2(n5044), .ZN(n4618) );
  INV_X1 U5282 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4619) );
  INV_X1 U5283 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5556) );
  INV_X1 U5284 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5502) );
  INV_X1 U5285 ( .A(n4799), .ZN(n4798) );
  OAI21_X1 U5286 ( .B1(n4423), .B2(n4800), .A(n5348), .ZN(n4799) );
  AND2_X1 U5287 ( .A1(n5275), .A2(n5290), .ZN(n8417) );
  CLKBUF_X1 U5288 ( .A(n5202), .Z(n5203) );
  AND2_X1 U5289 ( .A1(n4892), .A2(n5001), .ZN(n4606) );
  NOR2_X1 U5290 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5000) );
  INV_X1 U5291 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4537) );
  NAND2_X1 U5292 ( .A1(n6506), .A2(n6508), .ZN(n4838) );
  INV_X1 U5293 ( .A(n7986), .ZN(n6508) );
  OR2_X1 U5294 ( .A1(n6505), .A2(n6504), .ZN(n6506) );
  INV_X1 U5295 ( .A(n8885), .ZN(n4461) );
  AND2_X1 U5296 ( .A1(n6482), .A2(n6481), .ZN(n7798) );
  AOI21_X1 U5297 ( .B1(n4832), .B2(n4487), .A(n4382), .ZN(n4486) );
  INV_X1 U5298 ( .A(n8902), .ZN(n4487) );
  INV_X1 U5299 ( .A(n4832), .ZN(n4488) );
  AND2_X1 U5300 ( .A1(n4845), .A2(n6488), .ZN(n4843) );
  NAND2_X1 U5301 ( .A1(n4842), .A2(n4841), .ZN(n4840) );
  INV_X1 U5302 ( .A(n6487), .ZN(n4842) );
  OR2_X1 U5303 ( .A1(n5866), .A2(n5865), .ZN(n5878) );
  NAND2_X1 U5304 ( .A1(n5601), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5973) );
  NAND2_X1 U5305 ( .A1(n9940), .A2(n6604), .ZN(n6466) );
  AND2_X1 U5306 ( .A1(n4847), .A2(n4846), .ZN(n7830) );
  NAND2_X1 U5307 ( .A1(n4848), .A2(n4849), .ZN(n4847) );
  NAND2_X1 U5308 ( .A1(n5831), .A2(n5830), .ZN(n6499) );
  NAND2_X1 U5309 ( .A1(n6555), .A2(n6554), .ZN(n8965) );
  AND2_X1 U5310 ( .A1(n6612), .A2(n6611), .ZN(n6620) );
  NAND2_X1 U5311 ( .A1(n6014), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6065) );
  INV_X1 U5312 ( .A(n5685), .ZN(n6050) );
  NAND2_X1 U5313 ( .A1(n5685), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5653) );
  OR2_X1 U5314 ( .A1(n5701), .A2(n5651), .ZN(n5652) );
  NAND2_X1 U5315 ( .A1(n6094), .A2(n6097), .ZN(n6647) );
  NAND2_X1 U5316 ( .A1(n6685), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6811) );
  NAND2_X1 U5317 ( .A1(n4703), .A2(n9142), .ZN(n6118) );
  INV_X1 U5318 ( .A(n9157), .ZN(n9145) );
  NAND2_X1 U5319 ( .A1(n4581), .A2(n4580), .ZN(n9392) );
  AND2_X1 U5320 ( .A1(n9166), .A2(n9144), .ZN(n9157) );
  NAND2_X1 U5321 ( .A1(n9180), .A2(n9138), .ZN(n9411) );
  AND2_X1 U5322 ( .A1(n6043), .A2(n9172), .ZN(n4701) );
  NOR2_X1 U5323 ( .A1(n4378), .A2(n4682), .ZN(n4681) );
  INV_X1 U5324 ( .A(n5943), .ZN(n4682) );
  AND2_X1 U5325 ( .A1(n5955), .A2(n4369), .ZN(n4683) );
  AND2_X1 U5326 ( .A1(n9126), .A2(n9467), .ZN(n9481) );
  OR2_X1 U5327 ( .A1(n4656), .A2(n4381), .ZN(n4653) );
  AOI21_X1 U5328 ( .B1(n4657), .B2(n4659), .A(n4401), .ZN(n4656) );
  INV_X1 U5329 ( .A(n4660), .ZN(n4657) );
  OR2_X1 U5330 ( .A1(n4658), .A2(n4381), .ZN(n4654) );
  INV_X1 U5331 ( .A(n4659), .ZN(n4658) );
  AND2_X1 U5332 ( .A1(n4662), .A2(n5886), .ZN(n4660) );
  AND2_X1 U5333 ( .A1(n9242), .A2(n9248), .ZN(n9544) );
  NOR2_X1 U5334 ( .A1(n9564), .A2(n4565), .ZN(n4564) );
  INV_X1 U5335 ( .A(n9237), .ZN(n4565) );
  NAND2_X1 U5336 ( .A1(n4563), .A2(n4561), .ZN(n9556) );
  NOR2_X1 U5337 ( .A1(n4562), .A2(n6038), .ZN(n4561) );
  INV_X1 U5338 ( .A(n9558), .ZN(n4562) );
  AND2_X1 U5339 ( .A1(n9241), .A2(n9240), .ZN(n9558) );
  NAND2_X1 U5340 ( .A1(n4567), .A2(n4384), .ZN(n8012) );
  AND2_X1 U5341 ( .A1(n9233), .A2(n9097), .ZN(n9036) );
  OAI22_X1 U5342 ( .A1(n7909), .A2(n5859), .B1(n7989), .B2(n9002), .ZN(n8009)
         );
  AND2_X1 U5343 ( .A1(n7767), .A2(n4699), .ZN(n7911) );
  NAND2_X1 U5344 ( .A1(n9907), .A2(n6035), .ZN(n7767) );
  NAND2_X1 U5345 ( .A1(n9908), .A2(n4687), .ZN(n9907) );
  INV_X1 U5346 ( .A(n4689), .ZN(n4688) );
  OAI21_X1 U5347 ( .B1(n7560), .B2(n4693), .A(n4692), .ZN(n4689) );
  OR2_X1 U5348 ( .A1(n7882), .A2(n9910), .ZN(n4692) );
  NOR2_X1 U5349 ( .A1(n7560), .A2(n6034), .ZN(n4690) );
  AND2_X1 U5350 ( .A1(n9081), .A2(n9082), .ZN(n7560) );
  AOI22_X1 U5351 ( .A1(n9924), .A2(n5769), .B1(n9981), .B2(n7836), .ZN(n7519)
         );
  AND2_X1 U5352 ( .A1(n9944), .A2(n9981), .ZN(n9941) );
  NOR2_X2 U5353 ( .A1(n7479), .A2(n7598), .ZN(n9944) );
  NAND2_X1 U5354 ( .A1(n6894), .A2(n9019), .ZN(n6893) );
  INV_X1 U5355 ( .A(n7913), .ZN(n9932) );
  OR2_X1 U5356 ( .A1(n9260), .A2(n6397), .ZN(n7917) );
  OR2_X1 U5357 ( .A1(n6608), .A2(n4351), .ZN(n7913) );
  OR2_X1 U5358 ( .A1(n6688), .A2(n6621), .ZN(n9515) );
  NAND2_X1 U5359 ( .A1(n5984), .A2(n5983), .ZN(n9420) );
  OR2_X1 U5360 ( .A1(n7122), .A2(n5887), .ZN(n5893) );
  XNOR2_X1 U5361 ( .A(n6174), .B(n6173), .ZN(n9015) );
  OAI21_X1 U5362 ( .B1(n6171), .B2(n6170), .A(n6169), .ZN(n6174) );
  NAND2_X1 U5363 ( .A1(n4905), .A2(P1_IR_REG_30__SCAN_IN), .ZN(n5618) );
  XNOR2_X1 U5364 ( .A(n6171), .B(n6170), .ZN(n9010) );
  NAND2_X1 U5365 ( .A1(n4523), .A2(n4521), .ZN(n5619) );
  INV_X1 U5366 ( .A(n4522), .ZN(n4521) );
  NAND2_X1 U5367 ( .A1(n6069), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4523) );
  OAI21_X1 U5368 ( .B1(n4851), .B2(n5800), .A(n5617), .ZN(n4522) );
  NAND2_X1 U5369 ( .A1(n4721), .A2(n4421), .ZN(n5483) );
  OR2_X1 U5370 ( .A1(n5430), .A2(n4727), .ZN(n4721) );
  INV_X1 U5371 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5636) );
  OAI21_X1 U5372 ( .B1(n5347), .B2(n5346), .A(n4982), .ZN(n5366) );
  NAND2_X1 U5373 ( .A1(n5901), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5902) );
  NOR2_X1 U5374 ( .A1(n4754), .A2(n5333), .ZN(n4753) );
  NAND2_X1 U5375 ( .A1(n5303), .A2(n4362), .ZN(n4752) );
  NAND2_X1 U5376 ( .A1(n4756), .A2(n4970), .ZN(n5321) );
  NAND2_X1 U5377 ( .A1(n4747), .A2(n4965), .ZN(n5289) );
  OAI21_X1 U5378 ( .B1(n4960), .B2(SI_12_), .A(n4961), .ZN(n5240) );
  NOR2_X1 U5379 ( .A1(n4770), .A2(n5240), .ZN(n4769) );
  INV_X1 U5380 ( .A(n4772), .ZN(n4770) );
  AOI21_X1 U5381 ( .B1(n4775), .B2(n4774), .A(n4773), .ZN(n4772) );
  NOR2_X1 U5382 ( .A1(n5224), .A2(SI_11_), .ZN(n4773) );
  NAND2_X1 U5383 ( .A1(n5209), .A2(n4774), .ZN(n4771) );
  XNOR2_X1 U5384 ( .A(n5187), .B(n5186), .ZN(n6690) );
  NAND2_X1 U5385 ( .A1(n4743), .A2(n4945), .ZN(n5187) );
  NAND2_X1 U5386 ( .A1(n4491), .A2(n4489), .ZN(n4743) );
  INV_X1 U5387 ( .A(n4490), .ZN(n4489) );
  AOI21_X1 U5388 ( .B1(n5162), .B2(n4493), .A(n4371), .ZN(n4495) );
  NAND2_X1 U5389 ( .A1(n6918), .A2(n6917), .ZN(n6916) );
  INV_X1 U5390 ( .A(n8367), .ZN(n7864) );
  NOR2_X1 U5391 ( .A1(n4358), .A2(n4424), .ZN(n4816) );
  INV_X1 U5392 ( .A(n8342), .ZN(n8321) );
  NAND2_X1 U5393 ( .A1(n5055), .A2(n5054), .ZN(n8612) );
  INV_X1 U5394 ( .A(n8052), .ZN(n8362) );
  NOR2_X1 U5395 ( .A1(n7451), .A2(n7786), .ZN(n7664) );
  NOR2_X1 U5396 ( .A1(n8472), .A2(n8783), .ZN(n8493) );
  OAI21_X1 U5397 ( .B1(n8518), .B2(n8517), .A(n8516), .ZN(n4450) );
  OAI21_X1 U5398 ( .B1(n8472), .B2(n4642), .A(n4641), .ZN(n8523) );
  NAND2_X1 U5399 ( .A1(n4643), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4642) );
  INV_X1 U5400 ( .A(n8495), .ZN(n4643) );
  NAND2_X1 U5401 ( .A1(n4585), .A2(n4584), .ZN(n6183) );
  OAI21_X1 U5402 ( .B1(n5522), .B2(n8666), .A(n5521), .ZN(n8554) );
  NOR2_X1 U5403 ( .A1(n5520), .A2(n5519), .ZN(n5521) );
  NOR2_X1 U5404 ( .A1(n6184), .A2(n8548), .ZN(n5519) );
  NAND2_X1 U5405 ( .A1(n5247), .A2(n5246), .ZN(n8041) );
  OR2_X1 U5406 ( .A1(n8755), .A2(n8745), .ZN(n8774) );
  INV_X1 U5407 ( .A(n8210), .ZN(n8805) );
  NAND2_X1 U5408 ( .A1(n5338), .A2(n5337), .ZN(n8854) );
  NAND2_X1 U5409 ( .A1(n8069), .A2(n8202), .ZN(n6786) );
  AND2_X1 U5410 ( .A1(n6591), .A2(n6590), .ZN(n6614) );
  OAI22_X1 U5411 ( .A1(n8946), .A2(n4398), .B1(n4828), .B2(n4354), .ZN(n6639)
         );
  NAND2_X1 U5412 ( .A1(n5923), .A2(n5922), .ZN(n9513) );
  NAND2_X1 U5413 ( .A1(n5934), .A2(n5933), .ZN(n9636) );
  INV_X1 U5414 ( .A(n4645), .ZN(n4644) );
  OAI22_X1 U5415 ( .A1(n5673), .A2(n6673), .B1(n5675), .B2(n6752), .ZN(n4645)
         );
  NAND2_X1 U5416 ( .A1(n5633), .A2(n5632), .ZN(n9445) );
  NAND2_X1 U5417 ( .A1(n4910), .A2(n6056), .ZN(n6057) );
  NOR2_X1 U5418 ( .A1(n6047), .A2(n9934), .ZN(n6058) );
  NAND2_X1 U5419 ( .A1(n6117), .A2(n9142), .ZN(n6059) );
  NAND2_X1 U5420 ( .A1(n5675), .A2(n4579), .ZN(n4578) );
  NOR2_X1 U5421 ( .A1(n6684), .A2(n6669), .ZN(n4579) );
  NAND2_X1 U5422 ( .A1(n4517), .A2(n4515), .ZN(n9061) );
  NAND2_X1 U5423 ( .A1(n9212), .A2(n4516), .ZN(n4515) );
  NAND2_X1 U5424 ( .A1(n9047), .A2(n9155), .ZN(n4517) );
  AOI21_X1 U5425 ( .B1(n6659), .B2(n6285), .A(n6337), .ZN(n6286) );
  OAI21_X1 U5426 ( .B1(n4526), .B2(n4525), .A(n4524), .ZN(n9098) );
  NAND2_X1 U5427 ( .A1(n9093), .A2(n9230), .ZN(n4525) );
  AND2_X1 U5428 ( .A1(n4501), .A2(n4418), .ZN(n4507) );
  NAND2_X1 U5429 ( .A1(n4502), .A2(n9467), .ZN(n4501) );
  AOI21_X1 U5430 ( .B1(n4500), .B2(n4391), .A(n4510), .ZN(n4509) );
  INV_X1 U5431 ( .A(n4502), .ZN(n4500) );
  NOR2_X1 U5432 ( .A1(n6312), .A2(n8580), .ZN(n4452) );
  NAND2_X1 U5433 ( .A1(n6314), .A2(n6313), .ZN(n4453) );
  NAND2_X1 U5434 ( .A1(n9137), .A2(n9136), .ZN(n9156) );
  NAND2_X1 U5435 ( .A1(n9135), .A2(n9155), .ZN(n9136) );
  INV_X1 U5436 ( .A(n5376), .ZN(n4985) );
  AOI21_X1 U5437 ( .B1(n5346), .B2(n4982), .A(SI_20_), .ZN(n4764) );
  NAND2_X1 U5438 ( .A1(n5346), .A2(n4366), .ZN(n4761) );
  INV_X1 U5439 ( .A(n5364), .ZN(n4762) );
  INV_X1 U5440 ( .A(n5301), .ZN(n4969) );
  INV_X1 U5441 ( .A(n4965), .ZN(n4746) );
  INV_X1 U5442 ( .A(n5268), .ZN(n4964) );
  INV_X1 U5443 ( .A(n4774), .ZN(n4767) );
  INV_X1 U5444 ( .A(n4914), .ZN(n4736) );
  INV_X1 U5445 ( .A(SI_11_), .ZN(n7321) );
  INV_X1 U5446 ( .A(SI_14_), .ZN(n7272) );
  INV_X1 U5447 ( .A(n4374), .ZN(n4811) );
  OR2_X1 U5448 ( .A1(n4584), .A2(n6323), .ZN(n4583) );
  OR2_X1 U5449 ( .A1(n5514), .A2(n7573), .ZN(n5071) );
  AND2_X1 U5450 ( .A1(n7004), .A2(n7441), .ZN(n7005) );
  NAND2_X1 U5451 ( .A1(n4542), .A2(n4710), .ZN(n4541) );
  NAND2_X1 U5452 ( .A1(n7708), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4710) );
  NAND2_X1 U5453 ( .A1(n5448), .A2(n5447), .ZN(n5474) );
  NOR2_X1 U5454 ( .A1(n5440), .A2(n4373), .ZN(n4870) );
  INV_X1 U5455 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n7181) );
  NAND2_X1 U5456 ( .A1(n4357), .A2(n4601), .ZN(n4599) );
  NOR2_X1 U5457 ( .A1(n6351), .A2(n4890), .ZN(n4889) );
  INV_X1 U5458 ( .A(n5194), .ZN(n4890) );
  INV_X1 U5459 ( .A(n5117), .ZN(n4864) );
  NOR2_X1 U5460 ( .A1(n8600), .A2(n4876), .ZN(n4875) );
  INV_X1 U5461 ( .A(n5424), .ZN(n4876) );
  INV_X1 U5462 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4801) );
  INV_X1 U5463 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n4817) );
  AND2_X1 U5464 ( .A1(n5212), .A2(n4820), .ZN(n4819) );
  INV_X1 U5465 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n4820) );
  NOR2_X1 U5466 ( .A1(n4467), .A2(n4464), .ZN(n4463) );
  INV_X1 U5467 ( .A(n8967), .ZN(n4464) );
  XNOR2_X1 U5468 ( .A(n6443), .B(n6601), .ZN(n6444) );
  NOR2_X1 U5469 ( .A1(n4359), .A2(n4446), .ZN(n4849) );
  AOI21_X1 U5470 ( .B1(n4361), .B2(n4488), .A(n4426), .ZN(n4482) );
  NAND2_X1 U5471 ( .A1(n4850), .A2(n4396), .ZN(n4844) );
  AND2_X1 U5472 ( .A1(n4850), .A2(n4849), .ZN(n4845) );
  AOI21_X1 U5473 ( .B1(n9197), .B2(n9389), .A(n9196), .ZN(n9199) );
  OAI21_X1 U5474 ( .B1(n9194), .B2(n4370), .A(n4730), .ZN(n9195) );
  OR2_X1 U5475 ( .A1(n9393), .A2(n9147), .ZN(n9148) );
  NAND2_X1 U5476 ( .A1(n9393), .A2(n9150), .ZN(n9160) );
  OR2_X1 U5477 ( .A1(n8135), .A2(n6115), .ZN(n9166) );
  OR2_X1 U5478 ( .A1(n9420), .A2(n6629), .ZN(n9180) );
  INV_X1 U5479 ( .A(n4681), .ZN(n4679) );
  OAI21_X1 U5480 ( .B1(n4653), .B2(n4650), .A(n4360), .ZN(n4649) );
  INV_X1 U5481 ( .A(n5921), .ZN(n4650) );
  INV_X1 U5482 ( .A(n4654), .ZN(n4652) );
  OR2_X1 U5483 ( .A1(n9667), .A2(n9672), .ZN(n4577) );
  NAND2_X1 U5484 ( .A1(n4576), .A2(n9570), .ZN(n4575) );
  INV_X1 U5485 ( .A(n4577), .ZN(n4576) );
  AND2_X1 U5486 ( .A1(n5594), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5789) );
  NOR2_X1 U5487 ( .A1(n7512), .A2(n7801), .ZN(n6029) );
  AND2_X1 U5488 ( .A1(n5593), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5759) );
  OR2_X1 U5489 ( .A1(n5683), .A2(n5659), .ZN(n5661) );
  OR2_X1 U5490 ( .A1(n5469), .A2(n5468), .ZN(n5470) );
  NAND2_X1 U5491 ( .A1(n5463), .A2(n4726), .ZN(n4725) );
  INV_X1 U5492 ( .A(n5463), .ZN(n4727) );
  INV_X1 U5493 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5610) );
  INV_X1 U5494 ( .A(SI_22_), .ZN(n7189) );
  INV_X1 U5495 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6008) );
  INV_X1 U5496 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6009) );
  NOR2_X1 U5497 ( .A1(n4493), .A2(n4371), .ZN(n4492) );
  INV_X1 U5498 ( .A(n4941), .ZN(n4493) );
  INV_X1 U5499 ( .A(SI_7_), .ZN(n7177) );
  INV_X1 U5500 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5604) );
  NOR2_X1 U5501 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n4646) );
  NOR2_X2 U5502 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5672) );
  INV_X1 U5503 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4719) );
  INV_X1 U5504 ( .A(SI_23_), .ZN(n7320) );
  INV_X1 U5505 ( .A(SI_25_), .ZN(n7293) );
  NOR2_X1 U5506 ( .A1(n8214), .A2(n4814), .ZN(n4813) );
  INV_X1 U5507 ( .A(n8148), .ZN(n4814) );
  NAND2_X1 U5508 ( .A1(n8145), .A2(n4374), .ZN(n4815) );
  AND2_X1 U5509 ( .A1(n8316), .A2(n8154), .ZN(n8273) );
  INV_X1 U5510 ( .A(n8698), .ZN(n8278) );
  INV_X1 U5511 ( .A(n4789), .ZN(n4788) );
  OAI21_X1 U5512 ( .B1(n4794), .B2(n4790), .A(n4387), .ZN(n4789) );
  INV_X1 U5513 ( .A(n8019), .ZN(n4790) );
  OR2_X1 U5514 ( .A1(n5151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5166) );
  NAND2_X1 U5515 ( .A1(n5560), .A2(n5013), .ZN(n5019) );
  NOR2_X1 U5516 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n5017) );
  OR2_X1 U5517 ( .A1(n6958), .A2(n7573), .ZN(n7016) );
  OAI22_X1 U5518 ( .A1(n6979), .A2(n7124), .B1(n6959), .B2(n6978), .ZN(n10036)
         );
  AOI22_X1 U5519 ( .A1(n10036), .A2(n10037), .B1(n6980), .B2(n10022), .ZN(
        n10050) );
  AND2_X1 U5520 ( .A1(n4529), .A2(n7489), .ZN(n10054) );
  NAND2_X1 U5521 ( .A1(n4530), .A2(n10046), .ZN(n4529) );
  NAND2_X1 U5522 ( .A1(n10054), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n10053) );
  NAND2_X1 U5523 ( .A1(n7019), .A2(n7488), .ZN(n7492) );
  NAND2_X1 U5524 ( .A1(n7430), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7431) );
  AND2_X1 U5525 ( .A1(n7024), .A2(n7025), .ZN(n7399) );
  OAI21_X1 U5526 ( .B1(n7399), .B2(n4709), .A(n4707), .ZN(n7450) );
  AOI21_X1 U5527 ( .B1(n7025), .B2(n4708), .A(n4448), .ZN(n4707) );
  INV_X1 U5528 ( .A(n7025), .ZN(n4709) );
  NAND2_X1 U5529 ( .A1(n7399), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7398) );
  OR2_X1 U5530 ( .A1(n7809), .A2(n5232), .ZN(n4634) );
  NAND2_X1 U5531 ( .A1(n7807), .A2(n4633), .ZN(n4632) );
  INV_X1 U5532 ( .A(n7809), .ZN(n4633) );
  OR2_X1 U5533 ( .A1(n7706), .A2(n5232), .ZN(n4636) );
  NAND2_X1 U5534 ( .A1(n8400), .A2(n4436), .ZN(n4630) );
  NAND2_X1 U5535 ( .A1(n4629), .A2(n4436), .ZN(n4628) );
  NOR2_X1 U5536 ( .A1(n8459), .A2(n8460), .ZN(n8464) );
  NOR2_X1 U5537 ( .A1(n8482), .A2(n8700), .ZN(n8497) );
  AND2_X1 U5538 ( .A1(n8534), .A2(n8533), .ZN(n8511) );
  NAND2_X1 U5539 ( .A1(n4554), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4553) );
  NAND2_X1 U5540 ( .A1(n8498), .A2(n4554), .ZN(n4552) );
  NAND2_X1 U5541 ( .A1(n8568), .A2(n4590), .ZN(n4584) );
  NOR2_X1 U5542 ( .A1(n8577), .A2(n8669), .ZN(n5520) );
  NAND2_X1 U5543 ( .A1(n5042), .A2(n8252), .ZN(n5433) );
  INV_X1 U5544 ( .A(n5418), .ZN(n5042) );
  OR2_X1 U5545 ( .A1(n5369), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5383) );
  NAND2_X1 U5546 ( .A1(n5037), .A2(n7316), .ZN(n5369) );
  INV_X1 U5547 ( .A(n5354), .ZN(n5037) );
  NAND2_X1 U5548 ( .A1(n5036), .A2(n5035), .ZN(n5339) );
  INV_X1 U5549 ( .A(n5327), .ZN(n5036) );
  NAND2_X1 U5550 ( .A1(n5034), .A2(n7181), .ZN(n5312) );
  INV_X1 U5551 ( .A(n5294), .ZN(n5034) );
  OR2_X1 U5552 ( .A1(n5278), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5294) );
  OR2_X1 U5553 ( .A1(n5261), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5278) );
  NAND2_X1 U5554 ( .A1(n5033), .A2(n5032), .ZN(n5261) );
  INV_X1 U5555 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5032) );
  INV_X1 U5556 ( .A(n5248), .ZN(n5033) );
  NAND2_X1 U5557 ( .A1(n7782), .A2(n5208), .ZN(n7887) );
  NAND2_X1 U5558 ( .A1(n5031), .A2(n5030), .ZN(n5218) );
  INV_X1 U5559 ( .A(n5195), .ZN(n5031) );
  NAND2_X1 U5560 ( .A1(n5029), .A2(n5028), .ZN(n5180) );
  INV_X1 U5561 ( .A(n5166), .ZN(n5029) );
  NAND2_X1 U5562 ( .A1(n4881), .A2(n5177), .ZN(n4880) );
  NOR2_X1 U5563 ( .A1(n5178), .A2(n4884), .ZN(n4883) );
  INV_X1 U5564 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5024) );
  OR2_X1 U5565 ( .A1(n5101), .A2(n5099), .ZN(n5102) );
  AND2_X1 U5566 ( .A1(n5566), .A2(n5565), .ZN(n6140) );
  AND3_X1 U5567 ( .A1(n6879), .A2(n6141), .A3(n6864), .ZN(n7371) );
  OR2_X1 U5568 ( .A1(n7369), .A2(n6146), .ZN(n7373) );
  NAND2_X1 U5569 ( .A1(n4877), .A2(n5424), .ZN(n8601) );
  AND2_X1 U5570 ( .A1(n6305), .A2(n5541), .ZN(n8600) );
  OAI21_X1 U5571 ( .B1(n4609), .B2(n4376), .A(n4608), .ZN(n4607) );
  INV_X1 U5572 ( .A(n6337), .ZN(n4608) );
  AOI21_X1 U5573 ( .B1(n4614), .B2(n6342), .A(n4613), .ZN(n4612) );
  AND2_X1 U5574 ( .A1(n6289), .A2(n8647), .ZN(n8664) );
  NAND2_X1 U5575 ( .A1(n4857), .A2(n4854), .ZN(n8677) );
  INV_X1 U5576 ( .A(n4855), .ZN(n4854) );
  OAI22_X1 U5577 ( .A1(n5345), .A2(n4856), .B1(n8854), .B2(n8698), .ZN(n4855)
         );
  AND2_X1 U5578 ( .A1(n6280), .A2(n6287), .ZN(n8676) );
  OR2_X1 U5579 ( .A1(n6343), .A2(n6342), .ZN(n8687) );
  AND2_X1 U5580 ( .A1(n6258), .A2(n6259), .ZN(n8113) );
  OAI21_X1 U5581 ( .B1(n5239), .B2(n4896), .A(n4894), .ZN(n5267) );
  INV_X1 U5582 ( .A(n4895), .ZN(n4894) );
  OAI21_X1 U5583 ( .B1(n4897), .B2(n4896), .A(n6345), .ZN(n4895) );
  AND2_X1 U5584 ( .A1(n5215), .A2(n5214), .ZN(n8053) );
  OR2_X1 U5585 ( .A1(n6142), .A2(n7570), .ZN(n6875) );
  MUX2_X1 U5586 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5559), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5561) );
  OAI21_X1 U5587 ( .B1(n5578), .B2(n5558), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5559) );
  XNOR2_X1 U5588 ( .A(n5580), .B(n5579), .ZN(n6865) );
  INV_X1 U5589 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5001) );
  INV_X1 U5590 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5090) );
  INV_X1 U5591 ( .A(n9445), .ZN(n6643) );
  AOI21_X1 U5592 ( .B1(n4825), .B2(n4827), .A(n4824), .ZN(n4823) );
  INV_X1 U5593 ( .A(n8917), .ZN(n4831) );
  INV_X1 U5594 ( .A(n6471), .ZN(n4456) );
  INV_X1 U5595 ( .A(n6420), .ZN(n6404) );
  NAND2_X1 U5596 ( .A1(n8925), .A2(n8927), .ZN(n8926) );
  OR2_X1 U5597 ( .A1(n5948), .A2(n5600), .ZN(n5960) );
  AND2_X1 U5598 ( .A1(n6574), .A2(n6573), .ZN(n8945) );
  NAND2_X1 U5599 ( .A1(n6438), .A2(n6437), .ZN(n6439) );
  NOR2_X1 U5600 ( .A1(n6411), .A2(n6406), .ZN(n6792) );
  AND2_X1 U5601 ( .A1(n6607), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6406) );
  AOI21_X1 U5602 ( .B1(n6843), .B2(n6603), .A(n6408), .ZN(n6409) );
  NAND2_X1 U5603 ( .A1(n5598), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5916) );
  INV_X1 U5604 ( .A(n5908), .ZN(n5598) );
  OR2_X1 U5605 ( .A1(n6543), .A2(n6542), .ZN(n6544) );
  INV_X1 U5606 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5832) );
  NAND2_X1 U5607 ( .A1(n4839), .A2(n4844), .ZN(n7873) );
  NAND2_X1 U5608 ( .A1(n4848), .A2(n4845), .ZN(n4839) );
  AOI21_X1 U5609 ( .B1(n9284), .B2(n6407), .A(n6425), .ZN(n6427) );
  INV_X1 U5610 ( .A(n5878), .ZN(n5597) );
  OR2_X1 U5611 ( .A1(n5895), .A2(n5894), .ZN(n5908) );
  NAND2_X1 U5612 ( .A1(n8916), .A2(n8917), .ZN(n8988) );
  NAND2_X1 U5613 ( .A1(n4472), .A2(n6515), .ZN(n8995) );
  NAND2_X1 U5614 ( .A1(n5596), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5866) );
  NAND2_X1 U5615 ( .A1(n9200), .A2(n9265), .ZN(n4519) );
  OR2_X1 U5616 ( .A1(n9153), .A2(n4732), .ZN(n9257) );
  NAND2_X1 U5617 ( .A1(n5897), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5680) );
  NAND2_X1 U5618 ( .A1(n6007), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5888) );
  INV_X1 U5619 ( .A(n4703), .ZN(n6117) );
  INV_X1 U5620 ( .A(n4581), .ZN(n6129) );
  AND2_X1 U5621 ( .A1(n9179), .A2(n9178), .ZN(n9434) );
  NAND2_X1 U5622 ( .A1(n4673), .A2(n5981), .ZN(n4672) );
  INV_X1 U5623 ( .A(n4670), .ZN(n4669) );
  NAND2_X1 U5624 ( .A1(n4702), .A2(n9172), .ZN(n9441) );
  NAND2_X1 U5625 ( .A1(n9512), .A2(n9495), .ZN(n9490) );
  NAND2_X1 U5626 ( .A1(n4557), .A2(n4555), .ZN(n9504) );
  NOR2_X1 U5627 ( .A1(n4556), .A2(n6040), .ZN(n4555) );
  INV_X1 U5628 ( .A(n9510), .ZN(n4556) );
  AND2_X1 U5629 ( .A1(n9118), .A2(n9117), .ZN(n9510) );
  AND2_X1 U5630 ( .A1(n4557), .A2(n9116), .ZN(n9505) );
  NAND2_X1 U5631 ( .A1(n6039), .A2(n9248), .ZN(n9531) );
  NOR2_X1 U5632 ( .A1(n8010), .A2(n4577), .ZN(n9589) );
  NOR2_X1 U5633 ( .A1(n8010), .A2(n9672), .ZN(n9588) );
  OR2_X1 U5634 ( .A1(n5833), .A2(n5832), .ZN(n5850) );
  OAI21_X1 U5635 ( .B1(n4688), .B2(n4687), .A(n4352), .ZN(n4686) );
  AND2_X1 U5636 ( .A1(n9227), .A2(n9230), .ZN(n9034) );
  NAND2_X1 U5637 ( .A1(n5789), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5820) );
  INV_X1 U5638 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5819) );
  NAND2_X1 U5639 ( .A1(n4560), .A2(n5788), .ZN(n7391) );
  NAND2_X1 U5640 ( .A1(n6701), .A2(n9014), .ZN(n4560) );
  NAND2_X1 U5641 ( .A1(n9941), .A2(n4571), .ZN(n7564) );
  AND2_X1 U5642 ( .A1(n9222), .A2(n6034), .ZN(n4566) );
  NAND2_X1 U5643 ( .A1(n4664), .A2(n4665), .ZN(n7471) );
  AOI21_X1 U5644 ( .B1(n7109), .B2(n4666), .A(n4399), .ZN(n4665) );
  INV_X1 U5645 ( .A(n5730), .ZN(n4666) );
  INV_X1 U5646 ( .A(n6848), .ZN(n4499) );
  NAND2_X1 U5647 ( .A1(n5638), .A2(n5637), .ZN(n9616) );
  NAND2_X1 U5648 ( .A1(n5972), .A2(n5971), .ZN(n9452) );
  NAND2_X1 U5649 ( .A1(n5958), .A2(n5957), .ZN(n9626) );
  INV_X1 U5650 ( .A(n10004), .ZN(n9680) );
  OAI21_X1 U5651 ( .B1(n9718), .B2(P1_D_REG_0__SCAN_IN), .A(n9721), .ZN(n6708)
         );
  INV_X1 U5652 ( .A(n6813), .ZN(n6843) );
  XNOR2_X1 U5653 ( .A(n5444), .B(n5460), .ZN(n8070) );
  NAND2_X1 U5654 ( .A1(n5443), .A2(n5467), .ZN(n5444) );
  XNOR2_X1 U5655 ( .A(n6082), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6097) );
  INV_X1 U5656 ( .A(n6072), .ZN(n6074) );
  NOR2_X1 U5657 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n6073) );
  OR2_X1 U5658 ( .A1(n6069), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n6078) );
  XNOR2_X1 U5659 ( .A(n5413), .B(n5412), .ZN(n5956) );
  XNOR2_X1 U5660 ( .A(n6068), .B(n6067), .ZN(n6685) );
  NAND2_X1 U5661 ( .A1(n6015), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6017) );
  XNOR2_X1 U5662 ( .A(n5209), .B(n4379), .ZN(n6701) );
  NAND2_X1 U5663 ( .A1(n4734), .A2(n4737), .ZN(n5201) );
  OR2_X1 U5664 ( .A1(n5174), .A2(n4740), .ZN(n4734) );
  CLKBUF_X1 U5665 ( .A(n5741), .Z(n5742) );
  OR2_X1 U5666 ( .A1(n7857), .A2(n7864), .ZN(n7858) );
  OAI21_X1 U5667 ( .B1(n8187), .B2(n4785), .A(n4782), .ZN(n8206) );
  NAND2_X1 U5668 ( .A1(n4815), .A2(n8148), .ZN(n8213) );
  INV_X1 U5669 ( .A(n8628), .ZN(n8253) );
  INV_X1 U5670 ( .A(n4778), .ZN(n4777) );
  OAI22_X1 U5671 ( .A1(n8205), .A2(n4779), .B1(n8190), .B2(n8589), .ZN(n4778)
         );
  NAND2_X1 U5672 ( .A1(n5473), .A2(n5472), .ZN(n8197) );
  NAND2_X1 U5673 ( .A1(n7953), .A2(n4794), .ZN(n8020) );
  NAND2_X1 U5674 ( .A1(n5023), .A2(n5022), .ZN(n8256) );
  NOR2_X1 U5675 ( .A1(n7363), .A2(n7578), .ZN(n4803) );
  AND2_X1 U5676 ( .A1(n4809), .A2(n4808), .ZN(n7537) );
  INV_X1 U5677 ( .A(n8351), .ZN(n8324) );
  NAND2_X1 U5678 ( .A1(n6874), .A2(n6873), .ZN(n8335) );
  NAND2_X1 U5679 ( .A1(n6916), .A2(n4375), .ZN(n6908) );
  AND2_X1 U5680 ( .A1(n6887), .A2(n6886), .ZN(n8342) );
  NAND2_X1 U5681 ( .A1(n6881), .A2(n10064), .ZN(n8339) );
  NAND2_X1 U5682 ( .A1(n8187), .A2(n8186), .ZN(n8334) );
  NAND2_X1 U5683 ( .A1(n5432), .A2(n5431), .ZN(n5542) );
  AND4_X1 U5684 ( .A1(n5317), .A2(n5316), .A3(n5315), .A4(n5314), .ZN(n8346)
         );
  NAND2_X1 U5685 ( .A1(n6912), .A2(n6877), .ZN(n8347) );
  OR2_X1 U5686 ( .A1(n8260), .A2(n8343), .ZN(n8344) );
  AND2_X1 U5687 ( .A1(n6912), .A2(n6911), .ZN(n8351) );
  XNOR2_X1 U5688 ( .A(n5500), .B(P2_IR_REG_22__SCAN_IN), .ZN(n6392) );
  AND2_X1 U5689 ( .A1(n6168), .A2(n6167), .ZN(n8549) );
  NAND2_X1 U5690 ( .A1(n5481), .A2(n5480), .ZN(n8357) );
  INV_X1 U5691 ( .A(n8312), .ZN(n8641) );
  OAI211_X1 U5692 ( .C1(n5514), .C2(n8643), .A(n5395), .B(n5394), .ZN(n8655)
         );
  CLKBUF_X1 U5693 ( .A(n6878), .Z(n8371) );
  NAND2_X1 U5694 ( .A1(n5405), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5063) );
  INV_X1 U5695 ( .A(n8359), .ZN(n8512) );
  NOR2_X1 U5696 ( .A1(n4639), .A2(n7650), .ZN(n7649) );
  NOR2_X1 U5697 ( .A1(n7650), .A2(n4637), .ZN(n7653) );
  INV_X1 U5698 ( .A(n4639), .ZN(n4637) );
  INV_X1 U5699 ( .A(n4542), .ZN(n4539) );
  INV_X1 U5700 ( .A(n4636), .ZN(n7808) );
  NAND2_X1 U5701 ( .A1(n4632), .A2(n4631), .ZN(n8383) );
  NAND2_X1 U5702 ( .A1(n4548), .A2(n4547), .ZN(n8387) );
  INV_X1 U5703 ( .A(n4714), .ZN(n8404) );
  AND2_X1 U5704 ( .A1(n4714), .A2(n4715), .ZN(n8407) );
  NAND2_X1 U5705 ( .A1(n4534), .A2(n4532), .ZN(n8426) );
  NOR2_X1 U5706 ( .A1(n8398), .A2(n8399), .ZN(n8401) );
  NAND2_X1 U5707 ( .A1(n6178), .A2(n6177), .ZN(n8741) );
  AOI21_X1 U5708 ( .B1(n9010), .B2(n6175), .A(n6160), .ZN(n8746) );
  OAI21_X1 U5709 ( .B1(n8567), .B2(n8666), .A(n8566), .ZN(n8748) );
  NOR2_X1 U5710 ( .A1(n8565), .A2(n8564), .ZN(n8566) );
  NOR2_X1 U5711 ( .A1(n8589), .A2(n8669), .ZN(n8564) );
  NAND2_X1 U5712 ( .A1(n5368), .A2(n5367), .ZN(n8773) );
  NAND2_X1 U5713 ( .A1(n5293), .A2(n5292), .ZN(n8792) );
  NAND2_X1 U5714 ( .A1(n5260), .A2(n5259), .ZN(n8077) );
  NAND2_X1 U5715 ( .A1(n7974), .A2(n5254), .ZN(n8002) );
  AND2_X1 U5716 ( .A1(n5239), .A2(n5238), .ZN(n7976) );
  NAND2_X1 U5717 ( .A1(n5532), .A2(n6230), .ZN(n7886) );
  AND3_X1 U5718 ( .A1(n5193), .A2(n5192), .A3(n5191), .ZN(n7954) );
  NAND2_X1 U5719 ( .A1(n7547), .A2(n6348), .ZN(n4885) );
  AND2_X1 U5720 ( .A1(n4595), .A2(n4597), .ZN(n7689) );
  NAND2_X1 U5721 ( .A1(n6945), .A2(n6946), .ZN(n6944) );
  NAND2_X1 U5722 ( .A1(n7626), .A2(n6199), .ZN(n6945) );
  NAND2_X1 U5723 ( .A1(n6880), .A2(n6879), .ZN(n10064) );
  NAND2_X1 U5724 ( .A1(n8715), .A2(n7571), .ZN(n8738) );
  INV_X1 U5725 ( .A(n8734), .ZN(n8715) );
  NOR2_X1 U5726 ( .A1(n8554), .A2(n5545), .ZN(n6149) );
  INV_X1 U5727 ( .A(n8197), .ZN(n8801) );
  INV_X1 U5728 ( .A(n5542), .ZN(n8807) );
  NAND2_X1 U5729 ( .A1(n4867), .A2(n4873), .ZN(n8586) );
  NAND2_X1 U5730 ( .A1(n4878), .A2(n4373), .ZN(n4867) );
  INV_X1 U5731 ( .A(n8256), .ZN(n8812) );
  NAND2_X1 U5732 ( .A1(n4611), .A2(n4376), .ZN(n8618) );
  NAND2_X1 U5733 ( .A1(n5402), .A2(n5401), .ZN(n8824) );
  NAND2_X1 U5734 ( .A1(n4611), .A2(n6292), .ZN(n8625) );
  NAND2_X1 U5735 ( .A1(n5391), .A2(n5390), .ZN(n8830) );
  NAND2_X1 U5736 ( .A1(n5380), .A2(n5379), .ZN(n8836) );
  NAND2_X1 U5737 ( .A1(n5353), .A2(n5352), .ZN(n8848) );
  NAND2_X1 U5738 ( .A1(n5326), .A2(n5325), .ZN(n8860) );
  NAND2_X1 U5739 ( .A1(n5311), .A2(n5310), .ZN(n8867) );
  NAND2_X1 U5740 ( .A1(n5277), .A2(n5276), .ZN(n8149) );
  INV_X1 U5741 ( .A(n8841), .ZN(n8866) );
  CLKBUF_X1 U5742 ( .A(n5523), .Z(n7905) );
  INV_X1 U5743 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5045) );
  INV_X1 U5744 ( .A(n5563), .ZN(n8069) );
  NAND2_X1 U5745 ( .A1(n5551), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5552) );
  NAND2_X1 U5746 ( .A1(n5547), .A2(n5546), .ZN(n5550) );
  AND2_X1 U5747 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5546) );
  XNOR2_X1 U5748 ( .A(n5503), .B(n5502), .ZN(n7846) );
  NAND2_X1 U5749 ( .A1(n5507), .A2(n5506), .ZN(n7687) );
  NAND2_X1 U5750 ( .A1(n4796), .A2(n4795), .ZN(n5351) );
  AOI21_X1 U5751 ( .B1(n4798), .B2(n4800), .A(n4800), .ZN(n4795) );
  INV_X1 U5752 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6699) );
  INV_X1 U5753 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6691) );
  OR2_X1 U5754 ( .A1(n5161), .A2(n5160), .ZN(n7419) );
  NOR2_X1 U5755 ( .A1(n5111), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5141) );
  NAND2_X1 U5756 ( .A1(n4537), .A2(n4800), .ZN(n4536) );
  INV_X1 U5757 ( .A(n9280), .ZN(n7478) );
  INV_X1 U5758 ( .A(n4838), .ZN(n4837) );
  NAND2_X1 U5759 ( .A1(n6506), .A2(n6509), .ZN(n7985) );
  INV_X1 U5760 ( .A(n8965), .ZN(n4462) );
  NAND2_X1 U5761 ( .A1(n5906), .A2(n5905), .ZN(n9652) );
  INV_X1 U5762 ( .A(n9931), .ZN(n7681) );
  OR2_X1 U5763 ( .A1(n8901), .A2(n4488), .ZN(n4485) );
  AND3_X1 U5764 ( .A1(n6619), .A2(n7513), .A3(n6620), .ZN(n8999) );
  AND2_X1 U5765 ( .A1(n5690), .A2(n5689), .ZN(n7077) );
  NAND2_X1 U5766 ( .A1(n5918), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5690) );
  NOR2_X1 U5767 ( .A1(n4386), .A2(n5688), .ZN(n5689) );
  NOR2_X1 U5768 ( .A1(n7829), .A2(n4457), .ZN(n7834) );
  INV_X1 U5769 ( .A(n7830), .ZN(n4458) );
  NAND2_X1 U5770 ( .A1(n4834), .A2(n6544), .ZN(n8953) );
  NAND2_X1 U5771 ( .A1(n8901), .A2(n8902), .ZN(n4834) );
  NAND2_X1 U5772 ( .A1(n7848), .A2(n7849), .ZN(n7847) );
  NAND2_X1 U5773 ( .A1(n7755), .A2(n6497), .ZN(n7848) );
  INV_X1 U5774 ( .A(n9008), .ZN(n8972) );
  NAND2_X1 U5775 ( .A1(n4479), .A2(n4478), .ZN(n4477) );
  INV_X1 U5776 ( .A(n8990), .ZN(n4478) );
  NAND2_X1 U5777 ( .A1(n8988), .A2(n8987), .ZN(n4479) );
  AND2_X1 U5778 ( .A1(n8989), .A2(n8997), .ZN(n4476) );
  INV_X1 U5779 ( .A(n9277), .ZN(n9002) );
  NAND2_X1 U5780 ( .A1(n6626), .A2(n9273), .ZN(n9004) );
  OAI21_X1 U5781 ( .B1(n4520), .B2(n4518), .A(n9206), .ZN(n9269) );
  NAND2_X1 U5782 ( .A1(n4519), .A2(n6096), .ZN(n4518) );
  AOI21_X1 U5783 ( .B1(n9205), .B2(n9381), .A(n9204), .ZN(n9206) );
  AOI21_X1 U5784 ( .B1(n9264), .B2(n6021), .A(n6397), .ZN(n4520) );
  NAND2_X1 U5785 ( .A1(n5994), .A2(n5993), .ZN(n9435) );
  OR2_X1 U5786 ( .A1(n6641), .A2(n6050), .ZN(n5994) );
  NAND2_X1 U5787 ( .A1(n5980), .A2(n5979), .ZN(n9471) );
  OR2_X1 U5788 ( .A1(n9454), .A2(n6050), .ZN(n5980) );
  NAND2_X1 U5789 ( .A1(n5970), .A2(n5969), .ZN(n9477) );
  INV_X1 U5790 ( .A(n7077), .ZN(n9283) );
  OR2_X1 U5791 ( .A1(n5683), .A2(n5650), .ZN(n5655) );
  OR2_X1 U5792 ( .A1(n9892), .A2(n9891), .ZN(n9901) );
  AOI21_X1 U5793 ( .B1(n6128), .B2(n9906), .A(n6127), .ZN(n8141) );
  NAND2_X1 U5794 ( .A1(n6126), .A2(n6125), .ZN(n6127) );
  NAND2_X1 U5795 ( .A1(n9415), .A2(n9906), .ZN(n4569) );
  OAI21_X1 U5796 ( .B1(n9489), .B2(n4676), .A(n4674), .ZN(n9448) );
  NAND2_X1 U5797 ( .A1(n4677), .A2(n4680), .ZN(n9460) );
  NAND2_X1 U5798 ( .A1(n9489), .A2(n4681), .ZN(n4677) );
  NAND2_X1 U5799 ( .A1(n9489), .A2(n5943), .ZN(n4684) );
  OAI21_X1 U5800 ( .B1(n9565), .B2(n4654), .A(n4653), .ZN(n9522) );
  NAND2_X1 U5801 ( .A1(n4655), .A2(n4659), .ZN(n9537) );
  NAND2_X1 U5802 ( .A1(n9565), .A2(n4660), .ZN(n4655) );
  AND2_X1 U5803 ( .A1(n4563), .A2(n9236), .ZN(n9557) );
  AND2_X1 U5804 ( .A1(n4661), .A2(n4663), .ZN(n9550) );
  NAND2_X1 U5805 ( .A1(n9565), .A2(n5886), .ZN(n4661) );
  NAND2_X1 U5806 ( .A1(n4694), .A2(n9237), .ZN(n9572) );
  AND2_X1 U5807 ( .A1(n4567), .A2(n4696), .ZN(n8013) );
  NAND2_X1 U5808 ( .A1(n7767), .A2(n9230), .ZN(n7912) );
  NAND2_X1 U5809 ( .A1(n4685), .A2(n4688), .ZN(n9916) );
  NAND2_X1 U5810 ( .A1(n7381), .A2(n4690), .ZN(n4685) );
  AOI21_X1 U5811 ( .B1(n7381), .B2(n9018), .A(n4691), .ZN(n7557) );
  NAND2_X1 U5812 ( .A1(n4481), .A2(n5758), .ZN(n9940) );
  NAND2_X1 U5813 ( .A1(n6690), .A2(n9014), .ZN(n4481) );
  NAND2_X1 U5814 ( .A1(n7110), .A2(n7109), .ZN(n7108) );
  NAND2_X1 U5815 ( .A1(n6893), .A2(n5730), .ZN(n7110) );
  OR2_X1 U5816 ( .A1(n9576), .A2(n6892), .ZN(n9601) );
  INV_X1 U5817 ( .A(n9405), .ZN(n9949) );
  NAND2_X1 U5818 ( .A1(n7941), .A2(n6397), .ZN(n6717) );
  INV_X1 U5819 ( .A(n9515), .ZN(n9952) );
  NAND2_X1 U5820 ( .A1(n5755), .A2(n4705), .ZN(n7598) );
  NAND2_X1 U5821 ( .A1(n4706), .A2(n9014), .ZN(n4705) );
  INV_X1 U5822 ( .A(n6681), .ZN(n4706) );
  INV_X1 U5823 ( .A(n10021), .ZN(n10019) );
  AND2_X1 U5824 ( .A1(n9017), .A2(n9016), .ZN(n9687) );
  NAND2_X1 U5825 ( .A1(n5997), .A2(n5996), .ZN(n9402) );
  INV_X1 U5826 ( .A(n9420), .ZN(n6061) );
  INV_X1 U5827 ( .A(n9452), .ZN(n9699) );
  INV_X1 U5828 ( .A(n9483), .ZN(n9704) );
  INV_X1 U5829 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5620) );
  INV_X1 U5830 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5634) );
  NAND2_X1 U5831 ( .A1(n5621), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5635) );
  OAI21_X1 U5832 ( .B1(n6069), .B2(n4365), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n4667) );
  NAND2_X1 U5833 ( .A1(n6076), .A2(n6075), .ZN(n7997) );
  OR2_X1 U5834 ( .A1(n6071), .A2(n6070), .ZN(n6076) );
  NOR2_X1 U5835 ( .A1(n6074), .A2(n6073), .ZN(n6075) );
  INV_X1 U5836 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6070) );
  AND2_X1 U5837 ( .A1(n4751), .A2(n4748), .ZN(n5335) );
  INV_X1 U5838 ( .A(n4753), .ZN(n4748) );
  NAND2_X1 U5839 ( .A1(n4771), .A2(n4769), .ZN(n5243) );
  NAND2_X1 U5840 ( .A1(n4771), .A2(n4772), .ZN(n5241) );
  INV_X1 U5841 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6693) );
  XNOR2_X1 U5842 ( .A(n5174), .B(n5173), .ZN(n6681) );
  NAND2_X1 U5843 ( .A1(n4942), .A2(n4941), .ZN(n5163) );
  AOI21_X1 U5844 ( .B1(n8519), .B2(n10056), .A(n4450), .ZN(n4449) );
  MUX2_X1 U5845 ( .A(n8802), .B(n8753), .S(n8755), .Z(n8754) );
  MUX2_X1 U5846 ( .A(n8803), .B(n8802), .S(n10088), .Z(n8804) );
  AND2_X1 U5847 ( .A1(n6615), .A2(n8997), .ZN(n6634) );
  NAND2_X1 U5848 ( .A1(n4475), .A2(n4473), .ZN(P1_U3240) );
  INV_X1 U5849 ( .A(n4474), .ZN(n4473) );
  NAND2_X1 U5850 ( .A1(n4477), .A2(n4476), .ZN(n4475) );
  OAI21_X1 U5851 ( .B1(n9431), .B2(n9008), .A(n8994), .ZN(n4474) );
  INV_X4 U5852 ( .A(n6507), .ZN(n6407) );
  OR2_X1 U5853 ( .A1(n9914), .A2(n9278), .ZN(n4352) );
  AND2_X1 U5854 ( .A1(n6234), .A2(n6230), .ZN(n6351) );
  AND2_X1 U5855 ( .A1(n4571), .A2(n4570), .ZN(n4353) );
  OR2_X1 U5856 ( .A1(n9662), .A2(n6037), .ZN(n9236) );
  OR2_X1 U5857 ( .A1(n9647), .A2(n8903), .ZN(n9116) );
  AND2_X2 U5858 ( .A1(n5626), .A2(n5623), .ZN(n5684) );
  INV_X1 U5859 ( .A(n8611), .ZN(n4878) );
  OR2_X1 U5860 ( .A1(n6598), .A2(n6597), .ZN(n4354) );
  AND2_X1 U5861 ( .A1(n7498), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4355) );
  OR2_X1 U5862 ( .A1(n9626), .A2(n9477), .ZN(n4356) );
  OR2_X1 U5863 ( .A1(n8082), .A2(n8360), .ZN(n4357) );
  NOR2_X1 U5864 ( .A1(n8171), .A2(n8240), .ZN(n4358) );
  INV_X1 U5865 ( .A(n6340), .ZN(n4862) );
  AND2_X1 U5866 ( .A1(n6454), .A2(n6453), .ZN(n4359) );
  OR2_X1 U5867 ( .A1(n9647), .A2(n9546), .ZN(n4360) );
  AND2_X1 U5868 ( .A1(n4486), .A2(n4484), .ZN(n4361) );
  AND2_X1 U5869 ( .A1(n4970), .A2(n4422), .ZN(n4362) );
  AND2_X1 U5870 ( .A1(n9393), .A2(n4732), .ZN(n4363) );
  AND2_X1 U5871 ( .A1(n6669), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4364) );
  NAND2_X1 U5872 ( .A1(n4915), .A2(n4852), .ZN(n4365) );
  NAND2_X1 U5873 ( .A1(n5818), .A2(n5817), .ZN(n9914) );
  INV_X1 U5874 ( .A(n9915), .ZN(n4687) );
  AND2_X1 U5875 ( .A1(n4982), .A2(SI_20_), .ZN(n4366) );
  INV_X1 U5876 ( .A(n8944), .ZN(n4467) );
  OR2_X1 U5877 ( .A1(n8406), .A2(n8377), .ZN(n4367) );
  NAND2_X1 U5878 ( .A1(n7736), .A2(n4889), .ZN(n7782) );
  NOR2_X1 U5879 ( .A1(n7664), .A2(n4712), .ZN(n4368) );
  NAND2_X1 U5880 ( .A1(n9013), .A2(n9012), .ZN(n9393) );
  OR2_X1 U5881 ( .A1(n9636), .A2(n9507), .ZN(n4369) );
  OR2_X1 U5882 ( .A1(n9168), .A2(n9167), .ZN(n4370) );
  AND2_X1 U5883 ( .A1(n4943), .A2(SI_6_), .ZN(n4371) );
  OAI211_X1 U5884 ( .C1(n5088), .C2(n10022), .A(n5098), .B(n5097), .ZN(n5099)
         );
  NAND2_X1 U5885 ( .A1(n4786), .A2(n4892), .ZN(n5159) );
  NAND3_X1 U5886 ( .A1(n4853), .A2(n5615), .A3(n5609), .ZN(n6069) );
  INV_X1 U5887 ( .A(n6339), .ZN(n4610) );
  OR2_X1 U5888 ( .A1(n8818), .A2(n8628), .ZN(n4372) );
  AND2_X1 U5889 ( .A1(n4879), .A2(n4372), .ZN(n4373) );
  NAND2_X1 U5890 ( .A1(n8146), .A2(n8144), .ZN(n4374) );
  OR2_X1 U5891 ( .A1(n6907), .A2(n8371), .ZN(n4375) );
  AND2_X1 U5892 ( .A1(n4610), .A2(n6292), .ZN(n4376) );
  INV_X1 U5893 ( .A(n7807), .ZN(n4635) );
  AND2_X1 U5894 ( .A1(n9657), .A2(n9574), .ZN(n4377) );
  NAND2_X1 U5895 ( .A1(n5658), .A2(n4578), .ZN(n6835) );
  AND2_X1 U5896 ( .A1(n9483), .A2(n9499), .ZN(n4378) );
  XNOR2_X1 U5897 ( .A(n8197), .B(n8357), .ZN(n8191) );
  INV_X1 U5898 ( .A(n8191), .ZN(n8568) );
  OR2_X1 U5899 ( .A1(n8558), .A2(n8563), .ZN(n6321) );
  NAND2_X1 U5900 ( .A1(n4485), .A2(n4486), .ZN(n8909) );
  XOR2_X1 U5901 ( .A(n4957), .B(SI_10_), .Z(n4379) );
  OR2_X1 U5902 ( .A1(n4964), .A2(n7272), .ZN(n4380) );
  AND2_X1 U5903 ( .A1(n9652), .A2(n9559), .ZN(n4381) );
  INV_X1 U5904 ( .A(n6878), .ZN(n7630) );
  NAND2_X1 U5905 ( .A1(n5675), .A2(n4350), .ZN(n5887) );
  INV_X2 U5906 ( .A(n5887), .ZN(n9014) );
  NAND2_X1 U5907 ( .A1(n5775), .A2(n5774), .ZN(n7512) );
  AND2_X1 U5908 ( .A1(n8955), .A2(n8954), .ZN(n4382) );
  NOR2_X1 U5909 ( .A1(n5111), .A2(n4893), .ZN(n5157) );
  NAND2_X1 U5910 ( .A1(n9476), .A2(n9481), .ZN(n9466) );
  NAND2_X1 U5911 ( .A1(n4891), .A2(n5362), .ZN(n8662) );
  AND2_X1 U5912 ( .A1(n4468), .A2(n8884), .ZN(n4383) );
  NAND2_X1 U5913 ( .A1(n8964), .A2(n8967), .ZN(n8884) );
  AND2_X1 U5914 ( .A1(n9123), .A2(n9124), .ZN(n9498) );
  INV_X1 U5915 ( .A(n9467), .ZN(n4510) );
  NAND2_X1 U5916 ( .A1(n4606), .A2(n4786), .ZN(n5189) );
  AND2_X1 U5917 ( .A1(n4696), .A2(n9036), .ZN(n4384) );
  NOR2_X1 U5918 ( .A1(n8955), .A2(n8954), .ZN(n4385) );
  NOR2_X1 U5919 ( .A1(n5683), .A2(n5682), .ZN(n4386) );
  NAND2_X1 U5920 ( .A1(n6114), .A2(n6113), .ZN(n8135) );
  INV_X1 U5921 ( .A(n8135), .ZN(n4580) );
  OR2_X1 U5922 ( .A1(n8018), .A2(n8365), .ZN(n4387) );
  AND2_X1 U5923 ( .A1(n4788), .A2(n8292), .ZN(n4388) );
  NOR2_X1 U5924 ( .A1(n8493), .A2(n8494), .ZN(n4389) );
  OR2_X1 U5925 ( .A1(n8741), .A2(n8549), .ZN(n4390) );
  NAND2_X1 U5926 ( .A1(n4503), .A2(n9498), .ZN(n4391) );
  OR2_X1 U5927 ( .A1(n9402), .A2(n6110), .ZN(n9142) );
  AND2_X1 U5928 ( .A1(n9626), .A2(n9477), .ZN(n4392) );
  NAND2_X1 U5929 ( .A1(n6370), .A2(n8741), .ZN(n4393) );
  OR3_X1 U5930 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .A3(
        P1_IR_REG_30__SCAN_IN), .ZN(n4394) );
  AND2_X1 U5931 ( .A1(n6258), .A2(n4599), .ZN(n4395) );
  INV_X1 U5932 ( .A(n4713), .ZN(n4712) );
  NAND2_X1 U5933 ( .A1(n7665), .A2(n7666), .ZN(n4713) );
  INV_X1 U5934 ( .A(n5177), .ZN(n5178) );
  NAND2_X1 U5935 ( .A1(n6474), .A2(n4846), .ZN(n4396) );
  AND2_X1 U5936 ( .A1(n8860), .A2(n8688), .ZN(n4397) );
  INV_X1 U5937 ( .A(n8405), .ZN(n4715) );
  OR2_X1 U5938 ( .A1(n4354), .A2(n4831), .ZN(n4398) );
  INV_X1 U5939 ( .A(n4592), .ZN(n4591) );
  NOR2_X1 U5940 ( .A1(n8589), .A2(n8210), .ZN(n4592) );
  INV_X1 U5941 ( .A(n6034), .ZN(n9018) );
  AND2_X1 U5942 ( .A1(n9080), .A2(n9076), .ZN(n6034) );
  AND2_X1 U5943 ( .A1(n7478), .A2(n9975), .ZN(n4399) );
  NOR2_X1 U5944 ( .A1(n4626), .A2(n4625), .ZN(n4400) );
  AND2_X1 U5945 ( .A1(n9542), .A2(n9112), .ZN(n4401) );
  AND2_X1 U5946 ( .A1(n4752), .A2(n4754), .ZN(n4402) );
  AND2_X1 U5947 ( .A1(n6501), .A2(n6502), .ZN(n4403) );
  NAND2_X1 U5948 ( .A1(n9452), .A2(n9471), .ZN(n4404) );
  INV_X1 U5949 ( .A(n4693), .ZN(n4691) );
  NAND2_X1 U5950 ( .A1(n9993), .A2(n7879), .ZN(n4693) );
  OR2_X1 U5951 ( .A1(n6369), .A2(n6317), .ZN(n4405) );
  NAND2_X1 U5952 ( .A1(n8053), .A2(n8024), .ZN(n4406) );
  INV_X1 U5953 ( .A(n4731), .ZN(n9254) );
  NAND2_X1 U5954 ( .A1(n9160), .A2(n9144), .ZN(n4731) );
  OR2_X1 U5955 ( .A1(n4683), .A2(n4378), .ZN(n4680) );
  OR2_X1 U5956 ( .A1(n5885), .A2(n4377), .ZN(n4407) );
  AND2_X1 U5957 ( .A1(n7109), .A2(n9019), .ZN(n4408) );
  AND2_X1 U5958 ( .A1(n4684), .A2(n4369), .ZN(n4409) );
  OR2_X1 U5959 ( .A1(n4959), .A2(n7321), .ZN(n4410) );
  AND2_X1 U5960 ( .A1(n4877), .A2(n4875), .ZN(n4411) );
  AND2_X1 U5961 ( .A1(n4690), .A2(n9915), .ZN(n4412) );
  INV_X1 U5962 ( .A(n9667), .ZN(n9596) );
  NAND2_X1 U5963 ( .A1(n5864), .A2(n5863), .ZN(n9667) );
  AND2_X1 U5964 ( .A1(n6299), .A2(n8637), .ZN(n4413) );
  AND2_X1 U5965 ( .A1(n4627), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4414) );
  AND2_X1 U5966 ( .A1(n5375), .A2(n5362), .ZN(n4415) );
  AND2_X1 U5967 ( .A1(n8515), .A2(n4449), .ZN(n4416) );
  AND2_X1 U5968 ( .A1(n9999), .A2(n4353), .ZN(n4417) );
  NAND2_X1 U5969 ( .A1(n9183), .A2(n4516), .ZN(n4418) );
  AND2_X1 U5970 ( .A1(n4852), .A2(n5636), .ZN(n4419) );
  AND2_X1 U5971 ( .A1(n4819), .A2(n4817), .ZN(n4420) );
  INV_X1 U5972 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5557) );
  INV_X1 U5973 ( .A(n4615), .ZN(n4614) );
  NAND2_X1 U5974 ( .A1(n8676), .A2(n4616), .ZN(n4615) );
  INV_X1 U5975 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4852) );
  XNOR2_X1 U5976 ( .A(n5351), .B(n5350), .ZN(n5543) );
  INV_X1 U5977 ( .A(n9155), .ZN(n4516) );
  AND2_X1 U5978 ( .A1(n5470), .A2(n4725), .ZN(n4421) );
  INV_X1 U5979 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n4708) );
  OR2_X1 U5980 ( .A1(n4972), .A2(SI_17_), .ZN(n4422) );
  XNOR2_X1 U5981 ( .A(n6156), .B(SI_29_), .ZN(n8879) );
  AND2_X1 U5982 ( .A1(n5322), .A2(n4801), .ZN(n4423) );
  OAI21_X1 U5983 ( .B1(n8005), .B2(n4601), .A(n4357), .ZN(n8110) );
  OAI21_X1 U5984 ( .B1(n5319), .B2(n4862), .A(n4860), .ZN(n8686) );
  INV_X1 U5985 ( .A(n8144), .ZN(n8360) );
  NAND2_X1 U5986 ( .A1(n8926), .A2(n6521), .ZN(n8934) );
  NAND2_X1 U5987 ( .A1(n5319), .A2(n5318), .ZN(n8697) );
  NAND2_X1 U5988 ( .A1(n4797), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5349) );
  INV_X1 U5989 ( .A(n6287), .ZN(n4613) );
  AND2_X1 U5990 ( .A1(n8172), .A2(n8667), .ZN(n4424) );
  INV_X1 U5991 ( .A(n9278), .ZN(n7852) );
  NOR3_X1 U5992 ( .A1(n8010), .A2(n9657), .A3(n4575), .ZN(n4573) );
  AND2_X1 U5993 ( .A1(n8151), .A2(n8150), .ZN(n4425) );
  AND2_X1 U5994 ( .A1(n6547), .A2(n6548), .ZN(n4426) );
  NOR2_X1 U5995 ( .A1(n9551), .A2(n9652), .ZN(n9523) );
  INV_X1 U5996 ( .A(n4572), .ZN(n9482) );
  NOR2_X1 U5997 ( .A1(n8401), .A2(n8400), .ZN(n4427) );
  AND2_X1 U5998 ( .A1(n4815), .A2(n4813), .ZN(n4428) );
  INV_X1 U5999 ( .A(n4574), .ZN(n9566) );
  NOR2_X1 U6000 ( .A1(n8010), .A2(n4575), .ZN(n4574) );
  AND2_X1 U6001 ( .A1(n4837), .A2(n6509), .ZN(n4429) );
  INV_X1 U6002 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n4800) );
  OR2_X1 U6003 ( .A1(n6150), .A2(n8841), .ZN(n4430) );
  OR2_X1 U6004 ( .A1(n6150), .A2(n8774), .ZN(n4431) );
  AND2_X1 U6005 ( .A1(n6515), .A2(n6516), .ZN(n4432) );
  AND2_X1 U6006 ( .A1(n4977), .A2(n4362), .ZN(n4433) );
  AND2_X1 U6007 ( .A1(n4551), .A2(n4550), .ZN(n4434) );
  AND2_X1 U6008 ( .A1(n4636), .A2(n4635), .ZN(n4435) );
  INV_X1 U6009 ( .A(n5885), .ZN(n4663) );
  XNOR2_X1 U6010 ( .A(n5635), .B(n5634), .ZN(n6048) );
  OAI22_X1 U6011 ( .A1(n7519), .A2(n7518), .B1(n7512), .B2(n9930), .ZN(n7381)
         );
  XNOR2_X1 U6012 ( .A(n6017), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6395) );
  NAND2_X1 U6013 ( .A1(n8427), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4436) );
  AND2_X1 U6014 ( .A1(n9941), .A2(n4353), .ZN(n4437) );
  OAI211_X1 U6015 ( .C1(n6947), .C2(n4865), .A(n4866), .B(n5134), .ZN(n7610)
         );
  NAND2_X1 U6016 ( .A1(n4885), .A2(n6347), .ZN(n7523) );
  OR2_X1 U6017 ( .A1(n7813), .A2(n8382), .ZN(n4438) );
  AND2_X1 U6018 ( .A1(n9941), .A2(n9989), .ZN(n4439) );
  AND2_X1 U6019 ( .A1(n7736), .A2(n5194), .ZN(n4440) );
  OR2_X1 U6020 ( .A1(n7814), .A2(n7935), .ZN(n4441) );
  AND2_X1 U6021 ( .A1(n4787), .A2(n4788), .ZN(n4442) );
  AND2_X1 U6022 ( .A1(n4539), .A2(n4538), .ZN(n4443) );
  NAND2_X1 U6023 ( .A1(n8427), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4444) );
  OR2_X1 U6024 ( .A1(n7813), .A2(n7979), .ZN(n4445) );
  INV_X1 U6025 ( .A(n9389), .ZN(n4732) );
  NAND2_X1 U6026 ( .A1(n6046), .A2(n9262), .ZN(n9906) );
  INV_X1 U6027 ( .A(n9906), .ZN(n9934) );
  NAND2_X1 U6028 ( .A1(n5063), .A2(n5062), .ZN(n7046) );
  NAND2_X1 U6029 ( .A1(n5803), .A2(n5802), .ZN(n7882) );
  INV_X1 U6030 ( .A(n7882), .ZN(n4570) );
  AND2_X1 U6031 ( .A1(n6459), .A2(n6458), .ZN(n4446) );
  NOR2_X1 U6032 ( .A1(n4621), .A2(n4623), .ZN(n4447) );
  XOR2_X1 U6033 ( .A(n7464), .B(P2_REG2_REG_8__SCAN_IN), .Z(n4448) );
  INV_X1 U6034 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n4836) );
  INV_X1 U6035 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n4625) );
  XNOR2_X1 U6036 ( .A(n8457), .B(n8458), .ZN(n8428) );
  XNOR2_X1 U6037 ( .A(n8445), .B(n8458), .ZN(n8425) );
  AOI21_X1 U6038 ( .B1(n8506), .B2(n8505), .A(n8504), .ZN(n8507) );
  OAI21_X1 U6039 ( .B1(n8375), .B2(n8374), .A(n8373), .ZN(n8381) );
  NAND2_X1 U6040 ( .A1(n7659), .A2(n7660), .ZN(n7710) );
  NOR2_X1 U6041 ( .A1(n7408), .A2(n6994), .ZN(n6996) );
  NOR2_X1 U6042 ( .A1(n8451), .A2(n8450), .ZN(n8474) );
  NOR2_X1 U6043 ( .A1(n8414), .A2(n8413), .ZN(n8415) );
  NOR2_X1 U6044 ( .A1(n8435), .A2(n8434), .ZN(n8436) );
  OAI21_X1 U6045 ( .B1(n7657), .B2(n7658), .A(n7656), .ZN(n7659) );
  NAND2_X1 U6046 ( .A1(n4451), .A2(n10051), .ZN(n8514) );
  INV_X1 U6047 ( .A(n8511), .ZN(n4451) );
  INV_X1 U6048 ( .A(n5202), .ZN(n4818) );
  MUX2_X1 U6049 ( .A(n6279), .B(n6278), .S(n6322), .Z(n6288) );
  AOI21_X2 U6050 ( .B1(n4453), .B2(n4452), .A(n4405), .ZN(n6320) );
  INV_X1 U6051 ( .A(n6327), .ZN(n6334) );
  AOI21_X1 U6052 ( .B1(n8197), .B2(n6328), .A(n6330), .ZN(n6326) );
  AOI211_X1 U6053 ( .C1(n6299), .C2(n6298), .A(n6297), .B(n6296), .ZN(n6300)
         );
  AOI21_X1 U6054 ( .B1(n4456), .B2(n6469), .A(n7831), .ZN(n6472) );
  XNOR2_X1 U6055 ( .A(n7830), .B(n4456), .ZN(n7676) );
  NOR2_X1 U6056 ( .A1(n4458), .A2(n6471), .ZN(n4457) );
  OAI21_X1 U6057 ( .B1(n6515), .B2(n4471), .A(n4825), .ZN(n4470) );
  OAI21_X2 U6058 ( .B1(n4469), .B2(n4470), .A(n4823), .ZN(n6534) );
  NAND2_X1 U6059 ( .A1(n8995), .A2(n6516), .ZN(n8925) );
  INV_X1 U6060 ( .A(n4844), .ZN(n4480) );
  INV_X1 U6061 ( .A(n6473), .ZN(n4850) );
  NAND2_X1 U6062 ( .A1(n8901), .A2(n4361), .ZN(n4483) );
  OAI21_X1 U6063 ( .B1(n5162), .B2(n4371), .A(n5173), .ZN(n4490) );
  NAND2_X1 U6064 ( .A1(n4942), .A2(n4492), .ZN(n4491) );
  INV_X1 U6065 ( .A(n5162), .ZN(n4494) );
  OAI21_X2 U6066 ( .B1(n4942), .B2(n4494), .A(n4495), .ZN(n5174) );
  AND2_X1 U6067 ( .A1(n5653), .A2(n5652), .ZN(n4496) );
  NAND2_X1 U6068 ( .A1(n6417), .A2(n6415), .ZN(n6413) );
  OAI211_X1 U6069 ( .C1(n6712), .C2(n4498), .A(n4497), .B(n9209), .ZN(n6025)
         );
  NAND2_X1 U6070 ( .A1(n6848), .A2(n6023), .ZN(n4497) );
  INV_X1 U6071 ( .A(n6023), .ZN(n4498) );
  NAND2_X1 U6072 ( .A1(n6845), .A2(n6023), .ZN(n7075) );
  NAND2_X1 U6073 ( .A1(n4499), .A2(n6712), .ZN(n6845) );
  NAND2_X1 U6074 ( .A1(n9122), .A2(n4509), .ZN(n4508) );
  OR2_X1 U6075 ( .A1(n9169), .A2(n4516), .ZN(n4513) );
  NAND3_X1 U6076 ( .A1(n4503), .A2(n4512), .A3(n9498), .ZN(n4511) );
  NAND2_X1 U6077 ( .A1(n9212), .A2(n9048), .ZN(n9047) );
  NAND2_X1 U6078 ( .A1(n7062), .A2(n9215), .ZN(n9212) );
  AND2_X1 U6079 ( .A1(n6028), .A2(n9208), .ZN(n7062) );
  INV_X1 U6080 ( .A(n6069), .ZN(n5616) );
  NAND2_X1 U6081 ( .A1(n5616), .A2(n4851), .ZN(n5621) );
  NAND3_X1 U6082 ( .A1(n9086), .A2(n9155), .A3(n9085), .ZN(n4528) );
  NAND2_X1 U6083 ( .A1(n4531), .A2(n7018), .ZN(n7489) );
  INV_X1 U6084 ( .A(n4531), .ZN(n4530) );
  NAND2_X1 U6085 ( .A1(n8405), .A2(n4533), .ZN(n4532) );
  NAND3_X1 U6086 ( .A1(n4713), .A2(n4710), .A3(n7451), .ZN(n4540) );
  NAND2_X1 U6087 ( .A1(n4713), .A2(n7451), .ZN(n4538) );
  NAND2_X1 U6088 ( .A1(n4541), .A2(n4540), .ZN(n7810) );
  INV_X1 U6089 ( .A(n4551), .ZN(n7811) );
  INV_X1 U6090 ( .A(n7812), .ZN(n4550) );
  NOR2_X1 U6091 ( .A1(n8497), .A2(n8498), .ZN(n8501) );
  OAI21_X1 U6092 ( .B1(n8482), .B2(n4553), .A(n4552), .ZN(n8527) );
  INV_X1 U6093 ( .A(n8500), .ZN(n4554) );
  XNOR2_X1 U6094 ( .A(n8496), .B(n8505), .ZN(n8482) );
  NAND2_X1 U6095 ( .A1(n6039), .A2(n4558), .ZN(n4557) );
  NAND2_X1 U6096 ( .A1(n4694), .A2(n4564), .ZN(n4563) );
  NAND2_X1 U6097 ( .A1(n9908), .A2(n4568), .ZN(n4567) );
  OAI211_X1 U6098 ( .C1(n6045), .C2(n9934), .A(n4569), .B(n9417), .ZN(n9610)
         );
  NOR2_X1 U6099 ( .A1(n7084), .A2(n8896), .ZN(n7067) );
  NOR2_X2 U6100 ( .A1(n9482), .A2(n9626), .ZN(n9461) );
  NOR2_X2 U6101 ( .A1(n9524), .A2(n9513), .ZN(n9512) );
  INV_X1 U6102 ( .A(n4573), .ZN(n9551) );
  NOR2_X2 U6103 ( .A1(n9449), .A2(n9616), .ZN(n9418) );
  NAND2_X1 U6104 ( .A1(n4593), .A2(n4591), .ZN(n8569) );
  NOR2_X1 U6105 ( .A1(n6181), .A2(n6182), .ZN(n4589) );
  NAND2_X1 U6106 ( .A1(n8357), .A2(n8801), .ZN(n4590) );
  NAND2_X1 U6107 ( .A1(n4598), .A2(n6213), .ZN(n4597) );
  NAND2_X1 U6108 ( .A1(n4595), .A2(n4594), .ZN(n7688) );
  INV_X1 U6109 ( .A(n6207), .ZN(n4598) );
  AND2_X1 U6110 ( .A1(n6213), .A2(n6207), .ZN(n6946) );
  NAND2_X1 U6111 ( .A1(n8005), .A2(n4357), .ZN(n4600) );
  NAND2_X1 U6112 ( .A1(n5532), .A2(n4602), .ZN(n7930) );
  NAND2_X1 U6113 ( .A1(n7930), .A2(n6243), .ZN(n5534) );
  NAND2_X1 U6114 ( .A1(n4604), .A2(n4786), .ZN(n5202) );
  AOI21_X1 U6115 ( .B1(n8634), .B2(n4413), .A(n4607), .ZN(n8599) );
  OAI21_X1 U6116 ( .B1(n8685), .B2(n4615), .A(n4612), .ZN(n8661) );
  OAI21_X1 U6117 ( .B1(n8685), .B2(n6343), .A(n6341), .ZN(n8675) );
  NAND2_X1 U6118 ( .A1(n6343), .A2(n6341), .ZN(n4616) );
  NAND2_X1 U6119 ( .A1(n5529), .A2(n6228), .ZN(n7735) );
  NAND2_X1 U6120 ( .A1(n4617), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5046) );
  NAND3_X1 U6121 ( .A1(n4898), .A2(n5211), .A3(n4618), .ZN(n4617) );
  NAND3_X1 U6122 ( .A1(n4898), .A2(n5211), .A3(n5044), .ZN(n8873) );
  NAND2_X1 U6123 ( .A1(n7430), .A2(n4414), .ZN(n4622) );
  INV_X1 U6124 ( .A(n4622), .ZN(n4621) );
  INV_X1 U6125 ( .A(n4624), .ZN(n7008) );
  INV_X1 U6126 ( .A(n7412), .ZN(n4627) );
  OAI21_X1 U6127 ( .B1(n8398), .B2(n4628), .A(n4630), .ZN(n8445) );
  OR2_X1 U6128 ( .A1(n4638), .A2(n7650), .ZN(n7457) );
  INV_X1 U6129 ( .A(n4640), .ZN(n4638) );
  NAND2_X1 U6130 ( .A1(n8494), .A2(n4643), .ZN(n4641) );
  INV_X1 U6131 ( .A(n7089), .ZN(n9965) );
  NAND2_X2 U6132 ( .A1(n5675), .A2(n6669), .ZN(n5673) );
  NAND3_X1 U6133 ( .A1(n5707), .A2(n4646), .A3(n5672), .ZN(n5739) );
  NAND4_X1 U6134 ( .A1(n5707), .A2(n4646), .A3(n5672), .A4(n5604), .ZN(n5741)
         );
  NOR2_X2 U6135 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n5707) );
  NAND2_X1 U6136 ( .A1(n6894), .A2(n4408), .ZN(n4664) );
  OAI21_X1 U6137 ( .B1(n9489), .B2(n4672), .A(n4669), .ZN(n4668) );
  AOI21_X1 U6138 ( .B1(n7381), .B2(n4412), .A(n4686), .ZN(n7770) );
  NOR2_X2 U6139 ( .A1(n5202), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5211) );
  NOR2_X1 U6140 ( .A1(n5614), .A2(n5613), .ZN(n5615) );
  INV_X1 U6141 ( .A(n7044), .ZN(n7043) );
  NAND2_X2 U6142 ( .A1(n6961), .A2(n5000), .ZN(n5111) );
  NAND2_X1 U6143 ( .A1(n4695), .A2(n9222), .ZN(n7382) );
  NAND2_X1 U6144 ( .A1(n4702), .A2(n4701), .ZN(n9443) );
  NOR2_X4 U6145 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6961) );
  NAND2_X1 U6146 ( .A1(n6961), .A2(n5090), .ZN(n5109) );
  NAND2_X2 U6147 ( .A1(n4718), .A2(n4716), .ZN(n4928) );
  NAND3_X1 U6148 ( .A1(n4717), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4716) );
  NAND3_X1 U6149 ( .A1(n9386), .A2(n4720), .A3(n4719), .ZN(n4718) );
  NAND2_X1 U6150 ( .A1(n5430), .A2(n4421), .ZN(n4724) );
  NAND2_X1 U6151 ( .A1(n5430), .A2(n5429), .ZN(n5464) );
  INV_X1 U6152 ( .A(n9393), .ZN(n9691) );
  NAND2_X1 U6153 ( .A1(n4733), .A2(n4735), .ZN(n4956) );
  NAND2_X1 U6154 ( .A1(n5174), .A2(n4737), .ZN(n4733) );
  NAND2_X1 U6155 ( .A1(n4747), .A2(n4745), .ZN(n4968) );
  INV_X1 U6156 ( .A(n5270), .ZN(n4744) );
  NAND2_X1 U6157 ( .A1(n5303), .A2(n4433), .ZN(n4751) );
  OR2_X1 U6158 ( .A1(n5303), .A2(n4971), .ZN(n4756) );
  OAI21_X1 U6159 ( .B1(n5209), .B2(n4775), .A(n4958), .ZN(n5226) );
  XNOR2_X1 U6160 ( .A(n6907), .B(n7630), .ZN(n6918) );
  NAND2_X1 U6161 ( .A1(n8187), .A2(n4780), .ZN(n4776) );
  NAND2_X1 U6162 ( .A1(n4776), .A2(n4777), .ZN(n8193) );
  NAND2_X1 U6163 ( .A1(n5323), .A2(n4798), .ZN(n4796) );
  INV_X1 U6164 ( .A(n7362), .ZN(n4804) );
  AOI21_X1 U6165 ( .B1(n4804), .B2(n4803), .A(n7580), .ZN(n4802) );
  NAND2_X1 U6166 ( .A1(n4806), .A2(n7579), .ZN(n4805) );
  INV_X1 U6167 ( .A(n4809), .ZN(n7532) );
  OAI21_X1 U6168 ( .B1(n8145), .B2(n4812), .A(n4810), .ZN(n8260) );
  NAND2_X2 U6169 ( .A1(n8168), .A2(n8231), .ZN(n8301) );
  NAND2_X1 U6170 ( .A1(n4818), .A2(n4819), .ZN(n5244) );
  NAND2_X1 U6171 ( .A1(n4818), .A2(n4420), .ZN(n5258) );
  NAND2_X1 U6172 ( .A1(n8946), .A2(n6574), .ZN(n8916) );
  AND2_X1 U6173 ( .A1(n4918), .A2(n4835), .ZN(n5658) );
  NAND2_X1 U6174 ( .A1(n4838), .A2(n6509), .ZN(n6514) );
  NOR2_X1 U6175 ( .A1(n7033), .A2(n4359), .ZN(n7134) );
  OAI21_X1 U6176 ( .B1(n8996), .B2(n4432), .A(n8995), .ZN(n8998) );
  NAND2_X1 U6177 ( .A1(n5616), .A2(n4915), .ZN(n6072) );
  NAND2_X1 U6178 ( .A1(n4853), .A2(n5609), .ZN(n5873) );
  NAND2_X1 U6179 ( .A1(n5319), .A2(n4858), .ZN(n4857) );
  INV_X1 U6180 ( .A(n5118), .ZN(n4863) );
  NAND2_X1 U6181 ( .A1(n4863), .A2(n5133), .ZN(n4865) );
  OAI21_X1 U6182 ( .B1(n6947), .B2(n5118), .A(n5117), .ZN(n7692) );
  NAND2_X1 U6183 ( .A1(n5179), .A2(n6347), .ZN(n4881) );
  NAND2_X1 U6184 ( .A1(n7547), .A2(n4883), .ZN(n4882) );
  NAND2_X1 U6185 ( .A1(n4882), .A2(n4880), .ZN(n7738) );
  OAI21_X1 U6186 ( .B1(n7736), .B2(n4888), .A(n4886), .ZN(n7933) );
  NAND2_X1 U6187 ( .A1(n4891), .A2(n4415), .ZN(n8650) );
  NOR2_X2 U6188 ( .A1(n4893), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n4892) );
  NAND2_X1 U6189 ( .A1(n6848), .A2(n6842), .ZN(n6841) );
  OR2_X1 U6190 ( .A1(n7083), .A2(n7089), .ZN(n7084) );
  INV_X1 U6191 ( .A(n6405), .ZN(n6713) );
  NAND2_X1 U6192 ( .A1(n6189), .A2(n6188), .ZN(n6190) );
  NAND2_X1 U6193 ( .A1(n6186), .A2(n6185), .ZN(n6191) );
  NAND2_X1 U6194 ( .A1(n5543), .A2(n7687), .ZN(n6903) );
  NAND2_X1 U6195 ( .A1(n5553), .A2(n8129), .ZN(n5562) );
  NAND2_X1 U6196 ( .A1(n5562), .A2(n5563), .ZN(n6782) );
  AOI21_X1 U6197 ( .B1(n5555), .B2(n5549), .A(n4903), .ZN(n5551) );
  NAND2_X1 U6198 ( .A1(n6879), .A2(n6782), .ZN(n6818) );
  OR2_X1 U6199 ( .A1(n6782), .A2(n5577), .ZN(n6141) );
  OR2_X1 U6200 ( .A1(n6782), .A2(P2_D_REG_1__SCAN_IN), .ZN(n5564) );
  OAI21_X1 U6201 ( .B1(n8599), .B2(n6306), .A(n6305), .ZN(n8592) );
  XNOR2_X1 U6202 ( .A(n6906), .B(n7905), .ZN(n6907) );
  NAND2_X1 U6203 ( .A1(n8891), .A2(n6439), .ZN(n6650) );
  NOR2_X1 U6204 ( .A1(n5666), .A2(n5665), .ZN(n6405) );
  OAI22_X1 U6205 ( .A1(n6405), .A2(n6551), .B1(n6404), .B2(n6813), .ZN(n6411)
         );
  NAND2_X2 U6206 ( .A1(n6048), .A2(n8108), .ZN(n5675) );
  NAND2_X1 U6207 ( .A1(n5626), .A2(n8130), .ZN(n5701) );
  INV_X1 U6208 ( .A(n5626), .ZN(n5624) );
  NOR2_X2 U6209 ( .A1(n7034), .A2(n7035), .ZN(n7033) );
  OR2_X1 U6210 ( .A1(n6149), .A2(n10091), .ZN(n5589) );
  NAND2_X1 U6211 ( .A1(n8639), .A2(n5398), .ZN(n8627) );
  OR2_X1 U6212 ( .A1(n5095), .A2(n6672), .ZN(n5098) );
  OR2_X1 U6213 ( .A1(n5095), .A2(n6684), .ZN(n5077) );
  INV_X2 U6214 ( .A(n5095), .ZN(n6175) );
  OR2_X1 U6215 ( .A1(n6905), .A2(n6145), .ZN(n7372) );
  OR2_X1 U6216 ( .A1(n5096), .A2(n6664), .ZN(n5097) );
  OAI22_X1 U6217 ( .A1(n8575), .A2(n5457), .B1(n8589), .B2(n8805), .ZN(n8562)
         );
  OR2_X1 U6218 ( .A1(n4411), .A2(n8602), .ZN(n8603) );
  NOR2_X2 U6219 ( .A1(n6650), .A2(n6651), .ZN(n6649) );
  NOR3_X2 U6220 ( .A1(n6649), .A2(n6451), .A3(n6450), .ZN(n6930) );
  INV_X1 U6221 ( .A(n9229), .ZN(n6036) );
  OAI21_X1 U6222 ( .B1(n8112), .B2(n5285), .A(n5284), .ZN(n8724) );
  OR2_X1 U6223 ( .A1(n6061), .A2(n9008), .ZN(n4899) );
  INV_X1 U6224 ( .A(n9709), .ZN(n6137) );
  INV_X1 U6225 ( .A(n9645), .ZN(n6101) );
  INV_X1 U6226 ( .A(n9418), .ZN(n9428) );
  AND2_X1 U6227 ( .A1(n8747), .A2(n8794), .ZN(n4900) );
  AND2_X1 U6228 ( .A1(n4431), .A2(n6151), .ZN(n4901) );
  OR2_X1 U6229 ( .A1(n10088), .A2(n5588), .ZN(n4902) );
  NOR2_X1 U6230 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4903) );
  INV_X1 U6231 ( .A(n9236), .ZN(n6038) );
  OR2_X1 U6232 ( .A1(n9596), .A2(n8939), .ZN(n4904) );
  NAND2_X1 U6233 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), 
        .ZN(n4905) );
  AND2_X1 U6234 ( .A1(n4430), .A2(n4902), .ZN(n4906) );
  OR2_X1 U6235 ( .A1(n4985), .A2(n4984), .ZN(n4907) );
  AND2_X1 U6236 ( .A1(n6319), .A2(n6318), .ZN(n4909) );
  XNOR2_X1 U6237 ( .A(n4925), .B(n4924), .ZN(n5072) );
  OR2_X1 U6238 ( .A1(n6629), .A2(n7913), .ZN(n4910) );
  AND3_X1 U6239 ( .A1(n6010), .A2(n6009), .A3(n6008), .ZN(n4911) );
  NOR2_X1 U6240 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n4912) );
  AND2_X1 U6241 ( .A1(n5620), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4913) );
  INV_X1 U6242 ( .A(n6395), .ZN(n6397) );
  INV_X1 U6243 ( .A(P2_U3893), .ZN(n8359) );
  NAND2_X1 U6244 ( .A1(n6200), .A2(n6199), .ZN(n6197) );
  INV_X1 U6245 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5030) );
  OR2_X1 U6246 ( .A1(n9576), .A2(n6895), .ZN(n9955) );
  INV_X1 U6247 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4923) );
  AND2_X1 U6248 ( .A1(n4955), .A2(n4954), .ZN(n4914) );
  INV_X1 U6249 ( .A(n9116), .ZN(n6040) );
  NAND2_X1 U6250 ( .A1(n9198), .A2(n4351), .ZN(n7914) );
  INV_X1 U6251 ( .A(n7914), .ZN(n7513) );
  INV_X1 U6252 ( .A(n6956), .ZN(n6959) );
  INV_X1 U6253 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5028) );
  INV_X1 U6254 ( .A(n9402), .ZN(n6109) );
  CLKBUF_X1 U6255 ( .A(n6665), .Z(n8878) );
  AND2_X1 U6256 ( .A1(n5587), .A2(n5586), .ZN(n10091) );
  INV_X1 U6257 ( .A(n9416), .ZN(n6110) );
  INV_X1 U6258 ( .A(n5684), .ZN(n5913) );
  AND2_X1 U6259 ( .A1(n7941), .A2(n6096), .ZN(n9155) );
  NOR2_X1 U6260 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n4915) );
  INV_X1 U6261 ( .A(n7598), .ZN(n5756) );
  INV_X1 U6262 ( .A(n6350), .ZN(n5179) );
  INV_X2 U6263 ( .A(n8066), .ZN(n8786) );
  INV_X1 U6264 ( .A(n5701), .ZN(n5918) );
  XOR2_X1 U6265 ( .A(n8524), .B(n8530), .Z(n4917) );
  INV_X1 U6266 ( .A(n7813), .ZN(n8388) );
  OR2_X1 U6267 ( .A1(n5675), .A2(n6753), .ZN(n4918) );
  OR2_X1 U6268 ( .A1(n8848), .A2(n8689), .ZN(n4919) );
  INV_X1 U6269 ( .A(n8363), .ZN(n8024) );
  INV_X1 U6270 ( .A(n8664), .ZN(n5375) );
  INV_X1 U6271 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5003) );
  INV_X1 U6272 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5612) );
  NAND2_X1 U6273 ( .A1(n8025), .A2(n8024), .ZN(n8026) );
  NAND2_X1 U6274 ( .A1(n6332), .A2(n6331), .ZN(n6333) );
  INV_X1 U6275 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8382) );
  INV_X1 U6276 ( .A(n6018), .ZN(n6012) );
  INV_X1 U6277 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n4950) );
  INV_X1 U6278 ( .A(n8028), .ZN(n5533) );
  INV_X1 U6279 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5554) );
  NAND2_X1 U6280 ( .A1(n6519), .A2(n6520), .ZN(n6521) );
  INV_X1 U6281 ( .A(n5791), .ZN(n5594) );
  INV_X1 U6282 ( .A(n5960), .ZN(n5601) );
  INV_X1 U6283 ( .A(n9435), .ZN(n6629) );
  AND2_X1 U6284 ( .A1(n9067), .A2(n9925), .ZN(n9052) );
  AND2_X1 U6285 ( .A1(n5462), .A2(n5465), .ZN(n5463) );
  INV_X1 U6286 ( .A(SI_24_), .ZN(n7308) );
  INV_X1 U6287 ( .A(SI_19_), .ZN(n7260) );
  INV_X1 U6288 ( .A(SI_16_), .ZN(n7329) );
  INV_X1 U6289 ( .A(SI_8_), .ZN(n7180) );
  INV_X1 U6290 ( .A(n7358), .ZN(n8163) );
  OR2_X1 U6291 ( .A1(n5474), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5490) );
  INV_X1 U6292 ( .A(n5082), .ZN(n5120) );
  NOR2_X1 U6293 ( .A1(n10026), .A2(n10025), .ZN(n10024) );
  INV_X1 U6294 ( .A(n8396), .ZN(n8397) );
  NOR2_X1 U6295 ( .A1(n5020), .A2(n5017), .ZN(n5018) );
  INV_X1 U6296 ( .A(n5383), .ZN(n5039) );
  OR2_X1 U6297 ( .A1(n5218), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5230) );
  AND2_X1 U6298 ( .A1(n6875), .A2(n8745), .ZN(n7376) );
  OR2_X1 U6299 ( .A1(n6872), .A2(n6390), .ZN(n6876) );
  INV_X1 U6300 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5497) );
  INV_X1 U6301 ( .A(n5850), .ZN(n5595) );
  AND2_X1 U6302 ( .A1(n6607), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n6408) );
  INV_X1 U6303 ( .A(n6553), .ZN(n6554) );
  OR2_X1 U6304 ( .A1(n5975), .A2(n5602), .ZN(n5987) );
  NAND2_X1 U6305 ( .A1(n5687), .A2(n5686), .ZN(n5688) );
  OR2_X1 U6306 ( .A1(n9909), .A2(n6499), .ZN(n5840) );
  NAND2_X1 U6307 ( .A1(n7077), .A2(n8896), .ZN(n6026) );
  INV_X1 U6308 ( .A(n6608), .ZN(n9198) );
  INV_X1 U6309 ( .A(SI_26_), .ZN(n7337) );
  NAND2_X1 U6310 ( .A1(n4995), .A2(n4994), .ZN(n5413) );
  INV_X1 U6311 ( .A(SI_17_), .ZN(n7292) );
  INV_X1 U6312 ( .A(n5088), .ZN(n5188) );
  INV_X1 U6313 ( .A(n8678), .ZN(n8246) );
  INV_X1 U6314 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5026) );
  NAND2_X1 U6315 ( .A1(n10042), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n10041) );
  INV_X1 U6316 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5044) );
  OR2_X1 U6317 ( .A1(n6970), .A2(n8106), .ZN(n7127) );
  OR2_X1 U6318 ( .A1(n5433), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5449) );
  NAND2_X1 U6319 ( .A1(n5039), .A2(n5038), .ZN(n5392) );
  OR2_X1 U6320 ( .A1(n7967), .A2(n8052), .ZN(n6354) );
  NAND2_X1 U6321 ( .A1(n5531), .A2(n6351), .ZN(n5532) );
  INV_X1 U6322 ( .A(n7046), .ZN(n6920) );
  OAI21_X1 U6323 ( .B1(n8706), .B2(n5538), .A(n6266), .ZN(n8696) );
  INV_X1 U6324 ( .A(n8669), .ZN(n8726) );
  AND2_X1 U6325 ( .A1(n6345), .A2(n6344), .ZN(n8004) );
  AND2_X1 U6326 ( .A1(n7545), .A2(n6215), .ZN(n7612) );
  INV_X1 U6327 ( .A(n7375), .ZN(n7730) );
  NAND2_X1 U6328 ( .A1(n5595), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5852) );
  NAND2_X1 U6329 ( .A1(n5597), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5895) );
  NAND2_X1 U6330 ( .A1(n5759), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5791) );
  AND2_X1 U6331 ( .A1(n5987), .A2(n5603), .ZN(n9429) );
  OR2_X1 U6332 ( .A1(n5916), .A2(n8957), .ZN(n5925) );
  OR2_X1 U6333 ( .A1(n9792), .A2(n9788), .ZN(n9851) );
  INV_X1 U6334 ( .A(n9590), .ZN(n9942) );
  NAND2_X1 U6335 ( .A1(n9416), .A2(n9932), .ZN(n6126) );
  NAND2_X1 U6336 ( .A1(n9523), .A2(n9529), .ZN(n9524) );
  INV_X1 U6337 ( .A(n9523), .ZN(n9538) );
  AND2_X1 U6338 ( .A1(n9662), .A2(n9586), .ZN(n5885) );
  OR2_X1 U6339 ( .A1(n5820), .A2(n5819), .ZN(n5833) );
  OR2_X1 U6340 ( .A1(n6717), .A2(n9260), .ZN(n6621) );
  OR2_X1 U6341 ( .A1(n6717), .A2(n6063), .ZN(n9590) );
  OR2_X1 U6342 ( .A1(n6717), .A2(n6100), .ZN(n10004) );
  OR2_X1 U6343 ( .A1(n6811), .A2(n6607), .ZN(n6688) );
  NAND2_X1 U6344 ( .A1(n6011), .A2(n4911), .ZN(n6018) );
  INV_X1 U6345 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5800) );
  XNOR2_X1 U6346 ( .A(n8177), .B(n8178), .ZN(n8224) );
  OR2_X1 U6347 ( .A1(n5180), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5195) );
  AND2_X1 U6348 ( .A1(n8344), .A2(n8261), .ZN(n8275) );
  INV_X1 U6349 ( .A(n8347), .ZN(n8327) );
  AND2_X1 U6350 ( .A1(n6168), .A2(n5517), .ZN(n6184) );
  AND3_X1 U6351 ( .A1(n5408), .A2(n5407), .A3(n5406), .ZN(n8312) );
  AND4_X1 U6352 ( .A1(n5332), .A2(n5331), .A3(n5330), .A4(n5329), .ZN(n8712)
         );
  AND4_X1 U6353 ( .A1(n5266), .A2(n5265), .A3(n5264), .A4(n5263), .ZN(n8144)
         );
  NOR2_X1 U6354 ( .A1(n7653), .A2(n7652), .ZN(n7705) );
  INV_X1 U6355 ( .A(n8542), .ZN(n10051) );
  INV_X1 U6356 ( .A(n7975), .ZN(n7973) );
  INV_X1 U6357 ( .A(n8738), .ZN(n8596) );
  INV_X1 U6358 ( .A(n10064), .ZN(n8719) );
  AND2_X1 U6359 ( .A1(n7892), .A2(n7899), .ZN(n8118) );
  INV_X1 U6360 ( .A(n8774), .ZN(n8788) );
  INV_X1 U6361 ( .A(n8118), .ZN(n8794) );
  INV_X1 U6362 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5212) );
  INV_X1 U6363 ( .A(n9001), .ZN(n8984) );
  AND2_X1 U6364 ( .A1(n6613), .A2(n6620), .ZN(n8997) );
  INV_X1 U6365 ( .A(n9899), .ZN(n9882) );
  INV_X1 U6366 ( .A(n9125), .ZN(n9468) );
  INV_X1 U6367 ( .A(n9955), .ZN(n9939) );
  INV_X1 U6368 ( .A(n9601), .ZN(n9959) );
  INV_X1 U6369 ( .A(n10007), .ZN(n9675) );
  NAND2_X1 U6370 ( .A1(n7910), .A2(n9979), .ZN(n10007) );
  NAND2_X1 U6371 ( .A1(n6083), .A2(n6097), .ZN(n9718) );
  INV_X1 U6372 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6019) );
  AND2_X1 U6373 ( .A1(n5828), .A2(n5816), .ZN(n9366) );
  OR3_X1 U6374 ( .A1(n8129), .A2(n8202), .A3(n8069), .ZN(n6866) );
  INV_X1 U6375 ( .A(n8335), .ZN(n8348) );
  INV_X1 U6376 ( .A(n8339), .ZN(n8354) );
  NAND2_X1 U6377 ( .A1(n5456), .A2(n5455), .ZN(n8358) );
  INV_X1 U6378 ( .A(n10047), .ZN(n10023) );
  INV_X1 U6379 ( .A(n10056), .ZN(n8486) );
  INV_X1 U6380 ( .A(n8735), .ZN(n8594) );
  INV_X1 U6381 ( .A(n10069), .ZN(n8734) );
  NAND2_X1 U6382 ( .A1(n7374), .A2(n10064), .ZN(n10069) );
  OR2_X1 U6383 ( .A1(n8755), .A2(n8118), .ZN(n8791) );
  NAND3_X1 U6384 ( .A1(n6148), .A2(n7371), .A3(n6147), .ZN(n8066) );
  NAND2_X1 U6385 ( .A1(n10088), .A2(n8793), .ZN(n8841) );
  NAND2_X1 U6386 ( .A1(n10088), .A2(n8794), .ZN(n8870) );
  INV_X2 U6387 ( .A(n10091), .ZN(n10088) );
  AND2_X1 U6388 ( .A1(n6865), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6788) );
  INV_X1 U6389 ( .A(n6392), .ZN(n7944) );
  INV_X1 U6390 ( .A(n8417), .ZN(n8427) );
  INV_X1 U6391 ( .A(n8876), .ZN(n8880) );
  INV_X1 U6392 ( .A(n9914), .ZN(n9999) );
  INV_X1 U6393 ( .A(n6499), .ZN(n10005) );
  INV_X1 U6394 ( .A(n8997), .ZN(n8974) );
  AND2_X1 U6395 ( .A1(n6617), .A2(n9515), .ZN(n9008) );
  NAND2_X1 U6396 ( .A1(n6005), .A2(n6004), .ZN(n9416) );
  INV_X1 U6397 ( .A(n9870), .ZN(n9905) );
  OR2_X1 U6398 ( .A1(n9576), .A2(n6096), .ZN(n9405) );
  AND2_X1 U6399 ( .A1(n6719), .A2(n9515), .ZN(n9576) );
  INV_X1 U6400 ( .A(n9576), .ZN(n9598) );
  AND2_X2 U6401 ( .A1(n6104), .A2(n6611), .ZN(n10021) );
  NAND2_X1 U6402 ( .A1(n9402), .A2(n6137), .ZN(n6107) );
  INV_X1 U6403 ( .A(n10010), .ZN(n10009) );
  AND2_X2 U6404 ( .A1(n6104), .A2(n6708), .ZN(n10010) );
  INV_X1 U6405 ( .A(n6021), .ZN(n7941) );
  INV_X1 U6406 ( .A(n7948), .ZN(n9732) );
  INV_X1 U6407 ( .A(n9285), .ZN(P1_U3973) );
  AND2_X1 U6408 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4920) );
  NAND2_X1 U6409 ( .A1(n4928), .A2(n4920), .ZN(n5669) );
  AND2_X1 U6410 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4921) );
  NAND2_X1 U6411 ( .A1(n6663), .A2(n4921), .ZN(n5066) );
  NAND2_X1 U6412 ( .A1(n5669), .A2(n5066), .ZN(n5073) );
  OAI21_X1 U6413 ( .B1(n4928), .B2(n4923), .A(n4922), .ZN(n4925) );
  INV_X1 U6414 ( .A(SI_1_), .ZN(n4924) );
  NAND2_X1 U6415 ( .A1(n5073), .A2(n5072), .ZN(n4927) );
  NAND2_X1 U6416 ( .A1(n4925), .A2(SI_1_), .ZN(n4926) );
  NAND2_X1 U6417 ( .A1(n4927), .A2(n4926), .ZN(n5094) );
  MUX2_X1 U6418 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n4928), .Z(n4930) );
  INV_X1 U6419 ( .A(SI_2_), .ZN(n4929) );
  XNOR2_X1 U6420 ( .A(n4930), .B(n4929), .ZN(n5093) );
  NAND2_X1 U6421 ( .A1(n5094), .A2(n5093), .ZN(n4932) );
  NAND2_X1 U6422 ( .A1(n4930), .A2(SI_2_), .ZN(n4931) );
  NAND2_X1 U6423 ( .A1(n4932), .A2(n4931), .ZN(n5114) );
  MUX2_X1 U6424 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n4928), .Z(n4934) );
  INV_X1 U6425 ( .A(SI_3_), .ZN(n4933) );
  XNOR2_X1 U6426 ( .A(n4934), .B(n4933), .ZN(n5113) );
  NAND2_X1 U6427 ( .A1(n5114), .A2(n5113), .ZN(n4936) );
  NAND2_X1 U6428 ( .A1(n4934), .A2(SI_3_), .ZN(n4935) );
  NAND2_X1 U6429 ( .A1(n4936), .A2(n4935), .ZN(n5130) );
  MUX2_X1 U6430 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n4350), .Z(n4937) );
  INV_X1 U6431 ( .A(SI_4_), .ZN(n7249) );
  XNOR2_X1 U6432 ( .A(n4937), .B(n7249), .ZN(n5129) );
  NAND2_X1 U6433 ( .A1(n5130), .A2(n5129), .ZN(n4939) );
  NAND2_X1 U6434 ( .A1(n4937), .A2(SI_4_), .ZN(n4938) );
  NAND2_X1 U6435 ( .A1(n4939), .A2(n4938), .ZN(n5145) );
  MUX2_X1 U6436 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n4350), .Z(n4940) );
  INV_X1 U6437 ( .A(SI_5_), .ZN(n7190) );
  XNOR2_X1 U6438 ( .A(n4940), .B(n7190), .ZN(n5144) );
  NAND2_X1 U6439 ( .A1(n5145), .A2(n5144), .ZN(n4942) );
  NAND2_X1 U6440 ( .A1(n4940), .A2(SI_5_), .ZN(n4941) );
  MUX2_X1 U6441 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n4350), .Z(n4943) );
  INV_X1 U6442 ( .A(SI_6_), .ZN(n7187) );
  XNOR2_X1 U6443 ( .A(n4943), .B(n7187), .ZN(n5162) );
  MUX2_X1 U6444 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n4350), .Z(n4944) );
  XNOR2_X1 U6445 ( .A(n4944), .B(n7177), .ZN(n5173) );
  NAND2_X1 U6446 ( .A1(n4944), .A2(SI_7_), .ZN(n4945) );
  MUX2_X1 U6447 ( .A(n6691), .B(n6693), .S(n4350), .Z(n4946) );
  NAND2_X1 U6448 ( .A1(n4946), .A2(n7180), .ZN(n4949) );
  INV_X1 U6449 ( .A(n4946), .ZN(n4947) );
  NAND2_X1 U6450 ( .A1(n4947), .A2(SI_8_), .ZN(n4948) );
  NAND2_X1 U6451 ( .A1(n4949), .A2(n4948), .ZN(n5186) );
  MUX2_X1 U6452 ( .A(n6699), .B(n4950), .S(n4350), .Z(n4952) );
  INV_X1 U6453 ( .A(SI_9_), .ZN(n4951) );
  NAND2_X1 U6454 ( .A1(n4952), .A2(n4951), .ZN(n4955) );
  INV_X1 U6455 ( .A(n4952), .ZN(n4953) );
  NAND2_X1 U6456 ( .A1(n4953), .A2(SI_9_), .ZN(n4954) );
  MUX2_X1 U6457 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n4350), .Z(n4957) );
  NAND2_X1 U6458 ( .A1(n4957), .A2(SI_10_), .ZN(n4958) );
  MUX2_X1 U6459 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n4350), .Z(n5224) );
  INV_X1 U6460 ( .A(n5224), .ZN(n4959) );
  MUX2_X1 U6461 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n4350), .Z(n4960) );
  MUX2_X1 U6462 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n4350), .Z(n5255) );
  NAND2_X1 U6463 ( .A1(n5257), .A2(SI_13_), .ZN(n4962) );
  NAND2_X1 U6464 ( .A1(n4963), .A2(n4962), .ZN(n5270) );
  MUX2_X1 U6465 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n4350), .Z(n5268) );
  NAND2_X1 U6466 ( .A1(n4964), .A2(n7272), .ZN(n4965) );
  MUX2_X1 U6467 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n4350), .Z(n5287) );
  NOR2_X1 U6468 ( .A1(n5287), .A2(SI_15_), .ZN(n4966) );
  NAND2_X1 U6469 ( .A1(n5287), .A2(SI_15_), .ZN(n4967) );
  NAND2_X1 U6470 ( .A1(n4968), .A2(n4967), .ZN(n5303) );
  MUX2_X1 U6471 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n4350), .Z(n5301) );
  NOR2_X1 U6472 ( .A1(n4969), .A2(n7329), .ZN(n4971) );
  NAND2_X1 U6473 ( .A1(n4969), .A2(n7329), .ZN(n4970) );
  MUX2_X1 U6474 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n4350), .Z(n4972) );
  MUX2_X1 U6475 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4350), .Z(n4973) );
  NAND2_X1 U6476 ( .A1(n4973), .A2(SI_18_), .ZN(n4978) );
  INV_X1 U6477 ( .A(n4973), .ZN(n4975) );
  INV_X1 U6478 ( .A(SI_18_), .ZN(n4974) );
  NAND2_X1 U6479 ( .A1(n4975), .A2(n4974), .ZN(n4976) );
  NAND2_X1 U6480 ( .A1(n4978), .A2(n4976), .ZN(n5333) );
  INV_X1 U6481 ( .A(n5333), .ZN(n4977) );
  INV_X1 U6482 ( .A(n5347), .ZN(n4979) );
  MUX2_X1 U6483 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n4350), .Z(n4980) );
  XNOR2_X1 U6484 ( .A(n4980), .B(SI_19_), .ZN(n5346) );
  INV_X1 U6485 ( .A(n4980), .ZN(n4981) );
  NAND2_X1 U6486 ( .A1(n4981), .A2(n7260), .ZN(n4982) );
  INV_X1 U6487 ( .A(SI_20_), .ZN(n5363) );
  MUX2_X1 U6488 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n4350), .Z(n5364) );
  INV_X1 U6489 ( .A(n5378), .ZN(n4983) );
  MUX2_X1 U6490 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n4350), .Z(n5376) );
  INV_X1 U6491 ( .A(SI_21_), .ZN(n4984) );
  NAND2_X1 U6492 ( .A1(n4983), .A2(n4907), .ZN(n4987) );
  NAND2_X1 U6493 ( .A1(n4985), .A2(n4984), .ZN(n4986) );
  NAND2_X1 U6494 ( .A1(n4987), .A2(n4986), .ZN(n5389) );
  MUX2_X1 U6495 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n4350), .Z(n4988) );
  XNOR2_X1 U6496 ( .A(n4988), .B(n7189), .ZN(n5388) );
  NAND2_X1 U6497 ( .A1(n5389), .A2(n5388), .ZN(n4991) );
  INV_X1 U6498 ( .A(n4988), .ZN(n4989) );
  NAND2_X1 U6499 ( .A1(n4989), .A2(n7189), .ZN(n4990) );
  NAND2_X1 U6500 ( .A1(n4991), .A2(n4990), .ZN(n5400) );
  MUX2_X1 U6501 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .S(n4350), .Z(n4992) );
  XNOR2_X1 U6502 ( .A(n4992), .B(n7320), .ZN(n5399) );
  NAND2_X1 U6503 ( .A1(n5400), .A2(n5399), .ZN(n4995) );
  INV_X1 U6504 ( .A(n4992), .ZN(n4993) );
  NAND2_X1 U6505 ( .A1(n4993), .A2(n7320), .ZN(n4994) );
  MUX2_X1 U6506 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n4350), .Z(n4996) );
  XNOR2_X1 U6507 ( .A(n4996), .B(n7308), .ZN(n5412) );
  NAND2_X1 U6508 ( .A1(n5413), .A2(n5412), .ZN(n4999) );
  INV_X1 U6509 ( .A(n4996), .ZN(n4997) );
  NAND2_X1 U6510 ( .A1(n4997), .A2(n7308), .ZN(n4998) );
  NAND2_X1 U6511 ( .A1(n4999), .A2(n4998), .ZN(n5426) );
  MUX2_X1 U6512 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(P2_DATAO_REG_25__SCAN_IN), 
        .S(n4350), .Z(n5427) );
  XNOR2_X1 U6513 ( .A(n5427), .B(n7293), .ZN(n5425) );
  XNOR2_X1 U6514 ( .A(n5426), .B(n5425), .ZN(n7995) );
  NOR2_X1 U6515 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5006) );
  NOR2_X1 U6516 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5005) );
  NOR2_X1 U6517 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5004) );
  NAND4_X1 U6518 ( .A1(n5007), .A2(n5006), .A3(n5005), .A4(n5004), .ZN(n5015)
         );
  NOR2_X2 U6519 ( .A1(n5244), .A2(n5015), .ZN(n5498) );
  NOR2_X1 U6520 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5010) );
  NOR2_X1 U6521 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n5009) );
  NOR2_X1 U6522 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5008) );
  NAND4_X1 U6523 ( .A1(n5010), .A2(n5009), .A3(n5008), .A4(n5554), .ZN(n5014)
         );
  INV_X1 U6524 ( .A(n5014), .ZN(n5011) );
  NAND2_X1 U6525 ( .A1(n5498), .A2(n5011), .ZN(n5560) );
  NAND2_X1 U6526 ( .A1(n5019), .A2(n5018), .ZN(n5509) );
  INV_X1 U6527 ( .A(n4350), .ZN(n6669) );
  NAND2_X2 U6528 ( .A1(n5088), .A2(n6669), .ZN(n5095) );
  NAND2_X1 U6529 ( .A1(n7995), .A2(n6175), .ZN(n5023) );
  NAND2_X2 U6530 ( .A1(n5088), .A2(n4350), .ZN(n5096) );
  NAND2_X1 U6531 ( .A1(n5471), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5022) );
  NAND2_X1 U6532 ( .A1(n5025), .A2(n5024), .ZN(n5135) );
  INV_X1 U6533 ( .A(n5135), .ZN(n5027) );
  NAND2_X1 U6534 ( .A1(n5027), .A2(n5026), .ZN(n5151) );
  OR2_X2 U6535 ( .A1(n5230), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5248) );
  OR2_X2 U6536 ( .A1(n5312), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5327) );
  INV_X1 U6537 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5035) );
  OR2_X2 U6538 ( .A1(n5339), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5354) );
  INV_X1 U6539 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n7316) );
  INV_X1 U6540 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5038) );
  OR2_X2 U6541 ( .A1(n5403), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5416) );
  INV_X1 U6542 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5040) );
  INV_X1 U6543 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8252) );
  NAND2_X1 U6544 ( .A1(n5418), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5043) );
  NAND2_X1 U6545 ( .A1(n5433), .A2(n5043), .ZN(n8608) );
  XNOR2_X1 U6546 ( .A(n5046), .B(n5045), .ZN(n5048) );
  NAND2_X1 U6547 ( .A1(n8608), .A2(n5491), .ZN(n5055) );
  INV_X1 U6548 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n5052) );
  XNOR2_X2 U6549 ( .A(n5047), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5056) );
  NAND2_X4 U6550 ( .A1(n5057), .A2(n5056), .ZN(n5514) );
  INV_X2 U6551 ( .A(n5120), .ZN(n6162) );
  NAND2_X1 U6552 ( .A1(n6162), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5051) );
  NAND2_X1 U6553 ( .A1(n6161), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5050) );
  OAI211_X1 U6554 ( .C1(n5052), .C2(n5514), .A(n5051), .B(n5050), .ZN(n5053)
         );
  INV_X1 U6555 ( .A(n5053), .ZN(n5054) );
  NAND2_X1 U6556 ( .A1(n5082), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5061) );
  NAND2_X1 U6557 ( .A1(n5491), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5060) );
  INV_X1 U6558 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6960) );
  OR2_X1 U6559 ( .A1(n6960), .A2(n5056), .ZN(n5058) );
  OR2_X1 U6560 ( .A1(n5058), .A2(n5057), .ZN(n5059) );
  AND3_X1 U6561 ( .A1(n5061), .A2(n5060), .A3(n5059), .ZN(n5062) );
  NAND2_X1 U6562 ( .A1(n6663), .A2(SI_0_), .ZN(n5065) );
  INV_X1 U6563 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5064) );
  NAND2_X1 U6564 ( .A1(n5065), .A2(n5064), .ZN(n5067) );
  AND2_X1 U6565 ( .A1(n5067), .A2(n5066), .ZN(n8883) );
  MUX2_X1 U6566 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8883), .S(n5088), .Z(n7375) );
  INV_X1 U6567 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7573) );
  NAND2_X1 U6568 ( .A1(n5081), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5070) );
  NAND2_X1 U6569 ( .A1(n5491), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5069) );
  NAND2_X1 U6570 ( .A1(n5082), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5068) );
  OR2_X1 U6571 ( .A1(n5096), .A2(n4923), .ZN(n5078) );
  XNOR2_X1 U6572 ( .A(n5072), .B(n5073), .ZN(n6684) );
  NAND2_X1 U6573 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5074) );
  INV_X1 U6574 ( .A(n6961), .ZN(n5075) );
  NAND2_X1 U6575 ( .A1(n5188), .A2(n6959), .ZN(n5076) );
  AND3_X2 U6576 ( .A1(n5078), .A2(n5077), .A3(n5076), .ZN(n5523) );
  NAND2_X1 U6577 ( .A1(n7045), .A2(n7044), .ZN(n5080) );
  NAND2_X1 U6578 ( .A1(n7630), .A2(n7905), .ZN(n5079) );
  NAND2_X1 U6579 ( .A1(n5080), .A2(n5079), .ZN(n7628) );
  NAND2_X1 U6580 ( .A1(n5081), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5087) );
  NAND2_X1 U6581 ( .A1(n5082), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5086) );
  NAND2_X1 U6582 ( .A1(n5491), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5085) );
  INV_X1 U6583 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5083) );
  OR2_X1 U6584 ( .A1(n5514), .A2(n5083), .ZN(n5084) );
  NOR2_X1 U6585 ( .A1(n6961), .A2(n5210), .ZN(n5091) );
  NAND2_X1 U6586 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5090), .ZN(n5089) );
  XNOR2_X1 U6587 ( .A(n5094), .B(n5093), .ZN(n6672) );
  INV_X1 U6588 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6664) );
  NAND2_X1 U6589 ( .A1(n5101), .A2(n10062), .ZN(n6200) );
  NAND2_X1 U6590 ( .A1(n7628), .A2(n6197), .ZN(n5103) );
  NAND2_X1 U6591 ( .A1(n5103), .A2(n5102), .ZN(n6947) );
  OR2_X1 U6592 ( .A1(n5356), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5108) );
  INV_X1 U6593 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5104) );
  OR2_X1 U6594 ( .A1(n5514), .A2(n5104), .ZN(n5107) );
  NAND2_X1 U6595 ( .A1(n6161), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5106) );
  NAND2_X1 U6596 ( .A1(n5082), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5105) );
  NAND2_X1 U6597 ( .A1(n5109), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5110) );
  MUX2_X1 U6598 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5110), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5112) );
  NAND2_X1 U6599 ( .A1(n5112), .A2(n5111), .ZN(n7018) );
  INV_X1 U6600 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6666) );
  OR2_X1 U6601 ( .A1(n5096), .A2(n6666), .ZN(n5116) );
  XNOR2_X1 U6602 ( .A(n5114), .B(n5113), .ZN(n6674) );
  OR2_X1 U6603 ( .A1(n5095), .A2(n6674), .ZN(n5115) );
  OAI211_X1 U6604 ( .C1(n5088), .C2(n7018), .A(n5116), .B(n5115), .ZN(n7924)
         );
  NOR2_X1 U6605 ( .A1(n8370), .A2(n7924), .ZN(n5118) );
  NAND2_X1 U6606 ( .A1(n8370), .A2(n7924), .ZN(n5117) );
  NAND2_X1 U6607 ( .A1(n6161), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5126) );
  INV_X1 U6608 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5119) );
  OR2_X1 U6609 ( .A1(n5120), .A2(n5119), .ZN(n5125) );
  NAND2_X1 U6610 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5121) );
  AND2_X1 U6611 ( .A1(n5135), .A2(n5121), .ZN(n7690) );
  OR2_X1 U6612 ( .A1(n5356), .A2(n7690), .ZN(n5124) );
  INV_X1 U6613 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n5122) );
  OR2_X1 U6614 ( .A1(n5514), .A2(n5122), .ZN(n5123) );
  AND4_X2 U6615 ( .A1(n5126), .A2(n5125), .A3(n5124), .A4(n5123), .ZN(n7614)
         );
  NAND2_X1 U6616 ( .A1(n5111), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5128) );
  INV_X1 U6617 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5127) );
  XNOR2_X1 U6618 ( .A(n5128), .B(n5127), .ZN(n7498) );
  XNOR2_X1 U6619 ( .A(n5130), .B(n5129), .ZN(n6670) );
  OR2_X1 U6620 ( .A1(n5095), .A2(n6670), .ZN(n5132) );
  INV_X1 U6621 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6667) );
  OR2_X1 U6622 ( .A1(n5096), .A2(n6667), .ZN(n5131) );
  OAI211_X1 U6623 ( .C1(n5088), .C2(n7498), .A(n5132), .B(n5131), .ZN(n7542)
         );
  INV_X1 U6624 ( .A(n7542), .ZN(n7743) );
  NAND2_X1 U6625 ( .A1(n7614), .A2(n7743), .ZN(n5133) );
  NAND2_X1 U6626 ( .A1(n8369), .A2(n7542), .ZN(n5134) );
  NAND2_X1 U6627 ( .A1(n6161), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5140) );
  NAND2_X1 U6628 ( .A1(n5135), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5136) );
  AND2_X1 U6629 ( .A1(n5151), .A2(n5136), .ZN(n7620) );
  OR2_X1 U6630 ( .A1(n5356), .A2(n7620), .ZN(n5139) );
  NAND2_X1 U6631 ( .A1(n6162), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5138) );
  NAND2_X1 U6632 ( .A1(n5405), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5137) );
  NAND4_X1 U6633 ( .A1(n5140), .A2(n5139), .A3(n5138), .A4(n5137), .ZN(n8368)
         );
  OR2_X1 U6634 ( .A1(n5141), .A2(n5210), .ZN(n5143) );
  XNOR2_X1 U6635 ( .A(n5143), .B(n5142), .ZN(n7020) );
  XNOR2_X1 U6636 ( .A(n5145), .B(n5144), .ZN(n6682) );
  OR2_X1 U6637 ( .A1(n5095), .A2(n6682), .ZN(n5147) );
  INV_X1 U6638 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6668) );
  OR2_X1 U6639 ( .A1(n5096), .A2(n6668), .ZN(n5146) );
  OAI211_X1 U6640 ( .C1(n5088), .C2(n7020), .A(n5147), .B(n5146), .ZN(n7585)
         );
  INV_X1 U6641 ( .A(n7585), .ZN(n7721) );
  NAND2_X1 U6642 ( .A1(n7642), .A2(n7721), .ZN(n5148) );
  NAND2_X1 U6643 ( .A1(n8368), .A2(n7585), .ZN(n5149) );
  NAND2_X1 U6644 ( .A1(n5150), .A2(n5149), .ZN(n7547) );
  NAND2_X1 U6645 ( .A1(n6162), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5156) );
  NAND2_X1 U6646 ( .A1(n5151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5152) );
  AND2_X1 U6647 ( .A1(n5166), .A2(n5152), .ZN(n7648) );
  OR2_X1 U6648 ( .A1(n5356), .A2(n7648), .ZN(n5155) );
  NAND2_X1 U6649 ( .A1(n6161), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5154) );
  NAND2_X1 U6650 ( .A1(n5405), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5153) );
  NAND4_X1 U6651 ( .A1(n5156), .A2(n5155), .A3(n5154), .A4(n5153), .ZN(n8367)
         );
  NOR2_X1 U6652 ( .A1(n5157), .A2(n5210), .ZN(n5158) );
  MUX2_X1 U6653 ( .A(n5210), .B(n5158), .S(P2_IR_REG_6__SCAN_IN), .Z(n5161) );
  INV_X1 U6654 ( .A(n5159), .ZN(n5160) );
  XNOR2_X1 U6655 ( .A(n5163), .B(n5162), .ZN(n6678) );
  OR2_X1 U6656 ( .A1(n5095), .A2(n6678), .ZN(n5165) );
  INV_X1 U6657 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6677) );
  OR2_X1 U6658 ( .A1(n5096), .A2(n6677), .ZN(n5164) );
  OAI211_X1 U6659 ( .C1(n5088), .C2(n7419), .A(n5165), .B(n5164), .ZN(n7645)
         );
  INV_X1 U6660 ( .A(n7645), .ZN(n7550) );
  NAND2_X1 U6661 ( .A1(n7864), .A2(n7550), .ZN(n6348) );
  NAND2_X1 U6662 ( .A1(n8367), .A2(n7645), .ZN(n6347) );
  OR2_X1 U6663 ( .A1(n5514), .A2(n4708), .ZN(n5171) );
  NAND2_X1 U6664 ( .A1(n5166), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5167) );
  AND2_X1 U6665 ( .A1(n5180), .A2(n5167), .ZN(n7749) );
  OR2_X1 U6666 ( .A1(n5356), .A2(n7749), .ZN(n5170) );
  NAND2_X1 U6667 ( .A1(n6162), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5169) );
  NAND2_X1 U6668 ( .A1(n6161), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5168) );
  NAND4_X1 U6669 ( .A1(n5171), .A2(n5170), .A3(n5169), .A4(n5168), .ZN(n8366)
         );
  NAND2_X1 U6670 ( .A1(n5159), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5172) );
  XNOR2_X1 U6671 ( .A(n5172), .B(n5001), .ZN(n7403) );
  OR2_X1 U6672 ( .A1(n5095), .A2(n6681), .ZN(n5176) );
  INV_X1 U6673 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6680) );
  OR2_X1 U6674 ( .A1(n5096), .A2(n6680), .ZN(n5175) );
  OAI211_X1 U6675 ( .C1(n5088), .C2(n7403), .A(n5176), .B(n5175), .ZN(n7927)
         );
  XNOR2_X1 U6676 ( .A(n8366), .B(n7927), .ZN(n6350) );
  INV_X1 U6677 ( .A(n8366), .ZN(n7960) );
  INV_X1 U6678 ( .A(n7927), .ZN(n7526) );
  NAND2_X1 U6679 ( .A1(n7960), .A2(n7526), .ZN(n5177) );
  NAND2_X1 U6680 ( .A1(n6162), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5185) );
  NAND2_X1 U6681 ( .A1(n5180), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5181) );
  AND2_X1 U6682 ( .A1(n5195), .A2(n5181), .ZN(n7966) );
  OR2_X1 U6683 ( .A1(n5356), .A2(n7966), .ZN(n5184) );
  NAND2_X1 U6684 ( .A1(n5405), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5183) );
  NAND2_X1 U6685 ( .A1(n6161), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5182) );
  NAND4_X1 U6686 ( .A1(n5185), .A2(n5184), .A3(n5183), .A4(n5182), .ZN(n8365)
         );
  INV_X1 U6687 ( .A(n8365), .ZN(n7955) );
  NAND2_X1 U6688 ( .A1(n6690), .A2(n6175), .ZN(n5193) );
  NAND2_X1 U6689 ( .A1(n5471), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n5192) );
  NAND2_X1 U6690 ( .A1(n5189), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5190) );
  XNOR2_X1 U6691 ( .A(n5190), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7464) );
  NAND2_X1 U6692 ( .A1(n6661), .A2(n7464), .ZN(n5191) );
  INV_X1 U6693 ( .A(n7954), .ZN(n7963) );
  NAND2_X1 U6694 ( .A1(n7955), .A2(n7963), .ZN(n6233) );
  NAND2_X1 U6695 ( .A1(n8365), .A2(n7954), .ZN(n6229) );
  NAND2_X1 U6696 ( .A1(n6233), .A2(n6229), .ZN(n7737) );
  NAND2_X1 U6697 ( .A1(n7738), .A2(n7737), .ZN(n7736) );
  NAND2_X1 U6698 ( .A1(n8365), .A2(n7963), .ZN(n5194) );
  NAND2_X1 U6699 ( .A1(n6161), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5200) );
  NAND2_X1 U6700 ( .A1(n5195), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5196) );
  AND2_X1 U6701 ( .A1(n5218), .A2(n5196), .ZN(n8295) );
  OR2_X1 U6702 ( .A1(n5356), .A2(n8295), .ZN(n5199) );
  NAND2_X1 U6703 ( .A1(n6162), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5198) );
  NAND2_X1 U6704 ( .A1(n5405), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5197) );
  NAND4_X1 U6705 ( .A1(n5200), .A2(n5199), .A3(n5198), .A4(n5197), .ZN(n8364)
         );
  INV_X1 U6706 ( .A(n8364), .ZN(n7959) );
  XNOR2_X2 U6707 ( .A(n5201), .B(n4914), .ZN(n6697) );
  NAND2_X1 U6708 ( .A1(n6697), .A2(n6175), .ZN(n5206) );
  NAND2_X1 U6709 ( .A1(n5203), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5204) );
  XNOR2_X1 U6710 ( .A(n5204), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7455) );
  AOI22_X1 U6711 ( .A1(n5471), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6661), .B2(
        n7455), .ZN(n5205) );
  NAND2_X1 U6712 ( .A1(n5206), .A2(n5205), .ZN(n8296) );
  NAND2_X1 U6713 ( .A1(n7959), .A2(n8296), .ZN(n6234) );
  INV_X1 U6714 ( .A(n8296), .ZN(n7790) );
  NAND2_X1 U6715 ( .A1(n7790), .A2(n8364), .ZN(n6230) );
  INV_X1 U6716 ( .A(n6351), .ZN(n5207) );
  NAND2_X1 U6717 ( .A1(n7959), .A2(n7790), .ZN(n5208) );
  NAND2_X1 U6718 ( .A1(n6701), .A2(n6175), .ZN(n5215) );
  OR2_X1 U6719 ( .A1(n5211), .A2(n5210), .ZN(n5213) );
  XNOR2_X1 U6720 ( .A(n5213), .B(n5212), .ZN(n7708) );
  INV_X1 U6721 ( .A(n7708), .ZN(n7654) );
  AOI22_X1 U6722 ( .A1(n5471), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6661), .B2(
        n7654), .ZN(n5214) );
  INV_X1 U6723 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n5217) );
  OR2_X1 U6724 ( .A1(n5216), .A2(n5217), .ZN(n5223) );
  NAND2_X1 U6725 ( .A1(n5218), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5219) );
  AND2_X1 U6726 ( .A1(n5230), .A2(n5219), .ZN(n8048) );
  OR2_X1 U6727 ( .A1(n5356), .A2(n8048), .ZN(n5222) );
  INV_X1 U6728 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7893) );
  OR2_X1 U6729 ( .A1(n5514), .A2(n7893), .ZN(n5221) );
  NAND2_X1 U6730 ( .A1(n6162), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5220) );
  NAND4_X1 U6731 ( .A1(n5223), .A2(n5222), .A3(n5221), .A4(n5220), .ZN(n8363)
         );
  INV_X1 U6732 ( .A(n8053), .ZN(n7895) );
  NAND2_X1 U6733 ( .A1(n7895), .A2(n8363), .ZN(n8030) );
  XNOR2_X1 U6734 ( .A(n5224), .B(SI_11_), .ZN(n5225) );
  XNOR2_X1 U6735 ( .A(n5226), .B(n5225), .ZN(n6705) );
  NAND2_X1 U6736 ( .A1(n6705), .A2(n6175), .ZN(n5229) );
  NAND2_X1 U6737 ( .A1(n5244), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5227) );
  XNOR2_X1 U6738 ( .A(n5227), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7820) );
  AOI22_X1 U6739 ( .A1(n5471), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6661), .B2(
        n7820), .ZN(n5228) );
  NAND2_X1 U6740 ( .A1(n5229), .A2(n5228), .ZN(n7967) );
  NAND2_X1 U6741 ( .A1(n6162), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5236) );
  INV_X1 U6742 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7935) );
  OR2_X1 U6743 ( .A1(n5514), .A2(n7935), .ZN(n5235) );
  NAND2_X1 U6744 ( .A1(n5230), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5231) );
  AND2_X1 U6745 ( .A1(n5248), .A2(n5231), .ZN(n8093) );
  OR2_X1 U6746 ( .A1(n5356), .A2(n8093), .ZN(n5234) );
  INV_X1 U6747 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n5232) );
  OR2_X1 U6748 ( .A1(n5216), .A2(n5232), .ZN(n5233) );
  AND2_X1 U6749 ( .A1(n7967), .A2(n8362), .ZN(n5237) );
  OR2_X1 U6750 ( .A1(n7933), .A2(n5237), .ZN(n5239) );
  OR2_X1 U6751 ( .A1(n7967), .A2(n8362), .ZN(n5238) );
  NAND2_X1 U6752 ( .A1(n5241), .A2(n5240), .ZN(n5242) );
  NAND2_X1 U6753 ( .A1(n5243), .A2(n5242), .ZN(n6732) );
  OR2_X1 U6754 ( .A1(n6732), .A2(n5095), .ZN(n5247) );
  NAND2_X1 U6755 ( .A1(n5258), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5245) );
  XNOR2_X1 U6756 ( .A(n5245), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7813) );
  AOI22_X1 U6757 ( .A1(n5471), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6661), .B2(
        n7813), .ZN(n5246) );
  OR2_X1 U6758 ( .A1(n5216), .A2(n8382), .ZN(n5253) );
  NAND2_X1 U6759 ( .A1(n5248), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5249) );
  AND2_X1 U6760 ( .A1(n5261), .A2(n5249), .ZN(n8038) );
  OR2_X1 U6761 ( .A1(n5356), .A2(n8038), .ZN(n5252) );
  INV_X1 U6762 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7979) );
  OR2_X1 U6763 ( .A1(n5514), .A2(n7979), .ZN(n5251) );
  NAND2_X1 U6764 ( .A1(n6162), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5250) );
  NAND4_X1 U6765 ( .A1(n5253), .A2(n5252), .A3(n5251), .A4(n5250), .ZN(n8361)
         );
  NAND2_X1 U6766 ( .A1(n8041), .A2(n8097), .ZN(n6250) );
  NAND2_X1 U6767 ( .A1(n6251), .A2(n6250), .ZN(n7975) );
  NAND2_X1 U6768 ( .A1(n8041), .A2(n8361), .ZN(n5254) );
  XNOR2_X1 U6769 ( .A(n5255), .B(SI_13_), .ZN(n5256) );
  XNOR2_X1 U6770 ( .A(n5257), .B(n5256), .ZN(n6809) );
  NAND2_X1 U6771 ( .A1(n6809), .A2(n6175), .ZN(n5260) );
  OR2_X1 U6772 ( .A1(n5308), .A2(n5210), .ZN(n5271) );
  XNOR2_X1 U6773 ( .A(n5271), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8403) );
  AOI22_X1 U6774 ( .A1(n5471), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6661), .B2(
        n8403), .ZN(n5259) );
  NAND2_X1 U6775 ( .A1(n6162), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5266) );
  INV_X1 U6776 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8376) );
  OR2_X1 U6777 ( .A1(n5216), .A2(n8376), .ZN(n5265) );
  NAND2_X1 U6778 ( .A1(n5261), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5262) );
  AND2_X1 U6779 ( .A1(n5278), .A2(n5262), .ZN(n8079) );
  OR2_X1 U6780 ( .A1(n5356), .A2(n8079), .ZN(n5264) );
  INV_X1 U6781 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8377) );
  OR2_X1 U6782 ( .A1(n5514), .A2(n8377), .ZN(n5263) );
  OR2_X1 U6783 ( .A1(n8077), .A2(n8360), .ZN(n6345) );
  NAND2_X1 U6784 ( .A1(n8077), .A2(n8360), .ZN(n6344) );
  NAND2_X1 U6785 ( .A1(n5267), .A2(n6344), .ZN(n8112) );
  XNOR2_X1 U6786 ( .A(n5268), .B(SI_14_), .ZN(n5269) );
  XNOR2_X1 U6787 ( .A(n5270), .B(n5269), .ZN(n6838) );
  NAND2_X1 U6788 ( .A1(n6838), .A2(n6175), .ZN(n5277) );
  INV_X1 U6789 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5306) );
  NAND2_X1 U6790 ( .A1(n5271), .A2(n5306), .ZN(n5272) );
  NAND2_X1 U6791 ( .A1(n5272), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5274) );
  INV_X1 U6792 ( .A(n5274), .ZN(n5273) );
  NAND2_X1 U6793 ( .A1(n5273), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n5275) );
  NAND2_X1 U6794 ( .A1(n5274), .A2(n5305), .ZN(n5290) );
  AOI22_X1 U6795 ( .A1(n5471), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8417), .B2(
        n6661), .ZN(n5276) );
  INV_X1 U6796 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8409) );
  OR2_X1 U6797 ( .A1(n5216), .A2(n8409), .ZN(n5283) );
  NAND2_X1 U6798 ( .A1(n5278), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5279) );
  AND2_X1 U6799 ( .A1(n5294), .A2(n5279), .ZN(n8215) );
  OR2_X1 U6800 ( .A1(n5356), .A2(n8215), .ZN(n5282) );
  INV_X1 U6801 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8410) );
  OR2_X1 U6802 ( .A1(n5514), .A2(n8410), .ZN(n5281) );
  NAND2_X1 U6803 ( .A1(n6162), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5280) );
  NAND4_X1 U6804 ( .A1(n5283), .A2(n5282), .A3(n5281), .A4(n5280), .ZN(n8727)
         );
  AND2_X1 U6805 ( .A1(n8149), .A2(n8727), .ZN(n5285) );
  OR2_X1 U6806 ( .A1(n8149), .A2(n8727), .ZN(n5284) );
  INV_X1 U6807 ( .A(SI_15_), .ZN(n5286) );
  XNOR2_X1 U6808 ( .A(n5287), .B(n5286), .ZN(n5288) );
  XNOR2_X1 U6809 ( .A(n5289), .B(n5288), .ZN(n6857) );
  NAND2_X1 U6810 ( .A1(n6857), .A2(n6175), .ZN(n5293) );
  NAND2_X1 U6811 ( .A1(n5290), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5291) );
  XNOR2_X1 U6812 ( .A(n5291), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8458) );
  AOI22_X1 U6813 ( .A1(n6661), .A2(n8458), .B1(n5471), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5292) );
  INV_X1 U6814 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8431) );
  OR2_X1 U6815 ( .A1(n5514), .A2(n8431), .ZN(n5299) );
  NAND2_X1 U6816 ( .A1(n5294), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5295) );
  AND2_X1 U6817 ( .A1(n5312), .A2(n5295), .ZN(n8732) );
  OR2_X1 U6818 ( .A1(n5356), .A2(n8732), .ZN(n5298) );
  INV_X1 U6819 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8430) );
  OR2_X1 U6820 ( .A1(n5216), .A2(n8430), .ZN(n5297) );
  NAND2_X1 U6821 ( .A1(n6162), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5296) );
  NAND4_X1 U6822 ( .A1(n5299), .A2(n5298), .A3(n5297), .A4(n5296), .ZN(n8709)
         );
  NOR2_X1 U6823 ( .A1(n8792), .A2(n8709), .ZN(n5300) );
  INV_X1 U6824 ( .A(n8709), .ZN(n8217) );
  INV_X1 U6825 ( .A(n8792), .ZN(n8355) );
  XNOR2_X1 U6826 ( .A(n5301), .B(SI_16_), .ZN(n5302) );
  XNOR2_X1 U6827 ( .A(n5303), .B(n5302), .ZN(n6926) );
  NAND2_X1 U6828 ( .A1(n6926), .A2(n6175), .ZN(n5311) );
  INV_X1 U6829 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5304) );
  AND3_X1 U6830 ( .A1(n5306), .A2(n5305), .A3(n5304), .ZN(n5307) );
  OR2_X1 U6831 ( .A1(n5323), .A2(n5210), .ZN(n5309) );
  XNOR2_X1 U6832 ( .A(n5309), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8461) );
  AOI22_X1 U6833 ( .A1(n5471), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6661), .B2(
        n8461), .ZN(n5310) );
  NAND2_X1 U6834 ( .A1(n6162), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5317) );
  INV_X1 U6835 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8787) );
  OR2_X1 U6836 ( .A1(n5216), .A2(n8787), .ZN(n5316) );
  NAND2_X1 U6837 ( .A1(n5312), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5313) );
  AND2_X1 U6838 ( .A1(n5327), .A2(n5313), .ZN(n8717) );
  OR2_X1 U6839 ( .A1(n5356), .A2(n8717), .ZN(n5315) );
  INV_X1 U6840 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8716) );
  OR2_X1 U6841 ( .A1(n5514), .A2(n8716), .ZN(n5314) );
  NAND2_X1 U6842 ( .A1(n8867), .A2(n8346), .ZN(n6267) );
  NAND2_X1 U6843 ( .A1(n6266), .A2(n6267), .ZN(n8705) );
  NAND2_X1 U6844 ( .A1(n8708), .A2(n8705), .ZN(n5319) );
  INV_X1 U6845 ( .A(n8346), .ZN(n8729) );
  NAND2_X1 U6846 ( .A1(n8867), .A2(n8729), .ZN(n5318) );
  XNOR2_X1 U6847 ( .A(n5321), .B(n5320), .ZN(n7103) );
  NAND2_X1 U6848 ( .A1(n7103), .A2(n6175), .ZN(n5326) );
  INV_X1 U6849 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5322) );
  NAND2_X1 U6850 ( .A1(n5336), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5324) );
  XNOR2_X1 U6851 ( .A(n5324), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8505) );
  AOI22_X1 U6852 ( .A1(n5471), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6661), .B2(
        n8505), .ZN(n5325) );
  NAND2_X1 U6853 ( .A1(n6162), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5332) );
  INV_X1 U6854 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8700) );
  OR2_X1 U6855 ( .A1(n5514), .A2(n8700), .ZN(n5331) );
  NAND2_X1 U6856 ( .A1(n5327), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5328) );
  AND2_X1 U6857 ( .A1(n5339), .A2(n5328), .ZN(n8701) );
  OR2_X1 U6858 ( .A1(n5356), .A2(n8701), .ZN(n5330) );
  INV_X1 U6859 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8783) );
  OR2_X1 U6860 ( .A1(n5216), .A2(n8783), .ZN(n5329) );
  NAND2_X1 U6861 ( .A1(n8860), .A2(n8712), .ZN(n6272) );
  NAND2_X1 U6862 ( .A1(n6274), .A2(n6272), .ZN(n6340) );
  INV_X1 U6863 ( .A(n8712), .ZN(n8688) );
  NAND2_X1 U6864 ( .A1(n4402), .A2(n5333), .ZN(n5334) );
  NAND2_X1 U6865 ( .A1(n5335), .A2(n5334), .ZN(n7122) );
  OR2_X1 U6866 ( .A1(n7122), .A2(n5095), .ZN(n5338) );
  XNOR2_X1 U6867 ( .A(n5349), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8532) );
  AOI22_X1 U6868 ( .A1(n5471), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8532), .B2(
        n6661), .ZN(n5337) );
  NAND2_X1 U6869 ( .A1(n6161), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5344) );
  NAND2_X1 U6870 ( .A1(n5339), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5340) );
  AND2_X1 U6871 ( .A1(n5354), .A2(n5340), .ZN(n8692) );
  OR2_X1 U6872 ( .A1(n5356), .A2(n8692), .ZN(n5343) );
  NAND2_X1 U6873 ( .A1(n6162), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5342) );
  NAND2_X1 U6874 ( .A1(n5405), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5341) );
  NAND4_X1 U6875 ( .A1(n5344), .A2(n5343), .A3(n5342), .A4(n5341), .ZN(n8698)
         );
  AND2_X1 U6876 ( .A1(n8854), .A2(n8698), .ZN(n5345) );
  INV_X1 U6877 ( .A(n8677), .ZN(n5361) );
  XNOR2_X1 U6878 ( .A(n5347), .B(n5346), .ZN(n7553) );
  NAND2_X1 U6879 ( .A1(n7553), .A2(n6175), .ZN(n5353) );
  INV_X1 U6880 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5350) );
  AOI22_X1 U6881 ( .A1(n8539), .A2(n6661), .B1(n5471), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n5352) );
  NAND2_X1 U6882 ( .A1(n5354), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5355) );
  AND2_X1 U6883 ( .A1(n5369), .A2(n5355), .ZN(n8681) );
  OR2_X1 U6884 ( .A1(n5356), .A2(n8681), .ZN(n5360) );
  INV_X1 U6885 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8680) );
  OR2_X1 U6886 ( .A1(n5514), .A2(n8680), .ZN(n5359) );
  NAND2_X1 U6887 ( .A1(n6161), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5358) );
  NAND2_X1 U6888 ( .A1(n6162), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5357) );
  NAND4_X1 U6889 ( .A1(n5360), .A2(n5359), .A3(n5358), .A4(n5357), .ZN(n8689)
         );
  NAND2_X1 U6890 ( .A1(n8848), .A2(n8689), .ZN(n5362) );
  XNOR2_X1 U6891 ( .A(n5364), .B(n5363), .ZN(n5365) );
  XNOR2_X1 U6892 ( .A(n5366), .B(n5365), .ZN(n7674) );
  NAND2_X1 U6893 ( .A1(n7674), .A2(n6175), .ZN(n5368) );
  NAND2_X1 U6894 ( .A1(n5471), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5367) );
  NAND2_X1 U6895 ( .A1(n6162), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5374) );
  NAND2_X1 U6896 ( .A1(n6161), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5373) );
  NAND2_X1 U6897 ( .A1(n5369), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5370) );
  NAND2_X1 U6898 ( .A1(n5383), .A2(n5370), .ZN(n8672) );
  NAND2_X1 U6899 ( .A1(n5491), .A2(n8672), .ZN(n5372) );
  NAND2_X1 U6900 ( .A1(n5405), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5371) );
  NAND4_X1 U6901 ( .A1(n5374), .A2(n5373), .A3(n5372), .A4(n5371), .ZN(n8678)
         );
  NAND2_X1 U6902 ( .A1(n8773), .A2(n8246), .ZN(n8647) );
  OR2_X1 U6903 ( .A1(n8773), .A2(n8678), .ZN(n8652) );
  NAND2_X1 U6904 ( .A1(n8650), .A2(n8652), .ZN(n5387) );
  XNOR2_X1 U6905 ( .A(n5376), .B(SI_21_), .ZN(n5377) );
  XNOR2_X1 U6906 ( .A(n5378), .B(n5377), .ZN(n7842) );
  NAND2_X1 U6907 ( .A1(n7842), .A2(n6175), .ZN(n5380) );
  NAND2_X1 U6908 ( .A1(n5471), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5379) );
  INV_X1 U6909 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8657) );
  NAND2_X1 U6910 ( .A1(n6162), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5382) );
  NAND2_X1 U6911 ( .A1(n6161), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5381) );
  AND2_X1 U6912 ( .A1(n5382), .A2(n5381), .ZN(n5386) );
  NAND2_X1 U6913 ( .A1(n5383), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5384) );
  NAND2_X1 U6914 ( .A1(n5392), .A2(n5384), .ZN(n8658) );
  NAND2_X1 U6915 ( .A1(n8658), .A2(n5491), .ZN(n5385) );
  OAI211_X1 U6916 ( .C1(n5514), .C2(n8657), .A(n5386), .B(n5385), .ZN(n8640)
         );
  INV_X1 U6917 ( .A(n8640), .ZN(n8667) );
  NAND2_X1 U6918 ( .A1(n8836), .A2(n8667), .ZN(n6294) );
  NAND2_X1 U6919 ( .A1(n6290), .A2(n6294), .ZN(n8651) );
  NAND2_X1 U6920 ( .A1(n5387), .A2(n8651), .ZN(n8635) );
  OR2_X1 U6921 ( .A1(n8836), .A2(n8640), .ZN(n8636) );
  NAND2_X1 U6922 ( .A1(n8635), .A2(n8636), .ZN(n5397) );
  XNOR2_X1 U6923 ( .A(n5389), .B(n5388), .ZN(n7939) );
  NAND2_X1 U6924 ( .A1(n7939), .A2(n6175), .ZN(n5391) );
  NAND2_X1 U6925 ( .A1(n5471), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5390) );
  INV_X1 U6926 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8643) );
  NAND2_X1 U6927 ( .A1(n5392), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5393) );
  NAND2_X1 U6928 ( .A1(n5403), .A2(n5393), .ZN(n8644) );
  NAND2_X1 U6929 ( .A1(n8644), .A2(n5491), .ZN(n5395) );
  AOI22_X1 U6930 ( .A1(n6161), .A2(P2_REG1_REG_22__SCAN_IN), .B1(n6162), .B2(
        P2_REG0_REG_22__SCAN_IN), .ZN(n5394) );
  INV_X1 U6931 ( .A(n8655), .ZN(n5396) );
  NAND2_X1 U6932 ( .A1(n8830), .A2(n5396), .ZN(n6284) );
  NAND2_X1 U6933 ( .A1(n6292), .A2(n6284), .ZN(n6362) );
  NAND2_X1 U6934 ( .A1(n5397), .A2(n6362), .ZN(n8639) );
  OR2_X1 U6935 ( .A1(n8830), .A2(n8655), .ZN(n5398) );
  XNOR2_X1 U6936 ( .A(n5400), .B(n5399), .ZN(n7949) );
  NAND2_X1 U6937 ( .A1(n7949), .A2(n6175), .ZN(n5402) );
  NAND2_X1 U6938 ( .A1(n5471), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5401) );
  NAND2_X1 U6939 ( .A1(n5403), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5404) );
  NAND2_X1 U6940 ( .A1(n5416), .A2(n5404), .ZN(n8631) );
  NAND2_X1 U6941 ( .A1(n8631), .A2(n5491), .ZN(n5408) );
  AOI22_X1 U6942 ( .A1(n6161), .A2(P2_REG1_REG_23__SCAN_IN), .B1(n6162), .B2(
        P2_REG0_REG_23__SCAN_IN), .ZN(n5407) );
  NAND2_X1 U6943 ( .A1(n5405), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5406) );
  NAND2_X1 U6944 ( .A1(n8824), .A2(n8641), .ZN(n5409) );
  NAND2_X1 U6945 ( .A1(n8627), .A2(n5409), .ZN(n5411) );
  OR2_X1 U6946 ( .A1(n8824), .A2(n8641), .ZN(n5410) );
  NAND2_X1 U6947 ( .A1(n5411), .A2(n5410), .ZN(n8611) );
  NAND2_X1 U6948 ( .A1(n5956), .A2(n6175), .ZN(n5415) );
  NAND2_X1 U6949 ( .A1(n5471), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5414) );
  NAND2_X1 U6950 ( .A1(n5416), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5417) );
  NAND2_X1 U6951 ( .A1(n5418), .A2(n5417), .ZN(n8614) );
  NAND2_X1 U6952 ( .A1(n8614), .A2(n5491), .ZN(n5423) );
  INV_X1 U6953 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8621) );
  NAND2_X1 U6954 ( .A1(n6162), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5420) );
  NAND2_X1 U6955 ( .A1(n6161), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5419) );
  OAI211_X1 U6956 ( .C1(n8621), .C2(n5514), .A(n5420), .B(n5419), .ZN(n5421)
         );
  INV_X1 U6957 ( .A(n5421), .ZN(n5422) );
  NAND2_X1 U6958 ( .A1(n8818), .A2(n8628), .ZN(n5424) );
  NAND2_X1 U6959 ( .A1(n8256), .A2(n8588), .ZN(n5541) );
  NAND2_X1 U6960 ( .A1(n5426), .A2(n5425), .ZN(n5430) );
  INV_X1 U6961 ( .A(n5427), .ZN(n5428) );
  NAND2_X1 U6962 ( .A1(n5428), .A2(n7293), .ZN(n5429) );
  MUX2_X1 U6963 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .S(n4350), .Z(n5441) );
  XNOR2_X1 U6964 ( .A(n5441), .B(n7337), .ZN(n5462) );
  XNOR2_X1 U6965 ( .A(n5464), .B(n5462), .ZN(n8059) );
  NAND2_X1 U6966 ( .A1(n8059), .A2(n6175), .ZN(n5432) );
  NAND2_X1 U6967 ( .A1(n5471), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5431) );
  NAND2_X1 U6968 ( .A1(n5433), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5434) );
  NAND2_X1 U6969 ( .A1(n5449), .A2(n5434), .ZN(n8590) );
  NAND2_X1 U6970 ( .A1(n8590), .A2(n5491), .ZN(n5439) );
  INV_X1 U6971 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8593) );
  NAND2_X1 U6972 ( .A1(n6161), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5436) );
  NAND2_X1 U6973 ( .A1(n6162), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5435) );
  OAI211_X1 U6974 ( .C1(n8593), .C2(n5514), .A(n5436), .B(n5435), .ZN(n5437)
         );
  INV_X1 U6975 ( .A(n5437), .ZN(n5438) );
  NOR2_X1 U6976 ( .A1(n8807), .A2(n8578), .ZN(n5440) );
  NAND2_X1 U6977 ( .A1(n5464), .A2(n5462), .ZN(n5443) );
  INV_X1 U6978 ( .A(n5441), .ZN(n5442) );
  NAND2_X1 U6979 ( .A1(n5442), .A2(n7337), .ZN(n5467) );
  MUX2_X1 U6980 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .S(n4350), .Z(n5458) );
  INV_X1 U6981 ( .A(SI_27_), .ZN(n7295) );
  XNOR2_X1 U6982 ( .A(n5458), .B(n7295), .ZN(n5460) );
  NAND2_X1 U6983 ( .A1(n8070), .A2(n6175), .ZN(n5446) );
  NAND2_X1 U6984 ( .A1(n5471), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5445) );
  INV_X1 U6985 ( .A(n5449), .ZN(n5448) );
  INV_X1 U6986 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5447) );
  NAND2_X1 U6987 ( .A1(n5449), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5450) );
  NAND2_X1 U6988 ( .A1(n5474), .A2(n5450), .ZN(n8581) );
  NAND2_X1 U6989 ( .A1(n8581), .A2(n5491), .ZN(n5456) );
  INV_X1 U6990 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n5453) );
  NAND2_X1 U6991 ( .A1(n6161), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5452) );
  NAND2_X1 U6992 ( .A1(n6162), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5451) );
  OAI211_X1 U6993 ( .C1(n5453), .C2(n5514), .A(n5452), .B(n5451), .ZN(n5454)
         );
  INV_X1 U6994 ( .A(n5454), .ZN(n5455) );
  NOR2_X1 U6995 ( .A1(n8210), .A2(n8358), .ZN(n5457) );
  INV_X2 U6996 ( .A(n8358), .ZN(n8589) );
  INV_X1 U6997 ( .A(n5458), .ZN(n5459) );
  NAND2_X1 U6998 ( .A1(n5459), .A2(n7295), .ZN(n5466) );
  INV_X1 U6999 ( .A(n5466), .ZN(n5461) );
  OR2_X1 U7000 ( .A1(n5461), .A2(n5460), .ZN(n5465) );
  INV_X1 U7001 ( .A(n5465), .ZN(n5469) );
  AND2_X1 U7002 ( .A1(n5467), .A2(n5466), .ZN(n5468) );
  MUX2_X1 U7003 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n4350), .Z(n5484) );
  INV_X1 U7004 ( .A(SI_28_), .ZN(n7335) );
  XNOR2_X1 U7005 ( .A(n5484), .B(n7335), .ZN(n5482) );
  XNOR2_X1 U7006 ( .A(n5483), .B(n5482), .ZN(n8104) );
  NAND2_X1 U7007 ( .A1(n8104), .A2(n6175), .ZN(n5473) );
  NAND2_X1 U7008 ( .A1(n5471), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5472) );
  NAND2_X1 U7009 ( .A1(n5474), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5475) );
  NAND2_X1 U7010 ( .A1(n5490), .A2(n5475), .ZN(n8570) );
  NAND2_X1 U7011 ( .A1(n8570), .A2(n5491), .ZN(n5481) );
  INV_X1 U7012 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n5478) );
  NAND2_X1 U7013 ( .A1(n6161), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5477) );
  NAND2_X1 U7014 ( .A1(n6162), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5476) );
  OAI211_X1 U7015 ( .C1(n5478), .C2(n5514), .A(n5477), .B(n5476), .ZN(n5479)
         );
  INV_X1 U7016 ( .A(n5479), .ZN(n5480) );
  AOI22_X1 U7017 ( .A1(n8562), .A2(n8568), .B1(n8197), .B2(n8357), .ZN(n5496)
         );
  INV_X1 U7018 ( .A(n5484), .ZN(n5485) );
  NAND2_X1 U7019 ( .A1(n5485), .A2(n7335), .ZN(n5486) );
  INV_X1 U7020 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8881) );
  INV_X1 U7021 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9730) );
  MUX2_X1 U7022 ( .A(n8881), .B(n9730), .S(n4350), .Z(n6153) );
  NAND2_X1 U7023 ( .A1(n8879), .A2(n6175), .ZN(n5489) );
  OR2_X1 U7024 ( .A1(n5096), .A2(n8881), .ZN(n5488) );
  NAND2_X1 U7025 ( .A1(n8547), .A2(n5491), .ZN(n6168) );
  INV_X1 U7026 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8556) );
  NAND2_X1 U7027 ( .A1(n6161), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5493) );
  NAND2_X1 U7028 ( .A1(n6162), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5492) );
  OAI211_X1 U7029 ( .C1(n8556), .C2(n5514), .A(n5493), .B(n5492), .ZN(n5494)
         );
  INV_X1 U7030 ( .A(n5494), .ZN(n5495) );
  NAND2_X1 U7031 ( .A1(n8558), .A2(n8563), .ZN(n6180) );
  XOR2_X1 U7032 ( .A(n5496), .B(n6369), .Z(n5522) );
  INV_X1 U7033 ( .A(n5555), .ZN(n5499) );
  NAND2_X1 U7034 ( .A1(n5499), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5500) );
  OR2_X1 U7035 ( .A1(n5543), .A2(n7944), .ZN(n5508) );
  INV_X1 U7036 ( .A(n5501), .ZN(n5506) );
  NAND2_X1 U7037 ( .A1(n5506), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5503) );
  INV_X1 U7038 ( .A(n5498), .ZN(n5504) );
  NAND2_X1 U7039 ( .A1(n5504), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5505) );
  MUX2_X1 U7040 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5505), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n5507) );
  INV_X1 U7041 ( .A(n7687), .ZN(n5582) );
  NAND2_X1 U7042 ( .A1(n6144), .A2(n5582), .ZN(n6187) );
  INV_X1 U7043 ( .A(n6968), .ZN(n6953) );
  INV_X1 U7044 ( .A(n8529), .ZN(n5510) );
  NAND2_X1 U7045 ( .A1(n6953), .A2(n5510), .ZN(n5511) );
  AND2_X1 U7046 ( .A1(n5088), .A2(n5511), .ZN(n6911) );
  NAND2_X2 U7047 ( .A1(n6392), .A2(n6144), .ZN(n6322) );
  INV_X2 U7048 ( .A(n6322), .ZN(n6659) );
  INV_X1 U7049 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n5515) );
  NAND2_X1 U7050 ( .A1(n6161), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5513) );
  NAND2_X1 U7051 ( .A1(n6162), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5512) );
  OAI211_X1 U7052 ( .C1(n5515), .C2(n5514), .A(n5513), .B(n5512), .ZN(n5516)
         );
  INV_X1 U7053 ( .A(n5516), .ZN(n5517) );
  NOR2_X2 U7054 ( .A1(n6911), .A2(n6322), .ZN(n8728) );
  NAND2_X1 U7055 ( .A1(n5088), .A2(P2_B_REG_SCAN_IN), .ZN(n5518) );
  NAND2_X1 U7056 ( .A1(n8728), .A2(n5518), .ZN(n8548) );
  NAND2_X1 U7057 ( .A1(n6920), .A2(n7375), .ZN(n7042) );
  NAND2_X1 U7058 ( .A1(n7043), .A2(n7042), .ZN(n5526) );
  NAND2_X1 U7059 ( .A1(n7046), .A2(n7730), .ZN(n6346) );
  NAND2_X1 U7060 ( .A1(n6878), .A2(n5523), .ZN(n5524) );
  NAND2_X1 U7061 ( .A1(n6346), .A2(n5524), .ZN(n6194) );
  INV_X1 U7062 ( .A(n5523), .ZN(n7574) );
  NAND2_X1 U7063 ( .A1(n7630), .A2(n7574), .ZN(n5525) );
  NAND2_X1 U7064 ( .A1(n6194), .A2(n5525), .ZN(n6192) );
  NAND2_X1 U7065 ( .A1(n5526), .A2(n6192), .ZN(n6193) );
  INV_X1 U7066 ( .A(n6193), .ZN(n7627) );
  NAND2_X1 U7067 ( .A1(n7627), .A2(n5527), .ZN(n7626) );
  INV_X1 U7068 ( .A(n8370), .ZN(n7629) );
  NAND2_X1 U7069 ( .A1(n7629), .A2(n7924), .ZN(n6213) );
  NAND2_X1 U7070 ( .A1(n8370), .A2(n7699), .ZN(n6207) );
  NAND2_X1 U7071 ( .A1(n8369), .A2(n7743), .ZN(n6214) );
  NAND2_X1 U7072 ( .A1(n7614), .A2(n7542), .ZN(n6208) );
  NAND2_X1 U7073 ( .A1(n7688), .A2(n6208), .ZN(n7613) );
  NAND2_X1 U7074 ( .A1(n7642), .A2(n7585), .ZN(n7545) );
  NAND2_X1 U7075 ( .A1(n8368), .A2(n7721), .ZN(n6215) );
  NAND2_X1 U7076 ( .A1(n7613), .A2(n7612), .ZN(n7611) );
  NAND2_X1 U7077 ( .A1(n7864), .A2(n7645), .ZN(n6209) );
  AND2_X1 U7078 ( .A1(n7545), .A2(n6209), .ZN(n6220) );
  NAND2_X1 U7079 ( .A1(n7611), .A2(n6220), .ZN(n5528) );
  NAND2_X1 U7080 ( .A1(n8367), .A2(n7550), .ZN(n6218) );
  NAND2_X1 U7081 ( .A1(n5528), .A2(n6218), .ZN(n7522) );
  NAND2_X1 U7082 ( .A1(n7522), .A2(n6350), .ZN(n5529) );
  NAND2_X1 U7083 ( .A1(n8366), .A2(n7526), .ZN(n6228) );
  INV_X1 U7084 ( .A(n6229), .ZN(n5530) );
  AND2_X1 U7085 ( .A1(n8053), .A2(n8363), .ZN(n8028) );
  NAND2_X1 U7086 ( .A1(n7967), .A2(n8052), .ZN(n6353) );
  OR2_X1 U7087 ( .A1(n8053), .A2(n8363), .ZN(n7931) );
  AND2_X1 U7088 ( .A1(n6353), .A2(n7931), .ZN(n6243) );
  NAND2_X1 U7089 ( .A1(n5534), .A2(n6354), .ZN(n7972) );
  NAND2_X1 U7090 ( .A1(n7972), .A2(n7973), .ZN(n5535) );
  INV_X1 U7091 ( .A(n8077), .ZN(n8082) );
  INV_X1 U7092 ( .A(n8727), .ZN(n8150) );
  NAND2_X1 U7093 ( .A1(n8149), .A2(n8150), .ZN(n6259) );
  NAND2_X1 U7094 ( .A1(n5536), .A2(n6259), .ZN(n8722) );
  OR2_X1 U7095 ( .A1(n8792), .A2(n8217), .ZN(n6263) );
  NAND2_X1 U7096 ( .A1(n8722), .A2(n6263), .ZN(n5537) );
  NAND2_X1 U7097 ( .A1(n8792), .A2(n8217), .ZN(n6262) );
  NAND2_X1 U7098 ( .A1(n5537), .A2(n6262), .ZN(n8706) );
  INV_X1 U7099 ( .A(n6267), .ZN(n5538) );
  NAND2_X1 U7100 ( .A1(n8696), .A2(n6272), .ZN(n5539) );
  NAND2_X1 U7101 ( .A1(n5539), .A2(n6274), .ZN(n8685) );
  NOR2_X1 U7102 ( .A1(n8854), .A2(n8278), .ZN(n6343) );
  NAND2_X1 U7103 ( .A1(n8854), .A2(n8278), .ZN(n6341) );
  INV_X1 U7104 ( .A(n8689), .ZN(n8668) );
  OR2_X1 U7105 ( .A1(n8848), .A2(n8668), .ZN(n6280) );
  NAND2_X1 U7106 ( .A1(n8848), .A2(n8668), .ZN(n6287) );
  NAND2_X1 U7107 ( .A1(n8661), .A2(n6289), .ZN(n8648) );
  AND2_X1 U7108 ( .A1(n6294), .A2(n8647), .ZN(n6282) );
  NAND2_X1 U7109 ( .A1(n8648), .A2(n6282), .ZN(n5540) );
  NAND2_X1 U7110 ( .A1(n5540), .A2(n6290), .ZN(n8634) );
  INV_X1 U7111 ( .A(n6362), .ZN(n8637) );
  NOR2_X1 U7112 ( .A1(n8824), .A2(n8312), .ZN(n6339) );
  NAND2_X1 U7113 ( .A1(n8818), .A2(n8253), .ZN(n6335) );
  NAND2_X1 U7114 ( .A1(n8824), .A2(n8312), .ZN(n8617) );
  AND2_X2 U7115 ( .A1(n6335), .A2(n8617), .ZN(n6299) );
  INV_X1 U7116 ( .A(n5541), .ZN(n6306) );
  NOR2_X1 U7117 ( .A1(n5542), .A2(n8578), .ZN(n6310) );
  NAND2_X1 U7118 ( .A1(n5542), .A2(n8578), .ZN(n6308) );
  XNOR2_X1 U7119 ( .A(n6183), .B(n6369), .ZN(n8561) );
  NAND2_X1 U7120 ( .A1(n5543), .A2(n6392), .ZN(n6142) );
  NAND2_X1 U7121 ( .A1(n6144), .A2(n7687), .ZN(n7570) );
  AND2_X1 U7122 ( .A1(n7944), .A2(n7846), .ZN(n8793) );
  NAND2_X1 U7123 ( .A1(n6903), .A2(n6142), .ZN(n5544) );
  NAND2_X1 U7124 ( .A1(n8539), .A2(n7687), .ZN(n6383) );
  NOR2_X1 U7125 ( .A1(n8561), .A2(n8118), .ZN(n5545) );
  AND2_X1 U7126 ( .A1(n5554), .A2(n5579), .ZN(n5548) );
  NAND2_X1 U7127 ( .A1(n5555), .A2(n5548), .ZN(n5547) );
  AND2_X1 U7128 ( .A1(n5548), .A2(n5557), .ZN(n5549) );
  XNOR2_X1 U7129 ( .A(n8202), .B(P2_B_REG_SCAN_IN), .ZN(n5553) );
  NAND2_X1 U7130 ( .A1(n5555), .A2(n5554), .ZN(n5578) );
  NAND3_X1 U7131 ( .A1(n5557), .A2(n5579), .A3(n5556), .ZN(n5558) );
  OAI21_X2 U7132 ( .B1(n6782), .B2(P2_D_REG_0__SCAN_IN), .A(n6786), .ZN(n6905)
         );
  INV_X1 U7133 ( .A(n6905), .ZN(n5566) );
  NAND2_X1 U7134 ( .A1(n8129), .A2(n8069), .ZN(n6783) );
  INV_X1 U7135 ( .A(n7369), .ZN(n5565) );
  NOR2_X1 U7136 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n5570) );
  NOR4_X1 U7137 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5569) );
  NOR4_X1 U7138 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n5568) );
  NOR4_X1 U7139 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n5567) );
  NAND4_X1 U7140 ( .A1(n5570), .A2(n5569), .A3(n5568), .A4(n5567), .ZN(n5576)
         );
  NOR4_X1 U7141 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n5574) );
  NOR4_X1 U7142 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n5573) );
  NOR4_X1 U7143 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5572) );
  NOR4_X1 U7144 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n5571) );
  NAND4_X1 U7145 ( .A1(n5574), .A2(n5573), .A3(n5572), .A4(n5571), .ZN(n5575)
         );
  NOR2_X1 U7146 ( .A1(n5576), .A2(n5575), .ZN(n5577) );
  NAND2_X1 U7147 ( .A1(n6140), .A2(n6141), .ZN(n6862) );
  INV_X1 U7148 ( .A(n6862), .ZN(n5581) );
  NAND2_X1 U7149 ( .A1(n5578), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5580) );
  NAND2_X1 U7150 ( .A1(n5581), .A2(n6879), .ZN(n6883) );
  NAND2_X1 U7151 ( .A1(n7846), .A2(n5582), .ZN(n6904) );
  NOR2_X1 U7152 ( .A1(n7944), .A2(n6904), .ZN(n5583) );
  NAND2_X1 U7153 ( .A1(n8539), .A2(n5583), .ZN(n6863) );
  AND2_X1 U7154 ( .A1(n6875), .A2(n6863), .ZN(n5584) );
  OR2_X1 U7155 ( .A1(n6883), .A2(n5584), .ZN(n5587) );
  NAND3_X1 U7156 ( .A1(n6905), .A2(n7369), .A3(n6141), .ZN(n6872) );
  NAND2_X1 U7157 ( .A1(n6383), .A2(n8793), .ZN(n10061) );
  AND2_X1 U7158 ( .A1(n6322), .A2(n8745), .ZN(n5585) );
  NAND2_X1 U7159 ( .A1(n6863), .A2(n5585), .ZN(n6882) );
  NAND2_X1 U7160 ( .A1(n10061), .A2(n6882), .ZN(n6861) );
  NAND2_X1 U7161 ( .A1(n6885), .A2(n6861), .ZN(n5586) );
  INV_X1 U7162 ( .A(n8558), .ZN(n6150) );
  INV_X1 U7163 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U7164 ( .A1(n5589), .A2(n4906), .ZN(P2_U3456) );
  NAND2_X1 U7165 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5718) );
  INV_X1 U7166 ( .A(n5718), .ZN(n5590) );
  NAND2_X1 U7167 ( .A1(n5590), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5732) );
  INV_X1 U7168 ( .A(n5732), .ZN(n5591) );
  NAND2_X1 U7169 ( .A1(n5591), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5746) );
  INV_X1 U7170 ( .A(n5746), .ZN(n5592) );
  NAND2_X1 U7171 ( .A1(n5592), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5761) );
  INV_X1 U7172 ( .A(n5761), .ZN(n5593) );
  INV_X1 U7173 ( .A(n5852), .ZN(n5596) );
  INV_X1 U7174 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5865) );
  INV_X1 U7175 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5894) );
  INV_X1 U7176 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8957) );
  NAND2_X1 U7177 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(P1_REG3_REG_23__SCAN_IN), 
        .ZN(n5600) );
  INV_X1 U7178 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8919) );
  INV_X1 U7179 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5602) );
  NAND2_X1 U7180 ( .A1(n5975), .A2(n5602), .ZN(n5603) );
  NOR2_X1 U7181 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5608) );
  NOR2_X1 U7182 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5607) );
  NOR2_X1 U7183 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5606) );
  NOR2_X1 U7184 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5605) );
  NAND4_X1 U7185 ( .A1(n5611), .A2(n5610), .A3(n6010), .A4(n6009), .ZN(n5614)
         );
  NAND4_X1 U7186 ( .A1(n6008), .A2(n5612), .A3(n6016), .A4(n6067), .ZN(n5613)
         );
  NAND2_X1 U7187 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n5617) );
  OR2_X1 U7188 ( .A1(n5621), .A2(n4394), .ZN(n9724) );
  NAND2_X1 U7189 ( .A1(n9429), .A2(n5685), .ZN(n5633) );
  INV_X1 U7190 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n5630) );
  NAND2_X2 U7191 ( .A1(n8130), .A2(n5624), .ZN(n5683) );
  INV_X1 U7192 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n5625) );
  OR2_X1 U7193 ( .A1(n5683), .A2(n5625), .ZN(n5629) );
  INV_X1 U7194 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n5627) );
  OR2_X1 U7195 ( .A1(n5963), .A2(n5627), .ZN(n5628) );
  OAI211_X1 U7196 ( .C1(n5913), .C2(n5630), .A(n5629), .B(n5628), .ZN(n5631)
         );
  INV_X1 U7197 ( .A(n5631), .ZN(n5632) );
  NAND2_X1 U7198 ( .A1(n8059), .A2(n9014), .ZN(n5638) );
  INV_X1 U7199 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8060) );
  OR2_X1 U7200 ( .A1(n5673), .A2(n8060), .ZN(n5637) );
  NAND2_X1 U7201 ( .A1(n5684), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5645) );
  INV_X1 U7202 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5639) );
  NAND2_X1 U7203 ( .A1(n5852), .A2(n5639), .ZN(n5640) );
  AND2_X1 U7204 ( .A1(n5866), .A2(n5640), .ZN(n9005) );
  NAND2_X1 U7205 ( .A1(n5685), .A2(n9005), .ZN(n5644) );
  INV_X1 U7206 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9853) );
  OR2_X1 U7207 ( .A1(n5683), .A2(n9853), .ZN(n5643) );
  INV_X1 U7208 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n5641) );
  OR2_X1 U7209 ( .A1(n5963), .A2(n5641), .ZN(n5642) );
  NAND4_X1 U7210 ( .A1(n5645), .A2(n5644), .A3(n5643), .A4(n5642), .ZN(n9587)
         );
  INV_X1 U7211 ( .A(n9587), .ZN(n8930) );
  NAND2_X1 U7212 ( .A1(n6857), .A2(n9014), .ZN(n5649) );
  NAND2_X1 U7213 ( .A1(n5873), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5646) );
  MUX2_X1 U7214 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5646), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n5647) );
  OR2_X1 U7215 ( .A1(n5873), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n5861) );
  NAND2_X1 U7216 ( .A1(n5647), .A2(n5861), .ZN(n9368) );
  INV_X1 U7217 ( .A(n9368), .ZN(n9860) );
  AOI22_X1 U7218 ( .A1(n5904), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5903), .B2(
        n9860), .ZN(n5648) );
  INV_X1 U7219 ( .A(n9672), .ZN(n9009) );
  INV_X1 U7220 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n5650) );
  NAND2_X1 U7221 ( .A1(n5684), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5654) );
  INV_X1 U7222 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5651) );
  INV_X1 U7223 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5657) );
  NAND2_X1 U7224 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5656) );
  XNOR2_X1 U7225 ( .A(n5657), .B(n5656), .ZN(n6753) );
  XNOR2_X2 U7226 ( .A(n6417), .B(n6060), .ZN(n6848) );
  INV_X1 U7227 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n5659) );
  NAND2_X1 U7228 ( .A1(n5685), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5660) );
  NAND2_X1 U7229 ( .A1(n5661), .A2(n5660), .ZN(n5666) );
  INV_X1 U7230 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5662) );
  OR2_X1 U7231 ( .A1(n5701), .A2(n5662), .ZN(n5664) );
  NAND2_X1 U7232 ( .A1(n5684), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5663) );
  NAND2_X1 U7233 ( .A1(n5664), .A2(n5663), .ZN(n5665) );
  INV_X1 U7234 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9789) );
  NAND2_X1 U7235 ( .A1(n4350), .A2(SI_0_), .ZN(n5668) );
  INV_X1 U7236 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5667) );
  NAND2_X1 U7237 ( .A1(n5668), .A2(n5667), .ZN(n5670) );
  NAND2_X1 U7238 ( .A1(n5670), .A2(n5669), .ZN(n9733) );
  MUX2_X1 U7239 ( .A(n9789), .B(n9733), .S(n5675), .Z(n6813) );
  NAND2_X1 U7240 ( .A1(n6713), .A2(n6843), .ZN(n6842) );
  OR2_X1 U7241 ( .A1(n5672), .A2(n5800), .ZN(n5709) );
  INV_X1 U7242 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5691) );
  XNOR2_X1 U7243 ( .A(n5709), .B(n5691), .ZN(n6752) );
  OR2_X1 U7244 ( .A1(n5887), .A2(n6672), .ZN(n5674) );
  INV_X1 U7245 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6673) );
  NAND2_X1 U7246 ( .A1(n5684), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5679) );
  NAND2_X1 U7247 ( .A1(n5685), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5678) );
  INV_X1 U7248 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5676) );
  OR2_X1 U7249 ( .A1(n5701), .A2(n5676), .ZN(n5677) );
  XNOR2_X1 U7250 ( .A(n9965), .B(n9284), .ZN(n7081) );
  NAND2_X1 U7251 ( .A1(n7082), .A2(n7081), .ZN(n7080) );
  INV_X1 U7252 ( .A(n9284), .ZN(n6850) );
  NAND2_X1 U7253 ( .A1(n6850), .A2(n9965), .ZN(n5681) );
  NAND2_X1 U7254 ( .A1(n7080), .A2(n5681), .ZN(n7052) );
  INV_X1 U7255 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n5682) );
  NAND2_X1 U7256 ( .A1(n5684), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5687) );
  INV_X1 U7257 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9951) );
  NAND2_X1 U7258 ( .A1(n5685), .A2(n9951), .ZN(n5686) );
  NAND2_X1 U7259 ( .A1(n5709), .A2(n5691), .ZN(n5692) );
  NAND2_X1 U7260 ( .A1(n5692), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5694) );
  INV_X1 U7261 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5693) );
  XNOR2_X1 U7262 ( .A(n5694), .B(n5693), .ZN(n6756) );
  OR2_X1 U7263 ( .A1(n5887), .A2(n6674), .ZN(n5696) );
  INV_X1 U7264 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6675) );
  OR2_X1 U7265 ( .A1(n5673), .A2(n6675), .ZN(n5695) );
  NAND2_X1 U7266 ( .A1(n9283), .A2(n9956), .ZN(n9208) );
  NAND2_X1 U7267 ( .A1(n6026), .A2(n9208), .ZN(n9023) );
  NAND2_X1 U7268 ( .A1(n7052), .A2(n9023), .ZN(n7051) );
  NAND2_X1 U7269 ( .A1(n7077), .A2(n9956), .ZN(n5697) );
  NAND2_X1 U7270 ( .A1(n7051), .A2(n5697), .ZN(n7065) );
  INV_X1 U7271 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5698) );
  OR2_X1 U7272 ( .A1(n5683), .A2(n5698), .ZN(n5706) );
  INV_X1 U7273 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5699) );
  NAND2_X1 U7274 ( .A1(n9951), .A2(n5699), .ZN(n5700) );
  AND2_X1 U7275 ( .A1(n5700), .A2(n5718), .ZN(n7068) );
  NAND2_X1 U7276 ( .A1(n5685), .A2(n7068), .ZN(n5705) );
  NAND2_X1 U7277 ( .A1(n5684), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5704) );
  INV_X1 U7278 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5702) );
  OR2_X1 U7279 ( .A1(n5963), .A2(n5702), .ZN(n5703) );
  NAND4_X1 U7280 ( .A1(n5706), .A2(n5705), .A3(n5704), .A4(n5703), .ZN(n9282)
         );
  INV_X1 U7281 ( .A(n9282), .ZN(n6939) );
  OR2_X1 U7282 ( .A1(n5707), .A2(n5800), .ZN(n5708) );
  AND2_X1 U7283 ( .A1(n5709), .A2(n5708), .ZN(n5711) );
  INV_X1 U7284 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5710) );
  NAND2_X1 U7285 ( .A1(n5711), .A2(n5710), .ZN(n5725) );
  INV_X1 U7286 ( .A(n5711), .ZN(n5712) );
  NAND2_X1 U7287 ( .A1(n5712), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5713) );
  NAND2_X1 U7288 ( .A1(n5725), .A2(n5713), .ZN(n9312) );
  OR2_X1 U7289 ( .A1(n5887), .A2(n6670), .ZN(n5715) );
  INV_X1 U7290 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6671) );
  OR2_X1 U7291 ( .A1(n5673), .A2(n6671), .ZN(n5714) );
  OAI211_X1 U7292 ( .C1(n6686), .C2(n9312), .A(n5715), .B(n5714), .ZN(n7069)
         );
  NAND2_X1 U7293 ( .A1(n6939), .A2(n7069), .ZN(n9048) );
  INV_X1 U7294 ( .A(n7069), .ZN(n9970) );
  NAND2_X1 U7295 ( .A1(n9282), .A2(n9970), .ZN(n9215) );
  NAND2_X1 U7296 ( .A1(n9048), .A2(n9215), .ZN(n9020) );
  NAND2_X1 U7297 ( .A1(n7065), .A2(n9020), .ZN(n7064) );
  NAND2_X1 U7298 ( .A1(n6939), .A2(n9970), .ZN(n5716) );
  NAND2_X1 U7299 ( .A1(n7064), .A2(n5716), .ZN(n6894) );
  NAND2_X1 U7300 ( .A1(n5684), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5724) );
  INV_X1 U7301 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5717) );
  NAND2_X1 U7302 ( .A1(n5718), .A2(n5717), .ZN(n5719) );
  AND2_X1 U7303 ( .A1(n5732), .A2(n5719), .ZN(n6936) );
  NAND2_X1 U7304 ( .A1(n5685), .A2(n6936), .ZN(n5723) );
  INV_X1 U7305 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6760) );
  OR2_X1 U7306 ( .A1(n5683), .A2(n6760), .ZN(n5722) );
  INV_X1 U7307 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5720) );
  OR2_X1 U7308 ( .A1(n5963), .A2(n5720), .ZN(n5721) );
  NAND4_X1 U7309 ( .A1(n5724), .A2(n5723), .A3(n5722), .A4(n5721), .ZN(n9281)
         );
  INV_X1 U7310 ( .A(n9281), .ZN(n7107) );
  NAND2_X1 U7311 ( .A1(n5725), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5727) );
  INV_X1 U7312 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5726) );
  XNOR2_X1 U7313 ( .A(n5727), .B(n5726), .ZN(n6761) );
  OR2_X1 U7314 ( .A1(n6682), .A2(n5887), .ZN(n5729) );
  INV_X1 U7315 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6683) );
  OR2_X1 U7316 ( .A1(n5673), .A2(n6683), .ZN(n5728) );
  OAI211_X1 U7317 ( .C1(n6686), .C2(n6761), .A(n5729), .B(n5728), .ZN(n6941)
         );
  NAND2_X1 U7318 ( .A1(n7107), .A2(n6941), .ZN(n9057) );
  NAND2_X1 U7319 ( .A1(n9281), .A2(n7099), .ZN(n9217) );
  NAND2_X1 U7320 ( .A1(n9057), .A2(n9217), .ZN(n9019) );
  NAND2_X1 U7321 ( .A1(n7107), .A2(n7099), .ZN(n5730) );
  INV_X1 U7322 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5731) );
  NAND2_X1 U7323 ( .A1(n5732), .A2(n5731), .ZN(n5733) );
  AND2_X1 U7324 ( .A1(n5746), .A2(n5733), .ZN(n7112) );
  NAND2_X1 U7325 ( .A1(n5685), .A2(n7112), .ZN(n5738) );
  NAND2_X1 U7326 ( .A1(n5684), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5737) );
  INV_X1 U7327 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6763) );
  OR2_X1 U7328 ( .A1(n5683), .A2(n6763), .ZN(n5736) );
  INV_X1 U7329 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5734) );
  OR2_X1 U7330 ( .A1(n5963), .A2(n5734), .ZN(n5735) );
  NAND4_X1 U7331 ( .A1(n5738), .A2(n5737), .A3(n5736), .A4(n5735), .ZN(n9280)
         );
  OR2_X1 U7332 ( .A1(n6678), .A2(n5887), .ZN(n5745) );
  NAND2_X1 U7333 ( .A1(n5739), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5740) );
  MUX2_X1 U7334 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5740), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n5743) );
  AND2_X1 U7335 ( .A1(n5743), .A2(n5742), .ZN(n6764) );
  AOI22_X1 U7336 ( .A1(n5904), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5903), .B2(
        n6764), .ZN(n5744) );
  NAND2_X1 U7337 ( .A1(n5745), .A2(n5744), .ZN(n7113) );
  NAND2_X1 U7338 ( .A1(n7478), .A2(n7113), .ZN(n9062) );
  INV_X1 U7339 ( .A(n7113), .ZN(n9975) );
  NAND2_X1 U7340 ( .A1(n9280), .A2(n9975), .ZN(n9049) );
  NAND2_X1 U7341 ( .A1(n9062), .A2(n9049), .ZN(n7109) );
  NAND2_X1 U7342 ( .A1(n5684), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5753) );
  INV_X1 U7343 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n7135) );
  NAND2_X1 U7344 ( .A1(n5746), .A2(n7135), .ZN(n5747) );
  AND2_X1 U7345 ( .A1(n5761), .A2(n5747), .ZN(n7480) );
  NAND2_X1 U7346 ( .A1(n5685), .A2(n7480), .ZN(n5752) );
  INV_X1 U7347 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n5748) );
  OR2_X1 U7348 ( .A1(n5683), .A2(n5748), .ZN(n5751) );
  INV_X1 U7349 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n5749) );
  OR2_X1 U7350 ( .A1(n5963), .A2(n5749), .ZN(n5750) );
  NAND4_X1 U7351 ( .A1(n5753), .A2(n5752), .A3(n5751), .A4(n5750), .ZN(n9931)
         );
  NAND2_X1 U7352 ( .A1(n5742), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5754) );
  XNOR2_X1 U7353 ( .A(n5754), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9341) );
  AOI22_X1 U7354 ( .A1(n5904), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5903), .B2(
        n9341), .ZN(n5755) );
  OR2_X1 U7355 ( .A1(n7681), .A2(n7598), .ZN(n9064) );
  NAND2_X1 U7356 ( .A1(n7681), .A2(n7598), .ZN(n9925) );
  NAND2_X1 U7357 ( .A1(n9064), .A2(n9925), .ZN(n7475) );
  NAND2_X1 U7358 ( .A1(n7471), .A2(n7475), .ZN(n7473) );
  NAND2_X1 U7359 ( .A1(n5756), .A2(n7681), .ZN(n5757) );
  NOR2_X1 U7360 ( .A1(n5742), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5786) );
  OR2_X1 U7361 ( .A1(n5786), .A2(n5800), .ZN(n5771) );
  XNOR2_X1 U7362 ( .A(n5771), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6767) );
  AOI22_X1 U7363 ( .A1(n5904), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5903), .B2(
        n6767), .ZN(n5758) );
  NAND2_X1 U7364 ( .A1(n5684), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5768) );
  INV_X1 U7365 ( .A(n5759), .ZN(n5777) );
  INV_X1 U7366 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5760) );
  NAND2_X1 U7367 ( .A1(n5761), .A2(n5760), .ZN(n5762) );
  AND2_X1 U7368 ( .A1(n5777), .A2(n5762), .ZN(n9938) );
  NAND2_X1 U7369 ( .A1(n5685), .A2(n9938), .ZN(n5767) );
  INV_X1 U7370 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n5763) );
  OR2_X1 U7371 ( .A1(n5683), .A2(n5763), .ZN(n5766) );
  INV_X1 U7372 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5764) );
  OR2_X1 U7373 ( .A1(n5963), .A2(n5764), .ZN(n5765) );
  NAND4_X1 U7374 ( .A1(n5768), .A2(n5767), .A3(n5766), .A4(n5765), .ZN(n9922)
         );
  NAND2_X1 U7375 ( .A1(n9940), .A2(n9922), .ZN(n5769) );
  INV_X1 U7376 ( .A(n9940), .ZN(n9981) );
  INV_X1 U7377 ( .A(n9922), .ZN(n7836) );
  NAND2_X1 U7378 ( .A1(n6697), .A2(n9014), .ZN(n5775) );
  INV_X1 U7379 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5770) );
  NAND2_X1 U7380 ( .A1(n5771), .A2(n5770), .ZN(n5772) );
  NAND2_X1 U7381 ( .A1(n5772), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5773) );
  XNOR2_X1 U7382 ( .A(n5773), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9764) );
  AOI22_X1 U7383 ( .A1(n5904), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5903), .B2(
        n9764), .ZN(n5774) );
  NAND2_X1 U7384 ( .A1(n5684), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5784) );
  INV_X1 U7385 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5776) );
  NAND2_X1 U7386 ( .A1(n5777), .A2(n5776), .ZN(n5778) );
  AND2_X1 U7387 ( .A1(n5791), .A2(n5778), .ZN(n7839) );
  NAND2_X1 U7388 ( .A1(n5685), .A2(n7839), .ZN(n5783) );
  INV_X1 U7389 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5779) );
  OR2_X1 U7390 ( .A1(n5683), .A2(n5779), .ZN(n5782) );
  INV_X1 U7391 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n5780) );
  OR2_X1 U7392 ( .A1(n5963), .A2(n5780), .ZN(n5781) );
  NAND4_X1 U7393 ( .A1(n5784), .A2(n5783), .A3(n5782), .A4(n5781), .ZN(n9930)
         );
  INV_X1 U7394 ( .A(n9930), .ZN(n7801) );
  AND2_X1 U7395 ( .A1(n7512), .A2(n7801), .ZN(n6030) );
  NOR2_X1 U7396 ( .A1(n6029), .A2(n6030), .ZN(n7518) );
  NOR2_X1 U7397 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5785) );
  AND2_X1 U7398 ( .A1(n5786), .A2(n5785), .ZN(n5799) );
  OR2_X1 U7399 ( .A1(n5799), .A2(n5800), .ZN(n5787) );
  XNOR2_X1 U7400 ( .A(n5787), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6770) );
  AOI22_X1 U7401 ( .A1(n5904), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5903), .B2(
        n6770), .ZN(n5788) );
  NAND2_X1 U7402 ( .A1(n5684), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5797) );
  INV_X1 U7403 ( .A(n5789), .ZN(n5805) );
  INV_X1 U7404 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5790) );
  NAND2_X1 U7405 ( .A1(n5791), .A2(n5790), .ZN(n5792) );
  AND2_X1 U7406 ( .A1(n5805), .A2(n5792), .ZN(n7803) );
  NAND2_X1 U7407 ( .A1(n5685), .A2(n7803), .ZN(n5796) );
  INV_X1 U7408 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6750) );
  OR2_X1 U7409 ( .A1(n5683), .A2(n6750), .ZN(n5795) );
  INV_X1 U7410 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5793) );
  OR2_X1 U7411 ( .A1(n5963), .A2(n5793), .ZN(n5794) );
  NAND4_X1 U7412 ( .A1(n5797), .A2(n5796), .A3(n5795), .A4(n5794), .ZN(n9279)
         );
  INV_X1 U7413 ( .A(n9279), .ZN(n7879) );
  OR2_X1 U7414 ( .A1(n7391), .A2(n7879), .ZN(n9080) );
  NAND2_X1 U7415 ( .A1(n7391), .A2(n7879), .ZN(n9076) );
  INV_X1 U7416 ( .A(n7391), .ZN(n9993) );
  NAND2_X1 U7417 ( .A1(n6705), .A2(n9014), .ZN(n5803) );
  INV_X1 U7418 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5798) );
  AND2_X1 U7419 ( .A1(n5799), .A2(n5798), .ZN(n5814) );
  OR2_X1 U7420 ( .A1(n5814), .A2(n5800), .ZN(n5801) );
  XNOR2_X1 U7421 ( .A(n5801), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6772) );
  AOI22_X1 U7422 ( .A1(n5904), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5903), .B2(
        n6772), .ZN(n5802) );
  INV_X1 U7423 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5804) );
  NAND2_X1 U7424 ( .A1(n5805), .A2(n5804), .ZN(n5806) );
  AND2_X1 U7425 ( .A1(n5820), .A2(n5806), .ZN(n7881) );
  NAND2_X1 U7426 ( .A1(n5685), .A2(n7881), .ZN(n5811) );
  NAND2_X1 U7427 ( .A1(n5684), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5810) );
  INV_X1 U7428 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6771) );
  OR2_X1 U7429 ( .A1(n5683), .A2(n6771), .ZN(n5809) );
  INV_X1 U7430 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n5807) );
  OR2_X1 U7431 ( .A1(n5963), .A2(n5807), .ZN(n5808) );
  NAND4_X1 U7432 ( .A1(n5811), .A2(n5810), .A3(n5809), .A4(n5808), .ZN(n9910)
         );
  INV_X1 U7433 ( .A(n9910), .ZN(n5812) );
  NAND2_X1 U7434 ( .A1(n7882), .A2(n5812), .ZN(n9082) );
  OR2_X1 U7435 ( .A1(n6732), .A2(n5887), .ZN(n5818) );
  INV_X1 U7436 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5813) );
  NAND2_X1 U7437 ( .A1(n5814), .A2(n5813), .ZN(n5844) );
  NAND2_X1 U7438 ( .A1(n5844), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5815) );
  INV_X1 U7439 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5842) );
  NAND2_X1 U7440 ( .A1(n5815), .A2(n5842), .ZN(n5828) );
  OR2_X1 U7441 ( .A1(n5815), .A2(n5842), .ZN(n5816) );
  AOI22_X1 U7442 ( .A1(n5904), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5903), .B2(
        n9366), .ZN(n5817) );
  NAND2_X1 U7443 ( .A1(n5684), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5827) );
  NAND2_X1 U7444 ( .A1(n5820), .A2(n5819), .ZN(n5821) );
  AND2_X1 U7445 ( .A1(n5833), .A2(n5821), .ZN(n9913) );
  NAND2_X1 U7446 ( .A1(n5685), .A2(n9913), .ZN(n5826) );
  INV_X1 U7447 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n5822) );
  OR2_X1 U7448 ( .A1(n5683), .A2(n5822), .ZN(n5825) );
  INV_X1 U7449 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n5823) );
  OR2_X1 U7450 ( .A1(n5963), .A2(n5823), .ZN(n5824) );
  NAND4_X1 U7451 ( .A1(n5827), .A2(n5826), .A3(n5825), .A4(n5824), .ZN(n9278)
         );
  NAND2_X1 U7452 ( .A1(n9914), .A2(n7852), .ZN(n9224) );
  NAND2_X1 U7453 ( .A1(n9085), .A2(n9224), .ZN(n9915) );
  NAND2_X1 U7454 ( .A1(n6809), .A2(n9014), .ZN(n5831) );
  NAND2_X1 U7455 ( .A1(n5828), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5829) );
  XNOR2_X1 U7456 ( .A(n5829), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9830) );
  AOI22_X1 U7457 ( .A1(n5904), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5903), .B2(
        n9830), .ZN(n5830) );
  NAND2_X1 U7458 ( .A1(n5684), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5839) );
  NAND2_X1 U7459 ( .A1(n5833), .A2(n5832), .ZN(n5834) );
  AND2_X1 U7460 ( .A1(n5850), .A2(n5834), .ZN(n7854) );
  NAND2_X1 U7461 ( .A1(n5685), .A2(n7854), .ZN(n5838) );
  INV_X1 U7462 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9364) );
  OR2_X1 U7463 ( .A1(n5683), .A2(n9364), .ZN(n5837) );
  INV_X1 U7464 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n5835) );
  OR2_X1 U7465 ( .A1(n5963), .A2(n5835), .ZN(n5836) );
  NAND4_X1 U7466 ( .A1(n5839), .A2(n5838), .A3(n5837), .A4(n5836), .ZN(n9909)
         );
  INV_X1 U7467 ( .A(n9909), .ZN(n7988) );
  OR2_X1 U7468 ( .A1(n6499), .A2(n7988), .ZN(n9227) );
  NAND2_X1 U7469 ( .A1(n6499), .A2(n7988), .ZN(n9230) );
  OAI21_X1 U7470 ( .B1(n7770), .B2(n9034), .A(n5840), .ZN(n7909) );
  NAND2_X1 U7471 ( .A1(n6838), .A2(n9014), .ZN(n5848) );
  INV_X1 U7472 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5841) );
  NAND2_X1 U7473 ( .A1(n5842), .A2(n5841), .ZN(n5843) );
  OAI21_X1 U7474 ( .B1(n5844), .B2(n5843), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5845) );
  MUX2_X1 U7475 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5845), .S(
        P1_IR_REG_14__SCAN_IN), .Z(n5846) );
  AND2_X1 U7476 ( .A1(n5846), .A2(n5873), .ZN(n9835) );
  AOI22_X1 U7477 ( .A1(n5904), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5903), .B2(
        n9835), .ZN(n5847) );
  NAND2_X1 U7478 ( .A1(n5684), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5858) );
  INV_X1 U7479 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5849) );
  NAND2_X1 U7480 ( .A1(n5850), .A2(n5849), .ZN(n5851) );
  AND2_X1 U7481 ( .A1(n5852), .A2(n5851), .ZN(n7992) );
  NAND2_X1 U7482 ( .A1(n5685), .A2(n7992), .ZN(n5857) );
  INV_X1 U7483 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n5853) );
  OR2_X1 U7484 ( .A1(n5683), .A2(n5853), .ZN(n5856) );
  INV_X1 U7485 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n5854) );
  OR2_X1 U7486 ( .A1(n5963), .A2(n5854), .ZN(n5855) );
  NAND4_X1 U7487 ( .A1(n5858), .A2(n5857), .A3(n5856), .A4(n5855), .ZN(n9277)
         );
  NOR2_X1 U7488 ( .A1(n9679), .A2(n9277), .ZN(n5859) );
  INV_X1 U7489 ( .A(n9679), .ZN(n7989) );
  AOI21_X1 U7490 ( .B1(n9672), .B2(n9587), .A(n8009), .ZN(n5860) );
  AOI21_X1 U7491 ( .B1(n8930), .B2(n9009), .A(n5860), .ZN(n9582) );
  NAND2_X1 U7492 ( .A1(n6926), .A2(n9014), .ZN(n5864) );
  NAND2_X1 U7493 ( .A1(n5861), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5862) );
  XNOR2_X1 U7494 ( .A(n5862), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9874) );
  AOI22_X1 U7495 ( .A1(n5904), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5903), .B2(
        n9874), .ZN(n5863) );
  NAND2_X1 U7496 ( .A1(n5684), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5872) );
  NAND2_X1 U7497 ( .A1(n5866), .A2(n5865), .ZN(n5867) );
  AND2_X1 U7498 ( .A1(n5878), .A2(n5867), .ZN(n9592) );
  NAND2_X1 U7499 ( .A1(n5685), .A2(n9592), .ZN(n5871) );
  INV_X1 U7500 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9363) );
  OR2_X1 U7501 ( .A1(n5683), .A2(n9363), .ZN(n5870) );
  INV_X1 U7502 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n5868) );
  OR2_X1 U7503 ( .A1(n5963), .A2(n5868), .ZN(n5869) );
  NAND4_X1 U7504 ( .A1(n5872), .A2(n5871), .A3(n5870), .A4(n5869), .ZN(n9575)
         );
  INV_X1 U7505 ( .A(n9575), .ZN(n8939) );
  OR2_X1 U7506 ( .A1(n9667), .A2(n8939), .ZN(n9232) );
  NAND2_X1 U7507 ( .A1(n9667), .A2(n8939), .ZN(n9237) );
  NAND2_X1 U7508 ( .A1(n9232), .A2(n9237), .ZN(n9581) );
  NAND2_X1 U7509 ( .A1(n9582), .A2(n9581), .ZN(n9580) );
  NAND2_X1 U7510 ( .A1(n9580), .A2(n4904), .ZN(n9565) );
  NAND2_X1 U7511 ( .A1(n7103), .A2(n9014), .ZN(n5876) );
  INV_X1 U7512 ( .A(n5873), .ZN(n5874) );
  NAND2_X1 U7513 ( .A1(n5874), .A2(n4912), .ZN(n6007) );
  XNOR2_X1 U7514 ( .A(n5888), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9883) );
  AOI22_X1 U7515 ( .A1(n5904), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5903), .B2(
        n9883), .ZN(n5875) );
  NAND2_X2 U7516 ( .A1(n5876), .A2(n5875), .ZN(n9662) );
  INV_X1 U7517 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5877) );
  NAND2_X1 U7518 ( .A1(n5878), .A2(n5877), .ZN(n5879) );
  AND2_X1 U7519 ( .A1(n5895), .A2(n5879), .ZN(n9568) );
  NAND2_X1 U7520 ( .A1(n9568), .A2(n5685), .ZN(n5884) );
  INV_X1 U7521 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9371) );
  OR2_X1 U7522 ( .A1(n5683), .A2(n9371), .ZN(n5883) );
  NAND2_X1 U7523 ( .A1(n5684), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5882) );
  INV_X1 U7524 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n5880) );
  OR2_X1 U7525 ( .A1(n5963), .A2(n5880), .ZN(n5881) );
  NAND4_X1 U7526 ( .A1(n5884), .A2(n5883), .A3(n5882), .A4(n5881), .ZN(n9586)
         );
  INV_X1 U7527 ( .A(n9586), .ZN(n6037) );
  NAND2_X1 U7528 ( .A1(n9570), .A2(n6037), .ZN(n5886) );
  NAND2_X1 U7529 ( .A1(n5888), .A2(n6009), .ZN(n5889) );
  NAND2_X1 U7530 ( .A1(n5889), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5890) );
  NAND2_X1 U7531 ( .A1(n5890), .A2(n6010), .ZN(n5901) );
  OR2_X1 U7532 ( .A1(n5890), .A2(n6010), .ZN(n5891) );
  AND2_X1 U7533 ( .A1(n5901), .A2(n5891), .ZN(n9372) );
  AOI22_X1 U7534 ( .A1(n5904), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5903), .B2(
        n9372), .ZN(n5892) );
  NAND2_X1 U7535 ( .A1(n5895), .A2(n5894), .ZN(n5896) );
  NAND2_X1 U7536 ( .A1(n5908), .A2(n5896), .ZN(n9552) );
  AOI22_X1 U7537 ( .A1(n5684), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n5897), .B2(
        P1_REG1_REG_18__SCAN_IN), .ZN(n5900) );
  INV_X1 U7538 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n5898) );
  OR2_X1 U7539 ( .A1(n5963), .A2(n5898), .ZN(n5899) );
  OAI211_X1 U7540 ( .C1(n9552), .C2(n6050), .A(n5900), .B(n5899), .ZN(n9574)
         );
  INV_X1 U7541 ( .A(n9574), .ZN(n9102) );
  INV_X1 U7542 ( .A(n9657), .ZN(n9555) );
  NAND2_X1 U7543 ( .A1(n7553), .A2(n9014), .ZN(n5906) );
  XNOR2_X2 U7544 ( .A(n5902), .B(P1_IR_REG_19__SCAN_IN), .ZN(n6096) );
  AOI22_X1 U7545 ( .A1(n5904), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n6096), .B2(
        n5903), .ZN(n5905) );
  INV_X1 U7546 ( .A(n9652), .ZN(n9542) );
  INV_X1 U7547 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n5912) );
  INV_X1 U7548 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5907) );
  NAND2_X1 U7549 ( .A1(n5908), .A2(n5907), .ZN(n5909) );
  NAND2_X1 U7550 ( .A1(n5916), .A2(n5909), .ZN(n9539) );
  OR2_X1 U7551 ( .A1(n9539), .A2(n6050), .ZN(n5911) );
  AOI22_X1 U7552 ( .A1(n5918), .A2(P1_REG0_REG_19__SCAN_IN), .B1(n5897), .B2(
        P1_REG1_REG_19__SCAN_IN), .ZN(n5910) );
  OAI211_X1 U7553 ( .C1(n5913), .C2(n5912), .A(n5911), .B(n5910), .ZN(n9559)
         );
  INV_X1 U7554 ( .A(n9559), .ZN(n9112) );
  NAND2_X1 U7555 ( .A1(n7674), .A2(n9014), .ZN(n5915) );
  INV_X1 U7556 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7675) );
  OR2_X1 U7557 ( .A1(n5673), .A2(n7675), .ZN(n5914) );
  NAND2_X1 U7558 ( .A1(n5916), .A2(n8957), .ZN(n5917) );
  NAND2_X1 U7559 ( .A1(n5925), .A2(n5917), .ZN(n9526) );
  AOI22_X1 U7560 ( .A1(n5918), .A2(P1_REG0_REG_20__SCAN_IN), .B1(n5897), .B2(
        P1_REG1_REG_20__SCAN_IN), .ZN(n5920) );
  NAND2_X1 U7561 ( .A1(n5684), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5919) );
  OAI211_X1 U7562 ( .C1(n9526), .C2(n6050), .A(n5920), .B(n5919), .ZN(n9546)
         );
  NAND2_X1 U7563 ( .A1(n9647), .A2(n9546), .ZN(n5921) );
  INV_X1 U7564 ( .A(n9647), .ZN(n9529) );
  INV_X1 U7565 ( .A(n9546), .ZN(n8903) );
  NAND2_X1 U7566 ( .A1(n7842), .A2(n9014), .ZN(n5923) );
  INV_X1 U7567 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7843) );
  OR2_X1 U7568 ( .A1(n5673), .A2(n7843), .ZN(n5922) );
  INV_X1 U7569 ( .A(n9513), .ZN(n9710) );
  INV_X1 U7570 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5924) );
  NAND2_X1 U7571 ( .A1(n5925), .A2(n5924), .ZN(n5926) );
  NAND2_X1 U7572 ( .A1(n5948), .A2(n5926), .ZN(n9516) );
  OR2_X1 U7573 ( .A1(n9516), .A2(n6050), .ZN(n5931) );
  INV_X1 U7574 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9514) );
  INV_X1 U7575 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9707) );
  OR2_X1 U7576 ( .A1(n5963), .A2(n9707), .ZN(n5928) );
  INV_X1 U7577 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9643) );
  OR2_X1 U7578 ( .A1(n5683), .A2(n9643), .ZN(n5927) );
  OAI211_X1 U7579 ( .C1(n5913), .C2(n9514), .A(n5928), .B(n5927), .ZN(n5929)
         );
  INV_X1 U7580 ( .A(n5929), .ZN(n5930) );
  NAND2_X1 U7581 ( .A1(n5931), .A2(n5930), .ZN(n9533) );
  INV_X1 U7582 ( .A(n9533), .ZN(n8958) );
  NAND2_X1 U7583 ( .A1(n9710), .A2(n8958), .ZN(n5932) );
  NAND2_X1 U7584 ( .A1(n7939), .A2(n9014), .ZN(n5934) );
  INV_X1 U7585 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7940) );
  OR2_X1 U7586 ( .A1(n5673), .A2(n7940), .ZN(n5933) );
  XNOR2_X1 U7587 ( .A(n5948), .B(P1_REG3_REG_22__SCAN_IN), .ZN(n9493) );
  NAND2_X1 U7588 ( .A1(n9493), .A2(n5685), .ZN(n5942) );
  INV_X1 U7589 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n5939) );
  INV_X1 U7590 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n5935) );
  OR2_X1 U7591 ( .A1(n5683), .A2(n5935), .ZN(n5938) );
  INV_X1 U7592 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n5936) );
  OR2_X1 U7593 ( .A1(n5963), .A2(n5936), .ZN(n5937) );
  OAI211_X1 U7594 ( .C1(n5913), .C2(n5939), .A(n5938), .B(n5937), .ZN(n5940)
         );
  INV_X1 U7595 ( .A(n5940), .ZN(n5941) );
  NAND2_X1 U7596 ( .A1(n5942), .A2(n5941), .ZN(n9507) );
  NAND2_X1 U7597 ( .A1(n9636), .A2(n9507), .ZN(n5943) );
  NAND2_X1 U7598 ( .A1(n7949), .A2(n9014), .ZN(n5945) );
  INV_X1 U7599 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7951) );
  OR2_X1 U7600 ( .A1(n5673), .A2(n7951), .ZN(n5944) );
  INV_X1 U7601 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5947) );
  INV_X1 U7602 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5946) );
  OAI21_X1 U7603 ( .B1(n5948), .B2(n5947), .A(n5946), .ZN(n5949) );
  NAND2_X1 U7604 ( .A1(n5949), .A2(n5960), .ZN(n9475) );
  OR2_X1 U7605 ( .A1(n9475), .A2(n6050), .ZN(n5954) );
  INV_X1 U7606 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9484) );
  INV_X1 U7607 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9702) );
  OR2_X1 U7608 ( .A1(n5963), .A2(n9702), .ZN(n5951) );
  INV_X1 U7609 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9633) );
  OR2_X1 U7610 ( .A1(n5683), .A2(n9633), .ZN(n5950) );
  OAI211_X1 U7611 ( .C1(n5913), .C2(n9484), .A(n5951), .B(n5950), .ZN(n5952)
         );
  INV_X1 U7612 ( .A(n5952), .ZN(n5953) );
  NAND2_X1 U7613 ( .A1(n5954), .A2(n5953), .ZN(n9499) );
  INV_X1 U7614 ( .A(n9499), .ZN(n8970) );
  NAND2_X1 U7615 ( .A1(n9704), .A2(n8970), .ZN(n5955) );
  NAND2_X1 U7616 ( .A1(n5956), .A2(n9014), .ZN(n5958) );
  INV_X1 U7617 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7983) );
  OR2_X1 U7618 ( .A1(n5673), .A2(n7983), .ZN(n5957) );
  INV_X1 U7619 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5959) );
  NAND2_X1 U7620 ( .A1(n5960), .A2(n5959), .ZN(n5961) );
  NAND2_X1 U7621 ( .A1(n5973), .A2(n5961), .ZN(n9462) );
  OR2_X1 U7622 ( .A1(n9462), .A2(n6050), .ZN(n5970) );
  INV_X1 U7623 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n5967) );
  INV_X1 U7624 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n5962) );
  OR2_X1 U7625 ( .A1(n5963), .A2(n5962), .ZN(n5966) );
  INV_X1 U7626 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n5964) );
  OR2_X1 U7627 ( .A1(n5683), .A2(n5964), .ZN(n5965) );
  OAI211_X1 U7628 ( .C1(n5913), .C2(n5967), .A(n5966), .B(n5965), .ZN(n5968)
         );
  INV_X1 U7629 ( .A(n5968), .ZN(n5969) );
  NAND2_X1 U7630 ( .A1(n7995), .A2(n9014), .ZN(n5972) );
  INV_X1 U7631 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7996) );
  OR2_X1 U7632 ( .A1(n5673), .A2(n7996), .ZN(n5971) );
  NAND2_X1 U7633 ( .A1(n5973), .A2(n8919), .ZN(n5974) );
  NAND2_X1 U7634 ( .A1(n5975), .A2(n5974), .ZN(n9454) );
  INV_X1 U7635 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9453) );
  INV_X1 U7636 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9697) );
  OR2_X1 U7637 ( .A1(n5963), .A2(n9697), .ZN(n5977) );
  INV_X1 U7638 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9623) );
  OR2_X1 U7639 ( .A1(n5683), .A2(n9623), .ZN(n5976) );
  OAI211_X1 U7640 ( .C1(n5913), .C2(n9453), .A(n5977), .B(n5976), .ZN(n5978)
         );
  INV_X1 U7641 ( .A(n5978), .ZN(n5979) );
  INV_X1 U7642 ( .A(n9471), .ZN(n8992) );
  NAND2_X1 U7643 ( .A1(n9699), .A2(n8992), .ZN(n5981) );
  INV_X1 U7644 ( .A(n9616), .ZN(n9431) );
  NAND2_X1 U7645 ( .A1(n9427), .A2(n4908), .ZN(n5982) );
  OAI21_X1 U7646 ( .B1(n9445), .B2(n9616), .A(n5982), .ZN(n9412) );
  NAND2_X1 U7647 ( .A1(n8070), .A2(n9014), .ZN(n5984) );
  INV_X1 U7648 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8107) );
  OR2_X1 U7649 ( .A1(n5673), .A2(n8107), .ZN(n5983) );
  INV_X1 U7650 ( .A(n5987), .ZN(n5985) );
  NAND2_X1 U7651 ( .A1(n5985), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n8133) );
  INV_X1 U7652 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5986) );
  NAND2_X1 U7653 ( .A1(n5987), .A2(n5986), .ZN(n5988) );
  NAND2_X1 U7654 ( .A1(n8133), .A2(n5988), .ZN(n6641) );
  INV_X1 U7655 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n5991) );
  INV_X1 U7656 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9693) );
  OR2_X1 U7657 ( .A1(n5963), .A2(n9693), .ZN(n5990) );
  INV_X1 U7658 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9613) );
  OR2_X1 U7659 ( .A1(n5683), .A2(n9613), .ZN(n5989) );
  OAI211_X1 U7660 ( .C1(n5913), .C2(n5991), .A(n5990), .B(n5989), .ZN(n5992)
         );
  INV_X1 U7661 ( .A(n5992), .ZN(n5993) );
  NAND2_X1 U7662 ( .A1(n9420), .A2(n6629), .ZN(n9138) );
  NOR2_X1 U7663 ( .A1(n9420), .A2(n9435), .ZN(n5995) );
  NAND2_X1 U7664 ( .A1(n8104), .A2(n9014), .ZN(n5997) );
  INV_X1 U7665 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8142) );
  OR2_X1 U7666 ( .A1(n5673), .A2(n8142), .ZN(n5996) );
  XNOR2_X1 U7667 ( .A(n8133), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n9401) );
  NAND2_X1 U7668 ( .A1(n9401), .A2(n5685), .ZN(n6005) );
  INV_X1 U7669 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n6002) );
  INV_X1 U7670 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n5998) );
  OR2_X1 U7671 ( .A1(n5683), .A2(n5998), .ZN(n6001) );
  INV_X1 U7672 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n5999) );
  OR2_X1 U7673 ( .A1(n5963), .A2(n5999), .ZN(n6000) );
  OAI211_X1 U7674 ( .C1(n5913), .C2(n6002), .A(n6001), .B(n6000), .ZN(n6003)
         );
  INV_X1 U7675 ( .A(n6003), .ZN(n6004) );
  NAND2_X1 U7676 ( .A1(n9402), .A2(n6110), .ZN(n9140) );
  NAND2_X1 U7677 ( .A1(n9142), .A2(n9140), .ZN(n6044) );
  NAND2_X1 U7678 ( .A1(n6006), .A2(n6044), .ZN(n6112) );
  OAI21_X1 U7679 ( .B1(n6006), .B2(n6044), .A(n6112), .ZN(n9410) );
  INV_X1 U7680 ( .A(n6007), .ZN(n6011) );
  NAND2_X1 U7681 ( .A1(n6012), .A2(n6019), .ZN(n6015) );
  INV_X1 U7682 ( .A(n6015), .ZN(n6013) );
  NAND2_X1 U7683 ( .A1(n6013), .A2(n6016), .ZN(n6014) );
  XNOR2_X1 U7684 ( .A(n6065), .B(P1_IR_REG_22__SCAN_IN), .ZN(n6021) );
  NAND2_X1 U7685 ( .A1(n6021), .A2(n6395), .ZN(n6608) );
  NAND2_X1 U7686 ( .A1(n6018), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6020) );
  NAND2_X2 U7687 ( .A1(n9381), .A2(n9204), .ZN(n9261) );
  OR2_X1 U7688 ( .A1(n6608), .A2(n9261), .ZN(n6714) );
  NAND2_X1 U7689 ( .A1(n6021), .A2(n9381), .ZN(n6399) );
  NAND2_X1 U7690 ( .A1(n6399), .A2(n9261), .ZN(n6022) );
  NAND3_X1 U7691 ( .A1(n6714), .A2(n6717), .A3(n6022), .ZN(n7910) );
  NAND2_X1 U7692 ( .A1(n9155), .A2(n9204), .ZN(n9979) );
  AND2_X1 U7693 ( .A1(n6405), .A2(n6843), .ZN(n6712) );
  INV_X1 U7694 ( .A(n6417), .ZN(n7076) );
  NAND2_X1 U7695 ( .A1(n7076), .A2(n6835), .ZN(n6023) );
  NAND2_X1 U7696 ( .A1(n9284), .A2(n9965), .ZN(n9209) );
  NAND2_X1 U7697 ( .A1(n6850), .A2(n7089), .ZN(n6024) );
  NAND2_X1 U7698 ( .A1(n6025), .A2(n6024), .ZN(n7053) );
  INV_X1 U7699 ( .A(n7053), .ZN(n6027) );
  NAND2_X1 U7700 ( .A1(n6027), .A2(n6026), .ZN(n6028) );
  INV_X1 U7701 ( .A(n6029), .ZN(n9078) );
  OR2_X1 U7702 ( .A1(n9940), .A2(n7836), .ZN(n9065) );
  NAND2_X1 U7703 ( .A1(n9078), .A2(n9065), .ZN(n9054) );
  NAND2_X1 U7704 ( .A1(n9940), .A2(n7836), .ZN(n9067) );
  INV_X1 U7705 ( .A(n6030), .ZN(n9071) );
  AND2_X1 U7706 ( .A1(n9071), .A2(n9062), .ZN(n6031) );
  NAND2_X1 U7707 ( .A1(n9064), .A2(n9049), .ZN(n6032) );
  OR2_X1 U7708 ( .A1(n9054), .A2(n6032), .ZN(n9029) );
  NAND3_X1 U7709 ( .A1(n6033), .A2(n9029), .A3(n9071), .ZN(n9222) );
  NAND2_X1 U7710 ( .A1(n7384), .A2(n9076), .ZN(n7558) );
  INV_X1 U7711 ( .A(n7560), .ZN(n9032) );
  INV_X1 U7712 ( .A(n9034), .ZN(n7764) );
  INV_X1 U7713 ( .A(n9085), .ZN(n7765) );
  NOR2_X1 U7714 ( .A1(n7764), .A2(n7765), .ZN(n6035) );
  NAND2_X1 U7715 ( .A1(n9679), .A2(n9002), .ZN(n9093) );
  NAND2_X1 U7716 ( .A1(n9229), .A2(n9093), .ZN(n9088) );
  OR2_X1 U7717 ( .A1(n9672), .A2(n8930), .ZN(n9233) );
  NAND2_X1 U7718 ( .A1(n9672), .A2(n8930), .ZN(n9097) );
  NAND2_X1 U7719 ( .A1(n8012), .A2(n9097), .ZN(n9583) );
  INV_X1 U7720 ( .A(n9581), .ZN(n9584) );
  NAND2_X1 U7721 ( .A1(n9662), .A2(n6037), .ZN(n9239) );
  NAND2_X1 U7722 ( .A1(n9236), .A2(n9239), .ZN(n9564) );
  OR2_X1 U7723 ( .A1(n9657), .A2(n9102), .ZN(n9241) );
  NAND2_X1 U7724 ( .A1(n9657), .A2(n9102), .ZN(n9240) );
  NAND2_X1 U7725 ( .A1(n9556), .A2(n9240), .ZN(n9543) );
  OR2_X1 U7726 ( .A1(n9652), .A2(n9112), .ZN(n9242) );
  NAND2_X1 U7727 ( .A1(n9652), .A2(n9112), .ZN(n9248) );
  NAND2_X1 U7728 ( .A1(n9543), .A2(n9544), .ZN(n6039) );
  NAND2_X1 U7729 ( .A1(n9647), .A2(n8903), .ZN(n9109) );
  NAND2_X1 U7730 ( .A1(n9116), .A2(n9109), .ZN(n9530) );
  OR2_X1 U7731 ( .A1(n9513), .A2(n8958), .ZN(n9118) );
  NAND2_X1 U7732 ( .A1(n9513), .A2(n8958), .ZN(n9117) );
  NAND2_X1 U7733 ( .A1(n9504), .A2(n9117), .ZN(n9497) );
  INV_X1 U7734 ( .A(n9507), .ZN(n6550) );
  OR2_X1 U7735 ( .A1(n9636), .A2(n6550), .ZN(n9123) );
  NAND2_X1 U7736 ( .A1(n9636), .A2(n6550), .ZN(n9124) );
  NAND2_X1 U7737 ( .A1(n9497), .A2(n9498), .ZN(n9496) );
  NAND2_X1 U7738 ( .A1(n9496), .A2(n9124), .ZN(n9476) );
  OR2_X1 U7739 ( .A1(n9483), .A2(n8970), .ZN(n9126) );
  NAND2_X1 U7740 ( .A1(n9483), .A2(n8970), .ZN(n9467) );
  INV_X1 U7741 ( .A(n9477), .ZN(n6041) );
  NAND2_X1 U7742 ( .A1(n9626), .A2(n6041), .ZN(n9181) );
  NAND2_X1 U7743 ( .A1(n9172), .A2(n9181), .ZN(n9125) );
  NOR2_X1 U7744 ( .A1(n9125), .A2(n4510), .ZN(n6042) );
  OR2_X1 U7745 ( .A1(n9452), .A2(n8992), .ZN(n9175) );
  NAND2_X1 U7746 ( .A1(n9452), .A2(n8992), .ZN(n9186) );
  NAND2_X1 U7747 ( .A1(n9175), .A2(n9186), .ZN(n9440) );
  NAND2_X1 U7748 ( .A1(n9443), .A2(n9186), .ZN(n9433) );
  OR2_X1 U7749 ( .A1(n9616), .A2(n6643), .ZN(n9179) );
  NAND2_X1 U7750 ( .A1(n9616), .A2(n6643), .ZN(n9178) );
  NAND2_X1 U7751 ( .A1(n9433), .A2(n9434), .ZN(n9432) );
  NAND2_X1 U7752 ( .A1(n9432), .A2(n9178), .ZN(n9414) );
  INV_X1 U7753 ( .A(n9411), .ZN(n9413) );
  NAND2_X1 U7754 ( .A1(n9414), .A2(n9413), .ZN(n6045) );
  NAND2_X1 U7755 ( .A1(n9140), .A2(n9138), .ZN(n9189) );
  INV_X1 U7756 ( .A(n6044), .ZN(n9045) );
  AOI21_X1 U7757 ( .B1(n6045), .B2(n9138), .A(n9045), .ZN(n6047) );
  NAND2_X1 U7758 ( .A1(n6021), .A2(n6096), .ZN(n6046) );
  OR2_X1 U7759 ( .A1(n6397), .A2(n9204), .ZN(n9262) );
  INV_X1 U7760 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6049) );
  OR3_X1 U7761 ( .A1(n8133), .A2(n6050), .A3(n6049), .ZN(n6055) );
  INV_X1 U7762 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6136) );
  NAND2_X1 U7763 ( .A1(n5684), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6052) );
  INV_X1 U7764 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6132) );
  OR2_X1 U7765 ( .A1(n5683), .A2(n6132), .ZN(n6051) );
  OAI211_X1 U7766 ( .C1(n6136), .C2(n5963), .A(n6052), .B(n6051), .ZN(n6053)
         );
  INV_X1 U7767 ( .A(n6053), .ZN(n6054) );
  NAND2_X1 U7768 ( .A1(n6055), .A2(n6054), .ZN(n9276) );
  NAND2_X1 U7769 ( .A1(n9276), .A2(n7513), .ZN(n6056) );
  INV_X1 U7770 ( .A(n9636), .ZN(n9495) );
  NAND2_X1 U7771 ( .A1(n6060), .A2(n6813), .ZN(n7083) );
  NAND2_X1 U7772 ( .A1(n6896), .A2(n7099), .ZN(n6897) );
  OR2_X2 U7773 ( .A1(n6897), .A2(n7113), .ZN(n7479) );
  INV_X1 U7774 ( .A(n7512), .ZN(n9989) );
  NAND2_X1 U7775 ( .A1(n9917), .A2(n10005), .ZN(n7919) );
  OR2_X2 U7776 ( .A1(n7919), .A2(n9679), .ZN(n8010) );
  NAND2_X1 U7777 ( .A1(n9699), .A2(n9461), .ZN(n9449) );
  INV_X1 U7778 ( .A(n6062), .ZN(n9419) );
  INV_X1 U7779 ( .A(n9204), .ZN(n6063) );
  OAI211_X1 U7780 ( .C1(n6109), .C2(n9419), .A(n6129), .B(n9942), .ZN(n9406)
         );
  OAI211_X1 U7781 ( .C1(n9410), .C2(n9675), .A(n9400), .B(n9406), .ZN(n6105)
         );
  INV_X1 U7782 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U7783 ( .A1(n6065), .A2(n6064), .ZN(n6066) );
  NAND2_X1 U7784 ( .A1(n6066), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U7785 ( .A1(n6078), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6071) );
  NAND2_X1 U7786 ( .A1(n7997), .A2(P1_B_REG_SCAN_IN), .ZN(n6081) );
  NAND2_X1 U7787 ( .A1(n6069), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6077) );
  MUX2_X1 U7788 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6077), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n6079) );
  NAND2_X1 U7789 ( .A1(n6079), .A2(n6078), .ZN(n7984) );
  INV_X1 U7790 ( .A(n7984), .ZN(n6080) );
  MUX2_X1 U7791 ( .A(n6081), .B(P1_B_REG_SCAN_IN), .S(n6080), .Z(n6083) );
  NAND2_X1 U7792 ( .A1(n6072), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6082) );
  NOR4_X1 U7793 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6092) );
  NOR4_X1 U7794 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6091) );
  OR4_X1 U7795 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6089) );
  NOR4_X1 U7796 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6087) );
  NOR4_X1 U7797 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6086) );
  NOR4_X1 U7798 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6085) );
  NOR4_X1 U7799 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6084) );
  NAND4_X1 U7800 ( .A1(n6087), .A2(n6086), .A3(n6085), .A4(n6084), .ZN(n6088)
         );
  NOR4_X1 U7801 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n6089), .A4(n6088), .ZN(n6090) );
  AND3_X1 U7802 ( .A1(n6092), .A2(n6091), .A3(n6090), .ZN(n6093) );
  NOR2_X1 U7803 ( .A1(n9718), .A2(n6093), .ZN(n6610) );
  NOR2_X1 U7804 ( .A1(n6811), .A2(n6610), .ZN(n6095) );
  NOR2_X1 U7805 ( .A1(n7997), .A2(n7984), .ZN(n6094) );
  AOI21_X1 U7806 ( .B1(n9198), .B2(n9261), .A(n6607), .ZN(n6623) );
  AND2_X1 U7807 ( .A1(n6095), .A2(n6623), .ZN(n6711) );
  NAND2_X1 U7808 ( .A1(n6096), .A2(n9204), .ZN(n9260) );
  INV_X1 U7809 ( .A(n6097), .ZN(n8061) );
  NAND2_X1 U7810 ( .A1(n8061), .A2(n7997), .ZN(n9720) );
  OAI21_X1 U7811 ( .B1(n9718), .B2(P1_D_REG_1__SCAN_IN), .A(n9720), .ZN(n6707)
         );
  AND2_X1 U7812 ( .A1(n6621), .A2(n6707), .ZN(n6098) );
  AND2_X1 U7813 ( .A1(n6711), .A2(n6098), .ZN(n6104) );
  NAND2_X1 U7814 ( .A1(n8061), .A2(n7984), .ZN(n9721) );
  INV_X1 U7815 ( .A(n6708), .ZN(n6611) );
  MUX2_X1 U7816 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n6105), .S(n10021), .Z(n6099) );
  INV_X1 U7817 ( .A(n6099), .ZN(n6103) );
  INV_X1 U7818 ( .A(n9261), .ZN(n6100) );
  NAND2_X1 U7819 ( .A1(n10021), .A2(n9680), .ZN(n9645) );
  NAND2_X1 U7820 ( .A1(n9402), .A2(n6101), .ZN(n6102) );
  NAND2_X1 U7821 ( .A1(n6103), .A2(n6102), .ZN(P1_U3550) );
  MUX2_X1 U7822 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n6105), .S(n10010), .Z(n6106) );
  INV_X1 U7823 ( .A(n6106), .ZN(n6108) );
  NAND2_X1 U7824 ( .A1(n10010), .A2(n9680), .ZN(n9709) );
  NAND2_X1 U7825 ( .A1(n6108), .A2(n6107), .ZN(P1_U3518) );
  NAND2_X1 U7826 ( .A1(n9402), .A2(n9416), .ZN(n6111) );
  NAND2_X1 U7827 ( .A1(n6112), .A2(n6111), .ZN(n6116) );
  NAND2_X1 U7828 ( .A1(n8879), .A2(n9014), .ZN(n6114) );
  OR2_X1 U7829 ( .A1(n5673), .A2(n9730), .ZN(n6113) );
  INV_X1 U7830 ( .A(n9276), .ZN(n6115) );
  NAND2_X1 U7831 ( .A1(n8135), .A2(n6115), .ZN(n9144) );
  XNOR2_X1 U7832 ( .A(n6116), .B(n9157), .ZN(n8139) );
  INV_X1 U7833 ( .A(n9142), .ZN(n9167) );
  XNOR2_X1 U7834 ( .A(n6118), .B(n9145), .ZN(n6128) );
  INV_X1 U7835 ( .A(P1_B_REG_SCAN_IN), .ZN(n6119) );
  OR2_X1 U7836 ( .A1(n8108), .A2(n6119), .ZN(n6120) );
  AND2_X1 U7837 ( .A1(n7513), .A2(n6120), .ZN(n9388) );
  INV_X1 U7838 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n6124) );
  NAND2_X1 U7839 ( .A1(n5684), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6123) );
  INV_X1 U7840 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n6121) );
  OR2_X1 U7841 ( .A1(n5683), .A2(n6121), .ZN(n6122) );
  OAI211_X1 U7842 ( .C1(n5963), .C2(n6124), .A(n6123), .B(n6122), .ZN(n9275)
         );
  NAND2_X1 U7843 ( .A1(n9388), .A2(n9275), .ZN(n6125) );
  AOI21_X1 U7844 ( .B1(n8135), .B2(n6129), .A(n9590), .ZN(n6130) );
  NAND2_X1 U7845 ( .A1(n6130), .A2(n9392), .ZN(n8137) );
  NAND2_X1 U7846 ( .A1(n8141), .A2(n8137), .ZN(n6131) );
  AOI21_X1 U7847 ( .B1(n8139), .B2(n10007), .A(n6131), .ZN(n6135) );
  MUX2_X1 U7848 ( .A(n6132), .B(n6135), .S(n10021), .Z(n6134) );
  NAND2_X1 U7849 ( .A1(n8135), .A2(n6101), .ZN(n6133) );
  NAND2_X1 U7850 ( .A1(n6134), .A2(n6133), .ZN(P1_U3551) );
  MUX2_X1 U7851 ( .A(n6136), .B(n6135), .S(n10010), .Z(n6139) );
  NAND2_X1 U7852 ( .A1(n8135), .A2(n6137), .ZN(n6138) );
  NAND2_X1 U7853 ( .A1(n6139), .A2(n6138), .ZN(P1_U3519) );
  INV_X1 U7854 ( .A(n6140), .ZN(n6148) );
  NAND2_X1 U7855 ( .A1(n6903), .A2(n6659), .ZN(n6864) );
  OR2_X1 U7856 ( .A1(n6142), .A2(n7687), .ZN(n6143) );
  NAND2_X1 U7857 ( .A1(n6143), .A2(n6322), .ZN(n6145) );
  INV_X1 U7858 ( .A(n6145), .ZN(n6146) );
  OAI21_X1 U7859 ( .B1(n7372), .B2(n6880), .A(n7373), .ZN(n6147) );
  OR2_X1 U7860 ( .A1(n6149), .A2(n8755), .ZN(n6152) );
  NAND2_X1 U7861 ( .A1(n8755), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6151) );
  NAND2_X1 U7862 ( .A1(n6152), .A2(n4901), .ZN(P2_U3488) );
  INV_X1 U7863 ( .A(SI_29_), .ZN(n7305) );
  INV_X1 U7864 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8203) );
  INV_X1 U7865 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9011) );
  MUX2_X1 U7866 ( .A(n8203), .B(n9011), .S(n4350), .Z(n6157) );
  NAND2_X1 U7867 ( .A1(n6157), .A2(n7330), .ZN(n6169) );
  INV_X1 U7868 ( .A(n6157), .ZN(n6158) );
  NAND2_X1 U7869 ( .A1(n6158), .A2(SI_30_), .ZN(n6159) );
  NAND2_X1 U7870 ( .A1(n6169), .A2(n6159), .ZN(n6170) );
  NOR2_X1 U7871 ( .A1(n5096), .A2(n8203), .ZN(n6160) );
  INV_X1 U7872 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n6165) );
  NAND2_X1 U7873 ( .A1(n6161), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6164) );
  NAND2_X1 U7874 ( .A1(n6162), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6163) );
  OAI211_X1 U7875 ( .C1(n6165), .C2(n5514), .A(n6164), .B(n6163), .ZN(n6166)
         );
  INV_X1 U7876 ( .A(n6166), .ZN(n6167) );
  MUX2_X1 U7877 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n4350), .Z(n6172) );
  INV_X1 U7878 ( .A(SI_31_), .ZN(n7338) );
  XNOR2_X1 U7879 ( .A(n6172), .B(n7338), .ZN(n6173) );
  NAND2_X1 U7880 ( .A1(n9015), .A2(n6175), .ZN(n6178) );
  INV_X1 U7881 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6176) );
  OR2_X1 U7882 ( .A1(n5096), .A2(n6176), .ZN(n6177) );
  AOI21_X1 U7883 ( .B1(n8746), .B2(n8549), .A(n8741), .ZN(n6182) );
  INV_X1 U7884 ( .A(n8746), .ZN(n6179) );
  NAND2_X1 U7885 ( .A1(n6179), .A2(n6184), .ZN(n6372) );
  AND2_X1 U7886 ( .A1(n6372), .A2(n6180), .ZN(n6329) );
  INV_X1 U7887 ( .A(n6329), .ZN(n6181) );
  INV_X1 U7888 ( .A(n6184), .ZN(n8356) );
  AND2_X1 U7889 ( .A1(n8746), .A2(n8356), .ZN(n6370) );
  INV_X1 U7890 ( .A(n6189), .ZN(n6186) );
  NOR3_X1 U7891 ( .A1(n6374), .A2(n8539), .A3(n6187), .ZN(n6185) );
  NOR2_X1 U7892 ( .A1(n5543), .A2(n6187), .ZN(n6188) );
  NAND2_X1 U7893 ( .A1(n6191), .A2(n6190), .ZN(n6389) );
  AOI21_X1 U7894 ( .B1(n6339), .B2(n6299), .A(n6337), .ZN(n6304) );
  INV_X1 U7895 ( .A(n6192), .ZN(n6196) );
  OAI21_X1 U7896 ( .B1(n6194), .B2(n7846), .A(n6193), .ZN(n6195) );
  MUX2_X1 U7897 ( .A(n6196), .B(n6195), .S(n6322), .Z(n6198) );
  NAND2_X1 U7898 ( .A1(n6198), .A2(n5527), .ZN(n6205) );
  NAND2_X1 U7899 ( .A1(n6213), .A2(n6199), .ZN(n6202) );
  NAND2_X1 U7900 ( .A1(n6207), .A2(n6200), .ZN(n6201) );
  MUX2_X1 U7901 ( .A(n6202), .B(n6201), .S(n6659), .Z(n6203) );
  INV_X1 U7902 ( .A(n6203), .ZN(n6204) );
  NAND2_X1 U7903 ( .A1(n6205), .A2(n6204), .ZN(n6206) );
  NAND2_X1 U7904 ( .A1(n6206), .A2(n7691), .ZN(n6217) );
  OAI211_X1 U7905 ( .C1(n6217), .C2(n4598), .A(n6208), .B(n7545), .ZN(n6212)
         );
  AND2_X1 U7906 ( .A1(n6215), .A2(n6218), .ZN(n6211) );
  INV_X1 U7907 ( .A(n6209), .ZN(n6210) );
  AOI21_X1 U7908 ( .B1(n6212), .B2(n6211), .A(n6210), .ZN(n6223) );
  INV_X1 U7909 ( .A(n6213), .ZN(n6216) );
  OAI211_X1 U7910 ( .C1(n6217), .C2(n6216), .A(n6215), .B(n6214), .ZN(n6221)
         );
  INV_X1 U7911 ( .A(n6218), .ZN(n6219) );
  AOI21_X1 U7912 ( .B1(n6221), .B2(n6220), .A(n6219), .ZN(n6222) );
  MUX2_X1 U7913 ( .A(n6223), .B(n6222), .S(n6659), .Z(n6227) );
  NAND2_X1 U7914 ( .A1(n6233), .A2(n6234), .ZN(n6225) );
  NAND2_X1 U7915 ( .A1(n6230), .A2(n6229), .ZN(n6224) );
  MUX2_X1 U7916 ( .A(n6225), .B(n6224), .S(n6659), .Z(n6236) );
  INV_X1 U7917 ( .A(n6236), .ZN(n6226) );
  NAND3_X1 U7918 ( .A1(n6227), .A2(n6226), .A3(n6350), .ZN(n6241) );
  AND2_X1 U7919 ( .A1(n6229), .A2(n6228), .ZN(n6231) );
  OAI211_X1 U7920 ( .C1(n6236), .C2(n6231), .A(n5533), .B(n6230), .ZN(n6238)
         );
  NAND2_X1 U7921 ( .A1(n7960), .A2(n7927), .ZN(n6232) );
  AND2_X1 U7922 ( .A1(n6233), .A2(n6232), .ZN(n6235) );
  OAI211_X1 U7923 ( .C1(n6236), .C2(n6235), .A(n6234), .B(n7931), .ZN(n6237)
         );
  MUX2_X1 U7924 ( .A(n6238), .B(n6237), .S(n6659), .Z(n6239) );
  INV_X1 U7925 ( .A(n6239), .ZN(n6240) );
  NAND2_X1 U7926 ( .A1(n6241), .A2(n6240), .ZN(n6246) );
  INV_X1 U7927 ( .A(n6354), .ZN(n6242) );
  AOI21_X1 U7928 ( .B1(n6246), .B2(n6243), .A(n6242), .ZN(n6248) );
  AND2_X1 U7929 ( .A1(n5533), .A2(n6354), .ZN(n6245) );
  INV_X1 U7930 ( .A(n6353), .ZN(n6244) );
  AOI21_X1 U7931 ( .B1(n6246), .B2(n6245), .A(n6244), .ZN(n6247) );
  MUX2_X1 U7932 ( .A(n6248), .B(n6247), .S(n6659), .Z(n6249) );
  NAND2_X1 U7933 ( .A1(n6249), .A2(n7973), .ZN(n6253) );
  MUX2_X1 U7934 ( .A(n6251), .B(n6250), .S(n6322), .Z(n6252) );
  MUX2_X1 U7935 ( .A(n8360), .B(n8077), .S(n6659), .Z(n6255) );
  AOI22_X1 U7936 ( .A1(n6253), .A2(n6252), .B1(n6344), .B2(n6255), .ZN(n6257)
         );
  INV_X1 U7937 ( .A(n6345), .ZN(n6254) );
  NOR2_X1 U7938 ( .A1(n6255), .A2(n6254), .ZN(n6256) );
  OAI21_X1 U7939 ( .B1(n6257), .B2(n6256), .A(n8113), .ZN(n6261) );
  XNOR2_X1 U7940 ( .A(n8792), .B(n8709), .ZN(n8723) );
  MUX2_X1 U7941 ( .A(n6259), .B(n6258), .S(n6659), .Z(n6260) );
  NAND3_X1 U7942 ( .A1(n6261), .A2(n8723), .A3(n6260), .ZN(n6265) );
  INV_X1 U7943 ( .A(n8705), .ZN(n8707) );
  MUX2_X1 U7944 ( .A(n6263), .B(n6262), .S(n6659), .Z(n6264) );
  NAND3_X1 U7945 ( .A1(n6265), .A2(n8707), .A3(n6264), .ZN(n6271) );
  MUX2_X1 U7946 ( .A(n6267), .B(n6266), .S(n6659), .Z(n6268) );
  INV_X1 U7947 ( .A(n6268), .ZN(n6269) );
  NOR2_X1 U7948 ( .A1(n6340), .A2(n6269), .ZN(n6270) );
  NAND2_X1 U7949 ( .A1(n6271), .A2(n6270), .ZN(n6276) );
  NAND3_X1 U7950 ( .A1(n6276), .A2(n6341), .A3(n6272), .ZN(n6273) );
  INV_X1 U7951 ( .A(n6343), .ZN(n6275) );
  NAND3_X1 U7952 ( .A1(n6273), .A2(n6275), .A3(n6280), .ZN(n6279) );
  NAND3_X1 U7953 ( .A1(n6276), .A2(n6275), .A3(n6274), .ZN(n6277) );
  NAND2_X1 U7954 ( .A1(n6277), .A2(n6341), .ZN(n6278) );
  OAI211_X1 U7955 ( .C1(n6288), .C2(n4613), .A(n6289), .B(n6280), .ZN(n6283)
         );
  INV_X1 U7956 ( .A(n6290), .ZN(n6281) );
  AOI21_X1 U7957 ( .B1(n6283), .B2(n6282), .A(n6281), .ZN(n6302) );
  NAND3_X1 U7958 ( .A1(n6299), .A2(n6322), .A3(n6284), .ZN(n6301) );
  OAI21_X1 U7959 ( .B1(n6659), .B2(n6292), .A(n4610), .ZN(n6298) );
  INV_X1 U7960 ( .A(n6284), .ZN(n6285) );
  OAI21_X1 U7961 ( .B1(n6299), .B2(n6322), .A(n6286), .ZN(n6297) );
  NAND3_X1 U7962 ( .A1(n6288), .A2(n6287), .A3(n8647), .ZN(n6291) );
  NAND3_X1 U7963 ( .A1(n6291), .A2(n6290), .A3(n6289), .ZN(n6295) );
  INV_X1 U7964 ( .A(n6292), .ZN(n6293) );
  AOI211_X1 U7965 ( .C1(n6295), .C2(n6294), .A(n6293), .B(n6322), .ZN(n6296)
         );
  OAI21_X1 U7966 ( .B1(n6302), .B2(n6301), .A(n6300), .ZN(n6303) );
  OAI211_X1 U7967 ( .C1(n6304), .C2(n6322), .A(n6303), .B(n8600), .ZN(n6314)
         );
  INV_X1 U7968 ( .A(n6305), .ZN(n6307) );
  MUX2_X1 U7969 ( .A(n6307), .B(n6306), .S(n6659), .Z(n6309) );
  INV_X1 U7970 ( .A(n6308), .ZN(n6311) );
  NOR2_X1 U7971 ( .A1(n6309), .A2(n8591), .ZN(n6313) );
  MUX2_X1 U7972 ( .A(n6311), .B(n6310), .S(n6659), .Z(n6312) );
  NOR2_X1 U7973 ( .A1(n8589), .A2(n6659), .ZN(n6316) );
  NOR2_X1 U7974 ( .A1(n8358), .A2(n6322), .ZN(n6315) );
  MUX2_X1 U7975 ( .A(n6316), .B(n6315), .S(n8210), .Z(n6317) );
  MUX2_X1 U7976 ( .A(n8357), .B(n8197), .S(n6322), .Z(n6318) );
  NAND2_X1 U7977 ( .A1(n6320), .A2(n6318), .ZN(n6328) );
  INV_X1 U7978 ( .A(n6369), .ZN(n6319) );
  INV_X1 U7979 ( .A(n6321), .ZN(n6323) );
  NAND2_X1 U7980 ( .A1(n6371), .A2(n6324), .ZN(n6325) );
  OAI211_X1 U7981 ( .C1(n6330), .C2(n8357), .A(n6329), .B(n6328), .ZN(n6332)
         );
  OAI21_X1 U7982 ( .B1(n6370), .B2(n6659), .A(n6372), .ZN(n6331) );
  INV_X1 U7983 ( .A(n6374), .ZN(n6379) );
  INV_X1 U7984 ( .A(n6335), .ZN(n6336) );
  INV_X1 U7985 ( .A(n8619), .ZN(n6364) );
  INV_X1 U7986 ( .A(n8617), .ZN(n6338) );
  OR2_X1 U7987 ( .A1(n6339), .A2(n6338), .ZN(n8626) );
  INV_X1 U7988 ( .A(n8626), .ZN(n8624) );
  INV_X1 U7989 ( .A(n6341), .ZN(n6342) );
  INV_X1 U7990 ( .A(n8113), .ZN(n8111) );
  AND2_X1 U7991 ( .A1(n6346), .A2(n7042), .ZN(n7728) );
  AND4_X1 U7992 ( .A1(n7691), .A2(n7728), .A3(n5527), .A4(n6946), .ZN(n6349)
         );
  NAND2_X1 U7993 ( .A1(n6348), .A2(n6347), .ZN(n7548) );
  NAND4_X1 U7994 ( .A1(n6349), .A2(n7612), .A3(n7043), .A4(n7548), .ZN(n6352)
         );
  NOR4_X1 U7995 ( .A1(n6352), .A2(n5179), .A3(n5207), .A4(n7737), .ZN(n6356)
         );
  NAND2_X1 U7996 ( .A1(n6354), .A2(n6353), .ZN(n8032) );
  INV_X1 U7997 ( .A(n8032), .ZN(n6355) );
  NAND4_X1 U7998 ( .A1(n6356), .A2(n6355), .A3(n7973), .A4(n7888), .ZN(n6357)
         );
  OR4_X1 U7999 ( .A1(n8705), .A2(n8004), .A3(n8111), .A4(n6357), .ZN(n6358) );
  INV_X1 U8000 ( .A(n8723), .ZN(n8725) );
  NOR3_X1 U8001 ( .A1(n8687), .A2(n6358), .A3(n8725), .ZN(n6359) );
  NAND4_X1 U8002 ( .A1(n8664), .A2(n8676), .A3(n4862), .A4(n6359), .ZN(n6360)
         );
  OR2_X1 U8003 ( .A1(n8651), .A2(n6360), .ZN(n6361) );
  NOR2_X1 U8004 ( .A1(n6362), .A2(n6361), .ZN(n6363) );
  NAND4_X1 U8005 ( .A1(n8600), .A2(n6364), .A3(n8624), .A4(n6363), .ZN(n6365)
         );
  NOR2_X1 U8006 ( .A1(n8591), .A2(n6365), .ZN(n6367) );
  INV_X1 U8007 ( .A(n8580), .ZN(n6366) );
  NAND3_X1 U8008 ( .A1(n8191), .A2(n6367), .A3(n6366), .ZN(n6368) );
  NOR2_X1 U8009 ( .A1(n6369), .A2(n6368), .ZN(n6373) );
  INV_X1 U8010 ( .A(n6370), .ZN(n6371) );
  NAND4_X1 U8011 ( .A1(n4390), .A2(n6373), .A3(n6372), .A4(n6371), .ZN(n6376)
         );
  OR4_X1 U8012 ( .A1(n6376), .A2(n8539), .A3(n6374), .A4(n6904), .ZN(n6378) );
  INV_X1 U8013 ( .A(n6904), .ZN(n6375) );
  NAND3_X1 U8014 ( .A1(n6376), .A2(n6375), .A3(n8539), .ZN(n6377) );
  OAI211_X1 U8015 ( .C1(n6379), .C2(n5543), .A(n6378), .B(n6377), .ZN(n6380)
         );
  NOR2_X1 U8016 ( .A1(n6381), .A2(n6380), .ZN(n6386) );
  INV_X1 U8017 ( .A(n6382), .ZN(n6384) );
  NAND2_X1 U8018 ( .A1(n6386), .A2(n6385), .ZN(n6388) );
  OR2_X1 U8019 ( .A1(n6865), .A2(P2_U3151), .ZN(n7946) );
  INV_X1 U8020 ( .A(n7946), .ZN(n6387) );
  OAI21_X1 U8021 ( .B1(n6389), .B2(n6388), .A(n6387), .ZN(n6394) );
  NOR2_X1 U8022 ( .A1(n6390), .A2(n6875), .ZN(n6871) );
  NAND3_X1 U8023 ( .A1(n6871), .A2(n6953), .A3(n8529), .ZN(n6391) );
  OAI211_X1 U8024 ( .C1(n6392), .C2(n7946), .A(n6391), .B(P2_B_REG_SCAN_IN), 
        .ZN(n6393) );
  NAND2_X1 U8025 ( .A1(n6394), .A2(n6393), .ZN(P2_U3296) );
  NAND2_X1 U8026 ( .A1(n6395), .A2(n9204), .ZN(n6398) );
  INV_X1 U8027 ( .A(n6398), .ZN(n6396) );
  INV_X2 U8028 ( .A(n6551), .ZN(n6415) );
  NAND2_X1 U8029 ( .A1(n9280), .A2(n6603), .ZN(n6402) );
  AND2_X1 U8030 ( .A1(n6647), .A2(n6398), .ZN(n6400) );
  NAND2_X2 U8031 ( .A1(n6507), .A2(n6423), .ZN(n6420) );
  CLKBUF_X3 U8032 ( .A(n6420), .Z(n6604) );
  NAND2_X1 U8033 ( .A1(n7113), .A2(n6604), .ZN(n6401) );
  NAND2_X1 U8034 ( .A1(n6402), .A2(n6401), .ZN(n6403) );
  INV_X2 U8035 ( .A(n6423), .ZN(n6434) );
  XNOR2_X1 U8036 ( .A(n6403), .B(n6601), .ZN(n6452) );
  INV_X1 U8037 ( .A(n6452), .ZN(n6454) );
  BUF_X8 U8038 ( .A(n6415), .Z(n6603) );
  AOI22_X1 U8039 ( .A1(n9280), .A2(n6407), .B1(n6603), .B2(n7113), .ZN(n6453)
         );
  NAND2_X1 U8040 ( .A1(n6713), .A2(n6407), .ZN(n6410) );
  AND2_X1 U8041 ( .A1(n6410), .A2(n6409), .ZN(n6791) );
  OAI21_X1 U8042 ( .B1(n6792), .B2(n6791), .A(n4916), .ZN(n6831) );
  NAND2_X1 U8043 ( .A1(n6835), .A2(n6420), .ZN(n6412) );
  NAND2_X1 U8044 ( .A1(n6413), .A2(n6412), .ZN(n6414) );
  XNOR2_X1 U8045 ( .A(n6414), .B(n6434), .ZN(n6419) );
  AND2_X1 U8046 ( .A1(n6415), .A2(n6835), .ZN(n6416) );
  XNOR2_X1 U8047 ( .A(n6419), .B(n6418), .ZN(n6830) );
  NOR2_X2 U8048 ( .A1(n6831), .A2(n6830), .ZN(n6829) );
  AND2_X1 U8049 ( .A1(n6419), .A2(n6418), .ZN(n6823) );
  NAND2_X1 U8050 ( .A1(n7089), .A2(n6420), .ZN(n6422) );
  NAND2_X1 U8051 ( .A1(n9284), .A2(n6603), .ZN(n6421) );
  NAND2_X1 U8052 ( .A1(n6422), .A2(n6421), .ZN(n6424) );
  XNOR2_X1 U8053 ( .A(n6424), .B(n6434), .ZN(n6426) );
  AND2_X1 U8054 ( .A1(n7089), .A2(n6603), .ZN(n6425) );
  NAND2_X1 U8055 ( .A1(n6426), .A2(n6427), .ZN(n6431) );
  INV_X1 U8056 ( .A(n6426), .ZN(n6429) );
  INV_X1 U8057 ( .A(n6427), .ZN(n6428) );
  NAND2_X1 U8058 ( .A1(n6429), .A2(n6428), .ZN(n6430) );
  AND2_X1 U8059 ( .A1(n6431), .A2(n6430), .ZN(n6822) );
  NAND2_X1 U8060 ( .A1(n6821), .A2(n6431), .ZN(n8892) );
  NAND2_X1 U8061 ( .A1(n9283), .A2(n6603), .ZN(n6433) );
  NAND2_X1 U8062 ( .A1(n8896), .A2(n6604), .ZN(n6432) );
  NAND2_X1 U8063 ( .A1(n6433), .A2(n6432), .ZN(n6435) );
  XNOR2_X1 U8064 ( .A(n6435), .B(n6601), .ZN(n6436) );
  AOI22_X1 U8065 ( .A1(n9283), .A2(n6407), .B1(n6603), .B2(n8896), .ZN(n6437)
         );
  XNOR2_X1 U8066 ( .A(n6436), .B(n6437), .ZN(n8893) );
  NAND2_X1 U8067 ( .A1(n8892), .A2(n8893), .ZN(n8891) );
  INV_X1 U8068 ( .A(n6436), .ZN(n6438) );
  AND2_X1 U8069 ( .A1(n7069), .A2(n6603), .ZN(n6440) );
  AOI21_X1 U8070 ( .B1(n9282), .B2(n6407), .A(n6440), .ZN(n6445) );
  NAND2_X1 U8071 ( .A1(n9282), .A2(n6603), .ZN(n6442) );
  NAND2_X1 U8072 ( .A1(n7069), .A2(n6604), .ZN(n6441) );
  NAND2_X1 U8073 ( .A1(n6442), .A2(n6441), .ZN(n6443) );
  XOR2_X1 U8074 ( .A(n6445), .B(n6444), .Z(n6651) );
  INV_X1 U8075 ( .A(n6444), .ZN(n6446) );
  NOR2_X1 U8076 ( .A1(n6446), .A2(n6445), .ZN(n6451) );
  NAND2_X1 U8077 ( .A1(n9281), .A2(n6415), .ZN(n6448) );
  NAND2_X1 U8078 ( .A1(n6941), .A2(n6604), .ZN(n6447) );
  NAND2_X1 U8079 ( .A1(n6448), .A2(n6447), .ZN(n6449) );
  XNOR2_X1 U8080 ( .A(n6449), .B(n6601), .ZN(n6450) );
  AOI22_X1 U8081 ( .A1(n9281), .A2(n6407), .B1(n6603), .B2(n6941), .ZN(n6933)
         );
  OAI21_X1 U8082 ( .B1(n6649), .B2(n6451), .A(n6450), .ZN(n6931) );
  OAI21_X1 U8083 ( .B1(n6930), .B2(n6933), .A(n6931), .ZN(n7034) );
  XOR2_X1 U8084 ( .A(n6453), .B(n6452), .Z(n7035) );
  NAND2_X1 U8085 ( .A1(n7598), .A2(n6604), .ZN(n6456) );
  NAND2_X1 U8086 ( .A1(n9931), .A2(n6603), .ZN(n6455) );
  NAND2_X1 U8087 ( .A1(n6456), .A2(n6455), .ZN(n6457) );
  XNOR2_X1 U8088 ( .A(n6457), .B(n6434), .ZN(n6459) );
  AOI22_X1 U8089 ( .A1(n7598), .A2(n6603), .B1(n9931), .B2(n6407), .ZN(n6458)
         );
  NOR2_X1 U8090 ( .A1(n6459), .A2(n6458), .ZN(n7132) );
  AOI22_X1 U8091 ( .A1(n7512), .A2(n6604), .B1(n6603), .B2(n9930), .ZN(n6460)
         );
  XOR2_X1 U8092 ( .A(n6601), .B(n6460), .Z(n7832) );
  NAND2_X1 U8093 ( .A1(n7512), .A2(n6603), .ZN(n6462) );
  NAND2_X1 U8094 ( .A1(n9930), .A2(n6407), .ZN(n6461) );
  NAND2_X1 U8095 ( .A1(n6462), .A2(n6461), .ZN(n6468) );
  NAND2_X1 U8096 ( .A1(n9940), .A2(n6603), .ZN(n6464) );
  NAND2_X1 U8097 ( .A1(n9922), .A2(n6407), .ZN(n6463) );
  NAND2_X1 U8098 ( .A1(n6464), .A2(n6463), .ZN(n7677) );
  NAND2_X1 U8099 ( .A1(n9922), .A2(n6603), .ZN(n6465) );
  NAND2_X1 U8100 ( .A1(n6466), .A2(n6465), .ZN(n6467) );
  XNOR2_X1 U8101 ( .A(n6467), .B(n6601), .ZN(n6471) );
  AOI22_X1 U8102 ( .A1(n7832), .A2(n6468), .B1(n7677), .B2(n6471), .ZN(n6474)
         );
  INV_X1 U8103 ( .A(n7677), .ZN(n6469) );
  INV_X1 U8104 ( .A(n6468), .ZN(n7831) );
  NAND2_X1 U8105 ( .A1(n7831), .A2(n6469), .ZN(n6470) );
  OAI22_X1 U8106 ( .A1(n7832), .A2(n6472), .B1(n6471), .B2(n6470), .ZN(n6473)
         );
  AOI22_X1 U8107 ( .A1(n7882), .A2(n6604), .B1(n6603), .B2(n9910), .ZN(n6475)
         );
  XNOR2_X1 U8108 ( .A(n6475), .B(n6601), .ZN(n7875) );
  NAND2_X1 U8109 ( .A1(n7882), .A2(n6603), .ZN(n6477) );
  NAND2_X1 U8110 ( .A1(n9910), .A2(n6407), .ZN(n6476) );
  AND2_X1 U8111 ( .A1(n6477), .A2(n6476), .ZN(n7874) );
  NAND2_X1 U8112 ( .A1(n7391), .A2(n6604), .ZN(n6479) );
  NAND2_X1 U8113 ( .A1(n9279), .A2(n6603), .ZN(n6478) );
  NAND2_X1 U8114 ( .A1(n6479), .A2(n6478), .ZN(n6480) );
  XNOR2_X1 U8115 ( .A(n6480), .B(n6434), .ZN(n7796) );
  NAND2_X1 U8116 ( .A1(n7391), .A2(n6603), .ZN(n6482) );
  NAND2_X1 U8117 ( .A1(n9279), .A2(n6407), .ZN(n6481) );
  AOI22_X1 U8118 ( .A1(n7875), .A2(n7874), .B1(n7796), .B2(n7798), .ZN(n6488)
         );
  INV_X1 U8119 ( .A(n7796), .ZN(n7872) );
  INV_X1 U8120 ( .A(n7798), .ZN(n6483) );
  INV_X1 U8121 ( .A(n7874), .ZN(n6484) );
  AOI21_X1 U8122 ( .B1(n7872), .B2(n6483), .A(n6484), .ZN(n6486) );
  NAND3_X1 U8123 ( .A1(n7872), .A2(n6484), .A3(n6483), .ZN(n6485) );
  OAI21_X1 U8124 ( .B1(n7875), .B2(n6486), .A(n6485), .ZN(n6487) );
  NAND2_X1 U8125 ( .A1(n9914), .A2(n6604), .ZN(n6490) );
  NAND2_X1 U8126 ( .A1(n9278), .A2(n6603), .ZN(n6489) );
  NAND2_X1 U8127 ( .A1(n6490), .A2(n6489), .ZN(n6491) );
  XNOR2_X1 U8128 ( .A(n6491), .B(n6601), .ZN(n6495) );
  NAND2_X1 U8129 ( .A1(n9914), .A2(n6603), .ZN(n6493) );
  NAND2_X1 U8130 ( .A1(n9278), .A2(n6407), .ZN(n6492) );
  NAND2_X1 U8131 ( .A1(n6493), .A2(n6492), .ZN(n6494) );
  NOR2_X1 U8132 ( .A1(n6495), .A2(n6494), .ZN(n6496) );
  AOI21_X1 U8133 ( .B1(n6495), .B2(n6494), .A(n6496), .ZN(n7757) );
  INV_X1 U8134 ( .A(n6496), .ZN(n6497) );
  AND2_X1 U8135 ( .A1(n9909), .A2(n6407), .ZN(n6498) );
  AOI21_X1 U8136 ( .B1(n6499), .B2(n6603), .A(n6498), .ZN(n6502) );
  AOI22_X1 U8137 ( .A1(n6499), .A2(n6604), .B1(n6603), .B2(n9909), .ZN(n6500)
         );
  XNOR2_X1 U8138 ( .A(n6500), .B(n6601), .ZN(n6501) );
  XOR2_X1 U8139 ( .A(n6502), .B(n6501), .Z(n7849) );
  AOI22_X1 U8140 ( .A1(n9679), .A2(n6604), .B1(n6603), .B2(n9277), .ZN(n6503)
         );
  XNOR2_X1 U8141 ( .A(n6503), .B(n6601), .ZN(n6504) );
  NAND2_X1 U8142 ( .A1(n6505), .A2(n6504), .ZN(n6509) );
  OAI22_X1 U8143 ( .A1(n7989), .A2(n6551), .B1(n9002), .B2(n6507), .ZN(n7986)
         );
  INV_X1 U8144 ( .A(n6514), .ZN(n6512) );
  AOI22_X1 U8145 ( .A1(n9672), .A2(n6604), .B1(n6603), .B2(n9587), .ZN(n6510)
         );
  XNOR2_X1 U8146 ( .A(n6510), .B(n6601), .ZN(n6513) );
  INV_X1 U8147 ( .A(n6513), .ZN(n6511) );
  NAND2_X1 U8148 ( .A1(n6512), .A2(n6511), .ZN(n6515) );
  NAND2_X1 U8149 ( .A1(n6514), .A2(n6513), .ZN(n6516) );
  AOI22_X1 U8150 ( .A1(n9672), .A2(n6603), .B1(n6407), .B2(n9587), .ZN(n8996)
         );
  AND2_X1 U8151 ( .A1(n9575), .A2(n6407), .ZN(n6517) );
  AOI21_X1 U8152 ( .B1(n9667), .B2(n6603), .A(n6517), .ZN(n6520) );
  AOI22_X1 U8153 ( .A1(n9667), .A2(n6604), .B1(n6603), .B2(n9575), .ZN(n6518)
         );
  XNOR2_X1 U8154 ( .A(n6518), .B(n6601), .ZN(n6519) );
  XOR2_X1 U8155 ( .A(n6520), .B(n6519), .Z(n8927) );
  NAND2_X1 U8156 ( .A1(n9662), .A2(n6604), .ZN(n6523) );
  NAND2_X1 U8157 ( .A1(n9586), .A2(n6603), .ZN(n6522) );
  NAND2_X1 U8158 ( .A1(n6523), .A2(n6522), .ZN(n6524) );
  XNOR2_X1 U8159 ( .A(n6524), .B(n6601), .ZN(n6527) );
  NAND2_X1 U8160 ( .A1(n9662), .A2(n6603), .ZN(n6526) );
  NAND2_X1 U8161 ( .A1(n9586), .A2(n6407), .ZN(n6525) );
  NAND2_X1 U8162 ( .A1(n6526), .A2(n6525), .ZN(n6528) );
  NAND2_X1 U8163 ( .A1(n6527), .A2(n6528), .ZN(n8936) );
  INV_X1 U8164 ( .A(n6527), .ZN(n6530) );
  INV_X1 U8165 ( .A(n6528), .ZN(n6529) );
  NAND2_X1 U8166 ( .A1(n6530), .A2(n6529), .ZN(n8935) );
  NAND2_X1 U8167 ( .A1(n9657), .A2(n6604), .ZN(n6532) );
  NAND2_X1 U8168 ( .A1(n9574), .A2(n6603), .ZN(n6531) );
  NAND2_X1 U8169 ( .A1(n6532), .A2(n6531), .ZN(n6533) );
  XNOR2_X1 U8170 ( .A(n6533), .B(n6601), .ZN(n6535) );
  XNOR2_X1 U8171 ( .A(n6534), .B(n6535), .ZN(n8976) );
  AOI22_X1 U8172 ( .A1(n9657), .A2(n6603), .B1(n6407), .B2(n9574), .ZN(n8978)
         );
  NAND2_X1 U8173 ( .A1(n8976), .A2(n8978), .ZN(n8977) );
  INV_X1 U8174 ( .A(n6534), .ZN(n6536) );
  OR2_X1 U8175 ( .A1(n6536), .A2(n6535), .ZN(n6537) );
  NAND2_X1 U8176 ( .A1(n8977), .A2(n6537), .ZN(n8901) );
  NAND2_X1 U8177 ( .A1(n9652), .A2(n6604), .ZN(n6539) );
  NAND2_X1 U8178 ( .A1(n9559), .A2(n6415), .ZN(n6538) );
  NAND2_X1 U8179 ( .A1(n6539), .A2(n6538), .ZN(n6540) );
  XNOR2_X1 U8180 ( .A(n6540), .B(n6601), .ZN(n6543) );
  AOI22_X1 U8181 ( .A1(n9652), .A2(n6603), .B1(n6407), .B2(n9559), .ZN(n6541)
         );
  XNOR2_X1 U8182 ( .A(n6543), .B(n6541), .ZN(n8902) );
  INV_X1 U8183 ( .A(n6541), .ZN(n6542) );
  AOI22_X1 U8184 ( .A1(n9647), .A2(n6604), .B1(n6603), .B2(n9546), .ZN(n6545)
         );
  XOR2_X1 U8185 ( .A(n6601), .B(n6545), .Z(n8955) );
  OAI22_X1 U8186 ( .A1(n9529), .A2(n6551), .B1(n8903), .B2(n6507), .ZN(n8954)
         );
  AOI22_X1 U8187 ( .A1(n9513), .A2(n6604), .B1(n6603), .B2(n9533), .ZN(n6546)
         );
  XNOR2_X1 U8188 ( .A(n6546), .B(n6423), .ZN(n6547) );
  AOI22_X1 U8189 ( .A1(n9513), .A2(n6603), .B1(n6407), .B2(n9533), .ZN(n6548)
         );
  XNOR2_X1 U8190 ( .A(n6547), .B(n6548), .ZN(n8910) );
  AOI22_X1 U8191 ( .A1(n9636), .A2(n6604), .B1(n6603), .B2(n9507), .ZN(n6549)
         );
  XNOR2_X1 U8192 ( .A(n6549), .B(n6423), .ZN(n6553) );
  OAI22_X1 U8193 ( .A1(n9495), .A2(n6551), .B1(n6550), .B2(n6507), .ZN(n8967)
         );
  NAND2_X1 U8194 ( .A1(n9483), .A2(n6604), .ZN(n6557) );
  NAND2_X1 U8195 ( .A1(n9499), .A2(n6415), .ZN(n6556) );
  NAND2_X1 U8196 ( .A1(n6557), .A2(n6556), .ZN(n6558) );
  XNOR2_X1 U8197 ( .A(n6558), .B(n6434), .ZN(n6560) );
  AND2_X1 U8198 ( .A1(n9499), .A2(n6407), .ZN(n6559) );
  AOI21_X1 U8199 ( .B1(n9483), .B2(n6603), .A(n6559), .ZN(n6561) );
  NAND2_X1 U8200 ( .A1(n6560), .A2(n6561), .ZN(n8944) );
  INV_X1 U8201 ( .A(n6560), .ZN(n6563) );
  INV_X1 U8202 ( .A(n6561), .ZN(n6562) );
  NAND2_X1 U8203 ( .A1(n6563), .A2(n6562), .ZN(n6564) );
  AND2_X1 U8204 ( .A1(n8944), .A2(n6564), .ZN(n8885) );
  NAND2_X1 U8205 ( .A1(n9626), .A2(n6604), .ZN(n6566) );
  NAND2_X1 U8206 ( .A1(n9477), .A2(n6415), .ZN(n6565) );
  NAND2_X1 U8207 ( .A1(n6566), .A2(n6565), .ZN(n6567) );
  XNOR2_X1 U8208 ( .A(n6567), .B(n6434), .ZN(n6569) );
  AND2_X1 U8209 ( .A1(n9477), .A2(n6407), .ZN(n6568) );
  AOI21_X1 U8210 ( .B1(n9626), .B2(n6603), .A(n6568), .ZN(n6570) );
  NAND2_X1 U8211 ( .A1(n6569), .A2(n6570), .ZN(n6574) );
  INV_X1 U8212 ( .A(n6569), .ZN(n6572) );
  INV_X1 U8213 ( .A(n6570), .ZN(n6571) );
  NAND2_X1 U8214 ( .A1(n6572), .A2(n6571), .ZN(n6573) );
  NAND2_X1 U8215 ( .A1(n9452), .A2(n6604), .ZN(n6576) );
  NAND2_X1 U8216 ( .A1(n9471), .A2(n6603), .ZN(n6575) );
  NAND2_X1 U8217 ( .A1(n6576), .A2(n6575), .ZN(n6577) );
  XNOR2_X1 U8218 ( .A(n6577), .B(n6423), .ZN(n6582) );
  AOI22_X1 U8219 ( .A1(n9452), .A2(n6603), .B1(n6407), .B2(n9471), .ZN(n6583)
         );
  XNOR2_X1 U8220 ( .A(n6582), .B(n6583), .ZN(n8917) );
  NAND2_X1 U8221 ( .A1(n9616), .A2(n6604), .ZN(n6579) );
  NAND2_X1 U8222 ( .A1(n9445), .A2(n6415), .ZN(n6578) );
  NAND2_X1 U8223 ( .A1(n6579), .A2(n6578), .ZN(n6580) );
  XNOR2_X1 U8224 ( .A(n6580), .B(n6423), .ZN(n6596) );
  AND2_X1 U8225 ( .A1(n9445), .A2(n6407), .ZN(n6581) );
  AOI21_X1 U8226 ( .B1(n9616), .B2(n6603), .A(n6581), .ZN(n6594) );
  XNOR2_X1 U8227 ( .A(n6596), .B(n6594), .ZN(n8990) );
  INV_X1 U8228 ( .A(n6582), .ZN(n6584) );
  NAND2_X1 U8229 ( .A1(n6584), .A2(n6583), .ZN(n8987) );
  NAND2_X1 U8230 ( .A1(n9420), .A2(n6604), .ZN(n6587) );
  NAND2_X1 U8231 ( .A1(n9435), .A2(n6415), .ZN(n6586) );
  NAND2_X1 U8232 ( .A1(n6587), .A2(n6586), .ZN(n6588) );
  XNOR2_X1 U8233 ( .A(n6588), .B(n6434), .ZN(n6591) );
  INV_X1 U8234 ( .A(n6591), .ZN(n6593) );
  AND2_X1 U8235 ( .A1(n9435), .A2(n6407), .ZN(n6589) );
  AOI21_X1 U8236 ( .B1(n9420), .B2(n6603), .A(n6589), .ZN(n6590) );
  INV_X1 U8237 ( .A(n6590), .ZN(n6592) );
  AOI21_X1 U8238 ( .B1(n6593), .B2(n6592), .A(n6614), .ZN(n6637) );
  INV_X1 U8239 ( .A(n6637), .ZN(n6598) );
  INV_X1 U8240 ( .A(n6594), .ZN(n6595) );
  NAND2_X1 U8241 ( .A1(n6596), .A2(n6595), .ZN(n6638) );
  INV_X1 U8242 ( .A(n6638), .ZN(n6597) );
  NAND2_X1 U8243 ( .A1(n9402), .A2(n6415), .ZN(n6600) );
  NAND2_X1 U8244 ( .A1(n9416), .A2(n6407), .ZN(n6599) );
  NAND2_X1 U8245 ( .A1(n6600), .A2(n6599), .ZN(n6602) );
  XNOR2_X1 U8246 ( .A(n6602), .B(n6601), .ZN(n6606) );
  AOI22_X1 U8247 ( .A1(n9402), .A2(n6604), .B1(n6603), .B2(n9416), .ZN(n6605)
         );
  XNOR2_X1 U8248 ( .A(n6606), .B(n6605), .ZN(n6615) );
  NAND2_X1 U8249 ( .A1(n10004), .A2(n6608), .ZN(n6609) );
  NOR2_X1 U8250 ( .A1(n6688), .A2(n6609), .ZN(n6613) );
  NOR2_X1 U8251 ( .A1(n6707), .A2(n6610), .ZN(n6612) );
  NAND3_X1 U8252 ( .A1(n6615), .A2(n8997), .A3(n6614), .ZN(n6632) );
  INV_X1 U8253 ( .A(n6688), .ZN(n9719) );
  OR2_X1 U8254 ( .A1(n6717), .A2(n9204), .ZN(n6895) );
  INV_X1 U8255 ( .A(n6895), .ZN(n6616) );
  NAND3_X1 U8256 ( .A1(n6620), .A2(n9719), .A3(n6616), .ZN(n6617) );
  OR2_X1 U8257 ( .A1(n6688), .A2(n9261), .ZN(n6618) );
  NOR2_X1 U8258 ( .A1(n6618), .A2(n7913), .ZN(n9270) );
  NAND2_X1 U8259 ( .A1(n9270), .A2(n6620), .ZN(n9001) );
  INV_X1 U8260 ( .A(n6618), .ZN(n6619) );
  AOI22_X1 U8261 ( .A1(n9276), .A2(n8999), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n6628) );
  INV_X1 U8262 ( .A(n6620), .ZN(n6622) );
  NAND2_X1 U8263 ( .A1(n6622), .A2(n6621), .ZN(n6624) );
  NAND2_X1 U8264 ( .A1(n6624), .A2(n6623), .ZN(n6812) );
  NAND2_X1 U8265 ( .A1(n6812), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6626) );
  INV_X1 U8266 ( .A(n6685), .ZN(n6625) );
  NAND2_X1 U8267 ( .A1(n6625), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9273) );
  NAND2_X1 U8268 ( .A1(n9401), .A2(n9004), .ZN(n6627) );
  OAI211_X1 U8269 ( .C1(n6629), .C2(n9001), .A(n6628), .B(n6627), .ZN(n6630)
         );
  AOI21_X1 U8270 ( .B1(n9402), .B2(n8972), .A(n6630), .ZN(n6631) );
  NAND2_X1 U8271 ( .A1(n6632), .A2(n6631), .ZN(n6633) );
  AOI21_X1 U8272 ( .B1(n6639), .B2(n6634), .A(n6633), .ZN(n6635) );
  NAND2_X1 U8273 ( .A1(n6636), .A2(n6635), .ZN(P1_U3220) );
  AOI21_X1 U8274 ( .B1(n8989), .B2(n6638), .A(n6637), .ZN(n6640) );
  OAI21_X1 U8275 ( .B1(n6640), .B2(n6639), .A(n8997), .ZN(n6646) );
  INV_X1 U8276 ( .A(n6641), .ZN(n9421) );
  AOI22_X1 U8277 ( .A1(n9421), .A2(n9004), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n6642) );
  OAI21_X1 U8278 ( .B1(n6643), .B2(n9001), .A(n6642), .ZN(n6644) );
  AOI21_X1 U8279 ( .B1(n8999), .B2(n9416), .A(n6644), .ZN(n6645) );
  NAND3_X1 U8280 ( .A1(n6646), .A2(n6645), .A3(n4899), .ZN(P1_U3214) );
  OR2_X2 U8281 ( .A1(n6811), .A2(n6647), .ZN(n9285) );
  INV_X1 U8282 ( .A(n6788), .ZN(n6648) );
  AOI211_X1 U8283 ( .C1(n6651), .C2(n6650), .A(n8974), .B(n6649), .ZN(n6657)
         );
  INV_X1 U8284 ( .A(n9004), .ZN(n8980) );
  INV_X1 U8285 ( .A(n7068), .ZN(n6652) );
  NOR2_X1 U8286 ( .A1(n8980), .A2(n6652), .ZN(n6656) );
  NOR2_X1 U8287 ( .A1(n9008), .A2(n9970), .ZN(n6655) );
  NAND2_X1 U8288 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9311) );
  NAND2_X1 U8289 ( .A1(n8999), .A2(n9281), .ZN(n6653) );
  OAI211_X1 U8290 ( .C1(n7077), .C2(n9001), .A(n9311), .B(n6653), .ZN(n6654)
         );
  OR4_X1 U8291 ( .A1(n6657), .A2(n6656), .A3(n6655), .A4(n6654), .ZN(P1_U3230)
         );
  INV_X1 U8292 ( .A(n6866), .ZN(n6658) );
  NAND2_X1 U8293 ( .A1(n6658), .A2(n6865), .ZN(n6971) );
  NAND2_X1 U8294 ( .A1(n6659), .A2(n6865), .ZN(n6660) );
  NAND2_X1 U8295 ( .A1(n6971), .A2(n6660), .ZN(n6970) );
  OR2_X1 U8296 ( .A1(n6970), .A2(n6661), .ZN(n6662) );
  NAND2_X1 U8297 ( .A1(n6662), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  AND2_X1 U8298 ( .A1(n4350), .A2(P2_U3151), .ZN(n8876) );
  NAND2_X1 U8299 ( .A1(n6663), .A2(P2_U3151), .ZN(n6665) );
  OAI222_X1 U8300 ( .A1(n8880), .A2(n6664), .B1(n8878), .B2(n6672), .C1(n10022), .C2(P2_U3151), .ZN(P2_U3293) );
  OAI222_X1 U8301 ( .A1(n8880), .A2(n6666), .B1(n8878), .B2(n6674), .C1(n7018), 
        .C2(P2_U3151), .ZN(P2_U3292) );
  OAI222_X1 U8302 ( .A1(n8880), .A2(n4923), .B1(n8878), .B2(n6684), .C1(n6956), 
        .C2(P2_U3151), .ZN(P2_U3294) );
  OAI222_X1 U8303 ( .A1(n7498), .A2(P2_U3151), .B1(n8878), .B2(n6670), .C1(
        n6667), .C2(n8880), .ZN(P2_U3291) );
  OAI222_X1 U8304 ( .A1(n7020), .A2(P2_U3151), .B1(n8878), .B2(n6682), .C1(
        n6668), .C2(n8880), .ZN(P2_U3290) );
  NAND2_X1 U8305 ( .A1(n4350), .A2(P1_U3086), .ZN(n9727) );
  OAI222_X1 U8306 ( .A1(n9729), .A2(n6671), .B1(n9727), .B2(n6670), .C1(
        P1_U3086), .C2(n9312), .ZN(P1_U3351) );
  OAI222_X1 U8307 ( .A1(n9729), .A2(n6673), .B1(n9727), .B2(n6672), .C1(
        P1_U3086), .C2(n6752), .ZN(P1_U3353) );
  OAI222_X1 U8308 ( .A1(n9729), .A2(n6675), .B1(n9727), .B2(n6674), .C1(
        P1_U3086), .C2(n6756), .ZN(P1_U3352) );
  INV_X1 U8309 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6676) );
  INV_X1 U8310 ( .A(n6764), .ZN(n9802) );
  OAI222_X1 U8311 ( .A1(n9729), .A2(n6676), .B1(n9727), .B2(n6678), .C1(
        P1_U3086), .C2(n9802), .ZN(P1_U3349) );
  OAI222_X1 U8312 ( .A1(n7419), .A2(P2_U3151), .B1(n8878), .B2(n6678), .C1(
        n6677), .C2(n8880), .ZN(P2_U3289) );
  INV_X1 U8313 ( .A(n9729), .ZN(n6839) );
  AOI22_X1 U8314 ( .A1(n9341), .A2(P1_STATE_REG_SCAN_IN), .B1(n6839), .B2(
        P2_DATAO_REG_7__SCAN_IN), .ZN(n6679) );
  OAI21_X1 U8315 ( .B1(n6681), .B2(n9727), .A(n6679), .ZN(P1_U3348) );
  OAI222_X1 U8316 ( .A1(n7403), .A2(P2_U3151), .B1(n8878), .B2(n6681), .C1(
        n6680), .C2(n8880), .ZN(P2_U3288) );
  INV_X1 U8317 ( .A(n9727), .ZN(n7948) );
  OAI222_X1 U8318 ( .A1(n9729), .A2(n6683), .B1(n9732), .B2(n6682), .C1(
        P1_U3086), .C2(n6761), .ZN(P1_U3350) );
  OAI222_X1 U8319 ( .A1(n9729), .A2(n4836), .B1(n9732), .B2(n6684), .C1(
        P1_U3086), .C2(n6753), .ZN(P1_U3354) );
  NAND2_X1 U8320 ( .A1(n9198), .A2(n6685), .ZN(n6687) );
  AND2_X1 U8321 ( .A1(n6687), .A2(n6686), .ZN(n6733) );
  INV_X1 U8322 ( .A(n6733), .ZN(n6689) );
  NAND2_X1 U8323 ( .A1(n6688), .A2(n9273), .ZN(n6734) );
  AND2_X1 U8324 ( .A1(n6689), .A2(n6734), .ZN(n9870) );
  NOR2_X1 U8325 ( .A1(n9870), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8326 ( .A(n7464), .ZN(n7454) );
  INV_X1 U8327 ( .A(n6690), .ZN(n6692) );
  OAI222_X1 U8328 ( .A1(n7454), .A2(P2_U3151), .B1(n8878), .B2(n6692), .C1(
        n6691), .C2(n8880), .ZN(P2_U3287) );
  INV_X1 U8329 ( .A(n6767), .ZN(n9759) );
  OAI222_X1 U8330 ( .A1(n9729), .A2(n6693), .B1(n9727), .B2(n6692), .C1(
        P1_U3086), .C2(n9759), .ZN(P1_U3347) );
  INV_X1 U8331 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9685) );
  NAND2_X1 U8332 ( .A1(n5684), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6695) );
  INV_X1 U8333 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9604) );
  OR2_X1 U8334 ( .A1(n5683), .A2(n9604), .ZN(n6694) );
  OAI211_X1 U8335 ( .C1(n5963), .C2(n9685), .A(n6695), .B(n6694), .ZN(n9389)
         );
  NAND2_X1 U8336 ( .A1(n9389), .A2(P1_U3973), .ZN(n6696) );
  OAI21_X1 U8337 ( .B1(P1_U3973), .B2(n6176), .A(n6696), .ZN(P1_U3585) );
  INV_X1 U8338 ( .A(n6697), .ZN(n6700) );
  AOI22_X1 U8339 ( .A1(n9764), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n6839), .ZN(n6698) );
  OAI21_X1 U8340 ( .B1(n6700), .B2(n9727), .A(n6698), .ZN(P1_U3346) );
  INV_X1 U8341 ( .A(n7455), .ZN(n7666) );
  OAI222_X1 U8342 ( .A1(P2_U3151), .A2(n7666), .B1(n8878), .B2(n6700), .C1(
        n6699), .C2(n8880), .ZN(P2_U3286) );
  INV_X1 U8343 ( .A(n6701), .ZN(n6704) );
  INV_X1 U8344 ( .A(n6770), .ZN(n9745) );
  INV_X1 U8345 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6702) );
  OAI222_X1 U8346 ( .A1(n9732), .A2(n6704), .B1(n9745), .B2(P1_U3086), .C1(
        n6702), .C2(n9729), .ZN(P1_U3345) );
  INV_X1 U8347 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6703) );
  OAI222_X1 U8348 ( .A1(P2_U3151), .A2(n7708), .B1(n8878), .B2(n6704), .C1(
        n6703), .C2(n8880), .ZN(P2_U3285) );
  INV_X1 U8349 ( .A(n6705), .ZN(n6723) );
  AOI22_X1 U8350 ( .A1(n7820), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n8876), .ZN(n6706) );
  OAI21_X1 U8351 ( .B1(n6723), .B2(n8878), .A(n6706), .ZN(P2_U3284) );
  INV_X1 U8352 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6790) );
  INV_X1 U8353 ( .A(n6707), .ZN(n6709) );
  AND2_X1 U8354 ( .A1(n6709), .A2(n6708), .ZN(n6710) );
  NAND2_X1 U8355 ( .A1(n6711), .A2(n6710), .ZN(n6719) );
  INV_X1 U8356 ( .A(n6712), .ZN(n6847) );
  NAND2_X1 U8357 ( .A1(n6713), .A2(n6813), .ZN(n9022) );
  AND2_X1 U8358 ( .A1(n6847), .A2(n9022), .ZN(n6726) );
  INV_X1 U8359 ( .A(n6714), .ZN(n6715) );
  INV_X1 U8360 ( .A(n6717), .ZN(n6729) );
  NOR3_X1 U8361 ( .A1(n6726), .A2(n6715), .A3(n6729), .ZN(n6716) );
  NOR2_X1 U8362 ( .A1(n7076), .A2(n7914), .ZN(n6728) );
  OAI21_X1 U8363 ( .B1(n6716), .B2(n6728), .A(n9598), .ZN(n6722) );
  INV_X1 U8364 ( .A(n9260), .ZN(n6718) );
  NOR4_X1 U8365 ( .A1(n6719), .A2(n6813), .A3(n6718), .A4(n6717), .ZN(n6720)
         );
  AOI21_X1 U8366 ( .B1(n9952), .B2(P1_REG3_REG_0__SCAN_IN), .A(n6720), .ZN(
        n6721) );
  OAI211_X1 U8367 ( .C1(n6790), .C2(n9598), .A(n6722), .B(n6721), .ZN(P1_U3293) );
  INV_X1 U8368 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6724) );
  INV_X1 U8369 ( .A(n6772), .ZN(n9817) );
  OAI222_X1 U8370 ( .A1(n9729), .A2(n6724), .B1(n9727), .B2(n6723), .C1(
        P1_U3086), .C2(n9817), .ZN(P1_U3344) );
  INV_X1 U8371 ( .A(n9366), .ZN(n6778) );
  INV_X1 U8372 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6725) );
  OAI222_X1 U8373 ( .A1(n9732), .A2(n6732), .B1(n6778), .B2(P1_U3086), .C1(
        n6725), .C2(n9729), .ZN(P1_U3343) );
  AOI21_X1 U8374 ( .B1(n9934), .B2(n9675), .A(n6726), .ZN(n6727) );
  AOI211_X1 U8375 ( .C1(n6729), .C2(n6843), .A(n6728), .B(n6727), .ZN(n9963)
         );
  NAND2_X1 U8376 ( .A1(n10019), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6730) );
  OAI21_X1 U8377 ( .B1(n9963), .B2(n10019), .A(n6730), .ZN(P1_U3522) );
  INV_X1 U8378 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6731) );
  OAI222_X1 U8379 ( .A1(P2_U3151), .A2(n8388), .B1(n6665), .B2(n6732), .C1(
        n6731), .C2(n8880), .ZN(P2_U3283) );
  NAND2_X1 U8380 ( .A1(n6734), .A2(n6733), .ZN(n9792) );
  OR2_X1 U8381 ( .A1(n4351), .A2(n8108), .ZN(n6735) );
  OR2_X1 U8382 ( .A1(n9792), .A2(n6735), .ZN(n9890) );
  INV_X1 U8383 ( .A(n9890), .ZN(n9885) );
  NOR2_X1 U8384 ( .A1(n9366), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6736) );
  AOI21_X1 U8385 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n9366), .A(n6736), .ZN(
        n6749) );
  INV_X1 U8386 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7389) );
  AOI22_X1 U8387 ( .A1(n6770), .A2(n7389), .B1(P1_REG2_REG_10__SCAN_IN), .B2(
        n9745), .ZN(n9736) );
  NOR2_X1 U8388 ( .A1(n9764), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6737) );
  AOI21_X1 U8389 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n9764), .A(n6737), .ZN(
        n9771) );
  INV_X1 U8390 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7087) );
  MUX2_X1 U8391 ( .A(n7087), .B(P1_REG2_REG_2__SCAN_IN), .S(n6752), .Z(n6798)
         );
  INV_X1 U8392 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7144) );
  MUX2_X1 U8393 ( .A(n7144), .B(P1_REG2_REG_1__SCAN_IN), .S(n6753), .Z(n9288)
         );
  NOR2_X1 U8394 ( .A1(n9789), .A2(n6790), .ZN(n9287) );
  NAND2_X1 U8395 ( .A1(n9288), .A2(n9287), .ZN(n9286) );
  INV_X1 U8396 ( .A(n6753), .ZN(n9292) );
  NAND2_X1 U8397 ( .A1(n9292), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6738) );
  NAND2_X1 U8398 ( .A1(n9286), .A2(n6738), .ZN(n6797) );
  NAND2_X1 U8399 ( .A1(n6798), .A2(n6797), .ZN(n6796) );
  INV_X1 U8400 ( .A(n6752), .ZN(n6802) );
  NAND2_X1 U8401 ( .A1(n6802), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6739) );
  NAND2_X1 U8402 ( .A1(n6796), .A2(n6739), .ZN(n9305) );
  XNOR2_X1 U8403 ( .A(n6756), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9306) );
  NAND2_X1 U8404 ( .A1(n9305), .A2(n9306), .ZN(n9304) );
  INV_X1 U8405 ( .A(n6756), .ZN(n9300) );
  NAND2_X1 U8406 ( .A1(n9300), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6740) );
  NAND2_X1 U8407 ( .A1(n9304), .A2(n6740), .ZN(n9315) );
  XNOR2_X1 U8408 ( .A(n9312), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n9316) );
  NAND2_X1 U8409 ( .A1(n9315), .A2(n9316), .ZN(n9314) );
  INV_X1 U8410 ( .A(n9312), .ZN(n6758) );
  NAND2_X1 U8411 ( .A1(n6758), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6741) );
  NAND2_X1 U8412 ( .A1(n9314), .A2(n6741), .ZN(n9332) );
  XNOR2_X1 U8413 ( .A(n6761), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n9333) );
  NAND2_X1 U8414 ( .A1(n9332), .A2(n9333), .ZN(n9331) );
  INV_X1 U8415 ( .A(n6761), .ZN(n9327) );
  NAND2_X1 U8416 ( .A1(n9327), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6742) );
  NAND2_X1 U8417 ( .A1(n9331), .A2(n6742), .ZN(n9795) );
  INV_X1 U8418 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6743) );
  XNOR2_X1 U8419 ( .A(n6764), .B(n6743), .ZN(n9796) );
  NAND2_X1 U8420 ( .A1(n9795), .A2(n9796), .ZN(n9794) );
  NAND2_X1 U8421 ( .A1(n6764), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6744) );
  NAND2_X1 U8422 ( .A1(n9794), .A2(n6744), .ZN(n9343) );
  INV_X1 U8423 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7482) );
  MUX2_X1 U8424 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n7482), .S(n9341), .Z(n9344)
         );
  NAND2_X1 U8425 ( .A1(n9343), .A2(n9344), .ZN(n9342) );
  NAND2_X1 U8426 ( .A1(n9341), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6745) );
  NAND2_X1 U8427 ( .A1(n9342), .A2(n6745), .ZN(n9752) );
  INV_X1 U8428 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6746) );
  MUX2_X1 U8429 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n6746), .S(n6767), .Z(n9753)
         );
  AND2_X1 U8430 ( .A1(n9752), .A2(n9753), .ZN(n9750) );
  AOI21_X1 U8431 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n6767), .A(n9750), .ZN(
        n9770) );
  NAND2_X1 U8432 ( .A1(n9771), .A2(n9770), .ZN(n9769) );
  OAI21_X1 U8433 ( .B1(n9764), .B2(P1_REG2_REG_9__SCAN_IN), .A(n9769), .ZN(
        n9737) );
  NOR2_X1 U8434 ( .A1(n9736), .A2(n9737), .ZN(n9735) );
  AOI21_X1 U8435 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n6770), .A(n9735), .ZN(
        n9808) );
  INV_X1 U8436 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6747) );
  AOI22_X1 U8437 ( .A1(n6772), .A2(n6747), .B1(P1_REG2_REG_11__SCAN_IN), .B2(
        n9817), .ZN(n9809) );
  NOR2_X1 U8438 ( .A1(n9808), .A2(n9809), .ZN(n9807) );
  AOI21_X1 U8439 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n6772), .A(n9807), .ZN(
        n6748) );
  NAND2_X1 U8440 ( .A1(n6749), .A2(n6748), .ZN(n9352) );
  OAI21_X1 U8441 ( .B1(n6749), .B2(n6748), .A(n9352), .ZN(n6780) );
  INV_X1 U8442 ( .A(n4351), .ZN(n6793) );
  OR2_X1 U8443 ( .A1(n9792), .A2(n6793), .ZN(n9899) );
  MUX2_X1 U8444 ( .A(n6750), .B(P1_REG1_REG_10__SCAN_IN), .S(n6770), .Z(n9741)
         );
  OR2_X1 U8445 ( .A1(n9764), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6769) );
  NOR2_X1 U8446 ( .A1(n9764), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6751) );
  AOI21_X1 U8447 ( .B1(n9764), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6751), .ZN(
        n9766) );
  INV_X1 U8448 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10011) );
  MUX2_X1 U8449 ( .A(n10011), .B(P1_REG1_REG_2__SCAN_IN), .S(n6752), .Z(n6801)
         );
  MUX2_X1 U8450 ( .A(n5650), .B(P1_REG1_REG_1__SCAN_IN), .S(n6753), .Z(n9291)
         );
  AND2_X1 U8451 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9290) );
  NAND2_X1 U8452 ( .A1(n9291), .A2(n9290), .ZN(n9289) );
  NAND2_X1 U8453 ( .A1(n9292), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6754) );
  NAND2_X1 U8454 ( .A1(n9289), .A2(n6754), .ZN(n6800) );
  NAND2_X1 U8455 ( .A1(n6801), .A2(n6800), .ZN(n6799) );
  NAND2_X1 U8456 ( .A1(n6802), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6755) );
  NAND2_X1 U8457 ( .A1(n6799), .A2(n6755), .ZN(n9302) );
  XNOR2_X1 U8458 ( .A(n6756), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n9303) );
  NAND2_X1 U8459 ( .A1(n9302), .A2(n9303), .ZN(n9301) );
  NAND2_X1 U8460 ( .A1(n9300), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6757) );
  NAND2_X1 U8461 ( .A1(n9301), .A2(n6757), .ZN(n9318) );
  XNOR2_X1 U8462 ( .A(n9312), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n9319) );
  NAND2_X1 U8463 ( .A1(n9318), .A2(n9319), .ZN(n9317) );
  NAND2_X1 U8464 ( .A1(n6758), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6759) );
  NAND2_X1 U8465 ( .A1(n9317), .A2(n6759), .ZN(n9329) );
  XNOR2_X1 U8466 ( .A(n6761), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n9330) );
  NAND2_X1 U8467 ( .A1(n9329), .A2(n9330), .ZN(n9328) );
  OR2_X1 U8468 ( .A1(n6761), .A2(n6760), .ZN(n6762) );
  NAND2_X1 U8469 ( .A1(n9328), .A2(n6762), .ZN(n9798) );
  XNOR2_X1 U8470 ( .A(n6764), .B(n6763), .ZN(n9799) );
  NAND2_X1 U8471 ( .A1(n9798), .A2(n9799), .ZN(n9797) );
  NAND2_X1 U8472 ( .A1(n6764), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6765) );
  NAND2_X1 U8473 ( .A1(n9797), .A2(n6765), .ZN(n9346) );
  MUX2_X1 U8474 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n5748), .S(n9341), .Z(n9347)
         );
  NAND2_X1 U8475 ( .A1(n9346), .A2(n9347), .ZN(n9345) );
  NAND2_X1 U8476 ( .A1(n9341), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6766) );
  NAND2_X1 U8477 ( .A1(n9345), .A2(n6766), .ZN(n9755) );
  MUX2_X1 U8478 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n5763), .S(n6767), .Z(n9756)
         );
  NAND2_X1 U8479 ( .A1(n9755), .A2(n9756), .ZN(n9754) );
  NAND2_X1 U8480 ( .A1(n6767), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6768) );
  AND2_X1 U8481 ( .A1(n9754), .A2(n6768), .ZN(n9767) );
  NAND2_X1 U8482 ( .A1(n9766), .A2(n9767), .ZN(n9765) );
  NAND2_X1 U8483 ( .A1(n6769), .A2(n9765), .ZN(n9740) );
  NOR2_X1 U8484 ( .A1(n9741), .A2(n9740), .ZN(n9739) );
  AOI21_X1 U8485 ( .B1(n6770), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9739), .ZN(
        n9812) );
  MUX2_X1 U8486 ( .A(n6771), .B(P1_REG1_REG_11__SCAN_IN), .S(n6772), .Z(n9813)
         );
  NOR2_X1 U8487 ( .A1(n9812), .A2(n9813), .ZN(n9811) );
  AOI21_X1 U8488 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n6772), .A(n9811), .ZN(
        n6774) );
  AOI22_X1 U8489 ( .A1(n9366), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n5822), .B2(
        n6778), .ZN(n6773) );
  NAND2_X1 U8490 ( .A1(n6774), .A2(n6773), .ZN(n9365) );
  OAI21_X1 U8491 ( .B1(n6774), .B2(n6773), .A(n9365), .ZN(n6775) );
  INV_X1 U8492 ( .A(n8108), .ZN(n9788) );
  INV_X1 U8493 ( .A(n9851), .ZN(n9893) );
  NAND2_X1 U8494 ( .A1(n6775), .A2(n9893), .ZN(n6777) );
  AND2_X1 U8495 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7759) );
  AOI21_X1 U8496 ( .B1(n9870), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n7759), .ZN(
        n6776) );
  OAI211_X1 U8497 ( .C1(n9899), .C2(n6778), .A(n6777), .B(n6776), .ZN(n6779)
         );
  AOI21_X1 U8498 ( .B1(n9885), .B2(n6780), .A(n6779), .ZN(n6781) );
  INV_X1 U8499 ( .A(n6781), .ZN(P1_U3255) );
  INV_X1 U8500 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6785) );
  INV_X1 U8501 ( .A(n6783), .ZN(n6784) );
  AOI22_X1 U8502 ( .A1(n6818), .A2(n6785), .B1(n6788), .B2(n6784), .ZN(
        P2_U3377) );
  INV_X1 U8503 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6789) );
  INV_X1 U8504 ( .A(n6786), .ZN(n6787) );
  AOI22_X1 U8505 ( .A1(n6818), .A2(n6789), .B1(n6788), .B2(n6787), .ZN(
        P2_U3376) );
  AOI21_X1 U8506 ( .B1(n9788), .B2(n6790), .A(n4351), .ZN(n9787) );
  XNOR2_X1 U8507 ( .A(n6792), .B(n6791), .ZN(n6817) );
  MUX2_X1 U8508 ( .A(n9287), .B(n6817), .S(n8108), .Z(n6794) );
  NAND2_X1 U8509 ( .A1(n6794), .A2(n6793), .ZN(n6795) );
  OAI211_X1 U8510 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n9787), .A(n6795), .B(
        P1_U3973), .ZN(n9323) );
  INV_X1 U8511 ( .A(n9323), .ZN(n6808) );
  OAI211_X1 U8512 ( .C1(n6798), .C2(n6797), .A(n9885), .B(n6796), .ZN(n6806)
         );
  OAI211_X1 U8513 ( .C1(n6801), .C2(n6800), .A(n9893), .B(n6799), .ZN(n6805)
         );
  AOI22_X1 U8514 ( .A1(n9870), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n6804) );
  NAND2_X1 U8515 ( .A1(n9882), .A2(n6802), .ZN(n6803) );
  NAND4_X1 U8516 ( .A1(n6806), .A2(n6805), .A3(n6804), .A4(n6803), .ZN(n6807)
         );
  OR2_X1 U8517 ( .A1(n6808), .A2(n6807), .ZN(P1_U3245) );
  INV_X1 U8518 ( .A(n6809), .ZN(n6820) );
  AOI22_X1 U8519 ( .A1(n9830), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n6839), .ZN(n6810) );
  OAI21_X1 U8520 ( .B1(n6820), .B2(n9727), .A(n6810), .ZN(P1_U3342) );
  NOR2_X1 U8521 ( .A1(n6812), .A2(n6811), .ZN(n6832) );
  INV_X1 U8522 ( .A(n6832), .ZN(n6815) );
  INV_X1 U8523 ( .A(n8999), .ZN(n8981) );
  OAI22_X1 U8524 ( .A1(n8981), .A2(n7076), .B1(n9008), .B2(n6813), .ZN(n6814)
         );
  AOI21_X1 U8525 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n6815), .A(n6814), .ZN(
        n6816) );
  OAI21_X1 U8526 ( .B1(n6817), .B2(n8974), .A(n6816), .ZN(P1_U3232) );
  AND2_X1 U8527 ( .A1(n6818), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8528 ( .A1(n6818), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8529 ( .A1(n6818), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8530 ( .A1(n6818), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8531 ( .A1(n6818), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8532 ( .A1(n6818), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8533 ( .A1(n6818), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8534 ( .A1(n6818), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8535 ( .A1(n6818), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8536 ( .A1(n6818), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8537 ( .A1(n6818), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8538 ( .A1(n6818), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8539 ( .A1(n6818), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8540 ( .A1(n6818), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8541 ( .A1(n6818), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8542 ( .A1(n6818), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8543 ( .A1(n6818), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8544 ( .A1(n6818), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8545 ( .A1(n6818), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8546 ( .A1(n6818), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8547 ( .A1(n6818), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8548 ( .A1(n6818), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8549 ( .A1(n6818), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8550 ( .A1(n6818), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8551 ( .A1(n6818), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8552 ( .A1(n6818), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8553 ( .A1(n6818), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8554 ( .A1(n6818), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8555 ( .A1(n6818), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8556 ( .A1(n6818), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  INV_X1 U8557 ( .A(n8403), .ZN(n8389) );
  INV_X1 U8558 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6819) );
  OAI222_X1 U8559 ( .A1(n8389), .A2(P2_U3151), .B1(n6665), .B2(n6820), .C1(
        n6819), .C2(n8880), .ZN(P2_U3282) );
  INV_X1 U8560 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7086) );
  INV_X1 U8561 ( .A(n6821), .ZN(n6825) );
  NOR3_X1 U8562 ( .A1(n6829), .A2(n6823), .A3(n6822), .ZN(n6824) );
  OAI21_X1 U8563 ( .B1(n6825), .B2(n6824), .A(n8997), .ZN(n6828) );
  OAI22_X1 U8564 ( .A1(n7077), .A2(n8981), .B1(n7076), .B2(n9001), .ZN(n6826)
         );
  AOI21_X1 U8565 ( .B1(n7089), .B2(n8972), .A(n6826), .ZN(n6827) );
  OAI211_X1 U8566 ( .C1(n6832), .C2(n7086), .A(n6828), .B(n6827), .ZN(P1_U3237) );
  AOI21_X1 U8567 ( .B1(n6831), .B2(n6830), .A(n6829), .ZN(n6837) );
  INV_X1 U8568 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7143) );
  NOR2_X1 U8569 ( .A1(n6832), .A2(n7143), .ZN(n6834) );
  OAI22_X1 U8570 ( .A1(n8981), .A2(n6850), .B1(n6405), .B2(n9001), .ZN(n6833)
         );
  AOI211_X1 U8571 ( .C1(n6835), .C2(n8972), .A(n6834), .B(n6833), .ZN(n6836)
         );
  OAI21_X1 U8572 ( .B1(n6837), .B2(n8974), .A(n6836), .ZN(P1_U3222) );
  INV_X1 U8573 ( .A(n6838), .ZN(n6856) );
  AOI22_X1 U8574 ( .A1(n9835), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n6839), .ZN(n6840) );
  OAI21_X1 U8575 ( .B1(n6856), .B2(n9727), .A(n6840), .ZN(P1_U3341) );
  OAI21_X1 U8576 ( .B1(n6842), .B2(n6848), .A(n6841), .ZN(n7141) );
  AOI21_X1 U8577 ( .B1(n6843), .B2(n6835), .A(n9590), .ZN(n6844) );
  AND2_X1 U8578 ( .A1(n6844), .A2(n7083), .ZN(n7147) );
  INV_X1 U8579 ( .A(n6845), .ZN(n6846) );
  AOI21_X1 U8580 ( .B1(n6848), .B2(n6847), .A(n6846), .ZN(n6849) );
  OAI222_X1 U8581 ( .A1(n7914), .A2(n6850), .B1(n7913), .B2(n6405), .C1(n9934), 
        .C2(n6849), .ZN(n7142) );
  AOI211_X1 U8582 ( .C1(n10007), .C2(n7141), .A(n7147), .B(n7142), .ZN(n6854)
         );
  OAI22_X1 U8583 ( .A1(n9709), .A2(n6060), .B1(n10010), .B2(n5651), .ZN(n6851)
         );
  INV_X1 U8584 ( .A(n6851), .ZN(n6852) );
  OAI21_X1 U8585 ( .B1(n6854), .B2(n10009), .A(n6852), .ZN(P1_U3456) );
  AOI22_X1 U8586 ( .A1(n6101), .A2(n6835), .B1(n10019), .B2(
        P1_REG1_REG_1__SCAN_IN), .ZN(n6853) );
  OAI21_X1 U8587 ( .B1(n6854), .B2(n10019), .A(n6853), .ZN(P1_U3523) );
  INV_X1 U8588 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6855) );
  OAI222_X1 U8589 ( .A1(n8427), .A2(P2_U3151), .B1(n6665), .B2(n6856), .C1(
        n6855), .C2(n8880), .ZN(P2_U3281) );
  INV_X1 U8590 ( .A(n6857), .ZN(n6860) );
  AOI22_X1 U8591 ( .A1(n8458), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n8876), .ZN(n6858) );
  OAI21_X1 U8592 ( .B1(n6860), .B2(n8878), .A(n6858), .ZN(P2_U3280) );
  INV_X1 U8593 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6859) );
  OAI222_X1 U8594 ( .A1(n9732), .A2(n6860), .B1(n9368), .B2(P1_U3086), .C1(
        n6859), .C2(n9729), .ZN(P1_U3340) );
  NAND2_X1 U8595 ( .A1(n6862), .A2(n6861), .ZN(n6869) );
  INV_X1 U8596 ( .A(n6863), .ZN(n6884) );
  NAND3_X1 U8597 ( .A1(n6866), .A2(n6865), .A3(n6864), .ZN(n6867) );
  AOI21_X1 U8598 ( .B1(n6872), .B2(n6884), .A(n6867), .ZN(n6868) );
  NAND2_X1 U8599 ( .A1(n6869), .A2(n6868), .ZN(n6870) );
  NAND2_X1 U8600 ( .A1(n6870), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6874) );
  NAND2_X1 U8601 ( .A1(n6872), .A2(n6871), .ZN(n6873) );
  NOR2_X1 U8602 ( .A1(n8335), .A2(P2_U3151), .ZN(n6925) );
  INV_X1 U8603 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6890) );
  NOR2_X1 U8604 ( .A1(n6876), .A2(n6875), .ZN(n6912) );
  INV_X1 U8605 ( .A(n6911), .ZN(n6877) );
  OR2_X1 U8606 ( .A1(n6883), .A2(n8745), .ZN(n6881) );
  OR2_X1 U8607 ( .A1(n6883), .A2(n6882), .ZN(n6887) );
  NAND2_X1 U8608 ( .A1(n6885), .A2(n6884), .ZN(n6886) );
  OAI22_X1 U8609 ( .A1(n8354), .A2(n7730), .B1(n8342), .B2(n7728), .ZN(n6888)
         );
  AOI21_X1 U8610 ( .B1(n8327), .B2(n8371), .A(n6888), .ZN(n6889) );
  OAI21_X1 U8611 ( .B1(n6925), .B2(n6890), .A(n6889), .ZN(P2_U3172) );
  XNOR2_X1 U8612 ( .A(n9047), .B(n9019), .ZN(n6891) );
  OAI222_X1 U8613 ( .A1(n7914), .A2(n7478), .B1(n6891), .B2(n9934), .C1(n7913), 
        .C2(n6939), .ZN(n7094) );
  INV_X1 U8614 ( .A(n7094), .ZN(n6902) );
  INV_X2 U8615 ( .A(n9598), .ZN(n9593) );
  AND2_X1 U8616 ( .A1(n7910), .A2(n7917), .ZN(n6892) );
  OAI21_X1 U8617 ( .B1(n6894), .B2(n9019), .A(n6893), .ZN(n7096) );
  INV_X1 U8618 ( .A(n6896), .ZN(n7066) );
  INV_X1 U8619 ( .A(n6897), .ZN(n7111) );
  AOI211_X1 U8620 ( .C1(n6941), .C2(n7066), .A(n9590), .B(n7111), .ZN(n7095)
         );
  NAND2_X1 U8621 ( .A1(n7095), .A2(n9949), .ZN(n6899) );
  AOI22_X1 U8622 ( .A1(n9593), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n6936), .B2(
        n9952), .ZN(n6898) );
  OAI211_X1 U8623 ( .C1(n7099), .C2(n9955), .A(n6899), .B(n6898), .ZN(n6900)
         );
  AOI21_X1 U8624 ( .B1(n9959), .B2(n7096), .A(n6900), .ZN(n6901) );
  OAI21_X1 U8625 ( .B1(n6902), .B2(n9593), .A(n6901), .ZN(P1_U3288) );
  INV_X1 U8626 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10063) );
  OAI211_X2 U8627 ( .C1(n6905), .C2(n6904), .A(n7570), .B(n6903), .ZN(n6906)
         );
  XNOR2_X1 U8628 ( .A(n6906), .B(n5099), .ZN(n7359) );
  XNOR2_X1 U8629 ( .A(n7359), .B(n5101), .ZN(n6909) );
  OAI21_X1 U8630 ( .B1(n8173), .B2(n7375), .A(n7042), .ZN(n6917) );
  NAND2_X1 U8631 ( .A1(n6908), .A2(n6909), .ZN(n7360) );
  OAI21_X1 U8632 ( .B1(n6909), .B2(n6908), .A(n7360), .ZN(n6910) );
  NAND2_X1 U8633 ( .A1(n6910), .A2(n8321), .ZN(n6915) );
  OAI22_X1 U8634 ( .A1(n7630), .A2(n8324), .B1(n8354), .B2(n10062), .ZN(n6913)
         );
  AOI21_X1 U8635 ( .B1(n8327), .B2(n8370), .A(n6913), .ZN(n6914) );
  OAI211_X1 U8636 ( .C1(n6925), .C2(n10063), .A(n6915), .B(n6914), .ZN(
        P2_U3177) );
  INV_X1 U8637 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6924) );
  OAI21_X1 U8638 ( .B1(n6918), .B2(n6917), .A(n6916), .ZN(n6919) );
  NAND2_X1 U8639 ( .A1(n6919), .A2(n8321), .ZN(n6923) );
  OAI22_X1 U8640 ( .A1(n6920), .A2(n8324), .B1(n8354), .B2(n7905), .ZN(n6921)
         );
  AOI21_X1 U8641 ( .B1(n8327), .B2(n5101), .A(n6921), .ZN(n6922) );
  OAI211_X1 U8642 ( .C1(n6925), .C2(n6924), .A(n6923), .B(n6922), .ZN(P2_U3162) );
  INV_X1 U8643 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6927) );
  INV_X1 U8644 ( .A(n6926), .ZN(n6929) );
  INV_X1 U8645 ( .A(n9874), .ZN(n9362) );
  OAI222_X1 U8646 ( .A1(n9729), .A2(n6927), .B1(n9732), .B2(n6929), .C1(
        P1_U3086), .C2(n9362), .ZN(P1_U3339) );
  INV_X1 U8647 ( .A(n8461), .ZN(n8481) );
  INV_X1 U8648 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6928) );
  OAI222_X1 U8649 ( .A1(n8481), .A2(P2_U3151), .B1(n6665), .B2(n6929), .C1(
        n6928), .C2(n8880), .ZN(P2_U3279) );
  INV_X1 U8650 ( .A(n6930), .ZN(n6932) );
  NAND2_X1 U8651 ( .A1(n6932), .A2(n6931), .ZN(n6934) );
  XNOR2_X1 U8652 ( .A(n6934), .B(n6933), .ZN(n6943) );
  NAND2_X1 U8653 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9324) );
  INV_X1 U8654 ( .A(n9324), .ZN(n6935) );
  AOI21_X1 U8655 ( .B1(n8999), .B2(n9280), .A(n6935), .ZN(n6938) );
  NAND2_X1 U8656 ( .A1(n9004), .A2(n6936), .ZN(n6937) );
  OAI211_X1 U8657 ( .C1(n6939), .C2(n9001), .A(n6938), .B(n6937), .ZN(n6940)
         );
  AOI21_X1 U8658 ( .B1(n6941), .B2(n8972), .A(n6940), .ZN(n6942) );
  OAI21_X1 U8659 ( .B1(n6943), .B2(n8974), .A(n6942), .ZN(P1_U3227) );
  OAI21_X1 U8660 ( .B1(n6945), .B2(n6946), .A(n6944), .ZN(n7703) );
  XNOR2_X1 U8661 ( .A(n6947), .B(n6946), .ZN(n6948) );
  OAI222_X1 U8662 ( .A1(n8711), .A2(n7614), .B1(n8669), .B2(n5100), .C1(n8666), 
        .C2(n6948), .ZN(n7700) );
  AOI21_X1 U8663 ( .B1(n8794), .B2(n7703), .A(n7700), .ZN(n7926) );
  INV_X1 U8664 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6949) );
  OAI22_X1 U8665 ( .A1(n8841), .A2(n7699), .B1(n6949), .B2(n10088), .ZN(n6950)
         );
  INV_X1 U8666 ( .A(n6950), .ZN(n6951) );
  OAI21_X1 U8667 ( .B1(n7926), .B2(n10091), .A(n6951), .ZN(P2_U3399) );
  NAND2_X1 U8668 ( .A1(n8512), .A2(n6968), .ZN(n8542) );
  MUX2_X1 U8669 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n8529), .Z(n6977) );
  XNOR2_X1 U8670 ( .A(n6956), .B(n6977), .ZN(n6979) );
  MUX2_X1 U8671 ( .A(P2_REG2_REG_0__SCAN_IN), .B(P2_REG1_REG_0__SCAN_IN), .S(
        n8529), .Z(n7125) );
  INV_X1 U8672 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7131) );
  NOR2_X1 U8673 ( .A1(n7125), .A2(n7131), .ZN(n7124) );
  XNOR2_X1 U8674 ( .A(n6979), .B(n7124), .ZN(n6976) );
  INV_X1 U8675 ( .A(n6971), .ZN(n6952) );
  NOR2_X2 U8676 ( .A1(P2_U3150), .A2(n6952), .ZN(n10045) );
  NAND2_X1 U8677 ( .A1(n6953), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8106) );
  NOR2_X1 U8678 ( .A1(n7127), .A2(n8529), .ZN(n10056) );
  INV_X1 U8679 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6954) );
  NOR2_X1 U8680 ( .A1(n6954), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6955) );
  NAND2_X1 U8681 ( .A1(n6961), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7015) );
  INV_X1 U8682 ( .A(n7016), .ZN(n6957) );
  AOI21_X1 U8683 ( .B1(n7573), .B2(n6958), .A(n6957), .ZN(n6966) );
  INV_X1 U8684 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7904) );
  NOR2_X1 U8685 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(n6960), .ZN(n6962) );
  NAND2_X1 U8686 ( .A1(n6961), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6997) );
  NOR2_X1 U8687 ( .A1(n6963), .A2(n7904), .ZN(n6999) );
  AOI21_X1 U8688 ( .B1(n7904), .B2(n6963), .A(n6999), .ZN(n6965) );
  INV_X1 U8689 ( .A(n7127), .ZN(n6964) );
  NAND2_X1 U8690 ( .A1(n6964), .A2(n8529), .ZN(n10032) );
  OAI22_X1 U8691 ( .A1(n8486), .A2(n6966), .B1(n6965), .B2(n10032), .ZN(n6967)
         );
  AOI21_X1 U8692 ( .B1(n10045), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n6967), .ZN(
        n6975) );
  NOR2_X1 U8693 ( .A1(n8529), .A2(P2_U3151), .ZN(n8071) );
  NAND2_X1 U8694 ( .A1(n8071), .A2(n6968), .ZN(n6969) );
  OR2_X1 U8695 ( .A1(n6970), .A2(n6969), .ZN(n6973) );
  OR2_X1 U8696 ( .A1(n6971), .A2(n8106), .ZN(n6972) );
  NAND2_X1 U8697 ( .A1(n6973), .A2(n6972), .ZN(n10047) );
  AOI22_X1 U8698 ( .A1(n10047), .A2(n6959), .B1(P2_U3151), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n6974) );
  OAI211_X1 U8699 ( .C1(n8542), .C2(n6976), .A(n6975), .B(n6974), .ZN(P2_U3183) );
  INV_X1 U8700 ( .A(n7498), .ZN(n6985) );
  MUX2_X1 U8701 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8529), .Z(n6983) );
  INV_X1 U8702 ( .A(n6983), .ZN(n6984) );
  INV_X1 U8703 ( .A(n6977), .ZN(n6978) );
  MUX2_X1 U8704 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8529), .Z(n6980) );
  XOR2_X1 U8705 ( .A(n10022), .B(n6980), .Z(n10037) );
  MUX2_X1 U8706 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8529), .Z(n6981) );
  XOR2_X1 U8707 ( .A(n7018), .B(n6981), .Z(n10049) );
  NAND2_X1 U8708 ( .A1(n10050), .A2(n10049), .ZN(n10048) );
  INV_X1 U8709 ( .A(n6981), .ZN(n6982) );
  INV_X1 U8710 ( .A(n7018), .ZN(n10046) );
  NAND2_X1 U8711 ( .A1(n6982), .A2(n10046), .ZN(n7502) );
  XOR2_X1 U8712 ( .A(n7498), .B(n6983), .Z(n7504) );
  NAND3_X1 U8713 ( .A1(n10048), .A2(n7502), .A3(n7504), .ZN(n7503) );
  OAI21_X1 U8714 ( .B1(n6985), .B2(n6984), .A(n7503), .ZN(n7442) );
  MUX2_X1 U8715 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8529), .Z(n6986) );
  INV_X1 U8716 ( .A(n7020), .ZN(n7441) );
  XNOR2_X1 U8717 ( .A(n6986), .B(n7441), .ZN(n7443) );
  MUX2_X1 U8718 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8529), .Z(n6987) );
  NOR2_X1 U8719 ( .A1(n6987), .A2(n7419), .ZN(n6988) );
  AOI21_X1 U8720 ( .B1(n6987), .B2(n7419), .A(n6988), .ZN(n7424) );
  NAND2_X1 U8721 ( .A1(n7425), .A2(n7424), .ZN(n7423) );
  INV_X1 U8722 ( .A(n6988), .ZN(n7406) );
  INV_X1 U8723 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6989) );
  MUX2_X1 U8724 ( .A(n4708), .B(n6989), .S(n8529), .Z(n6990) );
  INV_X1 U8725 ( .A(n7403), .ZN(n7007) );
  NAND2_X1 U8726 ( .A1(n6990), .A2(n7007), .ZN(n6993) );
  INV_X1 U8727 ( .A(n6990), .ZN(n6991) );
  NAND2_X1 U8728 ( .A1(n6991), .A2(n7403), .ZN(n6992) );
  NAND2_X1 U8729 ( .A1(n6993), .A2(n6992), .ZN(n7405) );
  AOI21_X1 U8730 ( .B1(n7423), .B2(n7406), .A(n7405), .ZN(n7408) );
  INV_X1 U8731 ( .A(n6993), .ZN(n6994) );
  MUX2_X1 U8732 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8529), .Z(n7461) );
  XOR2_X1 U8733 ( .A(n7464), .B(n7461), .Z(n6995) );
  NOR2_X1 U8734 ( .A1(n6996), .A2(n6995), .ZN(n7462) );
  AOI21_X1 U8735 ( .B1(n6996), .B2(n6995), .A(n7462), .ZN(n7032) );
  INV_X1 U8736 ( .A(n6997), .ZN(n6998) );
  NOR2_X1 U8737 ( .A1(n6999), .A2(n6998), .ZN(n10026) );
  INV_X1 U8738 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7000) );
  MUX2_X1 U8739 ( .A(n7000), .B(P2_REG1_REG_2__SCAN_IN), .S(n10022), .Z(n10025) );
  AOI21_X1 U8740 ( .B1(P2_REG1_REG_2__SCAN_IN), .B2(n10022), .A(n10024), .ZN(
        n7001) );
  NOR2_X1 U8741 ( .A1(n7001), .A2(n10046), .ZN(n7002) );
  AOI21_X1 U8742 ( .B1(n7001), .B2(n10046), .A(n7002), .ZN(n10042) );
  INV_X1 U8743 ( .A(n7002), .ZN(n7494) );
  INV_X1 U8744 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7003) );
  MUX2_X1 U8745 ( .A(n7003), .B(P2_REG1_REG_4__SCAN_IN), .S(n7498), .Z(n7495)
         );
  AOI21_X1 U8746 ( .B1(n10041), .B2(n7494), .A(n7495), .ZN(n7493) );
  AOI21_X1 U8747 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(n7498), .A(n7493), .ZN(
        n7004) );
  INV_X1 U8748 ( .A(n7006), .ZN(n7411) );
  XNOR2_X1 U8749 ( .A(n7419), .B(P2_REG1_REG_6__SCAN_IN), .ZN(n7412) );
  AOI21_X1 U8750 ( .B1(n7008), .B2(n7007), .A(n7009), .ZN(n7397) );
  NAND2_X1 U8751 ( .A1(n7397), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7396) );
  INV_X1 U8752 ( .A(n7009), .ZN(n7011) );
  INV_X1 U8753 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7010) );
  XNOR2_X1 U8754 ( .A(n7464), .B(n7010), .ZN(n7012) );
  AOI21_X1 U8755 ( .B1(n7396), .B2(n7011), .A(n7012), .ZN(n7453) );
  INV_X1 U8756 ( .A(n7453), .ZN(n7014) );
  NAND3_X1 U8757 ( .A1(n7396), .A2(n7012), .A3(n7011), .ZN(n7013) );
  AOI21_X1 U8758 ( .B1(n7014), .B2(n7013), .A(n10032), .ZN(n7030) );
  MUX2_X1 U8759 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n5083), .S(n10022), .Z(n10029) );
  NAND2_X1 U8760 ( .A1(n7016), .A2(n7015), .ZN(n10028) );
  NAND2_X1 U8761 ( .A1(n10029), .A2(n10028), .ZN(n10027) );
  NAND2_X1 U8762 ( .A1(n10022), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7017) );
  NAND2_X1 U8763 ( .A1(n10053), .A2(n7489), .ZN(n7019) );
  MUX2_X1 U8764 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n5122), .S(n7498), .Z(n7488)
         );
  NAND2_X1 U8765 ( .A1(n7434), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7435) );
  NAND2_X1 U8766 ( .A1(n7435), .A2(n7415), .ZN(n7021) );
  INV_X1 U8767 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7590) );
  XNOR2_X1 U8768 ( .A(n7419), .B(n7590), .ZN(n7414) );
  NAND2_X1 U8769 ( .A1(n7021), .A2(n7414), .ZN(n7418) );
  NAND2_X1 U8770 ( .A1(n7419), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7022) );
  NAND2_X1 U8771 ( .A1(n7418), .A2(n7022), .ZN(n7023) );
  OR2_X1 U8772 ( .A1(n7023), .A2(n7403), .ZN(n7024) );
  NAND2_X1 U8773 ( .A1(n7023), .A2(n7403), .ZN(n7025) );
  NAND3_X1 U8774 ( .A1(n7398), .A2(n4448), .A3(n7025), .ZN(n7026) );
  AOI21_X1 U8775 ( .B1(n7450), .B2(n7026), .A(n8486), .ZN(n7029) );
  NAND2_X1 U8776 ( .A1(n10045), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n7027) );
  NAND2_X1 U8777 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7958) );
  OAI211_X1 U8778 ( .C1(n10023), .C2(n7454), .A(n7027), .B(n7958), .ZN(n7028)
         );
  NOR3_X1 U8779 ( .A1(n7030), .A2(n7029), .A3(n7028), .ZN(n7031) );
  OAI21_X1 U8780 ( .B1(n7032), .B2(n8542), .A(n7031), .ZN(P2_U3190) );
  AOI21_X1 U8781 ( .B1(n7035), .B2(n7034), .A(n7033), .ZN(n7041) );
  NAND2_X1 U8782 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9804) );
  INV_X1 U8783 ( .A(n9804), .ZN(n7036) );
  AOI21_X1 U8784 ( .B1(n8999), .B2(n9931), .A(n7036), .ZN(n7038) );
  NAND2_X1 U8785 ( .A1(n9004), .A2(n7112), .ZN(n7037) );
  OAI211_X1 U8786 ( .C1(n7107), .C2(n9001), .A(n7038), .B(n7037), .ZN(n7039)
         );
  AOI21_X1 U8787 ( .B1(n7113), .B2(n8972), .A(n7039), .ZN(n7040) );
  OAI21_X1 U8788 ( .B1(n7041), .B2(n8974), .A(n7040), .ZN(P1_U3239) );
  XNOR2_X1 U8789 ( .A(n7043), .B(n7042), .ZN(n7577) );
  XNOR2_X1 U8790 ( .A(n7044), .B(n7045), .ZN(n7047) );
  AOI222_X1 U8791 ( .A1(n8731), .A2(n7047), .B1(n5101), .B2(n8728), .C1(n7046), 
        .C2(n8726), .ZN(n7572) );
  OAI21_X1 U8792 ( .B1(n8118), .B2(n7577), .A(n7572), .ZN(n7907) );
  INV_X1 U8793 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n7048) );
  OAI22_X1 U8794 ( .A1(n8841), .A2(n7905), .B1(n7048), .B2(n10088), .ZN(n7049)
         );
  AOI21_X1 U8795 ( .B1(n10088), .B2(n7907), .A(n7049), .ZN(n7050) );
  INV_X1 U8796 ( .A(n7050), .ZN(P2_U3393) );
  OAI21_X1 U8797 ( .B1(n7052), .B2(n9023), .A(n7051), .ZN(n9958) );
  AOI211_X1 U8798 ( .C1(n8896), .C2(n7084), .A(n9590), .B(n7067), .ZN(n9950)
         );
  XOR2_X1 U8799 ( .A(n7053), .B(n9023), .Z(n7054) );
  AOI222_X1 U8800 ( .A1(n9284), .A2(n9932), .B1(n9282), .B2(n7513), .C1(n9906), 
        .C2(n7054), .ZN(n9961) );
  INV_X1 U8801 ( .A(n9961), .ZN(n7055) );
  AOI211_X1 U8802 ( .C1(n10007), .C2(n9958), .A(n9950), .B(n7055), .ZN(n7061)
         );
  OAI22_X1 U8803 ( .A1(n9645), .A2(n9956), .B1(n10021), .B2(n5682), .ZN(n7056)
         );
  INV_X1 U8804 ( .A(n7056), .ZN(n7057) );
  OAI21_X1 U8805 ( .B1(n7061), .B2(n10019), .A(n7057), .ZN(P1_U3525) );
  INV_X1 U8806 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n7058) );
  OAI22_X1 U8807 ( .A1(n9709), .A2(n9956), .B1(n10010), .B2(n7058), .ZN(n7059)
         );
  INV_X1 U8808 ( .A(n7059), .ZN(n7060) );
  OAI21_X1 U8809 ( .B1(n7061), .B2(n10009), .A(n7060), .ZN(P1_U3462) );
  XNOR2_X1 U8810 ( .A(n7062), .B(n9020), .ZN(n7063) );
  OAI222_X1 U8811 ( .A1(n7914), .A2(n7107), .B1(n7913), .B2(n7077), .C1(n9934), 
        .C2(n7063), .ZN(n9971) );
  INV_X1 U8812 ( .A(n9971), .ZN(n7074) );
  OAI21_X1 U8813 ( .B1(n7065), .B2(n9020), .A(n7064), .ZN(n9973) );
  OAI211_X1 U8814 ( .C1(n9970), .C2(n7067), .A(n7066), .B(n9942), .ZN(n9969)
         );
  AOI22_X1 U8815 ( .A1(n9593), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7068), .B2(
        n9952), .ZN(n7071) );
  NAND2_X1 U8816 ( .A1(n9939), .A2(n7069), .ZN(n7070) );
  OAI211_X1 U8817 ( .C1(n9969), .C2(n9405), .A(n7071), .B(n7070), .ZN(n7072)
         );
  AOI21_X1 U8818 ( .B1(n9973), .B2(n9959), .A(n7072), .ZN(n7073) );
  OAI21_X1 U8819 ( .B1(n7074), .B2(n9593), .A(n7073), .ZN(P1_U3289) );
  NOR2_X1 U8820 ( .A1(n7075), .A2(n7081), .ZN(n9027) );
  AOI211_X1 U8821 ( .C1(n7081), .C2(n7075), .A(n9934), .B(n9027), .ZN(n7079)
         );
  OAI22_X1 U8822 ( .A1(n7077), .A2(n7914), .B1(n7076), .B2(n7913), .ZN(n7078)
         );
  OR2_X1 U8823 ( .A1(n7079), .A2(n7078), .ZN(n9966) );
  INV_X1 U8824 ( .A(n9966), .ZN(n7093) );
  OAI21_X1 U8825 ( .B1(n7082), .B2(n7081), .A(n7080), .ZN(n9968) );
  INV_X1 U8826 ( .A(n7083), .ZN(n7085) );
  OAI211_X1 U8827 ( .C1(n7085), .C2(n9965), .A(n9942), .B(n7084), .ZN(n9964)
         );
  OAI22_X1 U8828 ( .A1(n9598), .A2(n7087), .B1(n7086), .B2(n9515), .ZN(n7088)
         );
  AOI21_X1 U8829 ( .B1(n9939), .B2(n7089), .A(n7088), .ZN(n7090) );
  OAI21_X1 U8830 ( .B1(n9405), .B2(n9964), .A(n7090), .ZN(n7091) );
  AOI21_X1 U8831 ( .B1(n9959), .B2(n9968), .A(n7091), .ZN(n7092) );
  OAI21_X1 U8832 ( .B1(n7093), .B2(n9593), .A(n7092), .ZN(P1_U3291) );
  AOI211_X1 U8833 ( .C1(n10007), .C2(n7096), .A(n7095), .B(n7094), .ZN(n7102)
         );
  OAI22_X1 U8834 ( .A1(n9645), .A2(n7099), .B1(n10021), .B2(n6760), .ZN(n7097)
         );
  INV_X1 U8835 ( .A(n7097), .ZN(n7098) );
  OAI21_X1 U8836 ( .B1(n7102), .B2(n10019), .A(n7098), .ZN(P1_U3527) );
  OAI22_X1 U8837 ( .A1(n9709), .A2(n7099), .B1(n10010), .B2(n5720), .ZN(n7100)
         );
  INV_X1 U8838 ( .A(n7100), .ZN(n7101) );
  OAI21_X1 U8839 ( .B1(n7102), .B2(n10009), .A(n7101), .ZN(P1_U3468) );
  INV_X1 U8840 ( .A(n7103), .ZN(n7120) );
  INV_X1 U8841 ( .A(n9883), .ZN(n9370) );
  INV_X1 U8842 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7104) );
  OAI222_X1 U8843 ( .A1(n9732), .A2(n7120), .B1(n9370), .B2(P1_U3086), .C1(
        n7104), .C2(n9729), .ZN(P1_U3338) );
  INV_X1 U8844 ( .A(n7105), .ZN(n7474) );
  XNOR2_X1 U8845 ( .A(n7474), .B(n7109), .ZN(n7106) );
  OAI222_X1 U8846 ( .A1(n7914), .A2(n7681), .B1(n7913), .B2(n7107), .C1(n9934), 
        .C2(n7106), .ZN(n9976) );
  INV_X1 U8847 ( .A(n9976), .ZN(n7118) );
  OAI21_X1 U8848 ( .B1(n7110), .B2(n7109), .A(n7108), .ZN(n9978) );
  OAI211_X1 U8849 ( .C1(n7111), .C2(n9975), .A(n9942), .B(n7479), .ZN(n9974)
         );
  AOI22_X1 U8850 ( .A1(n9593), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7112), .B2(
        n9952), .ZN(n7115) );
  NAND2_X1 U8851 ( .A1(n9939), .A2(n7113), .ZN(n7114) );
  OAI211_X1 U8852 ( .C1(n9974), .C2(n9405), .A(n7115), .B(n7114), .ZN(n7116)
         );
  AOI21_X1 U8853 ( .B1(n9978), .B2(n9959), .A(n7116), .ZN(n7117) );
  OAI21_X1 U8854 ( .B1(n7118), .B2(n9593), .A(n7117), .ZN(P1_U3287) );
  INV_X1 U8855 ( .A(n8505), .ZN(n8476) );
  INV_X1 U8856 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7119) );
  OAI222_X1 U8857 ( .A1(P2_U3151), .A2(n8476), .B1(n6665), .B2(n7120), .C1(
        n7119), .C2(n8880), .ZN(P2_U3278) );
  INV_X1 U8858 ( .A(n9372), .ZN(n9898) );
  INV_X1 U8859 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7121) );
  OAI222_X1 U8860 ( .A1(n9732), .A2(n7122), .B1(n9898), .B2(P1_U3086), .C1(
        n7121), .C2(n9729), .ZN(P1_U3337) );
  INV_X1 U8861 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7123) );
  INV_X1 U8862 ( .A(n8532), .ZN(n8499) );
  OAI222_X1 U8863 ( .A1(n8880), .A2(n7123), .B1(n6665), .B2(n7122), .C1(
        P2_U3151), .C2(n8499), .ZN(P2_U3277) );
  AOI21_X1 U8864 ( .B1(n7131), .B2(n7125), .A(n7124), .ZN(n7126) );
  AOI21_X1 U8865 ( .B1(n7127), .B2(n8542), .A(n7126), .ZN(n7128) );
  AOI21_X1 U8866 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .A(n7128), .ZN(
        n7130) );
  NAND2_X1 U8867 ( .A1(n10045), .A2(P2_ADDR_REG_0__SCAN_IN), .ZN(n7129) );
  OAI211_X1 U8868 ( .C1(n10023), .C2(n7131), .A(n7130), .B(n7129), .ZN(
        P2_U3182) );
  NOR2_X1 U8869 ( .A1(n7132), .A2(n4446), .ZN(n7133) );
  XNOR2_X1 U8870 ( .A(n7134), .B(n7133), .ZN(n7140) );
  NOR2_X1 U8871 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7135), .ZN(n9337) );
  AOI21_X1 U8872 ( .B1(n8999), .B2(n9922), .A(n9337), .ZN(n7137) );
  NAND2_X1 U8873 ( .A1(n9004), .A2(n7480), .ZN(n7136) );
  OAI211_X1 U8874 ( .C1(n7478), .C2(n9001), .A(n7137), .B(n7136), .ZN(n7138)
         );
  AOI21_X1 U8875 ( .B1(n7598), .B2(n8972), .A(n7138), .ZN(n7139) );
  OAI21_X1 U8876 ( .B1(n7140), .B2(n8974), .A(n7139), .ZN(P1_U3213) );
  INV_X1 U8877 ( .A(n7141), .ZN(n7150) );
  NAND2_X1 U8878 ( .A1(n7142), .A2(n9598), .ZN(n7149) );
  NOR2_X1 U8879 ( .A1(n9955), .A2(n6060), .ZN(n7146) );
  OAI22_X1 U8880 ( .A1(n9598), .A2(n7144), .B1(n7143), .B2(n9515), .ZN(n7145)
         );
  AOI211_X1 U8881 ( .C1(n7147), .C2(n9949), .A(n7146), .B(n7145), .ZN(n7148)
         );
  OAI211_X1 U8882 ( .C1(n9601), .C2(n7150), .A(n7149), .B(n7148), .ZN(P1_U3292) );
  INV_X1 U8883 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10098) );
  INV_X1 U8884 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9889) );
  INV_X1 U8885 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8479) );
  AOI22_X1 U8886 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .B1(n9889), .B2(n8479), .ZN(n10103) );
  NOR2_X1 U8887 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7151) );
  AOI21_X1 U8888 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7151), .ZN(n10106) );
  NOR2_X1 U8889 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7152) );
  AOI21_X1 U8890 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7152), .ZN(n10109) );
  NOR2_X1 U8891 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7153) );
  AOI21_X1 U8892 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7153), .ZN(n10112) );
  NOR2_X1 U8893 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7154) );
  AOI21_X1 U8894 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7154), .ZN(n10115) );
  NOR2_X1 U8895 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7155) );
  AOI21_X1 U8896 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7155), .ZN(n10118) );
  NOR2_X1 U8897 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7156) );
  AOI21_X1 U8898 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7156), .ZN(n10121) );
  NOR2_X1 U8899 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7157) );
  AOI21_X1 U8900 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7157), .ZN(n10124) );
  NOR2_X1 U8901 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7158) );
  AOI21_X1 U8902 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7158), .ZN(n10130) );
  NOR2_X1 U8903 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7159) );
  AOI21_X1 U8904 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7159), .ZN(n10133) );
  NOR2_X1 U8905 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7160) );
  AOI21_X1 U8906 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7160), .ZN(n10136) );
  NOR2_X1 U8907 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7161) );
  AOI21_X1 U8908 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n7161), .ZN(n10139) );
  NOR2_X1 U8909 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(P2_ADDR_REG_5__SCAN_IN), 
        .ZN(n7162) );
  AOI21_X1 U8910 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n7162), .ZN(n10142) );
  AND2_X1 U8911 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7163) );
  NOR2_X1 U8912 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7163), .ZN(n10093) );
  INV_X1 U8913 ( .A(n10093), .ZN(n10094) );
  INV_X1 U8914 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10096) );
  NAND3_X1 U8915 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10095) );
  NAND2_X1 U8916 ( .A1(n10096), .A2(n10095), .ZN(n10092) );
  NAND2_X1 U8917 ( .A1(n10094), .A2(n10092), .ZN(n10127) );
  NAND2_X1 U8918 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7164) );
  OAI21_X1 U8919 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7164), .ZN(n10126) );
  NOR2_X1 U8920 ( .A1(n10127), .A2(n10126), .ZN(n10125) );
  AOI21_X1 U8921 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10125), .ZN(n10145) );
  NAND2_X1 U8922 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7165) );
  OAI21_X1 U8923 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n7165), .ZN(n10144) );
  NOR2_X1 U8924 ( .A1(n10145), .A2(n10144), .ZN(n10143) );
  AOI21_X1 U8925 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10143), .ZN(n10148) );
  NOR2_X1 U8926 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7166) );
  AOI21_X1 U8927 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7166), .ZN(n10147) );
  NAND2_X1 U8928 ( .A1(n10148), .A2(n10147), .ZN(n10146) );
  OAI21_X1 U8929 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10146), .ZN(n10141) );
  NAND2_X1 U8930 ( .A1(n10142), .A2(n10141), .ZN(n10140) );
  OAI21_X1 U8931 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n10140), .ZN(n10138) );
  NAND2_X1 U8932 ( .A1(n10139), .A2(n10138), .ZN(n10137) );
  OAI21_X1 U8933 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10137), .ZN(n10135) );
  NAND2_X1 U8934 ( .A1(n10136), .A2(n10135), .ZN(n10134) );
  OAI21_X1 U8935 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10134), .ZN(n10132) );
  NAND2_X1 U8936 ( .A1(n10133), .A2(n10132), .ZN(n10131) );
  OAI21_X1 U8937 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10131), .ZN(n10129) );
  NAND2_X1 U8938 ( .A1(n10130), .A2(n10129), .ZN(n10128) );
  OAI21_X1 U8939 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10128), .ZN(n10123) );
  NAND2_X1 U8940 ( .A1(n10124), .A2(n10123), .ZN(n10122) );
  OAI21_X1 U8941 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10122), .ZN(n10120) );
  NAND2_X1 U8942 ( .A1(n10121), .A2(n10120), .ZN(n10119) );
  OAI21_X1 U8943 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10119), .ZN(n10117) );
  NAND2_X1 U8944 ( .A1(n10118), .A2(n10117), .ZN(n10116) );
  OAI21_X1 U8945 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10116), .ZN(n10114) );
  NAND2_X1 U8946 ( .A1(n10115), .A2(n10114), .ZN(n10113) );
  OAI21_X1 U8947 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10113), .ZN(n10111) );
  NAND2_X1 U8948 ( .A1(n10112), .A2(n10111), .ZN(n10110) );
  OAI21_X1 U8949 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10110), .ZN(n10108) );
  NAND2_X1 U8950 ( .A1(n10109), .A2(n10108), .ZN(n10107) );
  OAI21_X1 U8951 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10107), .ZN(n10105) );
  NAND2_X1 U8952 ( .A1(n10106), .A2(n10105), .ZN(n10104) );
  OAI21_X1 U8953 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10104), .ZN(n10102) );
  NAND2_X1 U8954 ( .A1(n10103), .A2(n10102), .ZN(n10101) );
  OAI21_X1 U8955 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10101), .ZN(n10099) );
  NAND2_X1 U8956 ( .A1(n10098), .A2(n10099), .ZN(n7167) );
  NOR2_X1 U8957 ( .A1(n10098), .A2(n10099), .ZN(n10097) );
  AOI21_X1 U8958 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n7167), .A(n10097), .ZN(
        n7357) );
  INV_X1 U8959 ( .A(P2_WR_REG_SCAN_IN), .ZN(n9786) );
  AOI22_X1 U8960 ( .A1(n9786), .A2(keyinput_g0), .B1(n5030), .B2(keyinput_g53), 
        .ZN(n7168) );
  OAI221_X1 U8961 ( .B1(n9786), .B2(keyinput_g0), .C1(n5030), .C2(keyinput_g53), .A(n7168), .ZN(n7175) );
  INV_X1 U8962 ( .A(SI_12_), .ZN(n7332) );
  AOI22_X1 U8963 ( .A1(n7337), .A2(keyinput_g6), .B1(keyinput_g20), .B2(n7332), 
        .ZN(n7169) );
  OAI221_X1 U8964 ( .B1(n7337), .B2(keyinput_g6), .C1(n7332), .C2(keyinput_g20), .A(n7169), .ZN(n7174) );
  INV_X1 U8965 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7661) );
  AOI22_X1 U8966 ( .A1(n5038), .A2(keyinput_g45), .B1(keyinput_g39), .B2(n7661), .ZN(n7170) );
  OAI221_X1 U8967 ( .B1(n5038), .B2(keyinput_g45), .C1(n7661), .C2(
        keyinput_g39), .A(n7170), .ZN(n7173) );
  AOI22_X1 U8968 ( .A1(n7320), .A2(keyinput_g9), .B1(n7293), .B2(keyinput_g7), 
        .ZN(n7171) );
  OAI221_X1 U8969 ( .B1(n7320), .B2(keyinput_g9), .C1(n7293), .C2(keyinput_g7), 
        .A(n7171), .ZN(n7172) );
  NOR4_X1 U8970 ( .A1(n7175), .A2(n7174), .A3(n7173), .A4(n7172), .ZN(n7353)
         );
  AOI22_X1 U8971 ( .A1(n7177), .A2(keyinput_g25), .B1(n5028), .B2(keyinput_g35), .ZN(n7176) );
  OAI221_X1 U8972 ( .B1(n7177), .B2(keyinput_g25), .C1(n5028), .C2(
        keyinput_g35), .A(n7176), .ZN(n7184) );
  AOI22_X1 U8973 ( .A1(n7260), .A2(keyinput_g13), .B1(keyinput_g21), .B2(n7321), .ZN(n7178) );
  OAI221_X1 U8974 ( .B1(n7260), .B2(keyinput_g13), .C1(n7321), .C2(
        keyinput_g21), .A(n7178), .ZN(n7183) );
  AOI22_X1 U8975 ( .A1(n7181), .A2(keyinput_g63), .B1(keyinput_g24), .B2(n7180), .ZN(n7179) );
  OAI221_X1 U8976 ( .B1(n7181), .B2(keyinput_g63), .C1(n7180), .C2(
        keyinput_g24), .A(n7179), .ZN(n7182) );
  NOR3_X1 U8977 ( .A1(n7184), .A2(n7183), .A3(n7182), .ZN(n7211) );
  AOI22_X1 U8978 ( .A1(n7272), .A2(keyinput_g18), .B1(n5025), .B2(keyinput_g52), .ZN(n7185) );
  OAI221_X1 U8979 ( .B1(n7272), .B2(keyinput_g18), .C1(n5025), .C2(
        keyinput_g52), .A(n7185), .ZN(n7193) );
  INV_X1 U8980 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8080) );
  AOI22_X1 U8981 ( .A1(n7187), .A2(keyinput_g26), .B1(n8080), .B2(keyinput_g56), .ZN(n7186) );
  OAI221_X1 U8982 ( .B1(n7187), .B2(keyinput_g26), .C1(n8080), .C2(
        keyinput_g56), .A(n7186), .ZN(n7192) );
  AOI22_X1 U8983 ( .A1(n7190), .A2(keyinput_g27), .B1(n7189), .B2(keyinput_g10), .ZN(n7188) );
  OAI221_X1 U8984 ( .B1(n7190), .B2(keyinput_g27), .C1(n7189), .C2(
        keyinput_g10), .A(n7188), .ZN(n7191) );
  NOR3_X1 U8985 ( .A1(n7193), .A2(n7192), .A3(n7191), .ZN(n7210) );
  INV_X1 U8986 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7290) );
  AOI22_X1 U8987 ( .A1(n7290), .A2(keyinput_g37), .B1(keyinput_g16), .B2(n7329), .ZN(n7194) );
  OAI221_X1 U8988 ( .B1(n7290), .B2(keyinput_g37), .C1(n7329), .C2(
        keyinput_g16), .A(n7194), .ZN(n7200) );
  XNOR2_X1 U8989 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_g48), .ZN(n7198)
         );
  XNOR2_X1 U8990 ( .A(SI_2_), .B(keyinput_g30), .ZN(n7197) );
  XNOR2_X1 U8991 ( .A(SI_3_), .B(keyinput_g29), .ZN(n7196) );
  XNOR2_X1 U8992 ( .A(SI_24_), .B(keyinput_g8), .ZN(n7195) );
  NAND4_X1 U8993 ( .A1(n7198), .A2(n7197), .A3(n7196), .A4(n7195), .ZN(n7199)
         );
  NOR2_X1 U8994 ( .A1(n7200), .A2(n7199), .ZN(n7209) );
  INV_X1 U8995 ( .A(SI_13_), .ZN(n7270) );
  AOI22_X1 U8996 ( .A1(n7270), .A2(keyinput_g19), .B1(n7305), .B2(keyinput_g3), 
        .ZN(n7201) );
  OAI221_X1 U8997 ( .B1(n7270), .B2(keyinput_g19), .C1(n7305), .C2(keyinput_g3), .A(n7201), .ZN(n7207) );
  XNOR2_X1 U8998 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput_g61), .ZN(n7205) );
  XNOR2_X1 U8999 ( .A(SI_1_), .B(keyinput_g31), .ZN(n7204) );
  XNOR2_X1 U9000 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput_g38), .ZN(n7203)
         );
  XNOR2_X1 U9001 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_g54), .ZN(n7202) );
  NAND4_X1 U9002 ( .A1(n7205), .A2(n7204), .A3(n7203), .A4(n7202), .ZN(n7206)
         );
  NOR2_X1 U9003 ( .A1(n7207), .A2(n7206), .ZN(n7208) );
  NAND4_X1 U9004 ( .A1(n7211), .A2(n7210), .A3(n7209), .A4(n7208), .ZN(n7248)
         );
  AOI22_X1 U9005 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(keyinput_g58), .B1(
        P2_REG3_REG_19__SCAN_IN), .B2(keyinput_g41), .ZN(n7212) );
  OAI221_X1 U9006 ( .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput_g58), .C1(
        P2_REG3_REG_19__SCAN_IN), .C2(keyinput_g41), .A(n7212), .ZN(n7219) );
  AOI22_X1 U9007 ( .A1(SI_17_), .A2(keyinput_g15), .B1(P2_REG3_REG_5__SCAN_IN), 
        .B2(keyinput_g49), .ZN(n7213) );
  OAI221_X1 U9008 ( .B1(SI_17_), .B2(keyinput_g15), .C1(P2_REG3_REG_5__SCAN_IN), .C2(keyinput_g49), .A(n7213), .ZN(n7218) );
  AOI22_X1 U9009 ( .A1(SI_31_), .A2(keyinput_g1), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(keyinput_g40), .ZN(n7214) );
  OAI221_X1 U9010 ( .B1(SI_31_), .B2(keyinput_g1), .C1(P2_REG3_REG_3__SCAN_IN), 
        .C2(keyinput_g40), .A(n7214), .ZN(n7217) );
  AOI22_X1 U9011 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_g44), .B1(
        P2_REG3_REG_26__SCAN_IN), .B2(keyinput_g62), .ZN(n7215) );
  OAI221_X1 U9012 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_g44), .C1(
        P2_REG3_REG_26__SCAN_IN), .C2(keyinput_g62), .A(n7215), .ZN(n7216) );
  NOR4_X1 U9013 ( .A1(n7219), .A2(n7218), .A3(n7217), .A4(n7216), .ZN(n7246)
         );
  INV_X1 U9014 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n7310) );
  XNOR2_X1 U9015 ( .A(n7310), .B(keyinput_g57), .ZN(n7226) );
  AOI22_X1 U9016 ( .A1(SI_20_), .A2(keyinput_g12), .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_g51), .ZN(n7220) );
  OAI221_X1 U9017 ( .B1(SI_20_), .B2(keyinput_g12), .C1(
        P2_REG3_REG_24__SCAN_IN), .C2(keyinput_g51), .A(n7220), .ZN(n7225) );
  AOI22_X1 U9018 ( .A1(SI_15_), .A2(keyinput_g17), .B1(SI_28_), .B2(
        keyinput_g4), .ZN(n7221) );
  OAI221_X1 U9019 ( .B1(SI_15_), .B2(keyinput_g17), .C1(SI_28_), .C2(
        keyinput_g4), .A(n7221), .ZN(n7224) );
  AOI22_X1 U9020 ( .A1(P2_RD_REG_SCAN_IN), .A2(keyinput_g33), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(keyinput_g50), .ZN(n7222) );
  OAI221_X1 U9021 ( .B1(P2_RD_REG_SCAN_IN), .B2(keyinput_g33), .C1(
        P2_REG3_REG_17__SCAN_IN), .C2(keyinput_g50), .A(n7222), .ZN(n7223) );
  NOR4_X1 U9022 ( .A1(n7226), .A2(n7225), .A3(n7224), .A4(n7223), .ZN(n7245)
         );
  AOI22_X1 U9023 ( .A1(SI_0_), .A2(keyinput_g32), .B1(P2_REG3_REG_12__SCAN_IN), 
        .B2(keyinput_g46), .ZN(n7227) );
  OAI221_X1 U9024 ( .B1(SI_0_), .B2(keyinput_g32), .C1(P2_REG3_REG_12__SCAN_IN), .C2(keyinput_g46), .A(n7227), .ZN(n7234) );
  AOI22_X1 U9025 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput_g47), .B1(
        P2_REG3_REG_27__SCAN_IN), .B2(keyinput_g36), .ZN(n7228) );
  OAI221_X1 U9026 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_g47), .C1(
        P2_REG3_REG_27__SCAN_IN), .C2(keyinput_g36), .A(n7228), .ZN(n7233) );
  AOI22_X1 U9027 ( .A1(SI_21_), .A2(keyinput_g11), .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .ZN(n7229) );
  OAI221_X1 U9028 ( .B1(SI_21_), .B2(keyinput_g11), .C1(
        P2_REG3_REG_18__SCAN_IN), .C2(keyinput_g60), .A(n7229), .ZN(n7232) );
  AOI22_X1 U9029 ( .A1(SI_30_), .A2(keyinput_g2), .B1(SI_10_), .B2(
        keyinput_g22), .ZN(n7230) );
  OAI221_X1 U9030 ( .B1(SI_30_), .B2(keyinput_g2), .C1(SI_10_), .C2(
        keyinput_g22), .A(n7230), .ZN(n7231) );
  NOR4_X1 U9031 ( .A1(n7234), .A2(n7233), .A3(n7232), .A4(n7231), .ZN(n7244)
         );
  AOI22_X1 U9032 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_g59), .B1(
        P2_REG3_REG_8__SCAN_IN), .B2(keyinput_g43), .ZN(n7235) );
  OAI221_X1 U9033 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_g59), .C1(
        P2_REG3_REG_8__SCAN_IN), .C2(keyinput_g43), .A(n7235), .ZN(n7242) );
  AOI22_X1 U9034 ( .A1(SI_27_), .A2(keyinput_g5), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(keyinput_g42), .ZN(n7236) );
  OAI221_X1 U9035 ( .B1(SI_27_), .B2(keyinput_g5), .C1(P2_REG3_REG_28__SCAN_IN), .C2(keyinput_g42), .A(n7236), .ZN(n7241) );
  AOI22_X1 U9036 ( .A1(P2_STATE_REG_SCAN_IN), .A2(keyinput_g34), .B1(
        P2_REG3_REG_20__SCAN_IN), .B2(keyinput_g55), .ZN(n7237) );
  OAI221_X1 U9037 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput_g34), .C1(
        P2_REG3_REG_20__SCAN_IN), .C2(keyinput_g55), .A(n7237), .ZN(n7240) );
  AOI22_X1 U9038 ( .A1(SI_9_), .A2(keyinput_g23), .B1(SI_18_), .B2(
        keyinput_g14), .ZN(n7238) );
  OAI221_X1 U9039 ( .B1(SI_9_), .B2(keyinput_g23), .C1(SI_18_), .C2(
        keyinput_g14), .A(n7238), .ZN(n7239) );
  NOR4_X1 U9040 ( .A1(n7242), .A2(n7241), .A3(n7240), .A4(n7239), .ZN(n7243)
         );
  NAND4_X1 U9041 ( .A1(n7246), .A2(n7245), .A3(n7244), .A4(n7243), .ZN(n7247)
         );
  NOR2_X1 U9042 ( .A1(n7248), .A2(n7247), .ZN(n7352) );
  XNOR2_X1 U9043 ( .A(n7249), .B(keyinput_g28), .ZN(n7351) );
  AOI22_X1 U9044 ( .A1(SI_20_), .A2(keyinput_f12), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(keyinput_f40), .ZN(n7250) );
  OAI221_X1 U9045 ( .B1(SI_20_), .B2(keyinput_f12), .C1(P2_REG3_REG_3__SCAN_IN), .C2(keyinput_f40), .A(n7250), .ZN(n7257) );
  AOI22_X1 U9046 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(keyinput_f58), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(keyinput_f63), .ZN(n7251) );
  OAI221_X1 U9047 ( .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput_f58), .C1(
        P2_REG3_REG_15__SCAN_IN), .C2(keyinput_f63), .A(n7251), .ZN(n7256) );
  AOI22_X1 U9048 ( .A1(SI_2_), .A2(keyinput_f30), .B1(SI_3_), .B2(keyinput_f29), .ZN(n7252) );
  OAI221_X1 U9049 ( .B1(SI_2_), .B2(keyinput_f30), .C1(SI_3_), .C2(
        keyinput_f29), .A(n7252), .ZN(n7255) );
  AOI22_X1 U9050 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(keyinput_f52), .B1(
        P2_REG3_REG_28__SCAN_IN), .B2(keyinput_f42), .ZN(n7253) );
  OAI221_X1 U9051 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput_f52), .C1(
        P2_REG3_REG_28__SCAN_IN), .C2(keyinput_f42), .A(n7253), .ZN(n7254) );
  NOR4_X1 U9052 ( .A1(n7257), .A2(n7256), .A3(n7255), .A4(n7254), .ZN(n7288)
         );
  INV_X1 U9053 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7258) );
  XOR2_X1 U9054 ( .A(n7258), .B(keyinput_f61), .Z(n7266) );
  AOI22_X1 U9055 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_f60), .B1(n7260), 
        .B2(keyinput_f13), .ZN(n7259) );
  OAI221_X1 U9056 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_f60), .C1(n7260), .C2(keyinput_f13), .A(n7259), .ZN(n7265) );
  AOI22_X1 U9057 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput_f46), .B1(
        P2_REG3_REG_24__SCAN_IN), .B2(keyinput_f51), .ZN(n7261) );
  OAI221_X1 U9058 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_f46), .C1(
        P2_REG3_REG_24__SCAN_IN), .C2(keyinput_f51), .A(n7261), .ZN(n7264) );
  AOI22_X1 U9059 ( .A1(SI_5_), .A2(keyinput_f27), .B1(SI_21_), .B2(
        keyinput_f11), .ZN(n7262) );
  OAI221_X1 U9060 ( .B1(SI_5_), .B2(keyinput_f27), .C1(SI_21_), .C2(
        keyinput_f11), .A(n7262), .ZN(n7263) );
  NOR4_X1 U9061 ( .A1(n7266), .A2(n7265), .A3(n7264), .A4(n7263), .ZN(n7287)
         );
  AOI22_X1 U9062 ( .A1(SI_6_), .A2(keyinput_f26), .B1(P2_REG3_REG_17__SCAN_IN), 
        .B2(keyinput_f50), .ZN(n7267) );
  OAI221_X1 U9063 ( .B1(SI_6_), .B2(keyinput_f26), .C1(P2_REG3_REG_17__SCAN_IN), .C2(keyinput_f50), .A(n7267), .ZN(n7276) );
  AOI22_X1 U9064 ( .A1(keyinput_f0), .A2(P2_WR_REG_SCAN_IN), .B1(
        P2_REG3_REG_27__SCAN_IN), .B2(keyinput_f36), .ZN(n7268) );
  OAI221_X1 U9065 ( .B1(keyinput_f0), .B2(P2_WR_REG_SCAN_IN), .C1(
        P2_REG3_REG_27__SCAN_IN), .C2(keyinput_f36), .A(n7268), .ZN(n7275) );
  AOI22_X1 U9066 ( .A1(n7270), .A2(keyinput_f19), .B1(n5030), .B2(keyinput_f53), .ZN(n7269) );
  OAI221_X1 U9067 ( .B1(n7270), .B2(keyinput_f19), .C1(n5030), .C2(
        keyinput_f53), .A(n7269), .ZN(n7274) );
  AOI22_X1 U9068 ( .A1(P2_STATE_REG_SCAN_IN), .A2(keyinput_f34), .B1(n7272), 
        .B2(keyinput_f18), .ZN(n7271) );
  OAI221_X1 U9069 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput_f34), .C1(n7272), 
        .C2(keyinput_f18), .A(n7271), .ZN(n7273) );
  NOR4_X1 U9070 ( .A1(n7276), .A2(n7275), .A3(n7274), .A4(n7273), .ZN(n7286)
         );
  AOI22_X1 U9071 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_f54), .B1(SI_22_), 
        .B2(keyinput_f10), .ZN(n7277) );
  OAI221_X1 U9072 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_f54), .C1(SI_22_), .C2(keyinput_f10), .A(n7277), .ZN(n7284) );
  AOI22_X1 U9073 ( .A1(SI_7_), .A2(keyinput_f25), .B1(SI_9_), .B2(keyinput_f23), .ZN(n7278) );
  OAI221_X1 U9074 ( .B1(SI_7_), .B2(keyinput_f25), .C1(SI_9_), .C2(
        keyinput_f23), .A(n7278), .ZN(n7283) );
  AOI22_X1 U9075 ( .A1(SI_18_), .A2(keyinput_f14), .B1(P2_REG3_REG_8__SCAN_IN), 
        .B2(keyinput_f43), .ZN(n7279) );
  OAI221_X1 U9076 ( .B1(SI_18_), .B2(keyinput_f14), .C1(P2_REG3_REG_8__SCAN_IN), .C2(keyinput_f43), .A(n7279), .ZN(n7282) );
  AOI22_X1 U9077 ( .A1(SI_10_), .A2(keyinput_f22), .B1(SI_15_), .B2(
        keyinput_f17), .ZN(n7280) );
  OAI221_X1 U9078 ( .B1(SI_10_), .B2(keyinput_f22), .C1(SI_15_), .C2(
        keyinput_f17), .A(n7280), .ZN(n7281) );
  NOR4_X1 U9079 ( .A1(n7284), .A2(n7283), .A3(n7282), .A4(n7281), .ZN(n7285)
         );
  NAND4_X1 U9080 ( .A1(n7288), .A2(n7287), .A3(n7286), .A4(n7285), .ZN(n7348)
         );
  AOI22_X1 U9081 ( .A1(n7290), .A2(keyinput_f37), .B1(keyinput_f33), .B2(n4717), .ZN(n7289) );
  OAI221_X1 U9082 ( .B1(n7290), .B2(keyinput_f37), .C1(n4717), .C2(
        keyinput_f33), .A(n7289), .ZN(n7301) );
  AOI22_X1 U9083 ( .A1(n7293), .A2(keyinput_f7), .B1(keyinput_f15), .B2(n7292), 
        .ZN(n7291) );
  OAI221_X1 U9084 ( .B1(n7293), .B2(keyinput_f7), .C1(n7292), .C2(keyinput_f15), .A(n7291), .ZN(n7300) );
  AOI22_X1 U9085 ( .A1(n7295), .A2(keyinput_f5), .B1(n8080), .B2(keyinput_f56), 
        .ZN(n7294) );
  OAI221_X1 U9086 ( .B1(n7295), .B2(keyinput_f5), .C1(n8080), .C2(keyinput_f56), .A(n7294), .ZN(n7299) );
  XNOR2_X1 U9087 ( .A(SI_1_), .B(keyinput_f31), .ZN(n7297) );
  XNOR2_X1 U9088 ( .A(SI_8_), .B(keyinput_f24), .ZN(n7296) );
  NAND2_X1 U9089 ( .A1(n7297), .A2(n7296), .ZN(n7298) );
  NOR4_X1 U9090 ( .A1(n7301), .A2(n7300), .A3(n7299), .A4(n7298), .ZN(n7346)
         );
  INV_X1 U9091 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n7303) );
  AOI22_X1 U9092 ( .A1(n7303), .A2(keyinput_f55), .B1(keyinput_f44), .B2(n6924), .ZN(n7302) );
  OAI221_X1 U9093 ( .B1(n7303), .B2(keyinput_f55), .C1(n6924), .C2(
        keyinput_f44), .A(n7302), .ZN(n7314) );
  INV_X1 U9094 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n7306) );
  AOI22_X1 U9095 ( .A1(n7306), .A2(keyinput_f38), .B1(keyinput_f3), .B2(n7305), 
        .ZN(n7304) );
  OAI221_X1 U9096 ( .B1(n7306), .B2(keyinput_f38), .C1(n7305), .C2(keyinput_f3), .A(n7304), .ZN(n7313) );
  AOI22_X1 U9097 ( .A1(n8252), .A2(keyinput_f47), .B1(keyinput_f8), .B2(n7308), 
        .ZN(n7307) );
  OAI221_X1 U9098 ( .B1(n8252), .B2(keyinput_f47), .C1(n7308), .C2(keyinput_f8), .A(n7307), .ZN(n7312) );
  AOI22_X1 U9099 ( .A1(n7310), .A2(keyinput_f57), .B1(keyinput_f45), .B2(n5038), .ZN(n7309) );
  OAI221_X1 U9100 ( .B1(n7310), .B2(keyinput_f57), .C1(n5038), .C2(
        keyinput_f45), .A(n7309), .ZN(n7311) );
  NOR4_X1 U9101 ( .A1(n7314), .A2(n7313), .A3(n7312), .A4(n7311), .ZN(n7345)
         );
  AOI22_X1 U9102 ( .A1(n7316), .A2(keyinput_f41), .B1(keyinput_f35), .B2(n5028), .ZN(n7315) );
  OAI221_X1 U9103 ( .B1(n7316), .B2(keyinput_f41), .C1(n5028), .C2(
        keyinput_f35), .A(n7315), .ZN(n7327) );
  INV_X1 U9104 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n7318) );
  AOI22_X1 U9105 ( .A1(n7318), .A2(keyinput_f62), .B1(keyinput_f49), .B2(n5026), .ZN(n7317) );
  OAI221_X1 U9106 ( .B1(n7318), .B2(keyinput_f62), .C1(n5026), .C2(
        keyinput_f49), .A(n7317), .ZN(n7326) );
  AOI22_X1 U9107 ( .A1(n7321), .A2(keyinput_f21), .B1(n7320), .B2(keyinput_f9), 
        .ZN(n7319) );
  OAI221_X1 U9108 ( .B1(n7321), .B2(keyinput_f21), .C1(n7320), .C2(keyinput_f9), .A(n7319), .ZN(n7325) );
  XNOR2_X1 U9109 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput_f39), .ZN(n7323)
         );
  XNOR2_X1 U9110 ( .A(SI_0_), .B(keyinput_f32), .ZN(n7322) );
  NAND2_X1 U9111 ( .A1(n7323), .A2(n7322), .ZN(n7324) );
  NOR4_X1 U9112 ( .A1(n7327), .A2(n7326), .A3(n7325), .A4(n7324), .ZN(n7344)
         );
  INV_X1 U9113 ( .A(SI_30_), .ZN(n7330) );
  AOI22_X1 U9114 ( .A1(n7330), .A2(keyinput_f2), .B1(n7329), .B2(keyinput_f16), 
        .ZN(n7328) );
  OAI221_X1 U9115 ( .B1(n7330), .B2(keyinput_f2), .C1(n7329), .C2(keyinput_f16), .A(n7328), .ZN(n7342) );
  INV_X1 U9116 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7333) );
  AOI22_X1 U9117 ( .A1(n7333), .A2(keyinput_f48), .B1(keyinput_f20), .B2(n7332), .ZN(n7331) );
  OAI221_X1 U9118 ( .B1(n7333), .B2(keyinput_f48), .C1(n7332), .C2(
        keyinput_f20), .A(n7331), .ZN(n7341) );
  AOI22_X1 U9119 ( .A1(n7335), .A2(keyinput_f4), .B1(keyinput_f59), .B2(n10063), .ZN(n7334) );
  OAI221_X1 U9120 ( .B1(n7335), .B2(keyinput_f4), .C1(n10063), .C2(
        keyinput_f59), .A(n7334), .ZN(n7340) );
  AOI22_X1 U9121 ( .A1(n7338), .A2(keyinput_f1), .B1(n7337), .B2(keyinput_f6), 
        .ZN(n7336) );
  OAI221_X1 U9122 ( .B1(n7338), .B2(keyinput_f1), .C1(n7337), .C2(keyinput_f6), 
        .A(n7336), .ZN(n7339) );
  NOR4_X1 U9123 ( .A1(n7342), .A2(n7341), .A3(n7340), .A4(n7339), .ZN(n7343)
         );
  NAND4_X1 U9124 ( .A1(n7346), .A2(n7345), .A3(n7344), .A4(n7343), .ZN(n7347)
         );
  OAI22_X1 U9125 ( .A1(n7348), .A2(n7347), .B1(keyinput_f28), .B2(SI_4_), .ZN(
        n7349) );
  AOI21_X1 U9126 ( .B1(keyinput_f28), .B2(SI_4_), .A(n7349), .ZN(n7350) );
  AOI211_X1 U9127 ( .C1(n7353), .C2(n7352), .A(n7351), .B(n7350), .ZN(n7355)
         );
  XNOR2_X1 U9128 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n7354) );
  XNOR2_X1 U9129 ( .A(n7355), .B(n7354), .ZN(n7356) );
  XNOR2_X1 U9130 ( .A(n7357), .B(n7356), .ZN(ADD_1068_U4) );
  XNOR2_X1 U9131 ( .A(n8173), .B(n7924), .ZN(n7531) );
  XOR2_X1 U9132 ( .A(n8370), .B(n7531), .Z(n7363) );
  INV_X1 U9133 ( .A(n7359), .ZN(n7361) );
  OAI21_X1 U9134 ( .B1(n7361), .B2(n5101), .A(n7360), .ZN(n7362) );
  AOI211_X1 U9135 ( .C1(n7363), .C2(n7362), .A(n8342), .B(n7532), .ZN(n7364)
         );
  INV_X1 U9136 ( .A(n7364), .ZN(n7368) );
  NAND2_X1 U9137 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n10059) );
  INV_X1 U9138 ( .A(n10059), .ZN(n7366) );
  OAI22_X1 U9139 ( .A1(n8324), .A2(n5100), .B1(n7614), .B2(n8347), .ZN(n7365)
         );
  AOI211_X1 U9140 ( .C1(n7924), .C2(n8339), .A(n7366), .B(n7365), .ZN(n7367)
         );
  OAI211_X1 U9141 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8348), .A(n7368), .B(
        n7367), .ZN(P2_U3158) );
  NAND2_X1 U9142 ( .A1(n6905), .A2(n7369), .ZN(n7370) );
  NAND4_X1 U9143 ( .A1(n7373), .A2(n7372), .A3(n7371), .A4(n7370), .ZN(n7374)
         );
  NOR2_X2 U9144 ( .A1(n7374), .A2(n10061), .ZN(n8735) );
  AOI22_X1 U9145 ( .A1(n8735), .A2(n7375), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n8719), .ZN(n7380) );
  INV_X1 U9146 ( .A(n7376), .ZN(n7377) );
  NAND2_X1 U9147 ( .A1(n8371), .A2(n8728), .ZN(n7729) );
  OAI21_X1 U9148 ( .B1(n7728), .B2(n7377), .A(n7729), .ZN(n7378) );
  NAND2_X1 U9149 ( .A1(n8715), .A2(n7378), .ZN(n7379) );
  OAI211_X1 U9150 ( .C1(n6954), .C2(n8715), .A(n7380), .B(n7379), .ZN(P2_U3233) );
  XNOR2_X1 U9151 ( .A(n7381), .B(n9018), .ZN(n9996) );
  INV_X1 U9152 ( .A(n9996), .ZN(n7395) );
  NAND2_X1 U9153 ( .A1(n7382), .A2(n9018), .ZN(n7383) );
  NAND2_X1 U9154 ( .A1(n7384), .A2(n7383), .ZN(n7385) );
  NAND2_X1 U9155 ( .A1(n7385), .A2(n9906), .ZN(n7387) );
  AOI22_X1 U9156 ( .A1(n9932), .A2(n9930), .B1(n9910), .B2(n7513), .ZN(n7386)
         );
  NAND2_X1 U9157 ( .A1(n7387), .A2(n7386), .ZN(n9995) );
  OAI211_X1 U9158 ( .C1(n4439), .C2(n9993), .A(n9942), .B(n7564), .ZN(n9992)
         );
  INV_X1 U9159 ( .A(n7803), .ZN(n7388) );
  OAI22_X1 U9160 ( .A1(n9598), .A2(n7389), .B1(n7388), .B2(n9515), .ZN(n7390)
         );
  AOI21_X1 U9161 ( .B1(n7391), .B2(n9939), .A(n7390), .ZN(n7392) );
  OAI21_X1 U9162 ( .B1(n9992), .B2(n9405), .A(n7392), .ZN(n7393) );
  AOI21_X1 U9163 ( .B1(n9995), .B2(n9598), .A(n7393), .ZN(n7394) );
  OAI21_X1 U9164 ( .B1(n7395), .B2(n9601), .A(n7394), .ZN(P1_U3283) );
  OAI21_X1 U9165 ( .B1(n7397), .B2(P2_REG1_REG_7__SCAN_IN), .A(n7396), .ZN(
        n7401) );
  INV_X1 U9166 ( .A(n10032), .ZN(n10043) );
  OAI21_X1 U9167 ( .B1(n7399), .B2(P2_REG2_REG_7__SCAN_IN), .A(n7398), .ZN(
        n7400) );
  AOI22_X1 U9168 ( .A1(n7401), .A2(n10043), .B1(n10056), .B2(n7400), .ZN(n7402) );
  NAND2_X1 U9169 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7863) );
  OAI211_X1 U9170 ( .C1(n10023), .C2(n7403), .A(n7402), .B(n7863), .ZN(n7404)
         );
  AOI21_X1 U9171 ( .B1(n10045), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n7404), .ZN(
        n7410) );
  AND3_X1 U9172 ( .A1(n7423), .A2(n7406), .A3(n7405), .ZN(n7407) );
  OAI21_X1 U9173 ( .B1(n7408), .B2(n7407), .A(n10051), .ZN(n7409) );
  NAND2_X1 U9174 ( .A1(n7410), .A2(n7409), .ZN(P2_U3189) );
  INV_X1 U9175 ( .A(n10045), .ZN(n8518) );
  INV_X1 U9176 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7429) );
  NAND3_X1 U9177 ( .A1(n7431), .A2(n7412), .A3(n7411), .ZN(n7413) );
  AOI21_X1 U9178 ( .B1(n4447), .B2(n7413), .A(n10032), .ZN(n7422) );
  INV_X1 U9179 ( .A(n7414), .ZN(n7416) );
  NAND3_X1 U9180 ( .A1(n7435), .A2(n7416), .A3(n7415), .ZN(n7417) );
  AOI21_X1 U9181 ( .B1(n7418), .B2(n7417), .A(n8486), .ZN(n7421) );
  NAND2_X1 U9182 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7641) );
  OAI21_X1 U9183 ( .B1(n10023), .B2(n7419), .A(n7641), .ZN(n7420) );
  NOR3_X1 U9184 ( .A1(n7422), .A2(n7421), .A3(n7420), .ZN(n7428) );
  OAI21_X1 U9185 ( .B1(n7425), .B2(n7424), .A(n7423), .ZN(n7426) );
  NAND2_X1 U9186 ( .A1(n7426), .A2(n10051), .ZN(n7427) );
  OAI211_X1 U9187 ( .C1(n8518), .C2(n7429), .A(n7428), .B(n7427), .ZN(P2_U3188) );
  INV_X1 U9188 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n7447) );
  NOR2_X1 U9189 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5026), .ZN(n7584) );
  INV_X1 U9190 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7727) );
  INV_X1 U9191 ( .A(n7430), .ZN(n7433) );
  INV_X1 U9192 ( .A(n7431), .ZN(n7432) );
  AOI21_X1 U9193 ( .B1(n7727), .B2(n7433), .A(n7432), .ZN(n7439) );
  INV_X1 U9194 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7619) );
  INV_X1 U9195 ( .A(n7434), .ZN(n7437) );
  INV_X1 U9196 ( .A(n7435), .ZN(n7436) );
  AOI21_X1 U9197 ( .B1(n7619), .B2(n7437), .A(n7436), .ZN(n7438) );
  OAI22_X1 U9198 ( .A1(n7439), .A2(n10032), .B1(n7438), .B2(n8486), .ZN(n7440)
         );
  AOI211_X1 U9199 ( .C1(n7441), .C2(n10047), .A(n7584), .B(n7440), .ZN(n7446)
         );
  XOR2_X1 U9200 ( .A(n7443), .B(n7442), .Z(n7444) );
  NAND2_X1 U9201 ( .A1(n7444), .A2(n10051), .ZN(n7445) );
  OAI211_X1 U9202 ( .C1(n7447), .C2(n8518), .A(n7446), .B(n7445), .ZN(P2_U3187) );
  INV_X1 U9203 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7786) );
  INV_X1 U9204 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7448) );
  OR2_X1 U9205 ( .A1(n7464), .A2(n7448), .ZN(n7449) );
  NAND2_X1 U9206 ( .A1(n7450), .A2(n7449), .ZN(n7665) );
  XNOR2_X1 U9207 ( .A(n7665), .B(n7666), .ZN(n7451) );
  AOI21_X1 U9208 ( .B1(n7786), .B2(n7451), .A(n7664), .ZN(n7470) );
  NOR2_X1 U9209 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5030), .ZN(n8294) );
  INV_X1 U9210 ( .A(n8294), .ZN(n7452) );
  OAI21_X1 U9211 ( .B1(n10023), .B2(n7666), .A(n7452), .ZN(n7460) );
  AOI21_X1 U9212 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n7454), .A(n7453), .ZN(
        n7456) );
  INV_X1 U9213 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7794) );
  AOI21_X1 U9214 ( .B1(n7457), .B2(n7794), .A(n7649), .ZN(n7458) );
  NOR2_X1 U9215 ( .A1(n7458), .A2(n10032), .ZN(n7459) );
  AOI211_X1 U9216 ( .C1(n10045), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n7460), .B(
        n7459), .ZN(n7469) );
  INV_X1 U9217 ( .A(n7461), .ZN(n7463) );
  AOI21_X1 U9218 ( .B1(n7464), .B2(n7463), .A(n7462), .ZN(n7657) );
  MUX2_X1 U9219 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8529), .Z(n7465) );
  OR2_X1 U9220 ( .A1(n7465), .A2(n7666), .ZN(n7656) );
  NAND2_X1 U9221 ( .A1(n7465), .A2(n7666), .ZN(n7655) );
  NAND2_X1 U9222 ( .A1(n7656), .A2(n7655), .ZN(n7466) );
  XNOR2_X1 U9223 ( .A(n7657), .B(n7466), .ZN(n7467) );
  NAND2_X1 U9224 ( .A1(n7467), .A2(n10051), .ZN(n7468) );
  OAI211_X1 U9225 ( .C1(n7470), .C2(n8486), .A(n7469), .B(n7468), .ZN(P2_U3191) );
  OR2_X1 U9226 ( .A1(n7471), .A2(n7475), .ZN(n7472) );
  NAND2_X1 U9227 ( .A1(n7473), .A2(n7472), .ZN(n7597) );
  INV_X1 U9228 ( .A(n7597), .ZN(n7487) );
  INV_X1 U9229 ( .A(n9062), .ZN(n9050) );
  AOI21_X1 U9230 ( .B1(n7474), .B2(n9049), .A(n9050), .ZN(n7476) );
  NOR2_X1 U9231 ( .A1(n7476), .A2(n7475), .ZN(n9927) );
  AOI21_X1 U9232 ( .B1(n7476), .B2(n7475), .A(n9927), .ZN(n7477) );
  OAI222_X1 U9233 ( .A1(n7914), .A2(n7836), .B1(n7913), .B2(n7478), .C1(n9934), 
        .C2(n7477), .ZN(n7595) );
  NAND2_X1 U9234 ( .A1(n7595), .A2(n9598), .ZN(n7486) );
  AOI211_X1 U9235 ( .C1(n7598), .C2(n7479), .A(n9590), .B(n9944), .ZN(n7596)
         );
  NOR2_X1 U9236 ( .A1(n9955), .A2(n5756), .ZN(n7484) );
  INV_X1 U9237 ( .A(n7480), .ZN(n7481) );
  OAI22_X1 U9238 ( .A1(n9598), .A2(n7482), .B1(n7481), .B2(n9515), .ZN(n7483)
         );
  AOI211_X1 U9239 ( .C1(n7596), .C2(n9949), .A(n7484), .B(n7483), .ZN(n7485)
         );
  OAI211_X1 U9240 ( .C1(n7487), .C2(n9601), .A(n7486), .B(n7485), .ZN(P1_U3286) );
  INV_X1 U9241 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7508) );
  INV_X1 U9242 ( .A(n7488), .ZN(n7490) );
  NAND3_X1 U9243 ( .A1(n10053), .A2(n7490), .A3(n7489), .ZN(n7491) );
  AOI21_X1 U9244 ( .B1(n7492), .B2(n7491), .A(n8486), .ZN(n7501) );
  INV_X1 U9245 ( .A(n7493), .ZN(n7497) );
  NAND3_X1 U9246 ( .A1(n10041), .A2(n7495), .A3(n7494), .ZN(n7496) );
  AOI21_X1 U9247 ( .B1(n7497), .B2(n7496), .A(n10032), .ZN(n7500) );
  NAND2_X1 U9248 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7539) );
  OAI21_X1 U9249 ( .B1(n10023), .B2(n7498), .A(n7539), .ZN(n7499) );
  NOR3_X1 U9250 ( .A1(n7501), .A2(n7500), .A3(n7499), .ZN(n7507) );
  AND2_X1 U9251 ( .A1(n10048), .A2(n7502), .ZN(n7505) );
  OAI211_X1 U9252 ( .C1(n7505), .C2(n7504), .A(n10051), .B(n7503), .ZN(n7506)
         );
  OAI211_X1 U9253 ( .C1(n8518), .C2(n7508), .A(n7507), .B(n7506), .ZN(P2_U3186) );
  INV_X1 U9254 ( .A(n9052), .ZN(n7509) );
  OAI21_X1 U9255 ( .B1(n9927), .B2(n7509), .A(n9065), .ZN(n7510) );
  XOR2_X1 U9256 ( .A(n7518), .B(n7510), .Z(n7511) );
  AOI22_X1 U9257 ( .A1(n7511), .A2(n9906), .B1(n9932), .B2(n9922), .ZN(n9988)
         );
  XNOR2_X1 U9258 ( .A(n9941), .B(n7512), .ZN(n7514) );
  AOI22_X1 U9259 ( .A1(n7514), .A2(n9942), .B1(n7513), .B2(n9279), .ZN(n9987)
         );
  INV_X1 U9260 ( .A(n9987), .ZN(n7517) );
  AOI22_X1 U9261 ( .A1(n9593), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7839), .B2(
        n9952), .ZN(n7515) );
  OAI21_X1 U9262 ( .B1(n9989), .B2(n9955), .A(n7515), .ZN(n7516) );
  AOI21_X1 U9263 ( .B1(n7517), .B2(n9949), .A(n7516), .ZN(n7521) );
  XNOR2_X1 U9264 ( .A(n7519), .B(n7518), .ZN(n9991) );
  NAND2_X1 U9265 ( .A1(n9991), .A2(n9959), .ZN(n7520) );
  OAI211_X1 U9266 ( .C1(n9988), .C2(n9576), .A(n7521), .B(n7520), .ZN(P1_U3284) );
  XNOR2_X1 U9267 ( .A(n7522), .B(n5179), .ZN(n7752) );
  XNOR2_X1 U9268 ( .A(n7523), .B(n5179), .ZN(n7524) );
  OAI222_X1 U9269 ( .A1(n8669), .A2(n7864), .B1(n8711), .B2(n7955), .C1(n8666), 
        .C2(n7524), .ZN(n7748) );
  AOI21_X1 U9270 ( .B1(n7752), .B2(n8794), .A(n7748), .ZN(n7929) );
  INV_X1 U9271 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7525) );
  OAI22_X1 U9272 ( .A1(n8841), .A2(n7526), .B1(n7525), .B2(n10088), .ZN(n7527)
         );
  INV_X1 U9273 ( .A(n7527), .ZN(n7528) );
  OAI21_X1 U9274 ( .B1(n7929), .B2(n10091), .A(n7528), .ZN(P2_U3411) );
  NAND2_X1 U9275 ( .A1(n8359), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n7529) );
  OAI21_X1 U9276 ( .B1(n8549), .B2(n8359), .A(n7529), .ZN(P2_U3522) );
  NAND2_X1 U9277 ( .A1(n8359), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7530) );
  OAI21_X1 U9278 ( .B1(n8563), .B2(n8359), .A(n7530), .ZN(P2_U3520) );
  INV_X1 U9279 ( .A(n7531), .ZN(n7533) );
  XNOR2_X1 U9280 ( .A(n8173), .B(n7542), .ZN(n7534) );
  INV_X1 U9281 ( .A(n7534), .ZN(n7535) );
  AND2_X1 U9282 ( .A1(n7534), .A2(n7614), .ZN(n7578) );
  AOI21_X1 U9283 ( .B1(n7535), .B2(n8369), .A(n7578), .ZN(n7536) );
  OAI21_X1 U9284 ( .B1(n7537), .B2(n7536), .A(n7581), .ZN(n7538) );
  NAND2_X1 U9285 ( .A1(n7538), .A2(n8321), .ZN(n7544) );
  INV_X1 U9286 ( .A(n7539), .ZN(n7541) );
  OAI22_X1 U9287 ( .A1(n8324), .A2(n7629), .B1(n7642), .B2(n8347), .ZN(n7540)
         );
  AOI211_X1 U9288 ( .C1(n7542), .C2(n8339), .A(n7541), .B(n7540), .ZN(n7543)
         );
  OAI211_X1 U9289 ( .C1(n7690), .C2(n8348), .A(n7544), .B(n7543), .ZN(P2_U3170) );
  NAND2_X1 U9290 ( .A1(n7611), .A2(n7545), .ZN(n7546) );
  XNOR2_X1 U9291 ( .A(n7546), .B(n7548), .ZN(n7588) );
  XNOR2_X1 U9292 ( .A(n7547), .B(n7548), .ZN(n7549) );
  AOI222_X1 U9293 ( .A1(n8731), .A2(n7549), .B1(n8366), .B2(n8728), .C1(n8368), 
        .C2(n8726), .ZN(n7589) );
  OAI21_X1 U9294 ( .B1(n7550), .B2(n8745), .A(n7589), .ZN(n7551) );
  AOI21_X1 U9295 ( .B1(n8794), .B2(n7588), .A(n7551), .ZN(n10078) );
  OR2_X1 U9296 ( .A1(n8786), .A2(n4625), .ZN(n7552) );
  OAI21_X1 U9297 ( .B1(n10078), .B2(n8066), .A(n7552), .ZN(P2_U3465) );
  INV_X1 U9298 ( .A(n7553), .ZN(n7555) );
  INV_X1 U9299 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7554) );
  OAI222_X1 U9300 ( .A1(n5543), .A2(P2_U3151), .B1(n6665), .B2(n7555), .C1(
        n7554), .C2(n8880), .ZN(P2_U3276) );
  INV_X1 U9301 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7556) );
  OAI222_X1 U9302 ( .A1(n9729), .A2(n7556), .B1(n9732), .B2(n7555), .C1(
        P1_U3086), .C2(n9381), .ZN(P1_U3336) );
  XNOR2_X1 U9303 ( .A(n7557), .B(n7560), .ZN(n7605) );
  INV_X1 U9304 ( .A(n7605), .ZN(n7569) );
  INV_X1 U9305 ( .A(n7558), .ZN(n7561) );
  OAI211_X1 U9306 ( .C1(n7561), .C2(n7560), .A(n9906), .B(n7559), .ZN(n7563)
         );
  AOI22_X1 U9307 ( .A1(n9932), .A2(n9279), .B1(n9278), .B2(n7513), .ZN(n7562)
         );
  NAND2_X1 U9308 ( .A1(n7563), .A2(n7562), .ZN(n7603) );
  AOI211_X1 U9309 ( .C1(n7882), .C2(n7564), .A(n9590), .B(n4437), .ZN(n7604)
         );
  NAND2_X1 U9310 ( .A1(n7604), .A2(n9949), .ZN(n7566) );
  AOI22_X1 U9311 ( .A1(n9593), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7881), .B2(
        n9952), .ZN(n7565) );
  OAI211_X1 U9312 ( .C1(n4570), .C2(n9955), .A(n7566), .B(n7565), .ZN(n7567)
         );
  AOI21_X1 U9313 ( .B1(n9598), .B2(n7603), .A(n7567), .ZN(n7568) );
  OAI21_X1 U9314 ( .B1(n7569), .B2(n9601), .A(n7568), .ZN(P1_U3282) );
  OR2_X1 U9315 ( .A1(n5543), .A2(n7570), .ZN(n7618) );
  NAND2_X1 U9316 ( .A1(n7892), .A2(n7618), .ZN(n7571) );
  MUX2_X1 U9317 ( .A(n7573), .B(n7572), .S(n8715), .Z(n7576) );
  AOI22_X1 U9318 ( .A1(n8735), .A2(n7574), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8719), .ZN(n7575) );
  OAI211_X1 U9319 ( .C1(n8738), .C2(n7577), .A(n7576), .B(n7575), .ZN(P2_U3232) );
  INV_X1 U9320 ( .A(n7578), .ZN(n7579) );
  XNOR2_X1 U9321 ( .A(n8173), .B(n7585), .ZN(n7638) );
  XOR2_X1 U9322 ( .A(n8368), .B(n7638), .Z(n7580) );
  AND3_X1 U9323 ( .A1(n7581), .A2(n7580), .A3(n7579), .ZN(n7582) );
  OAI21_X1 U9324 ( .B1(n7637), .B2(n7582), .A(n8321), .ZN(n7587) );
  OAI22_X1 U9325 ( .A1(n8324), .A2(n7614), .B1(n7864), .B2(n8347), .ZN(n7583)
         );
  AOI211_X1 U9326 ( .C1(n7585), .C2(n8339), .A(n7584), .B(n7583), .ZN(n7586)
         );
  OAI211_X1 U9327 ( .C1(n7620), .C2(n8348), .A(n7587), .B(n7586), .ZN(P2_U3167) );
  INV_X1 U9328 ( .A(n7588), .ZN(n7594) );
  MUX2_X1 U9329 ( .A(n7590), .B(n7589), .S(n8715), .Z(n7593) );
  INV_X1 U9330 ( .A(n7648), .ZN(n7591) );
  AOI22_X1 U9331 ( .A1(n8735), .A2(n7645), .B1(n8719), .B2(n7591), .ZN(n7592)
         );
  OAI211_X1 U9332 ( .C1(n7594), .C2(n8738), .A(n7593), .B(n7592), .ZN(P2_U3227) );
  AOI211_X1 U9333 ( .C1(n10007), .C2(n7597), .A(n7596), .B(n7595), .ZN(n7602)
         );
  AOI22_X1 U9334 ( .A1(n6101), .A2(n7598), .B1(n10019), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n7599) );
  OAI21_X1 U9335 ( .B1(n7602), .B2(n10019), .A(n7599), .ZN(P1_U3529) );
  OAI22_X1 U9336 ( .A1(n9709), .A2(n5756), .B1(n10010), .B2(n5749), .ZN(n7600)
         );
  INV_X1 U9337 ( .A(n7600), .ZN(n7601) );
  OAI21_X1 U9338 ( .B1(n7602), .B2(n10009), .A(n7601), .ZN(P1_U3474) );
  AOI211_X1 U9339 ( .C1(n7605), .C2(n10007), .A(n7604), .B(n7603), .ZN(n7609)
         );
  AOI22_X1 U9340 ( .A1(n7882), .A2(n6101), .B1(n10019), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n7606) );
  OAI21_X1 U9341 ( .B1(n7609), .B2(n10019), .A(n7606), .ZN(P1_U3533) );
  NOR2_X1 U9342 ( .A1(n10010), .A2(n5807), .ZN(n7607) );
  AOI21_X1 U9343 ( .B1(n7882), .B2(n6137), .A(n7607), .ZN(n7608) );
  OAI21_X1 U9344 ( .B1(n7609), .B2(n10009), .A(n7608), .ZN(P1_U3486) );
  XOR2_X1 U9345 ( .A(n7610), .B(n7612), .Z(n7617) );
  OAI21_X1 U9346 ( .B1(n7613), .B2(n7612), .A(n7611), .ZN(n7724) );
  INV_X1 U9347 ( .A(n7892), .ZN(n7632) );
  OAI22_X1 U9348 ( .A1(n7864), .A2(n8711), .B1(n7614), .B2(n8669), .ZN(n7615)
         );
  AOI21_X1 U9349 ( .B1(n7724), .B2(n7632), .A(n7615), .ZN(n7616) );
  OAI21_X1 U9350 ( .B1(n8666), .B2(n7617), .A(n7616), .ZN(n7722) );
  INV_X1 U9351 ( .A(n7722), .ZN(n7625) );
  INV_X1 U9352 ( .A(n7618), .ZN(n10068) );
  NAND2_X1 U9353 ( .A1(n8715), .A2(n10068), .ZN(n7898) );
  INV_X1 U9354 ( .A(n7898), .ZN(n7623) );
  NOR2_X1 U9355 ( .A1(n8715), .A2(n7619), .ZN(n7622) );
  OAI22_X1 U9356 ( .A1(n8594), .A2(n7721), .B1(n7620), .B2(n10064), .ZN(n7621)
         );
  AOI211_X1 U9357 ( .C1(n7724), .C2(n7623), .A(n7622), .B(n7621), .ZN(n7624)
         );
  OAI21_X1 U9358 ( .B1(n7625), .B2(n8734), .A(n7624), .ZN(P2_U3228) );
  INV_X1 U9359 ( .A(n7899), .ZN(n7725) );
  OAI21_X1 U9360 ( .B1(n7627), .B2(n5527), .A(n7626), .ZN(n10067) );
  NOR2_X1 U9361 ( .A1(n10062), .A2(n8745), .ZN(n7635) );
  XNOR2_X1 U9362 ( .A(n7628), .B(n5527), .ZN(n7634) );
  OAI22_X1 U9363 ( .A1(n7630), .A2(n8669), .B1(n7629), .B2(n8711), .ZN(n7631)
         );
  AOI21_X1 U9364 ( .B1(n10067), .B2(n7632), .A(n7631), .ZN(n7633) );
  OAI21_X1 U9365 ( .B1(n8666), .B2(n7634), .A(n7633), .ZN(n10065) );
  AOI211_X1 U9366 ( .C1(n7725), .C2(n10067), .A(n7635), .B(n10065), .ZN(n10073) );
  NAND2_X1 U9367 ( .A1(n8755), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7636) );
  OAI21_X1 U9368 ( .B1(n10073), .B2(n8066), .A(n7636), .ZN(P2_U3461) );
  AOI21_X1 U9369 ( .B1(n7642), .B2(n7638), .A(n7637), .ZN(n7640) );
  XNOR2_X1 U9370 ( .A(n8173), .B(n7645), .ZN(n7857) );
  XNOR2_X1 U9371 ( .A(n7857), .B(n8367), .ZN(n7639) );
  NAND2_X1 U9372 ( .A1(n7640), .A2(n7639), .ZN(n7859) );
  OAI211_X1 U9373 ( .C1(n7640), .C2(n7639), .A(n7859), .B(n8321), .ZN(n7647)
         );
  INV_X1 U9374 ( .A(n7641), .ZN(n7644) );
  OAI22_X1 U9375 ( .A1(n8324), .A2(n7642), .B1(n7960), .B2(n8347), .ZN(n7643)
         );
  AOI211_X1 U9376 ( .C1(n7645), .C2(n8339), .A(n7644), .B(n7643), .ZN(n7646)
         );
  OAI211_X1 U9377 ( .C1(n7648), .C2(n8348), .A(n7647), .B(n7646), .ZN(P2_U3179) );
  NAND2_X1 U9378 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n7708), .ZN(n7651) );
  OAI21_X1 U9379 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n7708), .A(n7651), .ZN(
        n7652) );
  AOI21_X1 U9380 ( .B1(n7653), .B2(n7652), .A(n7705), .ZN(n7673) );
  MUX2_X1 U9381 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8529), .Z(n7709) );
  XNOR2_X1 U9382 ( .A(n7709), .B(n7654), .ZN(n7660) );
  INV_X1 U9383 ( .A(n7655), .ZN(n7658) );
  OAI21_X1 U9384 ( .B1(n7660), .B2(n7659), .A(n7710), .ZN(n7662) );
  NOR2_X1 U9385 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7661), .ZN(n8049) );
  AOI21_X1 U9386 ( .B1(n10051), .B2(n7662), .A(n8049), .ZN(n7663) );
  OAI21_X1 U9387 ( .B1(n10023), .B2(n7708), .A(n7663), .ZN(n7671) );
  NAND2_X1 U9388 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n7708), .ZN(n7667) );
  OAI21_X1 U9389 ( .B1(n7708), .B2(P2_REG2_REG_10__SCAN_IN), .A(n7667), .ZN(
        n7668) );
  AOI21_X1 U9390 ( .B1(n4368), .B2(n7668), .A(n4443), .ZN(n7669) );
  NOR2_X1 U9391 ( .A1(n7669), .A2(n8486), .ZN(n7670) );
  AOI211_X1 U9392 ( .C1(n10045), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n7671), .B(
        n7670), .ZN(n7672) );
  OAI21_X1 U9393 ( .B1(n7673), .B2(n10032), .A(n7672), .ZN(P2_U3192) );
  INV_X1 U9394 ( .A(n7674), .ZN(n7686) );
  OAI222_X1 U9395 ( .A1(n9732), .A2(n7686), .B1(n9204), .B2(P1_U3086), .C1(
        n7675), .C2(n9729), .ZN(P1_U3335) );
  NOR2_X1 U9396 ( .A1(n7676), .A2(n7677), .ZN(n7829) );
  AOI21_X1 U9397 ( .B1(n7677), .B2(n7676), .A(n7829), .ZN(n7684) );
  NAND2_X1 U9398 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9761) );
  INV_X1 U9399 ( .A(n9761), .ZN(n7678) );
  AOI21_X1 U9400 ( .B1(n8999), .B2(n9930), .A(n7678), .ZN(n7680) );
  NAND2_X1 U9401 ( .A1(n9004), .A2(n9938), .ZN(n7679) );
  OAI211_X1 U9402 ( .C1(n7681), .C2(n9001), .A(n7680), .B(n7679), .ZN(n7682)
         );
  AOI21_X1 U9403 ( .B1(n9940), .B2(n8972), .A(n7682), .ZN(n7683) );
  OAI21_X1 U9404 ( .B1(n7684), .B2(n8974), .A(n7683), .ZN(P1_U3221) );
  INV_X1 U9405 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7685) );
  OAI222_X1 U9406 ( .A1(P2_U3151), .A2(n7687), .B1(n6665), .B2(n7686), .C1(
        n7685), .C2(n8880), .ZN(P2_U3275) );
  OAI21_X1 U9407 ( .B1(n7689), .B2(n7691), .A(n7688), .ZN(n7746) );
  OAI22_X1 U9408 ( .A1(n8594), .A2(n7743), .B1(n7690), .B2(n10064), .ZN(n7697)
         );
  XNOR2_X1 U9409 ( .A(n7692), .B(n7691), .ZN(n7693) );
  NAND2_X1 U9410 ( .A1(n7693), .A2(n8731), .ZN(n7695) );
  AOI22_X1 U9411 ( .A1(n8726), .A2(n8370), .B1(n8368), .B2(n8728), .ZN(n7694)
         );
  NAND2_X1 U9412 ( .A1(n7695), .A2(n7694), .ZN(n7744) );
  MUX2_X1 U9413 ( .A(n7744), .B(P2_REG2_REG_4__SCAN_IN), .S(n8734), .Z(n7696)
         );
  AOI211_X1 U9414 ( .C1(n8596), .C2(n7746), .A(n7697), .B(n7696), .ZN(n7698)
         );
  INV_X1 U9415 ( .A(n7698), .ZN(P2_U3229) );
  OAI22_X1 U9416 ( .A1(n8594), .A2(n7699), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n10064), .ZN(n7702) );
  MUX2_X1 U9417 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n7700), .S(n8715), .Z(n7701)
         );
  AOI211_X1 U9418 ( .C1(n8596), .C2(n7703), .A(n7702), .B(n7701), .ZN(n7704)
         );
  INV_X1 U9419 ( .A(n7704), .ZN(P2_U3230) );
  XNOR2_X1 U9420 ( .A(n7806), .B(n7820), .ZN(n7706) );
  AOI21_X1 U9421 ( .B1(n5232), .B2(n7706), .A(n7808), .ZN(n7720) );
  XNOR2_X1 U9422 ( .A(n7820), .B(n7810), .ZN(n7707) );
  AOI21_X1 U9423 ( .B1(n7707), .B2(n7935), .A(n7811), .ZN(n7717) );
  MUX2_X1 U9424 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8529), .Z(n7819) );
  XNOR2_X1 U9425 ( .A(n7819), .B(n7820), .ZN(n7713) );
  OR2_X1 U9426 ( .A1(n7709), .A2(n7708), .ZN(n7711) );
  NAND2_X1 U9427 ( .A1(n7711), .A2(n7710), .ZN(n7712) );
  NAND2_X1 U9428 ( .A1(n7713), .A2(n7712), .ZN(n7822) );
  OAI21_X1 U9429 ( .B1(n7713), .B2(n7712), .A(n7822), .ZN(n7714) );
  AND2_X1 U9430 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8094) );
  AOI21_X1 U9431 ( .B1(n10051), .B2(n7714), .A(n8094), .ZN(n7716) );
  NAND2_X1 U9432 ( .A1(n10047), .A2(n7820), .ZN(n7715) );
  OAI211_X1 U9433 ( .C1(n8486), .C2(n7717), .A(n7716), .B(n7715), .ZN(n7718)
         );
  AOI21_X1 U9434 ( .B1(n10045), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n7718), .ZN(
        n7719) );
  OAI21_X1 U9435 ( .B1(n7720), .B2(n10032), .A(n7719), .ZN(P2_U3193) );
  NOR2_X1 U9436 ( .A1(n7721), .A2(n8745), .ZN(n7723) );
  AOI211_X1 U9437 ( .C1(n7725), .C2(n7724), .A(n7723), .B(n7722), .ZN(n10076)
         );
  OR2_X1 U9438 ( .A1(n10076), .A2(n8755), .ZN(n7726) );
  OAI21_X1 U9439 ( .B1(n8786), .B2(n7727), .A(n7726), .ZN(P2_U3464) );
  INV_X1 U9440 ( .A(n7728), .ZN(n7733) );
  NAND2_X1 U9441 ( .A1(n8118), .A2(n8666), .ZN(n7732) );
  OAI21_X1 U9442 ( .B1(n7730), .B2(n8745), .A(n7729), .ZN(n7731) );
  AOI21_X1 U9443 ( .B1(n7733), .B2(n7732), .A(n7731), .ZN(n10071) );
  OR2_X1 U9444 ( .A1(n10071), .A2(n8755), .ZN(n7734) );
  OAI21_X1 U9445 ( .B1(n8786), .B2(n6960), .A(n7734), .ZN(P2_U3459) );
  XNOR2_X1 U9446 ( .A(n7735), .B(n7737), .ZN(n7779) );
  NOR2_X1 U9447 ( .A1(n7954), .A2(n8745), .ZN(n7741) );
  OAI211_X1 U9448 ( .C1(n7738), .C2(n7737), .A(n7736), .B(n8731), .ZN(n7740)
         );
  AOI22_X1 U9449 ( .A1(n8726), .A2(n8366), .B1(n8364), .B2(n8728), .ZN(n7739)
         );
  NAND2_X1 U9450 ( .A1(n7740), .A2(n7739), .ZN(n7776) );
  AOI211_X1 U9451 ( .C1(n8794), .C2(n7779), .A(n7741), .B(n7776), .ZN(n10080)
         );
  OR2_X1 U9452 ( .A1(n10080), .A2(n8755), .ZN(n7742) );
  OAI21_X1 U9453 ( .B1(n8786), .B2(n7010), .A(n7742), .ZN(P2_U3467) );
  NOR2_X1 U9454 ( .A1(n7743), .A2(n8745), .ZN(n7745) );
  AOI211_X1 U9455 ( .C1(n8794), .C2(n7746), .A(n7745), .B(n7744), .ZN(n10075)
         );
  OR2_X1 U9456 ( .A1(n10075), .A2(n8755), .ZN(n7747) );
  OAI21_X1 U9457 ( .B1(n8786), .B2(n7003), .A(n7747), .ZN(P2_U3463) );
  INV_X1 U9458 ( .A(n7748), .ZN(n7754) );
  INV_X1 U9459 ( .A(n7749), .ZN(n7867) );
  AOI22_X1 U9460 ( .A1(n8735), .A2(n7927), .B1(n8719), .B2(n7867), .ZN(n7750)
         );
  OAI21_X1 U9461 ( .B1(n4708), .B2(n10069), .A(n7750), .ZN(n7751) );
  AOI21_X1 U9462 ( .B1(n7752), .B2(n8596), .A(n7751), .ZN(n7753) );
  OAI21_X1 U9463 ( .B1(n7754), .B2(n8734), .A(n7753), .ZN(P2_U3226) );
  OAI21_X1 U9464 ( .B1(n7757), .B2(n7756), .A(n7755), .ZN(n7758) );
  NAND2_X1 U9465 ( .A1(n7758), .A2(n8997), .ZN(n7763) );
  AOI21_X1 U9466 ( .B1(n8984), .B2(n9910), .A(n7759), .ZN(n7760) );
  OAI21_X1 U9467 ( .B1(n7988), .B2(n8981), .A(n7760), .ZN(n7761) );
  AOI21_X1 U9468 ( .B1(n9913), .B2(n9004), .A(n7761), .ZN(n7762) );
  OAI211_X1 U9469 ( .C1(n9999), .C2(n9008), .A(n7763), .B(n7762), .ZN(P1_U3224) );
  INV_X1 U9470 ( .A(n9907), .ZN(n7766) );
  OAI21_X1 U9471 ( .B1(n7766), .B2(n7765), .A(n7764), .ZN(n7768) );
  NAND2_X1 U9472 ( .A1(n7768), .A2(n7767), .ZN(n7769) );
  AOI222_X1 U9473 ( .A1(n9906), .A2(n7769), .B1(n9277), .B2(n7513), .C1(n9278), 
        .C2(n9932), .ZN(n10003) );
  XNOR2_X1 U9474 ( .A(n7770), .B(n9034), .ZN(n10008) );
  NAND2_X1 U9475 ( .A1(n10008), .A2(n9959), .ZN(n7775) );
  OAI211_X1 U9476 ( .C1(n9917), .C2(n10005), .A(n9942), .B(n7919), .ZN(n10002)
         );
  INV_X1 U9477 ( .A(n10002), .ZN(n7773) );
  AOI22_X1 U9478 ( .A1(n9593), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7854), .B2(
        n9952), .ZN(n7771) );
  OAI21_X1 U9479 ( .B1(n10005), .B2(n9955), .A(n7771), .ZN(n7772) );
  AOI21_X1 U9480 ( .B1(n7773), .B2(n9949), .A(n7772), .ZN(n7774) );
  OAI211_X1 U9481 ( .C1(n9593), .C2(n10003), .A(n7775), .B(n7774), .ZN(
        P1_U3280) );
  OAI22_X1 U9482 ( .A1(n8594), .A2(n7954), .B1(n7966), .B2(n10064), .ZN(n7778)
         );
  MUX2_X1 U9483 ( .A(n7776), .B(P2_REG2_REG_8__SCAN_IN), .S(n8734), .Z(n7777)
         );
  AOI211_X1 U9484 ( .C1(n8596), .C2(n7779), .A(n7778), .B(n7777), .ZN(n7780)
         );
  INV_X1 U9485 ( .A(n7780), .ZN(P2_U3225) );
  XNOR2_X1 U9486 ( .A(n7781), .B(n5207), .ZN(n7791) );
  OAI21_X1 U9487 ( .B1(n4440), .B2(n5207), .A(n7782), .ZN(n7784) );
  OAI22_X1 U9488 ( .A1(n7955), .A2(n8669), .B1(n8024), .B2(n8711), .ZN(n7783)
         );
  AOI21_X1 U9489 ( .B1(n7784), .B2(n8731), .A(n7783), .ZN(n7785) );
  OAI21_X1 U9490 ( .B1(n7791), .B2(n7892), .A(n7785), .ZN(n7793) );
  NAND2_X1 U9491 ( .A1(n7793), .A2(n10069), .ZN(n7789) );
  OAI22_X1 U9492 ( .A1(n8715), .A2(n7786), .B1(n8295), .B2(n10064), .ZN(n7787)
         );
  AOI21_X1 U9493 ( .B1(n8735), .B2(n8296), .A(n7787), .ZN(n7788) );
  OAI211_X1 U9494 ( .C1(n7791), .C2(n7898), .A(n7789), .B(n7788), .ZN(P2_U3224) );
  OAI22_X1 U9495 ( .A1(n7791), .A2(n7899), .B1(n7790), .B2(n8745), .ZN(n7792)
         );
  NOR2_X1 U9496 ( .A1(n7793), .A2(n7792), .ZN(n10082) );
  OR2_X1 U9497 ( .A1(n8786), .A2(n7794), .ZN(n7795) );
  OAI21_X1 U9498 ( .B1(n10082), .B2(n8755), .A(n7795), .ZN(P2_U3468) );
  XNOR2_X1 U9499 ( .A(n7873), .B(n7796), .ZN(n7797) );
  NAND2_X1 U9500 ( .A1(n7797), .A2(n7798), .ZN(n7871) );
  OAI21_X1 U9501 ( .B1(n7798), .B2(n7797), .A(n7871), .ZN(n7799) );
  NAND2_X1 U9502 ( .A1(n7799), .A2(n8997), .ZN(n7805) );
  NAND2_X1 U9503 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n9747) );
  NAND2_X1 U9504 ( .A1(n8999), .A2(n9910), .ZN(n7800) );
  OAI211_X1 U9505 ( .C1(n7801), .C2(n9001), .A(n9747), .B(n7800), .ZN(n7802)
         );
  AOI21_X1 U9506 ( .B1(n7803), .B2(n9004), .A(n7802), .ZN(n7804) );
  OAI211_X1 U9507 ( .C1(n9993), .C2(n9008), .A(n7805), .B(n7804), .ZN(P1_U3217) );
  NOR2_X1 U9508 ( .A1(n7820), .A2(n7806), .ZN(n7807) );
  AOI22_X1 U9509 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n7813), .B1(n8388), .B2(
        n8382), .ZN(n7809) );
  AOI21_X1 U9510 ( .B1(n4435), .B2(n7809), .A(n8383), .ZN(n7828) );
  NAND2_X1 U9511 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8039) );
  OAI21_X1 U9512 ( .B1(n10023), .B2(n8388), .A(n8039), .ZN(n7817) );
  NOR2_X1 U9513 ( .A1(n7820), .A2(n7810), .ZN(n7812) );
  MUX2_X1 U9514 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n7979), .S(n7813), .Z(n7814)
         );
  AOI21_X1 U9515 ( .B1(n4434), .B2(n7814), .A(n8387), .ZN(n7815) );
  NOR2_X1 U9516 ( .A1(n7815), .A2(n8486), .ZN(n7816) );
  AOI211_X1 U9517 ( .C1(n10045), .C2(P2_ADDR_REG_12__SCAN_IN), .A(n7817), .B(
        n7816), .ZN(n7827) );
  MUX2_X1 U9518 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8529), .Z(n7818) );
  AND2_X1 U9519 ( .A1(n7818), .A2(n8388), .ZN(n8372) );
  NOR2_X1 U9520 ( .A1(n7818), .A2(n8388), .ZN(n8375) );
  NOR2_X1 U9521 ( .A1(n8372), .A2(n8375), .ZN(n7824) );
  INV_X1 U9522 ( .A(n7819), .ZN(n7821) );
  NAND2_X1 U9523 ( .A1(n7821), .A2(n7820), .ZN(n7823) );
  NAND2_X1 U9524 ( .A1(n7823), .A2(n7822), .ZN(n8374) );
  XNOR2_X1 U9525 ( .A(n7824), .B(n8374), .ZN(n7825) );
  NAND2_X1 U9526 ( .A1(n7825), .A2(n10051), .ZN(n7826) );
  OAI211_X1 U9527 ( .C1(n7828), .C2(n10032), .A(n7827), .B(n7826), .ZN(
        P2_U3194) );
  XNOR2_X1 U9528 ( .A(n7832), .B(n7831), .ZN(n7833) );
  XNOR2_X1 U9529 ( .A(n7834), .B(n7833), .ZN(n7841) );
  NAND2_X1 U9530 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n9777) );
  NAND2_X1 U9531 ( .A1(n8999), .A2(n9279), .ZN(n7835) );
  OAI211_X1 U9532 ( .C1(n7836), .C2(n9001), .A(n9777), .B(n7835), .ZN(n7838)
         );
  NOR2_X1 U9533 ( .A1(n9989), .A2(n9008), .ZN(n7837) );
  AOI211_X1 U9534 ( .C1(n7839), .C2(n9004), .A(n7838), .B(n7837), .ZN(n7840)
         );
  OAI21_X1 U9535 ( .B1(n7841), .B2(n8974), .A(n7840), .ZN(P1_U3231) );
  INV_X1 U9536 ( .A(n7842), .ZN(n7845) );
  OAI222_X1 U9537 ( .A1(n9729), .A2(n7843), .B1(n9732), .B2(n7845), .C1(n6397), 
        .C2(P1_U3086), .ZN(P1_U3334) );
  INV_X1 U9538 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7844) );
  OAI222_X1 U9539 ( .A1(n7846), .A2(P2_U3151), .B1(n6665), .B2(n7845), .C1(
        n7844), .C2(n8880), .ZN(P2_U3274) );
  OAI21_X1 U9540 ( .B1(n7849), .B2(n7848), .A(n7847), .ZN(n7850) );
  NAND2_X1 U9541 ( .A1(n7850), .A2(n8997), .ZN(n7856) );
  AND2_X1 U9542 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9831) );
  AOI21_X1 U9543 ( .B1(n8999), .B2(n9277), .A(n9831), .ZN(n7851) );
  OAI21_X1 U9544 ( .B1(n7852), .B2(n9001), .A(n7851), .ZN(n7853) );
  AOI21_X1 U9545 ( .B1(n7854), .B2(n9004), .A(n7853), .ZN(n7855) );
  OAI211_X1 U9546 ( .C1(n10005), .C2(n9008), .A(n7856), .B(n7855), .ZN(
        P1_U3234) );
  XNOR2_X1 U9547 ( .A(n8173), .B(n7927), .ZN(n7952) );
  XOR2_X1 U9548 ( .A(n8366), .B(n7952), .Z(n7862) );
  NAND2_X1 U9549 ( .A1(n7859), .A2(n7858), .ZN(n7861) );
  INV_X1 U9550 ( .A(n7953), .ZN(n7860) );
  AOI21_X1 U9551 ( .B1(n7862), .B2(n7861), .A(n7860), .ZN(n7870) );
  INV_X1 U9552 ( .A(n7863), .ZN(n7866) );
  OAI22_X1 U9553 ( .A1(n8324), .A2(n7864), .B1(n7955), .B2(n8347), .ZN(n7865)
         );
  AOI211_X1 U9554 ( .C1(n7927), .C2(n8339), .A(n7866), .B(n7865), .ZN(n7869)
         );
  NAND2_X1 U9555 ( .A1(n8335), .A2(n7867), .ZN(n7868) );
  OAI211_X1 U9556 ( .C1(n7870), .C2(n8342), .A(n7869), .B(n7868), .ZN(P2_U3153) );
  OAI21_X1 U9557 ( .B1(n7873), .B2(n7872), .A(n7871), .ZN(n7877) );
  XNOR2_X1 U9558 ( .A(n7875), .B(n7874), .ZN(n7876) );
  XNOR2_X1 U9559 ( .A(n7877), .B(n7876), .ZN(n7885) );
  NAND2_X1 U9560 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9819) );
  NAND2_X1 U9561 ( .A1(n8999), .A2(n9278), .ZN(n7878) );
  OAI211_X1 U9562 ( .C1(n7879), .C2(n9001), .A(n9819), .B(n7878), .ZN(n7880)
         );
  AOI21_X1 U9563 ( .B1(n7881), .B2(n9004), .A(n7880), .ZN(n7884) );
  NAND2_X1 U9564 ( .A1(n7882), .A2(n8972), .ZN(n7883) );
  OAI211_X1 U9565 ( .C1(n7885), .C2(n8974), .A(n7884), .B(n7883), .ZN(P1_U3236) );
  XNOR2_X1 U9566 ( .A(n7886), .B(n7888), .ZN(n7900) );
  XOR2_X1 U9567 ( .A(n7888), .B(n7887), .Z(n7890) );
  OAI22_X1 U9568 ( .A1(n7959), .A2(n8669), .B1(n8052), .B2(n8711), .ZN(n7889)
         );
  AOI21_X1 U9569 ( .B1(n7890), .B2(n8731), .A(n7889), .ZN(n7891) );
  OAI21_X1 U9570 ( .B1(n7900), .B2(n7892), .A(n7891), .ZN(n7902) );
  NAND2_X1 U9571 ( .A1(n7902), .A2(n10069), .ZN(n7897) );
  OAI22_X1 U9572 ( .A1(n8715), .A2(n7893), .B1(n8048), .B2(n10064), .ZN(n7894)
         );
  AOI21_X1 U9573 ( .B1(n8735), .B2(n7895), .A(n7894), .ZN(n7896) );
  OAI211_X1 U9574 ( .C1(n7900), .C2(n7898), .A(n7897), .B(n7896), .ZN(P2_U3223) );
  OAI22_X1 U9575 ( .A1(n7900), .A2(n7899), .B1(n8053), .B2(n8745), .ZN(n7901)
         );
  NOR2_X1 U9576 ( .A1(n7902), .A2(n7901), .ZN(n10084) );
  OR2_X1 U9577 ( .A1(n8786), .A2(n5217), .ZN(n7903) );
  OAI21_X1 U9578 ( .B1(n10084), .B2(n8066), .A(n7903), .ZN(P2_U3469) );
  OAI22_X1 U9579 ( .A1(n7905), .A2(n8774), .B1(n8786), .B2(n7904), .ZN(n7906)
         );
  AOI21_X1 U9580 ( .B1(n7907), .B2(n8786), .A(n7906), .ZN(n7908) );
  INV_X1 U9581 ( .A(n7908), .ZN(P2_U3460) );
  XNOR2_X1 U9582 ( .A(n7909), .B(n9088), .ZN(n9677) );
  INV_X1 U9583 ( .A(n7910), .ZN(n9937) );
  AOI211_X1 U9584 ( .C1(n9088), .C2(n7912), .A(n9934), .B(n7911), .ZN(n7916)
         );
  OAI22_X1 U9585 ( .A1(n8930), .A2(n7914), .B1(n7988), .B2(n7913), .ZN(n7915)
         );
  AOI211_X1 U9586 ( .C1(n9677), .C2(n9937), .A(n7916), .B(n7915), .ZN(n9682)
         );
  NOR2_X1 U9587 ( .A1(n9593), .A2(n7917), .ZN(n9946) );
  INV_X1 U9588 ( .A(n8010), .ZN(n7918) );
  AOI211_X1 U9589 ( .C1(n9679), .C2(n7919), .A(n9590), .B(n7918), .ZN(n9678)
         );
  NAND2_X1 U9590 ( .A1(n9678), .A2(n9949), .ZN(n7921) );
  AOI22_X1 U9591 ( .A1(n9593), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n7992), .B2(
        n9952), .ZN(n7920) );
  OAI211_X1 U9592 ( .C1(n7989), .C2(n9955), .A(n7921), .B(n7920), .ZN(n7922)
         );
  AOI21_X1 U9593 ( .B1(n9677), .B2(n9946), .A(n7922), .ZN(n7923) );
  OAI21_X1 U9594 ( .B1(n9682), .B2(n9593), .A(n7923), .ZN(P1_U3279) );
  AOI22_X1 U9595 ( .A1(n8788), .A2(n7924), .B1(n8755), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n7925) );
  OAI21_X1 U9596 ( .B1(n7926), .B2(n8066), .A(n7925), .ZN(P2_U3462) );
  AOI22_X1 U9597 ( .A1(n8788), .A2(n7927), .B1(n8755), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n7928) );
  OAI21_X1 U9598 ( .B1(n7929), .B2(n8066), .A(n7928), .ZN(P2_U3466) );
  NAND2_X1 U9599 ( .A1(n7930), .A2(n7931), .ZN(n7932) );
  XNOR2_X1 U9600 ( .A(n7932), .B(n8032), .ZN(n7968) );
  XNOR2_X1 U9601 ( .A(n7933), .B(n8032), .ZN(n7934) );
  OAI222_X1 U9602 ( .A1(n8669), .A2(n8024), .B1(n8711), .B2(n8097), .C1(n7934), 
        .C2(n8666), .ZN(n7970) );
  NAND2_X1 U9603 ( .A1(n7970), .A2(n10069), .ZN(n7938) );
  OAI22_X1 U9604 ( .A1(n8715), .A2(n7935), .B1(n8093), .B2(n10064), .ZN(n7936)
         );
  AOI21_X1 U9605 ( .B1(n8735), .B2(n7967), .A(n7936), .ZN(n7937) );
  OAI211_X1 U9606 ( .C1(n7968), .C2(n8738), .A(n7938), .B(n7937), .ZN(P2_U3222) );
  INV_X1 U9607 ( .A(n7939), .ZN(n7943) );
  OAI222_X1 U9608 ( .A1(n9732), .A2(n7943), .B1(P1_U3086), .B2(n7941), .C1(
        n7940), .C2(n9729), .ZN(P1_U3333) );
  INV_X1 U9609 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7942) );
  OAI222_X1 U9610 ( .A1(P2_U3151), .A2(n7944), .B1(n8878), .B2(n7943), .C1(
        n7942), .C2(n8880), .ZN(P2_U3273) );
  INV_X1 U9611 ( .A(n7949), .ZN(n7947) );
  NAND2_X1 U9612 ( .A1(n8876), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7945) );
  OAI211_X1 U9613 ( .C1(n7947), .C2(n8878), .A(n7946), .B(n7945), .ZN(P2_U3272) );
  NAND2_X1 U9614 ( .A1(n7949), .A2(n7948), .ZN(n7950) );
  OAI211_X1 U9615 ( .C1(n7951), .C2(n9729), .A(n7950), .B(n9273), .ZN(P1_U3332) );
  XNOR2_X1 U9616 ( .A(n8173), .B(n7954), .ZN(n8018) );
  XNOR2_X1 U9617 ( .A(n8018), .B(n7955), .ZN(n7956) );
  XNOR2_X1 U9618 ( .A(n8020), .B(n7956), .ZN(n7957) );
  NAND2_X1 U9619 ( .A1(n7957), .A2(n8321), .ZN(n7965) );
  INV_X1 U9620 ( .A(n7958), .ZN(n7962) );
  OAI22_X1 U9621 ( .A1(n8324), .A2(n7960), .B1(n7959), .B2(n8347), .ZN(n7961)
         );
  AOI211_X1 U9622 ( .C1(n7963), .C2(n8339), .A(n7962), .B(n7961), .ZN(n7964)
         );
  OAI211_X1 U9623 ( .C1(n7966), .C2(n8348), .A(n7965), .B(n7964), .ZN(P2_U3161) );
  INV_X1 U9624 ( .A(n7967), .ZN(n8098) );
  OAI22_X1 U9625 ( .A1(n7968), .A2(n8118), .B1(n8098), .B2(n8745), .ZN(n7969)
         );
  NOR2_X1 U9626 ( .A1(n7970), .A2(n7969), .ZN(n10086) );
  NAND2_X1 U9627 ( .A1(n8755), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7971) );
  OAI21_X1 U9628 ( .B1(n10086), .B2(n8755), .A(n7971), .ZN(P2_U3470) );
  XNOR2_X1 U9629 ( .A(n7972), .B(n7973), .ZN(n7998) );
  OAI211_X1 U9630 ( .C1(n7976), .C2(n7975), .A(n7974), .B(n8731), .ZN(n7978)
         );
  AOI22_X1 U9631 ( .A1(n8728), .A2(n8360), .B1(n8362), .B2(n8726), .ZN(n7977)
         );
  NAND2_X1 U9632 ( .A1(n7978), .A2(n7977), .ZN(n7999) );
  NAND2_X1 U9633 ( .A1(n7999), .A2(n10069), .ZN(n7982) );
  OAI22_X1 U9634 ( .A1(n8715), .A2(n7979), .B1(n8038), .B2(n10064), .ZN(n7980)
         );
  AOI21_X1 U9635 ( .B1(n8735), .B2(n8041), .A(n7980), .ZN(n7981) );
  OAI211_X1 U9636 ( .C1(n7998), .C2(n8738), .A(n7982), .B(n7981), .ZN(P2_U3221) );
  INV_X1 U9637 ( .A(n5956), .ZN(n8201) );
  OAI222_X1 U9638 ( .A1(n9732), .A2(n8201), .B1(P1_U3086), .B2(n7984), .C1(
        n7983), .C2(n9729), .ZN(P1_U3331) );
  AOI21_X1 U9639 ( .B1(n7986), .B2(n7985), .A(n4429), .ZN(n7994) );
  NAND2_X1 U9640 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9848) );
  NAND2_X1 U9641 ( .A1(n8999), .A2(n9587), .ZN(n7987) );
  OAI211_X1 U9642 ( .C1(n7988), .C2(n9001), .A(n9848), .B(n7987), .ZN(n7991)
         );
  NOR2_X1 U9643 ( .A1(n7989), .A2(n9008), .ZN(n7990) );
  AOI211_X1 U9644 ( .C1(n7992), .C2(n9004), .A(n7991), .B(n7990), .ZN(n7993)
         );
  OAI21_X1 U9645 ( .B1(n7994), .B2(n8974), .A(n7993), .ZN(P1_U3215) );
  INV_X1 U9646 ( .A(n7995), .ZN(n8128) );
  OAI222_X1 U9647 ( .A1(n9732), .A2(n8128), .B1(P1_U3086), .B2(n7997), .C1(
        n7996), .C2(n9729), .ZN(P1_U3330) );
  NOR2_X1 U9648 ( .A1(n7998), .A2(n8118), .ZN(n8000) );
  AOI211_X1 U9649 ( .C1(n8793), .C2(n8041), .A(n8000), .B(n7999), .ZN(n10089)
         );
  NAND2_X1 U9650 ( .A1(n8755), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n8001) );
  OAI21_X1 U9651 ( .B1(n10089), .B2(n8755), .A(n8001), .ZN(P2_U3471) );
  INV_X1 U9652 ( .A(n10061), .ZN(n8615) );
  XNOR2_X1 U9653 ( .A(n8002), .B(n8004), .ZN(n8003) );
  OAI222_X1 U9654 ( .A1(n8711), .A2(n8150), .B1(n8669), .B2(n8097), .C1(n8666), 
        .C2(n8003), .ZN(n8062) );
  AOI21_X1 U9655 ( .B1(n8615), .B2(n8077), .A(n8062), .ZN(n8008) );
  XNOR2_X1 U9656 ( .A(n8005), .B(n8004), .ZN(n8064) );
  OAI22_X1 U9657 ( .A1(n8715), .A2(n8377), .B1(n8079), .B2(n10064), .ZN(n8006)
         );
  AOI21_X1 U9658 ( .B1(n8064), .B2(n8596), .A(n8006), .ZN(n8007) );
  OAI21_X1 U9659 ( .B1(n8008), .B2(n8734), .A(n8007), .ZN(P2_U3220) );
  XOR2_X1 U9660 ( .A(n9036), .B(n8009), .Z(n9676) );
  AOI211_X1 U9661 ( .C1(n9672), .C2(n8010), .A(n9590), .B(n9588), .ZN(n9671)
         );
  AOI22_X1 U9662 ( .A1(n9593), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9005), .B2(
        n9952), .ZN(n8011) );
  OAI21_X1 U9663 ( .B1(n9009), .B2(n9955), .A(n8011), .ZN(n8016) );
  OAI21_X1 U9664 ( .B1(n9036), .B2(n8013), .A(n8012), .ZN(n8014) );
  AOI222_X1 U9665 ( .A1(n9906), .A2(n8014), .B1(n9575), .B2(n7513), .C1(n9277), 
        .C2(n9932), .ZN(n9674) );
  NOR2_X1 U9666 ( .A1(n9674), .A2(n9593), .ZN(n8015) );
  AOI211_X1 U9667 ( .C1(n9671), .C2(n9949), .A(n8016), .B(n8015), .ZN(n8017)
         );
  OAI21_X1 U9668 ( .B1(n9676), .B2(n9601), .A(n8017), .ZN(P1_U3278) );
  NAND2_X1 U9669 ( .A1(n8018), .A2(n8365), .ZN(n8019) );
  XNOR2_X1 U9670 ( .A(n8173), .B(n8296), .ZN(n8021) );
  XNOR2_X1 U9671 ( .A(n8021), .B(n8364), .ZN(n8292) );
  INV_X1 U9672 ( .A(n8021), .ZN(n8022) );
  NAND2_X1 U9673 ( .A1(n8022), .A2(n8364), .ZN(n8023) );
  NAND2_X1 U9674 ( .A1(n8291), .A2(n8023), .ZN(n8088) );
  XOR2_X1 U9675 ( .A(n8163), .B(n8032), .Z(n8092) );
  XNOR2_X1 U9676 ( .A(n8173), .B(n8053), .ZN(n8089) );
  INV_X1 U9677 ( .A(n8089), .ZN(n8025) );
  AND2_X1 U9678 ( .A1(n8092), .A2(n8026), .ZN(n8027) );
  NAND2_X1 U9679 ( .A1(n8088), .A2(n8027), .ZN(n8035) );
  MUX2_X1 U9680 ( .A(n8362), .B(n8028), .S(n8163), .Z(n8033) );
  NAND2_X1 U9681 ( .A1(n8163), .A2(n8362), .ZN(n8029) );
  OAI211_X1 U9682 ( .C1(n8163), .C2(n8030), .A(n8032), .B(n8029), .ZN(n8031)
         );
  OAI21_X1 U9683 ( .B1(n8033), .B2(n8032), .A(n8031), .ZN(n8034) );
  NAND2_X1 U9684 ( .A1(n8035), .A2(n8034), .ZN(n8036) );
  XNOR2_X1 U9685 ( .A(n8041), .B(n8163), .ZN(n8073) );
  XNOR2_X1 U9686 ( .A(n8073), .B(n8361), .ZN(n8037) );
  NAND2_X1 U9687 ( .A1(n8036), .A2(n8037), .ZN(n8076) );
  OAI211_X1 U9688 ( .C1(n8036), .C2(n8037), .A(n8076), .B(n8321), .ZN(n8047)
         );
  INV_X1 U9689 ( .A(n8038), .ZN(n8045) );
  NAND2_X1 U9690 ( .A1(n8351), .A2(n8362), .ZN(n8040) );
  OAI211_X1 U9691 ( .C1(n8144), .C2(n8347), .A(n8040), .B(n8039), .ZN(n8044)
         );
  INV_X1 U9692 ( .A(n8041), .ZN(n8042) );
  NOR2_X1 U9693 ( .A1(n8354), .A2(n8042), .ZN(n8043) );
  AOI211_X1 U9694 ( .C1(n8045), .C2(n8335), .A(n8044), .B(n8043), .ZN(n8046)
         );
  NAND2_X1 U9695 ( .A1(n8047), .A2(n8046), .ZN(P2_U3164) );
  XNOR2_X1 U9696 ( .A(n8088), .B(n8363), .ZN(n8090) );
  XOR2_X1 U9697 ( .A(n8089), .B(n8090), .Z(n8058) );
  INV_X1 U9698 ( .A(n8048), .ZN(n8056) );
  NAND2_X1 U9699 ( .A1(n8351), .A2(n8364), .ZN(n8051) );
  INV_X1 U9700 ( .A(n8049), .ZN(n8050) );
  OAI211_X1 U9701 ( .C1(n8052), .C2(n8347), .A(n8051), .B(n8050), .ZN(n8055)
         );
  NOR2_X1 U9702 ( .A1(n8354), .A2(n8053), .ZN(n8054) );
  AOI211_X1 U9703 ( .C1(n8056), .C2(n8335), .A(n8055), .B(n8054), .ZN(n8057)
         );
  OAI21_X1 U9704 ( .B1(n8058), .B2(n8342), .A(n8057), .ZN(P2_U3157) );
  INV_X1 U9705 ( .A(n8059), .ZN(n8068) );
  OAI222_X1 U9706 ( .A1(n9727), .A2(n8068), .B1(P1_U3086), .B2(n8061), .C1(
        n8060), .C2(n9729), .ZN(P1_U3329) );
  NOR2_X1 U9707 ( .A1(n8082), .A2(n8745), .ZN(n8063) );
  AOI211_X1 U9708 ( .C1(n8064), .C2(n8794), .A(n8063), .B(n8062), .ZN(n9784)
         );
  NAND2_X1 U9709 ( .A1(n8755), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8065) );
  OAI21_X1 U9710 ( .B1(n9784), .B2(n8066), .A(n8065), .ZN(P2_U3472) );
  INV_X1 U9711 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8067) );
  OAI222_X1 U9712 ( .A1(n8069), .A2(P2_U3151), .B1(n8878), .B2(n8068), .C1(
        n8067), .C2(n8880), .ZN(P2_U3269) );
  INV_X1 U9713 ( .A(n8070), .ZN(n8109) );
  AOI21_X1 U9714 ( .B1(n8876), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n8071), .ZN(
        n8072) );
  OAI21_X1 U9715 ( .B1(n8109), .B2(n8878), .A(n8072), .ZN(P2_U3268) );
  INV_X1 U9716 ( .A(n8073), .ZN(n8074) );
  NAND2_X1 U9717 ( .A1(n8074), .A2(n8361), .ZN(n8075) );
  XNOR2_X1 U9718 ( .A(n8077), .B(n8163), .ZN(n8146) );
  XNOR2_X1 U9719 ( .A(n8146), .B(n8360), .ZN(n8078) );
  XNOR2_X1 U9720 ( .A(n8145), .B(n8078), .ZN(n8087) );
  INV_X1 U9721 ( .A(n8079), .ZN(n8085) );
  NAND2_X1 U9722 ( .A1(n8351), .A2(n8361), .ZN(n8081) );
  OR2_X1 U9723 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8080), .ZN(n8391) );
  OAI211_X1 U9724 ( .C1(n8150), .C2(n8347), .A(n8081), .B(n8391), .ZN(n8084)
         );
  NOR2_X1 U9725 ( .A1(n8354), .A2(n8082), .ZN(n8083) );
  AOI211_X1 U9726 ( .C1(n8085), .C2(n8335), .A(n8084), .B(n8083), .ZN(n8086)
         );
  OAI21_X1 U9727 ( .B1(n8087), .B2(n8342), .A(n8086), .ZN(P2_U3174) );
  OAI22_X1 U9728 ( .A1(n8090), .A2(n8089), .B1(n8363), .B2(n8088), .ZN(n8091)
         );
  XOR2_X1 U9729 ( .A(n8092), .B(n8091), .Z(n8103) );
  INV_X1 U9730 ( .A(n8093), .ZN(n8101) );
  NAND2_X1 U9731 ( .A1(n8351), .A2(n8363), .ZN(n8096) );
  INV_X1 U9732 ( .A(n8094), .ZN(n8095) );
  OAI211_X1 U9733 ( .C1(n8097), .C2(n8347), .A(n8096), .B(n8095), .ZN(n8100)
         );
  NOR2_X1 U9734 ( .A1(n8354), .A2(n8098), .ZN(n8099) );
  AOI211_X1 U9735 ( .C1(n8101), .C2(n8335), .A(n8100), .B(n8099), .ZN(n8102)
         );
  OAI21_X1 U9736 ( .B1(n8103), .B2(n8342), .A(n8102), .ZN(P2_U3176) );
  INV_X1 U9737 ( .A(n8104), .ZN(n8143) );
  NAND2_X1 U9738 ( .A1(n8876), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8105) );
  OAI211_X1 U9739 ( .C1(n8143), .C2(n8878), .A(n8106), .B(n8105), .ZN(P2_U3267) );
  OAI222_X1 U9740 ( .A1(n9727), .A2(n8109), .B1(P1_U3086), .B2(n8108), .C1(
        n8107), .C2(n9729), .ZN(P1_U3328) );
  XNOR2_X1 U9741 ( .A(n8110), .B(n8111), .ZN(n8126) );
  INV_X1 U9742 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8115) );
  XNOR2_X1 U9743 ( .A(n8112), .B(n8113), .ZN(n8114) );
  AOI222_X1 U9744 ( .A1(n8731), .A2(n8114), .B1(n8709), .B2(n8728), .C1(n8360), 
        .C2(n8726), .ZN(n8121) );
  MUX2_X1 U9745 ( .A(n8115), .B(n8121), .S(n10088), .Z(n8117) );
  NAND2_X1 U9746 ( .A1(n8866), .A2(n8149), .ZN(n8116) );
  OAI211_X1 U9747 ( .C1(n8126), .C2(n8870), .A(n8117), .B(n8116), .ZN(P2_U3432) );
  MUX2_X1 U9748 ( .A(n8409), .B(n8121), .S(n8786), .Z(n8120) );
  NAND2_X1 U9749 ( .A1(n8149), .A2(n8788), .ZN(n8119) );
  OAI211_X1 U9750 ( .C1(n8791), .C2(n8126), .A(n8120), .B(n8119), .ZN(P2_U3473) );
  INV_X1 U9751 ( .A(n8121), .ZN(n8123) );
  INV_X1 U9752 ( .A(n8149), .ZN(n8218) );
  OAI22_X1 U9753 ( .A1(n8218), .A2(n10061), .B1(n8215), .B2(n10064), .ZN(n8122) );
  OAI21_X1 U9754 ( .B1(n8123), .B2(n8122), .A(n8715), .ZN(n8125) );
  NAND2_X1 U9755 ( .A1(n8734), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8124) );
  OAI211_X1 U9756 ( .C1(n8126), .C2(n8738), .A(n8125), .B(n8124), .ZN(P2_U3219) );
  INV_X1 U9757 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8127) );
  OAI222_X1 U9758 ( .A1(n8129), .A2(P2_U3151), .B1(n8878), .B2(n8128), .C1(
        n8127), .C2(n8880), .ZN(P2_U3270) );
  INV_X1 U9759 ( .A(n9010), .ZN(n8204) );
  OAI222_X1 U9760 ( .A1(n9729), .A2(n9011), .B1(n9727), .B2(n8204), .C1(
        P1_U3086), .C2(n8130), .ZN(P1_U3325) );
  NAND2_X1 U9761 ( .A1(n9952), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n8132) );
  INV_X1 U9762 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n8131) );
  OAI22_X1 U9763 ( .A1(n8133), .A2(n8132), .B1(n8131), .B2(n9598), .ZN(n8134)
         );
  AOI21_X1 U9764 ( .B1(n8135), .B2(n9939), .A(n8134), .ZN(n8136) );
  OAI21_X1 U9765 ( .B1(n8137), .B2(n9405), .A(n8136), .ZN(n8138) );
  AOI21_X1 U9766 ( .B1(n8139), .B2(n9959), .A(n8138), .ZN(n8140) );
  OAI21_X1 U9767 ( .B1(n8141), .B2(n9593), .A(n8140), .ZN(P1_U3356) );
  OAI222_X1 U9768 ( .A1(n9727), .A2(n8143), .B1(P1_U3086), .B2(n4351), .C1(
        n8142), .C2(n9729), .ZN(P1_U3327) );
  XNOR2_X1 U9769 ( .A(n8773), .B(n8163), .ZN(n8170) );
  XOR2_X1 U9770 ( .A(n8678), .B(n8170), .Z(n8302) );
  XNOR2_X1 U9771 ( .A(n8836), .B(n8163), .ZN(n8172) );
  XNOR2_X1 U9772 ( .A(n8172), .B(n8640), .ZN(n8243) );
  INV_X1 U9773 ( .A(n8243), .ZN(n8171) );
  OR2_X1 U9774 ( .A1(n8302), .A2(n8171), .ZN(n8169) );
  INV_X1 U9775 ( .A(n8146), .ZN(n8147) );
  NAND2_X1 U9776 ( .A1(n8147), .A2(n8360), .ZN(n8148) );
  XNOR2_X1 U9777 ( .A(n8149), .B(n8163), .ZN(n8151) );
  XOR2_X1 U9778 ( .A(n8727), .B(n8151), .Z(n8214) );
  XNOR2_X1 U9779 ( .A(n8792), .B(n8163), .ZN(n8157) );
  XOR2_X1 U9780 ( .A(n8709), .B(n8157), .Z(n8343) );
  XNOR2_X1 U9781 ( .A(n8860), .B(n8163), .ZN(n8152) );
  NAND2_X1 U9782 ( .A1(n8152), .A2(n8712), .ZN(n8316) );
  INV_X1 U9783 ( .A(n8152), .ZN(n8153) );
  NAND2_X1 U9784 ( .A1(n8153), .A2(n8688), .ZN(n8154) );
  INV_X1 U9785 ( .A(n8273), .ZN(n8155) );
  XNOR2_X1 U9786 ( .A(n8867), .B(n8163), .ZN(n8156) );
  NAND2_X1 U9787 ( .A1(n8156), .A2(n8346), .ZN(n8272) );
  NOR2_X1 U9788 ( .A1(n8155), .A2(n8272), .ZN(n8160) );
  OR2_X1 U9789 ( .A1(n8343), .A2(n8160), .ZN(n8162) );
  OAI21_X1 U9790 ( .B1(n8156), .B2(n8346), .A(n8272), .ZN(n8263) );
  INV_X1 U9791 ( .A(n8157), .ZN(n8158) );
  AND2_X1 U9792 ( .A1(n8158), .A2(n8709), .ZN(n8262) );
  NOR2_X1 U9793 ( .A1(n8263), .A2(n8262), .ZN(n8261) );
  AND2_X1 U9794 ( .A1(n8261), .A2(n8273), .ZN(n8159) );
  OR2_X1 U9795 ( .A1(n8160), .A2(n8159), .ZN(n8161) );
  OAI21_X1 U9796 ( .B1(n8260), .B2(n8162), .A(n8161), .ZN(n8276) );
  NAND2_X1 U9797 ( .A1(n8276), .A2(n8316), .ZN(n8164) );
  XNOR2_X1 U9798 ( .A(n8854), .B(n8163), .ZN(n8165) );
  XNOR2_X1 U9799 ( .A(n8165), .B(n8698), .ZN(n8317) );
  NAND2_X1 U9800 ( .A1(n8164), .A2(n8317), .ZN(n8320) );
  NAND2_X1 U9801 ( .A1(n8165), .A2(n8278), .ZN(n8166) );
  NAND2_X1 U9802 ( .A1(n8320), .A2(n8166), .ZN(n8234) );
  XNOR2_X1 U9803 ( .A(n8848), .B(n7358), .ZN(n8167) );
  NOR2_X1 U9804 ( .A1(n8167), .A2(n8689), .ZN(n8230) );
  NAND2_X1 U9805 ( .A1(n8167), .A2(n8689), .ZN(n8231) );
  NAND2_X1 U9806 ( .A1(n8170), .A2(n8246), .ZN(n8240) );
  XOR2_X1 U9807 ( .A(n8173), .B(n8830), .Z(n8175) );
  INV_X1 U9808 ( .A(n8175), .ZN(n8174) );
  XNOR2_X1 U9809 ( .A(n8174), .B(n8655), .ZN(n8309) );
  NOR2_X1 U9810 ( .A1(n8175), .A2(n8655), .ZN(n8176) );
  AOI21_X2 U9811 ( .B1(n8308), .B2(n8309), .A(n8176), .ZN(n8177) );
  XNOR2_X1 U9812 ( .A(n8824), .B(n8163), .ZN(n8178) );
  NAND2_X1 U9813 ( .A1(n8224), .A2(n8312), .ZN(n8181) );
  INV_X1 U9814 ( .A(n8177), .ZN(n8179) );
  NAND2_X1 U9815 ( .A1(n8179), .A2(n8178), .ZN(n8180) );
  NAND2_X1 U9816 ( .A1(n8181), .A2(n8180), .ZN(n8284) );
  XNOR2_X1 U9817 ( .A(n8818), .B(n8163), .ZN(n8182) );
  XNOR2_X1 U9818 ( .A(n8182), .B(n8628), .ZN(n8285) );
  NAND2_X1 U9819 ( .A1(n8284), .A2(n8285), .ZN(n8184) );
  NAND2_X1 U9820 ( .A1(n8182), .A2(n8253), .ZN(n8183) );
  XNOR2_X1 U9821 ( .A(n8256), .B(n8163), .ZN(n8185) );
  XNOR2_X1 U9822 ( .A(n8185), .B(n8612), .ZN(n8251) );
  NAND2_X1 U9823 ( .A1(n8250), .A2(n8251), .ZN(n8187) );
  NAND2_X1 U9824 ( .A1(n8185), .A2(n8588), .ZN(n8186) );
  XNOR2_X1 U9825 ( .A(n5542), .B(n7358), .ZN(n8188) );
  NAND2_X1 U9826 ( .A1(n8188), .A2(n8604), .ZN(n8331) );
  INV_X1 U9827 ( .A(n8188), .ZN(n8189) );
  NAND2_X1 U9828 ( .A1(n8189), .A2(n8578), .ZN(n8332) );
  XNOR2_X1 U9829 ( .A(n8210), .B(n8163), .ZN(n8190) );
  XOR2_X1 U9830 ( .A(n8358), .B(n8190), .Z(n8205) );
  XNOR2_X1 U9831 ( .A(n8191), .B(n8163), .ZN(n8192) );
  XNOR2_X1 U9832 ( .A(n8193), .B(n8192), .ZN(n8199) );
  AOI22_X1 U9833 ( .A1(n8358), .A2(n8351), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8195) );
  NAND2_X1 U9834 ( .A1(n8335), .A2(n8570), .ZN(n8194) );
  OAI211_X1 U9835 ( .C1(n8563), .C2(n8347), .A(n8195), .B(n8194), .ZN(n8196)
         );
  AOI21_X1 U9836 ( .B1(n8197), .B2(n8339), .A(n8196), .ZN(n8198) );
  OAI21_X1 U9837 ( .B1(n8199), .B2(n8342), .A(n8198), .ZN(P2_U3160) );
  INV_X1 U9838 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8200) );
  OAI222_X1 U9839 ( .A1(n8202), .A2(P2_U3151), .B1(n8878), .B2(n8201), .C1(
        n8200), .C2(n8880), .ZN(P2_U3271) );
  OAI222_X1 U9840 ( .A1(n5048), .A2(P2_U3151), .B1(n8878), .B2(n8204), .C1(
        n8203), .C2(n8880), .ZN(P2_U3265) );
  XNOR2_X1 U9841 ( .A(n8206), .B(n8205), .ZN(n8212) );
  AOI22_X1 U9842 ( .A1(n8351), .A2(n8604), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8208) );
  NAND2_X1 U9843 ( .A1(n8335), .A2(n8581), .ZN(n8207) );
  OAI211_X1 U9844 ( .C1(n8577), .C2(n8347), .A(n8208), .B(n8207), .ZN(n8209)
         );
  AOI21_X1 U9845 ( .B1(n8210), .B2(n8339), .A(n8209), .ZN(n8211) );
  OAI21_X1 U9846 ( .B1(n8212), .B2(n8342), .A(n8211), .ZN(P2_U3154) );
  AOI21_X1 U9847 ( .B1(n8214), .B2(n8213), .A(n4428), .ZN(n8223) );
  INV_X1 U9848 ( .A(n8215), .ZN(n8221) );
  NAND2_X1 U9849 ( .A1(n8351), .A2(n8360), .ZN(n8216) );
  NAND2_X1 U9850 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8418) );
  OAI211_X1 U9851 ( .C1(n8217), .C2(n8347), .A(n8216), .B(n8418), .ZN(n8220)
         );
  NOR2_X1 U9852 ( .A1(n8218), .A2(n8354), .ZN(n8219) );
  AOI211_X1 U9853 ( .C1(n8221), .C2(n8335), .A(n8220), .B(n8219), .ZN(n8222)
         );
  OAI21_X1 U9854 ( .B1(n8223), .B2(n8342), .A(n8222), .ZN(P2_U3155) );
  XNOR2_X1 U9855 ( .A(n8224), .B(n8641), .ZN(n8229) );
  AOI22_X1 U9856 ( .A1(n8351), .A2(n8655), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8226) );
  NAND2_X1 U9857 ( .A1(n8335), .A2(n8631), .ZN(n8225) );
  OAI211_X1 U9858 ( .C1(n8253), .C2(n8347), .A(n8226), .B(n8225), .ZN(n8227)
         );
  AOI21_X1 U9859 ( .B1(n8824), .B2(n8339), .A(n8227), .ZN(n8228) );
  OAI21_X1 U9860 ( .B1(n8229), .B2(n8342), .A(n8228), .ZN(P2_U3156) );
  INV_X1 U9861 ( .A(n8230), .ZN(n8232) );
  NAND2_X1 U9862 ( .A1(n8232), .A2(n8231), .ZN(n8233) );
  XNOR2_X1 U9863 ( .A(n8234), .B(n8233), .ZN(n8239) );
  AND2_X1 U9864 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8538) );
  NOR2_X1 U9865 ( .A1(n8347), .A2(n8246), .ZN(n8235) );
  AOI211_X1 U9866 ( .C1(n8351), .C2(n8698), .A(n8538), .B(n8235), .ZN(n8236)
         );
  OAI21_X1 U9867 ( .B1(n8681), .B2(n8348), .A(n8236), .ZN(n8237) );
  AOI21_X1 U9868 ( .B1(n8848), .B2(n8339), .A(n8237), .ZN(n8238) );
  OAI21_X1 U9869 ( .B1(n8239), .B2(n8342), .A(n8238), .ZN(P2_U3159) );
  OR2_X1 U9870 ( .A1(n8301), .A2(n8302), .ZN(n8241) );
  NAND2_X1 U9871 ( .A1(n8241), .A2(n8240), .ZN(n8242) );
  XOR2_X1 U9872 ( .A(n8243), .B(n8242), .Z(n8249) );
  AOI22_X1 U9873 ( .A1(n8327), .A2(n8655), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8245) );
  NAND2_X1 U9874 ( .A1(n8335), .A2(n8658), .ZN(n8244) );
  OAI211_X1 U9875 ( .C1(n8246), .C2(n8324), .A(n8245), .B(n8244), .ZN(n8247)
         );
  AOI21_X1 U9876 ( .B1(n8836), .B2(n8339), .A(n8247), .ZN(n8248) );
  OAI21_X1 U9877 ( .B1(n8249), .B2(n8342), .A(n8248), .ZN(P2_U3163) );
  XOR2_X1 U9878 ( .A(n8251), .B(n8250), .Z(n8259) );
  OAI22_X1 U9879 ( .A1(n8578), .A2(n8347), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8252), .ZN(n8255) );
  NOR2_X1 U9880 ( .A1(n8324), .A2(n8253), .ZN(n8254) );
  AOI211_X1 U9881 ( .C1(n8608), .C2(n8335), .A(n8255), .B(n8254), .ZN(n8258)
         );
  NAND2_X1 U9882 ( .A1(n8256), .A2(n8339), .ZN(n8257) );
  OAI211_X1 U9883 ( .C1(n8259), .C2(n8342), .A(n8258), .B(n8257), .ZN(P2_U3165) );
  INV_X1 U9884 ( .A(n8867), .ZN(n8271) );
  INV_X1 U9885 ( .A(n8262), .ZN(n8265) );
  INV_X1 U9886 ( .A(n8263), .ZN(n8264) );
  AOI21_X1 U9887 ( .B1(n8344), .B2(n8265), .A(n8264), .ZN(n8266) );
  OAI21_X1 U9888 ( .B1(n8275), .B2(n8266), .A(n8321), .ZN(n8270) );
  NAND2_X1 U9889 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8455) );
  OAI21_X1 U9890 ( .B1(n8347), .B2(n8712), .A(n8455), .ZN(n8268) );
  NOR2_X1 U9891 ( .A1(n8348), .A2(n8717), .ZN(n8267) );
  AOI211_X1 U9892 ( .C1(n8351), .C2(n8709), .A(n8268), .B(n8267), .ZN(n8269)
         );
  OAI211_X1 U9893 ( .C1(n8271), .C2(n8354), .A(n8270), .B(n8269), .ZN(P2_U3166) );
  INV_X1 U9894 ( .A(n8860), .ZN(n8283) );
  INV_X1 U9895 ( .A(n8272), .ZN(n8274) );
  NOR3_X1 U9896 ( .A1(n8275), .A2(n8274), .A3(n8273), .ZN(n8277) );
  INV_X1 U9897 ( .A(n8276), .ZN(n8319) );
  OAI21_X1 U9898 ( .B1(n8277), .B2(n8319), .A(n8321), .ZN(n8282) );
  NAND2_X1 U9899 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8484) );
  OAI21_X1 U9900 ( .B1(n8347), .B2(n8278), .A(n8484), .ZN(n8280) );
  NOR2_X1 U9901 ( .A1(n8348), .A2(n8701), .ZN(n8279) );
  AOI211_X1 U9902 ( .C1(n8351), .C2(n8729), .A(n8280), .B(n8279), .ZN(n8281)
         );
  OAI211_X1 U9903 ( .C1(n8283), .C2(n8354), .A(n8282), .B(n8281), .ZN(P2_U3168) );
  XOR2_X1 U9904 ( .A(n8285), .B(n8284), .Z(n8290) );
  AOI22_X1 U9905 ( .A1(n8327), .A2(n8612), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8287) );
  NAND2_X1 U9906 ( .A1(n8335), .A2(n8614), .ZN(n8286) );
  OAI211_X1 U9907 ( .C1(n8312), .C2(n8324), .A(n8287), .B(n8286), .ZN(n8288)
         );
  AOI21_X1 U9908 ( .B1(n8818), .B2(n8339), .A(n8288), .ZN(n8289) );
  OAI21_X1 U9909 ( .B1(n8290), .B2(n8342), .A(n8289), .ZN(P2_U3169) );
  OAI211_X1 U9910 ( .C1(n4442), .C2(n8292), .A(n8291), .B(n8321), .ZN(n8300)
         );
  NOR2_X1 U9911 ( .A1(n8347), .A2(n8024), .ZN(n8293) );
  AOI211_X1 U9912 ( .C1(n8351), .C2(n8365), .A(n8294), .B(n8293), .ZN(n8299)
         );
  INV_X1 U9913 ( .A(n8295), .ZN(n8297) );
  AOI22_X1 U9914 ( .A1(n8297), .A2(n8335), .B1(n8339), .B2(n8296), .ZN(n8298)
         );
  NAND3_X1 U9915 ( .A1(n8300), .A2(n8299), .A3(n8298), .ZN(P2_U3171) );
  XOR2_X1 U9916 ( .A(n8302), .B(n8301), .Z(n8307) );
  AOI22_X1 U9917 ( .A1(n8327), .A2(n8640), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8304) );
  NAND2_X1 U9918 ( .A1(n8335), .A2(n8672), .ZN(n8303) );
  OAI211_X1 U9919 ( .C1(n8668), .C2(n8324), .A(n8304), .B(n8303), .ZN(n8305)
         );
  AOI21_X1 U9920 ( .B1(n8773), .B2(n8339), .A(n8305), .ZN(n8306) );
  OAI21_X1 U9921 ( .B1(n8307), .B2(n8342), .A(n8306), .ZN(P2_U3173) );
  XOR2_X1 U9922 ( .A(n8309), .B(n8308), .Z(n8315) );
  AOI22_X1 U9923 ( .A1(n8351), .A2(n8640), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8311) );
  NAND2_X1 U9924 ( .A1(n8335), .A2(n8644), .ZN(n8310) );
  OAI211_X1 U9925 ( .C1(n8312), .C2(n8347), .A(n8311), .B(n8310), .ZN(n8313)
         );
  AOI21_X1 U9926 ( .B1(n8830), .B2(n8339), .A(n8313), .ZN(n8314) );
  OAI21_X1 U9927 ( .B1(n8315), .B2(n8342), .A(n8314), .ZN(P2_U3175) );
  INV_X1 U9928 ( .A(n8854), .ZN(n8330) );
  INV_X1 U9929 ( .A(n8316), .ZN(n8318) );
  NOR3_X1 U9930 ( .A1(n8319), .A2(n8318), .A3(n8317), .ZN(n8323) );
  INV_X1 U9931 ( .A(n8320), .ZN(n8322) );
  OAI21_X1 U9932 ( .B1(n8323), .B2(n8322), .A(n8321), .ZN(n8329) );
  NOR2_X1 U9933 ( .A1(n8348), .A2(n8692), .ZN(n8326) );
  NAND2_X1 U9934 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8516) );
  OAI21_X1 U9935 ( .B1(n8324), .B2(n8712), .A(n8516), .ZN(n8325) );
  AOI211_X1 U9936 ( .C1(n8327), .C2(n8689), .A(n8326), .B(n8325), .ZN(n8328)
         );
  OAI211_X1 U9937 ( .C1(n8330), .C2(n8354), .A(n8329), .B(n8328), .ZN(P2_U3178) );
  NAND2_X1 U9938 ( .A1(n8332), .A2(n8331), .ZN(n8333) );
  XNOR2_X1 U9939 ( .A(n8334), .B(n8333), .ZN(n8341) );
  AOI22_X1 U9940 ( .A1(n8351), .A2(n8612), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8337) );
  NAND2_X1 U9941 ( .A1(n8335), .A2(n8590), .ZN(n8336) );
  OAI211_X1 U9942 ( .C1(n8589), .C2(n8347), .A(n8337), .B(n8336), .ZN(n8338)
         );
  AOI21_X1 U9943 ( .B1(n5542), .B2(n8339), .A(n8338), .ZN(n8340) );
  OAI21_X1 U9944 ( .B1(n8341), .B2(n8342), .A(n8340), .ZN(P2_U3180) );
  AOI21_X1 U9945 ( .B1(n8260), .B2(n8343), .A(n8342), .ZN(n8345) );
  NAND2_X1 U9946 ( .A1(n8345), .A2(n8344), .ZN(n8353) );
  NAND2_X1 U9947 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8438) );
  OAI21_X1 U9948 ( .B1(n8347), .B2(n8346), .A(n8438), .ZN(n8350) );
  NOR2_X1 U9949 ( .A1(n8348), .A2(n8732), .ZN(n8349) );
  AOI211_X1 U9950 ( .C1(n8351), .C2(n8727), .A(n8350), .B(n8349), .ZN(n8352)
         );
  OAI211_X1 U9951 ( .C1(n8355), .C2(n8354), .A(n8353), .B(n8352), .ZN(P2_U3181) );
  MUX2_X1 U9952 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8356), .S(n8512), .Z(
        P2_U3521) );
  MUX2_X1 U9953 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8357), .S(n8512), .Z(
        P2_U3519) );
  MUX2_X1 U9954 ( .A(n8358), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8359), .Z(
        P2_U3518) );
  MUX2_X1 U9955 ( .A(n8604), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8359), .Z(
        P2_U3517) );
  MUX2_X1 U9956 ( .A(n8612), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8359), .Z(
        P2_U3516) );
  MUX2_X1 U9957 ( .A(n8628), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8359), .Z(
        P2_U3515) );
  MUX2_X1 U9958 ( .A(n8641), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8359), .Z(
        P2_U3514) );
  MUX2_X1 U9959 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8655), .S(n8512), .Z(
        P2_U3513) );
  MUX2_X1 U9960 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8640), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9961 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8678), .S(n8512), .Z(
        P2_U3511) );
  MUX2_X1 U9962 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8689), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9963 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8698), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U9964 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8688), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9965 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8729), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9966 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8709), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U9967 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8727), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U9968 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8360), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U9969 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8361), .S(P2_U3893), .Z(
        P2_U3503) );
  MUX2_X1 U9970 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8362), .S(n8512), .Z(
        P2_U3502) );
  MUX2_X1 U9971 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8363), .S(n8512), .Z(
        P2_U3501) );
  MUX2_X1 U9972 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8364), .S(n8512), .Z(
        P2_U3500) );
  MUX2_X1 U9973 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8365), .S(n8512), .Z(
        P2_U3499) );
  MUX2_X1 U9974 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8366), .S(n8512), .Z(
        P2_U3498) );
  MUX2_X1 U9975 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8367), .S(n8512), .Z(
        P2_U3497) );
  MUX2_X1 U9976 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8368), .S(n8512), .Z(
        P2_U3496) );
  MUX2_X1 U9977 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8369), .S(n8512), .Z(
        P2_U3495) );
  MUX2_X1 U9978 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8370), .S(n8512), .Z(
        P2_U3494) );
  MUX2_X1 U9979 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n5101), .S(n8512), .Z(
        P2_U3493) );
  MUX2_X1 U9980 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n8371), .S(n8512), .Z(
        P2_U3492) );
  MUX2_X1 U9981 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n7046), .S(n8512), .Z(
        P2_U3491) );
  INV_X1 U9982 ( .A(n8372), .ZN(n8373) );
  MUX2_X1 U9983 ( .A(n8377), .B(n8376), .S(n8529), .Z(n8379) );
  AND2_X1 U9984 ( .A1(n8379), .A2(n8403), .ZN(n8414) );
  INV_X1 U9985 ( .A(n8414), .ZN(n8378) );
  OAI21_X1 U9986 ( .B1(n8403), .B2(n8379), .A(n8378), .ZN(n8380) );
  NOR2_X1 U9987 ( .A1(n8381), .A2(n8380), .ZN(n8413) );
  AOI21_X1 U9988 ( .B1(n8381), .B2(n8380), .A(n8413), .ZN(n8386) );
  NOR2_X1 U9989 ( .A1(n8384), .A2(n8376), .ZN(n8398) );
  AOI21_X1 U9990 ( .B1(n8376), .B2(n8384), .A(n8398), .ZN(n8385) );
  OAI22_X1 U9991 ( .A1(n8386), .A2(n8542), .B1(n8385), .B2(n10032), .ZN(n8395)
         );
  AOI21_X1 U9992 ( .B1(n8377), .B2(n8390), .A(n8404), .ZN(n8393) );
  AOI22_X1 U9993 ( .A1(n10047), .A2(n8403), .B1(n10045), .B2(
        P2_ADDR_REG_13__SCAN_IN), .ZN(n8392) );
  OAI211_X1 U9994 ( .C1(n8393), .C2(n8486), .A(n8392), .B(n8391), .ZN(n8394)
         );
  OR2_X1 U9995 ( .A1(n8395), .A2(n8394), .ZN(P2_U3195) );
  NOR2_X1 U9996 ( .A1(n8403), .A2(n8397), .ZN(n8399) );
  AOI22_X1 U9997 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8417), .B1(n8427), .B2(
        n8409), .ZN(n8400) );
  AOI21_X1 U9998 ( .B1(n8401), .B2(n8400), .A(n4427), .ZN(n8424) );
  NOR2_X1 U9999 ( .A1(n8403), .A2(n8402), .ZN(n8405) );
  AOI22_X1 U10000 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8417), .B1(n8427), .B2(
        n8410), .ZN(n8406) );
  AOI21_X1 U10001 ( .B1(n8407), .B2(n8406), .A(n8426), .ZN(n8408) );
  NOR2_X1 U10002 ( .A1(n8408), .A2(n8486), .ZN(n8422) );
  MUX2_X1 U10003 ( .A(n8410), .B(n8409), .S(n8529), .Z(n8412) );
  AND2_X1 U10004 ( .A1(n8412), .A2(n8417), .ZN(n8435) );
  INV_X1 U10005 ( .A(n8435), .ZN(n8411) );
  OAI21_X1 U10006 ( .B1(n8417), .B2(n8412), .A(n8411), .ZN(n8416) );
  NOR2_X1 U10007 ( .A1(n8415), .A2(n8416), .ZN(n8434) );
  AOI21_X1 U10008 ( .B1(n8416), .B2(n8415), .A(n8434), .ZN(n8420) );
  AOI22_X1 U10009 ( .A1(n10047), .A2(n8417), .B1(n10045), .B2(
        P2_ADDR_REG_14__SCAN_IN), .ZN(n8419) );
  OAI211_X1 U10010 ( .C1(n8420), .C2(n8542), .A(n8419), .B(n8418), .ZN(n8421)
         );
  NOR2_X1 U10011 ( .A1(n8422), .A2(n8421), .ZN(n8423) );
  OAI21_X1 U10012 ( .B1(n8424), .B2(n10032), .A(n8423), .ZN(P2_U3196) );
  NOR2_X1 U10013 ( .A1(n8425), .A2(n8430), .ZN(n8446) );
  AOI21_X1 U10014 ( .B1(n8430), .B2(n8425), .A(n8446), .ZN(n8444) );
  AOI21_X1 U10015 ( .B1(n8431), .B2(n8428), .A(n8459), .ZN(n8429) );
  NOR2_X1 U10016 ( .A1(n8429), .A2(n8486), .ZN(n8442) );
  MUX2_X1 U10017 ( .A(n8431), .B(n8430), .S(n8529), .Z(n8433) );
  AND2_X1 U10018 ( .A1(n8458), .A2(n8433), .ZN(n8451) );
  INV_X1 U10019 ( .A(n8451), .ZN(n8432) );
  OAI21_X1 U10020 ( .B1(n8458), .B2(n8433), .A(n8432), .ZN(n8437) );
  NOR2_X1 U10021 ( .A1(n8436), .A2(n8437), .ZN(n8450) );
  AOI21_X1 U10022 ( .B1(n8437), .B2(n8436), .A(n8450), .ZN(n8440) );
  AOI22_X1 U10023 ( .A1(n10047), .A2(n8458), .B1(n10045), .B2(
        P2_ADDR_REG_15__SCAN_IN), .ZN(n8439) );
  OAI211_X1 U10024 ( .C1(n8440), .C2(n8542), .A(n8439), .B(n8438), .ZN(n8441)
         );
  NOR2_X1 U10025 ( .A1(n8442), .A2(n8441), .ZN(n8443) );
  OAI21_X1 U10026 ( .B1(n8444), .B2(n10032), .A(n8443), .ZN(P2_U3197) );
  NOR2_X1 U10027 ( .A1(n8458), .A2(n8445), .ZN(n8447) );
  NOR2_X1 U10028 ( .A1(n8447), .A2(n8446), .ZN(n8449) );
  AOI22_X1 U10029 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8461), .B1(n8481), .B2(
        n8787), .ZN(n8448) );
  NOR2_X1 U10030 ( .A1(n8449), .A2(n8448), .ZN(n8471) );
  AOI21_X1 U10031 ( .B1(n8449), .B2(n8448), .A(n8471), .ZN(n8470) );
  MUX2_X1 U10032 ( .A(n8716), .B(n8787), .S(n8529), .Z(n8452) );
  NAND2_X1 U10033 ( .A1(n8452), .A2(n8461), .ZN(n8473) );
  NOR2_X1 U10034 ( .A1(n8452), .A2(n8461), .ZN(n8475) );
  INV_X1 U10035 ( .A(n8475), .ZN(n8453) );
  NAND2_X1 U10036 ( .A1(n8473), .A2(n8453), .ZN(n8454) );
  XNOR2_X1 U10037 ( .A(n8474), .B(n8454), .ZN(n8468) );
  NAND2_X1 U10038 ( .A1(n10045), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n8456) );
  OAI211_X1 U10039 ( .C1(n10023), .C2(n8481), .A(n8456), .B(n8455), .ZN(n8467)
         );
  NOR2_X1 U10040 ( .A1(n8458), .A2(n8457), .ZN(n8460) );
  MUX2_X1 U10041 ( .A(n8716), .B(P2_REG2_REG_16__SCAN_IN), .S(n8461), .Z(n8462) );
  INV_X1 U10042 ( .A(n8462), .ZN(n8463) );
  NOR2_X1 U10043 ( .A1(n8464), .A2(n8463), .ZN(n8480) );
  AOI21_X1 U10044 ( .B1(n8464), .B2(n8463), .A(n8480), .ZN(n8465) );
  NOR2_X1 U10045 ( .A1(n8465), .A2(n8486), .ZN(n8466) );
  AOI211_X1 U10046 ( .C1(n10051), .C2(n8468), .A(n8467), .B(n8466), .ZN(n8469)
         );
  OAI21_X1 U10047 ( .B1(n8470), .B2(n10032), .A(n8469), .ZN(P2_U3198) );
  AOI21_X1 U10048 ( .B1(n8783), .B2(n8472), .A(n8493), .ZN(n8491) );
  OAI21_X1 U10049 ( .B1(n8475), .B2(n8474), .A(n8473), .ZN(n8478) );
  MUX2_X1 U10050 ( .A(n8700), .B(n8783), .S(n8529), .Z(n8506) );
  XNOR2_X1 U10051 ( .A(n8476), .B(n8506), .ZN(n8477) );
  NAND2_X1 U10052 ( .A1(n8477), .A2(n8478), .ZN(n8503) );
  OAI21_X1 U10053 ( .B1(n8478), .B2(n8477), .A(n8503), .ZN(n8489) );
  NOR2_X1 U10054 ( .A1(n8518), .A2(n8479), .ZN(n8488) );
  AOI21_X1 U10055 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n8481), .A(n8480), .ZN(
        n8496) );
  AOI21_X1 U10056 ( .B1(n8482), .B2(n8700), .A(n8497), .ZN(n8485) );
  NAND2_X1 U10057 ( .A1(n10047), .A2(n8505), .ZN(n8483) );
  OAI211_X1 U10058 ( .C1(n8486), .C2(n8485), .A(n8484), .B(n8483), .ZN(n8487)
         );
  AOI211_X1 U10059 ( .C1(n8489), .C2(n10051), .A(n8488), .B(n8487), .ZN(n8490)
         );
  OAI21_X1 U10060 ( .B1(n8491), .B2(n10032), .A(n8490), .ZN(P2_U3199) );
  NOR2_X1 U10061 ( .A1(n8505), .A2(n8492), .ZN(n8494) );
  NAND2_X1 U10062 ( .A1(n8499), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8521) );
  OAI21_X1 U10063 ( .B1(n8499), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8521), .ZN(
        n8495) );
  AOI21_X1 U10064 ( .B1(n4389), .B2(n8495), .A(n8523), .ZN(n8520) );
  NOR2_X1 U10065 ( .A1(n8505), .A2(n8496), .ZN(n8498) );
  NAND2_X1 U10066 ( .A1(n8499), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8525) );
  OAI21_X1 U10067 ( .B1(n8499), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8525), .ZN(
        n8500) );
  AOI21_X1 U10068 ( .B1(n8501), .B2(n8500), .A(n8527), .ZN(n8502) );
  INV_X1 U10069 ( .A(n8502), .ZN(n8519) );
  INV_X1 U10070 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8517) );
  INV_X1 U10071 ( .A(n8503), .ZN(n8504) );
  MUX2_X1 U10072 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8529), .Z(n8508) );
  NAND2_X1 U10073 ( .A1(n8507), .A2(n8508), .ZN(n8533) );
  INV_X1 U10074 ( .A(n8507), .ZN(n8510) );
  INV_X1 U10075 ( .A(n8508), .ZN(n8509) );
  NAND2_X1 U10076 ( .A1(n8510), .A2(n8509), .ZN(n8534) );
  AOI21_X1 U10077 ( .B1(n8512), .B2(n8511), .A(n10047), .ZN(n8513) );
  MUX2_X1 U10078 ( .A(n8514), .B(n8513), .S(n8532), .Z(n8515) );
  OAI21_X1 U10079 ( .B1(n8520), .B2(n10032), .A(n4416), .ZN(P2_U3200) );
  INV_X1 U10080 ( .A(n8521), .ZN(n8522) );
  NOR2_X1 U10081 ( .A1(n8523), .A2(n8522), .ZN(n8524) );
  XNOR2_X1 U10082 ( .A(n5543), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8530) );
  INV_X1 U10083 ( .A(n8525), .ZN(n8526) );
  NOR2_X1 U10084 ( .A1(n8527), .A2(n8526), .ZN(n8528) );
  MUX2_X1 U10085 ( .A(n8680), .B(P2_REG2_REG_19__SCAN_IN), .S(n5543), .Z(n8531) );
  XNOR2_X1 U10086 ( .A(n8528), .B(n8531), .ZN(n8545) );
  MUX2_X1 U10087 ( .A(n8531), .B(n8530), .S(n8529), .Z(n8537) );
  NAND2_X1 U10088 ( .A1(n8533), .A2(n8532), .ZN(n8535) );
  NAND2_X1 U10089 ( .A1(n8535), .A2(n8534), .ZN(n8536) );
  XNOR2_X1 U10090 ( .A(n8537), .B(n8536), .ZN(n8543) );
  NAND2_X1 U10091 ( .A1(n10045), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8541) );
  AOI21_X1 U10092 ( .B1(n10047), .B2(n8539), .A(n8538), .ZN(n8540) );
  OAI211_X1 U10093 ( .C1(n8543), .C2(n8542), .A(n8541), .B(n8540), .ZN(n8544)
         );
  AOI21_X1 U10094 ( .B1(n8545), .B2(n10056), .A(n8544), .ZN(n8546) );
  OAI21_X1 U10095 ( .B1(n4917), .B2(n10032), .A(n8546), .ZN(P2_U3201) );
  INV_X1 U10096 ( .A(n8741), .ZN(n8551) );
  NAND2_X1 U10097 ( .A1(n8547), .A2(n8719), .ZN(n8555) );
  AOI21_X1 U10098 ( .B1(n8555), .B2(n8744), .A(n8734), .ZN(n8552) );
  AOI21_X1 U10099 ( .B1(n8734), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8552), .ZN(
        n8550) );
  OAI21_X1 U10100 ( .B1(n8551), .B2(n8594), .A(n8550), .ZN(P2_U3202) );
  AOI21_X1 U10101 ( .B1(n8734), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8552), .ZN(
        n8553) );
  OAI21_X1 U10102 ( .B1(n8746), .B2(n8594), .A(n8553), .ZN(P2_U3203) );
  NAND2_X1 U10103 ( .A1(n8554), .A2(n10069), .ZN(n8560) );
  OAI21_X1 U10104 ( .B1(n8715), .B2(n8556), .A(n8555), .ZN(n8557) );
  AOI21_X1 U10105 ( .B1(n8558), .B2(n8735), .A(n8557), .ZN(n8559) );
  OAI211_X1 U10106 ( .C1(n8561), .C2(n8738), .A(n8560), .B(n8559), .ZN(
        P2_U3204) );
  XNOR2_X1 U10107 ( .A(n8562), .B(n8568), .ZN(n8567) );
  NOR2_X1 U10108 ( .A1(n8711), .A2(n8563), .ZN(n8565) );
  INV_X1 U10109 ( .A(n8748), .ZN(n8574) );
  XNOR2_X1 U10110 ( .A(n8569), .B(n8568), .ZN(n8747) );
  AOI22_X1 U10111 ( .A1(n8570), .A2(n8719), .B1(n8734), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n8571) );
  OAI21_X1 U10112 ( .B1(n8801), .B2(n8594), .A(n8571), .ZN(n8572) );
  AOI21_X1 U10113 ( .B1(n8747), .B2(n8596), .A(n8572), .ZN(n8573) );
  OAI21_X1 U10114 ( .B1(n8574), .B2(n8734), .A(n8573), .ZN(P2_U3205) );
  XOR2_X1 U10115 ( .A(n8580), .B(n8575), .Z(n8576) );
  OAI222_X1 U10116 ( .A1(n8669), .A2(n8578), .B1(n8711), .B2(n8577), .C1(n8576), .C2(n8666), .ZN(n8751) );
  INV_X1 U10117 ( .A(n8751), .ZN(n8585) );
  XOR2_X1 U10118 ( .A(n8580), .B(n8579), .Z(n8752) );
  AOI22_X1 U10119 ( .A1(n8734), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8581), .B2(
        n8719), .ZN(n8582) );
  OAI21_X1 U10120 ( .B1(n8805), .B2(n8594), .A(n8582), .ZN(n8583) );
  AOI21_X1 U10121 ( .B1(n8752), .B2(n8596), .A(n8583), .ZN(n8584) );
  OAI21_X1 U10122 ( .B1(n8585), .B2(n8734), .A(n8584), .ZN(P2_U3206) );
  XNOR2_X1 U10123 ( .A(n8586), .B(n8591), .ZN(n8587) );
  OAI222_X1 U10124 ( .A1(n8711), .A2(n8589), .B1(n8669), .B2(n8588), .C1(n8666), .C2(n8587), .ZN(n8806) );
  AOI21_X1 U10125 ( .B1(n8719), .B2(n8590), .A(n8806), .ZN(n8598) );
  XNOR2_X1 U10126 ( .A(n8592), .B(n8591), .ZN(n8756) );
  OAI22_X1 U10127 ( .A1(n8807), .A2(n8594), .B1(n8593), .B2(n10069), .ZN(n8595) );
  AOI21_X1 U10128 ( .B1(n8756), .B2(n8596), .A(n8595), .ZN(n8597) );
  OAI21_X1 U10129 ( .B1(n8598), .B2(n8734), .A(n8597), .ZN(P2_U3207) );
  XOR2_X1 U10130 ( .A(n8599), .B(n8600), .Z(n8813) );
  AND2_X1 U10131 ( .A1(n8601), .A2(n8600), .ZN(n8602) );
  NAND2_X1 U10132 ( .A1(n8603), .A2(n8731), .ZN(n8606) );
  AOI22_X1 U10133 ( .A1(n8604), .A2(n8728), .B1(n8726), .B2(n8628), .ZN(n8605)
         );
  NAND2_X1 U10134 ( .A1(n8606), .A2(n8605), .ZN(n8811) );
  NOR2_X1 U10135 ( .A1(n8812), .A2(n10061), .ZN(n8607) );
  OAI21_X1 U10136 ( .B1(n8811), .B2(n8607), .A(n8715), .ZN(n8610) );
  AOI22_X1 U10137 ( .A1(n8734), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8719), .B2(
        n8608), .ZN(n8609) );
  OAI211_X1 U10138 ( .C1(n8813), .C2(n8738), .A(n8610), .B(n8609), .ZN(
        P2_U3208) );
  XNOR2_X1 U10139 ( .A(n8611), .B(n8619), .ZN(n8613) );
  AOI222_X1 U10140 ( .A1(n8731), .A2(n8613), .B1(n8641), .B2(n8726), .C1(n8612), .C2(n8728), .ZN(n8816) );
  AOI22_X1 U10141 ( .A1(n8818), .A2(n8615), .B1(n8719), .B2(n8614), .ZN(n8616)
         );
  AOI21_X1 U10142 ( .B1(n8816), .B2(n8616), .A(n8734), .ZN(n8623) );
  NAND2_X1 U10143 ( .A1(n8618), .A2(n8617), .ZN(n8620) );
  XNOR2_X1 U10144 ( .A(n8620), .B(n8619), .ZN(n8821) );
  OAI22_X1 U10145 ( .A1(n8821), .A2(n8738), .B1(n8621), .B2(n10069), .ZN(n8622) );
  OR2_X1 U10146 ( .A1(n8623), .A2(n8622), .ZN(P2_U3209) );
  XNOR2_X1 U10147 ( .A(n8625), .B(n8624), .ZN(n8827) );
  INV_X1 U10148 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8630) );
  XNOR2_X1 U10149 ( .A(n8627), .B(n8626), .ZN(n8629) );
  AOI222_X1 U10150 ( .A1(n8731), .A2(n8629), .B1(n8655), .B2(n8726), .C1(n8628), .C2(n8728), .ZN(n8822) );
  MUX2_X1 U10151 ( .A(n8630), .B(n8822), .S(n10069), .Z(n8633) );
  AOI22_X1 U10152 ( .A1(n8824), .A2(n8735), .B1(n8719), .B2(n8631), .ZN(n8632)
         );
  OAI211_X1 U10153 ( .C1(n8827), .C2(n8738), .A(n8633), .B(n8632), .ZN(
        P2_U3210) );
  XNOR2_X1 U10154 ( .A(n8634), .B(n8637), .ZN(n8833) );
  NAND3_X1 U10155 ( .A1(n8635), .A2(n8637), .A3(n8636), .ZN(n8638) );
  NAND2_X1 U10156 ( .A1(n8639), .A2(n8638), .ZN(n8642) );
  AOI222_X1 U10157 ( .A1(n8731), .A2(n8642), .B1(n8641), .B2(n8728), .C1(n8640), .C2(n8726), .ZN(n8828) );
  MUX2_X1 U10158 ( .A(n8643), .B(n8828), .S(n8715), .Z(n8646) );
  AOI22_X1 U10159 ( .A1(n8830), .A2(n8735), .B1(n8719), .B2(n8644), .ZN(n8645)
         );
  OAI211_X1 U10160 ( .C1(n8833), .C2(n8738), .A(n8646), .B(n8645), .ZN(
        P2_U3211) );
  NAND2_X1 U10161 ( .A1(n8648), .A2(n8647), .ZN(n8649) );
  XNOR2_X1 U10162 ( .A(n8649), .B(n8651), .ZN(n8839) );
  INV_X1 U10163 ( .A(n8651), .ZN(n8653) );
  NAND3_X1 U10164 ( .A1(n8650), .A2(n8653), .A3(n8652), .ZN(n8654) );
  NAND2_X1 U10165 ( .A1(n8635), .A2(n8654), .ZN(n8656) );
  AOI222_X1 U10166 ( .A1(n8731), .A2(n8656), .B1(n8678), .B2(n8726), .C1(n8655), .C2(n8728), .ZN(n8834) );
  MUX2_X1 U10167 ( .A(n8657), .B(n8834), .S(n8715), .Z(n8660) );
  AOI22_X1 U10168 ( .A1(n8836), .A2(n8735), .B1(n8719), .B2(n8658), .ZN(n8659)
         );
  OAI211_X1 U10169 ( .C1(n8839), .C2(n8738), .A(n8660), .B(n8659), .ZN(
        P2_U3212) );
  XOR2_X1 U10170 ( .A(n8661), .B(n8664), .Z(n8843) );
  INV_X1 U10171 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8671) );
  INV_X1 U10172 ( .A(n8650), .ZN(n8663) );
  AOI21_X1 U10173 ( .B1(n8664), .B2(n8662), .A(n8663), .ZN(n8665) );
  OAI222_X1 U10174 ( .A1(n8669), .A2(n8668), .B1(n8711), .B2(n8667), .C1(n8666), .C2(n8665), .ZN(n8840) );
  INV_X1 U10175 ( .A(n8840), .ZN(n8670) );
  MUX2_X1 U10176 ( .A(n8671), .B(n8670), .S(n8715), .Z(n8674) );
  AOI22_X1 U10177 ( .A1(n8773), .A2(n8735), .B1(n8719), .B2(n8672), .ZN(n8673)
         );
  OAI211_X1 U10178 ( .C1(n8843), .C2(n8738), .A(n8674), .B(n8673), .ZN(
        P2_U3213) );
  XOR2_X1 U10179 ( .A(n8675), .B(n8676), .Z(n8851) );
  XOR2_X1 U10180 ( .A(n8677), .B(n8676), .Z(n8679) );
  AOI222_X1 U10181 ( .A1(n8731), .A2(n8679), .B1(n8678), .B2(n8728), .C1(n8698), .C2(n8726), .ZN(n8846) );
  MUX2_X1 U10182 ( .A(n8680), .B(n8846), .S(n8715), .Z(n8684) );
  INV_X1 U10183 ( .A(n8681), .ZN(n8682) );
  AOI22_X1 U10184 ( .A1(n8848), .A2(n8735), .B1(n8719), .B2(n8682), .ZN(n8683)
         );
  OAI211_X1 U10185 ( .C1(n8851), .C2(n8738), .A(n8684), .B(n8683), .ZN(
        P2_U3214) );
  XOR2_X1 U10186 ( .A(n8687), .B(n8685), .Z(n8857) );
  INV_X1 U10187 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8691) );
  XOR2_X1 U10188 ( .A(n8686), .B(n8687), .Z(n8690) );
  AOI222_X1 U10189 ( .A1(n8731), .A2(n8690), .B1(n8689), .B2(n8728), .C1(n8688), .C2(n8726), .ZN(n8852) );
  MUX2_X1 U10190 ( .A(n8691), .B(n8852), .S(n10069), .Z(n8695) );
  INV_X1 U10191 ( .A(n8692), .ZN(n8693) );
  AOI22_X1 U10192 ( .A1(n8854), .A2(n8735), .B1(n8719), .B2(n8693), .ZN(n8694)
         );
  OAI211_X1 U10193 ( .C1(n8857), .C2(n8738), .A(n8695), .B(n8694), .ZN(
        P2_U3215) );
  XNOR2_X1 U10194 ( .A(n8696), .B(n4862), .ZN(n8863) );
  XNOR2_X1 U10195 ( .A(n8697), .B(n4862), .ZN(n8699) );
  AOI222_X1 U10196 ( .A1(n8731), .A2(n8699), .B1(n8729), .B2(n8726), .C1(n8698), .C2(n8728), .ZN(n8858) );
  MUX2_X1 U10197 ( .A(n8700), .B(n8858), .S(n8715), .Z(n8704) );
  INV_X1 U10198 ( .A(n8701), .ZN(n8702) );
  AOI22_X1 U10199 ( .A1(n8860), .A2(n8735), .B1(n8719), .B2(n8702), .ZN(n8703)
         );
  OAI211_X1 U10200 ( .C1(n8863), .C2(n8738), .A(n8704), .B(n8703), .ZN(
        P2_U3216) );
  XNOR2_X1 U10201 ( .A(n8706), .B(n8705), .ZN(n8871) );
  XNOR2_X1 U10202 ( .A(n8708), .B(n8707), .ZN(n8714) );
  NAND2_X1 U10203 ( .A1(n8709), .A2(n8726), .ZN(n8710) );
  OAI21_X1 U10204 ( .B1(n8712), .B2(n8711), .A(n8710), .ZN(n8713) );
  AOI21_X1 U10205 ( .B1(n8714), .B2(n8731), .A(n8713), .ZN(n8864) );
  MUX2_X1 U10206 ( .A(n8716), .B(n8864), .S(n8715), .Z(n8721) );
  INV_X1 U10207 ( .A(n8717), .ZN(n8718) );
  AOI22_X1 U10208 ( .A1(n8867), .A2(n8735), .B1(n8719), .B2(n8718), .ZN(n8720)
         );
  OAI211_X1 U10209 ( .C1(n8871), .C2(n8738), .A(n8721), .B(n8720), .ZN(
        P2_U3217) );
  XNOR2_X1 U10210 ( .A(n8722), .B(n8723), .ZN(n8795) );
  INV_X1 U10211 ( .A(n8795), .ZN(n8739) );
  XNOR2_X1 U10212 ( .A(n8724), .B(n8725), .ZN(n8730) );
  AOI222_X1 U10213 ( .A1(n8731), .A2(n8730), .B1(n8729), .B2(n8728), .C1(n8727), .C2(n8726), .ZN(n8797) );
  OAI21_X1 U10214 ( .B1(n8732), .B2(n10064), .A(n8797), .ZN(n8733) );
  NAND2_X1 U10215 ( .A1(n8733), .A2(n10069), .ZN(n8737) );
  AOI22_X1 U10216 ( .A1(n8792), .A2(n8735), .B1(P2_REG2_REG_15__SCAN_IN), .B2(
        n8734), .ZN(n8736) );
  OAI211_X1 U10217 ( .C1(n8739), .C2(n8738), .A(n8737), .B(n8736), .ZN(
        P2_U3218) );
  INV_X1 U10218 ( .A(n8744), .ZN(n8740) );
  AOI21_X1 U10219 ( .B1(n8741), .B2(n8793), .A(n8740), .ZN(n9780) );
  INV_X1 U10220 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8742) );
  OR2_X1 U10221 ( .A1(n8786), .A2(n8742), .ZN(n8743) );
  OAI21_X1 U10222 ( .B1(n9780), .B2(n8755), .A(n8743), .ZN(P2_U3490) );
  OAI21_X1 U10223 ( .B1(n8746), .B2(n8745), .A(n8744), .ZN(n9782) );
  MUX2_X1 U10224 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9782), .S(n8786), .Z(
        P2_U3489) );
  NOR2_X1 U10225 ( .A1(n8748), .A2(n4900), .ZN(n8798) );
  INV_X1 U10226 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8749) );
  OAI21_X1 U10227 ( .B1(n8801), .B2(n8774), .A(n8750), .ZN(P2_U3487) );
  AOI21_X1 U10228 ( .B1(n8794), .B2(n8752), .A(n8751), .ZN(n8802) );
  INV_X1 U10229 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8753) );
  OAI21_X1 U10230 ( .B1(n8805), .B2(n8774), .A(n8754), .ZN(P2_U3486) );
  MUX2_X1 U10231 ( .A(n8806), .B(P2_REG1_REG_26__SCAN_IN), .S(n8755), .Z(n8758) );
  INV_X1 U10232 ( .A(n8756), .ZN(n8808) );
  OAI22_X1 U10233 ( .A1(n8808), .A2(n8791), .B1(n8807), .B2(n8774), .ZN(n8757)
         );
  OR2_X1 U10234 ( .A1(n8758), .A2(n8757), .ZN(P2_U3485) );
  MUX2_X1 U10235 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8811), .S(n8786), .Z(n8760) );
  OAI22_X1 U10236 ( .A1(n8813), .A2(n8791), .B1(n8812), .B2(n8774), .ZN(n8759)
         );
  OR2_X1 U10237 ( .A1(n8760), .A2(n8759), .ZN(P2_U3484) );
  INV_X1 U10238 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8761) );
  MUX2_X1 U10239 ( .A(n8761), .B(n8816), .S(n8786), .Z(n8763) );
  NAND2_X1 U10240 ( .A1(n8818), .A2(n8788), .ZN(n8762) );
  OAI211_X1 U10241 ( .C1(n8791), .C2(n8821), .A(n8763), .B(n8762), .ZN(
        P2_U3483) );
  INV_X1 U10242 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8764) );
  MUX2_X1 U10243 ( .A(n8764), .B(n8822), .S(n8786), .Z(n8766) );
  NAND2_X1 U10244 ( .A1(n8824), .A2(n8788), .ZN(n8765) );
  OAI211_X1 U10245 ( .C1(n8827), .C2(n8791), .A(n8766), .B(n8765), .ZN(
        P2_U3482) );
  INV_X1 U10246 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8767) );
  MUX2_X1 U10247 ( .A(n8767), .B(n8828), .S(n8786), .Z(n8769) );
  NAND2_X1 U10248 ( .A1(n8830), .A2(n8788), .ZN(n8768) );
  OAI211_X1 U10249 ( .C1(n8833), .C2(n8791), .A(n8769), .B(n8768), .ZN(
        P2_U3481) );
  INV_X1 U10250 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8770) );
  MUX2_X1 U10251 ( .A(n8770), .B(n8834), .S(n8786), .Z(n8772) );
  NAND2_X1 U10252 ( .A1(n8836), .A2(n8788), .ZN(n8771) );
  OAI211_X1 U10253 ( .C1(n8791), .C2(n8839), .A(n8772), .B(n8771), .ZN(
        P2_U3480) );
  MUX2_X1 U10254 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8840), .S(n8786), .Z(n8776) );
  INV_X1 U10255 ( .A(n8773), .ZN(n8842) );
  OAI22_X1 U10256 ( .A1(n8843), .A2(n8791), .B1(n8842), .B2(n8774), .ZN(n8775)
         );
  OR2_X1 U10257 ( .A1(n8776), .A2(n8775), .ZN(P2_U3479) );
  INV_X1 U10258 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8777) );
  MUX2_X1 U10259 ( .A(n8777), .B(n8846), .S(n8786), .Z(n8779) );
  NAND2_X1 U10260 ( .A1(n8848), .A2(n8788), .ZN(n8778) );
  OAI211_X1 U10261 ( .C1(n8791), .C2(n8851), .A(n8779), .B(n8778), .ZN(
        P2_U3478) );
  INV_X1 U10262 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8780) );
  MUX2_X1 U10263 ( .A(n8780), .B(n8852), .S(n8786), .Z(n8782) );
  NAND2_X1 U10264 ( .A1(n8854), .A2(n8788), .ZN(n8781) );
  OAI211_X1 U10265 ( .C1(n8857), .C2(n8791), .A(n8782), .B(n8781), .ZN(
        P2_U3477) );
  MUX2_X1 U10266 ( .A(n8783), .B(n8858), .S(n8786), .Z(n8785) );
  NAND2_X1 U10267 ( .A1(n8860), .A2(n8788), .ZN(n8784) );
  OAI211_X1 U10268 ( .C1(n8863), .C2(n8791), .A(n8785), .B(n8784), .ZN(
        P2_U3476) );
  MUX2_X1 U10269 ( .A(n8787), .B(n8864), .S(n8786), .Z(n8790) );
  NAND2_X1 U10270 ( .A1(n8867), .A2(n8788), .ZN(n8789) );
  OAI211_X1 U10271 ( .C1(n8791), .C2(n8871), .A(n8790), .B(n8789), .ZN(
        P2_U3475) );
  AOI22_X1 U10272 ( .A1(n8795), .A2(n8794), .B1(n8793), .B2(n8792), .ZN(n8796)
         );
  NAND2_X1 U10273 ( .A1(n8797), .A2(n8796), .ZN(n8872) );
  MUX2_X1 U10274 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8872), .S(n8786), .Z(
        P2_U3474) );
  INV_X1 U10275 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8799) );
  OAI21_X1 U10276 ( .B1(n8801), .B2(n8841), .A(n8800), .ZN(P2_U3455) );
  INV_X1 U10277 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8803) );
  OAI21_X1 U10278 ( .B1(n8805), .B2(n8841), .A(n8804), .ZN(P2_U3454) );
  MUX2_X1 U10279 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8806), .S(n10088), .Z(
        n8810) );
  OAI22_X1 U10280 ( .A1(n8808), .A2(n8870), .B1(n8807), .B2(n8841), .ZN(n8809)
         );
  OR2_X1 U10281 ( .A1(n8810), .A2(n8809), .ZN(P2_U3453) );
  MUX2_X1 U10282 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8811), .S(n10088), .Z(
        n8815) );
  OAI22_X1 U10283 ( .A1(n8813), .A2(n8870), .B1(n8812), .B2(n8841), .ZN(n8814)
         );
  OR2_X1 U10284 ( .A1(n8815), .A2(n8814), .ZN(P2_U3452) );
  INV_X1 U10285 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8817) );
  MUX2_X1 U10286 ( .A(n8817), .B(n8816), .S(n10088), .Z(n8820) );
  NAND2_X1 U10287 ( .A1(n8818), .A2(n8866), .ZN(n8819) );
  OAI211_X1 U10288 ( .C1(n8821), .C2(n8870), .A(n8820), .B(n8819), .ZN(
        P2_U3451) );
  INV_X1 U10289 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8823) );
  MUX2_X1 U10290 ( .A(n8823), .B(n8822), .S(n10088), .Z(n8826) );
  NAND2_X1 U10291 ( .A1(n8824), .A2(n8866), .ZN(n8825) );
  OAI211_X1 U10292 ( .C1(n8827), .C2(n8870), .A(n8826), .B(n8825), .ZN(
        P2_U3450) );
  INV_X1 U10293 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8829) );
  MUX2_X1 U10294 ( .A(n8829), .B(n8828), .S(n10088), .Z(n8832) );
  NAND2_X1 U10295 ( .A1(n8830), .A2(n8866), .ZN(n8831) );
  OAI211_X1 U10296 ( .C1(n8833), .C2(n8870), .A(n8832), .B(n8831), .ZN(
        P2_U3449) );
  INV_X1 U10297 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8835) );
  MUX2_X1 U10298 ( .A(n8835), .B(n8834), .S(n10088), .Z(n8838) );
  NAND2_X1 U10299 ( .A1(n8836), .A2(n8866), .ZN(n8837) );
  OAI211_X1 U10300 ( .C1(n8839), .C2(n8870), .A(n8838), .B(n8837), .ZN(
        P2_U3448) );
  MUX2_X1 U10301 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8840), .S(n10088), .Z(
        n8845) );
  OAI22_X1 U10302 ( .A1(n8843), .A2(n8870), .B1(n8842), .B2(n8841), .ZN(n8844)
         );
  OR2_X1 U10303 ( .A1(n8845), .A2(n8844), .ZN(P2_U3447) );
  INV_X1 U10304 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8847) );
  MUX2_X1 U10305 ( .A(n8847), .B(n8846), .S(n10088), .Z(n8850) );
  NAND2_X1 U10306 ( .A1(n8848), .A2(n8866), .ZN(n8849) );
  OAI211_X1 U10307 ( .C1(n8851), .C2(n8870), .A(n8850), .B(n8849), .ZN(
        P2_U3446) );
  INV_X1 U10308 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8853) );
  MUX2_X1 U10309 ( .A(n8853), .B(n8852), .S(n10088), .Z(n8856) );
  NAND2_X1 U10310 ( .A1(n8854), .A2(n8866), .ZN(n8855) );
  OAI211_X1 U10311 ( .C1(n8857), .C2(n8870), .A(n8856), .B(n8855), .ZN(
        P2_U3444) );
  INV_X1 U10312 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8859) );
  MUX2_X1 U10313 ( .A(n8859), .B(n8858), .S(n10088), .Z(n8862) );
  NAND2_X1 U10314 ( .A1(n8860), .A2(n8866), .ZN(n8861) );
  OAI211_X1 U10315 ( .C1(n8863), .C2(n8870), .A(n8862), .B(n8861), .ZN(
        P2_U3441) );
  INV_X1 U10316 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8865) );
  MUX2_X1 U10317 ( .A(n8865), .B(n8864), .S(n10088), .Z(n8869) );
  NAND2_X1 U10318 ( .A1(n8867), .A2(n8866), .ZN(n8868) );
  OAI211_X1 U10319 ( .C1(n8871), .C2(n8870), .A(n8869), .B(n8868), .ZN(
        P2_U3438) );
  MUX2_X1 U10320 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8872), .S(n10088), .Z(
        P2_U3435) );
  INV_X1 U10321 ( .A(n9015), .ZN(n9728) );
  OR2_X1 U10322 ( .A1(n8873), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n8874) );
  NOR4_X1 U10323 ( .A1(n8874), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n4800), .ZN(n8875) );
  AOI21_X1 U10324 ( .B1(n8876), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8875), .ZN(
        n8877) );
  OAI21_X1 U10325 ( .B1(n9728), .B2(n8878), .A(n8877), .ZN(P2_U3264) );
  INV_X1 U10326 ( .A(n8879), .ZN(n9731) );
  OAI222_X1 U10327 ( .A1(P2_U3151), .A2(n5056), .B1(n6665), .B2(n9731), .C1(
        n8881), .C2(n8880), .ZN(P2_U3266) );
  MUX2_X1 U10328 ( .A(n8883), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  AOI21_X1 U10329 ( .B1(n8884), .B2(n8965), .A(n8885), .ZN(n8886) );
  OAI21_X1 U10330 ( .B1(n4383), .B2(n8886), .A(n8997), .ZN(n8890) );
  AOI22_X1 U10331 ( .A1(n9477), .A2(n8999), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n8887) );
  OAI21_X1 U10332 ( .B1(n8980), .B2(n9475), .A(n8887), .ZN(n8888) );
  AOI21_X1 U10333 ( .B1(n8984), .B2(n9507), .A(n8888), .ZN(n8889) );
  OAI211_X1 U10334 ( .C1(n9704), .C2(n9008), .A(n8890), .B(n8889), .ZN(
        P1_U3216) );
  OAI21_X1 U10335 ( .B1(n8893), .B2(n8892), .A(n8891), .ZN(n8894) );
  NAND2_X1 U10336 ( .A1(n8894), .A2(n8997), .ZN(n8900) );
  NAND2_X1 U10337 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9297) );
  INV_X1 U10338 ( .A(n9297), .ZN(n8895) );
  AOI21_X1 U10339 ( .B1(n8999), .B2(n9282), .A(n8895), .ZN(n8899) );
  AOI22_X1 U10340 ( .A1(n8984), .A2(n9284), .B1(n8972), .B2(n8896), .ZN(n8898)
         );
  NAND2_X1 U10341 ( .A1(n9004), .A2(n9951), .ZN(n8897) );
  NAND4_X1 U10342 ( .A1(n8900), .A2(n8899), .A3(n8898), .A4(n8897), .ZN(
        P1_U3218) );
  XOR2_X1 U10343 ( .A(n8902), .B(n8901), .Z(n8908) );
  NAND2_X1 U10344 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9384) );
  OAI21_X1 U10345 ( .B1(n8903), .B2(n8981), .A(n9384), .ZN(n8904) );
  AOI21_X1 U10346 ( .B1(n8984), .B2(n9574), .A(n8904), .ZN(n8905) );
  OAI21_X1 U10347 ( .B1(n8980), .B2(n9539), .A(n8905), .ZN(n8906) );
  AOI21_X1 U10348 ( .B1(n9652), .B2(n8972), .A(n8906), .ZN(n8907) );
  OAI21_X1 U10349 ( .B1(n8908), .B2(n8974), .A(n8907), .ZN(P1_U3219) );
  XOR2_X1 U10350 ( .A(n8909), .B(n8910), .Z(n8915) );
  NAND2_X1 U10351 ( .A1(n9507), .A2(n8999), .ZN(n8912) );
  AOI22_X1 U10352 ( .A1(n9546), .A2(n8984), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n8911) );
  OAI211_X1 U10353 ( .C1(n8980), .C2(n9516), .A(n8912), .B(n8911), .ZN(n8913)
         );
  AOI21_X1 U10354 ( .B1(n9513), .B2(n8972), .A(n8913), .ZN(n8914) );
  OAI21_X1 U10355 ( .B1(n8915), .B2(n8974), .A(n8914), .ZN(P1_U3223) );
  OAI21_X1 U10356 ( .B1(n8917), .B2(n8916), .A(n8988), .ZN(n8918) );
  NAND2_X1 U10357 ( .A1(n8918), .A2(n8997), .ZN(n8924) );
  NOR2_X1 U10358 ( .A1(n8919), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8920) );
  AOI21_X1 U10359 ( .B1(n9477), .B2(n8984), .A(n8920), .ZN(n8921) );
  OAI21_X1 U10360 ( .B1(n8980), .B2(n9454), .A(n8921), .ZN(n8922) );
  AOI21_X1 U10361 ( .B1(n8999), .B2(n9445), .A(n8922), .ZN(n8923) );
  OAI211_X1 U10362 ( .C1(n9699), .C2(n9008), .A(n8924), .B(n8923), .ZN(
        P1_U3225) );
  OAI21_X1 U10363 ( .B1(n8927), .B2(n8925), .A(n8926), .ZN(n8928) );
  NAND2_X1 U10364 ( .A1(n8928), .A2(n8997), .ZN(n8933) );
  AND2_X1 U10365 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9869) );
  AOI21_X1 U10366 ( .B1(n8999), .B2(n9586), .A(n9869), .ZN(n8929) );
  OAI21_X1 U10367 ( .B1(n8930), .B2(n9001), .A(n8929), .ZN(n8931) );
  AOI21_X1 U10368 ( .B1(n9592), .B2(n9004), .A(n8931), .ZN(n8932) );
  OAI211_X1 U10369 ( .C1(n9596), .C2(n9008), .A(n8933), .B(n8932), .ZN(
        P1_U3226) );
  NAND2_X1 U10370 ( .A1(n8936), .A2(n8935), .ZN(n8937) );
  XNOR2_X1 U10371 ( .A(n8934), .B(n8937), .ZN(n8943) );
  NAND2_X1 U10372 ( .A1(n9574), .A2(n8999), .ZN(n8938) );
  NAND2_X1 U10373 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9887) );
  OAI211_X1 U10374 ( .C1(n8939), .C2(n9001), .A(n8938), .B(n9887), .ZN(n8941)
         );
  NOR2_X1 U10375 ( .A1(n9570), .A2(n9008), .ZN(n8940) );
  AOI211_X1 U10376 ( .C1(n9568), .C2(n9004), .A(n8941), .B(n8940), .ZN(n8942)
         );
  OAI21_X1 U10377 ( .B1(n8943), .B2(n8974), .A(n8942), .ZN(P1_U3228) );
  INV_X1 U10378 ( .A(n9626), .ZN(n9465) );
  NOR3_X1 U10379 ( .A1(n4383), .A2(n4467), .A3(n8945), .ZN(n8948) );
  INV_X1 U10380 ( .A(n8946), .ZN(n8947) );
  OAI21_X1 U10381 ( .B1(n8948), .B2(n8947), .A(n8997), .ZN(n8952) );
  AOI22_X1 U10382 ( .A1(n9499), .A2(n8984), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n8949) );
  OAI21_X1 U10383 ( .B1(n8980), .B2(n9462), .A(n8949), .ZN(n8950) );
  AOI21_X1 U10384 ( .B1(n8999), .B2(n9471), .A(n8950), .ZN(n8951) );
  OAI211_X1 U10385 ( .C1(n9465), .C2(n9008), .A(n8952), .B(n8951), .ZN(
        P1_U3229) );
  XNOR2_X1 U10386 ( .A(n8955), .B(n8954), .ZN(n8956) );
  XNOR2_X1 U10387 ( .A(n8953), .B(n8956), .ZN(n8963) );
  OAI22_X1 U10388 ( .A1(n8958), .A2(n8981), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8957), .ZN(n8959) );
  AOI21_X1 U10389 ( .B1(n8984), .B2(n9559), .A(n8959), .ZN(n8960) );
  OAI21_X1 U10390 ( .B1(n8980), .B2(n9526), .A(n8960), .ZN(n8961) );
  AOI21_X1 U10391 ( .B1(n9647), .B2(n8972), .A(n8961), .ZN(n8962) );
  OAI21_X1 U10392 ( .B1(n8963), .B2(n8974), .A(n8962), .ZN(P1_U3233) );
  NAND2_X1 U10393 ( .A1(n8965), .A2(n8964), .ZN(n8966) );
  XOR2_X1 U10394 ( .A(n8967), .B(n8966), .Z(n8975) );
  AOI22_X1 U10395 ( .A1(n9533), .A2(n8984), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n8969) );
  NAND2_X1 U10396 ( .A1(n9493), .A2(n9004), .ZN(n8968) );
  OAI211_X1 U10397 ( .C1(n8970), .C2(n8981), .A(n8969), .B(n8968), .ZN(n8971)
         );
  AOI21_X1 U10398 ( .B1(n9636), .B2(n8972), .A(n8971), .ZN(n8973) );
  OAI21_X1 U10399 ( .B1(n8975), .B2(n8974), .A(n8973), .ZN(P1_U3235) );
  OAI21_X1 U10400 ( .B1(n8978), .B2(n8976), .A(n8977), .ZN(n8979) );
  NAND2_X1 U10401 ( .A1(n8979), .A2(n8997), .ZN(n8986) );
  NOR2_X1 U10402 ( .A1(n8980), .A2(n9552), .ZN(n8983) );
  NAND2_X1 U10403 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9903) );
  OAI21_X1 U10404 ( .B1(n9112), .B2(n8981), .A(n9903), .ZN(n8982) );
  AOI211_X1 U10405 ( .C1(n8984), .C2(n9586), .A(n8983), .B(n8982), .ZN(n8985)
         );
  OAI211_X1 U10406 ( .C1(n9555), .C2(n9008), .A(n8986), .B(n8985), .ZN(
        P1_U3238) );
  AOI22_X1 U10407 ( .A1(n9429), .A2(n9004), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n8991) );
  OAI21_X1 U10408 ( .B1(n8992), .B2(n9001), .A(n8991), .ZN(n8993) );
  AOI21_X1 U10409 ( .B1(n8999), .B2(n9435), .A(n8993), .ZN(n8994) );
  NAND2_X1 U10410 ( .A1(n8998), .A2(n8997), .ZN(n9007) );
  AND2_X1 U10411 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9862) );
  AOI21_X1 U10412 ( .B1(n8999), .B2(n9575), .A(n9862), .ZN(n9000) );
  OAI21_X1 U10413 ( .B1(n9002), .B2(n9001), .A(n9000), .ZN(n9003) );
  AOI21_X1 U10414 ( .B1(n9005), .B2(n9004), .A(n9003), .ZN(n9006) );
  OAI211_X1 U10415 ( .C1(n9009), .C2(n9008), .A(n9007), .B(n9006), .ZN(
        P1_U3241) );
  NAND2_X1 U10416 ( .A1(n9010), .A2(n9014), .ZN(n9013) );
  OR2_X1 U10417 ( .A1(n5673), .A2(n9011), .ZN(n9012) );
  INV_X1 U10418 ( .A(n9275), .ZN(n9150) );
  NAND2_X1 U10419 ( .A1(n9015), .A2(n9014), .ZN(n9017) );
  INV_X1 U10420 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9722) );
  OR2_X1 U10421 ( .A1(n5673), .A2(n9722), .ZN(n9016) );
  INV_X1 U10422 ( .A(n9687), .ZN(n9153) );
  OR2_X1 U10423 ( .A1(n9393), .A2(n9150), .ZN(n9255) );
  INV_X1 U10424 ( .A(n9564), .ZN(n9571) );
  INV_X1 U10425 ( .A(n9088), .ZN(n9035) );
  INV_X1 U10426 ( .A(n9019), .ZN(n9026) );
  INV_X1 U10427 ( .A(n9020), .ZN(n9025) );
  NAND2_X1 U10428 ( .A1(n6417), .A2(n6060), .ZN(n9021) );
  NAND2_X1 U10429 ( .A1(n9022), .A2(n9021), .ZN(n9207) );
  NOR3_X1 U10430 ( .A1(n9207), .A2(n9023), .A3(n6395), .ZN(n9024) );
  NAND4_X1 U10431 ( .A1(n9027), .A2(n9026), .A3(n9025), .A4(n9024), .ZN(n9028)
         );
  NOR2_X1 U10432 ( .A1(n9029), .A2(n9028), .ZN(n9030) );
  NAND3_X1 U10433 ( .A1(n9218), .A2(n6034), .A3(n9030), .ZN(n9031) );
  NOR3_X1 U10434 ( .A1(n9915), .A2(n9032), .A3(n9031), .ZN(n9033) );
  NAND4_X1 U10435 ( .A1(n9036), .A2(n9035), .A3(n9034), .A4(n9033), .ZN(n9037)
         );
  NOR2_X1 U10436 ( .A1(n9581), .A2(n9037), .ZN(n9038) );
  NAND4_X1 U10437 ( .A1(n9544), .A2(n9571), .A3(n9558), .A4(n9038), .ZN(n9039)
         );
  NOR2_X1 U10438 ( .A1(n9530), .A2(n9039), .ZN(n9040) );
  NAND4_X1 U10439 ( .A1(n9481), .A2(n9498), .A3(n9510), .A4(n9040), .ZN(n9041)
         );
  NOR2_X1 U10440 ( .A1(n9125), .A2(n9041), .ZN(n9042) );
  NAND3_X1 U10441 ( .A1(n9434), .A2(n6043), .A3(n9042), .ZN(n9043) );
  NOR2_X1 U10442 ( .A1(n9411), .A2(n9043), .ZN(n9044) );
  AND4_X1 U10443 ( .A1(n9255), .A2(n9045), .A3(n9044), .A4(n9166), .ZN(n9046)
         );
  AND3_X1 U10444 ( .A1(n9254), .A2(n9257), .A3(n9046), .ZN(n9200) );
  NAND2_X1 U10445 ( .A1(n9153), .A2(n4732), .ZN(n9265) );
  AND2_X1 U10446 ( .A1(n9048), .A2(n9057), .ZN(n9211) );
  NAND2_X1 U10447 ( .A1(n9049), .A2(n9217), .ZN(n9058) );
  AOI21_X1 U10448 ( .B1(n9061), .B2(n9211), .A(n9058), .ZN(n9051) );
  OAI21_X1 U10449 ( .B1(n9051), .B2(n9050), .A(n9064), .ZN(n9053) );
  NAND2_X1 U10450 ( .A1(n9053), .A2(n9052), .ZN(n9056) );
  INV_X1 U10451 ( .A(n9054), .ZN(n9055) );
  NAND2_X1 U10452 ( .A1(n9056), .A2(n9055), .ZN(n9070) );
  INV_X1 U10453 ( .A(n9057), .ZN(n9060) );
  INV_X1 U10454 ( .A(n9058), .ZN(n9059) );
  OAI21_X1 U10455 ( .B1(n9061), .B2(n9060), .A(n9059), .ZN(n9063) );
  NAND3_X1 U10456 ( .A1(n9063), .A2(n9925), .A3(n9062), .ZN(n9066) );
  NAND3_X1 U10457 ( .A1(n9066), .A2(n9065), .A3(n9064), .ZN(n9068) );
  NAND3_X1 U10458 ( .A1(n9068), .A2(n9067), .A3(n9071), .ZN(n9069) );
  MUX2_X1 U10459 ( .A(n9070), .B(n9069), .S(n9155), .Z(n9079) );
  AND2_X1 U10460 ( .A1(n9082), .A2(n9076), .ZN(n9072) );
  NAND3_X1 U10461 ( .A1(n9079), .A2(n9072), .A3(n9071), .ZN(n9075) );
  INV_X1 U10462 ( .A(n9072), .ZN(n9221) );
  OAI211_X1 U10463 ( .C1(n9080), .C2(n9221), .A(n9085), .B(n9081), .ZN(n9225)
         );
  INV_X1 U10464 ( .A(n9225), .ZN(n9074) );
  INV_X1 U10465 ( .A(n9224), .ZN(n9073) );
  AOI21_X1 U10466 ( .B1(n9075), .B2(n9074), .A(n9073), .ZN(n9087) );
  INV_X1 U10467 ( .A(n9076), .ZN(n9077) );
  AOI21_X1 U10468 ( .B1(n9079), .B2(n9078), .A(n9077), .ZN(n9084) );
  NAND2_X1 U10469 ( .A1(n9081), .A2(n9080), .ZN(n9083) );
  OAI211_X1 U10470 ( .C1(n9084), .C2(n9083), .A(n9224), .B(n9082), .ZN(n9086)
         );
  INV_X1 U10471 ( .A(n9095), .ZN(n9089) );
  INV_X1 U10472 ( .A(n9227), .ZN(n9094) );
  AOI211_X1 U10473 ( .C1(n9089), .C2(n9230), .A(n9094), .B(n9088), .ZN(n9090)
         );
  NAND2_X1 U10474 ( .A1(n9097), .A2(n9093), .ZN(n9234) );
  OAI21_X1 U10475 ( .B1(n9090), .B2(n9234), .A(n9233), .ZN(n9092) );
  NAND4_X1 U10476 ( .A1(n9241), .A2(n9155), .A3(n9236), .A4(n9232), .ZN(n9091)
         );
  AOI21_X1 U10477 ( .B1(n9092), .B2(n9237), .A(n9091), .ZN(n9115) );
  INV_X1 U10478 ( .A(n9232), .ZN(n9096) );
  AOI21_X1 U10479 ( .B1(n9098), .B2(n9097), .A(n9096), .ZN(n9108) );
  NAND4_X1 U10480 ( .A1(n9240), .A2(n4516), .A3(n9237), .A4(n9239), .ZN(n9107)
         );
  NAND2_X1 U10481 ( .A1(n9102), .A2(n9155), .ZN(n9099) );
  OAI21_X1 U10482 ( .B1(n9239), .B2(n4516), .A(n9099), .ZN(n9105) );
  NAND2_X1 U10483 ( .A1(n9574), .A2(n4516), .ZN(n9100) );
  OAI22_X1 U10484 ( .A1(n9236), .A2(n9100), .B1(n9239), .B2(n9099), .ZN(n9104)
         );
  OAI211_X1 U10485 ( .C1(n9574), .C2(n9239), .A(n9555), .B(n4516), .ZN(n9101)
         );
  AOI21_X1 U10486 ( .B1(n9102), .B2(n9571), .A(n9101), .ZN(n9103) );
  AOI211_X1 U10487 ( .C1(n9657), .C2(n9105), .A(n9104), .B(n9103), .ZN(n9106)
         );
  OAI211_X1 U10488 ( .C1(n9108), .C2(n9107), .A(n9544), .B(n9106), .ZN(n9114)
         );
  INV_X1 U10489 ( .A(n9109), .ZN(n9119) );
  INV_X1 U10490 ( .A(n9242), .ZN(n9111) );
  AOI21_X1 U10491 ( .B1(n9109), .B2(n9542), .A(n9155), .ZN(n9110) );
  OAI33_X1 U10492 ( .A1(n9155), .A2(n9112), .A3(n9119), .B1(n9111), .B2(n9110), 
        .B3(n6040), .ZN(n9113) );
  OAI211_X1 U10493 ( .C1(n9115), .C2(n9114), .A(n9113), .B(n9118), .ZN(n9122)
         );
  AND2_X1 U10494 ( .A1(n9118), .A2(n9116), .ZN(n9176) );
  INV_X1 U10495 ( .A(n9117), .ZN(n9120) );
  OAI21_X1 U10496 ( .B1(n9120), .B2(n9119), .A(n9118), .ZN(n9182) );
  AND2_X1 U10497 ( .A1(n9126), .A2(n9123), .ZN(n9169) );
  NAND2_X1 U10498 ( .A1(n9467), .A2(n9124), .ZN(n9183) );
  OAI21_X1 U10499 ( .B1(n9155), .B2(n9126), .A(n9468), .ZN(n9128) );
  MUX2_X1 U10500 ( .A(n9181), .B(n9172), .S(n9155), .Z(n9127) );
  INV_X1 U10501 ( .A(n9186), .ZN(n9129) );
  OAI211_X1 U10502 ( .C1(n9133), .C2(n9129), .A(n9179), .B(n9175), .ZN(n9130)
         );
  NAND2_X1 U10503 ( .A1(n9130), .A2(n9178), .ZN(n9131) );
  NAND2_X1 U10504 ( .A1(n9131), .A2(n4516), .ZN(n9137) );
  INV_X1 U10505 ( .A(n9175), .ZN(n9132) );
  OAI211_X1 U10506 ( .C1(n9133), .C2(n9132), .A(n9178), .B(n9186), .ZN(n9134)
         );
  NAND2_X1 U10507 ( .A1(n9134), .A2(n9179), .ZN(n9135) );
  INV_X1 U10508 ( .A(n9180), .ZN(n9139) );
  OAI21_X1 U10509 ( .B1(n9156), .B2(n9139), .A(n9138), .ZN(n9143) );
  INV_X1 U10510 ( .A(n9140), .ZN(n9141) );
  AOI21_X1 U10511 ( .B1(n9143), .B2(n9142), .A(n9141), .ZN(n9146) );
  OAI21_X1 U10512 ( .B1(n9146), .B2(n9145), .A(n9144), .ZN(n9149) );
  NAND2_X1 U10513 ( .A1(n9275), .A2(n9389), .ZN(n9147) );
  NAND3_X1 U10514 ( .A1(n9149), .A2(n9148), .A3(n9155), .ZN(n9165) );
  NAND2_X1 U10515 ( .A1(n9275), .A2(n4516), .ZN(n9152) );
  NAND3_X1 U10516 ( .A1(n9393), .A2(n9155), .A3(n9150), .ZN(n9151) );
  OAI211_X1 U10517 ( .C1(n9393), .C2(n9152), .A(n9151), .B(n9389), .ZN(n9154)
         );
  AOI22_X1 U10518 ( .A1(n4363), .A2(n9155), .B1(n9154), .B2(n9153), .ZN(n9164)
         );
  AOI21_X1 U10519 ( .B1(n9156), .B2(n9180), .A(n9189), .ZN(n9158) );
  OAI21_X1 U10520 ( .B1(n9158), .B2(n9167), .A(n9157), .ZN(n9159) );
  NAND2_X1 U10521 ( .A1(n9159), .A2(n9166), .ZN(n9162) );
  OAI21_X1 U10522 ( .B1(n9393), .B2(n9389), .A(n9687), .ZN(n9161) );
  NAND4_X1 U10523 ( .A1(n9162), .A2(n4516), .A3(n9161), .A4(n9160), .ZN(n9163)
         );
  NAND3_X1 U10524 ( .A1(n9165), .A2(n9164), .A3(n9163), .ZN(n9264) );
  INV_X1 U10525 ( .A(n9255), .ZN(n9197) );
  INV_X1 U10526 ( .A(n9166), .ZN(n9168) );
  INV_X1 U10527 ( .A(n9169), .ZN(n9170) );
  NAND2_X1 U10528 ( .A1(n9170), .A2(n9467), .ZN(n9171) );
  NAND2_X1 U10529 ( .A1(n9172), .A2(n9171), .ZN(n9173) );
  NAND2_X1 U10530 ( .A1(n9173), .A2(n9181), .ZN(n9174) );
  NAND2_X1 U10531 ( .A1(n9175), .A2(n9174), .ZN(n9187) );
  INV_X1 U10532 ( .A(n9176), .ZN(n9177) );
  NOR2_X1 U10533 ( .A1(n9187), .A2(n9177), .ZN(n9245) );
  INV_X1 U10534 ( .A(n9178), .ZN(n9250) );
  AOI21_X1 U10535 ( .B1(n9245), .B2(n9531), .A(n9250), .ZN(n9192) );
  AND2_X1 U10536 ( .A1(n9180), .A2(n9179), .ZN(n9249) );
  INV_X1 U10537 ( .A(n9249), .ZN(n9191) );
  INV_X1 U10538 ( .A(n9181), .ZN(n9185) );
  INV_X1 U10539 ( .A(n9182), .ZN(n9184) );
  NOR3_X1 U10540 ( .A1(n9185), .A2(n9184), .A3(n9183), .ZN(n9188) );
  OAI21_X1 U10541 ( .B1(n9188), .B2(n9187), .A(n9186), .ZN(n9190) );
  AOI21_X1 U10542 ( .B1(n9249), .B2(n9190), .A(n9189), .ZN(n9253) );
  OAI21_X1 U10543 ( .B1(n9192), .B2(n9191), .A(n9253), .ZN(n9193) );
  INV_X1 U10544 ( .A(n9193), .ZN(n9194) );
  INV_X1 U10545 ( .A(n9195), .ZN(n9196) );
  INV_X1 U10546 ( .A(n9257), .ZN(n9263) );
  OAI21_X1 U10547 ( .B1(n9199), .B2(n9263), .A(n9198), .ZN(n9203) );
  INV_X1 U10548 ( .A(n9200), .ZN(n9202) );
  INV_X1 U10549 ( .A(n9265), .ZN(n9201) );
  AOI21_X1 U10550 ( .B1(n9203), .B2(n9202), .A(n9201), .ZN(n9205) );
  INV_X1 U10551 ( .A(n9207), .ZN(n9210) );
  AND4_X1 U10552 ( .A1(n6395), .A2(n9210), .A3(n9209), .A4(n9208), .ZN(n9216)
         );
  INV_X1 U10553 ( .A(n9211), .ZN(n9214) );
  INV_X1 U10554 ( .A(n9212), .ZN(n9213) );
  AOI211_X1 U10555 ( .C1(n9216), .C2(n9215), .A(n9214), .B(n9213), .ZN(n9220)
         );
  INV_X1 U10556 ( .A(n9217), .ZN(n9219) );
  OAI21_X1 U10557 ( .B1(n9220), .B2(n9219), .A(n9218), .ZN(n9223) );
  AOI21_X1 U10558 ( .B1(n9223), .B2(n9222), .A(n9221), .ZN(n9226) );
  OAI21_X1 U10559 ( .B1(n9226), .B2(n9225), .A(n9224), .ZN(n9228) );
  NAND2_X1 U10560 ( .A1(n9228), .A2(n9227), .ZN(n9231) );
  AOI21_X1 U10561 ( .B1(n9231), .B2(n9230), .A(n6036), .ZN(n9235) );
  OAI211_X1 U10562 ( .C1(n9235), .C2(n9234), .A(n9233), .B(n9232), .ZN(n9238)
         );
  AOI21_X1 U10563 ( .B1(n9238), .B2(n9237), .A(n6038), .ZN(n9244) );
  NAND2_X1 U10564 ( .A1(n9240), .A2(n9239), .ZN(n9243) );
  OAI211_X1 U10565 ( .C1(n9244), .C2(n9243), .A(n9242), .B(n9241), .ZN(n9247)
         );
  INV_X1 U10566 ( .A(n9245), .ZN(n9246) );
  AOI21_X1 U10567 ( .B1(n9248), .B2(n9247), .A(n9246), .ZN(n9251) );
  OAI21_X1 U10568 ( .B1(n9251), .B2(n9250), .A(n9249), .ZN(n9252) );
  AOI21_X1 U10569 ( .B1(n9253), .B2(n9252), .A(n4370), .ZN(n9256) );
  OAI211_X1 U10570 ( .C1(n9256), .C2(n4731), .A(n9265), .B(n9255), .ZN(n9258)
         );
  NAND2_X1 U10571 ( .A1(n9258), .A2(n9257), .ZN(n9259) );
  MUX2_X1 U10572 ( .A(n9261), .B(n9260), .S(n9259), .Z(n9268) );
  AOI211_X1 U10573 ( .C1(n9263), .C2(n6096), .A(n6021), .B(n9262), .ZN(n9267)
         );
  OAI21_X1 U10574 ( .B1(n4516), .B2(n9265), .A(n9264), .ZN(n9266) );
  AOI22_X1 U10575 ( .A1(n9269), .A2(n9268), .B1(n9267), .B2(n9266), .ZN(n9274)
         );
  NAND2_X1 U10576 ( .A1(n9270), .A2(n9788), .ZN(n9271) );
  OAI211_X1 U10577 ( .C1(n6021), .C2(n9273), .A(n9271), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9272) );
  OAI21_X1 U10578 ( .B1(n9274), .B2(n9273), .A(n9272), .ZN(P1_U3242) );
  MUX2_X1 U10579 ( .A(n9275), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9285), .Z(
        P1_U3584) );
  MUX2_X1 U10580 ( .A(n9276), .B(P1_DATAO_REG_29__SCAN_IN), .S(n9285), .Z(
        P1_U3583) );
  MUX2_X1 U10581 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9416), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10582 ( .A(n9435), .B(P1_DATAO_REG_27__SCAN_IN), .S(n9285), .Z(
        P1_U3581) );
  MUX2_X1 U10583 ( .A(n9445), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9285), .Z(
        P1_U3580) );
  MUX2_X1 U10584 ( .A(n9471), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9285), .Z(
        P1_U3579) );
  MUX2_X1 U10585 ( .A(n9477), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9285), .Z(
        P1_U3578) );
  MUX2_X1 U10586 ( .A(n9499), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9285), .Z(
        P1_U3577) );
  MUX2_X1 U10587 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9507), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10588 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9533), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10589 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9546), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10590 ( .A(n9559), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9285), .Z(
        P1_U3573) );
  MUX2_X1 U10591 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9574), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10592 ( .A(n9586), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9285), .Z(
        P1_U3571) );
  MUX2_X1 U10593 ( .A(n9575), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9285), .Z(
        P1_U3570) );
  MUX2_X1 U10594 ( .A(n9587), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9285), .Z(
        P1_U3569) );
  MUX2_X1 U10595 ( .A(n9277), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9285), .Z(
        P1_U3568) );
  MUX2_X1 U10596 ( .A(n9909), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9285), .Z(
        P1_U3567) );
  MUX2_X1 U10597 ( .A(n9278), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9285), .Z(
        P1_U3566) );
  MUX2_X1 U10598 ( .A(n9910), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9285), .Z(
        P1_U3565) );
  MUX2_X1 U10599 ( .A(n9279), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9285), .Z(
        P1_U3564) );
  MUX2_X1 U10600 ( .A(n9930), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9285), .Z(
        P1_U3563) );
  MUX2_X1 U10601 ( .A(n9922), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9285), .Z(
        P1_U3562) );
  MUX2_X1 U10602 ( .A(n9931), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9285), .Z(
        P1_U3561) );
  MUX2_X1 U10603 ( .A(n9280), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9285), .Z(
        P1_U3560) );
  MUX2_X1 U10604 ( .A(n9281), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9285), .Z(
        P1_U3559) );
  MUX2_X1 U10605 ( .A(n9282), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9285), .Z(
        P1_U3558) );
  MUX2_X1 U10606 ( .A(n9283), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9285), .Z(
        P1_U3557) );
  MUX2_X1 U10607 ( .A(n9284), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9285), .Z(
        P1_U3556) );
  MUX2_X1 U10608 ( .A(n6417), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9285), .Z(
        P1_U3555) );
  MUX2_X1 U10609 ( .A(n6713), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9285), .Z(
        P1_U3554) );
  OAI211_X1 U10610 ( .C1(n9288), .C2(n9287), .A(n9885), .B(n9286), .ZN(n9296)
         );
  OAI211_X1 U10611 ( .C1(n9291), .C2(n9290), .A(n9893), .B(n9289), .ZN(n9295)
         );
  AOI22_X1 U10612 ( .A1(n9870), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9294) );
  NAND2_X1 U10613 ( .A1(n9882), .A2(n9292), .ZN(n9293) );
  NAND4_X1 U10614 ( .A1(n9296), .A2(n9295), .A3(n9294), .A4(n9293), .ZN(
        P1_U3244) );
  INV_X1 U10615 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9298) );
  OAI21_X1 U10616 ( .B1(n9905), .B2(n9298), .A(n9297), .ZN(n9299) );
  AOI21_X1 U10617 ( .B1(n9300), .B2(n9882), .A(n9299), .ZN(n9309) );
  OAI211_X1 U10618 ( .C1(n9303), .C2(n9302), .A(n9893), .B(n9301), .ZN(n9308)
         );
  OAI211_X1 U10619 ( .C1(n9306), .C2(n9305), .A(n9885), .B(n9304), .ZN(n9307)
         );
  NAND3_X1 U10620 ( .A1(n9309), .A2(n9308), .A3(n9307), .ZN(P1_U3246) );
  NAND2_X1 U10621 ( .A1(n9870), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n9310) );
  OAI211_X1 U10622 ( .C1(n9899), .C2(n9312), .A(n9311), .B(n9310), .ZN(n9313)
         );
  INV_X1 U10623 ( .A(n9313), .ZN(n9322) );
  OAI211_X1 U10624 ( .C1(n9316), .C2(n9315), .A(n9885), .B(n9314), .ZN(n9321)
         );
  OAI211_X1 U10625 ( .C1(n9319), .C2(n9318), .A(n9893), .B(n9317), .ZN(n9320)
         );
  NAND4_X1 U10626 ( .A1(n9323), .A2(n9322), .A3(n9321), .A4(n9320), .ZN(
        P1_U3247) );
  INV_X1 U10627 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9325) );
  OAI21_X1 U10628 ( .B1(n9905), .B2(n9325), .A(n9324), .ZN(n9326) );
  AOI21_X1 U10629 ( .B1(n9327), .B2(n9882), .A(n9326), .ZN(n9336) );
  OAI211_X1 U10630 ( .C1(n9330), .C2(n9329), .A(n9893), .B(n9328), .ZN(n9335)
         );
  OAI211_X1 U10631 ( .C1(n9333), .C2(n9332), .A(n9885), .B(n9331), .ZN(n9334)
         );
  NAND3_X1 U10632 ( .A1(n9336), .A2(n9335), .A3(n9334), .ZN(P1_U3248) );
  INV_X1 U10633 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9339) );
  INV_X1 U10634 ( .A(n9337), .ZN(n9338) );
  OAI21_X1 U10635 ( .B1(n9905), .B2(n9339), .A(n9338), .ZN(n9340) );
  AOI21_X1 U10636 ( .B1(n9341), .B2(n9882), .A(n9340), .ZN(n9350) );
  OAI211_X1 U10637 ( .C1(n9344), .C2(n9343), .A(n9885), .B(n9342), .ZN(n9349)
         );
  OAI211_X1 U10638 ( .C1(n9347), .C2(n9346), .A(n9893), .B(n9345), .ZN(n9348)
         );
  NAND3_X1 U10639 ( .A1(n9350), .A2(n9349), .A3(n9348), .ZN(P1_U3250) );
  NAND2_X1 U10640 ( .A1(n9830), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9351) );
  OAI21_X1 U10641 ( .B1(n9830), .B2(P1_REG2_REG_13__SCAN_IN), .A(n9351), .ZN(
        n9826) );
  OAI21_X1 U10642 ( .B1(n9366), .B2(P1_REG2_REG_12__SCAN_IN), .A(n9352), .ZN(
        n9827) );
  NOR2_X1 U10643 ( .A1(n9826), .A2(n9827), .ZN(n9825) );
  AOI21_X1 U10644 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n9830), .A(n9825), .ZN(
        n9837) );
  NAND2_X1 U10645 ( .A1(n9835), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9353) );
  OAI21_X1 U10646 ( .B1(n9835), .B2(P1_REG2_REG_14__SCAN_IN), .A(n9353), .ZN(
        n9838) );
  NOR2_X1 U10647 ( .A1(n9837), .A2(n9838), .ZN(n9836) );
  AOI21_X1 U10648 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n9835), .A(n9836), .ZN(
        n9354) );
  NOR2_X1 U10649 ( .A1(n9354), .A2(n9368), .ZN(n9355) );
  INV_X1 U10650 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9856) );
  XNOR2_X1 U10651 ( .A(n9354), .B(n9368), .ZN(n9857) );
  NOR2_X1 U10652 ( .A1(n9856), .A2(n9857), .ZN(n9855) );
  NOR2_X1 U10653 ( .A1(n9355), .A2(n9855), .ZN(n9867) );
  NAND2_X1 U10654 ( .A1(n9874), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9356) );
  OAI21_X1 U10655 ( .B1(n9874), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9356), .ZN(
        n9866) );
  NOR2_X1 U10656 ( .A1(n9867), .A2(n9866), .ZN(n9865) );
  AOI21_X1 U10657 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n9874), .A(n9865), .ZN(
        n9879) );
  INV_X1 U10658 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9357) );
  XNOR2_X1 U10659 ( .A(n9883), .B(n9357), .ZN(n9878) );
  NAND2_X1 U10660 ( .A1(n9879), .A2(n9878), .ZN(n9359) );
  OR2_X1 U10661 ( .A1(n9883), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9358) );
  NAND2_X1 U10662 ( .A1(n9359), .A2(n9358), .ZN(n9892) );
  NAND2_X1 U10663 ( .A1(n9372), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9360) );
  OAI21_X1 U10664 ( .B1(n9372), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9360), .ZN(
        n9891) );
  NAND2_X1 U10665 ( .A1(n9901), .A2(n9360), .ZN(n9361) );
  XNOR2_X1 U10666 ( .A(n9361), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9378) );
  AOI22_X1 U10667 ( .A1(n9874), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n9363), .B2(
        n9362), .ZN(n9873) );
  MUX2_X1 U10668 ( .A(n9364), .B(P1_REG1_REG_13__SCAN_IN), .S(n9830), .Z(n9823) );
  OAI21_X1 U10669 ( .B1(n9366), .B2(P1_REG1_REG_12__SCAN_IN), .A(n9365), .ZN(
        n9824) );
  NOR2_X1 U10670 ( .A1(n9823), .A2(n9824), .ZN(n9822) );
  AOI21_X1 U10671 ( .B1(n9830), .B2(P1_REG1_REG_13__SCAN_IN), .A(n9822), .ZN(
        n9842) );
  XNOR2_X1 U10672 ( .A(n9835), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n9841) );
  NOR2_X1 U10673 ( .A1(n9842), .A2(n9841), .ZN(n9840) );
  AOI21_X1 U10674 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n9835), .A(n9840), .ZN(
        n9367) );
  NOR2_X1 U10675 ( .A1(n9367), .A2(n9368), .ZN(n9369) );
  XNOR2_X1 U10676 ( .A(n9368), .B(n9367), .ZN(n9854) );
  NOR2_X1 U10677 ( .A1(n9853), .A2(n9854), .ZN(n9852) );
  NOR2_X1 U10678 ( .A1(n9369), .A2(n9852), .ZN(n9872) );
  NAND2_X1 U10679 ( .A1(n9873), .A2(n9872), .ZN(n9871) );
  OAI21_X1 U10680 ( .B1(P1_REG1_REG_16__SCAN_IN), .B2(n9874), .A(n9871), .ZN(
        n9881) );
  XNOR2_X1 U10681 ( .A(n9883), .B(n9371), .ZN(n9880) );
  AOI22_X1 U10682 ( .A1(n9881), .A2(n9880), .B1(n9371), .B2(n9370), .ZN(n9896)
         );
  INV_X1 U10683 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9373) );
  AND2_X1 U10684 ( .A1(n9372), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9374) );
  AOI21_X1 U10685 ( .B1(n9373), .B2(n9898), .A(n9374), .ZN(n9895) );
  NAND2_X1 U10686 ( .A1(n9896), .A2(n9895), .ZN(n9894) );
  INV_X1 U10687 ( .A(n9374), .ZN(n9375) );
  NAND2_X1 U10688 ( .A1(n9894), .A2(n9375), .ZN(n9376) );
  XOR2_X1 U10689 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9376), .Z(n9379) );
  OAI21_X1 U10690 ( .B1(n9379), .B2(n9851), .A(n9899), .ZN(n9377) );
  AOI21_X1 U10691 ( .B1(n9885), .B2(n9378), .A(n9377), .ZN(n9383) );
  INV_X1 U10692 ( .A(n9378), .ZN(n9380) );
  AOI22_X1 U10693 ( .A1(n9380), .A2(n9885), .B1(n9893), .B2(n9379), .ZN(n9382)
         );
  MUX2_X1 U10694 ( .A(n9383), .B(n9382), .S(n9381), .Z(n9385) );
  OAI211_X1 U10695 ( .C1(n9386), .C2(n9905), .A(n9385), .B(n9384), .ZN(
        P1_U3262) );
  XNOR2_X1 U10696 ( .A(n9687), .B(n9396), .ZN(n9387) );
  NOR2_X2 U10697 ( .A1(n9387), .A2(n9590), .ZN(n9603) );
  NAND2_X1 U10698 ( .A1(n9603), .A2(n9949), .ZN(n9391) );
  AND2_X1 U10699 ( .A1(n9389), .A2(n9388), .ZN(n9602) );
  INV_X1 U10700 ( .A(n9602), .ZN(n9606) );
  NOR2_X1 U10701 ( .A1(n9606), .A2(n9593), .ZN(n9398) );
  AOI21_X1 U10702 ( .B1(n9593), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9398), .ZN(
        n9390) );
  OAI211_X1 U10703 ( .C1(n9687), .C2(n9955), .A(n9391), .B(n9390), .ZN(
        P1_U3263) );
  NAND2_X1 U10704 ( .A1(n9393), .A2(n9392), .ZN(n9394) );
  NAND2_X1 U10705 ( .A1(n9394), .A2(n9942), .ZN(n9395) );
  NOR2_X1 U10706 ( .A1(n9691), .A2(n9955), .ZN(n9397) );
  AOI211_X1 U10707 ( .C1(n9593), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9398), .B(
        n9397), .ZN(n9399) );
  OAI21_X1 U10708 ( .B1(n9607), .B2(n9405), .A(n9399), .ZN(P1_U3264) );
  INV_X1 U10709 ( .A(n9400), .ZN(n9408) );
  AOI22_X1 U10710 ( .A1(n9401), .A2(n9952), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9593), .ZN(n9404) );
  NAND2_X1 U10711 ( .A1(n9402), .A2(n9939), .ZN(n9403) );
  OAI211_X1 U10712 ( .C1(n9406), .C2(n9405), .A(n9404), .B(n9403), .ZN(n9407)
         );
  AOI21_X1 U10713 ( .B1(n9408), .B2(n9598), .A(n9407), .ZN(n9409) );
  OAI21_X1 U10714 ( .B1(n9410), .B2(n9601), .A(n9409), .ZN(P1_U3265) );
  XNOR2_X1 U10715 ( .A(n9412), .B(n9411), .ZN(n9612) );
  INV_X1 U10716 ( .A(n9612), .ZN(n9426) );
  NOR2_X1 U10717 ( .A1(n9414), .A2(n9413), .ZN(n9415) );
  AOI22_X1 U10718 ( .A1(n9416), .A2(n7513), .B1(n9932), .B2(n9445), .ZN(n9417)
         );
  AOI211_X1 U10719 ( .C1(n9420), .C2(n9428), .A(n9590), .B(n9419), .ZN(n9611)
         );
  NAND2_X1 U10720 ( .A1(n9611), .A2(n9949), .ZN(n9423) );
  AOI22_X1 U10721 ( .A1(n9421), .A2(n9952), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9593), .ZN(n9422) );
  OAI211_X1 U10722 ( .C1(n6061), .C2(n9955), .A(n9423), .B(n9422), .ZN(n9424)
         );
  AOI21_X1 U10723 ( .B1(n9610), .B2(n9598), .A(n9424), .ZN(n9425) );
  OAI21_X1 U10724 ( .B1(n9426), .B2(n9601), .A(n9425), .ZN(P1_U3266) );
  XNOR2_X1 U10725 ( .A(n9427), .B(n9434), .ZN(n9619) );
  AOI211_X1 U10726 ( .C1(n9616), .C2(n9449), .A(n9590), .B(n9418), .ZN(n9615)
         );
  AOI22_X1 U10727 ( .A1(n9429), .A2(n9952), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9593), .ZN(n9430) );
  OAI21_X1 U10728 ( .B1(n9431), .B2(n9955), .A(n9430), .ZN(n9438) );
  OAI21_X1 U10729 ( .B1(n9434), .B2(n9433), .A(n9432), .ZN(n9436) );
  AOI222_X1 U10730 ( .A1(n9906), .A2(n9436), .B1(n9435), .B2(n7513), .C1(n9471), .C2(n9932), .ZN(n9618) );
  NOR2_X1 U10731 ( .A1(n9618), .A2(n9576), .ZN(n9437) );
  AOI211_X1 U10732 ( .C1(n9615), .C2(n9949), .A(n9438), .B(n9437), .ZN(n9439)
         );
  OAI21_X1 U10733 ( .B1(n9619), .B2(n9601), .A(n9439), .ZN(P1_U3267) );
  NAND2_X1 U10734 ( .A1(n9441), .A2(n9440), .ZN(n9442) );
  NAND2_X1 U10735 ( .A1(n9443), .A2(n9442), .ZN(n9444) );
  NAND2_X1 U10736 ( .A1(n9444), .A2(n9906), .ZN(n9447) );
  AOI22_X1 U10737 ( .A1(n9445), .A2(n7513), .B1(n9932), .B2(n9477), .ZN(n9446)
         );
  NAND2_X1 U10738 ( .A1(n9447), .A2(n9446), .ZN(n9620) );
  INV_X1 U10739 ( .A(n9620), .ZN(n9459) );
  XNOR2_X1 U10740 ( .A(n9448), .B(n6043), .ZN(n9622) );
  NAND2_X1 U10741 ( .A1(n9622), .A2(n9959), .ZN(n9458) );
  INV_X1 U10742 ( .A(n9461), .ZN(n9451) );
  INV_X1 U10743 ( .A(n9449), .ZN(n9450) );
  AOI211_X1 U10744 ( .C1(n9452), .C2(n9451), .A(n9590), .B(n9450), .ZN(n9621)
         );
  NOR2_X1 U10745 ( .A1(n9699), .A2(n9955), .ZN(n9456) );
  OAI22_X1 U10746 ( .A1(n9454), .A2(n9515), .B1(n9453), .B2(n9598), .ZN(n9455)
         );
  AOI211_X1 U10747 ( .C1(n9621), .C2(n9949), .A(n9456), .B(n9455), .ZN(n9457)
         );
  OAI211_X1 U10748 ( .C1(n9593), .C2(n9459), .A(n9458), .B(n9457), .ZN(
        P1_U3268) );
  XNOR2_X1 U10749 ( .A(n9460), .B(n9468), .ZN(n9629) );
  AOI211_X1 U10750 ( .C1(n9626), .C2(n9482), .A(n9590), .B(n9461), .ZN(n9625)
         );
  INV_X1 U10751 ( .A(n9462), .ZN(n9463) );
  AOI22_X1 U10752 ( .A1(n9463), .A2(n9952), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9593), .ZN(n9464) );
  OAI21_X1 U10753 ( .B1(n9465), .B2(n9955), .A(n9464), .ZN(n9473) );
  NAND2_X1 U10754 ( .A1(n9466), .A2(n9467), .ZN(n9469) );
  XNOR2_X1 U10755 ( .A(n9469), .B(n9468), .ZN(n9470) );
  AOI222_X1 U10756 ( .A1(n9499), .A2(n9932), .B1(n9471), .B2(n7513), .C1(n9906), .C2(n9470), .ZN(n9628) );
  NOR2_X1 U10757 ( .A1(n9628), .A2(n9576), .ZN(n9472) );
  AOI211_X1 U10758 ( .C1(n9625), .C2(n9949), .A(n9473), .B(n9472), .ZN(n9474)
         );
  OAI21_X1 U10759 ( .B1(n9629), .B2(n9601), .A(n9474), .ZN(P1_U3269) );
  INV_X1 U10760 ( .A(n9475), .ZN(n9480) );
  OAI21_X1 U10761 ( .B1(n9481), .B2(n9476), .A(n9466), .ZN(n9478) );
  AOI222_X1 U10762 ( .A1(n9906), .A2(n9478), .B1(n9477), .B2(n7513), .C1(n9507), .C2(n9932), .ZN(n9479) );
  INV_X1 U10763 ( .A(n9479), .ZN(n9630) );
  AOI21_X1 U10764 ( .B1(n9480), .B2(n9952), .A(n9630), .ZN(n9488) );
  XNOR2_X1 U10765 ( .A(n4409), .B(n9481), .ZN(n9632) );
  NAND2_X1 U10766 ( .A1(n9632), .A2(n9959), .ZN(n9487) );
  AOI211_X1 U10767 ( .C1(n9483), .C2(n9490), .A(n9590), .B(n4572), .ZN(n9631)
         );
  OAI22_X1 U10768 ( .A1(n9704), .A2(n9955), .B1(n9598), .B2(n9484), .ZN(n9485)
         );
  AOI21_X1 U10769 ( .B1(n9631), .B2(n9949), .A(n9485), .ZN(n9486) );
  OAI211_X1 U10770 ( .C1(n9576), .C2(n9488), .A(n9487), .B(n9486), .ZN(
        P1_U3270) );
  XNOR2_X1 U10771 ( .A(n9489), .B(n9498), .ZN(n9639) );
  INV_X1 U10772 ( .A(n9512), .ZN(n9492) );
  INV_X1 U10773 ( .A(n9490), .ZN(n9491) );
  AOI211_X1 U10774 ( .C1(n9636), .C2(n9492), .A(n9590), .B(n9491), .ZN(n9635)
         );
  AOI22_X1 U10775 ( .A1(n9493), .A2(n9952), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n9593), .ZN(n9494) );
  OAI21_X1 U10776 ( .B1(n9495), .B2(n9955), .A(n9494), .ZN(n9502) );
  OAI21_X1 U10777 ( .B1(n9498), .B2(n9497), .A(n9496), .ZN(n9500) );
  AOI222_X1 U10778 ( .A1(n9906), .A2(n9500), .B1(n9499), .B2(n7513), .C1(n9533), .C2(n9932), .ZN(n9638) );
  NOR2_X1 U10779 ( .A1(n9638), .A2(n9576), .ZN(n9501) );
  AOI211_X1 U10780 ( .C1(n9635), .C2(n9949), .A(n9502), .B(n9501), .ZN(n9503)
         );
  OAI21_X1 U10781 ( .B1(n9639), .B2(n9601), .A(n9503), .ZN(P1_U3271) );
  OAI21_X1 U10782 ( .B1(n9510), .B2(n9505), .A(n9504), .ZN(n9506) );
  NAND2_X1 U10783 ( .A1(n9506), .A2(n9906), .ZN(n9509) );
  AOI22_X1 U10784 ( .A1(n9507), .A2(n7513), .B1(n9932), .B2(n9546), .ZN(n9508)
         );
  NAND2_X1 U10785 ( .A1(n9509), .A2(n9508), .ZN(n9640) );
  INV_X1 U10786 ( .A(n9640), .ZN(n9521) );
  XNOR2_X1 U10787 ( .A(n9511), .B(n9510), .ZN(n9642) );
  NAND2_X1 U10788 ( .A1(n9642), .A2(n9959), .ZN(n9520) );
  AOI211_X1 U10789 ( .C1(n9513), .C2(n9524), .A(n9590), .B(n9512), .ZN(n9641)
         );
  NOR2_X1 U10790 ( .A1(n9710), .A2(n9955), .ZN(n9518) );
  OAI22_X1 U10791 ( .A1(n9516), .A2(n9515), .B1(n9514), .B2(n9598), .ZN(n9517)
         );
  AOI211_X1 U10792 ( .C1(n9641), .C2(n9949), .A(n9518), .B(n9517), .ZN(n9519)
         );
  OAI211_X1 U10793 ( .C1(n9593), .C2(n9521), .A(n9520), .B(n9519), .ZN(
        P1_U3272) );
  XOR2_X1 U10794 ( .A(n9530), .B(n9522), .Z(n9650) );
  INV_X1 U10795 ( .A(n9524), .ZN(n9525) );
  AOI211_X1 U10796 ( .C1(n9647), .C2(n9538), .A(n9590), .B(n9525), .ZN(n9646)
         );
  INV_X1 U10797 ( .A(n9526), .ZN(n9527) );
  AOI22_X1 U10798 ( .A1(n9527), .A2(n9952), .B1(P1_REG2_REG_20__SCAN_IN), .B2(
        n9593), .ZN(n9528) );
  OAI21_X1 U10799 ( .B1(n9529), .B2(n9955), .A(n9528), .ZN(n9535) );
  XOR2_X1 U10800 ( .A(n9531), .B(n9530), .Z(n9532) );
  AOI222_X1 U10801 ( .A1(n9559), .A2(n9932), .B1(n9533), .B2(n7513), .C1(n9906), .C2(n9532), .ZN(n9649) );
  NOR2_X1 U10802 ( .A1(n9649), .A2(n9576), .ZN(n9534) );
  AOI211_X1 U10803 ( .C1(n9646), .C2(n9949), .A(n9535), .B(n9534), .ZN(n9536)
         );
  OAI21_X1 U10804 ( .B1(n9650), .B2(n9601), .A(n9536), .ZN(P1_U3273) );
  XOR2_X1 U10805 ( .A(n9537), .B(n9544), .Z(n9655) );
  AOI211_X1 U10806 ( .C1(n9652), .C2(n9551), .A(n9590), .B(n9523), .ZN(n9651)
         );
  INV_X1 U10807 ( .A(n9539), .ZN(n9540) );
  AOI22_X1 U10808 ( .A1(n9540), .A2(n9952), .B1(n9593), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n9541) );
  OAI21_X1 U10809 ( .B1(n9542), .B2(n9955), .A(n9541), .ZN(n9548) );
  XNOR2_X1 U10810 ( .A(n9543), .B(n9544), .ZN(n9545) );
  AOI222_X1 U10811 ( .A1(n9574), .A2(n9932), .B1(n9546), .B2(n7513), .C1(n9906), .C2(n9545), .ZN(n9654) );
  NOR2_X1 U10812 ( .A1(n9654), .A2(n9576), .ZN(n9547) );
  AOI211_X1 U10813 ( .C1(n9651), .C2(n9949), .A(n9548), .B(n9547), .ZN(n9549)
         );
  OAI21_X1 U10814 ( .B1(n9655), .B2(n9601), .A(n9549), .ZN(P1_U3274) );
  XNOR2_X1 U10815 ( .A(n9550), .B(n9558), .ZN(n9660) );
  AOI211_X1 U10816 ( .C1(n9657), .C2(n9566), .A(n9590), .B(n4573), .ZN(n9656)
         );
  INV_X1 U10817 ( .A(n9552), .ZN(n9553) );
  AOI22_X1 U10818 ( .A1(n9593), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9553), .B2(
        n9952), .ZN(n9554) );
  OAI21_X1 U10819 ( .B1(n9555), .B2(n9955), .A(n9554), .ZN(n9562) );
  OAI21_X1 U10820 ( .B1(n9558), .B2(n9557), .A(n9556), .ZN(n9560) );
  AOI222_X1 U10821 ( .A1(n9906), .A2(n9560), .B1(n9559), .B2(n7513), .C1(n9586), .C2(n9932), .ZN(n9659) );
  NOR2_X1 U10822 ( .A1(n9659), .A2(n9576), .ZN(n9561) );
  AOI211_X1 U10823 ( .C1(n9656), .C2(n9949), .A(n9562), .B(n9561), .ZN(n9563)
         );
  OAI21_X1 U10824 ( .B1(n9660), .B2(n9601), .A(n9563), .ZN(P1_U3275) );
  XNOR2_X1 U10825 ( .A(n9565), .B(n9564), .ZN(n9665) );
  INV_X1 U10826 ( .A(n9589), .ZN(n9567) );
  AOI211_X1 U10827 ( .C1(n9662), .C2(n9567), .A(n9590), .B(n4574), .ZN(n9661)
         );
  AOI22_X1 U10828 ( .A1(n9593), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9568), .B2(
        n9952), .ZN(n9569) );
  OAI21_X1 U10829 ( .B1(n9570), .B2(n9955), .A(n9569), .ZN(n9578) );
  XNOR2_X1 U10830 ( .A(n9572), .B(n9571), .ZN(n9573) );
  AOI222_X1 U10831 ( .A1(n9575), .A2(n9932), .B1(n9574), .B2(n7513), .C1(n9906), .C2(n9573), .ZN(n9664) );
  NOR2_X1 U10832 ( .A1(n9664), .A2(n9576), .ZN(n9577) );
  AOI211_X1 U10833 ( .C1(n9661), .C2(n9949), .A(n9578), .B(n9577), .ZN(n9579)
         );
  OAI21_X1 U10834 ( .B1(n9665), .B2(n9601), .A(n9579), .ZN(P1_U3276) );
  OAI21_X1 U10835 ( .B1(n9582), .B2(n9581), .A(n9580), .ZN(n9670) );
  XNOR2_X1 U10836 ( .A(n9583), .B(n9584), .ZN(n9585) );
  AOI222_X1 U10837 ( .A1(n9587), .A2(n9932), .B1(n9586), .B2(n7513), .C1(n9906), .C2(n9585), .ZN(n9669) );
  INV_X1 U10838 ( .A(n9669), .ZN(n9599) );
  INV_X1 U10839 ( .A(n9588), .ZN(n9591) );
  AOI211_X1 U10840 ( .C1(n9667), .C2(n9591), .A(n9590), .B(n9589), .ZN(n9666)
         );
  NAND2_X1 U10841 ( .A1(n9666), .A2(n9949), .ZN(n9595) );
  AOI22_X1 U10842 ( .A1(n9593), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9592), .B2(
        n9952), .ZN(n9594) );
  OAI211_X1 U10843 ( .C1(n9596), .C2(n9955), .A(n9595), .B(n9594), .ZN(n9597)
         );
  AOI21_X1 U10844 ( .B1(n9599), .B2(n9598), .A(n9597), .ZN(n9600) );
  OAI21_X1 U10845 ( .B1(n9670), .B2(n9601), .A(n9600), .ZN(P1_U3277) );
  NOR2_X1 U10846 ( .A1(n9603), .A2(n9602), .ZN(n9684) );
  MUX2_X1 U10847 ( .A(n9604), .B(n9684), .S(n10021), .Z(n9605) );
  OAI21_X1 U10848 ( .B1(n9687), .B2(n9645), .A(n9605), .ZN(P1_U3553) );
  NAND2_X1 U10849 ( .A1(n9607), .A2(n9606), .ZN(n9688) );
  MUX2_X1 U10850 ( .A(n9688), .B(P1_REG1_REG_30__SCAN_IN), .S(n10019), .Z(
        n9608) );
  INV_X1 U10851 ( .A(n9608), .ZN(n9609) );
  OAI21_X1 U10852 ( .B1(n9691), .B2(n9645), .A(n9609), .ZN(P1_U3552) );
  AOI211_X1 U10853 ( .C1(n9612), .C2(n10007), .A(n9611), .B(n9610), .ZN(n9692)
         );
  MUX2_X1 U10854 ( .A(n9613), .B(n9692), .S(n10021), .Z(n9614) );
  OAI21_X1 U10855 ( .B1(n6061), .B2(n9645), .A(n9614), .ZN(P1_U3549) );
  AOI21_X1 U10856 ( .B1(n9680), .B2(n9616), .A(n9615), .ZN(n9617) );
  OAI211_X1 U10857 ( .C1(n9619), .C2(n9675), .A(n9618), .B(n9617), .ZN(n9695)
         );
  MUX2_X1 U10858 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9695), .S(n10021), .Z(
        P1_U3548) );
  AOI211_X1 U10859 ( .C1(n9622), .C2(n10007), .A(n9621), .B(n9620), .ZN(n9696)
         );
  MUX2_X1 U10860 ( .A(n9623), .B(n9696), .S(n10021), .Z(n9624) );
  OAI21_X1 U10861 ( .B1(n9699), .B2(n9645), .A(n9624), .ZN(P1_U3547) );
  AOI21_X1 U10862 ( .B1(n9680), .B2(n9626), .A(n9625), .ZN(n9627) );
  OAI211_X1 U10863 ( .C1(n9629), .C2(n9675), .A(n9628), .B(n9627), .ZN(n9700)
         );
  MUX2_X1 U10864 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9700), .S(n10021), .Z(
        P1_U3546) );
  AOI211_X1 U10865 ( .C1(n9632), .C2(n10007), .A(n9631), .B(n9630), .ZN(n9701)
         );
  MUX2_X1 U10866 ( .A(n9633), .B(n9701), .S(n10021), .Z(n9634) );
  OAI21_X1 U10867 ( .B1(n9704), .B2(n9645), .A(n9634), .ZN(P1_U3545) );
  AOI21_X1 U10868 ( .B1(n9680), .B2(n9636), .A(n9635), .ZN(n9637) );
  OAI211_X1 U10869 ( .C1(n9639), .C2(n9675), .A(n9638), .B(n9637), .ZN(n9705)
         );
  MUX2_X1 U10870 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9705), .S(n10021), .Z(
        P1_U3544) );
  AOI211_X1 U10871 ( .C1(n9642), .C2(n10007), .A(n9641), .B(n9640), .ZN(n9706)
         );
  MUX2_X1 U10872 ( .A(n9643), .B(n9706), .S(n10021), .Z(n9644) );
  OAI21_X1 U10873 ( .B1(n9710), .B2(n9645), .A(n9644), .ZN(P1_U3543) );
  AOI21_X1 U10874 ( .B1(n9680), .B2(n9647), .A(n9646), .ZN(n9648) );
  OAI211_X1 U10875 ( .C1(n9650), .C2(n9675), .A(n9649), .B(n9648), .ZN(n9711)
         );
  MUX2_X1 U10876 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9711), .S(n10021), .Z(
        P1_U3542) );
  AOI21_X1 U10877 ( .B1(n9680), .B2(n9652), .A(n9651), .ZN(n9653) );
  OAI211_X1 U10878 ( .C1(n9655), .C2(n9675), .A(n9654), .B(n9653), .ZN(n9712)
         );
  MUX2_X1 U10879 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9712), .S(n10021), .Z(
        P1_U3541) );
  AOI21_X1 U10880 ( .B1(n9680), .B2(n9657), .A(n9656), .ZN(n9658) );
  OAI211_X1 U10881 ( .C1(n9660), .C2(n9675), .A(n9659), .B(n9658), .ZN(n9713)
         );
  MUX2_X1 U10882 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9713), .S(n10021), .Z(
        P1_U3540) );
  AOI21_X1 U10883 ( .B1(n9680), .B2(n9662), .A(n9661), .ZN(n9663) );
  OAI211_X1 U10884 ( .C1(n9665), .C2(n9675), .A(n9664), .B(n9663), .ZN(n9714)
         );
  MUX2_X1 U10885 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9714), .S(n10021), .Z(
        P1_U3539) );
  AOI21_X1 U10886 ( .B1(n9680), .B2(n9667), .A(n9666), .ZN(n9668) );
  OAI211_X1 U10887 ( .C1(n9670), .C2(n9675), .A(n9669), .B(n9668), .ZN(n9715)
         );
  MUX2_X1 U10888 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9715), .S(n10021), .Z(
        P1_U3538) );
  AOI21_X1 U10889 ( .B1(n9680), .B2(n9672), .A(n9671), .ZN(n9673) );
  OAI211_X1 U10890 ( .C1(n9676), .C2(n9675), .A(n9674), .B(n9673), .ZN(n9716)
         );
  MUX2_X1 U10891 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9716), .S(n10021), .Z(
        P1_U3537) );
  INV_X1 U10892 ( .A(n9677), .ZN(n9683) );
  AOI21_X1 U10893 ( .B1(n9680), .B2(n9679), .A(n9678), .ZN(n9681) );
  OAI211_X1 U10894 ( .C1(n9683), .C2(n9979), .A(n9682), .B(n9681), .ZN(n9717)
         );
  MUX2_X1 U10895 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9717), .S(n10021), .Z(
        P1_U3536) );
  MUX2_X1 U10896 ( .A(n9685), .B(n9684), .S(n10010), .Z(n9686) );
  OAI21_X1 U10897 ( .B1(n9687), .B2(n9709), .A(n9686), .ZN(P1_U3521) );
  MUX2_X1 U10898 ( .A(n9688), .B(P1_REG0_REG_30__SCAN_IN), .S(n10009), .Z(
        n9689) );
  INV_X1 U10899 ( .A(n9689), .ZN(n9690) );
  OAI21_X1 U10900 ( .B1(n9691), .B2(n9709), .A(n9690), .ZN(P1_U3520) );
  MUX2_X1 U10901 ( .A(n9693), .B(n9692), .S(n10010), .Z(n9694) );
  OAI21_X1 U10902 ( .B1(n6061), .B2(n9709), .A(n9694), .ZN(P1_U3517) );
  MUX2_X1 U10903 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9695), .S(n10010), .Z(
        P1_U3516) );
  MUX2_X1 U10904 ( .A(n9697), .B(n9696), .S(n10010), .Z(n9698) );
  OAI21_X1 U10905 ( .B1(n9699), .B2(n9709), .A(n9698), .ZN(P1_U3515) );
  MUX2_X1 U10906 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9700), .S(n10010), .Z(
        P1_U3514) );
  MUX2_X1 U10907 ( .A(n9702), .B(n9701), .S(n10010), .Z(n9703) );
  OAI21_X1 U10908 ( .B1(n9704), .B2(n9709), .A(n9703), .ZN(P1_U3513) );
  MUX2_X1 U10909 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9705), .S(n10010), .Z(
        P1_U3512) );
  MUX2_X1 U10910 ( .A(n9707), .B(n9706), .S(n10010), .Z(n9708) );
  OAI21_X1 U10911 ( .B1(n9710), .B2(n9709), .A(n9708), .ZN(P1_U3511) );
  MUX2_X1 U10912 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9711), .S(n10010), .Z(
        P1_U3510) );
  MUX2_X1 U10913 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9712), .S(n10010), .Z(
        P1_U3509) );
  MUX2_X1 U10914 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9713), .S(n10010), .Z(
        P1_U3507) );
  MUX2_X1 U10915 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9714), .S(n10010), .Z(
        P1_U3504) );
  MUX2_X1 U10916 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9715), .S(n10010), .Z(
        P1_U3501) );
  MUX2_X1 U10917 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9716), .S(n10010), .Z(
        P1_U3498) );
  MUX2_X1 U10918 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9717), .S(n10010), .Z(
        P1_U3495) );
  MUX2_X1 U10919 ( .A(n9720), .B(P1_D_REG_1__SCAN_IN), .S(n4349), .Z(P1_U3440)
         );
  MUX2_X1 U10920 ( .A(n9721), .B(P1_D_REG_0__SCAN_IN), .S(n4349), .Z(P1_U3439)
         );
  NAND2_X1 U10921 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_STATE_REG_SCAN_IN), 
        .ZN(n9723) );
  OAI22_X1 U10922 ( .A1(n9724), .A2(n9723), .B1(n9722), .B2(n9729), .ZN(n9725)
         );
  INV_X1 U10923 ( .A(n9725), .ZN(n9726) );
  OAI21_X1 U10924 ( .B1(n9728), .B2(n9727), .A(n9726), .ZN(P1_U3324) );
  OAI222_X1 U10925 ( .A1(n9732), .A2(n9731), .B1(P1_U3086), .B2(n5626), .C1(
        n9730), .C2(n9729), .ZN(P1_U3326) );
  INV_X1 U10926 ( .A(n9733), .ZN(n9734) );
  MUX2_X1 U10927 ( .A(n9734), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U10928 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9749) );
  AOI21_X1 U10929 ( .B1(n9737), .B2(n9736), .A(n9735), .ZN(n9738) );
  NAND2_X1 U10930 ( .A1(n9885), .A2(n9738), .ZN(n9744) );
  AOI21_X1 U10931 ( .B1(n9741), .B2(n9740), .A(n9739), .ZN(n9742) );
  NAND2_X1 U10932 ( .A1(n9893), .A2(n9742), .ZN(n9743) );
  OAI211_X1 U10933 ( .C1(n9899), .C2(n9745), .A(n9744), .B(n9743), .ZN(n9746)
         );
  INV_X1 U10934 ( .A(n9746), .ZN(n9748) );
  OAI211_X1 U10935 ( .C1(n9905), .C2(n9749), .A(n9748), .B(n9747), .ZN(
        P1_U3253) );
  INV_X1 U10936 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9763) );
  INV_X1 U10937 ( .A(n9750), .ZN(n9751) );
  OAI211_X1 U10938 ( .C1(n9753), .C2(n9752), .A(n9885), .B(n9751), .ZN(n9758)
         );
  OAI211_X1 U10939 ( .C1(n9756), .C2(n9755), .A(n9893), .B(n9754), .ZN(n9757)
         );
  OAI211_X1 U10940 ( .C1(n9899), .C2(n9759), .A(n9758), .B(n9757), .ZN(n9760)
         );
  INV_X1 U10941 ( .A(n9760), .ZN(n9762) );
  OAI211_X1 U10942 ( .C1(n9905), .C2(n9763), .A(n9762), .B(n9761), .ZN(
        P1_U3251) );
  INV_X1 U10943 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9779) );
  INV_X1 U10944 ( .A(n9764), .ZN(n9775) );
  OAI21_X1 U10945 ( .B1(n9767), .B2(n9766), .A(n9765), .ZN(n9768) );
  NAND2_X1 U10946 ( .A1(n9768), .A2(n9893), .ZN(n9774) );
  OAI21_X1 U10947 ( .B1(n9771), .B2(n9770), .A(n9769), .ZN(n9772) );
  NAND2_X1 U10948 ( .A1(n9885), .A2(n9772), .ZN(n9773) );
  OAI211_X1 U10949 ( .C1(n9899), .C2(n9775), .A(n9774), .B(n9773), .ZN(n9776)
         );
  INV_X1 U10950 ( .A(n9776), .ZN(n9778) );
  OAI211_X1 U10951 ( .C1(n9905), .C2(n9779), .A(n9778), .B(n9777), .ZN(
        P1_U3252) );
  INV_X1 U10952 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n9781) );
  AOI22_X1 U10953 ( .A1(n10091), .A2(n9781), .B1(n9780), .B2(n10088), .ZN(
        P2_U3458) );
  OAI22_X1 U10954 ( .A1(n10088), .A2(P2_REG0_REG_30__SCAN_IN), .B1(n9782), 
        .B2(n10091), .ZN(n9783) );
  INV_X1 U10955 ( .A(n9783), .ZN(P2_U3457) );
  INV_X1 U10956 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9785) );
  AOI22_X1 U10957 ( .A1(n10091), .A2(n9785), .B1(n9784), .B2(n10088), .ZN(
        P2_U3429) );
  XOR2_X1 U10958 ( .A(n9786), .B(P1_WR_REG_SCAN_IN), .Z(U123) );
  XOR2_X1 U10959 ( .A(n4717), .B(P1_RD_REG_SCAN_IN), .Z(U126) );
  OAI21_X1 U10960 ( .B1(n9788), .B2(P1_REG1_REG_0__SCAN_IN), .A(n9787), .ZN(
        n9790) );
  XNOR2_X1 U10961 ( .A(n9790), .B(n9789), .ZN(n9793) );
  AOI22_X1 U10962 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n9870), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9791) );
  OAI21_X1 U10963 ( .B1(n9793), .B2(n9792), .A(n9791), .ZN(P1_U3243) );
  INV_X1 U10964 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9806) );
  OAI211_X1 U10965 ( .C1(n9796), .C2(n9795), .A(n9885), .B(n9794), .ZN(n9801)
         );
  OAI211_X1 U10966 ( .C1(n9799), .C2(n9798), .A(n9893), .B(n9797), .ZN(n9800)
         );
  OAI211_X1 U10967 ( .C1(n9899), .C2(n9802), .A(n9801), .B(n9800), .ZN(n9803)
         );
  INV_X1 U10968 ( .A(n9803), .ZN(n9805) );
  OAI211_X1 U10969 ( .C1(n9905), .C2(n9806), .A(n9805), .B(n9804), .ZN(
        P1_U3249) );
  INV_X1 U10970 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9821) );
  AOI21_X1 U10971 ( .B1(n9809), .B2(n9808), .A(n9807), .ZN(n9810) );
  NAND2_X1 U10972 ( .A1(n9885), .A2(n9810), .ZN(n9816) );
  AOI21_X1 U10973 ( .B1(n9813), .B2(n9812), .A(n9811), .ZN(n9814) );
  NAND2_X1 U10974 ( .A1(n9893), .A2(n9814), .ZN(n9815) );
  OAI211_X1 U10975 ( .C1(n9899), .C2(n9817), .A(n9816), .B(n9815), .ZN(n9818)
         );
  INV_X1 U10976 ( .A(n9818), .ZN(n9820) );
  OAI211_X1 U10977 ( .C1(n9905), .C2(n9821), .A(n9820), .B(n9819), .ZN(
        P1_U3254) );
  INV_X1 U10978 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9834) );
  AOI211_X1 U10979 ( .C1(n9824), .C2(n9823), .A(n9822), .B(n9851), .ZN(n9829)
         );
  AOI211_X1 U10980 ( .C1(n9827), .C2(n9826), .A(n9825), .B(n9890), .ZN(n9828)
         );
  AOI211_X1 U10981 ( .C1(n9882), .C2(n9830), .A(n9829), .B(n9828), .ZN(n9833)
         );
  INV_X1 U10982 ( .A(n9831), .ZN(n9832) );
  OAI211_X1 U10983 ( .C1(n9905), .C2(n9834), .A(n9833), .B(n9832), .ZN(
        P1_U3256) );
  INV_X1 U10984 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9850) );
  INV_X1 U10985 ( .A(n9835), .ZN(n9846) );
  AOI21_X1 U10986 ( .B1(n9838), .B2(n9837), .A(n9836), .ZN(n9839) );
  NAND2_X1 U10987 ( .A1(n9885), .A2(n9839), .ZN(n9845) );
  AOI21_X1 U10988 ( .B1(n9842), .B2(n9841), .A(n9840), .ZN(n9843) );
  NAND2_X1 U10989 ( .A1(n9893), .A2(n9843), .ZN(n9844) );
  OAI211_X1 U10990 ( .C1(n9899), .C2(n9846), .A(n9845), .B(n9844), .ZN(n9847)
         );
  INV_X1 U10991 ( .A(n9847), .ZN(n9849) );
  OAI211_X1 U10992 ( .C1(n9905), .C2(n9850), .A(n9849), .B(n9848), .ZN(
        P1_U3257) );
  AOI211_X1 U10993 ( .C1(n9854), .C2(n9853), .A(n9852), .B(n9851), .ZN(n9859)
         );
  AOI211_X1 U10994 ( .C1(n9857), .C2(n9856), .A(n9855), .B(n9890), .ZN(n9858)
         );
  AOI211_X1 U10995 ( .C1(n9882), .C2(n9860), .A(n9859), .B(n9858), .ZN(n9861)
         );
  INV_X1 U10996 ( .A(n9861), .ZN(n9863) );
  AOI211_X1 U10997 ( .C1(n9870), .C2(P1_ADDR_REG_15__SCAN_IN), .A(n9863), .B(
        n9862), .ZN(n9864) );
  INV_X1 U10998 ( .A(n9864), .ZN(P1_U3258) );
  AOI211_X1 U10999 ( .C1(n9867), .C2(n9866), .A(n9865), .B(n9890), .ZN(n9868)
         );
  AOI211_X1 U11000 ( .C1(n9870), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n9869), .B(
        n9868), .ZN(n9877) );
  OAI21_X1 U11001 ( .B1(n9873), .B2(n9872), .A(n9871), .ZN(n9875) );
  AOI22_X1 U11002 ( .A1(n9875), .A2(n9893), .B1(n9874), .B2(n9882), .ZN(n9876)
         );
  NAND2_X1 U11003 ( .A1(n9877), .A2(n9876), .ZN(P1_U3259) );
  XNOR2_X1 U11004 ( .A(n9879), .B(n9878), .ZN(n9886) );
  XNOR2_X1 U11005 ( .A(n9881), .B(n9880), .ZN(n9884) );
  AOI222_X1 U11006 ( .A1(n9886), .A2(n9885), .B1(n9893), .B2(n9884), .C1(n9883), .C2(n9882), .ZN(n9888) );
  OAI211_X1 U11007 ( .C1(n9905), .C2(n9889), .A(n9888), .B(n9887), .ZN(
        P1_U3260) );
  AOI21_X1 U11008 ( .B1(n9892), .B2(n9891), .A(n9890), .ZN(n9902) );
  OAI211_X1 U11009 ( .C1(n9896), .C2(n9895), .A(n9894), .B(n9893), .ZN(n9897)
         );
  OAI21_X1 U11010 ( .B1(n9899), .B2(n9898), .A(n9897), .ZN(n9900) );
  AOI21_X1 U11011 ( .B1(n9902), .B2(n9901), .A(n9900), .ZN(n9904) );
  OAI211_X1 U11012 ( .C1(n9905), .C2(n10098), .A(n9904), .B(n9903), .ZN(
        P1_U3261) );
  OAI211_X1 U11013 ( .C1(n4687), .C2(n9908), .A(n9907), .B(n9906), .ZN(n9912)
         );
  AOI22_X1 U11014 ( .A1(n9932), .A2(n9910), .B1(n9909), .B2(n7513), .ZN(n9911)
         );
  AND2_X1 U11015 ( .A1(n9912), .A2(n9911), .ZN(n9998) );
  AOI222_X1 U11016 ( .A1(n9914), .A2(n9939), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n9593), .C1(n9952), .C2(n9913), .ZN(n9921) );
  XNOR2_X1 U11017 ( .A(n9916), .B(n9915), .ZN(n10001) );
  INV_X1 U11018 ( .A(n9917), .ZN(n9918) );
  OAI211_X1 U11019 ( .C1(n9999), .C2(n4437), .A(n9918), .B(n9942), .ZN(n9997)
         );
  INV_X1 U11020 ( .A(n9997), .ZN(n9919) );
  AOI22_X1 U11021 ( .A1(n10001), .A2(n9959), .B1(n9949), .B2(n9919), .ZN(n9920) );
  OAI211_X1 U11022 ( .C1(n9593), .C2(n9998), .A(n9921), .B(n9920), .ZN(
        P1_U3281) );
  XNOR2_X1 U11023 ( .A(n9940), .B(n9922), .ZN(n9928) );
  INV_X1 U11024 ( .A(n9928), .ZN(n9923) );
  XNOR2_X1 U11025 ( .A(n9924), .B(n9923), .ZN(n9985) );
  INV_X1 U11026 ( .A(n9925), .ZN(n9926) );
  NOR2_X1 U11027 ( .A1(n9927), .A2(n9926), .ZN(n9929) );
  XNOR2_X1 U11028 ( .A(n9929), .B(n9928), .ZN(n9935) );
  AOI22_X1 U11029 ( .A1(n9932), .A2(n9931), .B1(n9930), .B2(n7513), .ZN(n9933)
         );
  OAI21_X1 U11030 ( .B1(n9935), .B2(n9934), .A(n9933), .ZN(n9936) );
  AOI21_X1 U11031 ( .B1(n9937), .B2(n9985), .A(n9936), .ZN(n9982) );
  AOI222_X1 U11032 ( .A1(n9940), .A2(n9939), .B1(n9938), .B2(n9952), .C1(
        P1_REG2_REG_8__SCAN_IN), .C2(n9593), .ZN(n9948) );
  INV_X1 U11033 ( .A(n9941), .ZN(n9943) );
  OAI211_X1 U11034 ( .C1(n9981), .C2(n9944), .A(n9943), .B(n9942), .ZN(n9980)
         );
  INV_X1 U11035 ( .A(n9980), .ZN(n9945) );
  AOI22_X1 U11036 ( .A1(n9985), .A2(n9946), .B1(n9949), .B2(n9945), .ZN(n9947)
         );
  OAI211_X1 U11037 ( .C1(n9593), .C2(n9982), .A(n9948), .B(n9947), .ZN(
        P1_U3285) );
  NAND2_X1 U11038 ( .A1(n9950), .A2(n9949), .ZN(n9954) );
  AOI22_X1 U11039 ( .A1(n9593), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9952), .B2(
        n9951), .ZN(n9953) );
  OAI211_X1 U11040 ( .C1(n9956), .C2(n9955), .A(n9954), .B(n9953), .ZN(n9957)
         );
  AOI21_X1 U11041 ( .B1(n9959), .B2(n9958), .A(n9957), .ZN(n9960) );
  OAI21_X1 U11042 ( .B1(n9576), .B2(n9961), .A(n9960), .ZN(P1_U3290) );
  AND2_X1 U11043 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n4349), .ZN(P1_U3294) );
  AND2_X1 U11044 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n4349), .ZN(P1_U3295) );
  AND2_X1 U11045 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n4349), .ZN(P1_U3296) );
  AND2_X1 U11046 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n4349), .ZN(P1_U3297) );
  AND2_X1 U11047 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n4349), .ZN(P1_U3298) );
  AND2_X1 U11048 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n4349), .ZN(P1_U3299) );
  AND2_X1 U11049 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n4349), .ZN(P1_U3300) );
  AND2_X1 U11050 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n4349), .ZN(P1_U3301) );
  AND2_X1 U11051 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n4349), .ZN(P1_U3302) );
  AND2_X1 U11052 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n4349), .ZN(P1_U3303) );
  AND2_X1 U11053 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n4349), .ZN(P1_U3304) );
  AND2_X1 U11054 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n4349), .ZN(P1_U3305) );
  AND2_X1 U11055 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n4349), .ZN(P1_U3306) );
  AND2_X1 U11056 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n4349), .ZN(P1_U3307) );
  AND2_X1 U11057 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n4349), .ZN(P1_U3308) );
  AND2_X1 U11058 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n4349), .ZN(P1_U3309) );
  AND2_X1 U11059 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n4349), .ZN(P1_U3310) );
  AND2_X1 U11060 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n4349), .ZN(P1_U3311) );
  AND2_X1 U11061 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n4349), .ZN(P1_U3312) );
  AND2_X1 U11062 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n4349), .ZN(P1_U3313) );
  AND2_X1 U11063 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n4349), .ZN(P1_U3314) );
  AND2_X1 U11064 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n4349), .ZN(P1_U3315) );
  AND2_X1 U11065 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n4349), .ZN(P1_U3316) );
  AND2_X1 U11066 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n4349), .ZN(P1_U3317) );
  AND2_X1 U11067 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n4349), .ZN(P1_U3318) );
  AND2_X1 U11068 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n4349), .ZN(P1_U3319) );
  AND2_X1 U11069 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n4349), .ZN(P1_U3320) );
  AND2_X1 U11070 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n4349), .ZN(P1_U3321) );
  AND2_X1 U11071 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n4349), .ZN(P1_U3322) );
  AND2_X1 U11072 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n4349), .ZN(P1_U3323) );
  AOI22_X1 U11073 ( .A1(n10010), .A2(n9963), .B1(n5662), .B2(n10009), .ZN(
        P1_U3453) );
  OAI21_X1 U11074 ( .B1(n9965), .B2(n10004), .A(n9964), .ZN(n9967) );
  AOI211_X1 U11075 ( .C1(n10007), .C2(n9968), .A(n9967), .B(n9966), .ZN(n10012) );
  AOI22_X1 U11076 ( .A1(n10010), .A2(n10012), .B1(n5676), .B2(n10009), .ZN(
        P1_U3459) );
  OAI21_X1 U11077 ( .B1(n9970), .B2(n10004), .A(n9969), .ZN(n9972) );
  AOI211_X1 U11078 ( .C1(n10007), .C2(n9973), .A(n9972), .B(n9971), .ZN(n10013) );
  AOI22_X1 U11079 ( .A1(n10010), .A2(n10013), .B1(n5702), .B2(n10009), .ZN(
        P1_U3465) );
  OAI21_X1 U11080 ( .B1(n9975), .B2(n10004), .A(n9974), .ZN(n9977) );
  AOI211_X1 U11081 ( .C1(n10007), .C2(n9978), .A(n9977), .B(n9976), .ZN(n10014) );
  AOI22_X1 U11082 ( .A1(n10010), .A2(n10014), .B1(n5734), .B2(n10009), .ZN(
        P1_U3471) );
  INV_X1 U11083 ( .A(n9979), .ZN(n9986) );
  OAI21_X1 U11084 ( .B1(n9981), .B2(n10004), .A(n9980), .ZN(n9984) );
  INV_X1 U11085 ( .A(n9982), .ZN(n9983) );
  AOI211_X1 U11086 ( .C1(n9986), .C2(n9985), .A(n9984), .B(n9983), .ZN(n10015)
         );
  AOI22_X1 U11087 ( .A1(n10010), .A2(n10015), .B1(n5764), .B2(n10009), .ZN(
        P1_U3477) );
  OAI211_X1 U11088 ( .C1(n9989), .C2(n10004), .A(n9988), .B(n9987), .ZN(n9990)
         );
  AOI21_X1 U11089 ( .B1(n10007), .B2(n9991), .A(n9990), .ZN(n10016) );
  AOI22_X1 U11090 ( .A1(n10010), .A2(n10016), .B1(n5780), .B2(n10009), .ZN(
        P1_U3480) );
  OAI21_X1 U11091 ( .B1(n9993), .B2(n10004), .A(n9992), .ZN(n9994) );
  AOI211_X1 U11092 ( .C1(n9996), .C2(n10007), .A(n9995), .B(n9994), .ZN(n10017) );
  AOI22_X1 U11093 ( .A1(n10010), .A2(n10017), .B1(n5793), .B2(n10009), .ZN(
        P1_U3483) );
  OAI211_X1 U11094 ( .C1(n9999), .C2(n10004), .A(n9998), .B(n9997), .ZN(n10000) );
  AOI21_X1 U11095 ( .B1(n10001), .B2(n10007), .A(n10000), .ZN(n10018) );
  AOI22_X1 U11096 ( .A1(n10010), .A2(n10018), .B1(n5823), .B2(n10009), .ZN(
        P1_U3489) );
  OAI211_X1 U11097 ( .C1(n10005), .C2(n10004), .A(n10003), .B(n10002), .ZN(
        n10006) );
  AOI21_X1 U11098 ( .B1(n10008), .B2(n10007), .A(n10006), .ZN(n10020) );
  AOI22_X1 U11099 ( .A1(n10010), .A2(n10020), .B1(n5835), .B2(n10009), .ZN(
        P1_U3492) );
  AOI22_X1 U11100 ( .A1(n10021), .A2(n10012), .B1(n10011), .B2(n10019), .ZN(
        P1_U3524) );
  AOI22_X1 U11101 ( .A1(n10021), .A2(n10013), .B1(n5698), .B2(n10019), .ZN(
        P1_U3526) );
  AOI22_X1 U11102 ( .A1(n10021), .A2(n10014), .B1(n6763), .B2(n10019), .ZN(
        P1_U3528) );
  AOI22_X1 U11103 ( .A1(n10021), .A2(n10015), .B1(n5763), .B2(n10019), .ZN(
        P1_U3530) );
  AOI22_X1 U11104 ( .A1(n10021), .A2(n10016), .B1(n5779), .B2(n10019), .ZN(
        P1_U3531) );
  AOI22_X1 U11105 ( .A1(n10021), .A2(n10017), .B1(n6750), .B2(n10019), .ZN(
        P1_U3532) );
  AOI22_X1 U11106 ( .A1(n10021), .A2(n10018), .B1(n5822), .B2(n10019), .ZN(
        P1_U3534) );
  AOI22_X1 U11107 ( .A1(n10021), .A2(n10020), .B1(n9364), .B2(n10019), .ZN(
        P1_U3535) );
  OAI22_X1 U11108 ( .A1(n10023), .A2(n10022), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10063), .ZN(n10035) );
  AOI21_X1 U11109 ( .B1(n10026), .B2(n10025), .A(n10024), .ZN(n10033) );
  OAI21_X1 U11110 ( .B1(n10029), .B2(n10028), .A(n10027), .ZN(n10030) );
  NAND2_X1 U11111 ( .A1(n10056), .A2(n10030), .ZN(n10031) );
  OAI21_X1 U11112 ( .B1(n10033), .B2(n10032), .A(n10031), .ZN(n10034) );
  AOI211_X1 U11113 ( .C1(n10045), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n10035), .B(
        n10034), .ZN(n10040) );
  XOR2_X1 U11114 ( .A(n10037), .B(n10036), .Z(n10038) );
  NAND2_X1 U11115 ( .A1(n10038), .A2(n10051), .ZN(n10039) );
  NAND2_X1 U11116 ( .A1(n10040), .A2(n10039), .ZN(P2_U3184) );
  OAI21_X1 U11117 ( .B1(n10042), .B2(P2_REG1_REG_3__SCAN_IN), .A(n10041), .ZN(
        n10044) );
  AOI222_X1 U11118 ( .A1(n10047), .A2(n10046), .B1(n10045), .B2(
        P2_ADDR_REG_3__SCAN_IN), .C1(n10044), .C2(n10043), .ZN(n10060) );
  OAI21_X1 U11119 ( .B1(n10050), .B2(n10049), .A(n10048), .ZN(n10052) );
  NAND2_X1 U11120 ( .A1(n10052), .A2(n10051), .ZN(n10058) );
  OAI21_X1 U11121 ( .B1(n10054), .B2(P2_REG2_REG_3__SCAN_IN), .A(n10053), .ZN(
        n10055) );
  NAND2_X1 U11122 ( .A1(n10056), .A2(n10055), .ZN(n10057) );
  NAND4_X1 U11123 ( .A1(n10060), .A2(n10059), .A3(n10058), .A4(n10057), .ZN(
        P2_U3185) );
  OAI22_X1 U11124 ( .A1(n10064), .A2(n10063), .B1(n10062), .B2(n10061), .ZN(
        n10066) );
  AOI211_X1 U11125 ( .C1(n10068), .C2(n10067), .A(n10066), .B(n10065), .ZN(
        n10070) );
  AOI22_X1 U11126 ( .A1(n8734), .A2(n5083), .B1(n10070), .B2(n10069), .ZN(
        P2_U3231) );
  INV_X1 U11127 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10072) );
  AOI22_X1 U11128 ( .A1(n10091), .A2(n10072), .B1(n10071), .B2(n10088), .ZN(
        P2_U3390) );
  INV_X1 U11129 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10074) );
  AOI22_X1 U11130 ( .A1(n10091), .A2(n10074), .B1(n10073), .B2(n10088), .ZN(
        P2_U3396) );
  AOI22_X1 U11131 ( .A1(n10091), .A2(n5119), .B1(n10075), .B2(n10088), .ZN(
        P2_U3402) );
  INV_X1 U11132 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10077) );
  AOI22_X1 U11133 ( .A1(n10091), .A2(n10077), .B1(n10076), .B2(n10088), .ZN(
        P2_U3405) );
  INV_X1 U11134 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10079) );
  AOI22_X1 U11135 ( .A1(n10091), .A2(n10079), .B1(n10078), .B2(n10088), .ZN(
        P2_U3408) );
  INV_X1 U11136 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10081) );
  AOI22_X1 U11137 ( .A1(n10091), .A2(n10081), .B1(n10080), .B2(n10088), .ZN(
        P2_U3414) );
  INV_X1 U11138 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10083) );
  AOI22_X1 U11139 ( .A1(n10091), .A2(n10083), .B1(n10082), .B2(n10088), .ZN(
        P2_U3417) );
  INV_X1 U11140 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10085) );
  AOI22_X1 U11141 ( .A1(n10091), .A2(n10085), .B1(n10084), .B2(n10088), .ZN(
        P2_U3420) );
  INV_X1 U11142 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10087) );
  AOI22_X1 U11143 ( .A1(n10091), .A2(n10087), .B1(n10086), .B2(n10088), .ZN(
        P2_U3423) );
  INV_X1 U11144 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10090) );
  AOI22_X1 U11145 ( .A1(n10091), .A2(n10090), .B1(n10089), .B2(n10088), .ZN(
        P2_U3426) );
  OAI222_X1 U11146 ( .A1(n10096), .A2(n10095), .B1(n10096), .B2(n10094), .C1(
        n10093), .C2(n10092), .ZN(ADD_1068_U5) );
  XOR2_X1 U11147 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  AOI21_X1 U11148 ( .B1(n10099), .B2(n10098), .A(n10097), .ZN(n10100) );
  XOR2_X1 U11149 ( .A(n10100), .B(P2_ADDR_REG_18__SCAN_IN), .Z(ADD_1068_U55)
         );
  OAI21_X1 U11150 ( .B1(n10103), .B2(n10102), .A(n10101), .ZN(ADD_1068_U56) );
  OAI21_X1 U11151 ( .B1(n10106), .B2(n10105), .A(n10104), .ZN(ADD_1068_U57) );
  OAI21_X1 U11152 ( .B1(n10109), .B2(n10108), .A(n10107), .ZN(ADD_1068_U58) );
  OAI21_X1 U11153 ( .B1(n10112), .B2(n10111), .A(n10110), .ZN(ADD_1068_U59) );
  OAI21_X1 U11154 ( .B1(n10115), .B2(n10114), .A(n10113), .ZN(ADD_1068_U60) );
  OAI21_X1 U11155 ( .B1(n10118), .B2(n10117), .A(n10116), .ZN(ADD_1068_U61) );
  OAI21_X1 U11156 ( .B1(n10121), .B2(n10120), .A(n10119), .ZN(ADD_1068_U62) );
  OAI21_X1 U11157 ( .B1(n10124), .B2(n10123), .A(n10122), .ZN(ADD_1068_U63) );
  AOI21_X1 U11158 ( .B1(n10127), .B2(n10126), .A(n10125), .ZN(ADD_1068_U54) );
  OAI21_X1 U11159 ( .B1(n10130), .B2(n10129), .A(n10128), .ZN(ADD_1068_U47) );
  OAI21_X1 U11160 ( .B1(n10133), .B2(n10132), .A(n10131), .ZN(ADD_1068_U48) );
  OAI21_X1 U11161 ( .B1(n10136), .B2(n10135), .A(n10134), .ZN(ADD_1068_U49) );
  OAI21_X1 U11162 ( .B1(n10139), .B2(n10138), .A(n10137), .ZN(ADD_1068_U50) );
  OAI21_X1 U11163 ( .B1(n10142), .B2(n10141), .A(n10140), .ZN(ADD_1068_U51) );
  AOI21_X1 U11164 ( .B1(n10145), .B2(n10144), .A(n10143), .ZN(ADD_1068_U53) );
  OAI21_X1 U11165 ( .B1(n10148), .B2(n10147), .A(n10146), .ZN(ADD_1068_U52) );
  CLKBUF_X1 U4862 ( .A(n5188), .Z(n6661) );
  CLKBUF_X1 U4876 ( .A(n5701), .Z(n5963) );
  AND2_X1 U4950 ( .A1(n9719), .A2(n9718), .ZN(n10152) );
endmodule

