

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput127, keyinput126, keyinput125, keyinput124, keyinput123, 
        keyinput122, keyinput121, keyinput120, keyinput119, keyinput118, 
        keyinput117, keyinput116, keyinput115, keyinput114, keyinput113, 
        keyinput112, keyinput111, keyinput110, keyinput109, keyinput108, 
        keyinput107, keyinput106, keyinput105, keyinput104, keyinput103, 
        keyinput102, keyinput101, keyinput100, keyinput99, keyinput98, 
        keyinput97, keyinput96, keyinput95, keyinput94, keyinput93, keyinput92, 
        keyinput91, keyinput90, keyinput89, keyinput88, keyinput87, keyinput86, 
        keyinput85, keyinput84, keyinput83, keyinput82, keyinput81, keyinput80, 
        keyinput79, keyinput78, keyinput77, keyinput76, keyinput75, keyinput74, 
        keyinput73, keyinput72, keyinput71, keyinput70, keyinput69, keyinput68, 
        keyinput67, keyinput66, keyinput65, keyinput64, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347;

  INV_X4 U4896 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  AND2_X1 U4897 ( .A1(n4631), .A2(n4465), .ZN(n4629) );
  CLKBUF_X2 U4898 ( .A(n7551), .Z(n9065) );
  AND2_X1 U4900 ( .A1(n4391), .A2(n7813), .ZN(n5210) );
  OR2_X1 U4901 ( .A1(n5033), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n5032) );
  AND3_X1 U4902 ( .A1(n4985), .A2(n4984), .A3(n4988), .ZN(n4750) );
  NOR2_X1 U4903 ( .A1(n5946), .A2(n5706), .ZN(n4390) );
  NOR2_X1 U4904 ( .A1(n5946), .A2(n5706), .ZN(n5707) );
  AND2_X1 U4905 ( .A1(n5222), .A2(n4986), .ZN(n4751) );
  OR2_X1 U4906 ( .A1(n5593), .A2(n4595), .ZN(n4590) );
  INV_X2 U4907 ( .A(n5184), .ZN(n5460) );
  INV_X1 U4908 ( .A(n8186), .ZN(n8171) );
  AND2_X1 U4909 ( .A1(n4432), .A2(n4991), .ZN(n4794) );
  NAND2_X1 U4910 ( .A1(n5770), .A2(n7813), .ZN(n5768) );
  CLKBUF_X2 U4911 ( .A(n6197), .Z(n8280) );
  NAND3_X1 U4912 ( .A1(n4590), .A2(n4589), .A3(n4591), .ZN(n5002) );
  INV_X1 U4913 ( .A(n4979), .ZN(n5763) );
  CLKBUF_X2 U4915 ( .A(n5770), .Z(n6361) );
  NAND2_X1 U4916 ( .A1(n4416), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6101) );
  NAND2_X1 U4917 ( .A1(n5001), .A2(n5002), .ZN(n5184) );
  NAND2_X1 U4918 ( .A1(n5032), .A2(n4969), .ZN(n5037) );
  OR2_X1 U4919 ( .A1(n8542), .A2(n10220), .ZN(n4855) );
  INV_X1 U4920 ( .A(n5850), .ZN(n4914) );
  NAND2_X2 U4921 ( .A1(n5496), .A2(n8657), .ZN(n8646) );
  OAI21_X2 U4922 ( .B1(n7915), .B2(n7904), .A(n7903), .ZN(n7908) );
  NAND2_X2 U4923 ( .A1(n9157), .A2(n8982), .ZN(n9035) );
  AND2_X2 U4924 ( .A1(n8042), .A2(n8040), .ZN(n8212) );
  NAND2_X2 U4925 ( .A1(n5037), .A2(n5036), .ZN(n7745) );
  XNOR2_X2 U4926 ( .A(n6101), .B(P1_IR_REG_21__SCAN_IN), .ZN(n7757) );
  NAND2_X1 U4927 ( .A1(n5001), .A2(n5002), .ZN(n4391) );
  AND2_X4 U4928 ( .A1(n5054), .A2(n5053), .ZN(n5062) );
  NAND2_X1 U4929 ( .A1(n5041), .A2(n7745), .ZN(n4392) );
  NAND2_X1 U4930 ( .A1(n5041), .A2(n7745), .ZN(n4393) );
  NAND2_X1 U4931 ( .A1(n5041), .A2(n7745), .ZN(n5200) );
  INV_X2 U4932 ( .A(n8413), .ZN(n6845) );
  INV_X1 U4933 ( .A(n7950), .ZN(n7947) );
  INV_X4 U4934 ( .A(n7541), .ZN(n4394) );
  CLKBUF_X2 U4935 ( .A(n5800), .Z(n6072) );
  CLKBUF_X2 U4936 ( .A(n5191), .Z(n5435) );
  BUF_X2 U4937 ( .A(n5190), .Z(n8179) );
  NAND2_X1 U4938 ( .A1(n4907), .A2(n4906), .ZN(n5683) );
  NOR2_X1 U4939 ( .A1(n8261), .A2(n8651), .ZN(n8346) );
  NAND2_X1 U4940 ( .A1(n4909), .A2(n4908), .ZN(n4907) );
  NAND2_X1 U4941 ( .A1(n9137), .A2(n8995), .ZN(n9106) );
  AOI21_X1 U4942 ( .B1(n4880), .B2(n4879), .A(n8006), .ZN(n4874) );
  AOI21_X1 U4943 ( .B1(n8592), .B2(n8584), .A(n8152), .ZN(n5674) );
  XNOR2_X1 U4944 ( .A(n8512), .B(n10214), .ZN(n10219) );
  OAI21_X1 U4945 ( .B1(n7935), .B2(n7942), .A(n7934), .ZN(n7936) );
  OAI21_X1 U4946 ( .B1(n7943), .B2(n7942), .A(n4435), .ZN(n4684) );
  OR2_X1 U4947 ( .A1(n8637), .A2(n8135), .ZN(n8624) );
  NOR2_X1 U4948 ( .A1(n7982), .A2(n7985), .ZN(n4881) );
  NOR2_X1 U4949 ( .A1(n10216), .A2(n10217), .ZN(n10215) );
  XNOR2_X1 U4950 ( .A(n4820), .B(n8517), .ZN(n10216) );
  NAND2_X1 U4951 ( .A1(n8843), .A2(n8607), .ZN(n4906) );
  OR2_X1 U4952 ( .A1(n8532), .A2(n4484), .ZN(n4820) );
  NOR2_X1 U4953 ( .A1(n8504), .A2(n8503), .ZN(n8532) );
  NAND2_X1 U4954 ( .A1(n6284), .A2(n8400), .ZN(n4908) );
  NOR2_X1 U4955 ( .A1(n8500), .A2(n8501), .ZN(n8504) );
  AND2_X1 U4956 ( .A1(n4829), .A2(n4425), .ZN(n8442) );
  AND2_X1 U4957 ( .A1(n8430), .A2(n8429), .ZN(n8438) );
  OR2_X1 U4958 ( .A1(n7415), .A2(n7414), .ZN(n8430) );
  AND2_X1 U4959 ( .A1(n4735), .A2(n7549), .ZN(n4734) );
  NAND2_X1 U4960 ( .A1(n4454), .A2(n4403), .ZN(n4738) );
  NAND2_X1 U4961 ( .A1(n4886), .A2(n4436), .ZN(n7216) );
  NAND2_X1 U4962 ( .A1(n5361), .A2(n5360), .ZN(n10282) );
  NOR2_X1 U4963 ( .A1(n6634), .A2(n6633), .ZN(n6698) );
  INV_X1 U4964 ( .A(n7185), .ZN(n7176) );
  XNOR2_X1 U4965 ( .A(n5300), .B(n5299), .ZN(n6346) );
  INV_X1 U4966 ( .A(n8212), .ZN(n6839) );
  CLKBUF_X1 U4967 ( .A(n6573), .Z(n6594) );
  NAND4_X1 U4968 ( .A1(n5767), .A2(n5766), .A3(n5765), .A4(n5764), .ZN(n5784)
         );
  OR2_X1 U4969 ( .A1(n5817), .A2(n5816), .ZN(n9228) );
  NOR2_X2 U4970 ( .A1(n6287), .A2(n8186), .ZN(n5047) );
  INV_X2 U4971 ( .A(n5863), .ZN(n7818) );
  NAND2_X1 U4973 ( .A1(n5732), .A2(n9960), .ZN(n7744) );
  XNOR2_X1 U4974 ( .A(n5720), .B(n9809), .ZN(n9342) );
  OR2_X1 U4975 ( .A1(n4392), .A2(n6849), .ZN(n5180) );
  NAND2_X1 U4976 ( .A1(n4809), .A2(n5726), .ZN(n5732) );
  XNOR2_X1 U4977 ( .A(n5459), .B(n9797), .ZN(n8555) );
  NAND2_X1 U4978 ( .A1(n4527), .A2(n5059), .ZN(n5207) );
  XNOR2_X1 U4979 ( .A(n5006), .B(n4795), .ZN(n8241) );
  NAND2_X1 U4980 ( .A1(n8914), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5039) );
  NOR2_X1 U4981 ( .A1(n5430), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n4622) );
  XNOR2_X1 U4982 ( .A(n5241), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6657) );
  NAND2_X1 U4983 ( .A1(n4839), .A2(n4646), .ZN(n10203) );
  OR2_X1 U4984 ( .A1(n5256), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5272) );
  BUF_X2 U4985 ( .A(n5062), .Z(n7813) );
  AND4_X1 U4986 ( .A1(n4983), .A2(n4982), .A3(n4981), .A4(n4980), .ZN(n4398)
         );
  NOR2_X1 U4987 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n4982) );
  NOR2_X1 U4988 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n4983) );
  NOR2_X1 U4989 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5701) );
  INV_X1 U4990 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5038) );
  NOR2_X1 U4991 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5702) );
  INV_X4 U4992 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  AND2_X1 U4993 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n9971) );
  INV_X1 U4994 ( .A(P2_RD_REG_SCAN_IN), .ZN(n9795) );
  INV_X1 U4995 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5700) );
  NOR2_X2 U4996 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n4706) );
  INV_X1 U4997 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5222) );
  INV_X1 U4998 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4984) );
  NOR2_X1 U4999 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n4981) );
  NOR2_X2 U5000 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5204) );
  NOR2_X1 U5001 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n4980) );
  NAND2_X2 U5002 ( .A1(n6839), .A2(n6843), .ZN(n8758) );
  NOR2_X1 U5003 ( .A1(n4970), .A2(n4424), .ZN(n5203) );
  OAI211_X1 U5004 ( .C1(n5234), .C2(n8864), .A(n5514), .B(n5513), .ZN(n8651)
         );
  NAND2_X2 U5005 ( .A1(n5735), .A2(n5747), .ZN(n6131) );
  XNOR2_X2 U5006 ( .A(n5784), .B(n6106), .ZN(n6108) );
  NOR2_X2 U5007 ( .A1(n7255), .A2(n7455), .ZN(n7279) );
  INV_X1 U5008 ( .A(n4564), .ZN(n4560) );
  AOI21_X1 U5009 ( .B1(n4564), .B2(n4563), .A(n4562), .ZN(n4561) );
  INV_X1 U5010 ( .A(n5093), .ZN(n4562) );
  INV_X1 U5011 ( .A(n5088), .ZN(n4563) );
  INV_X1 U5012 ( .A(n8317), .ZN(n4774) );
  OR2_X1 U5013 ( .A1(n8901), .A2(n7644), .ZN(n8104) );
  NAND2_X1 U5014 ( .A1(n10154), .A2(n7552), .ZN(n4963) );
  AND2_X1 U5015 ( .A1(n5563), .A2(n5175), .ZN(n5561) );
  NAND2_X1 U5016 ( .A1(n4872), .A2(n5122), .ZN(n5428) );
  AOI21_X1 U5017 ( .B1(n4870), .B2(n4554), .A(n4452), .ZN(n4553) );
  INV_X1 U5018 ( .A(n8588), .ZN(n8156) );
  OR2_X1 U5019 ( .A1(n8304), .A2(n6230), .ZN(n4397) );
  INV_X1 U5020 ( .A(n5435), .ZN(n5574) );
  INV_X1 U5021 ( .A(n5200), .ZN(n5575) );
  AND4_X1 U5022 ( .A1(n5282), .A2(n5281), .A3(n5280), .A4(n5279), .ZN(n6215)
         );
  INV_X1 U5023 ( .A(n7744), .ZN(n5735) );
  INV_X1 U5024 ( .A(n6063), .ZN(n4922) );
  OAI21_X1 U5025 ( .B1(n9450), .B2(n6041), .A(n6042), .ZN(n9434) );
  AOI21_X1 U5026 ( .B1(n4580), .B2(n8210), .A(n4577), .ZN(n8095) );
  INV_X1 U5027 ( .A(n8638), .ZN(n4574) );
  INV_X1 U5028 ( .A(n8134), .ZN(n8136) );
  INV_X1 U5029 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4986) );
  NOR2_X1 U5030 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n4987) );
  NAND2_X1 U5031 ( .A1(n5678), .A2(n5677), .ZN(n7742) );
  NOR2_X1 U5032 ( .A1(n5454), .A2(n4867), .ZN(n4866) );
  INV_X1 U5033 ( .A(n5133), .ZN(n4867) );
  INV_X1 U5034 ( .A(n6250), .ZN(n4787) );
  OAI21_X1 U5035 ( .B1(n6560), .B2(n4832), .A(n4830), .ZN(n6659) );
  OR2_X1 U5036 ( .A1(n4836), .A2(n10291), .ZN(n4832) );
  INV_X1 U5037 ( .A(n4831), .ZN(n4830) );
  INV_X1 U5038 ( .A(n6756), .ZN(n4854) );
  INV_X1 U5039 ( .A(n6755), .ZN(n4850) );
  NAND2_X1 U5040 ( .A1(n6845), .A2(n10240), .ZN(n6853) );
  OR2_X1 U5041 ( .A1(n8859), .A2(n8614), .ZN(n8208) );
  OR2_X1 U5042 ( .A1(n8871), .A2(n8264), .ZN(n8129) );
  OR2_X1 U5043 ( .A1(n8883), .A2(n8693), .ZN(n8119) );
  INV_X1 U5044 ( .A(n4899), .ZN(n4898) );
  OAI21_X1 U5045 ( .B1(n7668), .B2(n4900), .A(n7666), .ZN(n4899) );
  NAND2_X1 U5046 ( .A1(n5370), .A2(n5369), .ZN(n4900) );
  OR2_X1 U5047 ( .A1(n10282), .A2(n7708), .ZN(n8030) );
  OR3_X1 U5048 ( .A1(n7532), .A2(n7530), .A3(n7531), .ZN(n4972) );
  INV_X1 U5049 ( .A(n6945), .ZN(n4723) );
  AND2_X1 U5050 ( .A1(n6606), .A2(n10092), .ZN(n6607) );
  NAND3_X1 U5051 ( .A1(n4968), .A2(n8007), .A3(n7009), .ZN(n6613) );
  AND2_X1 U5052 ( .A1(n6779), .A2(n6780), .ZN(n4724) );
  NOR2_X1 U5053 ( .A1(n9649), .A2(n9374), .ZN(n4879) );
  INV_X1 U5054 ( .A(n9213), .ZN(n9160) );
  NAND2_X1 U5055 ( .A1(n4511), .A2(n7765), .ZN(n4510) );
  AND2_X1 U5056 ( .A1(n6118), .A2(n4512), .ZN(n4511) );
  INV_X1 U5057 ( .A(n7964), .ZN(n4512) );
  NAND2_X1 U5058 ( .A1(n4954), .A2(n4953), .ZN(n7596) );
  AOI21_X1 U5059 ( .B1(n4404), .B2(n4957), .A(n4474), .ZN(n4953) );
  AND2_X1 U5060 ( .A1(n4542), .A2(n4540), .ZN(n4539) );
  INV_X1 U5061 ( .A(n5497), .ZN(n4540) );
  INV_X1 U5062 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5708) );
  NOR2_X1 U5063 ( .A1(n5117), .A2(n4871), .ZN(n4870) );
  INV_X1 U5064 ( .A(n5111), .ZN(n4871) );
  AOI21_X1 U5065 ( .B1(n4664), .B2(n4666), .A(n5372), .ZN(n4663) );
  OAI21_X1 U5066 ( .B1(n5300), .B2(n4560), .A(n4561), .ZN(n5323) );
  OAI21_X1 U5067 ( .B1(n5062), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n4528), .ZN(
        n5057) );
  NAND2_X1 U5068 ( .A1(n5062), .A2(n6331), .ZN(n4528) );
  XNOR2_X1 U5069 ( .A(n8288), .B(n8588), .ZN(n8279) );
  AND2_X1 U5070 ( .A1(n4774), .A2(n4765), .ZN(n4764) );
  NAND2_X1 U5071 ( .A1(n4766), .A2(n8318), .ZN(n4765) );
  INV_X1 U5072 ( .A(n8407), .ZN(n6219) );
  AND2_X1 U5073 ( .A1(n4778), .A2(n6233), .ZN(n4419) );
  OR2_X1 U5074 ( .A1(n4779), .A2(n4397), .ZN(n4778) );
  NOR2_X1 U5075 ( .A1(n6231), .A2(n4780), .ZN(n4779) );
  OR2_X1 U5076 ( .A1(n8183), .A2(n8288), .ZN(n4588) );
  INV_X1 U5077 ( .A(n8241), .ZN(n8204) );
  NOR2_X1 U5078 ( .A1(n8288), .A2(n8588), .ZN(n5682) );
  OR2_X1 U5079 ( .A1(n5501), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5511) );
  OAI21_X1 U5080 ( .B1(n8727), .B2(n5636), .A(n8104), .ZN(n8720) );
  OAI21_X1 U5081 ( .B1(n7191), .B2(n4606), .A(n4602), .ZN(n7474) );
  AOI21_X1 U5082 ( .B1(n4605), .B2(n4604), .A(n4603), .ZN(n4602) );
  INV_X1 U5083 ( .A(n8064), .ZN(n4603) );
  INV_X1 U5084 ( .A(n4611), .ZN(n4604) );
  AOI21_X1 U5085 ( .B1(n8056), .B2(n4611), .A(n4610), .ZN(n4609) );
  INV_X1 U5086 ( .A(n8078), .ZN(n4610) );
  INV_X1 U5087 ( .A(n5210), .ZN(n5290) );
  OR2_X1 U5088 ( .A1(n8889), .A2(n8357), .ZN(n8670) );
  INV_X1 U5089 ( .A(n5047), .ZN(n8762) );
  OR2_X1 U5090 ( .A1(n8894), .A2(n8692), .ZN(n8683) );
  INV_X1 U5091 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5588) );
  INV_X1 U5092 ( .A(n8997), .ZN(n9068) );
  AND2_X1 U5093 ( .A1(n4724), .A2(n4723), .ZN(n4717) );
  NAND2_X1 U5094 ( .A1(n4723), .A2(n4716), .ZN(n4715) );
  INV_X1 U5095 ( .A(n6944), .ZN(n4716) );
  INV_X1 U5096 ( .A(n6035), .ZN(n6033) );
  NAND2_X1 U5097 ( .A1(n6769), .A2(n6768), .ZN(n6803) );
  OR3_X1 U5098 ( .A1(n6992), .A2(n6602), .A3(n6601), .ZN(n6619) );
  OR2_X1 U5099 ( .A1(n8012), .A2(n7998), .ZN(n6603) );
  AND2_X1 U5100 ( .A1(n4718), .A2(n4715), .ZN(n4713) );
  NAND2_X1 U5101 ( .A1(n4722), .A2(n7096), .ZN(n4718) );
  OAI21_X1 U5102 ( .B1(n8001), .B2(n4532), .A(n4531), .ZN(n4530) );
  OAI21_X1 U5103 ( .B1(n8000), .B2(n4532), .A(n9342), .ZN(n4531) );
  NOR2_X1 U5104 ( .A1(n7983), .A2(n4533), .ZN(n4532) );
  AOI21_X1 U5105 ( .B1(n4878), .B2(n4652), .A(n4651), .ZN(n8001) );
  AND4_X1 U5106 ( .A1(n5899), .A2(n5898), .A3(n5897), .A4(n5896), .ZN(n7542)
         );
  NAND2_X1 U5107 ( .A1(n9590), .A2(n9209), .ZN(n4925) );
  NAND2_X1 U5108 ( .A1(n4921), .A2(n6064), .ZN(n4919) );
  INV_X1 U5109 ( .A(n4507), .ZN(n4506) );
  OAI21_X1 U5110 ( .B1(n4508), .B2(n7909), .A(n7910), .ZN(n4507) );
  OAI21_X1 U5111 ( .B1(n9468), .B2(n6030), .A(n6029), .ZN(n9450) );
  OR2_X1 U5112 ( .A1(n7561), .A2(n7552), .ZN(n7870) );
  INV_X1 U5113 ( .A(n7820), .ZN(n5986) );
  INV_X1 U5114 ( .A(n6361), .ZN(n5985) );
  NAND2_X1 U5115 ( .A1(n5770), .A2(n6325), .ZN(n5863) );
  XNOR2_X1 U5116 ( .A(n7817), .B(n7816), .ZN(n8912) );
  NAND2_X1 U5117 ( .A1(n7812), .A2(n7811), .ZN(n7817) );
  NAND2_X1 U5118 ( .A1(n4805), .A2(n4806), .ZN(n5734) );
  XNOR2_X1 U5119 ( .A(n5562), .B(n5561), .ZN(n7564) );
  NAND2_X1 U5120 ( .A1(n4862), .A2(n5171), .ZN(n5562) );
  XNOR2_X1 U5121 ( .A(n6140), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6167) );
  NOR2_X1 U5122 ( .A1(n6280), .A2(n6281), .ZN(n8277) );
  AND2_X1 U5123 ( .A1(n8182), .A2(n5051), .ZN(n8286) );
  OAI21_X1 U5124 ( .B1(n6210), .B2(n4793), .A(n4790), .ZN(n6218) );
  AOI21_X1 U5125 ( .B1(n4792), .B2(n7143), .A(n4791), .ZN(n4790) );
  INV_X1 U5126 ( .A(n7320), .ZN(n4791) );
  INV_X1 U5127 ( .A(n8400), .ZN(n8607) );
  OR2_X1 U5128 ( .A1(n8487), .A2(n8486), .ZN(n4645) );
  AND2_X1 U5129 ( .A1(n9342), .A2(n7108), .ZN(n8012) );
  AND2_X1 U5130 ( .A1(n4878), .A2(n4877), .ZN(n8009) );
  INV_X1 U5131 ( .A(n7836), .ZN(n4494) );
  INV_X1 U5132 ( .A(n7828), .ZN(n4496) );
  NAND2_X1 U5133 ( .A1(n8066), .A2(n8080), .ZN(n4582) );
  NAND2_X1 U5134 ( .A1(n4583), .A2(n4581), .ZN(n4580) );
  NAND2_X1 U5135 ( .A1(n4584), .A2(n8171), .ZN(n4583) );
  NAND2_X1 U5136 ( .A1(n4582), .A2(n8186), .ZN(n4581) );
  OAI21_X1 U5137 ( .B1(n8085), .B2(n8084), .A(n8083), .ZN(n4584) );
  AND2_X1 U5138 ( .A1(n4574), .A2(n4571), .ZN(n4570) );
  OR2_X1 U5139 ( .A1(n8125), .A2(n4572), .ZN(n4568) );
  OR2_X1 U5140 ( .A1(n9342), .A2(n7757), .ZN(n4968) );
  AND2_X1 U5141 ( .A1(n4678), .A2(n4677), .ZN(n7949) );
  INV_X1 U5142 ( .A(n7946), .ZN(n4677) );
  NAND2_X1 U5143 ( .A1(n5763), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5764) );
  NAND2_X1 U5144 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), 
        .ZN(n4595) );
  AND2_X1 U5145 ( .A1(n4993), .A2(n9810), .ZN(n4594) );
  OAI21_X1 U5146 ( .B1(n4993), .B2(n4595), .A(n4593), .ZN(n4592) );
  NAND2_X1 U5147 ( .A1(n8913), .A2(n9810), .ZN(n4593) );
  NAND2_X1 U5148 ( .A1(n6540), .A2(n6520), .ZN(n6522) );
  OR2_X1 U5149 ( .A1(n8288), .A2(n8156), .ZN(n4617) );
  AND2_X1 U5150 ( .A1(n4618), .A2(n8141), .ZN(n4615) );
  NOR2_X1 U5151 ( .A1(n5673), .A2(n8591), .ZN(n4618) );
  OR2_X1 U5152 ( .A1(n7314), .A2(n10267), .ZN(n8064) );
  OR2_X1 U5153 ( .A1(n7736), .A2(n7507), .ZN(n8097) );
  NAND2_X1 U5154 ( .A1(n5185), .A2(n10203), .ZN(n5186) );
  INV_X1 U5155 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4749) );
  INV_X1 U5156 ( .A(n4729), .ZN(n4728) );
  OAI21_X1 U5157 ( .B1(n9148), .B2(n4730), .A(n9098), .ZN(n4729) );
  INV_X1 U5158 ( .A(n8968), .ZN(n4730) );
  AND2_X1 U5159 ( .A1(n4403), .A2(n4478), .ZN(n4739) );
  NAND2_X1 U5160 ( .A1(n6945), .A2(n6944), .ZN(n4722) );
  AND2_X1 U5161 ( .A1(n9383), .A2(n9207), .ZN(n7945) );
  NOR2_X1 U5162 ( .A1(n9383), .A2(n9207), .ZN(n7944) );
  INV_X1 U5163 ( .A(n4800), .ZN(n4799) );
  OAI21_X1 U5164 ( .B1(n6128), .B2(n4801), .A(n9409), .ZN(n4800) );
  INV_X1 U5165 ( .A(n7794), .ZN(n4801) );
  NOR3_X1 U5166 ( .A1(n9452), .A2(n4700), .A3(n9389), .ZN(n4704) );
  NAND2_X1 U5167 ( .A1(n9663), .A2(n4703), .ZN(n4702) );
  NAND2_X1 U5168 ( .A1(n4929), .A2(n6009), .ZN(n4928) );
  INV_X1 U5169 ( .A(n4930), .ZN(n4929) );
  NOR2_X1 U5170 ( .A1(n9625), .A2(n9531), .ZN(n4697) );
  INV_X1 U5171 ( .A(n5995), .ZN(n4945) );
  NOR2_X1 U5172 ( .A1(n4395), .A2(n5995), .ZN(n4944) );
  INV_X1 U5173 ( .A(n6122), .ZN(n4812) );
  NAND2_X1 U5174 ( .A1(n4656), .A2(n4655), .ZN(n7893) );
  NAND2_X1 U5175 ( .A1(n9202), .A2(n8920), .ZN(n7891) );
  AND2_X1 U5176 ( .A1(n4815), .A2(n7880), .ZN(n4814) );
  INV_X1 U5177 ( .A(n7971), .ZN(n4815) );
  NOR2_X1 U5178 ( .A1(n4939), .A2(n4936), .ZN(n4935) );
  INV_X1 U5179 ( .A(n7840), .ZN(n4936) );
  INV_X1 U5180 ( .A(n7115), .ZN(n4939) );
  INV_X1 U5181 ( .A(n5866), .ZN(n4938) );
  INV_X1 U5182 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n9750) );
  OR2_X1 U5183 ( .A1(n7333), .A2(n7867), .ZN(n7967) );
  NOR2_X1 U5184 ( .A1(n4422), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n5712) );
  OAI21_X1 U5185 ( .B1(n7740), .B2(SI_29_), .A(n7743), .ZN(n7808) );
  XNOR2_X1 U5186 ( .A(n7742), .B(n7741), .ZN(n7740) );
  AOI21_X1 U5187 ( .B1(n4863), .B2(n4865), .A(n4860), .ZN(n4859) );
  INV_X1 U5188 ( .A(n5563), .ZN(n4860) );
  AND2_X1 U5189 ( .A1(n5171), .A2(n5170), .ZN(n5543) );
  AND2_X1 U5190 ( .A1(n5167), .A2(n5166), .ZN(n5531) );
  INV_X1 U5191 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5705) );
  INV_X1 U5192 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5704) );
  AOI21_X1 U5193 ( .B1(n4672), .B2(n4670), .A(n4669), .ZN(n4668) );
  INV_X1 U5194 ( .A(n5101), .ZN(n4669) );
  NOR2_X1 U5195 ( .A1(n5337), .A2(n4671), .ZN(n4670) );
  INV_X1 U5196 ( .A(n5096), .ZN(n4671) );
  INV_X1 U5197 ( .A(n5322), .ZN(n4672) );
  AND2_X1 U5198 ( .A1(n5903), .A2(n9750), .ZN(n5912) );
  NAND2_X1 U5199 ( .A1(n9971), .A2(n9795), .ZN(n5053) );
  INV_X1 U5200 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5052) );
  AOI21_X1 U5201 ( .B1(n4784), .B2(n4783), .A(n4782), .ZN(n4781) );
  INV_X1 U5202 ( .A(n4421), .ZN(n4783) );
  NOR2_X1 U5203 ( .A1(n8326), .A2(n4759), .ZN(n4758) );
  INV_X1 U5204 ( .A(n6243), .ZN(n4759) );
  OR2_X1 U5205 ( .A1(n8268), .A2(n8357), .ZN(n4789) );
  NAND2_X1 U5206 ( .A1(n6193), .A2(n6729), .ZN(n6730) );
  NAND2_X1 U5207 ( .A1(n6210), .A2(n6209), .ZN(n7140) );
  OR4_X1 U5208 ( .A1(n8239), .A2(n8238), .A3(n8237), .A4(n8236), .ZN(n8247) );
  OAI21_X1 U5209 ( .B1(n8202), .B2(n8201), .A(n8200), .ZN(n8250) );
  NAND2_X1 U5210 ( .A1(n8199), .A2(n8831), .ZN(n8200) );
  NAND2_X1 U5211 ( .A1(n8197), .A2(n8196), .ZN(n8201) );
  NOR2_X1 U5212 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n4989) );
  NAND2_X1 U5213 ( .A1(n5189), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n4576) );
  NOR2_X1 U5214 ( .A1(n5234), .A2(n9705), .ZN(n4970) );
  NAND2_X1 U5215 ( .A1(n6541), .A2(n6542), .ZN(n6540) );
  NAND2_X1 U5216 ( .A1(n4824), .A2(n4823), .ZN(n6542) );
  NAND2_X1 U5217 ( .A1(n6519), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4823) );
  OR2_X1 U5218 ( .A1(n6519), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4824) );
  NAND2_X1 U5219 ( .A1(n4634), .A2(n6508), .ZN(n6558) );
  AND2_X1 U5220 ( .A1(n6510), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4634) );
  NAND2_X1 U5221 ( .A1(n4852), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6757) );
  OR2_X1 U5222 ( .A1(n4431), .A2(n6915), .ZN(n4845) );
  NAND2_X1 U5223 ( .A1(n4850), .A2(n4409), .ZN(n4846) );
  NAND2_X1 U5224 ( .A1(n4401), .A2(n4853), .ZN(n4847) );
  NAND2_X1 U5225 ( .A1(n4850), .A2(n4854), .ZN(n4849) );
  NAND2_X1 U5226 ( .A1(n4852), .A2(n4401), .ZN(n4851) );
  NAND2_X1 U5227 ( .A1(n4643), .A2(n6915), .ZN(n4642) );
  INV_X1 U5228 ( .A(n6920), .ZN(n4643) );
  NAND2_X1 U5229 ( .A1(n6920), .A2(n4853), .ZN(n7053) );
  NAND2_X1 U5230 ( .A1(n4640), .A2(n7053), .ZN(n7055) );
  INV_X1 U5231 ( .A(n4641), .ZN(n4640) );
  OR2_X1 U5232 ( .A1(n7430), .A2(n7429), .ZN(n8417) );
  NAND2_X1 U5233 ( .A1(n8430), .A2(n4466), .ZN(n4825) );
  NAND2_X1 U5234 ( .A1(n5614), .A2(n5613), .ZN(n6501) );
  NOR2_X1 U5235 ( .A1(n8535), .A2(n10215), .ZN(n8538) );
  INV_X1 U5236 ( .A(n4820), .ZN(n8534) );
  INV_X1 U5237 ( .A(n5573), .ZN(n8571) );
  OR2_X1 U5238 ( .A1(n5547), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5549) );
  NAND2_X1 U5239 ( .A1(n5025), .A2(n5024), .ZN(n5535) );
  INV_X1 U5240 ( .A(n5522), .ZN(n5025) );
  NAND2_X1 U5241 ( .A1(n5023), .A2(n5022), .ZN(n5501) );
  INV_X1 U5242 ( .A(n5492), .ZN(n5023) );
  NOR2_X1 U5243 ( .A1(n8087), .A2(n4621), .ZN(n4620) );
  INV_X1 U5244 ( .A(n8032), .ZN(n4621) );
  AND4_X1 U5245 ( .A1(n5383), .A2(n5382), .A3(n5381), .A4(n5380), .ZN(n8308)
         );
  NOR2_X1 U5246 ( .A1(n4423), .A2(n4888), .ZN(n4887) );
  INV_X1 U5247 ( .A(n8086), .ZN(n7394) );
  OR2_X1 U5248 ( .A1(n5329), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5346) );
  NOR2_X1 U5249 ( .A1(n5629), .A2(n4612), .ZN(n4611) );
  INV_X1 U5250 ( .A(n8060), .ZN(n4612) );
  OR2_X1 U5251 ( .A1(n5291), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5305) );
  OR2_X1 U5252 ( .A1(n5263), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5277) );
  AND4_X1 U5253 ( .A1(n5195), .A2(n5194), .A3(n5193), .A4(n5192), .ZN(n6844)
         );
  INV_X1 U5254 ( .A(n8279), .ZN(n5673) );
  NAND2_X1 U5255 ( .A1(n5644), .A2(n8208), .ZN(n8617) );
  NAND2_X1 U5256 ( .A1(n4596), .A2(n4597), .ZN(n8637) );
  INV_X1 U5257 ( .A(n4598), .ZN(n4597) );
  OAI21_X1 U5258 ( .B1(n8120), .B2(n4599), .A(n8129), .ZN(n4598) );
  INV_X1 U5259 ( .A(n8118), .ZN(n4601) );
  OR2_X1 U5260 ( .A1(n8877), .A2(n6257), .ZN(n8120) );
  AND2_X1 U5261 ( .A1(n5485), .A2(n4904), .ZN(n4903) );
  INV_X1 U5262 ( .A(n8555), .ZN(n5618) );
  AND3_X1 U5263 ( .A1(n5484), .A2(n5483), .A3(n5482), .ZN(n8693) );
  NAND2_X1 U5264 ( .A1(n6287), .A2(n8171), .ZN(n8761) );
  OAI21_X1 U5265 ( .B1(n8720), .B2(n5637), .A(n5640), .ZN(n8685) );
  AOI21_X1 U5266 ( .B1(n4895), .B2(n4894), .A(n4444), .ZN(n4893) );
  INV_X1 U5267 ( .A(n4901), .ZN(n4894) );
  NAND2_X1 U5268 ( .A1(n4897), .A2(n4898), .ZN(n7722) );
  NAND2_X1 U5269 ( .A1(n7513), .A2(n4901), .ZN(n4897) );
  OAI21_X1 U5270 ( .B1(n7665), .B2(n8092), .A(n8090), .ZN(n7721) );
  INV_X1 U5271 ( .A(n8761), .ZN(n8741) );
  NAND2_X1 U5272 ( .A1(n5214), .A2(n5213), .ZN(n10240) );
  AND2_X1 U5273 ( .A1(n5212), .A2(n5211), .ZN(n5213) );
  INV_X1 U5274 ( .A(n8629), .ZN(n8765) );
  INV_X1 U5275 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5585) );
  AND2_X1 U5276 ( .A1(n4989), .A2(n4990), .ZN(n4884) );
  INV_X1 U5277 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4990) );
  AND2_X1 U5278 ( .A1(n5400), .A2(n5390), .ZN(n8455) );
  OR2_X1 U5279 ( .A1(n5297), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5341) );
  INV_X1 U5280 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n9815) );
  INV_X1 U5281 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4648) );
  INV_X1 U5282 ( .A(n7439), .ZN(n4740) );
  INV_X1 U5283 ( .A(n7550), .ZN(n4737) );
  INV_X1 U5284 ( .A(n4722), .ZN(n4721) );
  NAND2_X1 U5285 ( .A1(n6802), .A2(n4724), .ZN(n6946) );
  INV_X1 U5286 ( .A(n6002), .ZN(n6000) );
  OR2_X1 U5287 ( .A1(n5893), .A2(n5892), .ZN(n5918) );
  AND2_X1 U5288 ( .A1(n8949), .A2(n8951), .ZN(n4743) );
  INV_X1 U5289 ( .A(n6802), .ZN(n4709) );
  INV_X1 U5290 ( .A(n4717), .ZN(n4711) );
  NAND2_X1 U5291 ( .A1(n4449), .A2(n4712), .ZN(n7174) );
  NAND2_X1 U5292 ( .A1(n4707), .A2(n6802), .ZN(n4712) );
  OR2_X1 U5293 ( .A1(n4719), .A2(n4717), .ZN(n4707) );
  NAND2_X1 U5294 ( .A1(n9107), .A2(n8994), .ZN(n4747) );
  NOR2_X1 U5295 ( .A1(n6619), .A2(n6618), .ZN(n6622) );
  INV_X1 U5296 ( .A(n9342), .ZN(n8005) );
  AND2_X1 U5297 ( .A1(n6090), .A2(n6089), .ZN(n9187) );
  AND2_X1 U5298 ( .A1(n6062), .A2(n6061), .ZN(n9186) );
  AND4_X1 U5299 ( .A1(n6007), .A2(n6006), .A3(n6005), .A4(n6004), .ZN(n9060)
         );
  AND4_X1 U5300 ( .A1(n5751), .A2(n5750), .A3(n5749), .A4(n5748), .ZN(n9175)
         );
  AND4_X1 U5301 ( .A1(n5945), .A2(n5944), .A3(n5943), .A4(n5942), .ZN(n7594)
         );
  AND4_X1 U5302 ( .A1(n5874), .A2(n5873), .A3(n5872), .A4(n5871), .ZN(n7441)
         );
  AND4_X1 U5303 ( .A1(n5861), .A2(n5860), .A3(n5859), .A4(n5858), .ZN(n7177)
         );
  AND4_X1 U5304 ( .A1(n5804), .A2(n5803), .A3(n5802), .A4(n5801), .ZN(n6781)
         );
  XNOR2_X1 U5305 ( .A(n6381), .B(n4689), .ZN(n9233) );
  INV_X1 U5306 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n4689) );
  NOR2_X1 U5307 ( .A1(n6400), .A2(n4685), .ZN(n10047) );
  NOR2_X1 U5308 ( .A1(n6399), .A2(n7024), .ZN(n4685) );
  NOR2_X1 U5309 ( .A1(n10047), .A2(n10046), .ZN(n10045) );
  NOR2_X1 U5310 ( .A1(n9581), .A2(n9377), .ZN(n9376) );
  OR2_X1 U5311 ( .A1(n9395), .A2(n4522), .ZN(n4521) );
  NAND2_X1 U5312 ( .A1(n4523), .A2(n9370), .ZN(n4522) );
  NAND2_X1 U5313 ( .A1(n4517), .A2(n10072), .ZN(n4516) );
  OAI21_X1 U5314 ( .B1(n4523), .B2(n9371), .A(n4518), .ZN(n4517) );
  OR2_X1 U5315 ( .A1(n6107), .A2(n9071), .ZN(n9377) );
  NAND2_X1 U5316 ( .A1(n9438), .A2(n6128), .ZN(n9420) );
  AOI21_X1 U5317 ( .B1(n9479), .B2(n4506), .A(n4504), .ZN(n4503) );
  NAND2_X1 U5318 ( .A1(n4505), .A2(n9459), .ZN(n4504) );
  NAND2_X1 U5319 ( .A1(n4506), .A2(n4508), .ZN(n4505) );
  OR2_X1 U5320 ( .A1(n9451), .A2(n6126), .ZN(n9452) );
  OR2_X1 U5321 ( .A1(n6012), .A2(n9101), .ZN(n6025) );
  AND2_X1 U5322 ( .A1(n7922), .A2(n7910), .ZN(n9469) );
  NAND2_X1 U5323 ( .A1(n6020), .A2(n6019), .ZN(n9468) );
  NAND2_X1 U5324 ( .A1(n9497), .A2(n4816), .ZN(n9479) );
  NOR2_X1 U5325 ( .A1(n4817), .A2(n9483), .ZN(n4816) );
  NAND2_X1 U5326 ( .A1(n6125), .A2(n4818), .ZN(n9497) );
  NOR2_X1 U5327 ( .A1(n7906), .A2(n7905), .ZN(n4818) );
  NAND2_X1 U5328 ( .A1(n9516), .A2(n4931), .ZN(n4930) );
  INV_X1 U5329 ( .A(n5996), .ZN(n4931) );
  OR2_X1 U5330 ( .A1(n5758), .A2(n9763), .ZN(n6002) );
  INV_X1 U5331 ( .A(n4501), .ZN(n4500) );
  OAI21_X1 U5332 ( .B1(n4502), .B2(n7898), .A(n7916), .ZN(n4501) );
  OR2_X1 U5333 ( .A1(n7693), .A2(n9126), .ZN(n4978) );
  NAND2_X1 U5334 ( .A1(n4947), .A2(n4399), .ZN(n4946) );
  INV_X1 U5335 ( .A(n4949), .ZN(n4947) );
  NOR2_X1 U5336 ( .A1(n9202), .A2(n4655), .ZN(n4950) );
  AND2_X1 U5337 ( .A1(n7897), .A2(n9547), .ZN(n7974) );
  NOR2_X1 U5338 ( .A1(n7974), .A2(n4950), .ZN(n4949) );
  NAND2_X1 U5339 ( .A1(n4952), .A2(n7879), .ZN(n4951) );
  OR2_X1 U5340 ( .A1(n10164), .A2(n7626), .ZN(n7774) );
  NAND2_X1 U5341 ( .A1(n5741), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5966) );
  INV_X1 U5342 ( .A(n5955), .ZN(n5741) );
  NAND2_X1 U5343 ( .A1(n7487), .A2(n4814), .ZN(n7621) );
  NOR2_X1 U5344 ( .A1(n7597), .A2(n10164), .ZN(n7630) );
  NAND2_X1 U5345 ( .A1(n7485), .A2(n6122), .ZN(n7487) );
  NAND2_X1 U5346 ( .A1(n4455), .A2(n4963), .ZN(n4956) );
  NAND2_X1 U5347 ( .A1(n4960), .A2(n4961), .ZN(n4959) );
  INV_X1 U5348 ( .A(n4962), .ZN(n4960) );
  NAND2_X1 U5349 ( .A1(n4963), .A2(n4961), .ZN(n4957) );
  NAND2_X1 U5350 ( .A1(n7343), .A2(n9221), .ZN(n4962) );
  NAND2_X1 U5351 ( .A1(n7277), .A2(n5908), .ZN(n7329) );
  NAND2_X1 U5352 ( .A1(n7962), .A2(n7032), .ZN(n6116) );
  OR2_X1 U5353 ( .A1(n5868), .A2(n5867), .ZN(n5877) );
  OR2_X1 U5354 ( .A1(n7111), .A2(n9564), .ZN(n7255) );
  NAND2_X1 U5355 ( .A1(n7031), .A2(n7840), .ZN(n7030) );
  NAND2_X1 U5356 ( .A1(n7020), .A2(n7021), .ZN(n4912) );
  NOR2_X1 U5357 ( .A1(n6109), .A2(n10095), .ZN(n10086) );
  NAND2_X2 U5358 ( .A1(n7304), .A2(n7952), .ZN(n7009) );
  AND2_X1 U5359 ( .A1(n6484), .A2(n6170), .ZN(n10165) );
  AND2_X1 U5360 ( .A1(n7950), .A2(n7108), .ZN(n10148) );
  NAND2_X1 U5361 ( .A1(n6166), .A2(n6603), .ZN(n6994) );
  INV_X1 U5362 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5728) );
  XNOR2_X1 U5363 ( .A(n7808), .B(n7807), .ZN(n8161) );
  XNOR2_X1 U5364 ( .A(n7740), .B(SI_29_), .ZN(n7747) );
  XNOR2_X1 U5365 ( .A(n5724), .B(n5728), .ZN(n6130) );
  NAND2_X1 U5366 ( .A1(n5727), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5724) );
  XNOR2_X1 U5367 ( .A(n5676), .B(n5675), .ZN(n7603) );
  XNOR2_X1 U5368 ( .A(n5544), .B(n5543), .ZN(n7500) );
  NAND2_X1 U5369 ( .A1(n4538), .A2(n4536), .ZN(n5508) );
  AOI21_X1 U5370 ( .B1(n4539), .B2(n4543), .A(n4537), .ZN(n4536) );
  INV_X1 U5371 ( .A(n5151), .ZN(n4537) );
  AND2_X1 U5372 ( .A1(n5156), .A2(n5155), .ZN(n5507) );
  XNOR2_X1 U5373 ( .A(n6151), .B(n6150), .ZN(n7311) );
  NAND2_X1 U5374 ( .A1(n4541), .A2(n4542), .ZN(n5498) );
  XNOR2_X1 U5375 ( .A(n5489), .B(n5488), .ZN(n7189) );
  NAND2_X1 U5376 ( .A1(n5472), .A2(n5139), .ZN(n5487) );
  XNOR2_X1 U5377 ( .A(n5475), .B(n5474), .ZN(n7107) );
  INV_X1 U5378 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9809) );
  INV_X1 U5379 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5718) );
  NAND2_X1 U5380 ( .A1(n4869), .A2(n5116), .ZN(n5412) );
  NAND2_X1 U5381 ( .A1(n5112), .A2(n4870), .ZN(n4869) );
  XNOR2_X1 U5382 ( .A(n4650), .B(n5399), .ZN(n6690) );
  NAND2_X1 U5383 ( .A1(n5112), .A2(n5111), .ZN(n4650) );
  AND2_X1 U5384 ( .A1(n5951), .A2(n5962), .ZN(n9261) );
  NAND2_X1 U5385 ( .A1(n5106), .A2(n5105), .ZN(n5385) );
  OAI21_X1 U5386 ( .B1(n5323), .B2(n4666), .A(n4664), .ZN(n5371) );
  NAND2_X1 U5387 ( .A1(n5218), .A2(n5068), .ZN(n4653) );
  NAND2_X1 U5388 ( .A1(n5178), .A2(n5177), .ZN(n6284) );
  NAND2_X1 U5389 ( .A1(n8346), .A2(n4763), .ZN(n4762) );
  NAND2_X1 U5390 ( .A1(n4761), .A2(n8384), .ZN(n4760) );
  AOI21_X1 U5391 ( .B1(n4419), .B2(n4397), .A(n4777), .ZN(n4776) );
  AND4_X1 U5392 ( .A1(n5352), .A2(n5351), .A3(n5350), .A4(n5349), .ZN(n8303)
         );
  NAND2_X1 U5393 ( .A1(n8346), .A2(n4770), .ZN(n4768) );
  NAND2_X1 U5394 ( .A1(n7323), .A2(n6221), .ZN(n7467) );
  AOI21_X1 U5395 ( .B1(n4586), .B2(n4585), .A(n8238), .ZN(n8191) );
  AOI21_X1 U5396 ( .B1(n4588), .B2(n4587), .A(n8188), .ZN(n4586) );
  NAND2_X1 U5397 ( .A1(n8190), .A2(n8189), .ZN(n4585) );
  NAND2_X1 U5398 ( .A1(n5046), .A2(n5045), .ZN(n8400) );
  OAI21_X1 U5399 ( .B1(n10203), .B2(n6503), .A(n6504), .ZN(n10208) );
  NOR2_X1 U5400 ( .A1(n8484), .A2(n8485), .ZN(n8487) );
  AND2_X1 U5401 ( .A1(n8538), .A2(n8537), .ZN(n8539) );
  AND2_X1 U5402 ( .A1(n8541), .A2(n8548), .ZN(n4857) );
  XNOR2_X1 U5403 ( .A(n8193), .B(n5684), .ZN(n8576) );
  NOR2_X1 U5404 ( .A1(n5693), .A2(n5692), .ZN(n5694) );
  NOR2_X1 U5405 ( .A1(n8169), .A2(n8569), .ZN(n5692) );
  INV_X1 U5406 ( .A(n8752), .ZN(n8619) );
  NAND2_X1 U5407 ( .A1(n10303), .A2(n10281), .ZN(n8797) );
  NAND2_X1 U5408 ( .A1(n5602), .A2(n5601), .ZN(n6349) );
  AND2_X1 U5409 ( .A1(n6152), .A2(n6153), .ZN(n6146) );
  INV_X1 U5410 ( .A(n7027), .ZN(n5810) );
  NAND2_X1 U5411 ( .A1(n5988), .A2(n5987), .ZN(n9636) );
  AND2_X1 U5412 ( .A1(n6614), .A2(n6321), .ZN(n8013) );
  NAND2_X1 U5413 ( .A1(n4529), .A2(n4660), .ZN(n4659) );
  AND2_X1 U5414 ( .A1(n8004), .A2(n4661), .ZN(n4660) );
  NAND2_X1 U5415 ( .A1(n8011), .A2(n8012), .ZN(n4661) );
  OR2_X1 U5416 ( .A1(n9405), .A2(n6131), .ZN(n6078) );
  AND3_X1 U5417 ( .A1(n6040), .A2(n6039), .A3(n6038), .ZN(n9161) );
  OR2_X1 U5418 ( .A1(n5994), .A2(n5993), .ZN(n9217) );
  AND2_X1 U5419 ( .A1(n5824), .A2(n5836), .ZN(n10051) );
  NAND2_X1 U5420 ( .A1(n4804), .A2(n4802), .ZN(n9579) );
  AOI21_X1 U5421 ( .B1(n9363), .B2(n9173), .A(n4803), .ZN(n4802) );
  NAND2_X1 U5422 ( .A1(n4521), .A2(n4515), .ZN(n4804) );
  NOR2_X1 U5423 ( .A1(n9374), .A2(n9375), .ZN(n4803) );
  AND2_X1 U5424 ( .A1(n9562), .A2(n9342), .ZN(n10081) );
  AND2_X1 U5425 ( .A1(n4526), .A2(n7821), .ZN(n9649) );
  NAND2_X1 U5426 ( .A1(n8912), .A2(n7818), .ZN(n4526) );
  AND2_X1 U5427 ( .A1(n9571), .A2(n9574), .ZN(n9647) );
  NAND2_X1 U5428 ( .A1(n10174), .A2(n10165), .ZN(n9956) );
  OAI211_X1 U5429 ( .C1(n4496), .C2(n4495), .A(n7835), .B(n4493), .ZN(n7847)
         );
  NAND2_X1 U5430 ( .A1(n4494), .A2(n7950), .ZN(n4493) );
  NAND2_X1 U5431 ( .A1(n7827), .A2(n4433), .ZN(n4495) );
  OAI21_X1 U5432 ( .B1(n4440), .B2(n8210), .A(n4578), .ZN(n4577) );
  AND2_X1 U5433 ( .A1(n8225), .A2(n4579), .ZN(n4578) );
  NAND2_X1 U5434 ( .A1(n8089), .A2(n8186), .ZN(n4579) );
  INV_X1 U5435 ( .A(n8131), .ZN(n4573) );
  OR2_X1 U5436 ( .A1(n4573), .A2(n8171), .ZN(n4569) );
  OR2_X1 U5437 ( .A1(n4573), .A2(n8186), .ZN(n4572) );
  OR2_X1 U5438 ( .A1(n4573), .A2(n8648), .ZN(n4571) );
  INV_X1 U5439 ( .A(n7932), .ZN(n4673) );
  OAI211_X1 U5440 ( .C1(n4676), .C2(n7947), .A(n7933), .B(n4675), .ZN(n4674)
         );
  OR2_X1 U5441 ( .A1(n9486), .A2(n9160), .ZN(n7788) );
  INV_X1 U5442 ( .A(n4680), .ZN(n4679) );
  OAI21_X1 U5443 ( .B1(n7937), .B2(n7947), .A(n4681), .ZN(n4680) );
  NAND2_X1 U5444 ( .A1(n4682), .A2(n7947), .ZN(n4681) );
  INV_X1 U5445 ( .A(n9367), .ZN(n4682) );
  AND2_X1 U5446 ( .A1(n4565), .A2(n5312), .ZN(n4564) );
  NAND2_X1 U5447 ( .A1(n9229), .A2(n5810), .ZN(n7829) );
  AOI21_X1 U5448 ( .B1(n5163), .B2(n4549), .A(n4547), .ZN(n4546) );
  NAND2_X1 U5449 ( .A1(n4863), .A2(n4548), .ZN(n4547) );
  NAND2_X1 U5450 ( .A1(n4549), .A2(n4551), .ZN(n4548) );
  INV_X1 U5451 ( .A(n4864), .ZN(n4863) );
  OAI21_X1 U5452 ( .B1(n5543), .B2(n4865), .A(n5561), .ZN(n4864) );
  INV_X1 U5453 ( .A(n5171), .ZN(n4865) );
  INV_X1 U5454 ( .A(n5531), .ZN(n4551) );
  INV_X1 U5455 ( .A(n4550), .ZN(n4549) );
  OAI21_X1 U5456 ( .B1(n5162), .B2(n4551), .A(n5167), .ZN(n4550) );
  INV_X1 U5457 ( .A(n4870), .ZN(n4555) );
  INV_X1 U5458 ( .A(n4556), .ZN(n4554) );
  INV_X1 U5459 ( .A(n5116), .ZN(n4868) );
  INV_X1 U5460 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5703) );
  NOR2_X1 U5461 ( .A1(n5384), .A2(n4557), .ZN(n4556) );
  INV_X1 U5462 ( .A(n5105), .ZN(n4557) );
  NAND2_X1 U5463 ( .A1(n4561), .A2(n4560), .ZN(n4558) );
  NAND2_X1 U5464 ( .A1(n5098), .A2(n5097), .ZN(n5101) );
  INV_X1 U5465 ( .A(SI_9_), .ZN(n5089) );
  INV_X1 U5466 ( .A(n8345), .ZN(n4766) );
  INV_X1 U5467 ( .A(n8354), .ZN(n4788) );
  INV_X1 U5468 ( .A(n6225), .ZN(n4780) );
  CLKBUF_X1 U5469 ( .A(n5204), .Z(n6516) );
  INV_X1 U5470 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n9747) );
  INV_X1 U5471 ( .A(n4629), .ZN(n4625) );
  NOR2_X1 U5472 ( .A1(n7164), .A2(n4632), .ZN(n4628) );
  NAND2_X1 U5473 ( .A1(n4633), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4632) );
  INV_X1 U5474 ( .A(n7239), .ZN(n4633) );
  AOI21_X1 U5475 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n8475), .A(n8474), .ZN(
        n8498) );
  NAND2_X1 U5476 ( .A1(n8533), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4644) );
  NOR2_X1 U5477 ( .A1(n5346), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5345) );
  INV_X1 U5478 ( .A(n5321), .ZN(n4888) );
  AND2_X1 U5479 ( .A1(n6364), .A2(n5612), .ZN(n5653) );
  NAND2_X1 U5480 ( .A1(n5470), .A2(n8703), .ZN(n4904) );
  NOR2_X1 U5481 ( .A1(n7668), .A2(n4902), .ZN(n4901) );
  INV_X1 U5482 ( .A(n5369), .ZN(n4902) );
  OR2_X1 U5483 ( .A1(n6296), .A2(n8028), .ZN(n6285) );
  OR2_X1 U5484 ( .A1(n6309), .A2(n5653), .ZN(n6290) );
  INV_X1 U5485 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n4988) );
  AND3_X1 U5486 ( .A1(n4751), .A2(n4987), .A3(n4985), .ZN(n4883) );
  AND2_X1 U5487 ( .A1(n9367), .A2(n7934), .ZN(n7986) );
  INV_X1 U5488 ( .A(n7951), .ZN(n4652) );
  INV_X1 U5489 ( .A(n4968), .ZN(n4651) );
  NAND2_X1 U5490 ( .A1(n4535), .A2(n4534), .ZN(n4533) );
  NOR2_X1 U5491 ( .A1(n7981), .A2(n7984), .ZN(n4535) );
  NAND2_X1 U5492 ( .A1(n9653), .A2(n7947), .ZN(n4875) );
  NAND2_X1 U5493 ( .A1(n9360), .A2(n7950), .ZN(n4876) );
  NAND2_X1 U5494 ( .A1(n5709), .A2(n4967), .ZN(n4966) );
  INV_X1 U5495 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4967) );
  NOR2_X1 U5496 ( .A1(n9368), .A2(n4918), .ZN(n4525) );
  NAND2_X1 U5497 ( .A1(n4523), .A2(n4519), .ZN(n4518) );
  NAND2_X1 U5498 ( .A1(n4520), .A2(n9370), .ZN(n4519) );
  INV_X1 U5499 ( .A(n4525), .ZN(n4520) );
  INV_X1 U5500 ( .A(n4524), .ZN(n4523) );
  OAI21_X1 U5501 ( .B1(n9368), .B2(n7934), .A(n9367), .ZN(n4524) );
  OR2_X1 U5502 ( .A1(n9071), .A2(n9372), .ZN(n7937) );
  NAND2_X1 U5503 ( .A1(n9408), .A2(n4701), .ZN(n4700) );
  INV_X1 U5504 ( .A(n4702), .ZN(n4701) );
  OR2_X1 U5505 ( .A1(n9443), .A2(n9037), .ZN(n9417) );
  AND2_X1 U5506 ( .A1(n9504), .A2(n9060), .ZN(n7906) );
  AOI21_X1 U5507 ( .B1(n9548), .B2(n4500), .A(n4498), .ZN(n4497) );
  NAND2_X1 U5508 ( .A1(n9512), .A2(n4499), .ZN(n4498) );
  NAND2_X1 U5509 ( .A1(n4500), .A2(n4502), .ZN(n4499) );
  NOR2_X1 U5510 ( .A1(n9049), .A2(n7343), .ZN(n4693) );
  AND2_X1 U5511 ( .A1(n6115), .A2(n7851), .ZN(n7962) );
  NOR2_X1 U5512 ( .A1(n9452), .A2(n9443), .ZN(n9442) );
  NAND2_X1 U5513 ( .A1(n7279), .A2(n4400), .ZN(n7494) );
  AND2_X1 U5514 ( .A1(n4807), .A2(n5723), .ZN(n4806) );
  OR2_X1 U5515 ( .A1(n5713), .A2(n4808), .ZN(n4807) );
  AND2_X1 U5516 ( .A1(n5677), .A2(n5568), .ZN(n5675) );
  AND2_X1 U5517 ( .A1(n5162), .A2(n5161), .ZN(n5518) );
  NAND2_X1 U5518 ( .A1(n4544), .A2(n4413), .ZN(n4542) );
  AND2_X1 U5519 ( .A1(n5486), .A2(n5145), .ZN(n5146) );
  NAND2_X1 U5520 ( .A1(n5139), .A2(n4413), .ZN(n4543) );
  NAND2_X1 U5521 ( .A1(n5715), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5984) );
  NAND2_X1 U5522 ( .A1(n5106), .A2(n4556), .ZN(n5112) );
  INV_X1 U5523 ( .A(SI_14_), .ZN(n5107) );
  AOI21_X1 U5524 ( .B1(n4402), .B2(n4665), .A(n4451), .ZN(n4664) );
  INV_X1 U5525 ( .A(n4670), .ZN(n4665) );
  INV_X1 U5526 ( .A(n4402), .ZN(n4666) );
  NAND2_X1 U5527 ( .A1(n4488), .A2(n4487), .ZN(n5072) );
  NAND2_X1 U5528 ( .A1(n6325), .A2(n9808), .ZN(n4487) );
  OR2_X1 U5529 ( .A1(n6325), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n4488) );
  OAI21_X1 U5530 ( .B1(n5779), .B2(P1_DATAO_REG_3__SCAN_IN), .A(n5063), .ZN(
        n5066) );
  NAND2_X1 U5531 ( .A1(n5779), .A2(n6342), .ZN(n5063) );
  INV_X1 U5532 ( .A(n4769), .ZN(n4761) );
  NOR2_X1 U5533 ( .A1(n4771), .A2(n4767), .ZN(n4763) );
  NAND2_X1 U5534 ( .A1(n8384), .A2(n8385), .ZN(n4773) );
  NAND2_X1 U5535 ( .A1(n6272), .A2(n6273), .ZN(n6274) );
  INV_X1 U5536 ( .A(n7503), .ZN(n4777) );
  INV_X1 U5537 ( .A(n6264), .ZN(n4753) );
  INV_X1 U5538 ( .A(n8406), .ZN(n7314) );
  NAND2_X1 U5539 ( .A1(n6251), .A2(n4421), .ZN(n4786) );
  NAND2_X1 U5540 ( .A1(n6223), .A2(n6222), .ZN(n7465) );
  NAND2_X1 U5541 ( .A1(n7465), .A2(n6225), .ZN(n7699) );
  XNOR2_X1 U5542 ( .A(n6197), .B(n10240), .ZN(n6195) );
  NOR3_X1 U5543 ( .A1(n8187), .A2(n8186), .A3(n8237), .ZN(n4587) );
  INV_X1 U5544 ( .A(n4592), .ZN(n4591) );
  AND2_X1 U5545 ( .A1(n8182), .A2(n8181), .ZN(n8570) );
  OR2_X1 U5546 ( .A1(n6522), .A2(n6521), .ZN(n6523) );
  NAND2_X1 U5547 ( .A1(n4834), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6562) );
  INV_X1 U5548 ( .A(n6560), .ZN(n4834) );
  NAND2_X1 U5549 ( .A1(n4635), .A2(n6509), .ZN(n6653) );
  NAND2_X1 U5550 ( .A1(n4642), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4641) );
  OR2_X1 U5551 ( .A1(n5341), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5314) );
  INV_X1 U5552 ( .A(n4628), .ZN(n4627) );
  NAND2_X1 U5553 ( .A1(n4630), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7240) );
  INV_X1 U5554 ( .A(n7164), .ZN(n4630) );
  AND2_X1 U5555 ( .A1(n4840), .A2(n7229), .ZN(n4844) );
  OAI211_X1 U5556 ( .C1(n4626), .C2(n4628), .A(n4624), .B(n4623), .ZN(n7367)
         );
  NAND2_X1 U5557 ( .A1(n4625), .A2(n7418), .ZN(n4624) );
  NAND2_X1 U5558 ( .A1(n4629), .A2(n7424), .ZN(n4626) );
  NAND2_X1 U5559 ( .A1(n4628), .A2(n7418), .ZN(n4623) );
  NOR2_X1 U5560 ( .A1(n7357), .A2(n4485), .ZN(n7409) );
  NOR2_X1 U5561 ( .A1(n7244), .A2(n5328), .ZN(n4485) );
  AND2_X1 U5562 ( .A1(n4828), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4826) );
  NOR2_X1 U5563 ( .A1(n8453), .A2(n8454), .ZN(n8457) );
  OR2_X1 U5564 ( .A1(n8570), .A2(n8569), .ZN(n8776) );
  OAI21_X1 U5565 ( .B1(n8600), .B2(n4614), .A(n4613), .ZN(n8193) );
  AOI21_X1 U5566 ( .B1(n4615), .B2(n8148), .A(n4616), .ZN(n4613) );
  INV_X1 U5567 ( .A(n4615), .ZN(n4614) );
  NOR2_X1 U5568 ( .A1(n8156), .A2(n8761), .ZN(n5693) );
  INV_X1 U5569 ( .A(n4909), .ZN(n8585) );
  INV_X1 U5570 ( .A(n5535), .ZN(n5027) );
  OR2_X1 U5571 ( .A1(n5511), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5522) );
  NAND2_X1 U5572 ( .A1(n5021), .A2(n5020), .ZN(n5492) );
  NAND2_X1 U5573 ( .A1(n5019), .A2(n5018), .ZN(n5464) );
  NAND2_X1 U5574 ( .A1(n5017), .A2(n5016), .ZN(n5419) );
  INV_X1 U5575 ( .A(n5404), .ZN(n5017) );
  OR2_X1 U5576 ( .A1(n5419), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5447) );
  OR2_X1 U5577 ( .A1(n5393), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5404) );
  NAND2_X1 U5578 ( .A1(n5015), .A2(n9783), .ZN(n5393) );
  INV_X1 U5579 ( .A(n5378), .ZN(n5015) );
  NAND2_X1 U5580 ( .A1(n5631), .A2(n5630), .ZN(n7472) );
  NAND2_X1 U5581 ( .A1(n7347), .A2(n5321), .ZN(n7475) );
  NAND2_X1 U5582 ( .A1(n5013), .A2(n5012), .ZN(n5329) );
  INV_X1 U5583 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5012) );
  INV_X1 U5584 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5010) );
  INV_X1 U5585 ( .A(n5277), .ZN(n5011) );
  NAND2_X1 U5586 ( .A1(n4886), .A2(n5276), .ZN(n7193) );
  INV_X1 U5587 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5008) );
  AND4_X1 U5588 ( .A1(n5269), .A2(n5268), .A3(n5267), .A4(n5266), .ZN(n7207)
         );
  AND2_X1 U5589 ( .A1(n8071), .A2(n8068), .ZN(n8214) );
  NAND2_X1 U5590 ( .A1(n8212), .A2(n5624), .ZN(n6840) );
  AND2_X1 U5591 ( .A1(n8141), .A2(n8147), .ZN(n8604) );
  INV_X1 U5592 ( .A(n8604), .ZN(n8599) );
  OR2_X1 U5593 ( .A1(n8142), .A2(n8140), .ZN(n8618) );
  OR2_X1 U5594 ( .A1(n8135), .A2(n8130), .ZN(n8638) );
  NAND2_X1 U5595 ( .A1(n8704), .A2(n5470), .ZN(n8690) );
  NAND2_X1 U5596 ( .A1(n7302), .A2(n5647), .ZN(n10268) );
  AND2_X1 U5597 ( .A1(n6318), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6708) );
  NOR2_X1 U5598 ( .A1(n4441), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n4892) );
  AND2_X1 U5599 ( .A1(n5591), .A2(n5595), .ZN(n5597) );
  INV_X1 U5600 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n9797) );
  CLKBUF_X1 U5601 ( .A(n5430), .Z(n5431) );
  NAND2_X1 U5602 ( .A1(n8913), .A2(n4984), .ZN(n4837) );
  NAND3_X1 U5603 ( .A1(n4839), .A2(P2_IR_REG_2__SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n4838) );
  INV_X1 U5604 ( .A(n4739), .ZN(n4736) );
  NAND2_X1 U5605 ( .A1(n4741), .A2(n7439), .ZN(n7526) );
  NAND2_X1 U5606 ( .A1(n4742), .A2(n4478), .ZN(n4741) );
  AOI21_X1 U5607 ( .B1(n4728), .B2(n4730), .A(n4450), .ZN(n4726) );
  NAND2_X1 U5608 ( .A1(n4733), .A2(n4738), .ZN(n7651) );
  NAND2_X1 U5609 ( .A1(n4742), .A2(n4739), .ZN(n4733) );
  XNOR2_X1 U5610 ( .A(n4731), .B(n8997), .ZN(n6634) );
  OAI21_X1 U5611 ( .B1(n8996), .B2(n6106), .A(n6630), .ZN(n4731) );
  OAI21_X1 U5612 ( .B1(n6699), .B2(n6698), .A(n6697), .ZN(n6769) );
  INV_X1 U5613 ( .A(n9350), .ZN(n9150) );
  NOR2_X1 U5614 ( .A1(n9649), .A2(n9353), .ZN(n8006) );
  OAI21_X1 U5615 ( .B1(n6102), .B2(n4966), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6148) );
  AND4_X1 U5616 ( .A1(n5934), .A2(n5933), .A3(n5932), .A4(n5931), .ZN(n7552)
         );
  AND4_X1 U5617 ( .A1(n5883), .A2(n5882), .A3(n5881), .A4(n5880), .ZN(n7445)
         );
  AND4_X1 U5618 ( .A1(n5847), .A2(n5846), .A3(n5845), .A4(n5844), .ZN(n7092)
         );
  AND4_X1 U5619 ( .A1(n5835), .A2(n5834), .A3(n5833), .A4(n5832), .ZN(n6947)
         );
  AND4_X1 U5620 ( .A1(n4426), .A2(n5794), .A3(n5793), .A4(n5792), .ZN(n6693)
         );
  OR2_X1 U5621 ( .A1(n4979), .A2(n5789), .ZN(n5794) );
  NOR2_X1 U5622 ( .A1(n9233), .A2(n9243), .ZN(n9232) );
  NOR2_X1 U5623 ( .A1(n6471), .A2(n4686), .ZN(n6474) );
  AND2_X1 U5624 ( .A1(n6472), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4686) );
  NAND2_X1 U5625 ( .A1(n6474), .A2(n6473), .ZN(n6670) );
  NOR2_X1 U5626 ( .A1(n6871), .A2(n4687), .ZN(n6873) );
  AND2_X1 U5627 ( .A1(n6872), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4687) );
  NAND2_X1 U5628 ( .A1(n6873), .A2(n6874), .ZN(n7076) );
  NOR2_X1 U5629 ( .A1(n9260), .A2(n4483), .ZN(n9279) );
  AND3_X1 U5630 ( .A1(n7804), .A2(n7803), .A3(n7802), .ZN(n9374) );
  AOI21_X1 U5631 ( .B1(n4915), .B2(n4396), .A(n4410), .ZN(n6099) );
  AOI21_X1 U5632 ( .B1(n9438), .B2(n4799), .A(n4797), .ZN(n4796) );
  NAND2_X1 U5633 ( .A1(n4798), .A2(n7795), .ZN(n4797) );
  NAND2_X1 U5634 ( .A1(n4799), .A2(n4801), .ZN(n4798) );
  NOR2_X1 U5635 ( .A1(n9452), .A2(n4702), .ZN(n9425) );
  NAND2_X1 U5636 ( .A1(n6023), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6035) );
  NAND2_X1 U5637 ( .A1(n9497), .A2(n9494), .ZN(n9477) );
  AND2_X1 U5638 ( .A1(n4927), .A2(n4926), .ZN(n9484) );
  AOI21_X1 U5639 ( .B1(n6009), .B2(n4933), .A(n6008), .ZN(n4926) );
  AND2_X1 U5640 ( .A1(n9539), .A2(n4696), .ZN(n9485) );
  AND2_X1 U5641 ( .A1(n9942), .A2(n4407), .ZN(n4696) );
  NAND2_X1 U5642 ( .A1(n6125), .A2(n7917), .ZN(n9495) );
  NAND2_X1 U5643 ( .A1(n9539), .A2(n9951), .ZN(n9528) );
  NAND2_X1 U5644 ( .A1(n9539), .A2(n4697), .ZN(n4975) );
  NAND2_X1 U5645 ( .A1(n4940), .A2(n4942), .ZN(n9525) );
  AOI21_X1 U5646 ( .B1(n4946), .B2(n4944), .A(n4943), .ZN(n4942) );
  NOR2_X1 U5647 ( .A1(n9544), .A2(n8941), .ZN(n4943) );
  NAND2_X1 U5648 ( .A1(n5744), .A2(n5743), .ZN(n5758) );
  OR2_X1 U5649 ( .A1(n5978), .A2(n9286), .ZN(n5991) );
  NAND2_X1 U5650 ( .A1(n5742), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5978) );
  INV_X1 U5651 ( .A(n5966), .ZN(n5742) );
  INV_X1 U5652 ( .A(n4814), .ZN(n4813) );
  NAND2_X1 U5653 ( .A1(n4812), .A2(n4814), .ZN(n4811) );
  OR2_X1 U5654 ( .A1(n5939), .A2(n7085), .ZN(n5955) );
  NAND2_X1 U5655 ( .A1(n5740), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5927) );
  INV_X1 U5656 ( .A(n5918), .ZN(n5740) );
  OR2_X1 U5657 ( .A1(n5927), .A2(n6876), .ZN(n5939) );
  OR2_X1 U5658 ( .A1(n7343), .A2(n7537), .ZN(n7866) );
  NAND2_X1 U5659 ( .A1(n7279), .A2(n4693), .ZN(n7388) );
  AND2_X1 U5660 ( .A1(n7279), .A2(n7296), .ZN(n7328) );
  NAND2_X1 U5661 ( .A1(n4510), .A2(n4509), .ZN(n7384) );
  NOR2_X1 U5662 ( .A1(n7867), .A2(n7769), .ZN(n4509) );
  NAND2_X1 U5663 ( .A1(n4510), .A2(n7863), .ZN(n7331) );
  NAND2_X1 U5664 ( .A1(n5739), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5893) );
  NAND2_X1 U5665 ( .A1(n4934), .A2(n4937), .ZN(n7253) );
  AOI21_X1 U5666 ( .B1(n7115), .B2(n4938), .A(n4446), .ZN(n4937) );
  OAI21_X1 U5667 ( .B1(n6979), .B2(n7956), .A(n4911), .ZN(n6962) );
  NAND2_X1 U5668 ( .A1(n6947), .A2(n10065), .ZN(n4911) );
  AND2_X1 U5669 ( .A1(n6980), .A2(n7102), .ZN(n7039) );
  NAND2_X1 U5670 ( .A1(n7126), .A2(n7836), .ZN(n6981) );
  AND2_X1 U5671 ( .A1(n7760), .A2(n7838), .ZN(n7956) );
  OAI21_X1 U5672 ( .B1(n7834), .B2(n7021), .A(n7830), .ZN(n7126) );
  OR2_X1 U5673 ( .A1(n5773), .A2(n6626), .ZN(n10093) );
  NOR2_X2 U5674 ( .A1(n10093), .A2(n5795), .ZN(n10077) );
  NAND2_X1 U5675 ( .A1(n6112), .A2(n6111), .ZN(n10076) );
  OR2_X1 U5676 ( .A1(n7009), .A2(n8002), .ZN(n9540) );
  INV_X1 U5677 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5725) );
  INV_X1 U5678 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4695) );
  XNOR2_X1 U5679 ( .A(n6141), .B(P1_IR_REG_25__SCAN_IN), .ZN(n6152) );
  NAND2_X1 U5680 ( .A1(n4418), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6141) );
  CLKBUF_X1 U5681 ( .A(n6142), .Z(n6143) );
  NAND2_X1 U5682 ( .A1(n4667), .A2(n4668), .ZN(n5357) );
  NAND2_X1 U5683 ( .A1(n5323), .A2(n4670), .ZN(n4667) );
  AND2_X1 U5684 ( .A1(n5905), .A2(n5904), .ZN(n6788) );
  NAND2_X1 U5685 ( .A1(n4654), .A2(n5071), .ZN(n5254) );
  NAND2_X1 U5686 ( .A1(n5182), .A2(n5183), .ZN(n4527) );
  XNOR2_X1 U5687 ( .A(n5057), .B(SI_1_), .ZN(n5183) );
  AND2_X1 U5688 ( .A1(n7140), .A2(n6213), .ZN(n7204) );
  OAI211_X1 U5689 ( .C1(n6261), .C2(n4757), .A(n4754), .B(n4752), .ZN(n8261)
         );
  AOI21_X1 U5690 ( .B1(n8361), .B2(n4756), .A(n4755), .ZN(n4754) );
  NAND2_X1 U5691 ( .A1(n6261), .A2(n4469), .ZN(n4752) );
  NOR2_X1 U5692 ( .A1(n6264), .A2(n6263), .ZN(n4755) );
  AND4_X1 U5693 ( .A1(n5238), .A2(n5237), .A3(n5236), .A4(n5235), .ZN(n6901)
         );
  NAND2_X1 U5694 ( .A1(n6251), .A2(n6250), .ZN(n8270) );
  AOI21_X1 U5695 ( .B1(n8278), .B2(n8400), .A(n8277), .ZN(n8282) );
  NAND2_X1 U5696 ( .A1(n8035), .A2(n6192), .ZN(n6729) );
  AND2_X1 U5697 ( .A1(n5528), .A2(n5527), .ZN(n8614) );
  NAND2_X1 U5698 ( .A1(n7639), .A2(n6243), .ZN(n8325) );
  AND4_X1 U5699 ( .A1(n5334), .A2(n5333), .A3(n5332), .A4(n5331), .ZN(n7701)
         );
  AND4_X1 U5700 ( .A1(n5469), .A2(n5468), .A3(n5467), .A4(n5466), .ZN(n8357)
         );
  NAND2_X1 U5701 ( .A1(n4786), .A2(n4789), .ZN(n8353) );
  OAI21_X1 U5702 ( .B1(n7465), .B2(n4397), .A(n4419), .ZN(n7505) );
  NAND2_X1 U5703 ( .A1(n6261), .A2(n6260), .ZN(n8363) );
  INV_X1 U5704 ( .A(n8731), .ZN(n8377) );
  OAI21_X1 U5705 ( .B1(n8386), .B2(n8385), .A(n8384), .ZN(n8383) );
  AOI21_X1 U5706 ( .B1(n6240), .B2(n6239), .A(n4973), .ZN(n7641) );
  NAND2_X1 U5707 ( .A1(n7641), .A2(n7640), .ZN(n7639) );
  INV_X1 U5708 ( .A(n8381), .ZN(n8387) );
  INV_X1 U5709 ( .A(n8250), .ZN(n8205) );
  XNOR2_X1 U5710 ( .A(n5582), .B(P2_IR_REG_20__SCAN_IN), .ZN(n8254) );
  NAND2_X1 U5711 ( .A1(n4885), .A2(n4989), .ZN(n5581) );
  OR2_X1 U5712 ( .A1(n8186), .A2(n6182), .ZN(n8027) );
  CLKBUF_X1 U5713 ( .A(n5001), .Z(n8026) );
  XNOR2_X1 U5714 ( .A(n5004), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8029) );
  AND2_X1 U5715 ( .A1(n8182), .A2(n5690), .ZN(n8169) );
  INV_X1 U5716 ( .A(n8631), .ZN(n8401) );
  INV_X1 U5717 ( .A(n8614), .ZN(n8640) );
  OAI211_X1 U5718 ( .C1(n5234), .C2(n8870), .A(n5504), .B(n5503), .ZN(n8664)
         );
  OAI211_X1 U5719 ( .C1(n5234), .C2(n8876), .A(n5495), .B(n5494), .ZN(n8676)
         );
  INV_X1 U5720 ( .A(n8357), .ZN(n8706) );
  INV_X1 U5721 ( .A(n8303), .ZN(n8404) );
  INV_X1 U5722 ( .A(n7701), .ZN(n8405) );
  AND2_X1 U5723 ( .A1(n5295), .A2(n4576), .ZN(n4575) );
  OR2_X1 U5724 ( .A1(n8179), .A2(n10289), .ZN(n5202) );
  OR2_X1 U5725 ( .A1(n6501), .A2(n6396), .ZN(n8527) );
  AND3_X1 U5726 ( .A1(n5256), .A2(n4822), .A3(n4821), .ZN(n6567) );
  NAND2_X1 U5727 ( .A1(n8913), .A2(n5222), .ZN(n4821) );
  NAND2_X1 U5728 ( .A1(n5221), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n4822) );
  NAND2_X1 U5729 ( .A1(n4851), .A2(n4849), .ZN(n6914) );
  NOR2_X1 U5730 ( .A1(n7057), .A2(n4429), .ZN(n6916) );
  AND2_X1 U5731 ( .A1(n4849), .A2(n4431), .ZN(n4848) );
  NAND2_X1 U5732 ( .A1(n4642), .A2(n7053), .ZN(n6921) );
  NOR2_X1 U5733 ( .A1(n7152), .A2(n10297), .ZN(n7226) );
  OAI21_X1 U5734 ( .B1(n7152), .B2(n4842), .A(n4841), .ZN(n7357) );
  NAND2_X1 U5735 ( .A1(n4843), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4842) );
  NAND2_X1 U5736 ( .A1(n4844), .A2(n4843), .ZN(n4841) );
  INV_X1 U5737 ( .A(n7227), .ZN(n4843) );
  XNOR2_X1 U5738 ( .A(n7409), .B(n7424), .ZN(n7358) );
  OAI211_X1 U5739 ( .C1(n8417), .C2(n8452), .A(n4636), .B(n4637), .ZN(n8418)
         );
  NAND2_X1 U5740 ( .A1(n4638), .A2(n4639), .ZN(n4637) );
  NAND2_X1 U5741 ( .A1(n8417), .A2(n4470), .ZN(n4636) );
  INV_X1 U5742 ( .A(n8416), .ZN(n4638) );
  NAND2_X1 U5743 ( .A1(n5434), .A2(n5433), .ZN(n8818) );
  OR2_X1 U5744 ( .A1(n10274), .A2(n5647), .ZN(n8632) );
  NAND2_X1 U5745 ( .A1(n7400), .A2(n8032), .ZN(n7516) );
  NAND2_X1 U5746 ( .A1(n5327), .A2(n5326), .ZN(n10272) );
  NAND2_X1 U5747 ( .A1(n4608), .A2(n4609), .ZN(n7346) );
  NAND2_X1 U5748 ( .A1(n7191), .A2(n4611), .ZN(n4608) );
  OAI21_X1 U5749 ( .B1(n7191), .B2(n8056), .A(n8060), .ZN(n7222) );
  INV_X1 U5750 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6860) );
  OR2_X1 U5751 ( .A1(n8725), .A2(n5667), .ZN(n8752) );
  INV_X1 U5752 ( .A(n8595), .ZN(n8749) );
  INV_X2 U5753 ( .A(n8725), .ZN(n8745) );
  INV_X1 U5754 ( .A(n5683), .ZN(n5681) );
  NAND2_X1 U5755 ( .A1(n8175), .A2(n8174), .ZN(n8831) );
  NAND2_X1 U5756 ( .A1(n8163), .A2(n8162), .ZN(n8835) );
  NAND2_X1 U5757 ( .A1(n5570), .A2(n5569), .ZN(n8288) );
  OR2_X1 U5758 ( .A1(n8783), .A2(n8910), .ZN(n5649) );
  INV_X1 U5759 ( .A(n6284), .ZN(n8843) );
  NAND2_X1 U5760 ( .A1(n5546), .A2(n5545), .ZN(n8846) );
  NAND2_X1 U5761 ( .A1(n5534), .A2(n5533), .ZN(n8853) );
  NAND2_X1 U5762 ( .A1(n5521), .A2(n5520), .ZN(n8859) );
  NAND2_X1 U5763 ( .A1(n5510), .A2(n5509), .ZN(n8865) );
  NAND2_X1 U5764 ( .A1(n5500), .A2(n5499), .ZN(n8871) );
  NAND2_X1 U5765 ( .A1(n4600), .A2(n8120), .ZN(n8645) );
  NAND2_X1 U5766 ( .A1(n5642), .A2(n4405), .ZN(n4600) );
  NAND2_X1 U5767 ( .A1(n5491), .A2(n5490), .ZN(n8877) );
  NAND2_X1 U5768 ( .A1(n5642), .A2(n8118), .ZN(n8658) );
  NAND2_X1 U5769 ( .A1(n5477), .A2(n5476), .ZN(n8883) );
  NAND2_X1 U5770 ( .A1(n5463), .A2(n5462), .ZN(n8889) );
  NAND2_X1 U5771 ( .A1(n5446), .A2(n5445), .ZN(n8894) );
  NAND2_X1 U5772 ( .A1(n5418), .A2(n5417), .ZN(n8901) );
  NAND2_X1 U5773 ( .A1(n5403), .A2(n5402), .ZN(n8907) );
  NAND2_X1 U5774 ( .A1(n5392), .A2(n5391), .ZN(n7736) );
  AND2_X1 U5775 ( .A1(n7725), .A2(n7724), .ZN(n7734) );
  NAND2_X1 U5776 ( .A1(n5377), .A2(n5376), .ZN(n7713) );
  OAI21_X1 U5777 ( .B1(n7513), .B2(n5370), .A(n5369), .ZN(n7669) );
  NOR2_X1 U5778 ( .A1(n5035), .A2(n5034), .ZN(n5036) );
  NOR2_X1 U5779 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n5034) );
  INV_X1 U5780 ( .A(n5597), .ZN(n7524) );
  NAND2_X1 U5781 ( .A1(n5587), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5589) );
  INV_X1 U5782 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n9756) );
  INV_X1 U5783 ( .A(n8029), .ZN(n7302) );
  INV_X1 U5784 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n9776) );
  INV_X1 U5785 ( .A(n8254), .ZN(n8203) );
  INV_X1 U5786 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n9924) );
  INV_X1 U5787 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7008) );
  INV_X1 U5788 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6930) );
  INV_X1 U5789 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6865) );
  INV_X1 U5790 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n9732) );
  INV_X1 U5791 ( .A(n8455), .ZN(n8475) );
  INV_X1 U5792 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6453) );
  INV_X1 U5793 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6395) );
  INV_X1 U5794 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6359) );
  INV_X1 U5795 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6356) );
  INV_X1 U5796 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9733) );
  XNOR2_X1 U5797 ( .A(n5298), .B(n9815), .ZN(n7160) );
  INV_X1 U5798 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6343) );
  INV_X1 U5799 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6333) );
  INV_X1 U5800 ( .A(n6743), .ZN(n6668) );
  INV_X1 U5801 ( .A(n6567), .ZN(n6521) );
  NAND2_X1 U5802 ( .A1(n4453), .A2(P2_IR_REG_1__SCAN_IN), .ZN(n4649) );
  NAND2_X1 U5803 ( .A1(n8913), .A2(n4648), .ZN(n4647) );
  NAND2_X1 U5804 ( .A1(n6081), .A2(n6080), .ZN(n9389) );
  NAND2_X1 U5805 ( .A1(n5953), .A2(n5952), .ZN(n10164) );
  NAND2_X1 U5806 ( .A1(n6032), .A2(n6031), .ZN(n6126) );
  NAND2_X1 U5807 ( .A1(n5722), .A2(n5721), .ZN(n9625) );
  AOI21_X1 U5808 ( .B1(n9137), .B2(n4415), .A(n4745), .ZN(n9075) );
  OAI21_X1 U5809 ( .B1(n4746), .B2(n9107), .A(n9023), .ZN(n4745) );
  INV_X1 U5810 ( .A(n4415), .ZN(n4746) );
  AND2_X1 U5811 ( .A1(n9016), .A2(n9015), .ZN(n9081) );
  OR4_X2 U5812 ( .A1(n9075), .A2(n9081), .A3(n9082), .A4(n9204), .ZN(n9086) );
  NAND2_X1 U5813 ( .A1(n4727), .A2(n8968), .ZN(n9097) );
  NAND2_X1 U5814 ( .A1(n9149), .A2(n9148), .ZN(n4727) );
  NAND2_X1 U5815 ( .A1(n4714), .A2(n4715), .ZN(n7095) );
  NAND2_X1 U5816 ( .A1(n6802), .A2(n4717), .ZN(n4714) );
  AND2_X1 U5817 ( .A1(n8938), .A2(n8937), .ZN(n8939) );
  AOI21_X1 U5818 ( .B1(n6605), .B2(n6604), .A(P1_U3086), .ZN(n9145) );
  AND2_X1 U5819 ( .A1(n6640), .A2(n6639), .ZN(n6699) );
  NAND2_X1 U5820 ( .A1(n4710), .A2(n4708), .ZN(n7097) );
  NAND2_X1 U5821 ( .A1(n4709), .A2(n4713), .ZN(n4708) );
  OAI21_X1 U5822 ( .B1(n9137), .B2(n4748), .A(n4415), .ZN(n9183) );
  AND2_X1 U5823 ( .A1(n6622), .A2(n6621), .ZN(n9184) );
  INV_X1 U5824 ( .A(n9143), .ZN(n9195) );
  NAND2_X1 U5825 ( .A1(n6625), .A2(n9559), .ZN(n9201) );
  INV_X1 U5826 ( .A(n8017), .ZN(n4658) );
  XNOR2_X1 U5827 ( .A(n6148), .B(P1_IR_REG_22__SCAN_IN), .ZN(n8015) );
  OR2_X1 U5828 ( .A1(n6017), .A2(n6016), .ZN(n9213) );
  AND4_X1 U5829 ( .A1(n5961), .A2(n5960), .A3(n5959), .A4(n5958), .ZN(n7626)
         );
  INV_X1 U5830 ( .A(n6947), .ZN(n9227) );
  OR2_X1 U5831 ( .A1(n5800), .A2(n5774), .ZN(n5775) );
  OR2_X1 U5832 ( .A1(n4979), .A2(n7015), .ZN(n5778) );
  OR2_X1 U5833 ( .A1(n6131), .A2(n6629), .ZN(n5777) );
  NOR2_X1 U5834 ( .A1(n10045), .A2(n4472), .ZN(n6404) );
  NOR2_X1 U5835 ( .A1(n6404), .A2(n6403), .ZN(n6418) );
  NOR2_X1 U5836 ( .A1(n6436), .A2(n4467), .ZN(n6439) );
  NOR2_X1 U5837 ( .A1(n6439), .A2(n6438), .ZN(n6471) );
  NOR2_X1 U5838 ( .A1(n6787), .A2(n4688), .ZN(n6791) );
  AND2_X1 U5839 ( .A1(n6788), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4688) );
  NOR2_X1 U5840 ( .A1(n6791), .A2(n6790), .ZN(n6871) );
  NOR2_X1 U5841 ( .A1(n7261), .A2(n4691), .ZN(n7265) );
  AND2_X1 U5842 ( .A1(n7262), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4691) );
  NOR2_X1 U5843 ( .A1(n7265), .A2(n7264), .ZN(n9260) );
  XNOR2_X1 U5844 ( .A(n9279), .B(n9278), .ZN(n9262) );
  OR2_X1 U5845 ( .A1(n10041), .A2(n6373), .ZN(n10044) );
  OR2_X1 U5846 ( .A1(n10041), .A2(n6371), .ZN(n9335) );
  INV_X1 U5847 ( .A(n9336), .ZN(n10057) );
  AOI21_X1 U5848 ( .B1(n7747), .B2(n7818), .A(n4477), .ZN(n9383) );
  NAND2_X1 U5849 ( .A1(n4916), .A2(n4417), .ZN(n9387) );
  NAND2_X1 U5850 ( .A1(n9420), .A2(n7794), .ZN(n9410) );
  NAND2_X1 U5851 ( .A1(n4923), .A2(n6063), .ZN(n9402) );
  NAND2_X1 U5852 ( .A1(n4915), .A2(n4924), .ZN(n4923) );
  OAI21_X1 U5853 ( .B1(n9479), .B2(n4508), .A(n4506), .ZN(n9458) );
  INV_X1 U5854 ( .A(n6126), .ZN(n9456) );
  NAND2_X1 U5855 ( .A1(n9479), .A2(n7909), .ZN(n9465) );
  NAND2_X1 U5856 ( .A1(n6022), .A2(n6021), .ZN(n9474) );
  NAND2_X1 U5857 ( .A1(n9622), .A2(n4932), .ZN(n9502) );
  OR2_X1 U5858 ( .A1(n5997), .A2(n4930), .ZN(n9622) );
  OAI21_X1 U5859 ( .B1(n9548), .B2(n4502), .A(n4500), .ZN(n9513) );
  NAND2_X1 U5860 ( .A1(n9548), .A2(n7898), .ZN(n9533) );
  NAND2_X1 U5861 ( .A1(n4941), .A2(n4946), .ZN(n9538) );
  NAND2_X1 U5862 ( .A1(n4952), .A2(n4395), .ZN(n4941) );
  NAND2_X1 U5863 ( .A1(n4951), .A2(n4948), .ZN(n7691) );
  INV_X1 U5864 ( .A(n4950), .ZN(n4948) );
  NAND2_X1 U5865 ( .A1(n5977), .A2(n5976), .ZN(n9126) );
  NAND2_X1 U5866 ( .A1(n7487), .A2(n7880), .ZN(n7592) );
  NAND2_X1 U5867 ( .A1(n4955), .A2(n4956), .ZN(n7492) );
  OR2_X1 U5868 ( .A1(n7329), .A2(n4957), .ZN(n4955) );
  NAND2_X1 U5869 ( .A1(n4958), .A2(n4961), .ZN(n7387) );
  NAND2_X1 U5870 ( .A1(n7329), .A2(n4962), .ZN(n4958) );
  NAND2_X1 U5871 ( .A1(n7765), .A2(n6118), .ZN(n7281) );
  NAND2_X1 U5872 ( .A1(n7110), .A2(n7115), .ZN(n7109) );
  NAND2_X1 U5873 ( .A1(n7030), .A2(n5866), .ZN(n7110) );
  NAND2_X1 U5874 ( .A1(n4912), .A2(n5811), .ZN(n7129) );
  INV_X1 U5875 ( .A(n9557), .ZN(n10082) );
  OR3_X1 U5876 ( .A1(n6994), .A2(n6993), .A3(n6992), .ZN(n6995) );
  AND2_X1 U5877 ( .A1(n8013), .A2(n6624), .ZN(n10091) );
  INV_X1 U5878 ( .A(n10091), .ZN(n9559) );
  INV_X1 U5879 ( .A(n10096), .ZN(n10074) );
  AND2_X1 U5880 ( .A1(n8018), .A2(n8020), .ZN(n6139) );
  NAND2_X1 U5881 ( .A1(n4514), .A2(n4513), .ZN(n9564) );
  AND2_X1 U5882 ( .A1(n5875), .A2(n4458), .ZN(n4513) );
  NAND2_X1 U5883 ( .A1(n6346), .A2(n7818), .ZN(n4514) );
  NOR2_X1 U5884 ( .A1(n4406), .A2(n9579), .ZN(n9582) );
  AND2_X1 U5885 ( .A1(n6054), .A2(n6053), .ZN(n9663) );
  INV_X1 U5886 ( .A(n9564), .ZN(n7437) );
  INV_X1 U5887 ( .A(n6969), .ZN(n7102) );
  NAND2_X1 U5888 ( .A1(n5731), .A2(n5730), .ZN(n9960) );
  NOR2_X1 U5889 ( .A1(n5729), .A2(P1_IR_REG_30__SCAN_IN), .ZN(n5730) );
  INV_X1 U5890 ( .A(n5727), .ZN(n5731) );
  INV_X1 U5892 ( .A(n6152), .ZN(n7408) );
  XNOR2_X1 U5893 ( .A(n5508), .B(n5507), .ZN(n7310) );
  INV_X1 U5894 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7306) );
  INV_X1 U5895 ( .A(n8015), .ZN(n7304) );
  INV_X1 U5896 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7190) );
  INV_X1 U5897 ( .A(n7757), .ZN(n7952) );
  INV_X1 U5898 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n9766) );
  INV_X1 U5899 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n9874) );
  NAND2_X1 U5900 ( .A1(n5719), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5720) );
  INV_X1 U5901 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6767) );
  INV_X1 U5902 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n9921) );
  INV_X1 U5903 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6598) );
  INV_X1 U5904 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6451) );
  INV_X1 U5905 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9869) );
  INV_X1 U5906 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9798) );
  INV_X1 U5907 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6348) );
  INV_X1 U5908 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6345) );
  INV_X1 U5909 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6336) );
  INV_X1 U5910 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9808) );
  AND2_X1 U5911 ( .A1(n4653), .A2(n4430), .ZN(n5240) );
  XNOR2_X1 U5912 ( .A(n4690), .B(n5769), .ZN(n6381) );
  NAND2_X1 U5913 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4690) );
  NOR2_X2 U5914 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n9972) );
  INV_X1 U5915 ( .A(n4645), .ZN(n8511) );
  NOR2_X1 U5916 ( .A1(n8540), .A2(n4857), .ZN(n4856) );
  OAI21_X1 U5917 ( .B1(n8539), .B2(n8562), .A(n10197), .ZN(n4858) );
  OAI22_X1 U5918 ( .A1(n8580), .A2(n8797), .B1(n10303), .B2(n6314), .ZN(n6315)
         );
  MUX2_X1 U5919 ( .A(n9572), .B(n9647), .S(n10186), .Z(n9573) );
  MUX2_X1 U5920 ( .A(n9926), .B(n9647), .S(n10174), .Z(n9648) );
  AND2_X1 U5921 ( .A1(n7879), .A2(n4399), .ZN(n4395) );
  AND2_X1 U5922 ( .A1(n4918), .A2(n4417), .ZN(n4396) );
  INV_X1 U5923 ( .A(n9221), .ZN(n7537) );
  INV_X2 U5924 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8913) );
  NAND2_X1 U5925 ( .A1(n9126), .A2(n9218), .ZN(n4399) );
  AND2_X1 U5926 ( .A1(n4693), .A2(n10154), .ZN(n4400) );
  AND2_X1 U5927 ( .A1(n4854), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4401) );
  AND2_X1 U5928 ( .A1(n4668), .A2(n5356), .ZN(n4402) );
  AND2_X1 U5929 ( .A1(n4972), .A2(n7535), .ZN(n4403) );
  AND2_X1 U5930 ( .A1(n4956), .A2(n7970), .ZN(n4404) );
  INV_X1 U5931 ( .A(n7168), .ZN(n7229) );
  NOR2_X1 U5932 ( .A1(n5643), .A2(n4601), .ZN(n4405) );
  OR2_X1 U5933 ( .A1(n9580), .A2(n4471), .ZN(n4406) );
  AND2_X1 U5934 ( .A1(n4697), .A2(n9946), .ZN(n4407) );
  AND2_X1 U5935 ( .A1(n4965), .A2(n4964), .ZN(n4408) );
  AND2_X1 U5936 ( .A1(n4854), .A2(n4853), .ZN(n4409) );
  OR2_X1 U5937 ( .A1(n5922), .A2(n5921), .ZN(n9221) );
  INV_X1 U5938 ( .A(n7348), .ZN(n4607) );
  OAI21_X1 U5939 ( .B1(n5673), .B2(n4619), .A(n4617), .ZN(n4616) );
  NAND2_X1 U5940 ( .A1(n4917), .A2(n4468), .ZN(n4410) );
  AND2_X1 U5941 ( .A1(n4400), .A2(n4692), .ZN(n4411) );
  OR2_X1 U5942 ( .A1(n6657), .A2(n6524), .ZN(n4412) );
  INV_X1 U5943 ( .A(n7440), .ZN(n4742) );
  AND4_X1 U5944 ( .A1(n5973), .A2(n5972), .A3(n5971), .A4(n5970), .ZN(n8920)
         );
  INV_X1 U5945 ( .A(n8920), .ZN(n4655) );
  AOI21_X1 U5946 ( .B1(n9076), .B2(n6098), .A(n6097), .ZN(n9372) );
  NAND2_X1 U5947 ( .A1(n5145), .A2(n5144), .ZN(n4413) );
  AND2_X1 U5948 ( .A1(n7304), .A2(n8005), .ZN(n7950) );
  NAND2_X1 U5949 ( .A1(n9965), .A2(n7744), .ZN(n5800) );
  NAND2_X2 U5950 ( .A1(n7744), .A2(n5747), .ZN(n5790) );
  AND2_X1 U5951 ( .A1(n8363), .A2(n4756), .ZN(n4414) );
  AND2_X1 U5952 ( .A1(n9006), .A2(n4747), .ZN(n4415) );
  OR2_X1 U5953 ( .A1(n6102), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n4416) );
  INV_X1 U5954 ( .A(n9532), .ZN(n4502) );
  NAND2_X1 U5955 ( .A1(n4861), .A2(n4859), .ZN(n5676) );
  AND2_X1 U5956 ( .A1(n4919), .A2(n4925), .ZN(n4417) );
  NAND3_X1 U5957 ( .A1(n4819), .A2(n4913), .A3(n4408), .ZN(n4418) );
  AND2_X1 U5958 ( .A1(n4786), .A2(n4784), .ZN(n4420) );
  NAND2_X1 U5959 ( .A1(n6614), .A2(n6607), .ZN(n7551) );
  INV_X2 U5960 ( .A(n5773), .ZN(n6106) );
  NOR2_X1 U5961 ( .A1(n7944), .A2(n7945), .ZN(n9370) );
  NOR2_X1 U5962 ( .A1(n6252), .A2(n4787), .ZN(n4421) );
  OR2_X1 U5963 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n4422) );
  NOR2_X1 U5964 ( .A1(n10272), .A2(n8405), .ZN(n4423) );
  NOR2_X1 U5965 ( .A1(n4393), .A2(n6505), .ZN(n4424) );
  INV_X1 U5966 ( .A(n7879), .ZN(n7973) );
  NAND2_X1 U5967 ( .A1(n7893), .A2(n7891), .ZN(n7879) );
  AND2_X1 U5968 ( .A1(n8060), .A2(n8077), .ZN(n8220) );
  OR2_X4 U5969 ( .A1(n7744), .A2(n5747), .ZN(n4979) );
  OAI21_X1 U5970 ( .B1(n8346), .B2(n4414), .A(n8345), .ZN(n8316) );
  OR2_X1 U5971 ( .A1(n8452), .A2(n8438), .ZN(n4425) );
  OR2_X1 U5972 ( .A1(n6131), .A2(n6705), .ZN(n4426) );
  INV_X1 U5973 ( .A(n8414), .ZN(n6188) );
  OR2_X1 U5974 ( .A1(n5190), .A2(n6490), .ZN(n4427) );
  OR2_X1 U5975 ( .A1(n9228), .A2(n7136), .ZN(n4428) );
  NAND2_X1 U5976 ( .A1(n7801), .A2(n7800), .ZN(n9360) );
  INV_X1 U5977 ( .A(n9360), .ZN(n9653) );
  INV_X1 U5978 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5285) );
  NAND2_X1 U5979 ( .A1(n5754), .A2(n5753), .ZN(n9531) );
  OAI21_X1 U5980 ( .B1(n9434), .B2(n6052), .A(n6051), .ZN(n9416) );
  AND3_X1 U5981 ( .A1(n4848), .A2(n4851), .A3(n6915), .ZN(n4429) );
  NAND2_X1 U5982 ( .A1(n5925), .A2(n5924), .ZN(n7561) );
  OR2_X1 U5983 ( .A1(n5067), .A2(n5219), .ZN(n4430) );
  OR2_X1 U5984 ( .A1(n6913), .A2(n6754), .ZN(n4431) );
  AND2_X1 U5985 ( .A1(n4884), .A2(n4795), .ZN(n4432) );
  NAND2_X1 U5986 ( .A1(n4819), .A2(n4913), .ZN(n6102) );
  INV_X1 U5987 ( .A(n4933), .ZN(n4932) );
  NAND2_X1 U5988 ( .A1(n5907), .A2(n5906), .ZN(n9049) );
  AND2_X1 U5989 ( .A1(n7829), .A2(n7947), .ZN(n4433) );
  AND2_X1 U5990 ( .A1(n4558), .A2(n4664), .ZN(n4434) );
  NAND2_X1 U5991 ( .A1(n4885), .A2(n4884), .ZN(n5005) );
  AND2_X1 U5992 ( .A1(n7986), .A2(n7950), .ZN(n4435) );
  INV_X1 U5993 ( .A(n6064), .ZN(n4924) );
  NAND2_X1 U5994 ( .A1(n9539), .A2(n4407), .ZN(n4698) );
  AND2_X1 U5995 ( .A1(n8056), .A2(n5276), .ZN(n4436) );
  AND2_X1 U5996 ( .A1(n9649), .A2(n9353), .ZN(n7982) );
  INV_X1 U5997 ( .A(n7982), .ZN(n4534) );
  NAND2_X1 U5998 ( .A1(n7736), .A2(n8742), .ZN(n4437) );
  INV_X1 U5999 ( .A(n8128), .ZN(n4599) );
  AND2_X1 U6000 ( .A1(n8417), .A2(n8416), .ZN(n4438) );
  AND2_X1 U6001 ( .A1(n7751), .A2(n7934), .ZN(n9394) );
  INV_X1 U6002 ( .A(n9394), .ZN(n4918) );
  OR2_X1 U6003 ( .A1(n7528), .A2(n7527), .ZN(n4439) );
  AND2_X1 U6004 ( .A1(n7882), .A2(n7880), .ZN(n7491) );
  INV_X1 U6005 ( .A(n9946), .ZN(n9504) );
  AND2_X1 U6006 ( .A1(n5999), .A2(n5998), .ZN(n9946) );
  OR2_X1 U6007 ( .A1(n8089), .A2(n8186), .ZN(n4440) );
  NAND3_X1 U6008 ( .A1(n4997), .A2(n9810), .A3(n4996), .ZN(n4441) );
  INV_X1 U6009 ( .A(n4699), .ZN(n9403) );
  NOR2_X1 U6010 ( .A1(n9452), .A2(n4700), .ZN(n4699) );
  AND2_X1 U6011 ( .A1(n8683), .A2(n8109), .ZN(n8703) );
  AND2_X1 U6012 ( .A1(n4974), .A2(P1_IR_REG_30__SCAN_IN), .ZN(n4442) );
  NAND2_X1 U6013 ( .A1(n10146), .A2(n7537), .ZN(n4961) );
  AND2_X1 U6014 ( .A1(n4627), .A2(n4629), .ZN(n4443) );
  INV_X1 U6015 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n9810) );
  NAND2_X1 U6016 ( .A1(n6066), .A2(n6065), .ZN(n9590) );
  INV_X1 U6017 ( .A(n6915), .ZN(n4853) );
  NOR2_X1 U6018 ( .A1(n7736), .A2(n8742), .ZN(n4444) );
  AND2_X1 U6019 ( .A1(n7343), .A2(n7537), .ZN(n7867) );
  INV_X1 U6020 ( .A(n7867), .ZN(n4810) );
  OR2_X1 U6021 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n4445) );
  AND2_X1 U6022 ( .A1(n7441), .A2(n7437), .ZN(n4446) );
  AND2_X1 U6023 ( .A1(n9803), .A2(n5031), .ZN(n4447) );
  NAND2_X1 U6024 ( .A1(n4885), .A2(n4432), .ZN(n4448) );
  AND2_X1 U6025 ( .A1(n4713), .A2(n7098), .ZN(n4449) );
  INV_X1 U6026 ( .A(n4793), .ZN(n4792) );
  NAND2_X1 U6027 ( .A1(n7203), .A2(n6213), .ZN(n4793) );
  AND2_X1 U6028 ( .A1(n8975), .A2(n8974), .ZN(n4450) );
  AND2_X1 U6029 ( .A1(n5103), .A2(SI_12_), .ZN(n4451) );
  INV_X1 U6030 ( .A(n4606), .ZN(n4605) );
  NAND2_X1 U6031 ( .A1(n4609), .A2(n4607), .ZN(n4606) );
  OR2_X1 U6032 ( .A1(n4868), .A2(n5411), .ZN(n4452) );
  AND2_X1 U6033 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4453) );
  INV_X1 U6034 ( .A(n10146), .ZN(n7343) );
  AND2_X1 U6035 ( .A1(n5915), .A2(n5914), .ZN(n10146) );
  INV_X1 U6036 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n9803) );
  OR2_X1 U6037 ( .A1(n4439), .A2(n4740), .ZN(n4454) );
  NAND2_X1 U6038 ( .A1(n7969), .A2(n4959), .ZN(n4455) );
  AND3_X1 U6039 ( .A1(n7889), .A2(n7887), .A3(n7888), .ZN(n4456) );
  AND2_X1 U6040 ( .A1(n4525), .A2(n9371), .ZN(n4457) );
  OR2_X1 U6041 ( .A1(n6361), .A2(n6467), .ZN(n4458) );
  NAND2_X1 U6042 ( .A1(n5593), .A2(n4993), .ZN(n5591) );
  INV_X1 U6043 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4964) );
  AND2_X1 U6044 ( .A1(n4946), .A2(n4945), .ZN(n4459) );
  AND2_X1 U6045 ( .A1(n7866), .A2(n7865), .ZN(n4460) );
  AND2_X1 U6046 ( .A1(n4738), .A2(n4737), .ZN(n4461) );
  NOR2_X1 U6047 ( .A1(n4445), .A2(n4966), .ZN(n4965) );
  INV_X1 U6048 ( .A(n9486), .ZN(n9942) );
  NAND2_X1 U6049 ( .A1(n6011), .A2(n6010), .ZN(n9486) );
  AND2_X1 U6050 ( .A1(n4806), .A2(n4442), .ZN(n4462) );
  AND2_X1 U6051 ( .A1(n4405), .A2(n8128), .ZN(n4463) );
  AND3_X1 U6052 ( .A1(n9809), .A2(n5716), .A3(n5718), .ZN(n4464) );
  OR2_X1 U6053 ( .A1(n7244), .A2(n7480), .ZN(n4465) );
  INV_X1 U6054 ( .A(n4785), .ZN(n4784) );
  NAND2_X1 U6055 ( .A1(n4788), .A2(n4789), .ZN(n4785) );
  INV_X1 U6056 ( .A(n4896), .ZN(n4895) );
  NAND2_X1 U6057 ( .A1(n4898), .A2(n4437), .ZN(n4896) );
  INV_X1 U6058 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n4808) );
  NAND2_X2 U6059 ( .A1(n8029), .A2(n8204), .ZN(n8186) );
  NAND2_X1 U6060 ( .A1(n5965), .A2(n5964), .ZN(n9202) );
  INV_X1 U6061 ( .A(n9202), .ZN(n4656) );
  AND2_X1 U6062 ( .A1(n8429), .A2(n8452), .ZN(n4466) );
  AOI22_X1 U6063 ( .A1(n7596), .A2(n7971), .B1(n7613), .B2(n7626), .ZN(n7628)
         );
  NAND2_X1 U6064 ( .A1(n7518), .A2(n8030), .ZN(n7665) );
  AND2_X1 U6065 ( .A1(n7925), .A2(n9435), .ZN(n9459) );
  INV_X1 U6066 ( .A(n9459), .ZN(n4491) );
  INV_X1 U6067 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4795) );
  INV_X1 U6068 ( .A(n9107), .ZN(n4748) );
  AND2_X1 U6069 ( .A1(n6437), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4467) );
  NAND2_X1 U6070 ( .A1(n7639), .A2(n4758), .ZN(n8324) );
  OR2_X1 U6071 ( .A1(n8846), .A2(n6273), .ZN(n8147) );
  NAND2_X1 U6072 ( .A1(n6092), .A2(n6091), .ZN(n9071) );
  NAND2_X1 U6073 ( .A1(n9658), .A2(n9187), .ZN(n4468) );
  NAND2_X1 U6074 ( .A1(n6044), .A2(n6043), .ZN(n9443) );
  INV_X1 U6075 ( .A(n9443), .ZN(n4703) );
  NAND2_X1 U6076 ( .A1(n4914), .A2(n4390), .ZN(n5974) );
  AND2_X1 U6077 ( .A1(n6260), .A2(n4753), .ZN(n4469) );
  AND2_X1 U6078 ( .A1(n8452), .A2(n8416), .ZN(n4470) );
  OR2_X1 U6079 ( .A1(n9504), .A2(n9060), .ZN(n9494) );
  INV_X1 U6080 ( .A(n9494), .ZN(n4817) );
  AND2_X1 U6081 ( .A1(n9581), .A2(n10165), .ZN(n4471) );
  INV_X1 U6082 ( .A(n8318), .ZN(n4772) );
  AND2_X1 U6083 ( .A1(n10051), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4472) );
  AND2_X1 U6084 ( .A1(n4951), .A2(n4949), .ZN(n4473) );
  INV_X1 U6085 ( .A(n8152), .ZN(n4619) );
  INV_X1 U6086 ( .A(n4771), .ZN(n4770) );
  NAND2_X1 U6087 ( .A1(n4774), .A2(n8345), .ZN(n4771) );
  NOR2_X1 U6088 ( .A1(n7589), .A2(n9219), .ZN(n4474) );
  INV_X1 U6089 ( .A(n5139), .ZN(n4545) );
  INV_X1 U6090 ( .A(n4757), .ZN(n4756) );
  NAND2_X1 U6091 ( .A1(n6263), .A2(n6264), .ZN(n4757) );
  OAI21_X1 U6092 ( .B1(n4866), .B2(n4545), .A(n5146), .ZN(n4544) );
  INV_X1 U6093 ( .A(n4921), .ZN(n4920) );
  NOR2_X1 U6094 ( .A1(n6079), .A2(n4922), .ZN(n4921) );
  INV_X1 U6095 ( .A(n8184), .ZN(n8580) );
  NAND2_X1 U6096 ( .A1(n5680), .A2(n5679), .ZN(n8184) );
  AND2_X1 U6097 ( .A1(n4773), .A2(n6274), .ZN(n4475) );
  NOR2_X1 U6098 ( .A1(n5997), .A2(n5996), .ZN(n4476) );
  OR3_X1 U6099 ( .A1(n6994), .A2(n6173), .A3(n6993), .ZN(n10173) );
  NAND2_X1 U6100 ( .A1(n7140), .A2(n4792), .ZN(n7202) );
  NAND2_X1 U6101 ( .A1(n5938), .A2(n5937), .ZN(n7589) );
  INV_X1 U6102 ( .A(n7589), .ZN(n4692) );
  NOR2_X1 U6103 ( .A1(n7820), .A2(n9967), .ZN(n4477) );
  XNOR2_X1 U6104 ( .A(n4840), .B(n7229), .ZN(n7152) );
  OR2_X1 U6105 ( .A1(n7179), .A2(n7178), .ZN(n4478) );
  INV_X1 U6106 ( .A(n8291), .ZN(n4782) );
  XNOR2_X1 U6107 ( .A(n5589), .B(n5588), .ZN(n5600) );
  NOR2_X1 U6108 ( .A1(n7226), .A2(n4844), .ZN(n4479) );
  NAND2_X1 U6109 ( .A1(n5320), .A2(n7348), .ZN(n7347) );
  AND2_X1 U6110 ( .A1(n4627), .A2(n4631), .ZN(n4480) );
  AND2_X1 U6111 ( .A1(n6946), .A2(n4721), .ZN(n4481) );
  NAND2_X1 U6112 ( .A1(n4885), .A2(n4794), .ZN(n4482) );
  INV_X1 U6113 ( .A(n4720), .ZN(n4719) );
  NAND2_X1 U6114 ( .A1(n4724), .A2(n7096), .ZN(n4720) );
  NAND2_X1 U6115 ( .A1(n6371), .A2(n6620), .ZN(n9373) );
  AND2_X1 U6116 ( .A1(n10189), .A2(n8551), .ZN(n10197) );
  AND2_X1 U6117 ( .A1(n7951), .A2(n8007), .ZN(n10087) );
  AND2_X1 U6118 ( .A1(n9261), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4483) );
  AND2_X1 U6119 ( .A1(n8533), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n4484) );
  INV_X1 U6120 ( .A(n6525), .ZN(n4836) );
  INV_X1 U6121 ( .A(n6986), .ZN(n10065) );
  OR2_X1 U6122 ( .A1(n6947), .A2(n6986), .ZN(n7760) );
  NOR2_X1 U6123 ( .A1(n7131), .A2(n6986), .ZN(n6980) );
  OR2_X1 U6124 ( .A1(n8430), .A2(n8452), .ZN(n4827) );
  OR2_X1 U6125 ( .A1(n8429), .A2(n8452), .ZN(n4828) );
  INV_X1 U6126 ( .A(n8452), .ZN(n4639) );
  NOR2_X1 U6127 ( .A1(n5272), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5286) );
  NOR2_X1 U6128 ( .A1(n7410), .A2(n7411), .ZN(n7415) );
  NAND2_X1 U6129 ( .A1(n4486), .A2(n4456), .ZN(n4490) );
  NAND4_X1 U6130 ( .A1(n7872), .A2(n7883), .A3(n7880), .A4(n7950), .ZN(n4486)
         );
  NAND2_X1 U6131 ( .A1(n4874), .A2(n4873), .ZN(n4878) );
  NAND2_X1 U6132 ( .A1(n4674), .A2(n4673), .ZN(n7941) );
  AOI21_X1 U6133 ( .B1(n7928), .B2(n7927), .A(n7926), .ZN(n4676) );
  INV_X1 U6134 ( .A(n6115), .ZN(n7859) );
  OAI21_X1 U6135 ( .B1(n8010), .B2(n4659), .A(n4658), .ZN(n4657) );
  XNOR2_X2 U6136 ( .A(n5313), .B(n5312), .ZN(n6354) );
  NAND2_X2 U6137 ( .A1(n7174), .A2(n7173), .ZN(n7440) );
  NAND2_X2 U6138 ( .A1(n8990), .A2(n9033), .ZN(n9138) );
  NAND2_X1 U6139 ( .A1(n9158), .A2(n9159), .ZN(n9157) );
  NAND2_X1 U6140 ( .A1(n9129), .A2(n9130), .ZN(n4744) );
  NAND2_X1 U6141 ( .A1(n9106), .A2(n9107), .ZN(n9179) );
  NAND2_X2 U6142 ( .A1(n8962), .A2(n9055), .ZN(n9149) );
  NAND2_X1 U6143 ( .A1(n4882), .A2(n4881), .ZN(n4873) );
  INV_X1 U6144 ( .A(n7941), .ZN(n7938) );
  NAND2_X1 U6145 ( .A1(n4489), .A2(n4460), .ZN(n7869) );
  NAND2_X1 U6146 ( .A1(n7864), .A2(n7863), .ZN(n4489) );
  NAND2_X1 U6147 ( .A1(n4657), .A2(n8016), .ZN(P1_U3242) );
  NAND2_X1 U6148 ( .A1(n4530), .A2(n8002), .ZN(n4529) );
  AOI21_X1 U6149 ( .B1(n4490), .B2(n7896), .A(n7895), .ZN(n7902) );
  AOI21_X2 U6150 ( .B1(n4492), .B2(n7947), .A(n4491), .ZN(n7928) );
  NAND2_X1 U6151 ( .A1(n7913), .A2(n7922), .ZN(n4492) );
  OR2_X1 U6152 ( .A1(n5768), .A2(n6328), .ZN(n5772) );
  AND2_X1 U6153 ( .A1(n7850), .A2(n7862), .ZN(n6115) );
  INV_X1 U6154 ( .A(n4497), .ZN(n6125) );
  INV_X1 U6155 ( .A(n4503), .ZN(n9457) );
  INV_X1 U6156 ( .A(n9469), .ZN(n4508) );
  AOI21_X1 U6157 ( .B1(n9395), .B2(n9394), .A(n6129), .ZN(n9369) );
  AOI21_X1 U6158 ( .B1(n9395), .B2(n4457), .A(n4516), .ZN(n4515) );
  OR2_X1 U6159 ( .A1(n5134), .A2(n4543), .ZN(n4541) );
  NAND2_X1 U6160 ( .A1(n5134), .A2(n4539), .ZN(n4538) );
  NAND2_X1 U6161 ( .A1(n5134), .A2(n4866), .ZN(n5472) );
  OAI21_X1 U6162 ( .B1(n5163), .B2(n4551), .A(n4549), .ZN(n5544) );
  INV_X1 U6163 ( .A(n4546), .ZN(n4861) );
  NAND2_X1 U6164 ( .A1(n5163), .A2(n5162), .ZN(n5532) );
  OR2_X1 U6165 ( .A1(n5106), .A2(n4555), .ZN(n4552) );
  NAND2_X1 U6166 ( .A1(n4552), .A2(n4553), .ZN(n4872) );
  NAND2_X1 U6167 ( .A1(n4559), .A2(n4434), .ZN(n4662) );
  NAND2_X1 U6168 ( .A1(n5300), .A2(n4561), .ZN(n4559) );
  NAND2_X1 U6169 ( .A1(n5299), .A2(n5088), .ZN(n4565) );
  OAI21_X2 U6170 ( .B1(n5300), .B2(n5299), .A(n5088), .ZN(n5313) );
  AND4_X2 U6171 ( .A1(n4750), .A2(n4751), .A3(n4987), .A4(n5204), .ZN(n4566)
         );
  NAND2_X1 U6172 ( .A1(n4566), .A2(n4398), .ZN(n5413) );
  NAND3_X2 U6173 ( .A1(n4566), .A2(n4398), .A3(n4749), .ZN(n5430) );
  OR2_X1 U6174 ( .A1(n8126), .A2(n4569), .ZN(n4567) );
  NAND3_X1 U6175 ( .A1(n4568), .A2(n4567), .A3(n4570), .ZN(n8134) );
  NAND3_X1 U6176 ( .A1(n5294), .A2(n5296), .A3(n4575), .ZN(n8407) );
  NAND4_X2 U6177 ( .A1(n4885), .A2(n4794), .A3(n4447), .A4(n4892), .ZN(n8914)
         );
  NAND3_X1 U6178 ( .A1(n4885), .A2(n4794), .A3(n4892), .ZN(n5033) );
  NAND2_X1 U6179 ( .A1(n5593), .A2(n4594), .ZN(n4589) );
  NAND2_X1 U6180 ( .A1(n5642), .A2(n4463), .ZN(n4596) );
  INV_X1 U6181 ( .A(n7474), .ZN(n5631) );
  AOI21_X1 U6182 ( .B1(n8600), .B2(n8147), .A(n8149), .ZN(n8592) );
  NAND2_X2 U6183 ( .A1(n6850), .A2(n6188), .ZN(n8042) );
  NAND2_X1 U6184 ( .A1(n7400), .A2(n4620), .ZN(n7518) );
  NAND2_X1 U6185 ( .A1(n4794), .A2(n4622), .ZN(n4994) );
  INV_X2 U6186 ( .A(n5430), .ZN(n4885) );
  OR2_X2 U6187 ( .A1(n7238), .A2(n7239), .ZN(n4631) );
  NAND2_X1 U6188 ( .A1(n6558), .A2(n6510), .ZN(n4635) );
  NAND2_X1 U6189 ( .A1(n6508), .A2(n6510), .ZN(n6556) );
  NOR2_X1 U6190 ( .A1(n8418), .A2(n8420), .ZN(n8453) );
  NAND2_X1 U6191 ( .A1(n4641), .A2(n7053), .ZN(n7051) );
  AND2_X2 U6192 ( .A1(n4645), .A2(n4644), .ZN(n8512) );
  AND2_X1 U6193 ( .A1(n4649), .A2(n4647), .ZN(n4646) );
  NAND3_X1 U6194 ( .A1(n4653), .A2(n4430), .A3(n5239), .ZN(n4654) );
  NAND2_X1 U6195 ( .A1(n5254), .A2(n5255), .ZN(n5075) );
  NAND2_X1 U6196 ( .A1(n4662), .A2(n4663), .ZN(n5106) );
  OAI21_X1 U6197 ( .B1(n5323), .B2(n4672), .A(n5096), .ZN(n5338) );
  OAI21_X1 U6198 ( .B1(n7928), .B2(n7914), .A(n7947), .ZN(n4675) );
  NAND4_X1 U6199 ( .A1(n4683), .A2(n4684), .A3(n9370), .A4(n4679), .ZN(n4678)
         );
  NAND3_X1 U6200 ( .A1(n7936), .A2(n7937), .A3(n7947), .ZN(n4683) );
  NAND2_X1 U6201 ( .A1(n7279), .A2(n4411), .ZN(n7597) );
  NAND2_X1 U6202 ( .A1(n4694), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6140) );
  NAND4_X1 U6203 ( .A1(n4819), .A2(n4913), .A3(n4695), .A4(n4408), .ZN(n4694)
         );
  INV_X1 U6204 ( .A(n4698), .ZN(n9503) );
  INV_X1 U6205 ( .A(n4704), .ZN(n6107) );
  NAND4_X2 U6206 ( .A1(n5818), .A2(n5787), .A3(n4706), .A4(n5700), .ZN(n5850)
         );
  NOR2_X4 U6207 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5787) );
  AND2_X2 U6208 ( .A1(n5806), .A2(n4705), .ZN(n5818) );
  INV_X2 U6209 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4705) );
  NAND3_X1 U6210 ( .A1(n5818), .A2(n5787), .A3(n4706), .ZN(n5848) );
  NAND3_X1 U6211 ( .A1(n4720), .A2(n4713), .A3(n4711), .ZN(n4710) );
  NAND2_X1 U6212 ( .A1(n9149), .A2(n4728), .ZN(n4725) );
  NAND2_X1 U6213 ( .A1(n4725), .A2(n4726), .ZN(n8979) );
  AND2_X4 U6214 ( .A1(n7551), .A2(n8997), .ZN(n8996) );
  NAND2_X1 U6215 ( .A1(n7440), .A2(n4461), .ZN(n4732) );
  NAND2_X2 U6216 ( .A1(n4732), .A2(n4734), .ZN(n7581) );
  NAND3_X1 U6217 ( .A1(n4736), .A2(n4738), .A3(n4737), .ZN(n4735) );
  NAND2_X1 U6218 ( .A1(n4744), .A2(n4743), .ZN(n9167) );
  NAND2_X1 U6219 ( .A1(n4744), .A2(n8949), .ZN(n8954) );
  NAND2_X2 U6220 ( .A1(n9138), .A2(n9139), .ZN(n9137) );
  AND2_X2 U6221 ( .A1(n5204), .A2(n4984), .ZN(n5205) );
  OAI21_X1 U6222 ( .B1(n4414), .B2(n4772), .A(n4764), .ZN(n4769) );
  NAND3_X1 U6223 ( .A1(n4762), .A2(n4475), .A3(n4760), .ZN(n6280) );
  NAND2_X1 U6224 ( .A1(n4768), .A2(n4769), .ZN(n8386) );
  INV_X1 U6225 ( .A(n8384), .ZN(n4767) );
  NAND2_X1 U6226 ( .A1(n7465), .A2(n4419), .ZN(n4775) );
  NAND2_X1 U6227 ( .A1(n4775), .A2(n4776), .ZN(n6236) );
  OAI21_X1 U6228 ( .B1(n6251), .B2(n4785), .A(n4781), .ZN(n6256) );
  NOR2_X2 U6229 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5900) );
  INV_X1 U6230 ( .A(n4796), .ZN(n9395) );
  NAND2_X1 U6231 ( .A1(n4805), .A2(n4462), .ZN(n4809) );
  OR2_X2 U6232 ( .A1(n5714), .A2(n4808), .ZN(n4805) );
  NAND2_X1 U6233 ( .A1(n5714), .A2(n5713), .ZN(n5727) );
  OAI211_X1 U6234 ( .C1(n7485), .C2(n4813), .A(n6123), .B(n4811), .ZN(n7623)
         );
  NAND2_X1 U6235 ( .A1(n6113), .A2(n6112), .ZN(n7834) );
  NAND3_X1 U6236 ( .A1(n4819), .A2(n4965), .A3(n4913), .ZN(n6142) );
  AND2_X2 U6237 ( .A1(n4914), .A2(n4464), .ZN(n4819) );
  NAND2_X1 U6238 ( .A1(n4913), .A2(n4914), .ZN(n5715) );
  NAND3_X1 U6239 ( .A1(n4827), .A2(n4828), .A3(n4825), .ZN(n8431) );
  NAND3_X1 U6240 ( .A1(n4827), .A2(n4826), .A3(n4825), .ZN(n4829) );
  INV_X1 U6241 ( .A(n4829), .ZN(n8439) );
  AOI21_X1 U6242 ( .B1(n6526), .B2(n10291), .A(n4836), .ZN(n4835) );
  OAI21_X1 U6243 ( .B1(n6526), .B2(n4836), .A(n4412), .ZN(n4831) );
  NAND2_X1 U6244 ( .A1(n4833), .A2(n4835), .ZN(n6658) );
  NAND2_X1 U6245 ( .A1(n6560), .A2(n6526), .ZN(n4833) );
  NAND2_X1 U6246 ( .A1(n4838), .A2(n4837), .ZN(n5206) );
  INV_X1 U6247 ( .A(n5204), .ZN(n4839) );
  INV_X1 U6248 ( .A(n7225), .ZN(n4840) );
  OAI211_X1 U6249 ( .C1(n6660), .C2(n4847), .A(n4846), .B(n4845), .ZN(n7057)
         );
  INV_X1 U6250 ( .A(n6660), .ZN(n4852) );
  NAND3_X1 U6251 ( .A1(n4858), .A2(n4856), .A3(n4855), .ZN(P2_U3200) );
  NAND2_X2 U6252 ( .A1(n5083), .A2(n5082), .ZN(n5300) );
  NAND2_X1 U6253 ( .A1(n5544), .A2(n5543), .ZN(n4862) );
  NAND2_X1 U6254 ( .A1(n5134), .A2(n5133), .ZN(n5455) );
  OAI21_X1 U6255 ( .B1(n7949), .B2(n9653), .A(n4875), .ZN(n4880) );
  OAI21_X1 U6256 ( .B1(n7949), .B2(n9360), .A(n4876), .ZN(n4882) );
  NAND2_X1 U6257 ( .A1(n8006), .A2(n8005), .ZN(n4877) );
  NAND3_X1 U6258 ( .A1(n4398), .A2(n5205), .A3(n4883), .ZN(n5414) );
  NAND2_X1 U6259 ( .A1(n6954), .A2(n8216), .ZN(n4886) );
  NAND2_X1 U6260 ( .A1(n7347), .A2(n4887), .ZN(n5336) );
  NAND3_X1 U6261 ( .A1(n4890), .A2(n5231), .A3(n4889), .ZN(n6821) );
  NAND2_X1 U6262 ( .A1(n5230), .A2(n4891), .ZN(n4889) );
  NAND3_X1 U6263 ( .A1(n5215), .A2(n5230), .A3(n5625), .ZN(n4890) );
  NAND2_X1 U6264 ( .A1(n8760), .A2(n5216), .ZN(n6857) );
  NAND2_X1 U6265 ( .A1(n5215), .A2(n5625), .ZN(n8760) );
  INV_X1 U6266 ( .A(n5216), .ZN(n4891) );
  OAI21_X1 U6267 ( .B1(n7513), .B2(n4896), .A(n4893), .ZN(n8740) );
  NAND2_X1 U6268 ( .A1(n5442), .A2(n5470), .ZN(n4905) );
  NAND2_X2 U6269 ( .A1(n4905), .A2(n4903), .ZN(n8659) );
  NAND2_X1 U6270 ( .A1(n8705), .A2(n5453), .ZN(n8704) );
  INV_X1 U6271 ( .A(n5442), .ZN(n8705) );
  OR2_X2 U6272 ( .A1(n5560), .A2(n5559), .ZN(n4909) );
  NAND2_X1 U6273 ( .A1(n4910), .A2(n5827), .ZN(n6979) );
  NAND3_X1 U6274 ( .A1(n4428), .A2(n5811), .A3(n4912), .ZN(n4910) );
  AND2_X2 U6275 ( .A1(n5707), .A2(n5708), .ZN(n4913) );
  NAND2_X1 U6276 ( .A1(n9416), .A2(n4921), .ZN(n4916) );
  INV_X1 U6277 ( .A(n9416), .ZN(n4915) );
  NAND3_X1 U6278 ( .A1(n4918), .A2(n4417), .A3(n4920), .ZN(n4917) );
  OR2_X1 U6279 ( .A1(n5997), .A2(n4928), .ZN(n4927) );
  NOR2_X1 U6280 ( .A1(n9518), .A2(n9175), .ZN(n4933) );
  NAND2_X1 U6281 ( .A1(n7031), .A2(n4935), .ZN(n4934) );
  INV_X1 U6282 ( .A(n7628), .ZN(n4952) );
  NAND2_X1 U6283 ( .A1(n7628), .A2(n4459), .ZN(n4940) );
  NAND2_X1 U6284 ( .A1(n7329), .A2(n4404), .ZN(n4954) );
  INV_X1 U6285 ( .A(n9071), .ZN(n9362) );
  NOR2_X4 U6286 ( .A1(n5206), .A2(n5205), .ZN(n6519) );
  NAND2_X1 U6287 ( .A1(n9972), .A2(n5052), .ZN(n5054) );
  NAND2_X1 U6288 ( .A1(n5461), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5212) );
  NAND3_X1 U6289 ( .A1(n5000), .A2(n5032), .A3(n4999), .ZN(n5001) );
  OR2_X1 U6290 ( .A1(n5593), .A2(n5585), .ZN(n5586) );
  INV_X1 U6291 ( .A(n8914), .ZN(n5035) );
  NAND2_X1 U6292 ( .A1(n4391), .A2(n6325), .ZN(n5188) );
  OR2_X1 U6293 ( .A1(n6305), .A2(n6304), .ZN(P2_U3154) );
  NAND2_X1 U6294 ( .A1(n8293), .A2(n6259), .ZN(n8362) );
  NAND2_X1 U6295 ( .A1(n5672), .A2(n4976), .ZN(P2_U3205) );
  INV_X1 U6296 ( .A(n9590), .ZN(n9408) );
  NAND2_X1 U6297 ( .A1(n9376), .A2(n9653), .ZN(n9356) );
  INV_X1 U6298 ( .A(n7745), .ZN(n5040) );
  OR2_X1 U6299 ( .A1(n8612), .A2(n8601), .ZN(n8603) );
  NAND2_X1 U6300 ( .A1(n8940), .A2(n8939), .ZN(n9129) );
  AND2_X2 U6301 ( .A1(n6185), .A2(n6184), .ZN(n6191) );
  NAND2_X1 U6302 ( .A1(n8954), .A2(n8953), .ZN(n9168) );
  INV_X1 U6303 ( .A(n6142), .ZN(n5714) );
  AOI21_X1 U6304 ( .B1(n8576), .B2(n10279), .A(n8577), .ZN(n6313) );
  NAND2_X1 U6305 ( .A1(n8260), .A2(n5040), .ZN(n5190) );
  INV_X1 U6306 ( .A(n8260), .ZN(n5041) );
  XNOR2_X1 U6307 ( .A(n6191), .B(n6186), .ZN(n6189) );
  INV_X1 U6308 ( .A(n10303), .ZN(n6312) );
  AND2_X2 U6309 ( .A1(n6995), .A2(n9559), .ZN(n10102) );
  INV_X2 U6310 ( .A(n10102), .ZN(n9562) );
  AND2_X1 U6311 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n4969) );
  OR2_X1 U6312 ( .A1(n5768), .A2(n6327), .ZN(n4971) );
  AND2_X1 U6313 ( .A1(n6238), .A2(n7507), .ZN(n4973) );
  NAND2_X2 U6314 ( .A1(n6167), .A2(n6146), .ZN(n6614) );
  NAND2_X1 U6315 ( .A1(n5554), .A2(n5553), .ZN(n8587) );
  INV_X1 U6316 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5031) );
  NAND2_X1 U6317 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), 
        .ZN(n4974) );
  INV_X1 U6318 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5867) );
  AND2_X1 U6319 ( .A1(n5671), .A2(n5670), .ZN(n4976) );
  AND2_X1 U6320 ( .A1(n5649), .A2(n5648), .ZN(n4977) );
  OR2_X1 U6321 ( .A1(n10287), .A2(n10274), .ZN(n8842) );
  INV_X1 U6322 ( .A(n8842), .ZN(n5698) );
  INV_X2 U6323 ( .A(n10287), .ZN(n10286) );
  INV_X1 U6324 ( .A(n5747), .ZN(n9965) );
  INV_X1 U6325 ( .A(n8703), .ZN(n5453) );
  INV_X1 U6326 ( .A(n8087), .ZN(n5633) );
  INV_X1 U6327 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n4985) );
  INV_X1 U6328 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n4991) );
  INV_X1 U6329 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5709) );
  INV_X1 U6330 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4996) );
  NAND2_X1 U6331 ( .A1(n6181), .A2(n6180), .ZN(n6185) );
  INV_X1 U6332 ( .A(n9372), .ZN(n9363) );
  AND2_X1 U6333 ( .A1(n5712), .A2(n4964), .ZN(n5713) );
  INV_X1 U6334 ( .A(n7468), .ZN(n6222) );
  NAND2_X1 U6335 ( .A1(n8573), .A2(n8835), .ZN(n8196) );
  INV_X1 U6336 ( .A(n5447), .ZN(n5019) );
  INV_X1 U6337 ( .A(n5305), .ZN(n5013) );
  OAI21_X1 U6338 ( .B1(n5599), .B2(P2_D_REG_0__SCAN_IN), .A(n6397), .ZN(n6178)
         );
  NAND2_X1 U6339 ( .A1(n5210), .A2(n5209), .ZN(n5211) );
  AND2_X1 U6340 ( .A1(n5592), .A2(n4996), .ZN(n4993) );
  INV_X1 U6341 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5892) );
  NAND2_X1 U6342 ( .A1(n7534), .A2(n7533), .ZN(n7535) );
  INV_X1 U6343 ( .A(n8953), .ZN(n8951) );
  OR3_X1 U6344 ( .A1(n6055), .A2(n9142), .A3(n9109), .ZN(n6068) );
  INV_X1 U6345 ( .A(n6025), .ZN(n6023) );
  INV_X1 U6346 ( .A(n5991), .ZN(n5744) );
  INV_X1 U6347 ( .A(n5877), .ZN(n5739) );
  AND2_X1 U6348 ( .A1(n5471), .A2(n5473), .ZN(n5139) );
  INV_X1 U6349 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5716) );
  INV_X1 U6350 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n5113) );
  INV_X1 U6351 ( .A(SI_11_), .ZN(n5097) );
  INV_X1 U6352 ( .A(n8587), .ZN(n6273) );
  INV_X1 U6353 ( .A(n6191), .ZN(n6197) );
  OR2_X1 U6354 ( .A1(n5655), .A2(n5653), .ZN(n6296) );
  OR2_X1 U6355 ( .A1(n5571), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5573) );
  NAND2_X1 U6356 ( .A1(n8913), .A2(n9803), .ZN(n4999) );
  INV_X1 U6357 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n9783) );
  AND2_X1 U6358 ( .A1(n8846), .A2(n6273), .ZN(n8149) );
  INV_X1 U6359 ( .A(n5480), .ZN(n5021) );
  NAND2_X1 U6360 ( .A1(n5345), .A2(n5014), .ZN(n5378) );
  NAND2_X1 U6361 ( .A1(n6853), .A2(n8048), .ZN(n5625) );
  INV_X1 U6362 ( .A(n8742), .ZN(n7507) );
  AND2_X1 U6363 ( .A1(n5618), .A2(n8203), .ZN(n5647) );
  OR2_X1 U6364 ( .A1(n5341), .A2(n5340), .ZN(n5358) );
  AND2_X1 U6365 ( .A1(n6634), .A2(n6633), .ZN(n6635) );
  OR2_X1 U6366 ( .A1(n8936), .A2(n9118), .ZN(n8938) );
  INV_X1 U6367 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7085) );
  NAND2_X1 U6368 ( .A1(n6000), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6012) );
  INV_X1 U6369 ( .A(n7998), .ZN(n6620) );
  INV_X1 U6370 ( .A(n5399), .ZN(n5117) );
  INV_X1 U6371 ( .A(n8714), .ZN(n8692) );
  INV_X1 U6372 ( .A(n8390), .ZN(n8376) );
  INV_X1 U6373 ( .A(n8743), .ZN(n7644) );
  OR2_X1 U6374 ( .A1(n8783), .A2(n8752), .ZN(n5671) );
  NAND2_X1 U6375 ( .A1(n5027), .A2(n5026), .ZN(n5547) );
  OR2_X1 U6376 ( .A1(n5464), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5480) );
  AND2_X1 U6377 ( .A1(n8051), .A2(n8039), .ZN(n8211) );
  INV_X1 U6378 ( .A(n8651), .ZN(n8630) );
  OR2_X1 U6379 ( .A1(n8720), .A2(n8721), .ZN(n8718) );
  INV_X1 U6380 ( .A(n8216), .ZN(n6956) );
  AND2_X1 U6381 ( .A1(n5616), .A2(n5583), .ZN(n8629) );
  OR2_X1 U6382 ( .A1(n7608), .A2(n7607), .ZN(n7609) );
  OR2_X1 U6383 ( .A1(n8981), .A2(n8980), .ZN(n8982) );
  NOR2_X1 U6384 ( .A1(n6635), .A2(n6698), .ZN(n6640) );
  NAND2_X1 U6385 ( .A1(n6033), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6055) );
  INV_X1 U6386 ( .A(n9145), .ZN(n9198) );
  INV_X1 U6387 ( .A(n5800), .ZN(n6133) );
  INV_X1 U6388 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6876) );
  NAND2_X1 U6389 ( .A1(n7937), .A2(n9367), .ZN(n9368) );
  INV_X1 U6390 ( .A(n10164), .ZN(n7613) );
  NAND2_X1 U6391 ( .A1(n9562), .A2(n6998), .ZN(n10096) );
  INV_X1 U6392 ( .A(n9383), .ZN(n9581) );
  INV_X1 U6393 ( .A(n7561), .ZN(n10154) );
  OAI21_X1 U6394 ( .B1(n6600), .B2(P1_D_REG_1__SCAN_IN), .A(n9958), .ZN(n6992)
         );
  NAND2_X1 U6395 ( .A1(n5725), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5726) );
  AND2_X1 U6396 ( .A1(n5127), .A2(n5126), .ZN(n5427) );
  XNOR2_X1 U6397 ( .A(n5114), .B(SI_15_), .ZN(n5399) );
  AND2_X1 U6398 ( .A1(n5093), .A2(n5092), .ZN(n5312) );
  NAND2_X1 U6399 ( .A1(n5011), .A2(n5010), .ZN(n5291) );
  NAND2_X1 U6400 ( .A1(n6288), .A2(n6286), .ZN(n8392) );
  INV_X1 U6401 ( .A(n6729), .ZN(n6733) );
  AND2_X1 U6402 ( .A1(n6288), .A2(n6287), .ZN(n8390) );
  INV_X1 U6403 ( .A(n8392), .ZN(n8372) );
  NAND2_X1 U6404 ( .A1(n6709), .A2(n8243), .ZN(n8394) );
  NAND2_X1 U6405 ( .A1(n6283), .A2(n8771), .ZN(n8379) );
  AND2_X1 U6406 ( .A1(n5542), .A2(n5541), .ZN(n8631) );
  INV_X1 U6407 ( .A(n10192), .ZN(n10212) );
  INV_X2 U6408 ( .A(n6488), .ZN(n8551) );
  OR2_X1 U6409 ( .A1(n8028), .A2(n6306), .ZN(n8771) );
  INV_X1 U6410 ( .A(n8771), .ZN(n8748) );
  INV_X1 U6411 ( .A(n8797), .ZN(n8826) );
  NAND2_X1 U6412 ( .A1(n7302), .A2(n8241), .ZN(n10274) );
  INV_X1 U6413 ( .A(n8209), .ZN(n8739) );
  NAND2_X1 U6414 ( .A1(n7479), .A2(n10268), .ZN(n10279) );
  INV_X1 U6415 ( .A(n5599), .ZN(n6364) );
  NAND2_X1 U6416 ( .A1(n6501), .A2(n6708), .ZN(n8028) );
  AND2_X1 U6417 ( .A1(n5317), .A2(n5324), .ZN(n7168) );
  AND2_X1 U6418 ( .A1(n7311), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6321) );
  AND4_X1 U6419 ( .A1(n5983), .A2(n5982), .A3(n5981), .A4(n5980), .ZN(n9132)
         );
  OR2_X1 U6420 ( .A1(n9321), .A2(n9320), .ZN(n9332) );
  XNOR2_X1 U6421 ( .A(n9356), .B(n9649), .ZN(n9349) );
  OR2_X1 U6422 ( .A1(n6099), .A2(n9368), .ZN(n6100) );
  INV_X1 U6423 ( .A(n10087), .ZN(n10072) );
  INV_X1 U6424 ( .A(n9540), .ZN(n10094) );
  OAI21_X1 U6425 ( .B1(n6600), .B2(P1_D_REG_0__SCAN_IN), .A(n9959), .ZN(n6602)
         );
  NAND2_X1 U6426 ( .A1(n7330), .A2(n10168), .ZN(n10161) );
  NAND2_X1 U6427 ( .A1(n6155), .A2(n6167), .ZN(n6600) );
  AND2_X1 U6428 ( .A1(n5913), .A2(n5935), .ZN(n6872) );
  INV_X1 U6429 ( .A(n8394), .ZN(n8339) );
  AND2_X1 U6430 ( .A1(n6279), .A2(n6278), .ZN(n8381) );
  INV_X1 U6431 ( .A(n8379), .ZN(n8397) );
  NAND2_X1 U6432 ( .A1(n5580), .A2(n5579), .ZN(n8588) );
  INV_X1 U6433 ( .A(n8308), .ZN(n8402) );
  OR2_X1 U6434 ( .A1(P2_U3150), .A2(n6502), .ZN(n10192) );
  INV_X1 U6435 ( .A(n10197), .ZN(n10229) );
  OR2_X1 U6436 ( .A1(n6514), .A2(n8551), .ZN(n10220) );
  AND2_X1 U6437 ( .A1(n5668), .A2(n8771), .ZN(n8725) );
  NAND2_X1 U6438 ( .A1(n5669), .A2(n8769), .ZN(n8595) );
  NAND2_X1 U6439 ( .A1(n10303), .A2(n10279), .ZN(n8829) );
  AND3_X2 U6440 ( .A1(n6311), .A2(n6310), .A3(n6309), .ZN(n10303) );
  AOI21_X1 U6441 ( .B1(n8184), .B2(n5698), .A(n5697), .ZN(n5699) );
  OR2_X1 U6442 ( .A1(n10287), .A2(n10247), .ZN(n8910) );
  AND2_X1 U6443 ( .A1(n5622), .A2(n5621), .ZN(n10287) );
  NOR2_X1 U6444 ( .A1(n6364), .A2(n8028), .ZN(n6573) );
  INV_X1 U6445 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7303) );
  INV_X1 U6446 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6596) );
  INV_X1 U6447 ( .A(n9201), .ZN(n9191) );
  INV_X1 U6448 ( .A(n9184), .ZN(n9204) );
  NAND2_X1 U6449 ( .A1(n6078), .A2(n6077), .ZN(n9209) );
  OR2_X1 U6450 ( .A1(n5761), .A2(n5760), .ZN(n9216) );
  OR2_X1 U6451 ( .A1(n10041), .A2(n10031), .ZN(n9336) );
  INV_X1 U6452 ( .A(n10081), .ZN(n10097) );
  NAND2_X1 U6453 ( .A1(n9562), .A2(n6996), .ZN(n9557) );
  AOI21_X1 U6454 ( .B1(n6176), .B2(n10186), .A(n6175), .ZN(n6177) );
  NAND2_X1 U6455 ( .A1(n10186), .A2(n10165), .ZN(n9646) );
  INV_X2 U6456 ( .A(n10184), .ZN(n10186) );
  INV_X1 U6457 ( .A(n9389), .ZN(n9658) );
  INV_X1 U6458 ( .A(n9531), .ZN(n9951) );
  AND2_X1 U6459 ( .A1(n10151), .A2(n10150), .ZN(n10181) );
  INV_X2 U6460 ( .A(n10173), .ZN(n10174) );
  INV_X1 U6461 ( .A(n10116), .ZN(n10118) );
  NAND2_X1 U6462 ( .A1(n8013), .A2(n6600), .ZN(n10116) );
  INV_X1 U6463 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6883) );
  INV_X1 U6464 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6393) );
  INV_X1 U6465 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10311) );
  INV_X1 U6466 ( .A(n8527), .ZN(P2_U3893) );
  OAI21_X1 U6467 ( .B1(n6313), .B2(n10287), .A(n5699), .ZN(P2_U3456) );
  NAND2_X1 U6468 ( .A1(n5650), .A2(n4977), .ZN(P2_U3455) );
  INV_X1 U6469 ( .A(n6177), .ZN(P1_U3550) );
  INV_X1 U6470 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n5623) );
  INV_X1 U6471 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n4992) );
  NAND2_X2 U6472 ( .A1(n4994), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5593) );
  NAND2_X1 U6473 ( .A1(n5585), .A2(n5588), .ZN(n4995) );
  NAND2_X1 U6474 ( .A1(n4995), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5592) );
  INV_X1 U6475 ( .A(n4995), .ZN(n4997) );
  NAND2_X1 U6476 ( .A1(n5033), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4998) );
  OR2_X1 U6477 ( .A1(n4998), .A2(n9803), .ZN(n5000) );
  INV_X1 U6478 ( .A(n8026), .ZN(n6497) );
  INV_X1 U6479 ( .A(n5002), .ZN(n6488) );
  NAND2_X1 U6480 ( .A1(n6497), .A2(n6488), .ZN(n5003) );
  AND2_X1 U6481 ( .A1(n5184), .A2(n5003), .ZN(n6287) );
  NAND2_X1 U6482 ( .A1(n4448), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5004) );
  NAND2_X1 U6483 ( .A1(n5005), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5006) );
  INV_X1 U6484 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5007) );
  NAND2_X1 U6485 ( .A1(n5007), .A2(n6860), .ZN(n5248) );
  INV_X1 U6486 ( .A(n5248), .ZN(n5009) );
  NAND2_X1 U6487 ( .A1(n5009), .A2(n5008), .ZN(n5263) );
  INV_X1 U6488 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5014) );
  INV_X1 U6489 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5016) );
  NOR2_X1 U6490 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_REG3_REG_18__SCAN_IN), 
        .ZN(n5018) );
  INV_X1 U6491 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n5020) );
  INV_X1 U6492 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5022) );
  INV_X1 U6493 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5024) );
  INV_X1 U6494 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5026) );
  INV_X1 U6495 ( .A(n5549), .ZN(n5029) );
  INV_X1 U6496 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5028) );
  NAND2_X1 U6497 ( .A1(n5029), .A2(n5028), .ZN(n5571) );
  NAND2_X1 U6498 ( .A1(n5549), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5030) );
  NAND2_X1 U6499 ( .A1(n5571), .A2(n5030), .ZN(n8593) );
  XNOR2_X2 U6500 ( .A(n5039), .B(n5038), .ZN(n8260) );
  NAND2_X1 U6501 ( .A1(n5040), .A2(n5041), .ZN(n5191) );
  NAND2_X1 U6502 ( .A1(n8593), .A2(n5574), .ZN(n5046) );
  INV_X1 U6503 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9900) );
  NAND2_X1 U6504 ( .A1(n5575), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5043) );
  AND2_X2 U6505 ( .A1(n8260), .A2(n7745), .ZN(n5189) );
  INV_X2 U6506 ( .A(n5189), .ZN(n5234) );
  NAND2_X1 U6507 ( .A1(n5189), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5042) );
  OAI211_X1 U6508 ( .C1(n8179), .C2(n9900), .A(n5043), .B(n5042), .ZN(n5044)
         );
  INV_X1 U6509 ( .A(n5044), .ZN(n5045) );
  NAND2_X1 U6510 ( .A1(n8571), .A2(n5574), .ZN(n8182) );
  INV_X1 U6511 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6314) );
  NAND2_X1 U6512 ( .A1(n5575), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5049) );
  NAND2_X1 U6513 ( .A1(n5189), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5048) );
  OAI211_X1 U6514 ( .C1(n8179), .C2(n6314), .A(n5049), .B(n5048), .ZN(n5050)
         );
  INV_X1 U6515 ( .A(n5050), .ZN(n5051) );
  INV_X1 U6516 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6328) );
  INV_X1 U6517 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6331) );
  AND2_X1 U6518 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5055) );
  NAND2_X1 U6519 ( .A1(n7813), .A2(n5055), .ZN(n5198) );
  INV_X2 U6520 ( .A(n5062), .ZN(n5779) );
  AND2_X1 U6521 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5056) );
  NAND2_X1 U6522 ( .A1(n5779), .A2(n5056), .ZN(n5782) );
  NAND2_X1 U6523 ( .A1(n5198), .A2(n5782), .ZN(n5182) );
  INV_X1 U6524 ( .A(n5057), .ZN(n5058) );
  NAND2_X1 U6525 ( .A1(n5058), .A2(SI_1_), .ZN(n5059) );
  INV_X1 U6526 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6327) );
  INV_X1 U6527 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6323) );
  MUX2_X1 U6528 ( .A(n6327), .B(n6323), .S(n5062), .Z(n5060) );
  XNOR2_X1 U6529 ( .A(n5060), .B(SI_2_), .ZN(n5208) );
  NAND2_X1 U6530 ( .A1(n5207), .A2(n5208), .ZN(n5218) );
  INV_X1 U6531 ( .A(n5060), .ZN(n5061) );
  NAND2_X1 U6532 ( .A1(n5061), .A2(SI_2_), .ZN(n5217) );
  INV_X4 U6533 ( .A(n5062), .ZN(n6325) );
  INV_X1 U6534 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6324) );
  INV_X1 U6535 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6342) );
  INV_X1 U6536 ( .A(n5066), .ZN(n5064) );
  NAND2_X1 U6537 ( .A1(n5064), .A2(SI_3_), .ZN(n5065) );
  AND2_X1 U6538 ( .A1(n5217), .A2(n5065), .ZN(n5068) );
  INV_X1 U6539 ( .A(n5065), .ZN(n5067) );
  XNOR2_X1 U6540 ( .A(n5066), .B(SI_3_), .ZN(n5219) );
  INV_X1 U6541 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6329) );
  INV_X1 U6542 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6339) );
  MUX2_X1 U6543 ( .A(n6329), .B(n6339), .S(n6325), .Z(n5069) );
  XNOR2_X1 U6544 ( .A(n5069), .B(SI_4_), .ZN(n5239) );
  INV_X1 U6545 ( .A(n5069), .ZN(n5070) );
  NAND2_X1 U6546 ( .A1(n5070), .A2(SI_4_), .ZN(n5071) );
  INV_X1 U6547 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6330) );
  XNOR2_X1 U6548 ( .A(n5072), .B(SI_5_), .ZN(n5255) );
  INV_X1 U6549 ( .A(n5072), .ZN(n5073) );
  NAND2_X1 U6550 ( .A1(n5073), .A2(SI_5_), .ZN(n5074) );
  NAND2_X1 U6551 ( .A1(n5075), .A2(n5074), .ZN(n5270) );
  MUX2_X1 U6552 ( .A(n6333), .B(n6336), .S(n6325), .Z(n5076) );
  XNOR2_X1 U6553 ( .A(n5076), .B(SI_6_), .ZN(n5271) );
  NAND2_X1 U6554 ( .A1(n5270), .A2(n5271), .ZN(n5079) );
  INV_X1 U6555 ( .A(n5076), .ZN(n5077) );
  NAND2_X1 U6556 ( .A1(n5077), .A2(SI_6_), .ZN(n5078) );
  NAND2_X1 U6557 ( .A1(n5079), .A2(n5078), .ZN(n5283) );
  MUX2_X1 U6558 ( .A(n6343), .B(n6345), .S(n5779), .Z(n5080) );
  XNOR2_X1 U6559 ( .A(n5080), .B(SI_7_), .ZN(n5284) );
  NAND2_X1 U6560 ( .A1(n5283), .A2(n5284), .ZN(n5083) );
  INV_X1 U6561 ( .A(n5080), .ZN(n5081) );
  NAND2_X1 U6562 ( .A1(n5081), .A2(SI_7_), .ZN(n5082) );
  MUX2_X1 U6563 ( .A(n9733), .B(n6348), .S(n6325), .Z(n5085) );
  INV_X1 U6564 ( .A(SI_8_), .ZN(n5084) );
  NAND2_X1 U6565 ( .A1(n5085), .A2(n5084), .ZN(n5088) );
  INV_X1 U6566 ( .A(n5085), .ZN(n5086) );
  NAND2_X1 U6567 ( .A1(n5086), .A2(SI_8_), .ZN(n5087) );
  NAND2_X1 U6568 ( .A1(n5088), .A2(n5087), .ZN(n5299) );
  MUX2_X1 U6569 ( .A(n6356), .B(n9798), .S(n6325), .Z(n5090) );
  NAND2_X1 U6570 ( .A1(n5090), .A2(n5089), .ZN(n5093) );
  INV_X1 U6571 ( .A(n5090), .ZN(n5091) );
  NAND2_X1 U6572 ( .A1(n5091), .A2(SI_9_), .ZN(n5092) );
  MUX2_X1 U6573 ( .A(n6359), .B(n9869), .S(n6325), .Z(n5094) );
  XNOR2_X1 U6574 ( .A(n5094), .B(SI_10_), .ZN(n5322) );
  INV_X1 U6575 ( .A(n5094), .ZN(n5095) );
  NAND2_X1 U6576 ( .A1(n5095), .A2(SI_10_), .ZN(n5096) );
  MUX2_X1 U6577 ( .A(n6395), .B(n6393), .S(n5779), .Z(n5098) );
  INV_X1 U6578 ( .A(n5098), .ZN(n5099) );
  NAND2_X1 U6579 ( .A1(n5099), .A2(SI_11_), .ZN(n5100) );
  NAND2_X1 U6580 ( .A1(n5101), .A2(n5100), .ZN(n5337) );
  MUX2_X1 U6581 ( .A(n6453), .B(n6451), .S(n6325), .Z(n5102) );
  XNOR2_X1 U6582 ( .A(n5102), .B(SI_12_), .ZN(n5356) );
  INV_X1 U6583 ( .A(n5102), .ZN(n5103) );
  MUX2_X1 U6584 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6325), .Z(n5104) );
  XNOR2_X1 U6585 ( .A(n5104), .B(SI_13_), .ZN(n5372) );
  NAND2_X1 U6586 ( .A1(n5104), .A2(SI_13_), .ZN(n5105) );
  MUX2_X1 U6587 ( .A(n6596), .B(n6598), .S(n6325), .Z(n5108) );
  NAND2_X1 U6588 ( .A1(n5108), .A2(n5107), .ZN(n5111) );
  INV_X1 U6589 ( .A(n5108), .ZN(n5109) );
  NAND2_X1 U6590 ( .A1(n5109), .A2(SI_14_), .ZN(n5110) );
  NAND2_X1 U6591 ( .A1(n5111), .A2(n5110), .ZN(n5384) );
  MUX2_X1 U6592 ( .A(n5113), .B(n9921), .S(n5779), .Z(n5114) );
  INV_X1 U6593 ( .A(n5114), .ZN(n5115) );
  NAND2_X1 U6594 ( .A1(n5115), .A2(SI_15_), .ZN(n5116) );
  MUX2_X1 U6595 ( .A(n9732), .B(n6767), .S(n5779), .Z(n5119) );
  INV_X1 U6596 ( .A(SI_16_), .ZN(n5118) );
  NAND2_X1 U6597 ( .A1(n5119), .A2(n5118), .ZN(n5122) );
  INV_X1 U6598 ( .A(n5119), .ZN(n5120) );
  NAND2_X1 U6599 ( .A1(n5120), .A2(SI_16_), .ZN(n5121) );
  NAND2_X1 U6600 ( .A1(n5122), .A2(n5121), .ZN(n5411) );
  MUX2_X1 U6601 ( .A(n6865), .B(n6883), .S(n6325), .Z(n5124) );
  INV_X1 U6602 ( .A(SI_17_), .ZN(n5123) );
  NAND2_X1 U6603 ( .A1(n5124), .A2(n5123), .ZN(n5127) );
  INV_X1 U6604 ( .A(n5124), .ZN(n5125) );
  NAND2_X1 U6605 ( .A1(n5125), .A2(SI_17_), .ZN(n5126) );
  NAND2_X1 U6606 ( .A1(n5428), .A2(n5427), .ZN(n5128) );
  NAND2_X1 U6607 ( .A1(n5128), .A2(n5127), .ZN(n5444) );
  INV_X1 U6608 ( .A(n5444), .ZN(n5130) );
  INV_X1 U6609 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n5129) );
  MUX2_X1 U6610 ( .A(n6930), .B(n5129), .S(n5779), .Z(n5131) );
  XNOR2_X1 U6611 ( .A(n5131), .B(SI_18_), .ZN(n5443) );
  NAND2_X1 U6612 ( .A1(n5130), .A2(n5443), .ZN(n5134) );
  INV_X1 U6613 ( .A(n5131), .ZN(n5132) );
  NAND2_X1 U6614 ( .A1(n5132), .A2(SI_18_), .ZN(n5133) );
  MUX2_X1 U6615 ( .A(n7008), .B(n9874), .S(n5779), .Z(n5136) );
  INV_X1 U6616 ( .A(SI_19_), .ZN(n5135) );
  NAND2_X1 U6617 ( .A1(n5136), .A2(n5135), .ZN(n5471) );
  INV_X1 U6618 ( .A(n5136), .ZN(n5137) );
  NAND2_X1 U6619 ( .A1(n5137), .A2(SI_19_), .ZN(n5138) );
  NAND2_X1 U6620 ( .A1(n5471), .A2(n5138), .ZN(n5454) );
  MUX2_X1 U6621 ( .A(n9924), .B(n9766), .S(n6325), .Z(n5140) );
  INV_X1 U6622 ( .A(SI_20_), .ZN(n9884) );
  NAND2_X1 U6623 ( .A1(n5140), .A2(n9884), .ZN(n5473) );
  INV_X1 U6624 ( .A(n5140), .ZN(n5141) );
  NAND2_X1 U6625 ( .A1(n5141), .A2(SI_20_), .ZN(n5486) );
  MUX2_X1 U6626 ( .A(n9776), .B(n7190), .S(n6325), .Z(n5143) );
  INV_X1 U6627 ( .A(n5143), .ZN(n5142) );
  NAND2_X1 U6628 ( .A1(n5142), .A2(SI_21_), .ZN(n5145) );
  XNOR2_X1 U6629 ( .A(n5143), .B(SI_21_), .ZN(n5488) );
  INV_X1 U6630 ( .A(n5488), .ZN(n5144) );
  MUX2_X1 U6631 ( .A(n7303), .B(n7306), .S(n6325), .Z(n5148) );
  INV_X1 U6632 ( .A(SI_22_), .ZN(n5147) );
  NAND2_X1 U6633 ( .A1(n5148), .A2(n5147), .ZN(n5151) );
  INV_X1 U6634 ( .A(n5148), .ZN(n5149) );
  NAND2_X1 U6635 ( .A1(n5149), .A2(SI_22_), .ZN(n5150) );
  NAND2_X1 U6636 ( .A1(n5151), .A2(n5150), .ZN(n5497) );
  INV_X1 U6637 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7313) );
  MUX2_X1 U6638 ( .A(n9756), .B(n7313), .S(n6325), .Z(n5153) );
  INV_X1 U6639 ( .A(SI_23_), .ZN(n5152) );
  NAND2_X1 U6640 ( .A1(n5153), .A2(n5152), .ZN(n5156) );
  INV_X1 U6641 ( .A(n5153), .ZN(n5154) );
  NAND2_X1 U6642 ( .A1(n5154), .A2(SI_23_), .ZN(n5155) );
  NAND2_X1 U6643 ( .A1(n5508), .A2(n5507), .ZN(n5157) );
  NAND2_X1 U6644 ( .A1(n5157), .A2(n5156), .ZN(n5519) );
  INV_X1 U6645 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7381) );
  INV_X1 U6646 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7379) );
  MUX2_X1 U6647 ( .A(n7381), .B(n7379), .S(n6325), .Z(n5159) );
  INV_X1 U6648 ( .A(SI_24_), .ZN(n5158) );
  NAND2_X1 U6649 ( .A1(n5159), .A2(n5158), .ZN(n5162) );
  INV_X1 U6650 ( .A(n5159), .ZN(n5160) );
  NAND2_X1 U6651 ( .A1(n5160), .A2(SI_24_), .ZN(n5161) );
  NAND2_X1 U6652 ( .A1(n5519), .A2(n5518), .ZN(n5163) );
  INV_X1 U6653 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7458) );
  INV_X1 U6654 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n9923) );
  MUX2_X1 U6655 ( .A(n7458), .B(n9923), .S(n5779), .Z(n5164) );
  NAND2_X1 U6656 ( .A1(n5164), .A2(n9753), .ZN(n5167) );
  INV_X1 U6657 ( .A(n5164), .ZN(n5165) );
  NAND2_X1 U6658 ( .A1(n5165), .A2(SI_25_), .ZN(n5166) );
  INV_X1 U6659 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7522) );
  INV_X1 U6660 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7501) );
  MUX2_X1 U6661 ( .A(n7522), .B(n7501), .S(n5779), .Z(n5168) );
  INV_X1 U6662 ( .A(SI_26_), .ZN(n9915) );
  NAND2_X1 U6663 ( .A1(n5168), .A2(n9915), .ZN(n5171) );
  INV_X1 U6664 ( .A(n5168), .ZN(n5169) );
  NAND2_X1 U6665 ( .A1(n5169), .A2(SI_26_), .ZN(n5170) );
  INV_X1 U6666 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5172) );
  INV_X1 U6667 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7635) );
  MUX2_X1 U6668 ( .A(n5172), .B(n7635), .S(n6325), .Z(n5173) );
  INV_X1 U6669 ( .A(SI_27_), .ZN(n9764) );
  NAND2_X1 U6670 ( .A1(n5173), .A2(n9764), .ZN(n5563) );
  INV_X1 U6671 ( .A(n5173), .ZN(n5174) );
  NAND2_X1 U6672 ( .A1(n5174), .A2(SI_27_), .ZN(n5175) );
  INV_X2 U6673 ( .A(n5290), .ZN(n5176) );
  NAND2_X1 U6674 ( .A1(n7564), .A2(n5176), .ZN(n5178) );
  NAND2_X1 U6675 ( .A1(n5461), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5177) );
  INV_X1 U6676 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6490) );
  INV_X1 U6677 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6734) );
  OR2_X1 U6678 ( .A1(n5191), .A2(n6734), .ZN(n5181) );
  INV_X1 U6679 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6849) );
  NAND2_X1 U6680 ( .A1(n5189), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5179) );
  NAND4_X2 U6681 ( .A1(n4427), .A2(n5181), .A3(n5180), .A4(n5179), .ZN(n8414)
         );
  XNOR2_X1 U6682 ( .A(n5183), .B(n5182), .ZN(n6332) );
  NAND2_X1 U6683 ( .A1(n5210), .A2(n6332), .ZN(n5187) );
  INV_X1 U6684 ( .A(n5184), .ZN(n5185) );
  OAI211_X1 U6685 ( .C1(n5188), .C2(P1_DATAO_REG_1__SCAN_IN), .A(n5187), .B(
        n5186), .ZN(n6186) );
  INV_X1 U6686 ( .A(n6186), .ZN(n6850) );
  NAND2_X1 U6687 ( .A1(n8414), .A2(n6186), .ZN(n8040) );
  NAND2_X1 U6688 ( .A1(n5189), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5195) );
  INV_X1 U6689 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6515) );
  OR2_X1 U6690 ( .A1(n5190), .A2(n6515), .ZN(n5194) );
  INV_X1 U6691 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6717) );
  OR2_X1 U6692 ( .A1(n4393), .A2(n6717), .ZN(n5193) );
  INV_X1 U6693 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6712) );
  OR2_X1 U6694 ( .A1(n5191), .A2(n6712), .ZN(n5192) );
  INV_X1 U6695 ( .A(n6844), .ZN(n8415) );
  NAND2_X1 U6696 ( .A1(n7813), .A2(SI_0_), .ZN(n5197) );
  INV_X1 U6697 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5196) );
  NAND2_X1 U6698 ( .A1(n5197), .A2(n5196), .ZN(n5199) );
  AND2_X1 U6699 ( .A1(n5199), .A2(n5198), .ZN(n8919) );
  MUX2_X1 U6700 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8919), .S(n5184), .Z(n6684) );
  NAND2_X1 U6701 ( .A1(n8415), .A2(n6684), .ZN(n6843) );
  NAND2_X1 U6702 ( .A1(n6187), .A2(n6186), .ZN(n8756) );
  NAND2_X1 U6703 ( .A1(n8758), .A2(n8756), .ZN(n5215) );
  INV_X1 U6704 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9705) );
  INV_X1 U6705 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6505) );
  INV_X1 U6706 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6728) );
  OR2_X1 U6707 ( .A1(n5435), .A2(n6728), .ZN(n5201) );
  NAND3_X2 U6708 ( .A1(n5203), .A2(n5202), .A3(n5201), .ZN(n8413) );
  NAND2_X1 U6709 ( .A1(n5460), .A2(n6519), .ZN(n5214) );
  XNOR2_X1 U6710 ( .A(n5207), .B(n5208), .ZN(n6326) );
  INV_X1 U6711 ( .A(n6326), .ZN(n5209) );
  INV_X1 U6712 ( .A(n10240), .ZN(n6720) );
  NAND2_X1 U6713 ( .A1(n6720), .A2(n8413), .ZN(n8048) );
  NAND2_X1 U6714 ( .A1(n6845), .A2(n6720), .ZN(n5216) );
  NAND2_X1 U6715 ( .A1(n5218), .A2(n5217), .ZN(n5220) );
  XNOR2_X1 U6716 ( .A(n5220), .B(n5219), .ZN(n6341) );
  NAND2_X1 U6717 ( .A1(n5461), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5224) );
  NOR2_X1 U6718 ( .A1(n5205), .A2(n8913), .ZN(n5221) );
  NAND2_X1 U6719 ( .A1(n5205), .A2(n5222), .ZN(n5256) );
  NAND2_X1 U6720 ( .A1(n5460), .A2(n6567), .ZN(n5223) );
  OAI211_X1 U6721 ( .C1(n5290), .C2(n6341), .A(n5224), .B(n5223), .ZN(n6861)
         );
  INV_X1 U6722 ( .A(n6861), .ZN(n10246) );
  INV_X2 U6723 ( .A(n8179), .ZN(n5537) );
  NAND2_X1 U6724 ( .A1(n5537), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5229) );
  INV_X1 U6725 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6859) );
  OR2_X1 U6726 ( .A1(n5200), .A2(n6859), .ZN(n5228) );
  OR2_X1 U6727 ( .A1(n5435), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5227) );
  INV_X1 U6728 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5225) );
  OR2_X1 U6729 ( .A1(n5234), .A2(n5225), .ZN(n5226) );
  AND4_X2 U6730 ( .A1(n5229), .A2(n5228), .A3(n5227), .A4(n5226), .ZN(n8763)
         );
  OR2_X1 U6731 ( .A1(n10246), .A2(n8763), .ZN(n5230) );
  NAND2_X1 U6732 ( .A1(n8763), .A2(n10246), .ZN(n5231) );
  NAND2_X1 U6733 ( .A1(n5537), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5238) );
  INV_X1 U6734 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6651) );
  OR2_X1 U6735 ( .A1(n5200), .A2(n6651), .ZN(n5237) );
  NAND2_X1 U6736 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5232) );
  AND2_X1 U6737 ( .A1(n5248), .A2(n5232), .ZN(n6972) );
  OR2_X1 U6738 ( .A1(n5435), .A2(n6972), .ZN(n5236) );
  INV_X1 U6739 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5233) );
  OR2_X1 U6740 ( .A1(n5234), .A2(n5233), .ZN(n5235) );
  XNOR2_X1 U6741 ( .A(n5240), .B(n5239), .ZN(n6338) );
  NAND2_X1 U6742 ( .A1(n5461), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5243) );
  NAND2_X1 U6743 ( .A1(n5256), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5241) );
  NAND2_X1 U6744 ( .A1(n5460), .A2(n6657), .ZN(n5242) );
  OAI211_X1 U6745 ( .C1(n5290), .C2(n6338), .A(n5243), .B(n5242), .ZN(n6833)
         );
  OR2_X1 U6746 ( .A1(n6901), .A2(n6833), .ZN(n8067) );
  NAND2_X1 U6747 ( .A1(n6901), .A2(n6833), .ZN(n8052) );
  NAND2_X1 U6748 ( .A1(n8067), .A2(n8052), .ZN(n6818) );
  NAND2_X1 U6749 ( .A1(n6821), .A2(n6818), .ZN(n5245) );
  INV_X1 U6750 ( .A(n6833), .ZN(n6973) );
  NAND2_X1 U6751 ( .A1(n6901), .A2(n6973), .ZN(n5244) );
  NAND2_X1 U6752 ( .A1(n5245), .A2(n5244), .ZN(n6899) );
  NAND2_X1 U6753 ( .A1(n5189), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5253) );
  INV_X1 U6754 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5246) );
  OR2_X1 U6755 ( .A1(n8179), .A2(n5246), .ZN(n5252) );
  INV_X1 U6756 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n5247) );
  OR2_X1 U6757 ( .A1(n5200), .A2(n5247), .ZN(n5251) );
  NAND2_X1 U6758 ( .A1(n5248), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5249) );
  AND2_X1 U6759 ( .A1(n5263), .A2(n5249), .ZN(n6933) );
  OR2_X1 U6760 ( .A1(n5435), .A2(n6933), .ZN(n5250) );
  NAND4_X1 U6761 ( .A1(n5253), .A2(n5252), .A3(n5251), .A4(n5250), .ZN(n8410)
         );
  XNOR2_X1 U6762 ( .A(n5254), .B(n5255), .ZN(n6340) );
  NAND2_X1 U6763 ( .A1(n5461), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5259) );
  NAND2_X1 U6764 ( .A1(n5272), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5257) );
  XNOR2_X1 U6765 ( .A(n5257), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6743) );
  NAND2_X1 U6766 ( .A1(n5460), .A2(n6743), .ZN(n5258) );
  OAI211_X1 U6767 ( .C1(n5290), .C2(n6340), .A(n5259), .B(n5258), .ZN(n6902)
         );
  NOR2_X1 U6768 ( .A1(n8410), .A2(n6902), .ZN(n5261) );
  NAND2_X1 U6769 ( .A1(n8410), .A2(n6902), .ZN(n5260) );
  OAI21_X2 U6770 ( .B1(n6899), .B2(n5261), .A(n5260), .ZN(n6954) );
  NAND2_X1 U6771 ( .A1(n5537), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5269) );
  INV_X1 U6772 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n5262) );
  OR2_X1 U6773 ( .A1(n5200), .A2(n5262), .ZN(n5268) );
  NAND2_X1 U6774 ( .A1(n5263), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5264) );
  AND2_X1 U6775 ( .A1(n5277), .A2(n5264), .ZN(n7148) );
  OR2_X1 U6776 ( .A1(n5435), .A2(n7148), .ZN(n5267) );
  INV_X1 U6777 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5265) );
  OR2_X1 U6778 ( .A1(n5234), .A2(n5265), .ZN(n5266) );
  XNOR2_X1 U6779 ( .A(n5270), .B(n5271), .ZN(n6335) );
  NAND2_X1 U6780 ( .A1(n5461), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n5275) );
  OR2_X1 U6781 ( .A1(n5286), .A2(n8913), .ZN(n5273) );
  XNOR2_X1 U6782 ( .A(n5273), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6913) );
  NAND2_X1 U6783 ( .A1(n5460), .A2(n6913), .ZN(n5274) );
  OAI211_X1 U6784 ( .C1(n5290), .C2(n6335), .A(n5275), .B(n5274), .ZN(n7145)
         );
  OR2_X1 U6785 ( .A1(n7207), .A2(n7145), .ZN(n8074) );
  NAND2_X1 U6786 ( .A1(n7207), .A2(n7145), .ZN(n8072) );
  NAND2_X1 U6787 ( .A1(n8074), .A2(n8072), .ZN(n8216) );
  INV_X1 U6788 ( .A(n7145), .ZN(n10252) );
  OR2_X1 U6789 ( .A1(n10252), .A2(n7207), .ZN(n5276) );
  NAND2_X1 U6790 ( .A1(n5189), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5282) );
  INV_X1 U6791 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6909) );
  OR2_X1 U6792 ( .A1(n5200), .A2(n6909), .ZN(n5281) );
  NAND2_X1 U6793 ( .A1(n5277), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5278) );
  AND2_X1 U6794 ( .A1(n5291), .A2(n5278), .ZN(n7212) );
  OR2_X1 U6795 ( .A1(n5435), .A2(n7212), .ZN(n5280) );
  INV_X1 U6796 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6908) );
  OR2_X1 U6797 ( .A1(n8179), .A2(n6908), .ZN(n5279) );
  XNOR2_X1 U6798 ( .A(n5283), .B(n5284), .ZN(n6344) );
  NAND2_X1 U6799 ( .A1(n5461), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n5289) );
  NAND2_X1 U6800 ( .A1(n5286), .A2(n5285), .ZN(n5297) );
  NAND2_X1 U6801 ( .A1(n5297), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5287) );
  XNOR2_X1 U6802 ( .A(n5287), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6915) );
  NAND2_X1 U6803 ( .A1(n5460), .A2(n6915), .ZN(n5288) );
  OAI211_X1 U6804 ( .C1(n5290), .C2(n6344), .A(n5289), .B(n5288), .ZN(n7199)
         );
  OR2_X1 U6805 ( .A1(n6215), .A2(n7199), .ZN(n8060) );
  NAND2_X1 U6806 ( .A1(n6215), .A2(n7199), .ZN(n8077) );
  INV_X1 U6807 ( .A(n7199), .ZN(n10255) );
  NAND2_X1 U6808 ( .A1(n6215), .A2(n10255), .ZN(n7215) );
  NAND2_X1 U6809 ( .A1(n7216), .A2(n7215), .ZN(n5303) );
  NAND2_X1 U6810 ( .A1(n5537), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5296) );
  INV_X1 U6811 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7219) );
  OR2_X1 U6812 ( .A1(n5200), .A2(n7219), .ZN(n5295) );
  NAND2_X1 U6813 ( .A1(n5291), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5292) );
  AND2_X1 U6814 ( .A1(n5305), .A2(n5292), .ZN(n7318) );
  OR2_X1 U6815 ( .A1(n5435), .A2(n7318), .ZN(n5294) );
  INV_X1 U6816 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5293) );
  NAND2_X1 U6817 ( .A1(n5341), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5298) );
  NAND2_X1 U6818 ( .A1(n6346), .A2(n5176), .ZN(n5302) );
  NAND2_X1 U6819 ( .A1(n5461), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n5301) );
  OAI211_X1 U6820 ( .C1(n5184), .C2(n7160), .A(n5302), .B(n5301), .ZN(n7326)
         );
  NAND2_X1 U6821 ( .A1(n6219), .A2(n7326), .ZN(n8078) );
  INV_X1 U6822 ( .A(n7326), .ZN(n10261) );
  NAND2_X1 U6823 ( .A1(n10261), .A2(n8407), .ZN(n8059) );
  NAND2_X1 U6824 ( .A1(n8078), .A2(n8059), .ZN(n7221) );
  NAND2_X1 U6825 ( .A1(n5303), .A2(n7221), .ZN(n7214) );
  NAND2_X1 U6826 ( .A1(n6219), .A2(n10261), .ZN(n7349) );
  NAND2_X1 U6827 ( .A1(n7214), .A2(n7349), .ZN(n5320) );
  NAND2_X1 U6828 ( .A1(n5537), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5311) );
  INV_X1 U6829 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n5304) );
  OR2_X1 U6830 ( .A1(n5200), .A2(n5304), .ZN(n5310) );
  NAND2_X1 U6831 ( .A1(n5305), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5306) );
  AND2_X1 U6832 ( .A1(n5329), .A2(n5306), .ZN(n7461) );
  OR2_X1 U6833 ( .A1(n5435), .A2(n7461), .ZN(n5309) );
  INV_X1 U6834 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5307) );
  OR2_X1 U6835 ( .A1(n5234), .A2(n5307), .ZN(n5308) );
  NAND4_X1 U6836 ( .A1(n5311), .A2(n5310), .A3(n5309), .A4(n5308), .ZN(n8406)
         );
  NAND2_X1 U6837 ( .A1(n6354), .A2(n5176), .ZN(n5319) );
  NAND2_X1 U6838 ( .A1(n5314), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5316) );
  INV_X1 U6839 ( .A(n5316), .ZN(n5315) );
  NAND2_X1 U6840 ( .A1(n5315), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5317) );
  NAND2_X1 U6841 ( .A1(n5316), .A2(n9747), .ZN(n5324) );
  AOI22_X1 U6842 ( .A1(n5461), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5460), .B2(
        n7168), .ZN(n5318) );
  NAND2_X1 U6843 ( .A1(n5319), .A2(n5318), .ZN(n10267) );
  NAND2_X1 U6844 ( .A1(n10267), .A2(n7314), .ZN(n8079) );
  NAND2_X1 U6845 ( .A1(n8064), .A2(n8079), .ZN(n7348) );
  OR2_X1 U6846 ( .A1(n10267), .A2(n8406), .ZN(n5321) );
  XNOR2_X1 U6847 ( .A(n5323), .B(n5322), .ZN(n6357) );
  NAND2_X1 U6848 ( .A1(n6357), .A2(n5176), .ZN(n5327) );
  NAND2_X1 U6849 ( .A1(n5324), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5325) );
  XNOR2_X1 U6850 ( .A(n5325), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7244) );
  AOI22_X1 U6851 ( .A1(n5461), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5460), .B2(
        n7244), .ZN(n5326) );
  NAND2_X1 U6852 ( .A1(n5189), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5334) );
  INV_X1 U6853 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n5328) );
  OR2_X1 U6854 ( .A1(n8179), .A2(n5328), .ZN(n5333) );
  INV_X1 U6855 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7480) );
  OR2_X1 U6856 ( .A1(n5200), .A2(n7480), .ZN(n5332) );
  NAND2_X1 U6857 ( .A1(n5329), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5330) );
  AND2_X1 U6858 ( .A1(n5346), .A2(n5330), .ZN(n7677) );
  OR2_X1 U6859 ( .A1(n5435), .A2(n7677), .ZN(n5331) );
  NAND2_X1 U6860 ( .A1(n10272), .A2(n8405), .ZN(n5335) );
  NAND2_X1 U6861 ( .A1(n5336), .A2(n5335), .ZN(n7395) );
  XNOR2_X1 U6862 ( .A(n5338), .B(n5337), .ZN(n6392) );
  NAND2_X1 U6863 ( .A1(n6392), .A2(n5176), .ZN(n5344) );
  INV_X1 U6864 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5339) );
  NAND3_X1 U6865 ( .A1(n9815), .A2(n9747), .A3(n5339), .ZN(n5340) );
  NAND2_X1 U6866 ( .A1(n5358), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5342) );
  XNOR2_X1 U6867 ( .A(n5342), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7424) );
  AOI22_X1 U6868 ( .A1(n5461), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5460), .B2(
        n7424), .ZN(n5343) );
  NAND2_X1 U6869 ( .A1(n5344), .A2(n5343), .ZN(n7401) );
  NAND2_X1 U6870 ( .A1(n5537), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5352) );
  INV_X1 U6871 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7360) );
  OR2_X1 U6872 ( .A1(n5200), .A2(n7360), .ZN(n5351) );
  INV_X1 U6873 ( .A(n5345), .ZN(n5362) );
  NAND2_X1 U6874 ( .A1(n5346), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5347) );
  AND2_X1 U6875 ( .A1(n5362), .A2(n5347), .ZN(n7402) );
  OR2_X1 U6876 ( .A1(n5435), .A2(n7402), .ZN(n5350) );
  INV_X1 U6877 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n5348) );
  OR2_X1 U6878 ( .A1(n5234), .A2(n5348), .ZN(n5349) );
  OR2_X1 U6879 ( .A1(n7401), .A2(n8404), .ZN(n5353) );
  NAND2_X1 U6880 ( .A1(n7395), .A2(n5353), .ZN(n5355) );
  NAND2_X1 U6881 ( .A1(n7401), .A2(n8404), .ZN(n5354) );
  NAND2_X2 U6882 ( .A1(n5355), .A2(n5354), .ZN(n7513) );
  XNOR2_X1 U6883 ( .A(n5357), .B(n5356), .ZN(n6450) );
  NAND2_X1 U6884 ( .A1(n6450), .A2(n5176), .ZN(n5361) );
  NOR2_X1 U6885 ( .A1(n5358), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n5374) );
  OR2_X1 U6886 ( .A1(n5374), .A2(n8913), .ZN(n5359) );
  XNOR2_X1 U6887 ( .A(n5359), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7427) );
  AOI22_X1 U6888 ( .A1(n5461), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5460), .B2(
        n7427), .ZN(n5360) );
  NAND2_X1 U6889 ( .A1(n5537), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5368) );
  INV_X1 U6890 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7428) );
  OR2_X1 U6891 ( .A1(n5200), .A2(n7428), .ZN(n5367) );
  NAND2_X1 U6892 ( .A1(n5362), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5363) );
  AND2_X1 U6893 ( .A1(n5378), .A2(n5363), .ZN(n8312) );
  OR2_X1 U6894 ( .A1(n5435), .A2(n8312), .ZN(n5366) );
  INV_X1 U6895 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n5364) );
  OR2_X1 U6896 ( .A1(n5234), .A2(n5364), .ZN(n5365) );
  NAND4_X1 U6897 ( .A1(n5368), .A2(n5367), .A3(n5366), .A4(n5365), .ZN(n8403)
         );
  AND2_X1 U6898 ( .A1(n10282), .A2(n8403), .ZN(n5370) );
  OR2_X1 U6899 ( .A1(n10282), .A2(n8403), .ZN(n5369) );
  XNOR2_X1 U6900 ( .A(n5371), .B(n5372), .ZN(n6570) );
  NAND2_X1 U6901 ( .A1(n6570), .A2(n5176), .ZN(n5377) );
  INV_X1 U6902 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5373) );
  NAND2_X1 U6903 ( .A1(n5374), .A2(n5373), .ZN(n5375) );
  NAND2_X1 U6904 ( .A1(n5375), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5387) );
  XNOR2_X1 U6905 ( .A(n5387), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8452) );
  AOI22_X1 U6906 ( .A1(n5461), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5460), .B2(
        n8452), .ZN(n5376) );
  NAND2_X1 U6907 ( .A1(n5189), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5383) );
  INV_X1 U6908 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8420) );
  OR2_X1 U6909 ( .A1(n5200), .A2(n8420), .ZN(n5382) );
  INV_X1 U6910 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9752) );
  OR2_X1 U6911 ( .A1(n8179), .A2(n9752), .ZN(n5381) );
  NAND2_X1 U6912 ( .A1(n5378), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5379) );
  AND2_X1 U6913 ( .A1(n5393), .A2(n5379), .ZN(n7714) );
  OR2_X1 U6914 ( .A1(n5435), .A2(n7714), .ZN(n5380) );
  NOR2_X1 U6915 ( .A1(n7713), .A2(n8402), .ZN(n7668) );
  NAND2_X1 U6916 ( .A1(n7713), .A2(n8402), .ZN(n7666) );
  XNOR2_X1 U6917 ( .A(n5385), .B(n5384), .ZN(n6595) );
  NAND2_X1 U6918 ( .A1(n6595), .A2(n5176), .ZN(n5392) );
  INV_X1 U6919 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5386) );
  NAND2_X1 U6920 ( .A1(n5387), .A2(n5386), .ZN(n5388) );
  NAND2_X1 U6921 ( .A1(n5388), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5389) );
  INV_X1 U6922 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n9771) );
  NAND2_X1 U6923 ( .A1(n5389), .A2(n9771), .ZN(n5400) );
  OR2_X1 U6924 ( .A1(n5389), .A2(n9771), .ZN(n5390) );
  AOI22_X1 U6925 ( .A1(n5461), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5460), .B2(
        n8455), .ZN(n5391) );
  NAND2_X1 U6926 ( .A1(n5189), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5398) );
  INV_X1 U6927 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8440) );
  OR2_X1 U6928 ( .A1(n8179), .A2(n8440), .ZN(n5397) );
  INV_X1 U6929 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n9911) );
  OR2_X1 U6930 ( .A1(n5200), .A2(n9911), .ZN(n5396) );
  NAND2_X1 U6931 ( .A1(n5393), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5394) );
  AND2_X1 U6932 ( .A1(n5404), .A2(n5394), .ZN(n7726) );
  OR2_X1 U6933 ( .A1(n5435), .A2(n7726), .ZN(n5395) );
  NAND4_X1 U6934 ( .A1(n5398), .A2(n5397), .A3(n5396), .A4(n5395), .ZN(n8742)
         );
  NAND2_X1 U6935 ( .A1(n6690), .A2(n5176), .ZN(n5403) );
  NAND2_X1 U6936 ( .A1(n5400), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5401) );
  XNOR2_X1 U6937 ( .A(n5401), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8499) );
  AOI22_X1 U6938 ( .A1(n5461), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5460), .B2(
        n8499), .ZN(n5402) );
  NAND2_X1 U6939 ( .A1(n5189), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5409) );
  INV_X1 U6940 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8825) );
  OR2_X1 U6941 ( .A1(n8179), .A2(n8825), .ZN(n5408) );
  INV_X1 U6942 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8746) );
  OR2_X1 U6943 ( .A1(n4393), .A2(n8746), .ZN(n5407) );
  NAND2_X1 U6944 ( .A1(n5404), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5405) );
  AND2_X1 U6945 ( .A1(n5419), .A2(n5405), .ZN(n7642) );
  OR2_X1 U6946 ( .A1(n5435), .A2(n7642), .ZN(n5406) );
  NAND4_X1 U6947 ( .A1(n5409), .A2(n5408), .A3(n5407), .A4(n5406), .ZN(n8730)
         );
  NOR2_X1 U6948 ( .A1(n8907), .A2(n8730), .ZN(n5410) );
  INV_X1 U6949 ( .A(n8730), .ZN(n7570) );
  INV_X1 U6950 ( .A(n8907), .ZN(n7648) );
  OAI22_X2 U6951 ( .A1(n8740), .A2(n5410), .B1(n7570), .B2(n7648), .ZN(n8729)
         );
  XNOR2_X1 U6952 ( .A(n5412), .B(n5411), .ZN(n6765) );
  NAND2_X1 U6953 ( .A1(n6765), .A2(n5176), .ZN(n5418) );
  NAND2_X1 U6954 ( .A1(n5414), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5415) );
  MUX2_X1 U6955 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5415), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n5416) );
  AND2_X1 U6956 ( .A1(n5413), .A2(n5416), .ZN(n8502) );
  AOI22_X1 U6957 ( .A1(n5461), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5460), .B2(
        n8502), .ZN(n5417) );
  NAND2_X1 U6958 ( .A1(n5189), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5424) );
  INV_X1 U6959 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8822) );
  OR2_X1 U6960 ( .A1(n8179), .A2(n8822), .ZN(n5423) );
  INV_X1 U6961 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8733) );
  OR2_X1 U6962 ( .A1(n5200), .A2(n8733), .ZN(n5422) );
  NAND2_X1 U6963 ( .A1(n5419), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5420) );
  AND2_X1 U6964 ( .A1(n5447), .A2(n5420), .ZN(n8734) );
  OR2_X1 U6965 ( .A1(n5435), .A2(n8734), .ZN(n5421) );
  NAND4_X1 U6966 ( .A1(n5424), .A2(n5423), .A3(n5422), .A4(n5421), .ZN(n8743)
         );
  NAND2_X1 U6967 ( .A1(n8901), .A2(n7644), .ZN(n8105) );
  NAND2_X1 U6968 ( .A1(n8104), .A2(n8105), .ZN(n8726) );
  NAND2_X1 U6969 ( .A1(n8729), .A2(n8726), .ZN(n5426) );
  NAND2_X1 U6970 ( .A1(n8901), .A2(n8743), .ZN(n5425) );
  NAND2_X1 U6971 ( .A1(n5426), .A2(n5425), .ZN(n8712) );
  XNOR2_X1 U6972 ( .A(n5428), .B(n5427), .ZN(n6864) );
  NAND2_X1 U6973 ( .A1(n6864), .A2(n5176), .ZN(n5434) );
  NAND2_X1 U6974 ( .A1(n5413), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5429) );
  MUX2_X1 U6975 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5429), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n5432) );
  NAND2_X1 U6976 ( .A1(n5432), .A2(n5431), .ZN(n8517) );
  INV_X1 U6977 ( .A(n8517), .ZN(n10214) );
  AOI22_X1 U6978 ( .A1(n5461), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5460), .B2(
        n10214), .ZN(n5433) );
  NAND2_X1 U6979 ( .A1(n5189), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5439) );
  INV_X1 U6980 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n10217) );
  OR2_X1 U6981 ( .A1(n8179), .A2(n10217), .ZN(n5438) );
  INV_X1 U6982 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8717) );
  OR2_X1 U6983 ( .A1(n4393), .A2(n8717), .ZN(n5437) );
  INV_X1 U6984 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n10234) );
  XNOR2_X1 U6985 ( .A(n5447), .B(n10234), .ZN(n8716) );
  OR2_X1 U6986 ( .A1(n5435), .A2(n8716), .ZN(n5436) );
  NAND4_X1 U6987 ( .A1(n5439), .A2(n5438), .A3(n5437), .A4(n5436), .ZN(n8731)
         );
  OR2_X1 U6988 ( .A1(n8818), .A2(n8377), .ZN(n8108) );
  NAND2_X1 U6989 ( .A1(n8818), .A2(n8377), .ZN(n8701) );
  NAND2_X1 U6990 ( .A1(n8108), .A2(n8701), .ZN(n8721) );
  NAND2_X1 U6991 ( .A1(n8712), .A2(n8721), .ZN(n5441) );
  NAND2_X1 U6992 ( .A1(n8818), .A2(n8731), .ZN(n5440) );
  NAND2_X1 U6993 ( .A1(n5441), .A2(n5440), .ZN(n5442) );
  XNOR2_X1 U6994 ( .A(n5444), .B(n5443), .ZN(n6895) );
  NAND2_X1 U6995 ( .A1(n6895), .A2(n5176), .ZN(n5446) );
  NAND2_X1 U6996 ( .A1(n5431), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5457) );
  XNOR2_X1 U6997 ( .A(n5457), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8548) );
  AOI22_X1 U6998 ( .A1(n5461), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5460), .B2(
        n8548), .ZN(n5445) );
  NAND2_X1 U6999 ( .A1(n5575), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5452) );
  INV_X1 U7000 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9796) );
  OR2_X1 U7001 ( .A1(n5234), .A2(n9796), .ZN(n5451) );
  OAI21_X1 U7002 ( .B1(n5447), .B2(P2_REG3_REG_17__SCAN_IN), .A(
        P2_REG3_REG_18__SCAN_IN), .ZN(n5448) );
  AND2_X1 U7003 ( .A1(n5464), .A2(n5448), .ZN(n8373) );
  OR2_X1 U7004 ( .A1(n5435), .A2(n8373), .ZN(n5450) );
  INV_X1 U7005 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8815) );
  OR2_X1 U7006 ( .A1(n8179), .A2(n8815), .ZN(n5449) );
  NAND4_X1 U7007 ( .A1(n5452), .A2(n5451), .A3(n5450), .A4(n5449), .ZN(n8714)
         );
  NAND2_X1 U7008 ( .A1(n8894), .A2(n8692), .ZN(n8109) );
  XNOR2_X1 U7009 ( .A(n5455), .B(n5454), .ZN(n7006) );
  NAND2_X1 U7010 ( .A1(n7006), .A2(n5176), .ZN(n5463) );
  INV_X1 U7011 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5456) );
  NAND2_X1 U7012 ( .A1(n5457), .A2(n5456), .ZN(n5458) );
  NAND2_X1 U7013 ( .A1(n5458), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5459) );
  AOI22_X1 U7014 ( .A1(n5461), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n5618), .B2(
        n5460), .ZN(n5462) );
  NAND2_X1 U7015 ( .A1(n5464), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5465) );
  NAND2_X1 U7016 ( .A1(n5480), .A2(n5465), .ZN(n8698) );
  NAND2_X1 U7017 ( .A1(n5574), .A2(n8698), .ZN(n5469) );
  INV_X1 U7018 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8697) );
  OR2_X1 U7019 ( .A1(n5200), .A2(n8697), .ZN(n5468) );
  INV_X1 U7020 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8888) );
  OR2_X1 U7021 ( .A1(n5234), .A2(n8888), .ZN(n5467) );
  INV_X1 U7022 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9730) );
  OR2_X1 U7023 ( .A1(n8179), .A2(n9730), .ZN(n5466) );
  NAND2_X1 U7024 ( .A1(n8889), .A2(n8357), .ZN(n8117) );
  NAND2_X1 U7025 ( .A1(n8670), .A2(n8117), .ZN(n8231) );
  OR2_X1 U7026 ( .A1(n8894), .A2(n8714), .ZN(n8687) );
  AND2_X1 U7027 ( .A1(n8231), .A2(n8687), .ZN(n5470) );
  NAND2_X1 U7028 ( .A1(n5472), .A2(n5471), .ZN(n5475) );
  AND2_X1 U7029 ( .A1(n5473), .A2(n5486), .ZN(n5474) );
  NAND2_X1 U7030 ( .A1(n7107), .A2(n5176), .ZN(n5477) );
  NAND2_X1 U7031 ( .A1(n5461), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5476) );
  INV_X1 U7032 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8810) );
  OR2_X1 U7033 ( .A1(n8179), .A2(n8810), .ZN(n5479) );
  INV_X1 U7034 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8678) );
  OR2_X1 U7035 ( .A1(n4393), .A2(n8678), .ZN(n5478) );
  AND2_X1 U7036 ( .A1(n5479), .A2(n5478), .ZN(n5484) );
  NAND2_X1 U7037 ( .A1(n5480), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5481) );
  NAND2_X1 U7038 ( .A1(n5492), .A2(n5481), .ZN(n8679) );
  NAND2_X1 U7039 ( .A1(n8679), .A2(n5574), .ZN(n5483) );
  NAND2_X1 U7040 ( .A1(n5189), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5482) );
  NAND2_X1 U7041 ( .A1(n8883), .A2(n8693), .ZN(n8118) );
  NAND2_X1 U7042 ( .A1(n8119), .A2(n8118), .ZN(n8674) );
  NAND2_X1 U7043 ( .A1(n8889), .A2(n8706), .ZN(n8673) );
  AND2_X1 U7044 ( .A1(n8674), .A2(n8673), .ZN(n5485) );
  INV_X1 U7045 ( .A(n8693), .ZN(n8663) );
  OR2_X1 U7046 ( .A1(n8883), .A2(n8663), .ZN(n8660) );
  NAND2_X1 U7047 ( .A1(n8659), .A2(n8660), .ZN(n5496) );
  AND2_X1 U7048 ( .A1(n5487), .A2(n5486), .ZN(n5489) );
  NAND2_X1 U7049 ( .A1(n7189), .A2(n5176), .ZN(n5491) );
  NAND2_X1 U7050 ( .A1(n5461), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5490) );
  INV_X1 U7051 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8876) );
  NAND2_X1 U7052 ( .A1(n5492), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5493) );
  NAND2_X1 U7053 ( .A1(n5501), .A2(n5493), .ZN(n8667) );
  NAND2_X1 U7054 ( .A1(n8667), .A2(n5574), .ZN(n5495) );
  AOI22_X1 U7055 ( .A1(n5537), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n5575), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n5494) );
  INV_X1 U7056 ( .A(n8676), .ZN(n6257) );
  NAND2_X1 U7057 ( .A1(n8877), .A2(n6257), .ZN(n8123) );
  NAND2_X1 U7058 ( .A1(n8120), .A2(n8123), .ZN(n8657) );
  OR2_X1 U7059 ( .A1(n8877), .A2(n8676), .ZN(n8647) );
  NAND2_X1 U7060 ( .A1(n8646), .A2(n8647), .ZN(n5505) );
  XNOR2_X1 U7061 ( .A(n5498), .B(n5497), .ZN(n7301) );
  NAND2_X1 U7062 ( .A1(n7301), .A2(n5176), .ZN(n5500) );
  NAND2_X1 U7063 ( .A1(n5461), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5499) );
  INV_X1 U7064 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8870) );
  NAND2_X1 U7065 ( .A1(n5501), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5502) );
  NAND2_X1 U7066 ( .A1(n5511), .A2(n5502), .ZN(n8654) );
  NAND2_X1 U7067 ( .A1(n8654), .A2(n5574), .ZN(n5504) );
  AOI22_X1 U7068 ( .A1(n5537), .A2(P2_REG1_REG_22__SCAN_IN), .B1(n5575), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n5503) );
  INV_X1 U7069 ( .A(n8664), .ZN(n8264) );
  NAND2_X1 U7070 ( .A1(n8871), .A2(n8264), .ZN(n8128) );
  NAND2_X1 U7071 ( .A1(n8129), .A2(n8128), .ZN(n8127) );
  NAND2_X1 U7072 ( .A1(n5505), .A2(n8127), .ZN(n8650) );
  OR2_X1 U7073 ( .A1(n8871), .A2(n8664), .ZN(n5506) );
  NAND2_X1 U7074 ( .A1(n8650), .A2(n5506), .ZN(n8639) );
  NAND2_X1 U7075 ( .A1(n7310), .A2(n5176), .ZN(n5510) );
  NAND2_X1 U7076 ( .A1(n5461), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5509) );
  INV_X1 U7077 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8864) );
  NAND2_X1 U7078 ( .A1(n5511), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5512) );
  NAND2_X1 U7079 ( .A1(n5522), .A2(n5512), .ZN(n8642) );
  NAND2_X1 U7080 ( .A1(n8642), .A2(n5574), .ZN(n5514) );
  AOI22_X1 U7081 ( .A1(n5537), .A2(P2_REG1_REG_23__SCAN_IN), .B1(n5575), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n5513) );
  NAND2_X1 U7082 ( .A1(n8865), .A2(n8651), .ZN(n5515) );
  NAND2_X1 U7083 ( .A1(n8639), .A2(n5515), .ZN(n5517) );
  OR2_X1 U7084 ( .A1(n8865), .A2(n8651), .ZN(n5516) );
  NAND2_X1 U7085 ( .A1(n5517), .A2(n5516), .ZN(n8626) );
  XNOR2_X1 U7086 ( .A(n5519), .B(n5518), .ZN(n7378) );
  NAND2_X1 U7087 ( .A1(n7378), .A2(n5176), .ZN(n5521) );
  NAND2_X1 U7088 ( .A1(n5461), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5520) );
  NAND2_X1 U7089 ( .A1(n5522), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5523) );
  NAND2_X1 U7090 ( .A1(n5535), .A2(n5523), .ZN(n8634) );
  NAND2_X1 U7091 ( .A1(n8634), .A2(n5574), .ZN(n5528) );
  INV_X1 U7092 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8858) );
  NAND2_X1 U7093 ( .A1(n5575), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5525) );
  NAND2_X1 U7094 ( .A1(n5537), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5524) );
  OAI211_X1 U7095 ( .C1(n8858), .C2(n5234), .A(n5525), .B(n5524), .ZN(n5526)
         );
  INV_X1 U7096 ( .A(n5526), .ZN(n5527) );
  NOR2_X1 U7097 ( .A1(n8859), .A2(n8640), .ZN(n5530) );
  NAND2_X1 U7098 ( .A1(n8859), .A2(n8640), .ZN(n5529) );
  OAI21_X2 U7099 ( .B1(n8626), .B2(n5530), .A(n5529), .ZN(n8612) );
  XNOR2_X1 U7100 ( .A(n5532), .B(n5531), .ZN(n7407) );
  NAND2_X1 U7101 ( .A1(n7407), .A2(n5176), .ZN(n5534) );
  NAND2_X1 U7102 ( .A1(n5461), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5533) );
  NAND2_X1 U7103 ( .A1(n5535), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5536) );
  NAND2_X1 U7104 ( .A1(n5547), .A2(n5536), .ZN(n8616) );
  NAND2_X1 U7105 ( .A1(n8616), .A2(n5574), .ZN(n5542) );
  INV_X1 U7106 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8852) );
  NAND2_X1 U7107 ( .A1(n5575), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5539) );
  NAND2_X1 U7108 ( .A1(n5537), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5538) );
  OAI211_X1 U7109 ( .C1(n8852), .C2(n5234), .A(n5539), .B(n5538), .ZN(n5540)
         );
  INV_X1 U7110 ( .A(n5540), .ZN(n5541) );
  AND2_X1 U7111 ( .A1(n8853), .A2(n8401), .ZN(n8601) );
  NAND2_X1 U7112 ( .A1(n7500), .A2(n5176), .ZN(n5546) );
  NAND2_X1 U7113 ( .A1(n5461), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5545) );
  NAND2_X1 U7114 ( .A1(n5547), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5548) );
  NAND2_X1 U7115 ( .A1(n5549), .A2(n5548), .ZN(n8609) );
  NAND2_X1 U7116 ( .A1(n8609), .A2(n5574), .ZN(n5554) );
  INV_X1 U7117 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8845) );
  NAND2_X1 U7118 ( .A1(n5537), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5551) );
  NAND2_X1 U7119 ( .A1(n5575), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5550) );
  OAI211_X1 U7120 ( .C1(n8845), .C2(n5234), .A(n5551), .B(n5550), .ZN(n5552)
         );
  INV_X1 U7121 ( .A(n5552), .ZN(n5553) );
  AND2_X1 U7122 ( .A1(n8846), .A2(n8587), .ZN(n5558) );
  OR2_X1 U7123 ( .A1(n8601), .A2(n5558), .ZN(n5555) );
  NOR2_X1 U7124 ( .A1(n8612), .A2(n5555), .ZN(n5560) );
  OR2_X1 U7125 ( .A1(n8846), .A2(n8587), .ZN(n5556) );
  OR2_X1 U7126 ( .A1(n8853), .A2(n8401), .ZN(n8602) );
  AND2_X1 U7127 ( .A1(n5556), .A2(n8602), .ZN(n5557) );
  NOR2_X1 U7128 ( .A1(n5558), .A2(n5557), .ZN(n5559) );
  INV_X1 U7129 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5564) );
  INV_X1 U7130 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7637) );
  MUX2_X1 U7131 ( .A(n5564), .B(n7637), .S(n5779), .Z(n5566) );
  INV_X1 U7132 ( .A(SI_28_), .ZN(n5565) );
  NAND2_X1 U7133 ( .A1(n5566), .A2(n5565), .ZN(n5677) );
  INV_X1 U7134 ( .A(n5566), .ZN(n5567) );
  NAND2_X1 U7135 ( .A1(n5567), .A2(SI_28_), .ZN(n5568) );
  NAND2_X1 U7136 ( .A1(n7603), .A2(n5176), .ZN(n5570) );
  NAND2_X1 U7137 ( .A1(n5461), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5569) );
  NAND2_X1 U7138 ( .A1(n5571), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5572) );
  NAND2_X1 U7139 ( .A1(n5573), .A2(n5572), .ZN(n8283) );
  NAND2_X1 U7140 ( .A1(n8283), .A2(n5574), .ZN(n5580) );
  NAND2_X1 U7141 ( .A1(n5537), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5577) );
  NAND2_X1 U7142 ( .A1(n5575), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5576) );
  OAI211_X1 U7143 ( .C1(n5623), .C2(n5234), .A(n5577), .B(n5576), .ZN(n5578)
         );
  INV_X1 U7144 ( .A(n5578), .ZN(n5579) );
  XNOR2_X1 U7145 ( .A(n5681), .B(n5673), .ZN(n5584) );
  NAND2_X1 U7146 ( .A1(n8029), .A2(n5618), .ZN(n5616) );
  NAND2_X1 U7147 ( .A1(n5581), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5582) );
  OR2_X1 U7148 ( .A1(n8241), .A2(n8203), .ZN(n5583) );
  OAI222_X1 U7149 ( .A1(n8761), .A2(n8607), .B1(n8762), .B2(n8286), .C1(n5584), 
        .C2(n8629), .ZN(n8781) );
  INV_X1 U7150 ( .A(n8781), .ZN(n5665) );
  NAND2_X1 U7151 ( .A1(n5593), .A2(n5585), .ZN(n5587) );
  NAND2_X1 U7152 ( .A1(n5586), .A2(n5587), .ZN(n5598) );
  XNOR2_X1 U7153 ( .A(n5598), .B(P2_B_REG_SCAN_IN), .ZN(n5590) );
  NAND2_X1 U7154 ( .A1(n5590), .A2(n5600), .ZN(n5596) );
  NAND2_X1 U7155 ( .A1(n5593), .A2(n5592), .ZN(n5594) );
  NAND2_X1 U7156 ( .A1(n5594), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n5595) );
  NAND2_X1 U7157 ( .A1(n5596), .A2(n5597), .ZN(n5599) );
  NAND2_X1 U7158 ( .A1(n7524), .A2(n5598), .ZN(n6397) );
  INV_X1 U7159 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6353) );
  NAND2_X1 U7160 ( .A1(n6364), .A2(n6353), .ZN(n5602) );
  NAND2_X1 U7161 ( .A1(n5600), .A2(n7524), .ZN(n5601) );
  NAND2_X1 U7162 ( .A1(n6178), .A2(n6349), .ZN(n5655) );
  NOR2_X1 U7163 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .ZN(
        n9700) );
  NOR4_X1 U7164 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n5605) );
  NOR4_X1 U7165 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_27__SCAN_IN), .ZN(n5604) );
  NOR4_X1 U7166 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_30__SCAN_IN), .ZN(n5603) );
  AND4_X1 U7167 ( .A1(n9700), .A2(n5605), .A3(n5604), .A4(n5603), .ZN(n5611)
         );
  NOR4_X1 U7168 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n5609) );
  NOR4_X1 U7169 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n5608) );
  NOR4_X1 U7170 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5607) );
  NOR4_X1 U7171 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n5606) );
  AND4_X1 U7172 ( .A1(n5609), .A2(n5608), .A3(n5607), .A4(n5606), .ZN(n5610)
         );
  NAND2_X1 U7173 ( .A1(n5611), .A2(n5610), .ZN(n5612) );
  NOR2_X1 U7174 ( .A1(n7524), .A2(n5598), .ZN(n5614) );
  INV_X1 U7175 ( .A(n5600), .ZN(n5613) );
  NAND2_X1 U7176 ( .A1(n4482), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5615) );
  XNOR2_X1 U7177 ( .A(n5615), .B(n4992), .ZN(n6318) );
  INV_X1 U7178 ( .A(n6285), .ZN(n6276) );
  AND2_X1 U7179 ( .A1(n8186), .A2(n10274), .ZN(n5617) );
  NAND2_X1 U7180 ( .A1(n8241), .A2(n8254), .ZN(n6179) );
  OR2_X1 U7181 ( .A1(n5616), .A2(n6179), .ZN(n6275) );
  NAND2_X1 U7182 ( .A1(n5617), .A2(n6275), .ZN(n6277) );
  NAND2_X1 U7183 ( .A1(n6277), .A2(n8632), .ZN(n6289) );
  NAND2_X1 U7184 ( .A1(n6276), .A2(n6289), .ZN(n5622) );
  OR2_X1 U7185 ( .A1(n6349), .A2(n6178), .ZN(n6309) );
  INV_X1 U7186 ( .A(n6290), .ZN(n5619) );
  INV_X1 U7187 ( .A(n8028), .ZN(n6352) );
  NAND2_X1 U7188 ( .A1(n5619), .A2(n6352), .ZN(n6282) );
  NAND2_X1 U7189 ( .A1(n8555), .A2(n8203), .ZN(n6182) );
  AND2_X1 U7190 ( .A1(n8027), .A2(n6275), .ZN(n5620) );
  OR2_X1 U7191 ( .A1(n6282), .A2(n5620), .ZN(n5621) );
  MUX2_X1 U7192 ( .A(n5623), .B(n5665), .S(n10286), .Z(n5650) );
  NAND2_X1 U7193 ( .A1(n6844), .A2(n6684), .ZN(n8035) );
  INV_X1 U7194 ( .A(n8035), .ZN(n5624) );
  NAND2_X1 U7195 ( .A1(n6840), .A2(n8042), .ZN(n8754) );
  INV_X1 U7196 ( .A(n5625), .ZN(n8757) );
  NAND2_X1 U7197 ( .A1(n8754), .A2(n8757), .ZN(n8753) );
  NAND2_X1 U7198 ( .A1(n8753), .A2(n6853), .ZN(n5626) );
  OR2_X1 U7199 ( .A1(n8763), .A2(n6861), .ZN(n8051) );
  NAND2_X1 U7200 ( .A1(n8763), .A2(n6861), .ZN(n8039) );
  NAND2_X1 U7201 ( .A1(n5626), .A2(n8211), .ZN(n6854) );
  NAND2_X1 U7202 ( .A1(n6854), .A2(n8039), .ZN(n5627) );
  INV_X1 U7203 ( .A(n6818), .ZN(n8213) );
  NAND2_X1 U7204 ( .A1(n5627), .A2(n8213), .ZN(n6820) );
  NAND2_X1 U7205 ( .A1(n6820), .A2(n8052), .ZN(n6898) );
  INV_X1 U7206 ( .A(n8410), .ZN(n6823) );
  NAND2_X1 U7207 ( .A1(n6823), .A2(n6902), .ZN(n8071) );
  INV_X1 U7208 ( .A(n6902), .ZN(n6934) );
  NAND2_X1 U7209 ( .A1(n6934), .A2(n8410), .ZN(n8068) );
  NAND2_X1 U7210 ( .A1(n6898), .A2(n8214), .ZN(n6897) );
  NAND2_X1 U7211 ( .A1(n6897), .A2(n8071), .ZN(n6957) );
  NAND2_X1 U7212 ( .A1(n6957), .A2(n6956), .ZN(n5628) );
  NAND2_X1 U7213 ( .A1(n5628), .A2(n8072), .ZN(n7191) );
  INV_X1 U7214 ( .A(n8220), .ZN(n8056) );
  INV_X1 U7215 ( .A(n8059), .ZN(n5629) );
  OR2_X1 U7216 ( .A1(n10272), .A2(n7701), .ZN(n8083) );
  NAND2_X1 U7217 ( .A1(n10272), .A2(n7701), .ZN(n8080) );
  NAND2_X1 U7218 ( .A1(n8083), .A2(n8080), .ZN(n8223) );
  INV_X1 U7219 ( .A(n8223), .ZN(n5630) );
  NAND2_X1 U7220 ( .A1(n7472), .A2(n8080), .ZN(n5632) );
  XNOR2_X1 U7221 ( .A(n7401), .B(n8303), .ZN(n8086) );
  NAND2_X1 U7222 ( .A1(n5632), .A2(n7394), .ZN(n7400) );
  NAND2_X1 U7223 ( .A1(n7401), .A2(n8303), .ZN(n8032) );
  INV_X1 U7224 ( .A(n8403), .ZN(n7708) );
  NAND2_X1 U7225 ( .A1(n10282), .A2(n7708), .ZN(n8033) );
  NAND2_X1 U7226 ( .A1(n8030), .A2(n8033), .ZN(n8087) );
  NOR2_X1 U7227 ( .A1(n7713), .A2(n8308), .ZN(n8092) );
  NAND2_X1 U7228 ( .A1(n7713), .A2(n8308), .ZN(n8090) );
  NAND2_X1 U7229 ( .A1(n7721), .A2(n8097), .ZN(n5634) );
  NAND2_X1 U7230 ( .A1(n7736), .A2(n7507), .ZN(n8096) );
  NAND2_X1 U7231 ( .A1(n5634), .A2(n8096), .ZN(n8738) );
  OR2_X1 U7232 ( .A1(n8907), .A2(n7570), .ZN(n8100) );
  NAND2_X1 U7233 ( .A1(n8738), .A2(n8100), .ZN(n5635) );
  NAND2_X1 U7234 ( .A1(n8907), .A2(n7570), .ZN(n8099) );
  NAND2_X1 U7235 ( .A1(n5635), .A2(n8099), .ZN(n8727) );
  INV_X1 U7236 ( .A(n8105), .ZN(n5636) );
  NOR2_X1 U7237 ( .A1(n8231), .A2(n8683), .ZN(n5639) );
  OR2_X1 U7238 ( .A1(n8721), .A2(n5639), .ZN(n5637) );
  AND2_X1 U7239 ( .A1(n8109), .A2(n8701), .ZN(n8682) );
  INV_X1 U7240 ( .A(n8231), .ZN(n8688) );
  AND2_X1 U7241 ( .A1(n8682), .A2(n8688), .ZN(n5638) );
  OR2_X1 U7242 ( .A1(n5639), .A2(n5638), .ZN(n5640) );
  AND2_X1 U7243 ( .A1(n8119), .A2(n8670), .ZN(n5641) );
  NAND2_X1 U7244 ( .A1(n8685), .A2(n5641), .ZN(n5642) );
  INV_X1 U7245 ( .A(n8123), .ZN(n5643) );
  NOR2_X1 U7246 ( .A1(n8865), .A2(n8630), .ZN(n8135) );
  NAND2_X1 U7247 ( .A1(n8859), .A2(n8614), .ZN(n8207) );
  NAND2_X1 U7248 ( .A1(n8865), .A2(n8630), .ZN(n8623) );
  AND2_X1 U7249 ( .A1(n8207), .A2(n8623), .ZN(n8133) );
  NAND2_X1 U7250 ( .A1(n8624), .A2(n8133), .ZN(n5644) );
  NAND2_X1 U7251 ( .A1(n8853), .A2(n8631), .ZN(n8144) );
  NOR2_X1 U7252 ( .A1(n8853), .A2(n8631), .ZN(n8142) );
  AOI21_X2 U7253 ( .B1(n8617), .B2(n8144), .A(n8142), .ZN(n8600) );
  XNOR2_X1 U7254 ( .A(n6284), .B(n8400), .ZN(n8584) );
  NOR2_X1 U7255 ( .A1(n6284), .A2(n8607), .ZN(n8152) );
  XNOR2_X1 U7256 ( .A(n5674), .B(n5673), .ZN(n8783) );
  NAND2_X1 U7257 ( .A1(n8204), .A2(n8203), .ZN(n6183) );
  INV_X1 U7258 ( .A(n6183), .ZN(n5645) );
  OR2_X1 U7259 ( .A1(n5645), .A2(n8029), .ZN(n5646) );
  AND2_X1 U7260 ( .A1(n5646), .A2(n8555), .ZN(n5657) );
  NAND2_X1 U7261 ( .A1(n5657), .A2(n8027), .ZN(n7479) );
  INV_X1 U7262 ( .A(n10279), .ZN(n10247) );
  NAND2_X1 U7263 ( .A1(n8288), .A2(n5698), .ZN(n5648) );
  INV_X1 U7264 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n5666) );
  INV_X1 U7265 ( .A(n6182), .ZN(n5651) );
  OR2_X1 U7266 ( .A1(n8186), .A2(n5651), .ZN(n6293) );
  INV_X1 U7267 ( .A(n6293), .ZN(n5652) );
  OR2_X1 U7268 ( .A1(n8028), .A2(n5652), .ZN(n5654) );
  OR2_X1 U7269 ( .A1(n5654), .A2(n5653), .ZN(n6308) );
  INV_X1 U7270 ( .A(n6308), .ZN(n5656) );
  AND2_X1 U7271 ( .A1(n5656), .A2(n5655), .ZN(n5664) );
  NAND2_X1 U7272 ( .A1(n5657), .A2(n8254), .ZN(n5658) );
  AND2_X1 U7273 ( .A1(n5658), .A2(n8186), .ZN(n5659) );
  OR2_X1 U7274 ( .A1(n6349), .A2(n5659), .ZN(n5662) );
  INV_X1 U7275 ( .A(n5659), .ZN(n5660) );
  OR2_X1 U7276 ( .A1(n6178), .A2(n5660), .ZN(n5661) );
  NAND2_X1 U7277 ( .A1(n5662), .A2(n5661), .ZN(n6310) );
  INV_X1 U7278 ( .A(n6310), .ZN(n5663) );
  NAND2_X1 U7279 ( .A1(n5664), .A2(n5663), .ZN(n5668) );
  OR2_X1 U7280 ( .A1(n10268), .A2(n8204), .ZN(n6306) );
  MUX2_X1 U7281 ( .A(n5666), .B(n5665), .S(n8745), .Z(n5672) );
  OR2_X1 U7282 ( .A1(n6183), .A2(n8555), .ZN(n6842) );
  AND2_X1 U7283 ( .A1(n7479), .A2(n6842), .ZN(n5667) );
  INV_X1 U7284 ( .A(n5668), .ZN(n5669) );
  INV_X1 U7285 ( .A(n8632), .ZN(n8769) );
  AOI22_X1 U7286 ( .A1(n8288), .A2(n8749), .B1(n8748), .B2(n8283), .ZN(n5670)
         );
  NAND2_X1 U7287 ( .A1(n5676), .A2(n5675), .ZN(n5678) );
  INV_X1 U7288 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7746) );
  INV_X1 U7289 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9967) );
  MUX2_X1 U7290 ( .A(n7746), .B(n9967), .S(n6325), .Z(n7741) );
  NAND2_X1 U7291 ( .A1(n7747), .A2(n5176), .ZN(n5680) );
  NAND2_X1 U7292 ( .A1(n5461), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n5679) );
  XNOR2_X1 U7293 ( .A(n8184), .B(n8286), .ZN(n5684) );
  INV_X1 U7294 ( .A(n8288), .ZN(n8782) );
  OAI22_X2 U7295 ( .A1(n5683), .A2(n5682), .B1(n8156), .B2(n8782), .ZN(n5685)
         );
  XNOR2_X1 U7296 ( .A(n5685), .B(n5684), .ZN(n5695) );
  INV_X1 U7297 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9895) );
  NAND2_X1 U7298 ( .A1(n5189), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5688) );
  INV_X1 U7299 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n5686) );
  OR2_X1 U7300 ( .A1(n5200), .A2(n5686), .ZN(n5687) );
  OAI211_X1 U7301 ( .C1(n8179), .C2(n9895), .A(n5688), .B(n5687), .ZN(n5689)
         );
  INV_X1 U7302 ( .A(n5689), .ZN(n5690) );
  NAND2_X1 U7303 ( .A1(n5184), .A2(P2_B_REG_SCAN_IN), .ZN(n5691) );
  NAND2_X1 U7304 ( .A1(n5047), .A2(n5691), .ZN(n8569) );
  OAI21_X1 U7305 ( .B1(n5695), .B2(n8629), .A(n5694), .ZN(n8577) );
  INV_X1 U7306 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n5696) );
  NOR2_X1 U7307 ( .A1(n10286), .A2(n5696), .ZN(n5697) );
  NAND3_X1 U7308 ( .A1(n5900), .A2(n5702), .A3(n5701), .ZN(n5946) );
  NAND3_X1 U7309 ( .A1(n5705), .A2(n5704), .A3(n5703), .ZN(n5706) );
  NAND2_X1 U7310 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .ZN(n5710) );
  NAND2_X1 U7311 ( .A1(n6140), .A2(n5710), .ZN(n5711) );
  XNOR2_X2 U7312 ( .A(n5711), .B(P1_IR_REG_27__SCAN_IN), .ZN(n6372) );
  NAND2_X2 U7313 ( .A1(n6372), .A2(n6130), .ZN(n5770) );
  NAND2_X1 U7314 ( .A1(n7006), .A2(n7818), .ZN(n5722) );
  NAND2_X1 U7315 ( .A1(n5984), .A2(n5716), .ZN(n5717) );
  NAND2_X1 U7316 ( .A1(n5717), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5752) );
  NAND2_X1 U7317 ( .A1(n5752), .A2(n5718), .ZN(n5719) );
  AOI22_X1 U7318 ( .A1(n5986), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n8005), .B2(
        n5985), .ZN(n5721) );
  INV_X1 U7319 ( .A(n9625), .ZN(n9518) );
  NAND2_X1 U7320 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n5723) );
  INV_X1 U7321 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5733) );
  NAND2_X1 U7322 ( .A1(n5728), .A2(n5733), .ZN(n5729) );
  XNOR2_X2 U7323 ( .A(n5734), .B(n5733), .ZN(n5747) );
  INV_X1 U7324 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9520) );
  OR2_X1 U7325 ( .A1(n4979), .A2(n9520), .ZN(n5751) );
  NAND2_X1 U7326 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5829) );
  INV_X1 U7327 ( .A(n5829), .ZN(n5736) );
  NAND2_X1 U7328 ( .A1(n5736), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5841) );
  INV_X1 U7329 ( .A(n5841), .ZN(n5737) );
  NAND2_X1 U7330 ( .A1(n5737), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5855) );
  INV_X1 U7331 ( .A(n5855), .ZN(n5738) );
  NAND2_X1 U7332 ( .A1(n5738), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5868) );
  INV_X1 U7333 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9286) );
  AND2_X1 U7334 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_17__SCAN_IN), 
        .ZN(n5743) );
  INV_X1 U7335 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9763) );
  NAND2_X1 U7336 ( .A1(n5758), .A2(n9763), .ZN(n5745) );
  NAND2_X1 U7337 ( .A1(n6002), .A2(n5745), .ZN(n9519) );
  OR2_X1 U7338 ( .A1(n6131), .A2(n9519), .ZN(n5750) );
  INV_X1 U7339 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n5746) );
  OR2_X1 U7340 ( .A1(n6072), .A2(n5746), .ZN(n5749) );
  INV_X1 U7341 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9333) );
  OR2_X1 U7342 ( .A1(n5790), .A2(n9333), .ZN(n5748) );
  NAND2_X1 U7343 ( .A1(n6895), .A2(n7818), .ZN(n5754) );
  XNOR2_X1 U7344 ( .A(n5752), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9330) );
  AOI22_X1 U7345 ( .A1(n5986), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5985), .B2(
        n9330), .ZN(n5753) );
  INV_X1 U7346 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9527) );
  INV_X1 U7347 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9949) );
  OR2_X1 U7348 ( .A1(n6072), .A2(n9949), .ZN(n5755) );
  OAI21_X1 U7349 ( .B1(n4979), .B2(n9527), .A(n5755), .ZN(n5761) );
  INV_X1 U7350 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5990) );
  INV_X1 U7351 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5756) );
  OAI21_X1 U7352 ( .B1(n5991), .B2(n5990), .A(n5756), .ZN(n5757) );
  NAND2_X1 U7353 ( .A1(n5758), .A2(n5757), .ZN(n9526) );
  INV_X1 U7354 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9633) );
  OR2_X1 U7355 ( .A1(n5790), .A2(n9633), .ZN(n5759) );
  OAI21_X1 U7356 ( .B1(n6131), .B2(n9526), .A(n5759), .ZN(n5760) );
  INV_X1 U7357 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6645) );
  OR2_X1 U7358 ( .A1(n6131), .A2(n6645), .ZN(n5767) );
  INV_X1 U7359 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5762) );
  OR2_X1 U7360 ( .A1(n5800), .A2(n5762), .ZN(n5766) );
  INV_X1 U7361 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10175) );
  OR2_X1 U7362 ( .A1(n5790), .A2(n10175), .ZN(n5765) );
  INV_X1 U7363 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5769) );
  OR2_X1 U7364 ( .A1(n5770), .A2(n6381), .ZN(n5771) );
  OAI211_X1 U7365 ( .C1(n5863), .C2(n6332), .A(n5772), .B(n5771), .ZN(n5773)
         );
  INV_X1 U7366 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7015) );
  INV_X1 U7367 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6629) );
  INV_X1 U7368 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6616) );
  OR2_X1 U7369 ( .A1(n5790), .A2(n6616), .ZN(n5776) );
  INV_X1 U7370 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5774) );
  NAND4_X2 U7371 ( .A1(n5778), .A2(n5777), .A3(n5776), .A4(n5775), .ZN(n6109)
         );
  NAND2_X1 U7372 ( .A1(n6325), .A2(SI_0_), .ZN(n5781) );
  INV_X1 U7373 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5780) );
  NAND2_X1 U7374 ( .A1(n5781), .A2(n5780), .ZN(n5783) );
  AND2_X1 U7375 ( .A1(n5783), .A2(n5782), .ZN(n9970) );
  MUX2_X1 U7376 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9970), .S(n6361), .Z(n6626) );
  NAND2_X1 U7377 ( .A1(n6109), .A2(n6626), .ZN(n10085) );
  NAND2_X1 U7378 ( .A1(n6108), .A2(n10085), .ZN(n5786) );
  INV_X1 U7379 ( .A(n5784), .ZN(n6702) );
  NAND2_X1 U7380 ( .A1(n6702), .A2(n6106), .ZN(n5785) );
  NAND2_X1 U7381 ( .A1(n5786), .A2(n5785), .ZN(n10075) );
  OR2_X1 U7382 ( .A1(n5787), .A2(n4808), .ZN(n5820) );
  XNOR2_X1 U7383 ( .A(n5820), .B(n4705), .ZN(n9255) );
  OR2_X1 U7384 ( .A1(n5863), .A2(n6326), .ZN(n5788) );
  OAI211_X1 U7385 ( .C1(n6361), .C2(n9255), .A(n4971), .B(n5788), .ZN(n5795)
         );
  INV_X1 U7386 ( .A(n5795), .ZN(n5796) );
  INV_X1 U7387 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6705) );
  INV_X1 U7388 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5789) );
  INV_X1 U7389 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6380) );
  OR2_X1 U7390 ( .A1(n5790), .A2(n6380), .ZN(n5793) );
  INV_X1 U7391 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5791) );
  OR2_X1 U7392 ( .A1(n5800), .A2(n5791), .ZN(n5792) );
  INV_X1 U7393 ( .A(n6693), .ZN(n6805) );
  NAND2_X1 U7394 ( .A1(n5796), .A2(n6805), .ZN(n6112) );
  NAND2_X1 U7395 ( .A1(n6693), .A2(n5795), .ZN(n6111) );
  NAND2_X1 U7396 ( .A1(n10075), .A2(n10076), .ZN(n5798) );
  NAND2_X1 U7397 ( .A1(n6693), .A2(n5796), .ZN(n5797) );
  NAND2_X1 U7398 ( .A1(n5798), .A2(n5797), .ZN(n7020) );
  INV_X1 U7399 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7024) );
  OR2_X1 U7400 ( .A1(n4979), .A2(n7024), .ZN(n5804) );
  OR2_X1 U7401 ( .A1(n6131), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5803) );
  INV_X1 U7402 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5799) );
  OR2_X1 U7403 ( .A1(n5800), .A2(n5799), .ZN(n5802) );
  INV_X1 U7404 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6376) );
  OR2_X1 U7405 ( .A1(n5790), .A2(n6376), .ZN(n5801) );
  NAND2_X1 U7406 ( .A1(n5820), .A2(n4705), .ZN(n5805) );
  NAND2_X1 U7407 ( .A1(n5805), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5807) );
  INV_X1 U7408 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5806) );
  XNOR2_X1 U7409 ( .A(n5807), .B(n5806), .ZN(n6399) );
  OR2_X1 U7410 ( .A1(n5768), .A2(n6342), .ZN(n5809) );
  OR2_X1 U7411 ( .A1(n5863), .A2(n6341), .ZN(n5808) );
  OAI211_X1 U7412 ( .C1(n6361), .C2(n6399), .A(n5809), .B(n5808), .ZN(n7027)
         );
  NAND2_X1 U7413 ( .A1(n6781), .A2(n7027), .ZN(n7830) );
  INV_X1 U7414 ( .A(n6781), .ZN(n9229) );
  NAND2_X1 U7415 ( .A1(n7830), .A2(n7829), .ZN(n7021) );
  NAND2_X1 U7416 ( .A1(n6781), .A2(n5810), .ZN(n5811) );
  INV_X1 U7417 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7134) );
  INV_X1 U7418 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5812) );
  OR2_X1 U7419 ( .A1(n5790), .A2(n5812), .ZN(n5813) );
  OAI21_X1 U7420 ( .B1(n4979), .B2(n7134), .A(n5813), .ZN(n5817) );
  OAI21_X1 U7421 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n5829), .ZN(n7133) );
  INV_X1 U7422 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5814) );
  OR2_X1 U7423 ( .A1(n5800), .A2(n5814), .ZN(n5815) );
  OAI21_X1 U7424 ( .B1(n6131), .B2(n7133), .A(n5815), .ZN(n5816) );
  OR2_X1 U7425 ( .A1(n5818), .A2(n4808), .ZN(n5819) );
  AND2_X1 U7426 ( .A1(n5820), .A2(n5819), .ZN(n5823) );
  INV_X1 U7427 ( .A(n5823), .ZN(n5821) );
  NAND2_X1 U7428 ( .A1(n5821), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5824) );
  INV_X1 U7429 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5822) );
  NAND2_X1 U7430 ( .A1(n5823), .A2(n5822), .ZN(n5836) );
  INV_X1 U7431 ( .A(n10051), .ZN(n6337) );
  OR2_X1 U7432 ( .A1(n5863), .A2(n6338), .ZN(n5826) );
  OR2_X1 U7433 ( .A1(n7820), .A2(n6339), .ZN(n5825) );
  OAI211_X1 U7434 ( .C1(n6361), .C2(n6337), .A(n5826), .B(n5825), .ZN(n7136)
         );
  NAND2_X1 U7435 ( .A1(n9228), .A2(n7136), .ZN(n5827) );
  INV_X1 U7436 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n5828) );
  OR2_X1 U7437 ( .A1(n4979), .A2(n5828), .ZN(n5835) );
  INV_X1 U7438 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6411) );
  NAND2_X1 U7439 ( .A1(n5829), .A2(n6411), .ZN(n5830) );
  NAND2_X1 U7440 ( .A1(n5841), .A2(n5830), .ZN(n6950) );
  OR2_X1 U7441 ( .A1(n6131), .A2(n6950), .ZN(n5834) );
  INV_X1 U7442 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5831) );
  OR2_X1 U7443 ( .A1(n6072), .A2(n5831), .ZN(n5833) );
  INV_X1 U7444 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6408) );
  OR2_X1 U7445 ( .A1(n5790), .A2(n6408), .ZN(n5832) );
  NAND2_X1 U7446 ( .A1(n5836), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5837) );
  XNOR2_X1 U7447 ( .A(n5837), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6423) );
  INV_X1 U7448 ( .A(n6423), .ZN(n6415) );
  OR2_X1 U7449 ( .A1(n5863), .A2(n6340), .ZN(n5839) );
  OR2_X1 U7450 ( .A1(n5768), .A2(n9808), .ZN(n5838) );
  OAI211_X1 U7451 ( .C1(n6361), .C2(n6415), .A(n5839), .B(n5838), .ZN(n6986)
         );
  NAND2_X1 U7452 ( .A1(n6947), .A2(n6986), .ZN(n7838) );
  INV_X1 U7453 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6999) );
  OR2_X1 U7454 ( .A1(n4979), .A2(n6999), .ZN(n5847) );
  INV_X1 U7455 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5840) );
  NAND2_X1 U7456 ( .A1(n5841), .A2(n5840), .ZN(n5842) );
  NAND2_X1 U7457 ( .A1(n5855), .A2(n5842), .ZN(n7101) );
  OR2_X1 U7458 ( .A1(n6131), .A2(n7101), .ZN(n5846) );
  INV_X1 U7459 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6422) );
  OR2_X1 U7460 ( .A1(n5790), .A2(n6422), .ZN(n5845) );
  INV_X1 U7461 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5843) );
  OR2_X1 U7462 ( .A1(n6072), .A2(n5843), .ZN(n5844) );
  NAND2_X1 U7463 ( .A1(n5848), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5849) );
  MUX2_X1 U7464 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5849), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n5851) );
  AND2_X1 U7465 ( .A1(n5850), .A2(n5851), .ZN(n6464) );
  INV_X1 U7466 ( .A(n6464), .ZN(n6334) );
  OR2_X1 U7467 ( .A1(n5863), .A2(n6335), .ZN(n5853) );
  OR2_X1 U7468 ( .A1(n7820), .A2(n6336), .ZN(n5852) );
  OAI211_X1 U7469 ( .C1(n6361), .C2(n6334), .A(n5853), .B(n5852), .ZN(n6969)
         );
  NAND2_X1 U7470 ( .A1(n7092), .A2(n6969), .ZN(n7848) );
  INV_X1 U7471 ( .A(n7092), .ZN(n9226) );
  NAND2_X1 U7472 ( .A1(n9226), .A2(n7102), .ZN(n7032) );
  NAND2_X1 U7473 ( .A1(n7848), .A2(n7032), .ZN(n6964) );
  NAND2_X1 U7474 ( .A1(n6962), .A2(n6964), .ZN(n6961) );
  NAND2_X1 U7475 ( .A1(n7092), .A2(n7102), .ZN(n5854) );
  NAND2_X1 U7476 ( .A1(n6961), .A2(n5854), .ZN(n7031) );
  INV_X1 U7477 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7042) );
  OR2_X1 U7478 ( .A1(n4979), .A2(n7042), .ZN(n5861) );
  INV_X1 U7479 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6430) );
  NAND2_X1 U7480 ( .A1(n5855), .A2(n6430), .ZN(n5856) );
  NAND2_X1 U7481 ( .A1(n5868), .A2(n5856), .ZN(n7183) );
  OR2_X1 U7482 ( .A1(n6131), .A2(n7183), .ZN(n5860) );
  INV_X1 U7483 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n5857) );
  OR2_X1 U7484 ( .A1(n6072), .A2(n5857), .ZN(n5859) );
  INV_X1 U7485 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6427) );
  OR2_X1 U7486 ( .A1(n5790), .A2(n6427), .ZN(n5858) );
  NAND2_X1 U7487 ( .A1(n5850), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5862) );
  XNOR2_X1 U7488 ( .A(n5862), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6437) );
  INV_X1 U7489 ( .A(n6437), .ZN(n6441) );
  OR2_X1 U7490 ( .A1(n5863), .A2(n6344), .ZN(n5865) );
  OR2_X1 U7491 ( .A1(n7820), .A2(n6345), .ZN(n5864) );
  OAI211_X1 U7492 ( .C1(n6361), .C2(n6441), .A(n5865), .B(n5864), .ZN(n7185)
         );
  NAND2_X1 U7493 ( .A1(n7177), .A2(n7185), .ZN(n7113) );
  INV_X1 U7494 ( .A(n7177), .ZN(n9225) );
  NAND2_X1 U7495 ( .A1(n9225), .A2(n7176), .ZN(n7851) );
  NAND2_X1 U7496 ( .A1(n7113), .A2(n7851), .ZN(n7840) );
  NAND2_X1 U7497 ( .A1(n7177), .A2(n7176), .ZN(n5866) );
  INV_X1 U7498 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n9561) );
  OR2_X1 U7499 ( .A1(n4979), .A2(n9561), .ZN(n5874) );
  NAND2_X1 U7500 ( .A1(n5868), .A2(n5867), .ZN(n5869) );
  NAND2_X1 U7501 ( .A1(n5877), .A2(n5869), .ZN(n9560) );
  OR2_X1 U7502 ( .A1(n6131), .A2(n9560), .ZN(n5873) );
  INV_X1 U7503 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5870) );
  OR2_X1 U7504 ( .A1(n6072), .A2(n5870), .ZN(n5872) );
  INV_X1 U7505 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6442) );
  OR2_X1 U7506 ( .A1(n5790), .A2(n6442), .ZN(n5871) );
  NOR2_X1 U7507 ( .A1(n5850), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5948) );
  OR2_X1 U7508 ( .A1(n5948), .A2(n4808), .ZN(n5885) );
  XNOR2_X1 U7509 ( .A(n5885), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6472) );
  INV_X1 U7510 ( .A(n6472), .ZN(n6467) );
  OR2_X1 U7511 ( .A1(n7820), .A2(n6348), .ZN(n5875) );
  NAND2_X1 U7512 ( .A1(n7441), .A2(n9564), .ZN(n7857) );
  INV_X1 U7513 ( .A(n7441), .ZN(n9224) );
  NAND2_X1 U7514 ( .A1(n9224), .A2(n7437), .ZN(n7850) );
  NAND2_X1 U7515 ( .A1(n7857), .A2(n7850), .ZN(n7115) );
  INV_X1 U7516 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7254) );
  OR2_X1 U7517 ( .A1(n4979), .A2(n7254), .ZN(n5883) );
  INV_X1 U7518 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5876) );
  NAND2_X1 U7519 ( .A1(n5877), .A2(n5876), .ZN(n5878) );
  NAND2_X1 U7520 ( .A1(n5893), .A2(n5878), .ZN(n7453) );
  OR2_X1 U7521 ( .A1(n6131), .A2(n7453), .ZN(n5882) );
  INV_X1 U7522 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n5879) );
  OR2_X1 U7523 ( .A1(n6072), .A2(n5879), .ZN(n5881) );
  INV_X1 U7524 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6468) );
  OR2_X1 U7525 ( .A1(n5790), .A2(n6468), .ZN(n5880) );
  NAND2_X1 U7526 ( .A1(n6354), .A2(n7818), .ZN(n5889) );
  INV_X1 U7527 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5884) );
  NAND2_X1 U7528 ( .A1(n5885), .A2(n5884), .ZN(n5886) );
  NAND2_X1 U7529 ( .A1(n5886), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5887) );
  XNOR2_X1 U7530 ( .A(n5887), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6671) );
  AOI22_X1 U7531 ( .A1(n5986), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5985), .B2(
        n6671), .ZN(n5888) );
  NAND2_X1 U7532 ( .A1(n5889), .A2(n5888), .ZN(n7455) );
  NAND2_X1 U7533 ( .A1(n7445), .A2(n7455), .ZN(n7874) );
  INV_X1 U7534 ( .A(n7455), .ZN(n10142) );
  INV_X1 U7535 ( .A(n7445), .ZN(n9223) );
  NAND2_X1 U7536 ( .A1(n10142), .A2(n9223), .ZN(n7862) );
  NAND2_X1 U7537 ( .A1(n7874), .A2(n7862), .ZN(n7252) );
  NAND2_X1 U7538 ( .A1(n7253), .A2(n7252), .ZN(n7251) );
  NAND2_X1 U7539 ( .A1(n7445), .A2(n10142), .ZN(n5890) );
  NAND2_X1 U7540 ( .A1(n7251), .A2(n5890), .ZN(n7278) );
  INV_X1 U7541 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n5891) );
  OR2_X1 U7542 ( .A1(n4979), .A2(n5891), .ZN(n5899) );
  NAND2_X1 U7543 ( .A1(n5893), .A2(n5892), .ZN(n5894) );
  NAND2_X1 U7544 ( .A1(n5918), .A2(n5894), .ZN(n7293) );
  OR2_X1 U7545 ( .A1(n6131), .A2(n7293), .ZN(n5898) );
  INV_X1 U7546 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5895) );
  OR2_X1 U7547 ( .A1(n6072), .A2(n5895), .ZN(n5897) );
  INV_X1 U7548 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6676) );
  OR2_X1 U7549 ( .A1(n5790), .A2(n6676), .ZN(n5896) );
  NAND2_X1 U7550 ( .A1(n6357), .A2(n7818), .ZN(n5907) );
  AND2_X1 U7551 ( .A1(n5948), .A2(n5900), .ZN(n5903) );
  NOR2_X1 U7552 ( .A1(n5903), .A2(n4808), .ZN(n5901) );
  MUX2_X1 U7553 ( .A(n4808), .B(n5901), .S(P1_IR_REG_10__SCAN_IN), .Z(n5902)
         );
  INV_X1 U7554 ( .A(n5902), .ZN(n5905) );
  INV_X1 U7555 ( .A(n5912), .ZN(n5904) );
  AOI22_X1 U7556 ( .A1(n5986), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5985), .B2(
        n6788), .ZN(n5906) );
  OR2_X1 U7557 ( .A1(n7542), .A2(n9049), .ZN(n7865) );
  NAND2_X1 U7558 ( .A1(n9049), .A2(n7542), .ZN(n7863) );
  NAND2_X1 U7559 ( .A1(n7865), .A2(n7863), .ZN(n7964) );
  NAND2_X1 U7560 ( .A1(n7278), .A2(n7964), .ZN(n7277) );
  INV_X1 U7561 ( .A(n7542), .ZN(n9222) );
  OR2_X1 U7562 ( .A1(n9049), .A2(n9222), .ZN(n5908) );
  NAND2_X1 U7563 ( .A1(n6392), .A2(n7818), .ZN(n5915) );
  NOR2_X1 U7564 ( .A1(n5912), .A2(n4808), .ZN(n5909) );
  MUX2_X1 U7565 ( .A(n4808), .B(n5909), .S(P1_IR_REG_11__SCAN_IN), .Z(n5910)
         );
  INV_X1 U7566 ( .A(n5910), .ZN(n5913) );
  INV_X1 U7567 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5911) );
  NAND2_X1 U7568 ( .A1(n5912), .A2(n5911), .ZN(n5935) );
  AOI22_X1 U7569 ( .A1(n5986), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5985), .B2(
        n6872), .ZN(n5914) );
  INV_X1 U7570 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7341) );
  INV_X1 U7571 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n5916) );
  OR2_X1 U7572 ( .A1(n6072), .A2(n5916), .ZN(n5917) );
  OAI21_X1 U7573 ( .B1(n4979), .B2(n7341), .A(n5917), .ZN(n5922) );
  INV_X1 U7574 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6797) );
  NAND2_X1 U7575 ( .A1(n5918), .A2(n6797), .ZN(n5919) );
  NAND2_X1 U7576 ( .A1(n5927), .A2(n5919), .ZN(n7660) );
  INV_X1 U7577 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6794) );
  OR2_X1 U7578 ( .A1(n5790), .A2(n6794), .ZN(n5920) );
  OAI21_X1 U7579 ( .B1(n6131), .B2(n7660), .A(n5920), .ZN(n5921) );
  NAND2_X1 U7580 ( .A1(n6450), .A2(n7818), .ZN(n5925) );
  NAND2_X1 U7581 ( .A1(n5935), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5923) );
  XNOR2_X1 U7582 ( .A(n5923), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7079) );
  AOI22_X1 U7583 ( .A1(n5986), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5985), .B2(
        n7079), .ZN(n5924) );
  INV_X1 U7584 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n5926) );
  OR2_X1 U7585 ( .A1(n4979), .A2(n5926), .ZN(n5934) );
  NAND2_X1 U7586 ( .A1(n5927), .A2(n6876), .ZN(n5928) );
  NAND2_X1 U7587 ( .A1(n5939), .A2(n5928), .ZN(n7559) );
  OR2_X1 U7588 ( .A1(n6131), .A2(n7559), .ZN(n5933) );
  INV_X1 U7589 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n5929) );
  OR2_X1 U7590 ( .A1(n6072), .A2(n5929), .ZN(n5932) );
  INV_X1 U7591 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n5930) );
  OR2_X1 U7592 ( .A1(n5790), .A2(n5930), .ZN(n5931) );
  NAND2_X1 U7593 ( .A1(n7561), .A2(n7552), .ZN(n7868) );
  NAND2_X1 U7594 ( .A1(n7870), .A2(n7868), .ZN(n7969) );
  NAND2_X1 U7595 ( .A1(n6570), .A2(n7818), .ZN(n5938) );
  OAI21_X1 U7596 ( .B1(n5935), .B2(P1_IR_REG_12__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5936) );
  XNOR2_X1 U7597 ( .A(n5936), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7262) );
  AOI22_X1 U7598 ( .A1(n5986), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5985), .B2(
        n7262), .ZN(n5937) );
  INV_X1 U7599 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7493) );
  OR2_X1 U7600 ( .A1(n4979), .A2(n7493), .ZN(n5945) );
  NAND2_X1 U7601 ( .A1(n5939), .A2(n7085), .ZN(n5940) );
  NAND2_X1 U7602 ( .A1(n5955), .A2(n5940), .ZN(n7587) );
  OR2_X1 U7603 ( .A1(n6131), .A2(n7587), .ZN(n5944) );
  INV_X1 U7604 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n5941) );
  OR2_X1 U7605 ( .A1(n6072), .A2(n5941), .ZN(n5943) );
  INV_X1 U7606 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7082) );
  OR2_X1 U7607 ( .A1(n5790), .A2(n7082), .ZN(n5942) );
  OR2_X1 U7608 ( .A1(n7589), .A2(n7594), .ZN(n7882) );
  NAND2_X1 U7609 ( .A1(n7589), .A2(n7594), .ZN(n7880) );
  INV_X1 U7610 ( .A(n7594), .ZN(n9219) );
  NAND2_X1 U7611 ( .A1(n6595), .A2(n7818), .ZN(n5953) );
  INV_X1 U7612 ( .A(n5946), .ZN(n5947) );
  NAND2_X1 U7613 ( .A1(n5948), .A2(n5947), .ZN(n5950) );
  NAND2_X1 U7614 ( .A1(n5950), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5949) );
  MUX2_X1 U7615 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5949), .S(
        P1_IR_REG_14__SCAN_IN), .Z(n5951) );
  OR2_X1 U7616 ( .A1(n5950), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n5962) );
  AOI22_X1 U7617 ( .A1(n5986), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5985), .B2(
        n9261), .ZN(n5952) );
  INV_X1 U7618 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5954) );
  NAND2_X1 U7619 ( .A1(n5955), .A2(n5954), .ZN(n5956) );
  NAND2_X1 U7620 ( .A1(n5966), .A2(n5956), .ZN(n7617) );
  OR2_X1 U7621 ( .A1(n6131), .A2(n7617), .ZN(n5961) );
  INV_X1 U7622 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7598) );
  OR2_X1 U7623 ( .A1(n4979), .A2(n7598), .ZN(n5960) );
  INV_X1 U7624 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7266) );
  OR2_X1 U7625 ( .A1(n5790), .A2(n7266), .ZN(n5959) );
  INV_X1 U7626 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n5957) );
  OR2_X1 U7627 ( .A1(n6072), .A2(n5957), .ZN(n5958) );
  NAND2_X1 U7628 ( .A1(n10164), .A2(n7626), .ZN(n7776) );
  NAND2_X1 U7629 ( .A1(n7774), .A2(n7776), .ZN(n7971) );
  NAND2_X1 U7630 ( .A1(n6690), .A2(n7818), .ZN(n5965) );
  NAND2_X1 U7631 ( .A1(n5962), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5963) );
  XNOR2_X1 U7632 ( .A(n5963), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9273) );
  AOI22_X1 U7633 ( .A1(n5986), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5985), .B2(
        n9273), .ZN(n5964) );
  INV_X1 U7634 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7629) );
  OR2_X1 U7635 ( .A1(n4979), .A2(n7629), .ZN(n5973) );
  INV_X1 U7636 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9266) );
  NAND2_X1 U7637 ( .A1(n5966), .A2(n9266), .ZN(n5967) );
  NAND2_X1 U7638 ( .A1(n5978), .A2(n5967), .ZN(n9199) );
  OR2_X1 U7639 ( .A1(n6131), .A2(n9199), .ZN(n5972) );
  INV_X1 U7640 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n5968) );
  OR2_X1 U7641 ( .A1(n6072), .A2(n5968), .ZN(n5971) );
  INV_X1 U7642 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n5969) );
  OR2_X1 U7643 ( .A1(n5790), .A2(n5969), .ZN(n5970) );
  NAND2_X1 U7644 ( .A1(n6765), .A2(n7818), .ZN(n5977) );
  NAND2_X1 U7645 ( .A1(n5974), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5975) );
  XNOR2_X1 U7646 ( .A(n5975), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9294) );
  AOI22_X1 U7647 ( .A1(n5986), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5985), .B2(
        n9294), .ZN(n5976) );
  INV_X1 U7648 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7692) );
  OR2_X1 U7649 ( .A1(n4979), .A2(n7692), .ZN(n5983) );
  NAND2_X1 U7650 ( .A1(n5978), .A2(n9286), .ZN(n5979) );
  NAND2_X1 U7651 ( .A1(n5991), .A2(n5979), .ZN(n9124) );
  OR2_X1 U7652 ( .A1(n6131), .A2(n9124), .ZN(n5982) );
  INV_X1 U7653 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9954) );
  OR2_X1 U7654 ( .A1(n6072), .A2(n9954), .ZN(n5981) );
  INV_X1 U7655 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9845) );
  OR2_X1 U7656 ( .A1(n5790), .A2(n9845), .ZN(n5980) );
  OR2_X1 U7657 ( .A1(n9126), .A2(n9132), .ZN(n7897) );
  NAND2_X1 U7658 ( .A1(n9126), .A2(n9132), .ZN(n9547) );
  INV_X1 U7659 ( .A(n9132), .ZN(n9218) );
  NAND2_X1 U7660 ( .A1(n6864), .A2(n7818), .ZN(n5988) );
  XNOR2_X1 U7661 ( .A(n5984), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9317) );
  AOI22_X1 U7662 ( .A1(n5986), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5985), .B2(
        n9317), .ZN(n5987) );
  INV_X1 U7663 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9292) );
  INV_X1 U7664 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9773) );
  OR2_X1 U7665 ( .A1(n6072), .A2(n9773), .ZN(n5989) );
  OAI21_X1 U7666 ( .B1(n4979), .B2(n9292), .A(n5989), .ZN(n5994) );
  XNOR2_X1 U7667 ( .A(n5991), .B(n5990), .ZN(n9541) );
  INV_X1 U7668 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9295) );
  OR2_X1 U7669 ( .A1(n5790), .A2(n9295), .ZN(n5992) );
  OAI21_X1 U7670 ( .B1(n6131), .B2(n9541), .A(n5992), .ZN(n5993) );
  NOR2_X1 U7671 ( .A1(n9636), .A2(n9217), .ZN(n5995) );
  INV_X1 U7672 ( .A(n9217), .ZN(n8941) );
  INV_X1 U7673 ( .A(n9636), .ZN(n9544) );
  AOI21_X1 U7674 ( .B1(n9531), .B2(n9216), .A(n9525), .ZN(n5997) );
  NOR2_X1 U7675 ( .A1(n9531), .A2(n9216), .ZN(n5996) );
  OR2_X1 U7676 ( .A1(n9625), .A2(n9175), .ZN(n7920) );
  NAND2_X1 U7677 ( .A1(n9625), .A2(n9175), .ZN(n7917) );
  NAND2_X1 U7678 ( .A1(n7920), .A2(n7917), .ZN(n9516) );
  NAND2_X1 U7679 ( .A1(n7107), .A2(n7818), .ZN(n5999) );
  OR2_X1 U7680 ( .A1(n7820), .A2(n9766), .ZN(n5998) );
  INV_X1 U7681 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n9506) );
  OR2_X1 U7682 ( .A1(n4979), .A2(n9506), .ZN(n6007) );
  INV_X1 U7683 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n6001) );
  NAND2_X1 U7684 ( .A1(n6002), .A2(n6001), .ZN(n6003) );
  NAND2_X1 U7685 ( .A1(n6012), .A2(n6003), .ZN(n9505) );
  OR2_X1 U7686 ( .A1(n6131), .A2(n9505), .ZN(n6006) );
  INV_X1 U7687 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9944) );
  OR2_X1 U7688 ( .A1(n6072), .A2(n9944), .ZN(n6005) );
  INV_X1 U7689 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9840) );
  OR2_X1 U7690 ( .A1(n5790), .A2(n9840), .ZN(n6004) );
  NAND2_X1 U7691 ( .A1(n9946), .A2(n9060), .ZN(n6009) );
  NOR2_X1 U7692 ( .A1(n9946), .A2(n9060), .ZN(n6008) );
  NAND2_X1 U7693 ( .A1(n7189), .A2(n7818), .ZN(n6011) );
  OR2_X1 U7694 ( .A1(n7820), .A2(n7190), .ZN(n6010) );
  INV_X1 U7695 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9101) );
  NAND2_X1 U7696 ( .A1(n6012), .A2(n9101), .ZN(n6013) );
  NAND2_X1 U7697 ( .A1(n6025), .A2(n6013), .ZN(n9487) );
  INV_X1 U7698 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9786) );
  OR2_X1 U7699 ( .A1(n5790), .A2(n9786), .ZN(n6014) );
  OAI21_X1 U7700 ( .B1(n9487), .B2(n6131), .A(n6014), .ZN(n6017) );
  INV_X1 U7701 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9488) );
  INV_X1 U7702 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9940) );
  OR2_X1 U7703 ( .A1(n6072), .A2(n9940), .ZN(n6015) );
  OAI21_X1 U7704 ( .B1(n4979), .B2(n9488), .A(n6015), .ZN(n6016) );
  NAND2_X1 U7705 ( .A1(n9486), .A2(n9213), .ZN(n6018) );
  NAND2_X1 U7706 ( .A1(n9484), .A2(n6018), .ZN(n6020) );
  NAND2_X1 U7707 ( .A1(n9942), .A2(n9160), .ZN(n6019) );
  NAND2_X1 U7708 ( .A1(n7301), .A2(n7818), .ZN(n6022) );
  OR2_X1 U7709 ( .A1(n7820), .A2(n7306), .ZN(n6021) );
  INV_X1 U7710 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9674) );
  INV_X1 U7711 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n6024) );
  NAND2_X1 U7712 ( .A1(n6025), .A2(n6024), .ZN(n6026) );
  NAND2_X1 U7713 ( .A1(n6035), .A2(n6026), .ZN(n9471) );
  OR2_X1 U7714 ( .A1(n9471), .A2(n6131), .ZN(n6028) );
  AOI22_X1 U7715 ( .A1(n5763), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n6133), .B2(
        P1_REG0_REG_22__SCAN_IN), .ZN(n6027) );
  OAI211_X1 U7716 ( .C1(n5790), .C2(n9674), .A(n6028), .B(n6027), .ZN(n9212)
         );
  NOR2_X1 U7717 ( .A1(n9474), .A2(n9212), .ZN(n6030) );
  NAND2_X1 U7718 ( .A1(n9474), .A2(n9212), .ZN(n6029) );
  NAND2_X1 U7719 ( .A1(n7310), .A2(n7818), .ZN(n6032) );
  OR2_X1 U7720 ( .A1(n7820), .A2(n7313), .ZN(n6031) );
  INV_X1 U7721 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6034) );
  NAND2_X1 U7722 ( .A1(n6035), .A2(n6034), .ZN(n6036) );
  NAND2_X1 U7723 ( .A1(n6055), .A2(n6036), .ZN(n9038) );
  OR2_X1 U7724 ( .A1(n9038), .A2(n6131), .ZN(n6040) );
  AOI22_X1 U7725 ( .A1(n5763), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n6133), .B2(
        P1_REG0_REG_23__SCAN_IN), .ZN(n6039) );
  INV_X1 U7726 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n6037) );
  OR2_X1 U7727 ( .A1(n5790), .A2(n6037), .ZN(n6038) );
  NOR2_X1 U7728 ( .A1(n9456), .A2(n9161), .ZN(n6041) );
  NAND2_X1 U7729 ( .A1(n9456), .A2(n9161), .ZN(n6042) );
  NAND2_X1 U7730 ( .A1(n7378), .A2(n7818), .ZN(n6044) );
  OR2_X1 U7731 ( .A1(n7820), .A2(n7379), .ZN(n6043) );
  XNOR2_X1 U7732 ( .A(n6055), .B(P1_REG3_REG_24__SCAN_IN), .ZN(n9444) );
  INV_X1 U7733 ( .A(n6131), .ZN(n6098) );
  NAND2_X1 U7734 ( .A1(n9444), .A2(n6098), .ZN(n6050) );
  INV_X1 U7735 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n6047) );
  INV_X1 U7736 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9665) );
  OR2_X1 U7737 ( .A1(n6072), .A2(n9665), .ZN(n6046) );
  INV_X1 U7738 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9602) );
  OR2_X1 U7739 ( .A1(n5790), .A2(n9602), .ZN(n6045) );
  OAI211_X1 U7740 ( .C1(n4979), .C2(n6047), .A(n6046), .B(n6045), .ZN(n6048)
         );
  INV_X1 U7741 ( .A(n6048), .ZN(n6049) );
  NAND2_X1 U7742 ( .A1(n6050), .A2(n6049), .ZN(n9211) );
  NOR2_X1 U7743 ( .A1(n9443), .A2(n9211), .ZN(n6052) );
  NAND2_X1 U7744 ( .A1(n9443), .A2(n9211), .ZN(n6051) );
  NAND2_X1 U7745 ( .A1(n7407), .A2(n7818), .ZN(n6054) );
  OR2_X1 U7746 ( .A1(n7820), .A2(n9923), .ZN(n6053) );
  INV_X1 U7747 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9142) );
  INV_X1 U7748 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9109) );
  OAI21_X1 U7749 ( .B1(n6055), .B2(n9142), .A(n9109), .ZN(n6056) );
  AND2_X1 U7750 ( .A1(n6056), .A2(n6068), .ZN(n9428) );
  NAND2_X1 U7751 ( .A1(n9428), .A2(n6098), .ZN(n6062) );
  INV_X1 U7752 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n6059) );
  INV_X1 U7753 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9661) );
  OR2_X1 U7754 ( .A1(n6072), .A2(n9661), .ZN(n6058) );
  INV_X1 U7755 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9597) );
  OR2_X1 U7756 ( .A1(n5790), .A2(n9597), .ZN(n6057) );
  OAI211_X1 U7757 ( .C1(n4979), .C2(n6059), .A(n6058), .B(n6057), .ZN(n6060)
         );
  INV_X1 U7758 ( .A(n6060), .ZN(n6061) );
  NOR2_X1 U7759 ( .A1(n9663), .A2(n9186), .ZN(n6064) );
  NAND2_X1 U7760 ( .A1(n9663), .A2(n9186), .ZN(n6063) );
  NAND2_X1 U7761 ( .A1(n7500), .A2(n7818), .ZN(n6066) );
  OR2_X1 U7762 ( .A1(n7820), .A2(n7501), .ZN(n6065) );
  INV_X1 U7763 ( .A(n6068), .ZN(n6067) );
  NAND2_X1 U7764 ( .A1(n6067), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6084) );
  INV_X1 U7765 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9775) );
  NAND2_X1 U7766 ( .A1(n6068), .A2(n9775), .ZN(n6069) );
  NAND2_X1 U7767 ( .A1(n6084), .A2(n6069), .ZN(n9405) );
  INV_X1 U7768 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n6075) );
  INV_X1 U7769 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n6070) );
  OR2_X1 U7770 ( .A1(n5790), .A2(n6070), .ZN(n6074) );
  INV_X1 U7771 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n6071) );
  OR2_X1 U7772 ( .A1(n6072), .A2(n6071), .ZN(n6073) );
  OAI211_X1 U7773 ( .C1(n4979), .C2(n6075), .A(n6074), .B(n6073), .ZN(n6076)
         );
  INV_X1 U7774 ( .A(n6076), .ZN(n6077) );
  NOR2_X1 U7775 ( .A1(n9590), .A2(n9209), .ZN(n6079) );
  INV_X1 U7776 ( .A(n9209), .ZN(n7749) );
  NAND2_X1 U7777 ( .A1(n7564), .A2(n7818), .ZN(n6081) );
  OR2_X1 U7778 ( .A1(n7820), .A2(n7635), .ZN(n6080) );
  INV_X1 U7779 ( .A(n6084), .ZN(n6082) );
  NAND2_X1 U7780 ( .A1(n6082), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n9379) );
  INV_X1 U7781 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6083) );
  NAND2_X1 U7782 ( .A1(n6084), .A2(n6083), .ZN(n6085) );
  NAND2_X1 U7783 ( .A1(n9379), .A2(n6085), .ZN(n9391) );
  OR2_X1 U7784 ( .A1(n9391), .A2(n6131), .ZN(n6090) );
  INV_X1 U7785 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n9390) );
  INV_X1 U7786 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9656) );
  OR2_X1 U7787 ( .A1(n6072), .A2(n9656), .ZN(n6087) );
  INV_X1 U7788 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9587) );
  OR2_X1 U7789 ( .A1(n5790), .A2(n9587), .ZN(n6086) );
  OAI211_X1 U7790 ( .C1(n4979), .C2(n9390), .A(n6087), .B(n6086), .ZN(n6088)
         );
  INV_X1 U7791 ( .A(n6088), .ZN(n6089) );
  OR2_X1 U7792 ( .A1(n9389), .A2(n9187), .ZN(n7751) );
  NAND2_X1 U7793 ( .A1(n9389), .A2(n9187), .ZN(n7934) );
  NAND2_X1 U7794 ( .A1(n7603), .A2(n7818), .ZN(n6092) );
  OR2_X1 U7795 ( .A1(n7820), .A2(n7637), .ZN(n6091) );
  XNOR2_X1 U7796 ( .A(n9379), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n9076) );
  INV_X1 U7797 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n6096) );
  INV_X1 U7798 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6093) );
  OR2_X1 U7799 ( .A1(n5790), .A2(n6093), .ZN(n6095) );
  INV_X1 U7800 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9740) );
  OR2_X1 U7801 ( .A1(n6072), .A2(n9740), .ZN(n6094) );
  OAI211_X1 U7802 ( .C1(n4979), .C2(n6096), .A(n6095), .B(n6094), .ZN(n6097)
         );
  NAND2_X1 U7803 ( .A1(n9071), .A2(n9372), .ZN(n9367) );
  NAND2_X1 U7804 ( .A1(n6099), .A2(n9368), .ZN(n9365) );
  NAND2_X1 U7805 ( .A1(n9365), .A2(n6100), .ZN(n8025) );
  NAND2_X1 U7806 ( .A1(n8015), .A2(n7757), .ZN(n7998) );
  NAND2_X1 U7807 ( .A1(n6102), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6103) );
  MUX2_X1 U7808 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6103), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n6104) );
  NAND2_X1 U7809 ( .A1(n6104), .A2(n4416), .ZN(n7108) );
  INV_X1 U7810 ( .A(n8012), .ZN(n6170) );
  OR2_X1 U7811 ( .A1(n7998), .A2(n6170), .ZN(n7010) );
  INV_X1 U7812 ( .A(n7108), .ZN(n8002) );
  AOI21_X1 U7813 ( .B1(n7304), .B2(n8002), .A(n8005), .ZN(n6105) );
  NAND3_X1 U7814 ( .A1(n7010), .A2(n6105), .A3(n7009), .ZN(n7330) );
  INV_X1 U7815 ( .A(n10148), .ZN(n10168) );
  INV_X1 U7816 ( .A(n10161), .ZN(n9639) );
  NAND2_X1 U7817 ( .A1(n10077), .A2(n5810), .ZN(n7130) );
  OR2_X1 U7818 ( .A1(n7130), .A2(n7136), .ZN(n7131) );
  NAND2_X1 U7819 ( .A1(n7039), .A2(n7176), .ZN(n7111) );
  INV_X1 U7820 ( .A(n9049), .ZN(n7296) );
  NAND2_X1 U7821 ( .A1(n7630), .A2(n4656), .ZN(n7693) );
  NOR2_X2 U7822 ( .A1(n4978), .A2(n9636), .ZN(n9539) );
  INV_X1 U7823 ( .A(n9474), .ZN(n9610) );
  NAND2_X1 U7824 ( .A1(n9485), .A2(n9610), .ZN(n9451) );
  INV_X1 U7825 ( .A(n6107), .ZN(n9388) );
  OAI211_X1 U7826 ( .C1(n9388), .C2(n9362), .A(n10094), .B(n9377), .ZN(n8018)
         );
  INV_X1 U7827 ( .A(n6108), .ZN(n7960) );
  INV_X1 U7828 ( .A(n6626), .ZN(n10095) );
  INV_X2 U7829 ( .A(n6702), .ZN(n9230) );
  NOR2_X1 U7830 ( .A1(n9230), .A2(n6106), .ZN(n6110) );
  AOI21_X1 U7831 ( .B1(n7960), .B2(n10086), .A(n6110), .ZN(n10070) );
  NAND2_X1 U7832 ( .A1(n10070), .A2(n6111), .ZN(n6113) );
  INV_X1 U7833 ( .A(n7136), .ZN(n10135) );
  NAND2_X1 U7834 ( .A1(n9228), .A2(n10135), .ZN(n7836) );
  INV_X1 U7835 ( .A(n9228), .ZN(n6949) );
  NAND2_X1 U7836 ( .A1(n6949), .A2(n7136), .ZN(n7831) );
  AND2_X1 U7837 ( .A1(n7831), .A2(n7838), .ZN(n7844) );
  NAND2_X1 U7838 ( .A1(n6981), .A2(n7844), .ZN(n7033) );
  NAND2_X1 U7839 ( .A1(n7033), .A2(n7760), .ZN(n6965) );
  NAND2_X1 U7840 ( .A1(n7113), .A2(n7857), .ZN(n7853) );
  NAND2_X1 U7841 ( .A1(n6115), .A2(n7853), .ZN(n6114) );
  NAND2_X1 U7842 ( .A1(n6114), .A2(n7874), .ZN(n7965) );
  INV_X1 U7843 ( .A(n7848), .ZN(n7839) );
  NOR2_X1 U7844 ( .A1(n7965), .A2(n7839), .ZN(n7763) );
  NAND2_X1 U7845 ( .A1(n6965), .A2(n7763), .ZN(n6118) );
  INV_X1 U7846 ( .A(n7965), .ZN(n6117) );
  INV_X1 U7847 ( .A(n7851), .ZN(n7841) );
  NAND2_X1 U7848 ( .A1(n6117), .A2(n6116), .ZN(n7765) );
  NAND2_X1 U7849 ( .A1(n7384), .A2(n7866), .ZN(n6120) );
  INV_X1 U7850 ( .A(n7969), .ZN(n6119) );
  NAND2_X1 U7851 ( .A1(n6120), .A2(n6119), .ZN(n7485) );
  INV_X1 U7852 ( .A(n7491), .ZN(n7970) );
  INV_X1 U7853 ( .A(n7870), .ZN(n6121) );
  NOR2_X1 U7854 ( .A1(n7970), .A2(n6121), .ZN(n6122) );
  INV_X1 U7855 ( .A(n7774), .ZN(n7890) );
  NOR2_X1 U7856 ( .A1(n7879), .A2(n7890), .ZN(n6123) );
  NAND2_X1 U7857 ( .A1(n7623), .A2(n7891), .ZN(n7688) );
  NAND2_X1 U7858 ( .A1(n7688), .A2(n7974), .ZN(n9545) );
  NAND2_X1 U7859 ( .A1(n9545), .A2(n9547), .ZN(n6124) );
  XNOR2_X1 U7860 ( .A(n9636), .B(n9217), .ZN(n9549) );
  NAND2_X1 U7861 ( .A1(n6124), .A2(n9549), .ZN(n9548) );
  NAND2_X1 U7862 ( .A1(n9636), .A2(n8941), .ZN(n7898) );
  XNOR2_X1 U7863 ( .A(n9531), .B(n9216), .ZN(n9532) );
  INV_X1 U7864 ( .A(n9216), .ZN(n7753) );
  NAND2_X1 U7865 ( .A1(n9531), .A2(n7753), .ZN(n7916) );
  INV_X1 U7866 ( .A(n9516), .ZN(n9512) );
  XNOR2_X1 U7867 ( .A(n9486), .B(n9160), .ZN(n9483) );
  NAND2_X1 U7868 ( .A1(n9486), .A2(n9160), .ZN(n7909) );
  INV_X1 U7869 ( .A(n9212), .ZN(n9036) );
  OR2_X1 U7870 ( .A1(n9474), .A2(n9036), .ZN(n7922) );
  NAND2_X1 U7871 ( .A1(n9474), .A2(n9036), .ZN(n7910) );
  OR2_X1 U7872 ( .A1(n6126), .A2(n9161), .ZN(n7925) );
  NAND2_X1 U7873 ( .A1(n6126), .A2(n9161), .ZN(n9435) );
  INV_X1 U7874 ( .A(n9211), .ZN(n9037) );
  NAND2_X1 U7875 ( .A1(n9443), .A2(n9037), .ZN(n7929) );
  NAND2_X1 U7876 ( .A1(n9417), .A2(n7929), .ZN(n9436) );
  INV_X1 U7877 ( .A(n9435), .ZN(n7914) );
  NOR2_X1 U7878 ( .A1(n9436), .A2(n7914), .ZN(n6127) );
  NAND2_X1 U7879 ( .A1(n9457), .A2(n6127), .ZN(n9438) );
  INV_X1 U7880 ( .A(n9663), .ZN(n9427) );
  OR2_X1 U7881 ( .A1(n9427), .A2(n9186), .ZN(n7940) );
  NAND2_X1 U7882 ( .A1(n9427), .A2(n9186), .ZN(n7794) );
  NAND2_X1 U7883 ( .A1(n7940), .A2(n7794), .ZN(n9418) );
  INV_X1 U7884 ( .A(n9417), .ZN(n7931) );
  NOR2_X1 U7885 ( .A1(n9418), .A2(n7931), .ZN(n6128) );
  XNOR2_X1 U7886 ( .A(n9590), .B(n9209), .ZN(n9409) );
  NAND2_X1 U7887 ( .A1(n9590), .A2(n7749), .ZN(n7795) );
  INV_X1 U7888 ( .A(n7934), .ZN(n6129) );
  XNOR2_X1 U7889 ( .A(n9369), .B(n9368), .ZN(n6138) );
  NAND2_X1 U7890 ( .A1(n8015), .A2(n8005), .ZN(n7951) );
  NAND2_X1 U7891 ( .A1(n7757), .A2(n8002), .ZN(n8007) );
  INV_X1 U7892 ( .A(n9246), .ZN(n6371) );
  INV_X1 U7893 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6136) );
  INV_X1 U7894 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9378) );
  OR2_X1 U7895 ( .A1(n6131), .A2(n9378), .ZN(n6132) );
  OR2_X1 U7896 ( .A1(n9379), .A2(n6132), .ZN(n6135) );
  AOI22_X1 U7897 ( .A1(n5763), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n6133), .B2(
        P1_REG0_REG_29__SCAN_IN), .ZN(n6134) );
  OAI211_X1 U7898 ( .C1(n5790), .C2(n6136), .A(n6135), .B(n6134), .ZN(n9207)
         );
  NAND2_X1 U7899 ( .A1(n9246), .A2(n6620), .ZN(n9350) );
  NAND2_X1 U7900 ( .A1(n9207), .A2(n9150), .ZN(n6137) );
  OAI21_X1 U7901 ( .B1(n9187), .B2(n9373), .A(n6137), .ZN(n9080) );
  AOI21_X1 U7902 ( .B1(n6138), .B2(n10072), .A(n9080), .ZN(n8020) );
  OAI21_X1 U7903 ( .B1(n8025), .B2(n9639), .A(n6139), .ZN(n6176) );
  NAND2_X1 U7904 ( .A1(n6143), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6144) );
  MUX2_X1 U7905 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6144), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n6145) );
  AND2_X1 U7906 ( .A1(n6145), .A2(n4418), .ZN(n6153) );
  INV_X1 U7907 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U7908 ( .A1(n6148), .A2(n6147), .ZN(n6149) );
  NAND2_X1 U7909 ( .A1(n6149), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6151) );
  INV_X1 U7910 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6150) );
  NAND2_X1 U7911 ( .A1(n7408), .A2(P1_B_REG_SCAN_IN), .ZN(n6154) );
  INV_X1 U7912 ( .A(n6153), .ZN(n7380) );
  MUX2_X1 U7913 ( .A(P1_B_REG_SCAN_IN), .B(n6154), .S(n7380), .Z(n6155) );
  NOR4_X1 U7914 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n9688) );
  NOR2_X1 U7915 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .ZN(
        n6158) );
  NOR4_X1 U7916 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6157) );
  NOR4_X1 U7917 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6156) );
  NAND4_X1 U7918 ( .A1(n9688), .A2(n6158), .A3(n6157), .A4(n6156), .ZN(n6164)
         );
  NOR4_X1 U7919 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6162) );
  NOR4_X1 U7920 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n6161) );
  NOR4_X1 U7921 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n6160) );
  NOR4_X1 U7922 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6159) );
  NAND4_X1 U7923 ( .A1(n6162), .A2(n6161), .A3(n6160), .A4(n6159), .ZN(n6163)
         );
  NOR2_X1 U7924 ( .A1(n6164), .A2(n6163), .ZN(n6599) );
  NAND2_X1 U7925 ( .A1(n8013), .A2(n6599), .ZN(n6165) );
  NAND2_X1 U7926 ( .A1(n10116), .A2(n6165), .ZN(n6166) );
  INV_X1 U7927 ( .A(n6167), .ZN(n7502) );
  NAND2_X1 U7928 ( .A1(n7502), .A2(n7408), .ZN(n9958) );
  NAND2_X1 U7929 ( .A1(n10148), .A2(n7952), .ZN(n6623) );
  NAND2_X1 U7930 ( .A1(n6992), .A2(n6623), .ZN(n6173) );
  NAND2_X1 U7931 ( .A1(n7502), .A2(n7380), .ZN(n9959) );
  INV_X1 U7932 ( .A(n6602), .ZN(n6993) );
  NAND2_X1 U7933 ( .A1(n6176), .A2(n10174), .ZN(n6169) );
  NAND2_X1 U7934 ( .A1(n10173), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6168) );
  NAND2_X1 U7935 ( .A1(n6169), .A2(n6168), .ZN(n6172) );
  INV_X1 U7936 ( .A(n7009), .ZN(n6484) );
  NOR2_X1 U7937 ( .A1(n9362), .A2(n9956), .ZN(n6171) );
  OR2_X1 U7938 ( .A1(n6172), .A2(n6171), .ZN(P1_U3518) );
  OR3_X2 U7939 ( .A1(n6994), .A2(n6173), .A3(n6602), .ZN(n10184) );
  NAND2_X1 U7940 ( .A1(n10184), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6174) );
  OAI21_X1 U7941 ( .B1(n9362), .B2(n9646), .A(n6174), .ZN(n6175) );
  INV_X1 U7942 ( .A(n6178), .ZN(n6181) );
  INV_X1 U7943 ( .A(n6179), .ZN(n6180) );
  AND2_X1 U7944 ( .A1(n6183), .A2(n6182), .ZN(n6184) );
  XNOR2_X1 U7945 ( .A(n6284), .B(n8280), .ZN(n8276) );
  XOR2_X1 U7946 ( .A(n8400), .B(n8276), .Z(n6281) );
  INV_X1 U7947 ( .A(n8414), .ZN(n6187) );
  OR2_X1 U7948 ( .A1(n6189), .A2(n6187), .ZN(n6190) );
  NAND2_X1 U7949 ( .A1(n6189), .A2(n6188), .ZN(n6194) );
  NAND2_X1 U7950 ( .A1(n6190), .A2(n6194), .ZN(n6732) );
  INV_X1 U7951 ( .A(n6732), .ZN(n6193) );
  INV_X1 U7952 ( .A(n6684), .ZN(n6719) );
  NAND2_X1 U7953 ( .A1(n6191), .A2(n6719), .ZN(n6192) );
  NAND2_X1 U7954 ( .A1(n6730), .A2(n6194), .ZN(n6723) );
  XNOR2_X1 U7955 ( .A(n6195), .B(n8413), .ZN(n6724) );
  NAND2_X1 U7956 ( .A1(n6723), .A2(n6724), .ZN(n6722) );
  NAND2_X1 U7957 ( .A1(n6195), .A2(n6845), .ZN(n6196) );
  NAND2_X1 U7958 ( .A1(n6722), .A2(n6196), .ZN(n6810) );
  INV_X1 U7959 ( .A(n6810), .ZN(n6199) );
  XNOR2_X1 U7960 ( .A(n6861), .B(n6197), .ZN(n6200) );
  XNOR2_X1 U7961 ( .A(n6200), .B(n8763), .ZN(n6813) );
  INV_X1 U7962 ( .A(n6813), .ZN(n6198) );
  NAND2_X1 U7963 ( .A1(n6199), .A2(n6198), .ZN(n6811) );
  INV_X1 U7964 ( .A(n6200), .ZN(n6201) );
  INV_X1 U7965 ( .A(n8763), .ZN(n8412) );
  NAND2_X1 U7966 ( .A1(n6201), .A2(n8412), .ZN(n6202) );
  AND2_X1 U7967 ( .A1(n6811), .A2(n6202), .ZN(n6830) );
  XNOR2_X1 U7968 ( .A(n6833), .B(n8280), .ZN(n6203) );
  NAND2_X1 U7969 ( .A1(n6203), .A2(n6901), .ZN(n6885) );
  INV_X1 U7970 ( .A(n6203), .ZN(n6204) );
  INV_X1 U7971 ( .A(n6901), .ZN(n8411) );
  NAND2_X1 U7972 ( .A1(n6204), .A2(n8411), .ZN(n6205) );
  AND2_X1 U7973 ( .A1(n6885), .A2(n6205), .ZN(n6829) );
  NAND2_X1 U7974 ( .A1(n6830), .A2(n6829), .ZN(n6828) );
  NAND2_X1 U7975 ( .A1(n6828), .A2(n6885), .ZN(n6206) );
  XNOR2_X1 U7976 ( .A(n6902), .B(n8280), .ZN(n6207) );
  XNOR2_X1 U7977 ( .A(n6207), .B(n8410), .ZN(n6884) );
  NAND2_X1 U7978 ( .A1(n6206), .A2(n6884), .ZN(n6888) );
  NAND2_X1 U7979 ( .A1(n6207), .A2(n6823), .ZN(n6208) );
  NAND2_X1 U7980 ( .A1(n6888), .A2(n6208), .ZN(n7142) );
  INV_X1 U7981 ( .A(n7142), .ZN(n6210) );
  XNOR2_X1 U7982 ( .A(n7145), .B(n8280), .ZN(n6211) );
  XNOR2_X1 U7983 ( .A(n6211), .B(n7207), .ZN(n7143) );
  INV_X1 U7984 ( .A(n7143), .ZN(n6209) );
  INV_X1 U7985 ( .A(n6211), .ZN(n6212) );
  INV_X1 U7986 ( .A(n7207), .ZN(n8409) );
  NAND2_X1 U7987 ( .A1(n6212), .A2(n8409), .ZN(n6213) );
  XNOR2_X1 U7988 ( .A(n7199), .B(n8280), .ZN(n6214) );
  NAND2_X1 U7989 ( .A1(n6214), .A2(n6215), .ZN(n7320) );
  INV_X1 U7990 ( .A(n6214), .ZN(n6216) );
  INV_X1 U7991 ( .A(n6215), .ZN(n8408) );
  NAND2_X1 U7992 ( .A1(n6216), .A2(n8408), .ZN(n6217) );
  AND2_X1 U7993 ( .A1(n7320), .A2(n6217), .ZN(n7203) );
  XNOR2_X1 U7994 ( .A(n7326), .B(n8280), .ZN(n6220) );
  XNOR2_X1 U7995 ( .A(n6220), .B(n8407), .ZN(n7319) );
  NAND2_X1 U7996 ( .A1(n6218), .A2(n7319), .ZN(n7323) );
  NAND2_X1 U7997 ( .A1(n6220), .A2(n6219), .ZN(n6221) );
  INV_X1 U7998 ( .A(n7467), .ZN(n6223) );
  XNOR2_X1 U7999 ( .A(n10267), .B(n6191), .ZN(n6224) );
  XNOR2_X1 U8000 ( .A(n6224), .B(n8406), .ZN(n7468) );
  NAND2_X1 U8001 ( .A1(n6224), .A2(n8406), .ZN(n6225) );
  XNOR2_X1 U8002 ( .A(n10272), .B(n8280), .ZN(n7681) );
  XNOR2_X1 U8003 ( .A(n7394), .B(n8280), .ZN(n8302) );
  OAI21_X1 U8004 ( .B1(n7701), .B2(n7681), .A(n8302), .ZN(n6231) );
  XNOR2_X1 U8005 ( .A(n10282), .B(n6191), .ZN(n6232) );
  XNOR2_X1 U8006 ( .A(n6232), .B(n8403), .ZN(n8304) );
  NAND3_X1 U8007 ( .A1(n10272), .A2(n7701), .A3(n8280), .ZN(n6226) );
  OAI21_X1 U8008 ( .B1(n8280), .B2(n8404), .A(n6226), .ZN(n6229) );
  NAND2_X1 U8009 ( .A1(n7701), .A2(n6191), .ZN(n6227) );
  OAI22_X1 U8010 ( .A1(n10272), .A2(n6227), .B1(n6191), .B2(n8404), .ZN(n6228)
         );
  MUX2_X1 U8011 ( .A(n6229), .B(n6228), .S(n8086), .Z(n6230) );
  NAND2_X1 U8012 ( .A1(n6232), .A2(n8403), .ZN(n6233) );
  XNOR2_X1 U8013 ( .A(n7713), .B(n8280), .ZN(n6234) );
  NAND2_X1 U8014 ( .A1(n6234), .A2(n8308), .ZN(n7503) );
  INV_X1 U8015 ( .A(n6234), .ZN(n6235) );
  NAND2_X1 U8016 ( .A1(n6235), .A2(n8402), .ZN(n7504) );
  NAND2_X1 U8017 ( .A1(n6236), .A2(n7504), .ZN(n7568) );
  INV_X1 U8018 ( .A(n7568), .ZN(n6240) );
  XNOR2_X1 U8019 ( .A(n7736), .B(n6191), .ZN(n6237) );
  XNOR2_X1 U8020 ( .A(n6237), .B(n8742), .ZN(n7569) );
  INV_X1 U8021 ( .A(n7569), .ZN(n6239) );
  INV_X1 U8022 ( .A(n6237), .ZN(n6238) );
  XNOR2_X1 U8023 ( .A(n8907), .B(n8280), .ZN(n6241) );
  XNOR2_X1 U8024 ( .A(n6241), .B(n8730), .ZN(n7640) );
  INV_X1 U8025 ( .A(n6241), .ZN(n6242) );
  NAND2_X1 U8026 ( .A1(n6242), .A2(n8730), .ZN(n6243) );
  XNOR2_X1 U8027 ( .A(n8901), .B(n6191), .ZN(n6244) );
  XNOR2_X1 U8028 ( .A(n6244), .B(n8743), .ZN(n8326) );
  INV_X1 U8029 ( .A(n6244), .ZN(n6245) );
  NAND2_X1 U8030 ( .A1(n6245), .A2(n7644), .ZN(n8332) );
  NAND2_X1 U8031 ( .A1(n8324), .A2(n8332), .ZN(n6246) );
  XNOR2_X1 U8032 ( .A(n8818), .B(n8280), .ZN(n6247) );
  XNOR2_X1 U8033 ( .A(n6247), .B(n8731), .ZN(n8333) );
  NAND2_X1 U8034 ( .A1(n6246), .A2(n8333), .ZN(n8336) );
  NAND2_X1 U8035 ( .A1(n6247), .A2(n8377), .ZN(n6248) );
  NAND2_X1 U8036 ( .A1(n8336), .A2(n6248), .ZN(n8371) );
  XNOR2_X1 U8037 ( .A(n8894), .B(n8280), .ZN(n6249) );
  XNOR2_X1 U8038 ( .A(n6249), .B(n8714), .ZN(n8370) );
  NAND2_X1 U8039 ( .A1(n8371), .A2(n8370), .ZN(n6251) );
  NAND2_X1 U8040 ( .A1(n6249), .A2(n8692), .ZN(n6250) );
  XNOR2_X1 U8041 ( .A(n8889), .B(n8280), .ZN(n8268) );
  AND2_X1 U8042 ( .A1(n8268), .A2(n8357), .ZN(n6252) );
  XNOR2_X1 U8043 ( .A(n8883), .B(n8280), .ZN(n6253) );
  NAND2_X1 U8044 ( .A1(n6253), .A2(n8693), .ZN(n8291) );
  INV_X1 U8045 ( .A(n6253), .ZN(n6254) );
  NAND2_X1 U8046 ( .A1(n6254), .A2(n8663), .ZN(n6255) );
  NAND2_X1 U8047 ( .A1(n8291), .A2(n6255), .ZN(n8354) );
  XNOR2_X1 U8048 ( .A(n8877), .B(n8280), .ZN(n6258) );
  XNOR2_X1 U8049 ( .A(n6258), .B(n8676), .ZN(n8292) );
  NAND2_X1 U8050 ( .A1(n6256), .A2(n8292), .ZN(n8293) );
  NAND2_X1 U8051 ( .A1(n6258), .A2(n6257), .ZN(n6259) );
  INV_X1 U8052 ( .A(n8362), .ZN(n6261) );
  XNOR2_X1 U8053 ( .A(n8871), .B(n6191), .ZN(n6262) );
  XNOR2_X1 U8054 ( .A(n6262), .B(n8664), .ZN(n8361) );
  INV_X1 U8055 ( .A(n8361), .ZN(n6260) );
  NAND2_X1 U8056 ( .A1(n6262), .A2(n8664), .ZN(n6263) );
  XNOR2_X1 U8057 ( .A(n8865), .B(n8280), .ZN(n6264) );
  XNOR2_X1 U8058 ( .A(n8859), .B(n8280), .ZN(n6265) );
  NAND2_X1 U8059 ( .A1(n6265), .A2(n8614), .ZN(n8318) );
  INV_X1 U8060 ( .A(n6265), .ZN(n6266) );
  NAND2_X1 U8061 ( .A1(n6266), .A2(n8640), .ZN(n6267) );
  AND2_X1 U8062 ( .A1(n8318), .A2(n6267), .ZN(n8345) );
  XNOR2_X1 U8063 ( .A(n8853), .B(n8280), .ZN(n6268) );
  NAND2_X1 U8064 ( .A1(n6268), .A2(n8631), .ZN(n6271) );
  INV_X1 U8065 ( .A(n6268), .ZN(n6269) );
  NAND2_X1 U8066 ( .A1(n6269), .A2(n8401), .ZN(n6270) );
  NAND2_X1 U8067 ( .A1(n6271), .A2(n6270), .ZN(n8317) );
  INV_X1 U8068 ( .A(n6271), .ZN(n8385) );
  XNOR2_X1 U8069 ( .A(n8846), .B(n8280), .ZN(n6272) );
  XNOR2_X1 U8070 ( .A(n6272), .B(n8587), .ZN(n8384) );
  INV_X1 U8071 ( .A(n6275), .ZN(n6291) );
  NAND2_X1 U8072 ( .A1(n6276), .A2(n6291), .ZN(n6279) );
  OR2_X1 U8073 ( .A1(n6282), .A2(n6277), .ZN(n6278) );
  AOI211_X1 U8074 ( .C1(n6281), .C2(n6280), .A(n8381), .B(n8277), .ZN(n6305)
         );
  OR2_X1 U8075 ( .A1(n6282), .A2(n10274), .ZN(n6283) );
  NAND2_X1 U8076 ( .A1(n6284), .A2(n8379), .ZN(n6303) );
  NOR2_X1 U8077 ( .A1(n6285), .A2(n8027), .ZN(n6288) );
  INV_X1 U8078 ( .A(n6287), .ZN(n6286) );
  AOI22_X1 U8079 ( .A1(n8587), .A2(n8390), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n6300) );
  NAND2_X1 U8080 ( .A1(n6290), .A2(n6289), .ZN(n6294) );
  NAND2_X1 U8081 ( .A1(n6296), .A2(n6291), .ZN(n6292) );
  NAND4_X1 U8082 ( .A1(n6294), .A2(n6501), .A3(n6293), .A4(n6292), .ZN(n6298)
         );
  NOR2_X1 U8083 ( .A1(n8028), .A2(n8027), .ZN(n6295) );
  AND2_X1 U8084 ( .A1(n6296), .A2(n6295), .ZN(n6297) );
  AOI21_X1 U8085 ( .B1(n6298), .B2(P2_STATE_REG_SCAN_IN), .A(n6297), .ZN(n6709) );
  INV_X1 U8086 ( .A(n6318), .ZN(n6500) );
  NAND2_X1 U8087 ( .A1(n6500), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8243) );
  NAND2_X1 U8088 ( .A1(n8593), .A2(n8394), .ZN(n6299) );
  OAI211_X1 U8089 ( .C1(n8156), .C2(n8392), .A(n6300), .B(n6299), .ZN(n6301)
         );
  INV_X1 U8090 ( .A(n6301), .ZN(n6302) );
  NAND2_X1 U8091 ( .A1(n6303), .A2(n6302), .ZN(n6304) );
  INV_X1 U8092 ( .A(n6306), .ZN(n6307) );
  NOR2_X1 U8093 ( .A1(n6308), .A2(n6307), .ZN(n6311) );
  OR2_X1 U8094 ( .A1(n6313), .A2(n6312), .ZN(n6317) );
  INV_X1 U8095 ( .A(n10274), .ZN(n10281) );
  INV_X1 U8096 ( .A(n6315), .ZN(n6316) );
  NAND2_X1 U8097 ( .A1(n6317), .A2(n6316), .ZN(P2_U3488) );
  NAND2_X1 U8098 ( .A1(n6501), .A2(n8186), .ZN(n6319) );
  NAND2_X1 U8099 ( .A1(n6319), .A2(n6318), .ZN(n6513) );
  NAND2_X1 U8100 ( .A1(n6513), .A2(n5184), .ZN(n6320) );
  NAND2_X1 U8101 ( .A1(n6320), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U8102 ( .A(n6321), .ZN(n6322) );
  NOR2_X2 U8103 ( .A1(n6614), .A2(n6322), .ZN(P1_U3973) );
  INV_X1 U8104 ( .A(n6708), .ZN(n6396) );
  XNOR2_X1 U8105 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  NOR2_X1 U8106 ( .A1(n7813), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8916) );
  INV_X2 U8107 ( .A(n8916), .ZN(n8258) );
  NAND2_X1 U8108 ( .A1(n7813), .A2(P2_U3151), .ZN(n8918) );
  INV_X1 U8109 ( .A(n6519), .ZN(n6535) );
  OAI222_X1 U8110 ( .A1(n8258), .A2(n6323), .B1(n8918), .B2(n6326), .C1(
        P2_U3151), .C2(n6535), .ZN(P2_U3293) );
  OAI222_X1 U8111 ( .A1(n8258), .A2(n6324), .B1(n8918), .B2(n6341), .C1(
        P2_U3151), .C2(n6521), .ZN(P2_U3292) );
  AND2_X1 U8112 ( .A1(n7813), .A2(P1_U3086), .ZN(n9962) );
  INV_X2 U8113 ( .A(n9962), .ZN(n9966) );
  AND2_X1 U8114 ( .A1(n6325), .A2(P1_U3086), .ZN(n7309) );
  INV_X2 U8115 ( .A(n7309), .ZN(n9969) );
  OAI222_X1 U8116 ( .A1(n9966), .A2(n6327), .B1(n9969), .B2(n6326), .C1(
        P1_U3086), .C2(n9255), .ZN(P1_U3353) );
  OAI222_X1 U8117 ( .A1(n9966), .A2(n6328), .B1(n9969), .B2(n6332), .C1(
        P1_U3086), .C2(n6381), .ZN(P1_U3354) );
  INV_X1 U8118 ( .A(n6657), .ZN(n6534) );
  OAI222_X1 U8119 ( .A1(n8258), .A2(n6329), .B1(n8918), .B2(n6338), .C1(
        P2_U3151), .C2(n6534), .ZN(P2_U3291) );
  OAI222_X1 U8120 ( .A1(n8258), .A2(n6330), .B1(n8918), .B2(n6340), .C1(
        P2_U3151), .C2(n6668), .ZN(P2_U3290) );
  INV_X1 U8121 ( .A(n8918), .ZN(n7307) );
  INV_X1 U8122 ( .A(n7307), .ZN(n7567) );
  OAI222_X1 U8123 ( .A1(n10203), .A2(P2_U3151), .B1(n7567), .B2(n6332), .C1(
        n6331), .C2(n8258), .ZN(P2_U3294) );
  INV_X1 U8124 ( .A(n6913), .ZN(n6917) );
  OAI222_X1 U8125 ( .A1(n8258), .A2(n6333), .B1(n8918), .B2(n6335), .C1(
        P2_U3151), .C2(n6917), .ZN(P2_U3289) );
  OAI222_X1 U8126 ( .A1(n9966), .A2(n6336), .B1(n9969), .B2(n6335), .C1(
        P1_U3086), .C2(n6334), .ZN(P1_U3349) );
  OAI222_X1 U8127 ( .A1(n9966), .A2(n6339), .B1(n9969), .B2(n6338), .C1(
        P1_U3086), .C2(n6337), .ZN(P1_U3351) );
  OAI222_X1 U8128 ( .A1(n9966), .A2(n9808), .B1(n9969), .B2(n6340), .C1(
        P1_U3086), .C2(n6415), .ZN(P1_U3350) );
  OAI222_X1 U8129 ( .A1(n9966), .A2(n6342), .B1(n9969), .B2(n6341), .C1(
        P1_U3086), .C2(n6399), .ZN(P1_U3352) );
  OAI222_X1 U8130 ( .A1(n8258), .A2(n6343), .B1(n8918), .B2(n6344), .C1(
        P2_U3151), .C2(n4853), .ZN(P2_U3288) );
  OAI222_X1 U8131 ( .A1(n9966), .A2(n6345), .B1(n9969), .B2(n6344), .C1(
        P1_U3086), .C2(n6441), .ZN(P1_U3348) );
  INV_X1 U8132 ( .A(n6346), .ZN(n6347) );
  OAI222_X1 U8133 ( .A1(n8258), .A2(n9733), .B1(n8918), .B2(n6347), .C1(
        P2_U3151), .C2(n7160), .ZN(P2_U3287) );
  OAI222_X1 U8134 ( .A1(n9966), .A2(n6348), .B1(n9969), .B2(n6347), .C1(
        P1_U3086), .C2(n6467), .ZN(P1_U3347) );
  INV_X1 U8135 ( .A(n6349), .ZN(n6350) );
  NAND2_X1 U8136 ( .A1(n6350), .A2(n6352), .ZN(n6351) );
  OAI21_X1 U8137 ( .B1(n6353), .B2(n6352), .A(n6351), .ZN(P2_U3377) );
  INV_X1 U8138 ( .A(n6354), .ZN(n6355) );
  INV_X1 U8139 ( .A(n6671), .ZN(n6675) );
  OAI222_X1 U8140 ( .A1(n9969), .A2(n6355), .B1(n6675), .B2(P1_U3086), .C1(
        n9798), .C2(n9966), .ZN(P1_U3346) );
  OAI222_X1 U8141 ( .A1(n8258), .A2(n6356), .B1(n7567), .B2(n6355), .C1(n7229), 
        .C2(P2_U3151), .ZN(P2_U3286) );
  INV_X1 U8142 ( .A(n6357), .ZN(n6358) );
  INV_X1 U8143 ( .A(n6788), .ZN(n6793) );
  OAI222_X1 U8144 ( .A1(n9969), .A2(n6358), .B1(n6793), .B2(P1_U3086), .C1(
        n9869), .C2(n9966), .ZN(P1_U3345) );
  INV_X1 U8145 ( .A(n7244), .ZN(n7366) );
  OAI222_X1 U8146 ( .A1(n8258), .A2(n6359), .B1(n7567), .B2(n6358), .C1(n7366), 
        .C2(P2_U3151), .ZN(P2_U3285) );
  NAND2_X1 U8147 ( .A1(n6620), .A2(n7311), .ZN(n6360) );
  NAND2_X1 U8148 ( .A1(n6361), .A2(n6360), .ZN(n6370) );
  INV_X1 U8149 ( .A(n6370), .ZN(n6363) );
  INV_X1 U8150 ( .A(n7311), .ZN(n6362) );
  OAI21_X1 U8151 ( .B1(n6614), .B2(n6362), .A(P1_STATE_REG_SCAN_IN), .ZN(n6369) );
  NOR2_X2 U8152 ( .A1(n6363), .A2(n6369), .ZN(n10043) );
  NOR2_X1 U8153 ( .A1(n10043), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8154 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n9875) );
  NOR2_X1 U8155 ( .A1(n6573), .A2(n9875), .ZN(P2_U3247) );
  INV_X1 U8156 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n6365) );
  NOR2_X1 U8157 ( .A1(n6573), .A2(n6365), .ZN(P2_U3258) );
  INV_X1 U8158 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n6366) );
  NOR2_X1 U8159 ( .A1(n6573), .A2(n6366), .ZN(P2_U3261) );
  INV_X1 U8160 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n6367) );
  NOR2_X1 U8161 ( .A1(n6573), .A2(n6367), .ZN(P2_U3260) );
  INV_X1 U8162 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n6368) );
  NOR2_X1 U8163 ( .A1(n6573), .A2(n6368), .ZN(P2_U3259) );
  OR2_X1 U8164 ( .A1(n6370), .A2(n6369), .ZN(n10041) );
  INV_X1 U8165 ( .A(n9255), .ZN(n6377) );
  INV_X1 U8166 ( .A(n6381), .ZN(n9235) );
  NAND2_X1 U8167 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9243) );
  AOI21_X1 U8168 ( .B1(P1_REG2_REG_1__SCAN_IN), .B2(n9235), .A(n9232), .ZN(
        n9250) );
  XOR2_X1 U8169 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n9255), .Z(n9249) );
  NOR2_X1 U8170 ( .A1(n9250), .A2(n9249), .ZN(n9248) );
  AOI21_X1 U8171 ( .B1(P1_REG2_REG_2__SCAN_IN), .B2(n6377), .A(n9248), .ZN(
        n6375) );
  XNOR2_X1 U8172 ( .A(n6399), .B(n7024), .ZN(n6374) );
  NOR2_X1 U8173 ( .A1(n6375), .A2(n6374), .ZN(n6400) );
  OR2_X1 U8174 ( .A1(n6372), .A2(n9246), .ZN(n6373) );
  AOI211_X1 U8175 ( .C1(n6375), .C2(n6374), .A(n6400), .B(n10044), .ZN(n6387)
         );
  MUX2_X1 U8176 ( .A(n6376), .B(P1_REG1_REG_3__SCAN_IN), .S(n6399), .Z(n6379)
         );
  NAND2_X1 U8177 ( .A1(n6377), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6384) );
  INV_X1 U8178 ( .A(n6384), .ZN(n6378) );
  NOR2_X1 U8179 ( .A1(n6379), .A2(n6378), .ZN(n6385) );
  MUX2_X1 U8180 ( .A(n6380), .B(P1_REG1_REG_2__SCAN_IN), .S(n9255), .Z(n9253)
         );
  XNOR2_X1 U8181 ( .A(n6381), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n9238) );
  AND2_X1 U8182 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9237) );
  NAND2_X1 U8183 ( .A1(n9238), .A2(n9237), .ZN(n9236) );
  NAND2_X1 U8184 ( .A1(n9235), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6382) );
  NAND2_X1 U8185 ( .A1(n9236), .A2(n6382), .ZN(n9252) );
  NAND2_X1 U8186 ( .A1(n9253), .A2(n9252), .ZN(n9251) );
  MUX2_X1 U8187 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6376), .S(n6399), .Z(n6383)
         );
  AOI21_X1 U8188 ( .B1(n9251), .B2(n6384), .A(n6383), .ZN(n6405) );
  INV_X1 U8189 ( .A(n6372), .ZN(n10031) );
  AOI211_X1 U8190 ( .C1(n6385), .C2(n9251), .A(n6405), .B(n9336), .ZN(n6386)
         );
  NOR2_X1 U8191 ( .A1(n6387), .A2(n6386), .ZN(n6391) );
  INV_X1 U8192 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6388) );
  NOR2_X1 U8193 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6388), .ZN(n6389) );
  AOI21_X1 U8194 ( .B1(n10043), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n6389), .ZN(
        n6390) );
  OAI211_X1 U8195 ( .C1(n6399), .C2(n9335), .A(n6391), .B(n6390), .ZN(P1_U3246) );
  INV_X1 U8196 ( .A(n6392), .ZN(n6394) );
  INV_X1 U8197 ( .A(n6872), .ZN(n6868) );
  OAI222_X1 U8198 ( .A1(n9966), .A2(n6393), .B1(n9969), .B2(n6394), .C1(
        P1_U3086), .C2(n6868), .ZN(P1_U3344) );
  INV_X1 U8199 ( .A(n7424), .ZN(n7418) );
  OAI222_X1 U8200 ( .A1(n8258), .A2(n6395), .B1(n7567), .B2(n6394), .C1(
        P2_U3151), .C2(n7418), .ZN(P2_U3284) );
  OAI22_X1 U8201 ( .A1(n6573), .A2(P2_D_REG_0__SCAN_IN), .B1(n6397), .B2(n6396), .ZN(n6398) );
  INV_X1 U8202 ( .A(n6398), .ZN(P2_U3376) );
  INV_X1 U8203 ( .A(n6399), .ZN(n6406) );
  NAND2_X1 U8204 ( .A1(n10051), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6401) );
  OAI21_X1 U8205 ( .B1(n10051), .B2(P1_REG2_REG_4__SCAN_IN), .A(n6401), .ZN(
        n10046) );
  NAND2_X1 U8206 ( .A1(n6423), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6402) );
  OAI21_X1 U8207 ( .B1(n6423), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6402), .ZN(
        n6403) );
  AOI211_X1 U8208 ( .C1(n6404), .C2(n6403), .A(n6418), .B(n10044), .ZN(n6417)
         );
  NAND2_X1 U8209 ( .A1(n10051), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6407) );
  AOI21_X1 U8210 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(n6406), .A(n6405), .ZN(
        n10054) );
  MUX2_X1 U8211 ( .A(n5812), .B(P1_REG1_REG_4__SCAN_IN), .S(n10051), .Z(n10053) );
  OR2_X1 U8212 ( .A1(n10054), .A2(n10053), .ZN(n10056) );
  NAND2_X1 U8213 ( .A1(n6407), .A2(n10056), .ZN(n6410) );
  MUX2_X1 U8214 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6408), .S(n6423), .Z(n6409)
         );
  NAND2_X1 U8215 ( .A1(n6409), .A2(n6410), .ZN(n6424) );
  OAI211_X1 U8216 ( .C1(n6410), .C2(n6409), .A(n10057), .B(n6424), .ZN(n6414)
         );
  NOR2_X1 U8217 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6411), .ZN(n6412) );
  AOI21_X1 U8218 ( .B1(n10043), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n6412), .ZN(
        n6413) );
  OAI211_X1 U8219 ( .C1(n9335), .C2(n6415), .A(n6414), .B(n6413), .ZN(n6416)
         );
  OR2_X1 U8220 ( .A1(n6417), .A2(n6416), .ZN(P1_U3248) );
  AOI21_X1 U8221 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n6423), .A(n6418), .ZN(
        n6461) );
  NAND2_X1 U8222 ( .A1(P1_REG2_REG_6__SCAN_IN), .A2(n6464), .ZN(n6419) );
  OAI21_X1 U8223 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n6464), .A(n6419), .ZN(
        n6460) );
  NOR2_X1 U8224 ( .A1(n6461), .A2(n6460), .ZN(n6459) );
  AOI21_X1 U8225 ( .B1(n6464), .B2(P1_REG2_REG_6__SCAN_IN), .A(n6459), .ZN(
        n6421) );
  AOI22_X1 U8226 ( .A1(n6437), .A2(n7042), .B1(P1_REG2_REG_7__SCAN_IN), .B2(
        n6441), .ZN(n6420) );
  NOR2_X1 U8227 ( .A1(n6421), .A2(n6420), .ZN(n6436) );
  AOI211_X1 U8228 ( .C1(n6421), .C2(n6420), .A(n6436), .B(n10044), .ZN(n6435)
         );
  NAND2_X1 U8229 ( .A1(P1_REG1_REG_6__SCAN_IN), .A2(n6464), .ZN(n6426) );
  MUX2_X1 U8230 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6422), .S(n6464), .Z(n6455)
         );
  NAND2_X1 U8231 ( .A1(n6423), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6425) );
  NAND2_X1 U8232 ( .A1(n6425), .A2(n6424), .ZN(n6456) );
  NAND2_X1 U8233 ( .A1(n6455), .A2(n6456), .ZN(n6454) );
  NAND2_X1 U8234 ( .A1(n6426), .A2(n6454), .ZN(n6429) );
  MUX2_X1 U8235 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n6427), .S(n6437), .Z(n6428)
         );
  NAND2_X1 U8236 ( .A1(n6428), .A2(n6429), .ZN(n6440) );
  OAI211_X1 U8237 ( .C1(n6429), .C2(n6428), .A(n10057), .B(n6440), .ZN(n6433)
         );
  NOR2_X1 U8238 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6430), .ZN(n6431) );
  AOI21_X1 U8239 ( .B1(n10043), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n6431), .ZN(
        n6432) );
  OAI211_X1 U8240 ( .C1(n9335), .C2(n6441), .A(n6433), .B(n6432), .ZN(n6434)
         );
  OR2_X1 U8241 ( .A1(n6435), .A2(n6434), .ZN(P1_U3250) );
  AOI22_X1 U8242 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n6467), .B1(n6472), .B2(
        n9561), .ZN(n6438) );
  AOI211_X1 U8243 ( .C1(n6439), .C2(n6438), .A(n6471), .B(n10044), .ZN(n6449)
         );
  OAI21_X1 U8244 ( .B1(n6441), .B2(n6427), .A(n6440), .ZN(n6444) );
  MUX2_X1 U8245 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n6442), .S(n6472), .Z(n6443)
         );
  NAND2_X1 U8246 ( .A1(n6443), .A2(n6444), .ZN(n6466) );
  OAI211_X1 U8247 ( .C1(n6444), .C2(n6443), .A(n10057), .B(n6466), .ZN(n6447)
         );
  NOR2_X1 U8248 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5867), .ZN(n6445) );
  AOI21_X1 U8249 ( .B1(n10043), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n6445), .ZN(
        n6446) );
  OAI211_X1 U8250 ( .C1(n9335), .C2(n6467), .A(n6447), .B(n6446), .ZN(n6448)
         );
  OR2_X1 U8251 ( .A1(n6449), .A2(n6448), .ZN(P1_U3251) );
  INV_X1 U8252 ( .A(n6450), .ZN(n6452) );
  INV_X1 U8253 ( .A(n7079), .ZN(n6877) );
  OAI222_X1 U8254 ( .A1(n9969), .A2(n6452), .B1(n6877), .B2(P1_U3086), .C1(
        n6451), .C2(n9966), .ZN(P1_U3343) );
  INV_X1 U8255 ( .A(n7427), .ZN(n8428) );
  OAI222_X1 U8256 ( .A1(n8258), .A2(n6453), .B1(n7567), .B2(n6452), .C1(n8428), 
        .C2(P2_U3151), .ZN(P2_U3283) );
  INV_X1 U8257 ( .A(n9335), .ZN(n10052) );
  INV_X1 U8258 ( .A(n10043), .ZN(n9347) );
  INV_X1 U8259 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6458) );
  OAI211_X1 U8260 ( .C1(n6456), .C2(n6455), .A(n10057), .B(n6454), .ZN(n6457)
         );
  NAND2_X1 U8261 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7099) );
  OAI211_X1 U8262 ( .C1(n9347), .C2(n6458), .A(n6457), .B(n7099), .ZN(n6463)
         );
  AOI211_X1 U8263 ( .C1(n6461), .C2(n6460), .A(n6459), .B(n10044), .ZN(n6462)
         );
  AOI211_X1 U8264 ( .C1(n10052), .C2(n6464), .A(n6463), .B(n6462), .ZN(n6465)
         );
  INV_X1 U8265 ( .A(n6465), .ZN(P1_U3249) );
  OAI21_X1 U8266 ( .B1(n6467), .B2(n6442), .A(n6466), .ZN(n6470) );
  MUX2_X1 U8267 ( .A(n6468), .B(P1_REG1_REG_9__SCAN_IN), .S(n6671), .Z(n6469)
         );
  NOR2_X1 U8268 ( .A1(n6469), .A2(n6470), .ZN(n6674) );
  AOI21_X1 U8269 ( .B1(n6470), .B2(n6469), .A(n6674), .ZN(n6480) );
  MUX2_X1 U8270 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n7254), .S(n6671), .Z(n6473)
         );
  OAI21_X1 U8271 ( .B1(n6474), .B2(n6473), .A(n6670), .ZN(n6475) );
  INV_X1 U8272 ( .A(n10044), .ZN(n9340) );
  NAND2_X1 U8273 ( .A1(n6475), .A2(n9340), .ZN(n6479) );
  INV_X1 U8274 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n6476) );
  NAND2_X1 U8275 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7451) );
  OAI21_X1 U8276 ( .B1(n9347), .B2(n6476), .A(n7451), .ZN(n6477) );
  AOI21_X1 U8277 ( .B1(n6671), .B2(n10052), .A(n6477), .ZN(n6478) );
  OAI211_X1 U8278 ( .C1(n6480), .C2(n9336), .A(n6479), .B(n6478), .ZN(P1_U3252) );
  INV_X2 U8279 ( .A(P1_U3973), .ZN(n9231) );
  NAND2_X1 U8280 ( .A1(n9231), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n6481) );
  OAI21_X1 U8281 ( .B1(n7626), .B2(n9231), .A(n6481), .ZN(P1_U3568) );
  NAND2_X1 U8282 ( .A1(n9231), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6482) );
  OAI21_X1 U8283 ( .B1(n9161), .B2(n9231), .A(n6482), .ZN(P1_U3577) );
  AND2_X1 U8284 ( .A1(n9230), .A2(n9150), .ZN(n7012) );
  AND2_X1 U8285 ( .A1(n6109), .A2(n10095), .ZN(n7755) );
  NOR2_X1 U8286 ( .A1(n10086), .A2(n7755), .ZN(n7955) );
  AOI21_X1 U8287 ( .B1(n9639), .B2(n10087), .A(n7955), .ZN(n6483) );
  AOI211_X1 U8288 ( .C1(n6484), .C2(n6626), .A(n7012), .B(n6483), .ZN(n6487)
         );
  NAND2_X1 U8289 ( .A1(n10173), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6485) );
  OAI21_X1 U8290 ( .B1(n6487), .B2(n10173), .A(n6485), .ZN(P1_U3453) );
  NAND2_X1 U8291 ( .A1(n10184), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6486) );
  OAI21_X1 U8292 ( .B1(n6487), .B2(n10184), .A(n6486), .ZN(P1_U3522) );
  NOR2_X1 U8293 ( .A1(n8551), .A2(P2_U3151), .ZN(n7565) );
  NAND2_X1 U8294 ( .A1(n7565), .A2(n6513), .ZN(n6489) );
  MUX2_X1 U8295 ( .A(n8527), .B(n6489), .S(n8026), .Z(n10204) );
  MUX2_X1 U8296 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8551), .Z(n6495) );
  INV_X1 U8297 ( .A(n6495), .ZN(n6496) );
  MUX2_X1 U8298 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8551), .Z(n6493) );
  INV_X1 U8299 ( .A(n6493), .ZN(n6494) );
  INV_X1 U8300 ( .A(n10203), .ZN(n6492) );
  MUX2_X1 U8301 ( .A(n6849), .B(n6490), .S(n8551), .Z(n6491) );
  XNOR2_X1 U8302 ( .A(n6491), .B(n10203), .ZN(n10200) );
  MUX2_X1 U8303 ( .A(n6717), .B(n6515), .S(n8551), .Z(n10187) );
  NAND2_X1 U8304 ( .A1(n10187), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n10199) );
  NAND2_X1 U8305 ( .A1(n10200), .A2(n10199), .ZN(n10198) );
  OAI21_X1 U8306 ( .B1(n6492), .B2(n6491), .A(n10198), .ZN(n6550) );
  XNOR2_X1 U8307 ( .A(n6493), .B(n6519), .ZN(n6549) );
  NAND2_X1 U8308 ( .A1(n6550), .A2(n6549), .ZN(n6548) );
  OAI21_X1 U8309 ( .B1(n6519), .B2(n6494), .A(n6548), .ZN(n6554) );
  XOR2_X1 U8310 ( .A(n6567), .B(n6495), .Z(n6555) );
  NOR2_X1 U8311 ( .A1(n6554), .A2(n6555), .ZN(n6553) );
  AOI21_X1 U8312 ( .B1(n6567), .B2(n6496), .A(n6553), .ZN(n6499) );
  MUX2_X1 U8313 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8551), .Z(n6646) );
  XNOR2_X1 U8314 ( .A(n6646), .B(n6657), .ZN(n6498) );
  NAND2_X1 U8315 ( .A1(n6499), .A2(n6498), .ZN(n6647) );
  NOR2_X2 U8316 ( .A1(n8527), .A2(n6497), .ZN(n10225) );
  OAI211_X1 U8317 ( .C1(n6499), .C2(n6498), .A(n6647), .B(n10225), .ZN(n6533)
         );
  NOR2_X1 U8318 ( .A1(n6501), .A2(n6500), .ZN(n6502) );
  MUX2_X1 U8319 ( .A(n6505), .B(P2_REG2_REG_2__SCAN_IN), .S(n6519), .Z(n6538)
         );
  NOR2_X1 U8320 ( .A1(n6717), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6503) );
  NAND2_X1 U8321 ( .A1(n6516), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6504) );
  OR2_X1 U8322 ( .A1(n10208), .A2(n6849), .ZN(n10206) );
  NAND2_X1 U8323 ( .A1(n10206), .A2(n6504), .ZN(n6537) );
  NAND2_X1 U8324 ( .A1(n6538), .A2(n6537), .ZN(n6536) );
  OR2_X1 U8325 ( .A1(n6519), .A2(n6505), .ZN(n6506) );
  NAND2_X1 U8326 ( .A1(n6536), .A2(n6506), .ZN(n6507) );
  NAND2_X1 U8327 ( .A1(n6507), .A2(n6521), .ZN(n6510) );
  OR2_X1 U8328 ( .A1(n6507), .A2(n6521), .ZN(n6508) );
  MUX2_X1 U8329 ( .A(n6651), .B(P2_REG2_REG_4__SCAN_IN), .S(n6657), .Z(n6509)
         );
  INV_X1 U8330 ( .A(n6509), .ZN(n6511) );
  NAND3_X1 U8331 ( .A1(n6558), .A2(n6511), .A3(n6510), .ZN(n6512) );
  AND2_X1 U8332 ( .A1(n6653), .A2(n6512), .ZN(n6530) );
  NOR2_X1 U8333 ( .A1(n8026), .A2(P2_U3151), .ZN(n7604) );
  AND2_X1 U8334 ( .A1(n6513), .A2(n7604), .ZN(n10189) );
  INV_X1 U8335 ( .A(n10189), .ZN(n6514) );
  INV_X1 U8336 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10289) );
  NOR2_X1 U8337 ( .A1(n6515), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6517) );
  NAND2_X1 U8338 ( .A1(n6516), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6518) );
  OAI21_X1 U8339 ( .B1(n10203), .B2(n6517), .A(n6518), .ZN(n10193) );
  OR2_X1 U8340 ( .A1(n10193), .A2(n6490), .ZN(n10194) );
  NAND2_X1 U8341 ( .A1(n10194), .A2(n6518), .ZN(n6541) );
  OR2_X1 U8342 ( .A1(n6519), .A2(n10289), .ZN(n6520) );
  NAND2_X1 U8343 ( .A1(n6522), .A2(n6521), .ZN(n6526) );
  NAND2_X1 U8344 ( .A1(n6526), .A2(n6523), .ZN(n6560) );
  INV_X1 U8345 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10291) );
  INV_X1 U8346 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6524) );
  MUX2_X1 U8347 ( .A(n6524), .B(P2_REG1_REG_4__SCAN_IN), .S(n6657), .Z(n6525)
         );
  NAND3_X1 U8348 ( .A1(n6562), .A2(n4836), .A3(n6526), .ZN(n6527) );
  NAND2_X1 U8349 ( .A1(n6658), .A2(n6527), .ZN(n6528) );
  NAND2_X1 U8350 ( .A1(n10197), .A2(n6528), .ZN(n6529) );
  NAND2_X1 U8351 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n6831) );
  OAI211_X1 U8352 ( .C1(n6530), .C2(n10220), .A(n6529), .B(n6831), .ZN(n6531)
         );
  AOI21_X1 U8353 ( .B1(n10212), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n6531), .ZN(
        n6532) );
  OAI211_X1 U8354 ( .C1(n10204), .C2(n6534), .A(n6533), .B(n6532), .ZN(
        P2_U3186) );
  NOR2_X1 U8355 ( .A1(n10204), .A2(n6535), .ZN(n6547) );
  INV_X1 U8356 ( .A(n10220), .ZN(n7368) );
  OAI21_X1 U8357 ( .B1(n6538), .B2(n6537), .A(n6536), .ZN(n6539) );
  NAND2_X1 U8358 ( .A1(n7368), .A2(n6539), .ZN(n6545) );
  OAI21_X1 U8359 ( .B1(n6542), .B2(n6541), .A(n6540), .ZN(n6543) );
  NAND2_X1 U8360 ( .A1(n10197), .A2(n6543), .ZN(n6544) );
  OAI211_X1 U8361 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n6728), .A(n6545), .B(n6544), .ZN(n6546) );
  AOI211_X1 U8362 ( .C1(n10212), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n6547), .B(
        n6546), .ZN(n6552) );
  OAI211_X1 U8363 ( .C1(n6550), .C2(n6549), .A(n6548), .B(n10225), .ZN(n6551)
         );
  NAND2_X1 U8364 ( .A1(n6552), .A2(n6551), .ZN(P2_U3184) );
  AOI21_X1 U8365 ( .B1(n6555), .B2(n6554), .A(n6553), .ZN(n6569) );
  INV_X1 U8366 ( .A(n10225), .ZN(n6928) );
  INV_X1 U8367 ( .A(n10204), .ZN(n10213) );
  INV_X1 U8368 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n9975) );
  NAND2_X1 U8369 ( .A1(n6556), .A2(n6859), .ZN(n6557) );
  NAND2_X1 U8370 ( .A1(n6558), .A2(n6557), .ZN(n6559) );
  AOI22_X1 U8371 ( .A1(n7368), .A2(n6559), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        P2_U3151), .ZN(n6565) );
  NAND2_X1 U8372 ( .A1(n6560), .A2(n10291), .ZN(n6561) );
  NAND2_X1 U8373 ( .A1(n6562), .A2(n6561), .ZN(n6563) );
  NAND2_X1 U8374 ( .A1(n10197), .A2(n6563), .ZN(n6564) );
  OAI211_X1 U8375 ( .C1(n9975), .C2(n10192), .A(n6565), .B(n6564), .ZN(n6566)
         );
  AOI21_X1 U8376 ( .B1(n6567), .B2(n10213), .A(n6566), .ZN(n6568) );
  OAI21_X1 U8377 ( .B1(n6569), .B2(n6928), .A(n6568), .ZN(P2_U3185) );
  INV_X1 U8378 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n9893) );
  INV_X1 U8379 ( .A(n6570), .ZN(n6571) );
  OAI222_X1 U8380 ( .A1(n8258), .A2(n9893), .B1(n7567), .B2(n6571), .C1(
        P2_U3151), .C2(n4639), .ZN(P2_U3282) );
  INV_X1 U8381 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6572) );
  INV_X1 U8382 ( .A(n7262), .ZN(n7269) );
  OAI222_X1 U8383 ( .A1(n9966), .A2(n6572), .B1(n9969), .B2(n6571), .C1(
        P1_U3086), .C2(n7269), .ZN(P1_U3342) );
  INV_X1 U8384 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n6574) );
  NOR2_X1 U8385 ( .A1(n6594), .A2(n6574), .ZN(P2_U3234) );
  INV_X1 U8386 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n6575) );
  NOR2_X1 U8387 ( .A1(n6594), .A2(n6575), .ZN(P2_U3262) );
  INV_X1 U8388 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n6576) );
  NOR2_X1 U8389 ( .A1(n6594), .A2(n6576), .ZN(P2_U3256) );
  INV_X1 U8390 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n6577) );
  NOR2_X1 U8391 ( .A1(n6594), .A2(n6577), .ZN(P2_U3263) );
  INV_X1 U8392 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n6578) );
  NOR2_X1 U8393 ( .A1(n6594), .A2(n6578), .ZN(P2_U3254) );
  INV_X1 U8394 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n6579) );
  NOR2_X1 U8395 ( .A1(n6594), .A2(n6579), .ZN(P2_U3253) );
  INV_X1 U8396 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n9899) );
  NOR2_X1 U8397 ( .A1(n6594), .A2(n9899), .ZN(P2_U3252) );
  INV_X1 U8398 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n6580) );
  NOR2_X1 U8399 ( .A1(n6594), .A2(n6580), .ZN(P2_U3255) );
  INV_X1 U8400 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n9721) );
  NOR2_X1 U8401 ( .A1(n6594), .A2(n9721), .ZN(P2_U3250) );
  INV_X1 U8402 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n6581) );
  NOR2_X1 U8403 ( .A1(n6594), .A2(n6581), .ZN(P2_U3249) );
  INV_X1 U8404 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n6582) );
  NOR2_X1 U8405 ( .A1(n6594), .A2(n6582), .ZN(P2_U3248) );
  INV_X1 U8406 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n6583) );
  NOR2_X1 U8407 ( .A1(n6594), .A2(n6583), .ZN(P2_U3251) );
  INV_X1 U8408 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n6584) );
  NOR2_X1 U8409 ( .A1(n6594), .A2(n6584), .ZN(P2_U3246) );
  INV_X1 U8410 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n9723) );
  NOR2_X1 U8411 ( .A1(n6594), .A2(n9723), .ZN(P2_U3245) );
  INV_X1 U8412 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n9871) );
  NOR2_X1 U8413 ( .A1(n6594), .A2(n9871), .ZN(P2_U3243) );
  INV_X1 U8414 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n9897) );
  NOR2_X1 U8415 ( .A1(n6594), .A2(n9897), .ZN(P2_U3242) );
  INV_X1 U8416 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n6585) );
  NOR2_X1 U8417 ( .A1(n6594), .A2(n6585), .ZN(P2_U3241) );
  INV_X1 U8418 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n6586) );
  NOR2_X1 U8419 ( .A1(n6594), .A2(n6586), .ZN(P2_U3240) );
  INV_X1 U8420 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n6587) );
  NOR2_X1 U8421 ( .A1(n6594), .A2(n6587), .ZN(P2_U3239) );
  INV_X1 U8422 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n6588) );
  NOR2_X1 U8423 ( .A1(n6594), .A2(n6588), .ZN(P2_U3238) );
  INV_X1 U8424 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n6589) );
  NOR2_X1 U8425 ( .A1(n6594), .A2(n6589), .ZN(P2_U3237) );
  INV_X1 U8426 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n6590) );
  NOR2_X1 U8427 ( .A1(n6594), .A2(n6590), .ZN(P2_U3236) );
  INV_X1 U8428 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n6591) );
  NOR2_X1 U8429 ( .A1(n6594), .A2(n6591), .ZN(P2_U3235) );
  INV_X1 U8430 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n6592) );
  NOR2_X1 U8431 ( .A1(n6594), .A2(n6592), .ZN(P2_U3257) );
  INV_X1 U8432 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n6593) );
  NOR2_X1 U8433 ( .A1(n6594), .A2(n6593), .ZN(P2_U3244) );
  INV_X1 U8434 ( .A(n6595), .ZN(n6597) );
  OAI222_X1 U8435 ( .A1(n8258), .A2(n6596), .B1(n7567), .B2(n6597), .C1(
        P2_U3151), .C2(n8475), .ZN(P2_U3281) );
  INV_X1 U8436 ( .A(n9261), .ZN(n9264) );
  OAI222_X1 U8437 ( .A1(n9966), .A2(n6598), .B1(n9969), .B2(n6597), .C1(
        P1_U3086), .C2(n9264), .ZN(P1_U3341) );
  NOR2_X1 U8438 ( .A1(n6600), .A2(n6599), .ZN(n6601) );
  NAND2_X1 U8439 ( .A1(n6619), .A2(n6623), .ZN(n6605) );
  AND3_X1 U8440 ( .A1(n6614), .A2(n7311), .A3(n6603), .ZN(n6604) );
  NOR2_X1 U8441 ( .A1(n9145), .A2(P1_U3086), .ZN(n6706) );
  NAND2_X1 U8442 ( .A1(n7304), .A2(n8012), .ZN(n6606) );
  NAND2_X1 U8443 ( .A1(n7757), .A2(n7108), .ZN(n6608) );
  OR2_X1 U8444 ( .A1(n6608), .A2(n9342), .ZN(n10092) );
  INV_X1 U8445 ( .A(n7551), .ZN(n9002) );
  NAND2_X1 U8446 ( .A1(n6109), .A2(n9002), .ZN(n6612) );
  INV_X1 U8447 ( .A(n6608), .ZN(n6609) );
  AND2_X2 U8448 ( .A1(n6614), .A2(n6609), .ZN(n7541) );
  INV_X1 U8449 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10034) );
  NOR2_X1 U8450 ( .A1(n6614), .A2(n10034), .ZN(n6610) );
  AOI21_X1 U8451 ( .B1(n6626), .B2(n7541), .A(n6610), .ZN(n6611) );
  NAND2_X1 U8452 ( .A1(n6612), .A2(n6611), .ZN(n6637) );
  INV_X1 U8453 ( .A(n6637), .ZN(n6617) );
  NAND2_X1 U8454 ( .A1(n6109), .A2(n7541), .ZN(n6615) );
  NAND2_X4 U8455 ( .A1(n6614), .A2(n6613), .ZN(n8997) );
  INV_X2 U8456 ( .A(n8996), .ZN(n9070) );
  NAND2_X1 U8457 ( .A1(n6626), .A2(n9070), .ZN(n6636) );
  OAI211_X1 U8458 ( .C1(n6616), .C2(n6614), .A(n6615), .B(n6636), .ZN(n6638)
         );
  XNOR2_X1 U8459 ( .A(n6617), .B(n6638), .ZN(n9244) );
  INV_X1 U8460 ( .A(n8013), .ZN(n6618) );
  NOR2_X1 U8461 ( .A1(n10165), .A2(n6620), .ZN(n6621) );
  NAND2_X1 U8462 ( .A1(n9244), .A2(n9184), .ZN(n6628) );
  NAND2_X1 U8463 ( .A1(n6622), .A2(n8012), .ZN(n9143) );
  NOR2_X1 U8464 ( .A1(n7009), .A2(n7108), .ZN(n6998) );
  NAND2_X1 U8465 ( .A1(n6622), .A2(n6998), .ZN(n6625) );
  INV_X1 U8466 ( .A(n6623), .ZN(n6624) );
  AOI22_X1 U8467 ( .A1(n9195), .A2(n7012), .B1(n9201), .B2(n6626), .ZN(n6627)
         );
  OAI211_X1 U8468 ( .C1(n6706), .C2(n6629), .A(n6628), .B(n6627), .ZN(P1_U3232) );
  NAND2_X1 U8469 ( .A1(n9230), .A2(n7541), .ZN(n6630) );
  NAND2_X1 U8470 ( .A1(n9230), .A2(n9002), .ZN(n6632) );
  OR2_X1 U8471 ( .A1(n6106), .A2(n4394), .ZN(n6631) );
  NAND2_X1 U8472 ( .A1(n6632), .A2(n6631), .ZN(n6633) );
  AOI22_X1 U8473 ( .A1(n6638), .A2(n6637), .B1(n9068), .B2(n6636), .ZN(n6639)
         );
  NOR2_X1 U8474 ( .A1(n6640), .A2(n6639), .ZN(n6641) );
  OAI21_X1 U8475 ( .B1(n6641), .B2(n6699), .A(n9184), .ZN(n6644) );
  INV_X1 U8476 ( .A(n6109), .ZN(n6642) );
  OAI22_X1 U8477 ( .A1(n6693), .A2(n9350), .B1(n6642), .B2(n9373), .ZN(n10090)
         );
  AOI22_X1 U8478 ( .A1(n10090), .A2(n9195), .B1(n5773), .B2(n9201), .ZN(n6643)
         );
  OAI211_X1 U8479 ( .C1(n6706), .C2(n6645), .A(n6644), .B(n6643), .ZN(P1_U3222) );
  INV_X1 U8480 ( .A(n6646), .ZN(n6648) );
  OAI21_X1 U8481 ( .B1(n6657), .B2(n6648), .A(n6647), .ZN(n6650) );
  MUX2_X1 U8482 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8551), .Z(n6740) );
  XNOR2_X1 U8483 ( .A(n6740), .B(n6743), .ZN(n6649) );
  NAND2_X1 U8484 ( .A1(n6650), .A2(n6649), .ZN(n6741) );
  OAI211_X1 U8485 ( .C1(n6650), .C2(n6649), .A(n6741), .B(n10225), .ZN(n6667)
         );
  OR2_X1 U8486 ( .A1(n6657), .A2(n6651), .ZN(n6652) );
  NAND2_X1 U8487 ( .A1(n6653), .A2(n6652), .ZN(n6654) );
  NAND2_X1 U8488 ( .A1(n6654), .A2(n6668), .ZN(n6748) );
  OAI21_X1 U8489 ( .B1(n6654), .B2(n6668), .A(n6748), .ZN(n6655) );
  OR2_X1 U8490 ( .A1(n6655), .A2(n5247), .ZN(n6750) );
  NAND2_X1 U8491 ( .A1(n6655), .A2(n5247), .ZN(n6656) );
  AND2_X1 U8492 ( .A1(n6750), .A2(n6656), .ZN(n6664) );
  NAND2_X1 U8493 ( .A1(n6659), .A2(n6668), .ZN(n6755) );
  OAI21_X1 U8494 ( .B1(n6659), .B2(n6668), .A(n6755), .ZN(n6660) );
  NAND2_X1 U8495 ( .A1(n6660), .A2(n5246), .ZN(n6661) );
  NAND2_X1 U8496 ( .A1(n6757), .A2(n6661), .ZN(n6662) );
  NAND2_X1 U8497 ( .A1(n10197), .A2(n6662), .ZN(n6663) );
  NAND2_X1 U8498 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6889) );
  OAI211_X1 U8499 ( .C1(n6664), .C2(n10220), .A(n6663), .B(n6889), .ZN(n6665)
         );
  AOI21_X1 U8500 ( .B1(n10212), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6665), .ZN(
        n6666) );
  OAI211_X1 U8501 ( .C1(n10204), .C2(n6668), .A(n6667), .B(n6666), .ZN(
        P2_U3187) );
  NAND2_X1 U8502 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n6788), .ZN(n6669) );
  OAI21_X1 U8503 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n6788), .A(n6669), .ZN(
        n6673) );
  OAI21_X1 U8504 ( .B1(n6671), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6670), .ZN(
        n6672) );
  NOR2_X1 U8505 ( .A1(n6673), .A2(n6672), .ZN(n6787) );
  AOI211_X1 U8506 ( .C1(n6673), .C2(n6672), .A(n6787), .B(n10044), .ZN(n6683)
         );
  AOI21_X1 U8507 ( .B1(n6468), .B2(n6675), .A(n6674), .ZN(n6678) );
  MUX2_X1 U8508 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6676), .S(n6788), .Z(n6677)
         );
  NAND2_X1 U8509 ( .A1(n6678), .A2(n6677), .ZN(n6792) );
  OAI211_X1 U8510 ( .C1(n6678), .C2(n6677), .A(n10057), .B(n6792), .ZN(n6681)
         );
  AND2_X1 U8511 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6679) );
  AOI21_X1 U8512 ( .B1(n10043), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n6679), .ZN(
        n6680) );
  OAI211_X1 U8513 ( .C1(n9335), .C2(n6793), .A(n6681), .B(n6680), .ZN(n6682)
         );
  OR2_X1 U8514 ( .A1(n6683), .A2(n6682), .ZN(P1_U3253) );
  INV_X1 U8515 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6689) );
  NOR2_X1 U8516 ( .A1(n6844), .A2(n6684), .ZN(n8034) );
  INV_X1 U8517 ( .A(n8034), .ZN(n8036) );
  AND2_X1 U8518 ( .A1(n8036), .A2(n8035), .ZN(n8215) );
  INV_X1 U8519 ( .A(n8215), .ZN(n6685) );
  OAI21_X1 U8520 ( .B1(n8765), .B2(n10279), .A(n6685), .ZN(n6687) );
  NOR2_X1 U8521 ( .A1(n6187), .A2(n8762), .ZN(n6715) );
  INV_X1 U8522 ( .A(n6715), .ZN(n6686) );
  OAI211_X1 U8523 ( .C1(n10274), .C2(n6719), .A(n6687), .B(n6686), .ZN(n8830)
         );
  NAND2_X1 U8524 ( .A1(n8830), .A2(n10286), .ZN(n6688) );
  OAI21_X1 U8525 ( .B1(n6689), .B2(n10286), .A(n6688), .ZN(P2_U3390) );
  INV_X1 U8526 ( .A(n6690), .ZN(n6707) );
  AOI22_X1 U8527 ( .A1(n8499), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n8916), .ZN(n6691) );
  OAI21_X1 U8528 ( .B1(n6707), .B2(n8918), .A(n6691), .ZN(P2_U3280) );
  OAI22_X1 U8529 ( .A1(n6693), .A2(n4394), .B1(n5796), .B2(n8996), .ZN(n6692)
         );
  XNOR2_X1 U8530 ( .A(n6692), .B(n8997), .ZN(n6695) );
  OAI22_X1 U8531 ( .A1(n6693), .A2(n9065), .B1(n5796), .B2(n4394), .ZN(n6694)
         );
  OR2_X1 U8532 ( .A1(n6695), .A2(n6694), .ZN(n6768) );
  NAND2_X1 U8533 ( .A1(n6695), .A2(n6694), .ZN(n6696) );
  AND2_X1 U8534 ( .A1(n6768), .A2(n6696), .ZN(n6697) );
  INV_X1 U8535 ( .A(n6769), .ZN(n6701) );
  NOR3_X1 U8536 ( .A1(n6699), .A2(n6698), .A3(n6697), .ZN(n6700) );
  OAI21_X1 U8537 ( .B1(n6701), .B2(n6700), .A(n9184), .ZN(n6704) );
  OAI22_X1 U8538 ( .A1(n6781), .A2(n9350), .B1(n6702), .B2(n9373), .ZN(n10071)
         );
  AOI22_X1 U8539 ( .A1(n10071), .A2(n9195), .B1(n5795), .B2(n9201), .ZN(n6703)
         );
  OAI211_X1 U8540 ( .C1(n6706), .C2(n6705), .A(n6704), .B(n6703), .ZN(P1_U3237) );
  INV_X1 U8541 ( .A(n9273), .ZN(n9278) );
  OAI222_X1 U8542 ( .A1(n9969), .A2(n6707), .B1(n9278), .B2(P1_U3086), .C1(
        n9921), .C2(n9966), .ZN(P1_U3340) );
  AND2_X1 U8543 ( .A1(n6709), .A2(n6708), .ZN(n6735) );
  OAI22_X1 U8544 ( .A1(n8397), .A2(n6719), .B1(n8381), .B2(n8215), .ZN(n6710)
         );
  AOI21_X1 U8545 ( .B1(n8372), .B2(n8414), .A(n6710), .ZN(n6711) );
  OAI21_X1 U8546 ( .B1(n6735), .B2(n6712), .A(n6711), .ZN(P2_U3172) );
  INV_X1 U8547 ( .A(n8027), .ZN(n6713) );
  NOR3_X1 U8548 ( .A1(n8215), .A2(n6713), .A3(n10281), .ZN(n6714) );
  AOI211_X1 U8549 ( .C1(n8748), .C2(P2_REG3_REG_0__SCAN_IN), .A(n6715), .B(
        n6714), .ZN(n6716) );
  MUX2_X1 U8550 ( .A(n6717), .B(n6716), .S(n8745), .Z(n6718) );
  OAI21_X1 U8551 ( .B1(n8595), .B2(n6719), .A(n6718), .ZN(P2_U3233) );
  OAI22_X1 U8552 ( .A1(n8376), .A2(n6187), .B1(n8397), .B2(n6720), .ZN(n6721)
         );
  AOI21_X1 U8553 ( .B1(n8372), .B2(n8412), .A(n6721), .ZN(n6727) );
  OAI21_X1 U8554 ( .B1(n6724), .B2(n6723), .A(n6722), .ZN(n6725) );
  NAND2_X1 U8555 ( .A1(n6725), .A2(n8387), .ZN(n6726) );
  OAI211_X1 U8556 ( .C1(n6735), .C2(n6728), .A(n6727), .B(n6726), .ZN(P2_U3177) );
  INV_X1 U8557 ( .A(n6730), .ZN(n6731) );
  AOI21_X1 U8558 ( .B1(n6733), .B2(n6732), .A(n6731), .ZN(n6739) );
  NOR2_X1 U8559 ( .A1(n6735), .A2(n6734), .ZN(n6737) );
  OAI22_X1 U8560 ( .A1(n8376), .A2(n6844), .B1(n8397), .B2(n6186), .ZN(n6736)
         );
  AOI211_X1 U8561 ( .C1(n8372), .C2(n8413), .A(n6737), .B(n6736), .ZN(n6738)
         );
  OAI21_X1 U8562 ( .B1(n8381), .B2(n6739), .A(n6738), .ZN(P2_U3162) );
  MUX2_X1 U8563 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8551), .Z(n6910) );
  XOR2_X1 U8564 ( .A(n6913), .B(n6910), .Z(n6745) );
  INV_X1 U8565 ( .A(n6740), .ZN(n6742) );
  OAI21_X1 U8566 ( .B1(n6743), .B2(n6742), .A(n6741), .ZN(n6744) );
  NOR2_X1 U8567 ( .A1(n6744), .A2(n6745), .ZN(n6911) );
  AOI21_X1 U8568 ( .B1(n6745), .B2(n6744), .A(n6911), .ZN(n6763) );
  INV_X1 U8569 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n9987) );
  NAND2_X1 U8570 ( .A1(n6750), .A2(n6748), .ZN(n6746) );
  MUX2_X1 U8571 ( .A(n5262), .B(P2_REG2_REG_6__SCAN_IN), .S(n6913), .Z(n6747)
         );
  NAND2_X1 U8572 ( .A1(n6746), .A2(n6747), .ZN(n6919) );
  INV_X1 U8573 ( .A(n6747), .ZN(n6749) );
  NAND3_X1 U8574 ( .A1(n6750), .A2(n6749), .A3(n6748), .ZN(n6751) );
  AOI21_X1 U8575 ( .B1(n6919), .B2(n6751), .A(n10220), .ZN(n6753) );
  INV_X1 U8576 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6752) );
  NOR2_X1 U8577 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6752), .ZN(n7144) );
  NOR2_X1 U8578 ( .A1(n6753), .A2(n7144), .ZN(n6760) );
  INV_X1 U8579 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6754) );
  MUX2_X1 U8580 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6754), .S(n6913), .Z(n6756)
         );
  AND3_X1 U8581 ( .A1(n6757), .A2(n6756), .A3(n6755), .ZN(n6758) );
  OAI21_X1 U8582 ( .B1(n6914), .B2(n6758), .A(n10197), .ZN(n6759) );
  OAI211_X1 U8583 ( .C1(n9987), .C2(n10192), .A(n6760), .B(n6759), .ZN(n6761)
         );
  AOI21_X1 U8584 ( .B1(n6913), .B2(n10213), .A(n6761), .ZN(n6762) );
  OAI21_X1 U8585 ( .B1(n6763), .B2(n6928), .A(n6762), .ZN(P2_U3188) );
  NAND2_X1 U8586 ( .A1(n9231), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6764) );
  OAI21_X1 U8587 ( .B1(n9372), .B2(n9231), .A(n6764), .ZN(P1_U3582) );
  INV_X1 U8588 ( .A(n6765), .ZN(n6766) );
  INV_X1 U8589 ( .A(n8502), .ZN(n8533) );
  OAI222_X1 U8590 ( .A1(n8258), .A2(n9732), .B1(n7567), .B2(n6766), .C1(
        P2_U3151), .C2(n8533), .ZN(P2_U3279) );
  INV_X1 U8591 ( .A(n9294), .ZN(n9297) );
  OAI222_X1 U8592 ( .A1(n9966), .A2(n6767), .B1(n9969), .B2(n6766), .C1(
        P1_U3086), .C2(n9297), .ZN(P1_U3339) );
  OAI22_X1 U8593 ( .A1(n6781), .A2(n9065), .B1(n5810), .B2(n4394), .ZN(n6776)
         );
  OAI22_X1 U8594 ( .A1(n6781), .A2(n4394), .B1(n5810), .B2(n8996), .ZN(n6770)
         );
  XNOR2_X1 U8595 ( .A(n6770), .B(n8997), .ZN(n6775) );
  XOR2_X1 U8596 ( .A(n6776), .B(n6775), .Z(n6804) );
  NAND2_X2 U8597 ( .A1(n6803), .A2(n6804), .ZN(n6802) );
  NAND2_X1 U8598 ( .A1(n9228), .A2(n7541), .ZN(n6772) );
  NAND2_X1 U8599 ( .A1(n7136), .A2(n9070), .ZN(n6771) );
  NAND2_X1 U8600 ( .A1(n6772), .A2(n6771), .ZN(n6773) );
  XNOR2_X1 U8601 ( .A(n6773), .B(n8997), .ZN(n6942) );
  AND2_X1 U8602 ( .A1(n7136), .A2(n7541), .ZN(n6774) );
  AOI21_X1 U8603 ( .B1(n9228), .B2(n9002), .A(n6774), .ZN(n6940) );
  XNOR2_X1 U8604 ( .A(n6942), .B(n6940), .ZN(n6779) );
  INV_X1 U8605 ( .A(n6775), .ZN(n6778) );
  INV_X1 U8606 ( .A(n6776), .ZN(n6777) );
  NAND2_X1 U8607 ( .A1(n6778), .A2(n6777), .ZN(n6780) );
  NAND2_X1 U8608 ( .A1(n6946), .A2(n9184), .ZN(n6786) );
  AOI21_X1 U8609 ( .B1(n6802), .B2(n6780), .A(n6779), .ZN(n6785) );
  OAI22_X1 U8610 ( .A1(n6947), .A2(n9350), .B1(n6781), .B2(n9373), .ZN(n7127)
         );
  AOI22_X1 U8611 ( .A1(n7127), .A2(n9195), .B1(P1_REG3_REG_4__SCAN_IN), .B2(
        P1_U3086), .ZN(n6784) );
  INV_X1 U8612 ( .A(n7133), .ZN(n6782) );
  AOI22_X1 U8613 ( .A1(n9201), .A2(n7136), .B1(n9145), .B2(n6782), .ZN(n6783)
         );
  OAI211_X1 U8614 ( .C1(n6786), .C2(n6785), .A(n6784), .B(n6783), .ZN(P1_U3230) );
  NAND2_X1 U8615 ( .A1(n6872), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6789) );
  OAI21_X1 U8616 ( .B1(n6872), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6789), .ZN(
        n6790) );
  AOI211_X1 U8617 ( .C1(n6791), .C2(n6790), .A(n6871), .B(n10044), .ZN(n6801)
         );
  OAI21_X1 U8618 ( .B1(n6676), .B2(n6793), .A(n6792), .ZN(n6796) );
  MUX2_X1 U8619 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n6794), .S(n6872), .Z(n6795)
         );
  NAND2_X1 U8620 ( .A1(n6795), .A2(n6796), .ZN(n6867) );
  OAI211_X1 U8621 ( .C1(n6796), .C2(n6795), .A(n10057), .B(n6867), .ZN(n6799)
         );
  NOR2_X1 U8622 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6797), .ZN(n7657) );
  AOI21_X1 U8623 ( .B1(n10043), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n7657), .ZN(
        n6798) );
  OAI211_X1 U8624 ( .C1(n9335), .C2(n6868), .A(n6799), .B(n6798), .ZN(n6800)
         );
  OR2_X1 U8625 ( .A1(n6801), .A2(n6800), .ZN(P1_U3254) );
  OAI21_X1 U8626 ( .B1(n6804), .B2(n6803), .A(n6802), .ZN(n6808) );
  MUX2_X1 U8627 ( .A(n9145), .B(P1_U3086), .S(P1_REG3_REG_3__SCAN_IN), .Z(
        n6807) );
  INV_X1 U8628 ( .A(n9373), .ZN(n9173) );
  AOI22_X1 U8629 ( .A1(n6805), .A2(n9173), .B1(n9150), .B2(n9228), .ZN(n7022)
         );
  OAI22_X1 U8630 ( .A1(n7022), .A2(n9143), .B1(n5810), .B2(n9191), .ZN(n6806)
         );
  AOI211_X1 U8631 ( .C1(n6808), .C2(n9184), .A(n6807), .B(n6806), .ZN(n6809)
         );
  INV_X1 U8632 ( .A(n6809), .ZN(P1_U3218) );
  INV_X1 U8633 ( .A(n6811), .ZN(n6812) );
  AOI211_X1 U8634 ( .C1(n6813), .C2(n6810), .A(n8381), .B(n6812), .ZN(n6817)
         );
  MUX2_X1 U8635 ( .A(n8339), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n6815) );
  AOI22_X1 U8636 ( .A1(n8390), .A2(n8413), .B1(n8379), .B2(n6861), .ZN(n6814)
         );
  OAI211_X1 U8637 ( .C1(n6901), .C2(n8392), .A(n6815), .B(n6814), .ZN(n6816)
         );
  OR2_X1 U8638 ( .A1(n6817), .A2(n6816), .ZN(P2_U3158) );
  NAND3_X1 U8639 ( .A1(n6854), .A2(n6818), .A3(n8039), .ZN(n6819) );
  NAND2_X1 U8640 ( .A1(n6820), .A2(n6819), .ZN(n6977) );
  XNOR2_X1 U8641 ( .A(n6821), .B(n8213), .ZN(n6822) );
  OAI222_X1 U8642 ( .A1(n8762), .A2(n6823), .B1(n8761), .B2(n8763), .C1(n8629), 
        .C2(n6822), .ZN(n6974) );
  AOI21_X1 U8643 ( .B1(n10279), .B2(n6977), .A(n6974), .ZN(n6827) );
  OAI22_X1 U8644 ( .A1(n6973), .A2(n8842), .B1(n10286), .B2(n5233), .ZN(n6824)
         );
  INV_X1 U8645 ( .A(n6824), .ZN(n6825) );
  OAI21_X1 U8646 ( .B1(n6827), .B2(n10287), .A(n6825), .ZN(P2_U3402) );
  AOI22_X1 U8647 ( .A1(n8826), .A2(n6833), .B1(n6312), .B2(
        P2_REG1_REG_4__SCAN_IN), .ZN(n6826) );
  OAI21_X1 U8648 ( .B1(n6827), .B2(n6312), .A(n6826), .ZN(P2_U3463) );
  OAI21_X1 U8649 ( .B1(n6830), .B2(n6829), .A(n6828), .ZN(n6837) );
  AOI22_X1 U8650 ( .A1(n8372), .A2(n8410), .B1(n8390), .B2(n8412), .ZN(n6835)
         );
  INV_X1 U8651 ( .A(n6831), .ZN(n6832) );
  AOI21_X1 U8652 ( .B1(n8379), .B2(n6833), .A(n6832), .ZN(n6834) );
  OAI211_X1 U8653 ( .C1(n6972), .C2(n8339), .A(n6835), .B(n6834), .ZN(n6836)
         );
  AOI21_X1 U8654 ( .B1(n6837), .B2(n8387), .A(n6836), .ZN(n6838) );
  INV_X1 U8655 ( .A(n6838), .ZN(P2_U3170) );
  INV_X1 U8656 ( .A(n6840), .ZN(n6841) );
  AOI21_X1 U8657 ( .B1(n6839), .B2(n8035), .A(n6841), .ZN(n10236) );
  INV_X1 U8658 ( .A(n6842), .ZN(n8773) );
  NAND2_X1 U8659 ( .A1(n8745), .A2(n8773), .ZN(n7484) );
  OAI21_X1 U8660 ( .B1(n6843), .B2(n6839), .A(n8758), .ZN(n6848) );
  OAI22_X1 U8661 ( .A1(n6845), .A2(n8762), .B1(n6844), .B2(n8761), .ZN(n6847)
         );
  NOR2_X1 U8662 ( .A1(n10236), .A2(n7479), .ZN(n6846) );
  AOI211_X1 U8663 ( .C1(n8765), .C2(n6848), .A(n6847), .B(n6846), .ZN(n10235)
         );
  MUX2_X1 U8664 ( .A(n6849), .B(n10235), .S(n8745), .Z(n6852) );
  AOI22_X1 U8665 ( .A1(n8749), .A2(n6850), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8748), .ZN(n6851) );
  OAI211_X1 U8666 ( .C1(n10236), .C2(n7484), .A(n6852), .B(n6851), .ZN(
        P2_U3232) );
  INV_X1 U8667 ( .A(n6853), .ZN(n8041) );
  NOR2_X1 U8668 ( .A1(n8211), .A2(n8041), .ZN(n6856) );
  INV_X1 U8669 ( .A(n6854), .ZN(n6855) );
  AOI21_X1 U8670 ( .B1(n6856), .B2(n8753), .A(n6855), .ZN(n10248) );
  XOR2_X1 U8671 ( .A(n8211), .B(n6857), .Z(n6858) );
  AOI222_X1 U8672 ( .A1(n8765), .A2(n6858), .B1(n8411), .B2(n5047), .C1(n8413), 
        .C2(n8741), .ZN(n10245) );
  MUX2_X1 U8673 ( .A(n6859), .B(n10245), .S(n8745), .Z(n6863) );
  AOI22_X1 U8674 ( .A1(n8749), .A2(n6861), .B1(n8748), .B2(n6860), .ZN(n6862)
         );
  OAI211_X1 U8675 ( .C1(n10248), .C2(n8752), .A(n6863), .B(n6862), .ZN(
        P2_U3230) );
  INV_X1 U8676 ( .A(n6864), .ZN(n6882) );
  OAI222_X1 U8677 ( .A1(n8258), .A2(n6865), .B1(n7567), .B2(n6882), .C1(n8517), 
        .C2(P2_U3151), .ZN(P2_U3278) );
  NAND2_X1 U8678 ( .A1(n8527), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n6866) );
  OAI21_X1 U8679 ( .B1(n8169), .B2(n8527), .A(n6866), .ZN(P2_U3521) );
  OAI21_X1 U8680 ( .B1(n6794), .B2(n6868), .A(n6867), .ZN(n6870) );
  AOI22_X1 U8681 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n6877), .B1(n7079), .B2(
        n5930), .ZN(n6869) );
  NOR2_X1 U8682 ( .A1(n6870), .A2(n6869), .ZN(n7081) );
  AOI21_X1 U8683 ( .B1(n6870), .B2(n6869), .A(n7081), .ZN(n6881) );
  AOI22_X1 U8684 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7079), .B1(n6877), .B2(
        n5926), .ZN(n6874) );
  OAI21_X1 U8685 ( .B1(n6874), .B2(n6873), .A(n7076), .ZN(n6875) );
  NAND2_X1 U8686 ( .A1(n6875), .A2(n9340), .ZN(n6880) );
  NOR2_X1 U8687 ( .A1(n6876), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7556) );
  NOR2_X1 U8688 ( .A1(n9335), .A2(n6877), .ZN(n6878) );
  AOI211_X1 U8689 ( .C1(n10043), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n7556), .B(
        n6878), .ZN(n6879) );
  OAI211_X1 U8690 ( .C1(n6881), .C2(n9336), .A(n6880), .B(n6879), .ZN(P1_U3255) );
  INV_X1 U8691 ( .A(n9317), .ZN(n9303) );
  OAI222_X1 U8692 ( .A1(n9966), .A2(n6883), .B1(n9303), .B2(P1_U3086), .C1(
        n9969), .C2(n6882), .ZN(P1_U3338) );
  INV_X1 U8693 ( .A(n6884), .ZN(n6886) );
  NAND3_X1 U8694 ( .A1(n6828), .A2(n6886), .A3(n6885), .ZN(n6887) );
  AOI21_X1 U8695 ( .B1(n6888), .B2(n6887), .A(n8381), .ZN(n6894) );
  AOI22_X1 U8696 ( .A1(n8372), .A2(n8409), .B1(n8390), .B2(n8411), .ZN(n6892)
         );
  INV_X1 U8697 ( .A(n6889), .ZN(n6890) );
  AOI21_X1 U8698 ( .B1(n8379), .B2(n6902), .A(n6890), .ZN(n6891) );
  OAI211_X1 U8699 ( .C1(n8339), .C2(n6933), .A(n6892), .B(n6891), .ZN(n6893)
         );
  OR2_X1 U8700 ( .A1(n6894), .A2(n6893), .ZN(P2_U3167) );
  INV_X1 U8701 ( .A(n6895), .ZN(n6931) );
  AOI22_X1 U8702 ( .A1(n9330), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9962), .ZN(n6896) );
  OAI21_X1 U8703 ( .B1(n6931), .B2(n9969), .A(n6896), .ZN(P1_U3337) );
  OAI21_X1 U8704 ( .B1(n6898), .B2(n8214), .A(n6897), .ZN(n6937) );
  XNOR2_X1 U8705 ( .A(n6899), .B(n8214), .ZN(n6900) );
  OAI222_X1 U8706 ( .A1(n8762), .A2(n7207), .B1(n8761), .B2(n6901), .C1(n8629), 
        .C2(n6900), .ZN(n6932) );
  AOI21_X1 U8707 ( .B1(n10279), .B2(n6937), .A(n6932), .ZN(n6907) );
  AOI22_X1 U8708 ( .A1(n8826), .A2(n6902), .B1(n6312), .B2(
        P2_REG1_REG_5__SCAN_IN), .ZN(n6903) );
  OAI21_X1 U8709 ( .B1(n6907), .B2(n6312), .A(n6903), .ZN(P2_U3464) );
  INV_X1 U8710 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n6904) );
  OAI22_X1 U8711 ( .A1(n6934), .A2(n8842), .B1(n10286), .B2(n6904), .ZN(n6905)
         );
  INV_X1 U8712 ( .A(n6905), .ZN(n6906) );
  OAI21_X1 U8713 ( .B1(n6907), .B2(n10287), .A(n6906), .ZN(P2_U3405) );
  MUX2_X1 U8714 ( .A(n6909), .B(n6908), .S(n8551), .Z(n7047) );
  XNOR2_X1 U8715 ( .A(n7047), .B(n6915), .ZN(n7049) );
  INV_X1 U8716 ( .A(n6910), .ZN(n6912) );
  AOI21_X1 U8717 ( .B1(n6913), .B2(n6912), .A(n6911), .ZN(n7050) );
  XOR2_X1 U8718 ( .A(n7049), .B(n7050), .Z(n6929) );
  NAND2_X1 U8719 ( .A1(n6916), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7060) );
  OAI21_X1 U8720 ( .B1(n6916), .B2(P2_REG1_REG_7__SCAN_IN), .A(n7060), .ZN(
        n6926) );
  NAND2_X1 U8721 ( .A1(n6917), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6918) );
  NAND2_X1 U8722 ( .A1(n6919), .A2(n6918), .ZN(n6920) );
  NAND2_X1 U8723 ( .A1(n6921), .A2(n6909), .ZN(n6922) );
  AOI21_X1 U8724 ( .B1(n7055), .B2(n6922), .A(n10220), .ZN(n6925) );
  NAND2_X1 U8725 ( .A1(n10212), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n6923) );
  NAND2_X1 U8726 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7206) );
  OAI211_X1 U8727 ( .C1(n10204), .C2(n4853), .A(n6923), .B(n7206), .ZN(n6924)
         );
  AOI211_X1 U8728 ( .C1(n6926), .C2(n10197), .A(n6925), .B(n6924), .ZN(n6927)
         );
  OAI21_X1 U8729 ( .B1(n6929), .B2(n6928), .A(n6927), .ZN(P2_U3189) );
  INV_X1 U8730 ( .A(n8548), .ZN(n8536) );
  OAI222_X1 U8731 ( .A1(P2_U3151), .A2(n8536), .B1(n7567), .B2(n6931), .C1(
        n6930), .C2(n8258), .ZN(P2_U3277) );
  INV_X1 U8732 ( .A(n6932), .ZN(n6939) );
  NOR2_X1 U8733 ( .A1(n8745), .A2(n5247), .ZN(n6936) );
  OAI22_X1 U8734 ( .A1(n8595), .A2(n6934), .B1(n6933), .B2(n8771), .ZN(n6935)
         );
  AOI211_X1 U8735 ( .C1(n6937), .C2(n8619), .A(n6936), .B(n6935), .ZN(n6938)
         );
  OAI21_X1 U8736 ( .B1(n6939), .B2(n8725), .A(n6938), .ZN(P2_U3228) );
  INV_X1 U8737 ( .A(n6940), .ZN(n6941) );
  NAND2_X1 U8738 ( .A1(n6942), .A2(n6941), .ZN(n6944) );
  OAI22_X1 U8739 ( .A1(n6947), .A2(n4394), .B1(n10065), .B2(n8996), .ZN(n6943)
         );
  XNOR2_X1 U8740 ( .A(n6943), .B(n9068), .ZN(n6945) );
  NOR2_X1 U8741 ( .A1(n7095), .A2(n4481), .ZN(n6948) );
  OAI22_X1 U8742 ( .A1(n6947), .A2(n9065), .B1(n10065), .B2(n4394), .ZN(n7096)
         );
  XNOR2_X1 U8743 ( .A(n6948), .B(n7096), .ZN(n6953) );
  OAI22_X1 U8744 ( .A1(n6949), .A2(n9373), .B1(n7092), .B2(n9350), .ZN(n6983)
         );
  AOI22_X1 U8745 ( .A1(n6983), .A2(n9195), .B1(P1_REG3_REG_5__SCAN_IN), .B2(
        P1_U3086), .ZN(n6952) );
  INV_X1 U8746 ( .A(n6950), .ZN(n10062) );
  AOI22_X1 U8747 ( .A1(n9201), .A2(n6986), .B1(n9145), .B2(n10062), .ZN(n6951)
         );
  OAI211_X1 U8748 ( .C1(n6953), .C2(n9204), .A(n6952), .B(n6951), .ZN(P1_U3227) );
  XNOR2_X1 U8749 ( .A(n6954), .B(n6956), .ZN(n6955) );
  AOI222_X1 U8750 ( .A1(n8765), .A2(n6955), .B1(n8408), .B2(n5047), .C1(n8410), 
        .C2(n8741), .ZN(n10251) );
  XNOR2_X1 U8751 ( .A(n6957), .B(n6956), .ZN(n10254) );
  NOR2_X1 U8752 ( .A1(n8745), .A2(n5262), .ZN(n6959) );
  OAI22_X1 U8753 ( .A1(n8595), .A2(n10252), .B1(n7148), .B2(n8771), .ZN(n6958)
         );
  AOI211_X1 U8754 ( .C1(n10254), .C2(n8619), .A(n6959), .B(n6958), .ZN(n6960)
         );
  OAI21_X1 U8755 ( .B1(n10251), .B2(n8725), .A(n6960), .ZN(P2_U3227) );
  OAI21_X1 U8756 ( .B1(n6962), .B2(n6964), .A(n6961), .ZN(n6991) );
  INV_X1 U8757 ( .A(n6980), .ZN(n6963) );
  AOI211_X1 U8758 ( .C1(n6969), .C2(n6963), .A(n9540), .B(n7039), .ZN(n7002)
         );
  INV_X1 U8759 ( .A(n6964), .ZN(n7961) );
  XNOR2_X1 U8760 ( .A(n6965), .B(n7961), .ZN(n6966) );
  AOI22_X1 U8761 ( .A1(n9173), .A2(n9227), .B1(n9225), .B2(n9150), .ZN(n7100)
         );
  OAI21_X1 U8762 ( .B1(n6966), .B2(n10087), .A(n7100), .ZN(n6997) );
  AOI211_X1 U8763 ( .C1(n10161), .C2(n6991), .A(n7002), .B(n6997), .ZN(n6971)
         );
  OAI22_X1 U8764 ( .A1(n9956), .A2(n7102), .B1(n10174), .B2(n5843), .ZN(n6967)
         );
  INV_X1 U8765 ( .A(n6967), .ZN(n6968) );
  OAI21_X1 U8766 ( .B1(n6971), .B2(n10173), .A(n6968), .ZN(P1_U3471) );
  INV_X1 U8767 ( .A(n9646), .ZN(n7286) );
  AOI22_X1 U8768 ( .A1(n7286), .A2(n6969), .B1(n10184), .B2(
        P1_REG1_REG_6__SCAN_IN), .ZN(n6970) );
  OAI21_X1 U8769 ( .B1(n6971), .B2(n10184), .A(n6970), .ZN(P1_U3528) );
  OAI22_X1 U8770 ( .A1(n8595), .A2(n6973), .B1(n6972), .B2(n8771), .ZN(n6976)
         );
  MUX2_X1 U8771 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6974), .S(n8745), .Z(n6975)
         );
  AOI211_X1 U8772 ( .C1(n8619), .C2(n6977), .A(n6976), .B(n6975), .ZN(n6978)
         );
  INV_X1 U8773 ( .A(n6978), .ZN(P2_U3229) );
  XNOR2_X1 U8774 ( .A(n6979), .B(n7956), .ZN(n10067) );
  AOI211_X1 U8775 ( .C1(n6986), .C2(n7131), .A(n9540), .B(n6980), .ZN(n10061)
         );
  NAND2_X1 U8776 ( .A1(n6981), .A2(n7831), .ZN(n6982) );
  XNOR2_X1 U8777 ( .A(n6982), .B(n7956), .ZN(n6984) );
  AOI21_X1 U8778 ( .B1(n6984), .B2(n10072), .A(n6983), .ZN(n10069) );
  INV_X1 U8779 ( .A(n10069), .ZN(n6985) );
  AOI211_X1 U8780 ( .C1(n10067), .C2(n10161), .A(n10061), .B(n6985), .ZN(n6990) );
  AOI22_X1 U8781 ( .A1(n7286), .A2(n6986), .B1(n10184), .B2(
        P1_REG1_REG_5__SCAN_IN), .ZN(n6987) );
  OAI21_X1 U8782 ( .B1(n6990), .B2(n10184), .A(n6987), .ZN(P1_U3527) );
  OAI22_X1 U8783 ( .A1(n9956), .A2(n10065), .B1(n10174), .B2(n5831), .ZN(n6988) );
  INV_X1 U8784 ( .A(n6988), .ZN(n6989) );
  OAI21_X1 U8785 ( .B1(n6990), .B2(n10173), .A(n6989), .ZN(P1_U3468) );
  INV_X1 U8786 ( .A(n6991), .ZN(n7005) );
  NAND2_X1 U8787 ( .A1(n7330), .A2(n10092), .ZN(n6996) );
  NAND2_X1 U8788 ( .A1(n6997), .A2(n9562), .ZN(n7004) );
  NOR2_X1 U8789 ( .A1(n10096), .A2(n7102), .ZN(n7001) );
  OAI22_X1 U8790 ( .A1(n9562), .A2(n6999), .B1(n7101), .B2(n9559), .ZN(n7000)
         );
  AOI211_X1 U8791 ( .C1(n7002), .C2(n10081), .A(n7001), .B(n7000), .ZN(n7003)
         );
  OAI211_X1 U8792 ( .C1(n7005), .C2(n9557), .A(n7004), .B(n7003), .ZN(P1_U3287) );
  INV_X1 U8793 ( .A(n7006), .ZN(n7007) );
  OAI222_X1 U8794 ( .A1(n9966), .A2(n9874), .B1(n9969), .B2(n7007), .C1(
        P1_U3086), .C2(n9342), .ZN(P1_U3336) );
  OAI222_X1 U8795 ( .A1(n8258), .A2(n7008), .B1(n7567), .B2(n7007), .C1(
        P2_U3151), .C2(n8555), .ZN(P2_U3276) );
  AOI21_X1 U8796 ( .B1(n10081), .B2(n10094), .A(n10074), .ZN(n7019) );
  INV_X1 U8797 ( .A(n7955), .ZN(n7011) );
  NAND3_X1 U8798 ( .A1(n7011), .A2(n7010), .A3(n7009), .ZN(n7014) );
  INV_X1 U8799 ( .A(n7012), .ZN(n7013) );
  OAI211_X1 U8800 ( .C1(n6629), .C2(n9559), .A(n7014), .B(n7013), .ZN(n7017)
         );
  NOR2_X1 U8801 ( .A1(n9562), .A2(n7015), .ZN(n7016) );
  AOI21_X1 U8802 ( .B1(n7017), .B2(n9562), .A(n7016), .ZN(n7018) );
  OAI21_X1 U8803 ( .B1(n7019), .B2(n10095), .A(n7018), .ZN(P1_U3293) );
  INV_X1 U8804 ( .A(n7021), .ZN(n7954) );
  XNOR2_X1 U8805 ( .A(n7020), .B(n7954), .ZN(n10129) );
  XNOR2_X1 U8806 ( .A(n7834), .B(n7954), .ZN(n7023) );
  OAI21_X1 U8807 ( .B1(n7023), .B2(n10087), .A(n7022), .ZN(n10131) );
  NAND2_X1 U8808 ( .A1(n10131), .A2(n9562), .ZN(n7029) );
  OAI22_X1 U8809 ( .A1(n9562), .A2(n7024), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9559), .ZN(n7026) );
  OAI211_X1 U8810 ( .C1(n10077), .C2(n5810), .A(n7130), .B(n10094), .ZN(n10130) );
  NOR2_X1 U8811 ( .A1(n10130), .A2(n10097), .ZN(n7025) );
  AOI211_X1 U8812 ( .C1(n10074), .C2(n7027), .A(n7026), .B(n7025), .ZN(n7028)
         );
  OAI211_X1 U8813 ( .C1(n10129), .C2(n9557), .A(n7029), .B(n7028), .ZN(
        P1_U3290) );
  INV_X1 U8814 ( .A(n10092), .ZN(n7038) );
  OAI21_X1 U8815 ( .B1(n7031), .B2(n7840), .A(n7030), .ZN(n7071) );
  INV_X1 U8816 ( .A(n7071), .ZN(n7037) );
  AOI22_X1 U8817 ( .A1(n9173), .A2(n9226), .B1(n9224), .B2(n9150), .ZN(n7181)
         );
  NAND2_X1 U8818 ( .A1(n7760), .A2(n7032), .ZN(n7837) );
  INV_X1 U8819 ( .A(n7837), .ZN(n7845) );
  NAND2_X1 U8820 ( .A1(n7033), .A2(n7845), .ZN(n7034) );
  AOI21_X1 U8821 ( .B1(n7034), .B2(n7848), .A(n7840), .ZN(n7248) );
  AND3_X1 U8822 ( .A1(n7034), .A2(n7848), .A3(n7840), .ZN(n7035) );
  OAI21_X1 U8823 ( .B1(n7248), .B2(n7035), .A(n10072), .ZN(n7036) );
  OAI211_X1 U8824 ( .C1(n7037), .C2(n7330), .A(n7181), .B(n7036), .ZN(n7069)
         );
  AOI21_X1 U8825 ( .B1(n7038), .B2(n7071), .A(n7069), .ZN(n7046) );
  INV_X1 U8826 ( .A(n7039), .ZN(n7041) );
  INV_X1 U8827 ( .A(n7111), .ZN(n7040) );
  AOI211_X1 U8828 ( .C1(n7185), .C2(n7041), .A(n9540), .B(n7040), .ZN(n7070)
         );
  NOR2_X1 U8829 ( .A1(n10096), .A2(n7176), .ZN(n7044) );
  OAI22_X1 U8830 ( .A1(n9562), .A2(n7042), .B1(n7183), .B2(n9559), .ZN(n7043)
         );
  AOI211_X1 U8831 ( .C1(n7070), .C2(n10081), .A(n7044), .B(n7043), .ZN(n7045)
         );
  OAI21_X1 U8832 ( .B1(n7046), .B2(n10102), .A(n7045), .ZN(P1_U3286) );
  INV_X1 U8833 ( .A(n7047), .ZN(n7048) );
  OAI22_X1 U8834 ( .A1(n7050), .A2(n7049), .B1(n4853), .B2(n7048), .ZN(n7157)
         );
  MUX2_X1 U8835 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8551), .Z(n7153) );
  XOR2_X1 U8836 ( .A(n7160), .B(n7153), .Z(n7156) );
  XNOR2_X1 U8837 ( .A(n7157), .B(n7156), .ZN(n7067) );
  XNOR2_X1 U8838 ( .A(n7160), .B(n7219), .ZN(n7052) );
  NAND2_X1 U8839 ( .A1(n7051), .A2(n7052), .ZN(n7162) );
  INV_X1 U8840 ( .A(n7052), .ZN(n7054) );
  NAND3_X1 U8841 ( .A1(n7055), .A2(n7054), .A3(n7053), .ZN(n7056) );
  AOI21_X1 U8842 ( .B1(n7162), .B2(n7056), .A(n10220), .ZN(n7066) );
  INV_X1 U8843 ( .A(n7057), .ZN(n7058) );
  XNOR2_X1 U8844 ( .A(n7160), .B(P2_REG1_REG_8__SCAN_IN), .ZN(n7059) );
  AOI21_X1 U8845 ( .B1(n7060), .B2(n7058), .A(n7059), .ZN(n7151) );
  AND3_X1 U8846 ( .A1(n7060), .A2(n7059), .A3(n7058), .ZN(n7061) );
  OAI21_X1 U8847 ( .B1(n7151), .B2(n7061), .A(n10197), .ZN(n7064) );
  INV_X1 U8848 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7062) );
  NOR2_X1 U8849 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7062), .ZN(n7316) );
  AOI21_X1 U8850 ( .B1(n10212), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n7316), .ZN(
        n7063) );
  OAI211_X1 U8851 ( .C1(n10204), .C2(n7160), .A(n7064), .B(n7063), .ZN(n7065)
         );
  AOI211_X1 U8852 ( .C1(n7067), .C2(n10225), .A(n7066), .B(n7065), .ZN(n7068)
         );
  INV_X1 U8853 ( .A(n7068), .ZN(P2_U3190) );
  AOI211_X1 U8854 ( .C1(n10148), .C2(n7071), .A(n7070), .B(n7069), .ZN(n7075)
         );
  OAI22_X1 U8855 ( .A1(n9956), .A2(n7176), .B1(n10174), .B2(n5857), .ZN(n7072)
         );
  INV_X1 U8856 ( .A(n7072), .ZN(n7073) );
  OAI21_X1 U8857 ( .B1(n7075), .B2(n10173), .A(n7073), .ZN(P1_U3474) );
  AOI22_X1 U8858 ( .A1(n7286), .A2(n7185), .B1(n10184), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n7074) );
  OAI21_X1 U8859 ( .B1(n7075), .B2(n10184), .A(n7074), .ZN(P1_U3529) );
  AOI22_X1 U8860 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n7269), .B1(n7262), .B2(
        n7493), .ZN(n7078) );
  OAI21_X1 U8861 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7079), .A(n7076), .ZN(
        n7077) );
  NOR2_X1 U8862 ( .A1(n7078), .A2(n7077), .ZN(n7261) );
  AOI211_X1 U8863 ( .C1(n7078), .C2(n7077), .A(n7261), .B(n10044), .ZN(n7090)
         );
  NOR2_X1 U8864 ( .A1(n7079), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7080) );
  NOR2_X1 U8865 ( .A1(n7081), .A2(n7080), .ZN(n7084) );
  MUX2_X1 U8866 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n7082), .S(n7262), .Z(n7083)
         );
  NAND2_X1 U8867 ( .A1(n7083), .A2(n7084), .ZN(n7268) );
  OAI211_X1 U8868 ( .C1(n7084), .C2(n7083), .A(n7268), .B(n10057), .ZN(n7088)
         );
  NOR2_X1 U8869 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7085), .ZN(n7086) );
  AOI21_X1 U8870 ( .B1(n10043), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n7086), .ZN(
        n7087) );
  OAI211_X1 U8871 ( .C1(n9335), .C2(n7269), .A(n7088), .B(n7087), .ZN(n7089)
         );
  OR2_X1 U8872 ( .A1(n7090), .A2(n7089), .ZN(P1_U3256) );
  OAI22_X1 U8873 ( .A1(n7092), .A2(n4394), .B1(n7102), .B2(n8996), .ZN(n7091)
         );
  XNOR2_X1 U8874 ( .A(n7091), .B(n8997), .ZN(n7094) );
  OAI22_X1 U8875 ( .A1(n7092), .A2(n9065), .B1(n7102), .B2(n4394), .ZN(n7093)
         );
  NOR2_X1 U8876 ( .A1(n7094), .A2(n7093), .ZN(n7172) );
  AOI21_X1 U8877 ( .B1(n7094), .B2(n7093), .A(n7172), .ZN(n7098) );
  OAI21_X1 U8878 ( .B1(n7098), .B2(n7097), .A(n7174), .ZN(n7105) );
  OAI21_X1 U8879 ( .B1(n7100), .B2(n9143), .A(n7099), .ZN(n7104) );
  OAI22_X1 U8880 ( .A1(n9191), .A2(n7102), .B1(n9198), .B2(n7101), .ZN(n7103)
         );
  AOI211_X1 U8881 ( .C1(n7105), .C2(n9184), .A(n7104), .B(n7103), .ZN(n7106)
         );
  INV_X1 U8882 ( .A(n7106), .ZN(P1_U3239) );
  INV_X1 U8883 ( .A(n7107), .ZN(n7125) );
  OAI222_X1 U8884 ( .A1(n9969), .A2(n7125), .B1(n7108), .B2(P1_U3086), .C1(
        n9766), .C2(n9966), .ZN(P1_U3335) );
  OAI21_X1 U8885 ( .B1(n7110), .B2(n7115), .A(n7109), .ZN(n9565) );
  AOI21_X1 U8886 ( .B1(n7111), .B2(n9564), .A(n9540), .ZN(n7112) );
  AND2_X1 U8887 ( .A1(n7112), .A2(n7255), .ZN(n9566) );
  INV_X1 U8888 ( .A(n7248), .ZN(n7114) );
  NAND2_X1 U8889 ( .A1(n7114), .A2(n7113), .ZN(n7116) );
  XNOR2_X1 U8890 ( .A(n7116), .B(n7115), .ZN(n7120) );
  OR2_X1 U8891 ( .A1(n7177), .A2(n9373), .ZN(n7118) );
  OR2_X1 U8892 ( .A1(n7445), .A2(n9350), .ZN(n7117) );
  NAND2_X1 U8893 ( .A1(n7118), .A2(n7117), .ZN(n9091) );
  INV_X1 U8894 ( .A(n9091), .ZN(n7119) );
  OAI21_X1 U8895 ( .B1(n7120), .B2(n10087), .A(n7119), .ZN(n9558) );
  AOI211_X1 U8896 ( .C1(n10161), .C2(n9565), .A(n9566), .B(n9558), .ZN(n7124)
         );
  AOI22_X1 U8897 ( .A1(n7286), .A2(n9564), .B1(n10184), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n7121) );
  OAI21_X1 U8898 ( .B1(n7124), .B2(n10184), .A(n7121), .ZN(P1_U3530) );
  OAI22_X1 U8899 ( .A1(n9956), .A2(n7437), .B1(n10174), .B2(n5870), .ZN(n7122)
         );
  INV_X1 U8900 ( .A(n7122), .ZN(n7123) );
  OAI21_X1 U8901 ( .B1(n7124), .B2(n10173), .A(n7123), .ZN(P1_U3477) );
  OAI222_X1 U8902 ( .A1(n8258), .A2(n9924), .B1(n7567), .B2(n7125), .C1(n8203), 
        .C2(P2_U3151), .ZN(P2_U3275) );
  AND2_X1 U8903 ( .A1(n7831), .A2(n7836), .ZN(n7827) );
  XNOR2_X1 U8904 ( .A(n7126), .B(n7827), .ZN(n7128) );
  AOI21_X1 U8905 ( .B1(n7128), .B2(n10072), .A(n7127), .ZN(n10136) );
  INV_X1 U8906 ( .A(n7827), .ZN(n7957) );
  XNOR2_X1 U8907 ( .A(n7129), .B(n7957), .ZN(n10139) );
  INV_X1 U8908 ( .A(n7130), .ZN(n7132) );
  OAI211_X1 U8909 ( .C1(n7132), .C2(n10135), .A(n10094), .B(n7131), .ZN(n10134) );
  OAI22_X1 U8910 ( .A1(n9562), .A2(n7134), .B1(n7133), .B2(n9559), .ZN(n7135)
         );
  AOI21_X1 U8911 ( .B1(n10074), .B2(n7136), .A(n7135), .ZN(n7137) );
  OAI21_X1 U8912 ( .B1(n10134), .B2(n10097), .A(n7137), .ZN(n7138) );
  AOI21_X1 U8913 ( .B1(n10139), .B2(n10082), .A(n7138), .ZN(n7139) );
  OAI21_X1 U8914 ( .B1(n10136), .B2(n10102), .A(n7139), .ZN(P1_U3289) );
  INV_X1 U8915 ( .A(n7140), .ZN(n7141) );
  AOI211_X1 U8916 ( .C1(n7143), .C2(n7142), .A(n8381), .B(n7141), .ZN(n7150)
         );
  AOI22_X1 U8917 ( .A1(n8372), .A2(n8408), .B1(n8390), .B2(n8410), .ZN(n7147)
         );
  AOI21_X1 U8918 ( .B1(n8379), .B2(n7145), .A(n7144), .ZN(n7146) );
  OAI211_X1 U8919 ( .C1(n8339), .C2(n7148), .A(n7147), .B(n7146), .ZN(n7149)
         );
  OR2_X1 U8920 ( .A1(n7150), .A2(n7149), .ZN(P2_U3179) );
  INV_X1 U8921 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10297) );
  AOI21_X1 U8922 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n7160), .A(n7151), .ZN(
        n7225) );
  AOI21_X1 U8923 ( .B1(n10297), .B2(n7152), .A(n7226), .ZN(n7171) );
  INV_X1 U8924 ( .A(n7160), .ZN(n7155) );
  INV_X1 U8925 ( .A(n7153), .ZN(n7154) );
  AOI22_X1 U8926 ( .A1(n7157), .A2(n7156), .B1(n7155), .B2(n7154), .ZN(n7232)
         );
  MUX2_X1 U8927 ( .A(n5304), .B(n10297), .S(n8551), .Z(n7228) );
  XNOR2_X1 U8928 ( .A(n7228), .B(n7168), .ZN(n7231) );
  XNOR2_X1 U8929 ( .A(n7232), .B(n7231), .ZN(n7158) );
  NAND2_X1 U8930 ( .A1(n7158), .A2(n10225), .ZN(n7170) );
  INV_X1 U8931 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n9995) );
  AND2_X1 U8932 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7460) );
  INV_X1 U8933 ( .A(n7460), .ZN(n7159) );
  OAI21_X1 U8934 ( .B1(n10192), .B2(n9995), .A(n7159), .ZN(n7167) );
  NAND2_X1 U8935 ( .A1(n7160), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7161) );
  NAND2_X1 U8936 ( .A1(n7162), .A2(n7161), .ZN(n7163) );
  NAND2_X1 U8937 ( .A1(n7163), .A2(n7229), .ZN(n7238) );
  OAI21_X1 U8938 ( .B1(n7163), .B2(n7229), .A(n7238), .ZN(n7164) );
  NAND2_X1 U8939 ( .A1(n7164), .A2(n5304), .ZN(n7165) );
  AOI21_X1 U8940 ( .B1(n7240), .B2(n7165), .A(n10220), .ZN(n7166) );
  AOI211_X1 U8941 ( .C1(n10213), .C2(n7168), .A(n7167), .B(n7166), .ZN(n7169)
         );
  OAI211_X1 U8942 ( .C1(n7171), .C2(n10229), .A(n7170), .B(n7169), .ZN(
        P2_U3191) );
  INV_X1 U8943 ( .A(n7172), .ZN(n7173) );
  OAI22_X1 U8944 ( .A1(n7177), .A2(n4394), .B1(n7176), .B2(n8996), .ZN(n7175)
         );
  XNOR2_X1 U8945 ( .A(n7175), .B(n8997), .ZN(n7179) );
  OAI22_X1 U8946 ( .A1(n7177), .A2(n9065), .B1(n7176), .B2(n4394), .ZN(n7178)
         );
  NAND2_X1 U8947 ( .A1(n7179), .A2(n7178), .ZN(n7439) );
  NAND2_X1 U8948 ( .A1(n4478), .A2(n7439), .ZN(n7180) );
  XNOR2_X1 U8949 ( .A(n7440), .B(n7180), .ZN(n7188) );
  INV_X1 U8950 ( .A(n7181), .ZN(n7182) );
  AOI22_X1 U8951 ( .A1(n7182), .A2(n9195), .B1(P1_REG3_REG_7__SCAN_IN), .B2(
        P1_U3086), .ZN(n7187) );
  INV_X1 U8952 ( .A(n7183), .ZN(n7184) );
  AOI22_X1 U8953 ( .A1(n9201), .A2(n7185), .B1(n9145), .B2(n7184), .ZN(n7186)
         );
  OAI211_X1 U8954 ( .C1(n7188), .C2(n9204), .A(n7187), .B(n7186), .ZN(P1_U3213) );
  INV_X1 U8955 ( .A(n7189), .ZN(n7213) );
  OAI222_X1 U8956 ( .A1(n9969), .A2(n7213), .B1(n7952), .B2(P1_U3086), .C1(
        n7190), .C2(n9966), .ZN(P1_U3334) );
  XNOR2_X1 U8957 ( .A(n7191), .B(n8220), .ZN(n7194) );
  INV_X1 U8958 ( .A(n7194), .ZN(n10256) );
  INV_X1 U8959 ( .A(n7216), .ZN(n7192) );
  AOI21_X1 U8960 ( .B1(n8220), .B2(n7193), .A(n7192), .ZN(n7197) );
  AOI22_X1 U8961 ( .A1(n8409), .A2(n8741), .B1(n5047), .B2(n8407), .ZN(n7196)
         );
  INV_X1 U8962 ( .A(n7479), .ZN(n8755) );
  NAND2_X1 U8963 ( .A1(n7194), .A2(n8755), .ZN(n7195) );
  OAI211_X1 U8964 ( .C1(n7197), .C2(n8629), .A(n7196), .B(n7195), .ZN(n10258)
         );
  NAND2_X1 U8965 ( .A1(n10258), .A2(n8745), .ZN(n7201) );
  OAI22_X1 U8966 ( .A1(n8745), .A2(n6909), .B1(n7212), .B2(n8771), .ZN(n7198)
         );
  AOI21_X1 U8967 ( .B1(n8749), .B2(n7199), .A(n7198), .ZN(n7200) );
  OAI211_X1 U8968 ( .C1(n10256), .C2(n7484), .A(n7201), .B(n7200), .ZN(
        P2_U3226) );
  OAI21_X1 U8969 ( .B1(n7204), .B2(n7203), .A(n7202), .ZN(n7205) );
  NAND2_X1 U8970 ( .A1(n7205), .A2(n8387), .ZN(n7211) );
  INV_X1 U8971 ( .A(n7206), .ZN(n7209) );
  OAI22_X1 U8972 ( .A1(n8376), .A2(n7207), .B1(n8397), .B2(n10255), .ZN(n7208)
         );
  AOI211_X1 U8973 ( .C1(n8372), .C2(n8407), .A(n7209), .B(n7208), .ZN(n7210)
         );
  OAI211_X1 U8974 ( .C1(n7212), .C2(n8339), .A(n7211), .B(n7210), .ZN(P2_U3153) );
  OAI222_X1 U8975 ( .A1(n8258), .A2(n9776), .B1(n7567), .B2(n7213), .C1(n8241), 
        .C2(P2_U3151), .ZN(P2_U3274) );
  INV_X1 U8976 ( .A(n7221), .ZN(n8219) );
  NAND3_X1 U8977 ( .A1(n7216), .A2(n8219), .A3(n7215), .ZN(n7217) );
  NAND2_X1 U8978 ( .A1(n7214), .A2(n7217), .ZN(n7218) );
  AOI222_X1 U8979 ( .A1(n8765), .A2(n7218), .B1(n8406), .B2(n5047), .C1(n8408), 
        .C2(n8741), .ZN(n10260) );
  OAI22_X1 U8980 ( .A1(n8745), .A2(n7219), .B1(n7318), .B2(n8771), .ZN(n7220)
         );
  AOI21_X1 U8981 ( .B1(n8749), .B2(n7326), .A(n7220), .ZN(n7224) );
  XNOR2_X1 U8982 ( .A(n7222), .B(n7221), .ZN(n10263) );
  NAND2_X1 U8983 ( .A1(n10263), .A2(n8619), .ZN(n7223) );
  OAI211_X1 U8984 ( .C1(n10260), .C2(n8725), .A(n7224), .B(n7223), .ZN(
        P2_U3225) );
  AOI22_X1 U8985 ( .A1(n7244), .A2(P2_REG1_REG_10__SCAN_IN), .B1(n5328), .B2(
        n7366), .ZN(n7227) );
  AOI21_X1 U8986 ( .B1(n4479), .B2(n7227), .A(n7357), .ZN(n7247) );
  INV_X1 U8987 ( .A(n7228), .ZN(n7230) );
  OAI22_X1 U8988 ( .A1(n7232), .A2(n7231), .B1(n7230), .B2(n7229), .ZN(n7235)
         );
  NAND2_X1 U8989 ( .A1(n8551), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7233) );
  OAI21_X1 U8990 ( .B1(n8551), .B2(n7480), .A(n7233), .ZN(n7361) );
  XNOR2_X1 U8991 ( .A(n7361), .B(n7244), .ZN(n7234) );
  NAND2_X1 U8992 ( .A1(n7234), .A2(n7235), .ZN(n7362) );
  OAI21_X1 U8993 ( .B1(n7235), .B2(n7234), .A(n7362), .ZN(n7236) );
  NAND2_X1 U8994 ( .A1(n7236), .A2(n10225), .ZN(n7246) );
  INV_X1 U8995 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n9998) );
  AND2_X1 U8996 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7676) );
  INV_X1 U8997 ( .A(n7676), .ZN(n7237) );
  OAI21_X1 U8998 ( .B1(n10192), .B2(n9998), .A(n7237), .ZN(n7243) );
  MUX2_X1 U8999 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n7480), .S(n7244), .Z(n7239)
         );
  NAND3_X1 U9000 ( .A1(n7240), .A2(n7239), .A3(n7238), .ZN(n7241) );
  AOI21_X1 U9001 ( .B1(n4480), .B2(n7241), .A(n10220), .ZN(n7242) );
  AOI211_X1 U9002 ( .C1(n10213), .C2(n7244), .A(n7243), .B(n7242), .ZN(n7245)
         );
  OAI211_X1 U9003 ( .C1(n7247), .C2(n10229), .A(n7246), .B(n7245), .ZN(
        P2_U3192) );
  OAI21_X1 U9004 ( .B1(n7248), .B2(n7853), .A(n7850), .ZN(n7249) );
  XNOR2_X1 U9005 ( .A(n7249), .B(n7252), .ZN(n7250) );
  NOR2_X1 U9006 ( .A1(n7441), .A2(n9373), .ZN(n7449) );
  AOI21_X1 U9007 ( .B1(n7250), .B2(n10072), .A(n7449), .ZN(n10141) );
  OAI21_X1 U9008 ( .B1(n7253), .B2(n7252), .A(n7251), .ZN(n10144) );
  NAND2_X1 U9009 ( .A1(n10144), .A2(n10082), .ZN(n7260) );
  OAI22_X1 U9010 ( .A1(n9562), .A2(n7254), .B1(n7453), .B2(n9559), .ZN(n7258)
         );
  XNOR2_X1 U9011 ( .A(n7255), .B(n10142), .ZN(n7256) );
  NOR2_X1 U9012 ( .A1(n7542), .A2(n9350), .ZN(n7450) );
  AOI21_X1 U9013 ( .B1(n7256), .B2(n10094), .A(n7450), .ZN(n10140) );
  NOR2_X1 U9014 ( .A1(n10140), .A2(n10097), .ZN(n7257) );
  AOI211_X1 U9015 ( .C1(n10074), .C2(n7455), .A(n7258), .B(n7257), .ZN(n7259)
         );
  OAI211_X1 U9016 ( .C1(n10102), .C2(n10141), .A(n7260), .B(n7259), .ZN(
        P1_U3284) );
  NAND2_X1 U9017 ( .A1(P1_REG2_REG_14__SCAN_IN), .A2(n9261), .ZN(n7263) );
  OAI21_X1 U9018 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n9261), .A(n7263), .ZN(
        n7264) );
  AOI211_X1 U9019 ( .C1(n7265), .C2(n7264), .A(n9260), .B(n10044), .ZN(n7276)
         );
  NOR2_X1 U9020 ( .A1(n9264), .A2(n7266), .ZN(n7267) );
  AOI21_X1 U9021 ( .B1(n7266), .B2(n9264), .A(n7267), .ZN(n7271) );
  OAI21_X1 U9022 ( .B1(n7269), .B2(n7082), .A(n7268), .ZN(n7270) );
  NAND2_X1 U9023 ( .A1(n7271), .A2(n7270), .ZN(n9263) );
  OAI211_X1 U9024 ( .C1(n7271), .C2(n7270), .A(n10057), .B(n9263), .ZN(n7274)
         );
  AND2_X1 U9025 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n7272) );
  AOI21_X1 U9026 ( .B1(n10043), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n7272), .ZN(
        n7273) );
  OAI211_X1 U9027 ( .C1(n9335), .C2(n9264), .A(n7274), .B(n7273), .ZN(n7275)
         );
  OR2_X1 U9028 ( .A1(n7276), .A2(n7275), .ZN(P1_U3257) );
  OAI21_X1 U9029 ( .B1(n7278), .B2(n7964), .A(n7277), .ZN(n7291) );
  INV_X1 U9030 ( .A(n7279), .ZN(n7280) );
  AOI211_X1 U9031 ( .C1(n9049), .C2(n7280), .A(n9540), .B(n7328), .ZN(n7292)
         );
  XOR2_X1 U9032 ( .A(n7964), .B(n7281), .Z(n7285) );
  OR2_X1 U9033 ( .A1(n7445), .A2(n9373), .ZN(n7283) );
  NAND2_X1 U9034 ( .A1(n9221), .A2(n9150), .ZN(n7282) );
  NAND2_X1 U9035 ( .A1(n7283), .A2(n7282), .ZN(n9048) );
  INV_X1 U9036 ( .A(n9048), .ZN(n7284) );
  OAI21_X1 U9037 ( .B1(n7285), .B2(n10087), .A(n7284), .ZN(n7298) );
  AOI211_X1 U9038 ( .C1(n7291), .C2(n10161), .A(n7292), .B(n7298), .ZN(n7290)
         );
  AOI22_X1 U9039 ( .A1(n9049), .A2(n7286), .B1(n10184), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n7287) );
  OAI21_X1 U9040 ( .B1(n7290), .B2(n10184), .A(n7287), .ZN(P1_U3532) );
  OAI22_X1 U9041 ( .A1(n7296), .A2(n9956), .B1(n10174), .B2(n5895), .ZN(n7288)
         );
  INV_X1 U9042 ( .A(n7288), .ZN(n7289) );
  OAI21_X1 U9043 ( .B1(n7290), .B2(n10173), .A(n7289), .ZN(P1_U3483) );
  INV_X1 U9044 ( .A(n7291), .ZN(n7300) );
  NAND2_X1 U9045 ( .A1(n7292), .A2(n10081), .ZN(n7295) );
  INV_X1 U9046 ( .A(n7293), .ZN(n9050) );
  AOI22_X1 U9047 ( .A1(n10102), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n9050), .B2(
        n10091), .ZN(n7294) );
  OAI211_X1 U9048 ( .C1(n7296), .C2(n10096), .A(n7295), .B(n7294), .ZN(n7297)
         );
  AOI21_X1 U9049 ( .B1(n9562), .B2(n7298), .A(n7297), .ZN(n7299) );
  OAI21_X1 U9050 ( .B1(n7300), .B2(n9557), .A(n7299), .ZN(P1_U3283) );
  INV_X1 U9051 ( .A(n7301), .ZN(n7305) );
  OAI222_X1 U9052 ( .A1(n8258), .A2(n7303), .B1(n7567), .B2(n7305), .C1(
        P2_U3151), .C2(n7302), .ZN(P2_U3273) );
  OAI222_X1 U9053 ( .A1(n9966), .A2(n7306), .B1(n9969), .B2(n7305), .C1(
        P1_U3086), .C2(n7304), .ZN(P1_U3333) );
  NAND2_X1 U9054 ( .A1(n7310), .A2(n7307), .ZN(n7308) );
  OAI211_X1 U9055 ( .C1(n9756), .C2(n8258), .A(n7308), .B(n8243), .ZN(P2_U3272) );
  NAND2_X1 U9056 ( .A1(n7310), .A2(n7309), .ZN(n7312) );
  OR2_X1 U9057 ( .A1(n7311), .A2(P1_U3086), .ZN(n8017) );
  OAI211_X1 U9058 ( .C1(n7313), .C2(n9966), .A(n7312), .B(n8017), .ZN(P1_U3332) );
  NOR2_X1 U9059 ( .A1(n8392), .A2(n7314), .ZN(n7315) );
  AOI211_X1 U9060 ( .C1(n8390), .C2(n8408), .A(n7316), .B(n7315), .ZN(n7317)
         );
  OAI21_X1 U9061 ( .B1(n7318), .B2(n8339), .A(n7317), .ZN(n7325) );
  INV_X1 U9062 ( .A(n7319), .ZN(n7321) );
  NAND3_X1 U9063 ( .A1(n7202), .A2(n7321), .A3(n7320), .ZN(n7322) );
  AOI21_X1 U9064 ( .B1(n7323), .B2(n7322), .A(n8381), .ZN(n7324) );
  AOI211_X1 U9065 ( .C1(n7326), .C2(n8379), .A(n7325), .B(n7324), .ZN(n7327)
         );
  INV_X1 U9066 ( .A(n7327), .ZN(P2_U3161) );
  OAI211_X1 U9067 ( .C1(n7328), .C2(n10146), .A(n10094), .B(n7388), .ZN(n10145) );
  INV_X1 U9068 ( .A(n7866), .ZN(n7333) );
  XNOR2_X1 U9069 ( .A(n7329), .B(n7967), .ZN(n10149) );
  INV_X1 U9070 ( .A(n10149), .ZN(n7339) );
  INV_X1 U9071 ( .A(n7330), .ZN(n10172) );
  AOI21_X1 U9072 ( .B1(n7331), .B2(n7967), .A(n10087), .ZN(n7332) );
  OAI21_X1 U9073 ( .B1(n7384), .B2(n7333), .A(n7332), .ZN(n7337) );
  OR2_X1 U9074 ( .A1(n7542), .A2(n9373), .ZN(n7335) );
  OR2_X1 U9075 ( .A1(n7552), .A2(n9350), .ZN(n7334) );
  NAND2_X1 U9076 ( .A1(n7335), .A2(n7334), .ZN(n7656) );
  INV_X1 U9077 ( .A(n7656), .ZN(n7336) );
  NAND2_X1 U9078 ( .A1(n7337), .A2(n7336), .ZN(n7338) );
  AOI21_X1 U9079 ( .B1(n10149), .B2(n10172), .A(n7338), .ZN(n10151) );
  OAI21_X1 U9080 ( .B1(n7339), .B2(n10092), .A(n10151), .ZN(n7340) );
  NAND2_X1 U9081 ( .A1(n7340), .A2(n9562), .ZN(n7345) );
  OAI22_X1 U9082 ( .A1(n9562), .A2(n7341), .B1(n7660), .B2(n9559), .ZN(n7342)
         );
  AOI21_X1 U9083 ( .B1(n7343), .B2(n10074), .A(n7342), .ZN(n7344) );
  OAI211_X1 U9084 ( .C1(n10097), .C2(n10145), .A(n7345), .B(n7344), .ZN(
        P1_U3282) );
  XNOR2_X1 U9085 ( .A(n7346), .B(n7348), .ZN(n10264) );
  AOI22_X1 U9086 ( .A1(n8405), .A2(n5047), .B1(n8741), .B2(n8407), .ZN(n7353)
         );
  INV_X1 U9087 ( .A(n7347), .ZN(n7351) );
  AND3_X1 U9088 ( .A1(n7214), .A2(n4607), .A3(n7349), .ZN(n7350) );
  OAI21_X1 U9089 ( .B1(n7351), .B2(n7350), .A(n8765), .ZN(n7352) );
  OAI211_X1 U9090 ( .C1(n10264), .C2(n7479), .A(n7353), .B(n7352), .ZN(n10265)
         );
  NAND2_X1 U9091 ( .A1(n10265), .A2(n8745), .ZN(n7356) );
  OAI22_X1 U9092 ( .A1(n8745), .A2(n5304), .B1(n7461), .B2(n8771), .ZN(n7354)
         );
  AOI21_X1 U9093 ( .B1(n8749), .B2(n10267), .A(n7354), .ZN(n7355) );
  OAI211_X1 U9094 ( .C1(n10264), .C2(n7484), .A(n7356), .B(n7355), .ZN(
        P2_U3224) );
  INV_X1 U9095 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10300) );
  NOR2_X1 U9096 ( .A1(n10300), .A2(n7358), .ZN(n7410) );
  AOI21_X1 U9097 ( .B1(n10300), .B2(n7358), .A(n7410), .ZN(n7377) );
  NAND2_X1 U9098 ( .A1(n8551), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7359) );
  OAI21_X1 U9099 ( .B1(n8551), .B2(n7360), .A(n7359), .ZN(n7417) );
  XNOR2_X1 U9100 ( .A(n7417), .B(n7424), .ZN(n7365) );
  OR2_X1 U9101 ( .A1(n7366), .A2(n7361), .ZN(n7363) );
  NAND2_X1 U9102 ( .A1(n7363), .A2(n7362), .ZN(n7364) );
  NAND2_X1 U9103 ( .A1(n7365), .A2(n7364), .ZN(n7419) );
  OAI21_X1 U9104 ( .B1(n7365), .B2(n7364), .A(n7419), .ZN(n7375) );
  NOR2_X1 U9105 ( .A1(n10204), .A2(n7418), .ZN(n7374) );
  INV_X1 U9106 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n10002) );
  NOR2_X1 U9107 ( .A1(n7360), .A2(n7367), .ZN(n7425) );
  AND2_X1 U9108 ( .A1(n7367), .A2(n7360), .ZN(n7369) );
  OAI21_X1 U9109 ( .B1(n7425), .B2(n7369), .A(n7368), .ZN(n7372) );
  INV_X1 U9110 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7370) );
  NOR2_X1 U9111 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7370), .ZN(n7704) );
  INV_X1 U9112 ( .A(n7704), .ZN(n7371) );
  OAI211_X1 U9113 ( .C1(n10002), .C2(n10192), .A(n7372), .B(n7371), .ZN(n7373)
         );
  AOI211_X1 U9114 ( .C1(n10225), .C2(n7375), .A(n7374), .B(n7373), .ZN(n7376)
         );
  OAI21_X1 U9115 ( .B1(n7377), .B2(n10229), .A(n7376), .ZN(P2_U3193) );
  INV_X1 U9116 ( .A(n7378), .ZN(n7382) );
  OAI222_X1 U9117 ( .A1(n9969), .A2(n7382), .B1(P1_U3086), .B2(n7380), .C1(
        n7379), .C2(n9966), .ZN(P1_U3331) );
  OAI222_X1 U9118 ( .A1(P2_U3151), .A2(n5598), .B1(n8918), .B2(n7382), .C1(
        n7381), .C2(n8258), .ZN(P2_U3271) );
  AND2_X1 U9119 ( .A1(n7969), .A2(n7866), .ZN(n7383) );
  AOI21_X1 U9120 ( .B1(n7384), .B2(n7383), .A(n10087), .ZN(n7386) );
  NAND2_X1 U9121 ( .A1(n9221), .A2(n9173), .ZN(n7385) );
  OAI21_X1 U9122 ( .B1(n7594), .B2(n9350), .A(n7385), .ZN(n7557) );
  AOI21_X1 U9123 ( .B1(n7485), .B2(n7386), .A(n7557), .ZN(n10153) );
  XNOR2_X1 U9124 ( .A(n7387), .B(n7969), .ZN(n10156) );
  NAND2_X1 U9125 ( .A1(n10156), .A2(n10082), .ZN(n7393) );
  OAI22_X1 U9126 ( .A1(n9562), .A2(n5926), .B1(n7559), .B2(n9559), .ZN(n7391)
         );
  INV_X1 U9127 ( .A(n7388), .ZN(n7389) );
  OAI211_X1 U9128 ( .C1(n7389), .C2(n10154), .A(n10094), .B(n7494), .ZN(n10152) );
  NOR2_X1 U9129 ( .A1(n10152), .A2(n10097), .ZN(n7390) );
  AOI211_X1 U9130 ( .C1(n10074), .C2(n7561), .A(n7391), .B(n7390), .ZN(n7392)
         );
  OAI211_X1 U9131 ( .C1(n10102), .C2(n10153), .A(n7393), .B(n7392), .ZN(
        P1_U3281) );
  XNOR2_X1 U9132 ( .A(n7395), .B(n7394), .ZN(n7396) );
  NAND2_X1 U9133 ( .A1(n7396), .A2(n8765), .ZN(n7398) );
  AOI22_X1 U9134 ( .A1(n8405), .A2(n8741), .B1(n5047), .B2(n8403), .ZN(n7397)
         );
  NAND2_X1 U9135 ( .A1(n7398), .A2(n7397), .ZN(n10276) );
  INV_X1 U9136 ( .A(n10276), .ZN(n7406) );
  NAND3_X1 U9137 ( .A1(n7472), .A2(n8086), .A3(n8080), .ZN(n7399) );
  NAND2_X1 U9138 ( .A1(n7400), .A2(n7399), .ZN(n10278) );
  INV_X1 U9139 ( .A(n7401), .ZN(n10275) );
  INV_X1 U9140 ( .A(n7402), .ZN(n7705) );
  AOI22_X1 U9141 ( .A1(n8725), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n8748), .B2(
        n7705), .ZN(n7403) );
  OAI21_X1 U9142 ( .B1(n10275), .B2(n8595), .A(n7403), .ZN(n7404) );
  AOI21_X1 U9143 ( .B1(n10278), .B2(n8619), .A(n7404), .ZN(n7405) );
  OAI21_X1 U9144 ( .B1(n7406), .B2(n8725), .A(n7405), .ZN(P2_U3222) );
  INV_X1 U9145 ( .A(n7407), .ZN(n7459) );
  OAI222_X1 U9146 ( .A1(n9969), .A2(n7459), .B1(P1_U3086), .B2(n7408), .C1(
        n9923), .C2(n9966), .ZN(P1_U3330) );
  NOR2_X1 U9147 ( .A1(n7424), .A2(n7409), .ZN(n7411) );
  INV_X1 U9148 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7412) );
  MUX2_X1 U9149 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n7412), .S(n7427), .Z(n7414)
         );
  INV_X1 U9150 ( .A(n8430), .ZN(n7413) );
  AOI21_X1 U9151 ( .B1(n7415), .B2(n7414), .A(n7413), .ZN(n7436) );
  NAND2_X1 U9152 ( .A1(n8551), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7416) );
  OAI21_X1 U9153 ( .B1(n8551), .B2(n7428), .A(n7416), .ZN(n8421) );
  XNOR2_X1 U9154 ( .A(n8421), .B(n7427), .ZN(n7422) );
  OR2_X1 U9155 ( .A1(n7418), .A2(n7417), .ZN(n7420) );
  NAND2_X1 U9156 ( .A1(n7420), .A2(n7419), .ZN(n7421) );
  NAND2_X1 U9157 ( .A1(n7422), .A2(n7421), .ZN(n8422) );
  OAI21_X1 U9158 ( .B1(n7422), .B2(n7421), .A(n8422), .ZN(n7434) );
  NAND2_X1 U9159 ( .A1(n10212), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n7423) );
  NAND2_X1 U9160 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3151), .ZN(n8306) );
  OAI211_X1 U9161 ( .C1(n10204), .C2(n8428), .A(n7423), .B(n8306), .ZN(n7433)
         );
  NOR2_X1 U9162 ( .A1(n7424), .A2(n4443), .ZN(n7426) );
  NOR2_X1 U9163 ( .A1(n7426), .A2(n7425), .ZN(n7430) );
  MUX2_X1 U9164 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n7428), .S(n7427), .Z(n7429)
         );
  NAND2_X1 U9165 ( .A1(n7430), .A2(n7429), .ZN(n7431) );
  AOI21_X1 U9166 ( .B1(n8417), .B2(n7431), .A(n10220), .ZN(n7432) );
  AOI211_X1 U9167 ( .C1(n10225), .C2(n7434), .A(n7433), .B(n7432), .ZN(n7435)
         );
  OAI21_X1 U9168 ( .B1(n7436), .B2(n10229), .A(n7435), .ZN(P2_U3194) );
  OAI22_X1 U9169 ( .A1(n7441), .A2(n4394), .B1(n7437), .B2(n8996), .ZN(n7438)
         );
  XNOR2_X1 U9170 ( .A(n7438), .B(n8997), .ZN(n7532) );
  XOR2_X1 U9171 ( .A(n7526), .B(n7532), .Z(n9089) );
  OR2_X1 U9172 ( .A1(n7441), .A2(n9065), .ZN(n7443) );
  NAND2_X1 U9173 ( .A1(n9564), .A2(n7541), .ZN(n7442) );
  NAND2_X1 U9174 ( .A1(n7443), .A2(n7442), .ZN(n7531) );
  INV_X1 U9175 ( .A(n7531), .ZN(n9088) );
  NAND2_X1 U9176 ( .A1(n9089), .A2(n9088), .ZN(n9087) );
  OAI21_X1 U9177 ( .B1(n7532), .B2(n7526), .A(n9087), .ZN(n7448) );
  NAND2_X1 U9178 ( .A1(n7455), .A2(n9070), .ZN(n7444) );
  OAI21_X1 U9179 ( .B1(n7445), .B2(n4394), .A(n7444), .ZN(n7446) );
  XNOR2_X1 U9180 ( .A(n7446), .B(n9068), .ZN(n7533) );
  AOI22_X1 U9181 ( .A1(n9223), .A2(n9002), .B1(n7541), .B2(n7455), .ZN(n7529)
         );
  XNOR2_X1 U9182 ( .A(n7533), .B(n7529), .ZN(n7447) );
  XNOR2_X1 U9183 ( .A(n7448), .B(n7447), .ZN(n7457) );
  OAI21_X1 U9184 ( .B1(n7450), .B2(n7449), .A(n9195), .ZN(n7452) );
  OAI211_X1 U9185 ( .C1(n9198), .C2(n7453), .A(n7452), .B(n7451), .ZN(n7454)
         );
  AOI21_X1 U9186 ( .B1(n7455), .B2(n9201), .A(n7454), .ZN(n7456) );
  OAI21_X1 U9187 ( .B1(n7457), .B2(n9204), .A(n7456), .ZN(P1_U3231) );
  OAI222_X1 U9188 ( .A1(P2_U3151), .A2(n5600), .B1(n8918), .B2(n7459), .C1(
        n7458), .C2(n8258), .ZN(P2_U3270) );
  AOI21_X1 U9189 ( .B1(n8390), .B2(n8407), .A(n7460), .ZN(n7464) );
  INV_X1 U9190 ( .A(n7461), .ZN(n7462) );
  NAND2_X1 U9191 ( .A1(n8394), .A2(n7462), .ZN(n7463) );
  OAI211_X1 U9192 ( .C1(n7701), .C2(n8392), .A(n7464), .B(n7463), .ZN(n7470)
         );
  INV_X1 U9193 ( .A(n7465), .ZN(n7466) );
  AOI211_X1 U9194 ( .C1(n7468), .C2(n7467), .A(n8381), .B(n7466), .ZN(n7469)
         );
  AOI211_X1 U9195 ( .C1(n10267), .C2(n8379), .A(n7470), .B(n7469), .ZN(n7471)
         );
  INV_X1 U9196 ( .A(n7471), .ZN(P2_U3171) );
  INV_X1 U9197 ( .A(n7472), .ZN(n7473) );
  AOI21_X1 U9198 ( .B1(n8223), .B2(n7474), .A(n7473), .ZN(n10269) );
  AOI22_X1 U9199 ( .A1(n8404), .A2(n5047), .B1(n8741), .B2(n8406), .ZN(n7478)
         );
  XNOR2_X1 U9200 ( .A(n7475), .B(n8223), .ZN(n7476) );
  NAND2_X1 U9201 ( .A1(n7476), .A2(n8765), .ZN(n7477) );
  OAI211_X1 U9202 ( .C1(n10269), .C2(n7479), .A(n7478), .B(n7477), .ZN(n10270)
         );
  NAND2_X1 U9203 ( .A1(n10270), .A2(n8745), .ZN(n7483) );
  OAI22_X1 U9204 ( .A1(n8745), .A2(n7480), .B1(n7677), .B2(n8771), .ZN(n7481)
         );
  AOI21_X1 U9205 ( .B1(n8749), .B2(n10272), .A(n7481), .ZN(n7482) );
  OAI211_X1 U9206 ( .C1(n10269), .C2(n7484), .A(n7483), .B(n7482), .ZN(
        P2_U3223) );
  NAND2_X1 U9207 ( .A1(n7485), .A2(n7870), .ZN(n7486) );
  NAND2_X1 U9208 ( .A1(n7486), .A2(n7970), .ZN(n7488) );
  NAND2_X1 U9209 ( .A1(n7488), .A2(n7487), .ZN(n7490) );
  OR2_X1 U9210 ( .A1(n7626), .A2(n9350), .ZN(n7489) );
  OAI21_X1 U9211 ( .B1(n7552), .B2(n9373), .A(n7489), .ZN(n7585) );
  AOI21_X1 U9212 ( .B1(n7490), .B2(n10072), .A(n7585), .ZN(n10158) );
  XNOR2_X1 U9213 ( .A(n7492), .B(n7491), .ZN(n10162) );
  NAND2_X1 U9214 ( .A1(n10162), .A2(n10082), .ZN(n7499) );
  OAI22_X1 U9215 ( .A1(n9562), .A2(n7493), .B1(n7587), .B2(n9559), .ZN(n7497)
         );
  INV_X1 U9216 ( .A(n7494), .ZN(n7495) );
  OAI211_X1 U9217 ( .C1(n7495), .C2(n4692), .A(n10094), .B(n7597), .ZN(n10157)
         );
  NOR2_X1 U9218 ( .A1(n10157), .A2(n10097), .ZN(n7496) );
  AOI211_X1 U9219 ( .C1(n10074), .C2(n7589), .A(n7497), .B(n7496), .ZN(n7498)
         );
  OAI211_X1 U9220 ( .C1(n10102), .C2(n10158), .A(n7499), .B(n7498), .ZN(
        P1_U3280) );
  INV_X1 U9221 ( .A(n7500), .ZN(n7523) );
  OAI222_X1 U9222 ( .A1(n9969), .A2(n7523), .B1(P1_U3086), .B2(n7502), .C1(
        n7501), .C2(n9966), .ZN(P1_U3329) );
  NAND2_X1 U9223 ( .A1(n7504), .A2(n7503), .ZN(n7506) );
  XOR2_X1 U9224 ( .A(n7506), .B(n7505), .Z(n7512) );
  OR2_X1 U9225 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9783), .ZN(n8426) );
  OAI21_X1 U9226 ( .B1(n8392), .B2(n7507), .A(n8426), .ZN(n7508) );
  AOI21_X1 U9227 ( .B1(n8390), .B2(n8403), .A(n7508), .ZN(n7509) );
  OAI21_X1 U9228 ( .B1(n7714), .B2(n8339), .A(n7509), .ZN(n7510) );
  AOI21_X1 U9229 ( .B1(n7713), .B2(n8379), .A(n7510), .ZN(n7511) );
  OAI21_X1 U9230 ( .B1(n7512), .B2(n8381), .A(n7511), .ZN(P2_U3174) );
  XNOR2_X1 U9231 ( .A(n7513), .B(n5633), .ZN(n7515) );
  OAI22_X1 U9232 ( .A1(n8308), .A2(n8762), .B1(n8303), .B2(n8761), .ZN(n7514)
         );
  AOI21_X1 U9233 ( .B1(n7515), .B2(n8765), .A(n7514), .ZN(n10284) );
  NAND2_X1 U9234 ( .A1(n7516), .A2(n8087), .ZN(n7517) );
  AND2_X1 U9235 ( .A1(n7518), .A2(n7517), .ZN(n10280) );
  NAND2_X1 U9236 ( .A1(n10280), .A2(n8619), .ZN(n7521) );
  OAI22_X1 U9237 ( .A1(n8745), .A2(n7428), .B1(n8312), .B2(n8771), .ZN(n7519)
         );
  AOI21_X1 U9238 ( .B1(n8749), .B2(n10282), .A(n7519), .ZN(n7520) );
  OAI211_X1 U9239 ( .C1(n10284), .C2(n8725), .A(n7521), .B(n7520), .ZN(
        P2_U3221) );
  OAI222_X1 U9240 ( .A1(P2_U3151), .A2(n7524), .B1(n8918), .B2(n7523), .C1(
        n7522), .C2(n8258), .ZN(P2_U3269) );
  NOR2_X1 U9241 ( .A1(n7533), .A2(n7529), .ZN(n7528) );
  AND2_X1 U9242 ( .A1(n7532), .A2(n7531), .ZN(n7527) );
  INV_X1 U9243 ( .A(n7529), .ZN(n7530) );
  OAI21_X1 U9244 ( .B1(n7532), .B2(n7531), .A(n7530), .ZN(n7534) );
  OAI22_X1 U9245 ( .A1(n10146), .A2(n8996), .B1(n7537), .B2(n4394), .ZN(n7536)
         );
  XNOR2_X1 U9246 ( .A(n7536), .B(n9068), .ZN(n7653) );
  OAI22_X1 U9247 ( .A1(n10146), .A2(n4394), .B1(n7537), .B2(n9065), .ZN(n7652)
         );
  INV_X1 U9248 ( .A(n7652), .ZN(n7545) );
  NAND2_X1 U9249 ( .A1(n9049), .A2(n9070), .ZN(n7539) );
  OR2_X1 U9250 ( .A1(n7542), .A2(n4394), .ZN(n7538) );
  NAND2_X1 U9251 ( .A1(n7539), .A2(n7538), .ZN(n7540) );
  XNOR2_X1 U9252 ( .A(n7540), .B(n8997), .ZN(n7650) );
  INV_X1 U9253 ( .A(n7650), .ZN(n7649) );
  NAND2_X1 U9254 ( .A1(n9049), .A2(n7541), .ZN(n7544) );
  OR2_X1 U9255 ( .A1(n7542), .A2(n9065), .ZN(n7543) );
  NAND2_X1 U9256 ( .A1(n7544), .A2(n7543), .ZN(n7546) );
  INV_X1 U9257 ( .A(n7546), .ZN(n9046) );
  OAI22_X1 U9258 ( .A1(n7653), .A2(n7545), .B1(n7649), .B2(n9046), .ZN(n7550)
         );
  OAI21_X1 U9259 ( .B1(n7650), .B2(n7546), .A(n7652), .ZN(n7548) );
  NOR3_X1 U9260 ( .A1(n7652), .A2(n7650), .A3(n7546), .ZN(n7547) );
  AOI21_X1 U9261 ( .B1(n7653), .B2(n7548), .A(n7547), .ZN(n7549) );
  OAI22_X1 U9262 ( .A1(n10154), .A2(n4394), .B1(n7552), .B2(n9065), .ZN(n7576)
         );
  NAND2_X1 U9263 ( .A1(n7561), .A2(n9070), .ZN(n7554) );
  INV_X1 U9264 ( .A(n7552), .ZN(n9220) );
  NAND2_X1 U9265 ( .A1(n9220), .A2(n7541), .ZN(n7553) );
  NAND2_X1 U9266 ( .A1(n7554), .A2(n7553), .ZN(n7555) );
  XNOR2_X1 U9267 ( .A(n7555), .B(n8997), .ZN(n7577) );
  XOR2_X1 U9268 ( .A(n7576), .B(n7577), .Z(n7580) );
  XOR2_X1 U9269 ( .A(n7581), .B(n7580), .Z(n7563) );
  AOI21_X1 U9270 ( .B1(n7557), .B2(n9195), .A(n7556), .ZN(n7558) );
  OAI21_X1 U9271 ( .B1(n7559), .B2(n9198), .A(n7558), .ZN(n7560) );
  AOI21_X1 U9272 ( .B1(n7561), .B2(n9201), .A(n7560), .ZN(n7562) );
  OAI21_X1 U9273 ( .B1(n7563), .B2(n9204), .A(n7562), .ZN(P1_U3224) );
  INV_X1 U9274 ( .A(n7564), .ZN(n7636) );
  AOI21_X1 U9275 ( .B1(n8916), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n7565), .ZN(
        n7566) );
  OAI21_X1 U9276 ( .B1(n7636), .B2(n7567), .A(n7566), .ZN(P2_U3268) );
  XOR2_X1 U9277 ( .A(n7568), .B(n7569), .Z(n7575) );
  NAND2_X1 U9278 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8450) );
  OAI21_X1 U9279 ( .B1(n8392), .B2(n7570), .A(n8450), .ZN(n7571) );
  AOI21_X1 U9280 ( .B1(n8390), .B2(n8402), .A(n7571), .ZN(n7572) );
  OAI21_X1 U9281 ( .B1(n7726), .B2(n8339), .A(n7572), .ZN(n7573) );
  AOI21_X1 U9282 ( .B1(n7736), .B2(n8379), .A(n7573), .ZN(n7574) );
  OAI21_X1 U9283 ( .B1(n7575), .B2(n8381), .A(n7574), .ZN(P2_U3155) );
  INV_X1 U9284 ( .A(n7576), .ZN(n7579) );
  INV_X1 U9285 ( .A(n7577), .ZN(n7578) );
  AOI22_X2 U9286 ( .A1(n7581), .A2(n7580), .B1(n7579), .B2(n7578), .ZN(n7611)
         );
  AOI22_X1 U9287 ( .A1(n7589), .A2(n7541), .B1(n9002), .B2(n9219), .ZN(n7606)
         );
  NAND2_X1 U9288 ( .A1(n7589), .A2(n9070), .ZN(n7583) );
  NAND2_X1 U9289 ( .A1(n9219), .A2(n7541), .ZN(n7582) );
  NAND2_X1 U9290 ( .A1(n7583), .A2(n7582), .ZN(n7584) );
  XNOR2_X1 U9291 ( .A(n7584), .B(n8997), .ZN(n7608) );
  XOR2_X1 U9292 ( .A(n7606), .B(n7608), .Z(n7610) );
  XOR2_X1 U9293 ( .A(n7611), .B(n7610), .Z(n7591) );
  AOI22_X1 U9294 ( .A1(n7585), .A2(n9195), .B1(P1_REG3_REG_13__SCAN_IN), .B2(
        P1_U3086), .ZN(n7586) );
  OAI21_X1 U9295 ( .B1(n7587), .B2(n9198), .A(n7586), .ZN(n7588) );
  AOI21_X1 U9296 ( .B1(n7589), .B2(n9201), .A(n7588), .ZN(n7590) );
  OAI21_X1 U9297 ( .B1(n7591), .B2(n9204), .A(n7590), .ZN(P1_U3234) );
  AOI21_X1 U9298 ( .B1(n7592), .B2(n7971), .A(n10087), .ZN(n7595) );
  OR2_X1 U9299 ( .A1(n8920), .A2(n9350), .ZN(n7593) );
  OAI21_X1 U9300 ( .B1(n7594), .B2(n9373), .A(n7593), .ZN(n7615) );
  AOI21_X1 U9301 ( .B1(n7595), .B2(n7621), .A(n7615), .ZN(n10167) );
  XOR2_X1 U9302 ( .A(n7596), .B(n7971), .Z(n10169) );
  INV_X1 U9303 ( .A(n10169), .ZN(n10171) );
  NAND2_X1 U9304 ( .A1(n10171), .A2(n10082), .ZN(n7602) );
  AOI211_X1 U9305 ( .C1(n10164), .C2(n7597), .A(n9540), .B(n7630), .ZN(n10163)
         );
  NOR2_X1 U9306 ( .A1(n7613), .A2(n10096), .ZN(n7600) );
  OAI22_X1 U9307 ( .A1(n9562), .A2(n7598), .B1(n7617), .B2(n9559), .ZN(n7599)
         );
  AOI211_X1 U9308 ( .C1(n10163), .C2(n10081), .A(n7600), .B(n7599), .ZN(n7601)
         );
  OAI211_X1 U9309 ( .C1(n10102), .C2(n10167), .A(n7602), .B(n7601), .ZN(
        P1_U3279) );
  INV_X1 U9310 ( .A(n7603), .ZN(n7638) );
  AOI21_X1 U9311 ( .B1(n8916), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n7604), .ZN(
        n7605) );
  OAI21_X1 U9312 ( .B1(n7638), .B2(n8918), .A(n7605), .ZN(P2_U3267) );
  INV_X1 U9313 ( .A(n7606), .ZN(n7607) );
  OAI21_X2 U9314 ( .B1(n7611), .B2(n7610), .A(n7609), .ZN(n8926) );
  OAI22_X1 U9315 ( .A1(n7613), .A2(n8996), .B1(n7626), .B2(n4394), .ZN(n7612)
         );
  XOR2_X1 U9316 ( .A(n8997), .B(n7612), .Z(n8925) );
  INV_X1 U9317 ( .A(n8925), .ZN(n8927) );
  OAI22_X1 U9318 ( .A1(n7613), .A2(n4394), .B1(n7626), .B2(n9065), .ZN(n8929)
         );
  XNOR2_X1 U9319 ( .A(n8927), .B(n8929), .ZN(n7614) );
  XNOR2_X1 U9320 ( .A(n8926), .B(n7614), .ZN(n7620) );
  AOI22_X1 U9321 ( .A1(n7615), .A2(n9195), .B1(P1_REG3_REG_14__SCAN_IN), .B2(
        P1_U3086), .ZN(n7616) );
  OAI21_X1 U9322 ( .B1(n7617), .B2(n9198), .A(n7616), .ZN(n7618) );
  AOI21_X1 U9323 ( .B1(n10164), .B2(n9201), .A(n7618), .ZN(n7619) );
  OAI21_X1 U9324 ( .B1(n7620), .B2(n9204), .A(n7619), .ZN(P1_U3215) );
  NAND2_X1 U9325 ( .A1(n7621), .A2(n7774), .ZN(n7622) );
  NAND2_X1 U9326 ( .A1(n7622), .A2(n7879), .ZN(n7624) );
  NAND2_X1 U9327 ( .A1(n7624), .A2(n7623), .ZN(n7627) );
  OR2_X1 U9328 ( .A1(n9132), .A2(n9350), .ZN(n7625) );
  OAI21_X1 U9329 ( .B1(n7626), .B2(n9373), .A(n7625), .ZN(n9196) );
  AOI21_X1 U9330 ( .B1(n7627), .B2(n10072), .A(n9196), .ZN(n10027) );
  XNOR2_X1 U9331 ( .A(n7628), .B(n7973), .ZN(n10029) );
  NAND2_X1 U9332 ( .A1(n10029), .A2(n10082), .ZN(n7634) );
  OAI22_X1 U9333 ( .A1(n9562), .A2(n7629), .B1(n9199), .B2(n9559), .ZN(n7632)
         );
  OAI211_X1 U9334 ( .C1(n7630), .C2(n4656), .A(n7693), .B(n10094), .ZN(n10026)
         );
  NOR2_X1 U9335 ( .A1(n10026), .A2(n10097), .ZN(n7631) );
  AOI211_X1 U9336 ( .C1(n10074), .C2(n9202), .A(n7632), .B(n7631), .ZN(n7633)
         );
  OAI211_X1 U9337 ( .C1(n10102), .C2(n10027), .A(n7634), .B(n7633), .ZN(
        P1_U3278) );
  OAI222_X1 U9338 ( .A1(n9969), .A2(n7636), .B1(P1_U3086), .B2(n6372), .C1(
        n7635), .C2(n9966), .ZN(P1_U3328) );
  OAI222_X1 U9339 ( .A1(n9969), .A2(n7638), .B1(n9246), .B2(P1_U3086), .C1(
        n7637), .C2(n9966), .ZN(P1_U3327) );
  OAI211_X1 U9340 ( .C1(n7641), .C2(n7640), .A(n7639), .B(n8387), .ZN(n7647)
         );
  INV_X1 U9341 ( .A(n7642), .ZN(n8747) );
  NAND2_X1 U9342 ( .A1(n8390), .A2(n8742), .ZN(n7643) );
  NAND2_X1 U9343 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8472) );
  OAI211_X1 U9344 ( .C1(n7644), .C2(n8392), .A(n7643), .B(n8472), .ZN(n7645)
         );
  AOI21_X1 U9345 ( .B1(n8747), .B2(n8394), .A(n7645), .ZN(n7646) );
  OAI211_X1 U9346 ( .C1(n7648), .C2(n8397), .A(n7647), .B(n7646), .ZN(P2_U3181) );
  XNOR2_X1 U9347 ( .A(n7651), .B(n7649), .ZN(n9045) );
  NAND2_X1 U9348 ( .A1(n9045), .A2(n9046), .ZN(n9044) );
  OAI21_X1 U9349 ( .B1(n7651), .B2(n7650), .A(n9044), .ZN(n7655) );
  XNOR2_X1 U9350 ( .A(n7653), .B(n7652), .ZN(n7654) );
  XNOR2_X1 U9351 ( .A(n7655), .B(n7654), .ZN(n7663) );
  NOR2_X1 U9352 ( .A1(n10146), .A2(n9191), .ZN(n7662) );
  NAND2_X1 U9353 ( .A1(n7656), .A2(n9195), .ZN(n7659) );
  INV_X1 U9354 ( .A(n7657), .ZN(n7658) );
  OAI211_X1 U9355 ( .C1(n9198), .C2(n7660), .A(n7659), .B(n7658), .ZN(n7661)
         );
  AOI211_X1 U9356 ( .C1(n7663), .C2(n9184), .A(n7662), .B(n7661), .ZN(n7664)
         );
  INV_X1 U9357 ( .A(n7664), .ZN(P1_U3236) );
  INV_X1 U9358 ( .A(n7666), .ZN(n7667) );
  OR2_X1 U9359 ( .A1(n7668), .A2(n7667), .ZN(n8225) );
  XNOR2_X1 U9360 ( .A(n7665), .B(n8225), .ZN(n7720) );
  INV_X1 U9361 ( .A(n8225), .ZN(n8088) );
  XNOR2_X1 U9362 ( .A(n7669), .B(n8088), .ZN(n7670) );
  AOI222_X1 U9363 ( .A1(n8765), .A2(n7670), .B1(n8742), .B2(n5047), .C1(n8403), 
        .C2(n8741), .ZN(n7712) );
  MUX2_X1 U9364 ( .A(n9752), .B(n7712), .S(n10303), .Z(n7672) );
  NAND2_X1 U9365 ( .A1(n7713), .A2(n8826), .ZN(n7671) );
  OAI211_X1 U9366 ( .C1(n8829), .C2(n7720), .A(n7672), .B(n7671), .ZN(P2_U3472) );
  INV_X1 U9367 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7673) );
  MUX2_X1 U9368 ( .A(n7673), .B(n7712), .S(n10286), .Z(n7675) );
  NAND2_X1 U9369 ( .A1(n7713), .A2(n5698), .ZN(n7674) );
  OAI211_X1 U9370 ( .C1(n7720), .C2(n8910), .A(n7675), .B(n7674), .ZN(P2_U3429) );
  AOI21_X1 U9371 ( .B1(n8390), .B2(n8406), .A(n7676), .ZN(n7680) );
  INV_X1 U9372 ( .A(n7677), .ZN(n7678) );
  NAND2_X1 U9373 ( .A1(n8394), .A2(n7678), .ZN(n7679) );
  OAI211_X1 U9374 ( .C1(n8303), .C2(n8392), .A(n7680), .B(n7679), .ZN(n7686)
         );
  INV_X1 U9375 ( .A(n7681), .ZN(n7683) );
  XNOR2_X1 U9376 ( .A(n7699), .B(n8405), .ZN(n7682) );
  NOR2_X1 U9377 ( .A1(n7682), .A2(n7683), .ZN(n7700) );
  AOI21_X1 U9378 ( .B1(n7683), .B2(n7682), .A(n7700), .ZN(n7684) );
  NOR2_X1 U9379 ( .A1(n7684), .A2(n8381), .ZN(n7685) );
  AOI211_X1 U9380 ( .C1(n10272), .C2(n8379), .A(n7686), .B(n7685), .ZN(n7687)
         );
  INV_X1 U9381 ( .A(n7687), .ZN(P2_U3157) );
  XNOR2_X1 U9382 ( .A(n7688), .B(n7974), .ZN(n7690) );
  NAND2_X1 U9383 ( .A1(n9217), .A2(n9150), .ZN(n7689) );
  OAI21_X1 U9384 ( .B1(n8920), .B2(n9373), .A(n7689), .ZN(n9122) );
  AOI21_X1 U9385 ( .B1(n7690), .B2(n10072), .A(n9122), .ZN(n9642) );
  AOI21_X1 U9386 ( .B1(n7974), .B2(n7691), .A(n4473), .ZN(n9644) );
  NAND2_X1 U9387 ( .A1(n9644), .A2(n10082), .ZN(n7698) );
  OAI22_X1 U9388 ( .A1(n9562), .A2(n7692), .B1(n9124), .B2(n9559), .ZN(n7696)
         );
  INV_X1 U9389 ( .A(n9126), .ZN(n9957) );
  INV_X1 U9390 ( .A(n7693), .ZN(n7694) );
  OAI211_X1 U9391 ( .C1(n9957), .C2(n7694), .A(n4978), .B(n10094), .ZN(n9641)
         );
  NOR2_X1 U9392 ( .A1(n9641), .A2(n10097), .ZN(n7695) );
  AOI211_X1 U9393 ( .C1(n10074), .C2(n9126), .A(n7696), .B(n7695), .ZN(n7697)
         );
  OAI211_X1 U9394 ( .C1(n10102), .C2(n9642), .A(n7698), .B(n7697), .ZN(
        P1_U3277) );
  INV_X1 U9395 ( .A(n7699), .ZN(n7702) );
  AOI21_X1 U9396 ( .B1(n7702), .B2(n7701), .A(n7700), .ZN(n7703) );
  NAND2_X1 U9397 ( .A1(n7703), .A2(n8302), .ZN(n8301) );
  OAI211_X1 U9398 ( .C1(n7703), .C2(n8302), .A(n8301), .B(n8387), .ZN(n7711)
         );
  AOI21_X1 U9399 ( .B1(n8390), .B2(n8405), .A(n7704), .ZN(n7707) );
  NAND2_X1 U9400 ( .A1(n8394), .A2(n7705), .ZN(n7706) );
  OAI211_X1 U9401 ( .C1(n7708), .C2(n8392), .A(n7707), .B(n7706), .ZN(n7709)
         );
  INV_X1 U9402 ( .A(n7709), .ZN(n7710) );
  OAI211_X1 U9403 ( .C1(n10275), .C2(n8397), .A(n7711), .B(n7710), .ZN(
        P2_U3176) );
  INV_X1 U9404 ( .A(n7712), .ZN(n7717) );
  INV_X1 U9405 ( .A(n7713), .ZN(n7715) );
  OAI22_X1 U9406 ( .A1(n7715), .A2(n8632), .B1(n7714), .B2(n8771), .ZN(n7716)
         );
  OAI21_X1 U9407 ( .B1(n7717), .B2(n7716), .A(n8745), .ZN(n7719) );
  NAND2_X1 U9408 ( .A1(n8725), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7718) );
  OAI211_X1 U9409 ( .C1(n7720), .C2(n8752), .A(n7719), .B(n7718), .ZN(P2_U3220) );
  NAND2_X1 U9410 ( .A1(n8097), .A2(n8096), .ZN(n8093) );
  XNOR2_X1 U9411 ( .A(n7721), .B(n8093), .ZN(n7739) );
  INV_X1 U9412 ( .A(n8093), .ZN(n8227) );
  XNOR2_X1 U9413 ( .A(n7722), .B(n8227), .ZN(n7723) );
  NAND2_X1 U9414 ( .A1(n7723), .A2(n8765), .ZN(n7725) );
  AOI22_X1 U9415 ( .A1(n8402), .A2(n8741), .B1(n5047), .B2(n8730), .ZN(n7724)
         );
  INV_X1 U9416 ( .A(n7734), .ZN(n7729) );
  INV_X1 U9417 ( .A(n7736), .ZN(n7727) );
  OAI22_X1 U9418 ( .A1(n7727), .A2(n8632), .B1(n7726), .B2(n8771), .ZN(n7728)
         );
  OAI21_X1 U9419 ( .B1(n7729), .B2(n7728), .A(n8745), .ZN(n7731) );
  NAND2_X1 U9420 ( .A1(n8725), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7730) );
  OAI211_X1 U9421 ( .C1(n7739), .C2(n8752), .A(n7731), .B(n7730), .ZN(P2_U3219) );
  MUX2_X1 U9422 ( .A(n8440), .B(n7734), .S(n10303), .Z(n7733) );
  NAND2_X1 U9423 ( .A1(n7736), .A2(n8826), .ZN(n7732) );
  OAI211_X1 U9424 ( .C1(n8829), .C2(n7739), .A(n7733), .B(n7732), .ZN(P2_U3473) );
  INV_X1 U9425 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7735) );
  MUX2_X1 U9426 ( .A(n7735), .B(n7734), .S(n10286), .Z(n7738) );
  NAND2_X1 U9427 ( .A1(n7736), .A2(n5698), .ZN(n7737) );
  OAI211_X1 U9428 ( .C1(n7739), .C2(n8910), .A(n7738), .B(n7737), .ZN(P2_U3432) );
  NAND2_X1 U9429 ( .A1(n7742), .A2(n7741), .ZN(n7743) );
  INV_X1 U9430 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n7799) );
  INV_X1 U9431 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9755) );
  MUX2_X1 U9432 ( .A(n7799), .B(n9755), .S(n7813), .Z(n7810) );
  XNOR2_X1 U9433 ( .A(n7810), .B(SI_30_), .ZN(n7807) );
  INV_X1 U9434 ( .A(n8161), .ZN(n8259) );
  OAI222_X1 U9435 ( .A1(n9969), .A2(n8259), .B1(n7744), .B2(P1_U3086), .C1(
        n7799), .C2(n9966), .ZN(P1_U3325) );
  INV_X1 U9436 ( .A(n7747), .ZN(n9968) );
  OAI222_X1 U9437 ( .A1(n8258), .A2(n7746), .B1(n8918), .B2(n9968), .C1(n7745), 
        .C2(P2_U3151), .ZN(P2_U3266) );
  INV_X1 U9438 ( .A(n7937), .ZN(n7748) );
  NOR2_X1 U9439 ( .A1(n7945), .A2(n7748), .ZN(n7991) );
  OR2_X1 U9440 ( .A1(n9590), .A2(n7749), .ZN(n7750) );
  NAND2_X1 U9441 ( .A1(n7751), .A2(n7750), .ZN(n7942) );
  NAND2_X1 U9442 ( .A1(n7929), .A2(n9435), .ZN(n7791) );
  AND2_X1 U9443 ( .A1(n7925), .A2(n7922), .ZN(n7752) );
  OAI211_X1 U9444 ( .C1(n7791), .C2(n7752), .A(n9417), .B(n7940), .ZN(n7793)
         );
  OR2_X1 U9445 ( .A1(n7942), .A2(n7793), .ZN(n7990) );
  NAND2_X1 U9446 ( .A1(n7788), .A2(n9494), .ZN(n7911) );
  INV_X1 U9447 ( .A(n7911), .ZN(n7987) );
  OR2_X1 U9448 ( .A1(n9531), .A2(n7753), .ZN(n7783) );
  NOR2_X1 U9449 ( .A1(n9636), .A2(n8941), .ZN(n7904) );
  INV_X1 U9450 ( .A(n7904), .ZN(n7754) );
  NAND2_X1 U9451 ( .A1(n7783), .A2(n7754), .ZN(n7918) );
  INV_X1 U9452 ( .A(n7918), .ZN(n7782) );
  NAND2_X1 U9453 ( .A1(n7834), .A2(n7830), .ZN(n7828) );
  INV_X1 U9454 ( .A(n7755), .ZN(n7758) );
  NAND2_X1 U9455 ( .A1(n9230), .A2(n6106), .ZN(n7756) );
  AND4_X1 U9456 ( .A1(n6112), .A2(n7758), .A3(n7757), .A4(n7756), .ZN(n7759)
         );
  OAI211_X1 U9457 ( .C1(n7828), .C2(n7759), .A(n7836), .B(n7829), .ZN(n7762)
         );
  INV_X1 U9458 ( .A(n7760), .ZN(n7761) );
  AOI21_X1 U9459 ( .B1(n7762), .B2(n7844), .A(n7761), .ZN(n7768) );
  INV_X1 U9460 ( .A(n7763), .ZN(n7767) );
  NAND2_X1 U9461 ( .A1(n7870), .A2(n7866), .ZN(n7770) );
  INV_X1 U9462 ( .A(n7865), .ZN(n7764) );
  OR2_X1 U9463 ( .A1(n7770), .A2(n7764), .ZN(n7873) );
  INV_X1 U9464 ( .A(n7873), .ZN(n7766) );
  OAI211_X1 U9465 ( .C1(n7768), .C2(n7767), .A(n7766), .B(n7765), .ZN(n7773)
         );
  INV_X1 U9466 ( .A(n7863), .ZN(n7769) );
  OR2_X1 U9467 ( .A1(n7770), .A2(n4509), .ZN(n7771) );
  NAND2_X1 U9468 ( .A1(n7771), .A2(n7868), .ZN(n7876) );
  INV_X1 U9469 ( .A(n7876), .ZN(n7772) );
  NAND3_X1 U9470 ( .A1(n7773), .A2(n7772), .A3(n7880), .ZN(n7775) );
  NAND3_X1 U9471 ( .A1(n7775), .A2(n7774), .A3(n7882), .ZN(n7777) );
  AND2_X1 U9472 ( .A1(n7891), .A2(n7776), .ZN(n7883) );
  NAND2_X1 U9473 ( .A1(n7777), .A2(n7883), .ZN(n7778) );
  NAND3_X1 U9474 ( .A1(n7778), .A2(n7893), .A3(n7897), .ZN(n7779) );
  NAND2_X1 U9475 ( .A1(n7779), .A2(n9547), .ZN(n7781) );
  AND2_X1 U9476 ( .A1(n7916), .A2(n7898), .ZN(n7903) );
  INV_X1 U9477 ( .A(n7903), .ZN(n7780) );
  AOI21_X1 U9478 ( .B1(n7782), .B2(n7781), .A(n7780), .ZN(n7785) );
  AND2_X1 U9479 ( .A1(n7920), .A2(n7783), .ZN(n7907) );
  INV_X1 U9480 ( .A(n7907), .ZN(n7784) );
  OAI21_X1 U9481 ( .B1(n7785), .B2(n7784), .A(n7917), .ZN(n7786) );
  NAND2_X1 U9482 ( .A1(n7987), .A2(n7786), .ZN(n7798) );
  INV_X1 U9483 ( .A(n7906), .ZN(n7787) );
  NAND2_X1 U9484 ( .A1(n7909), .A2(n7787), .ZN(n7789) );
  NAND2_X1 U9485 ( .A1(n7789), .A2(n7788), .ZN(n7790) );
  NAND2_X1 U9486 ( .A1(n7910), .A2(n7790), .ZN(n7923) );
  NOR2_X1 U9487 ( .A1(n7791), .A2(n7923), .ZN(n7792) );
  NOR2_X1 U9488 ( .A1(n7793), .A2(n7792), .ZN(n7796) );
  NAND2_X1 U9489 ( .A1(n7795), .A2(n7794), .ZN(n7939) );
  NOR2_X1 U9490 ( .A1(n7796), .A2(n7939), .ZN(n7797) );
  OR2_X1 U9491 ( .A1(n7942), .A2(n7797), .ZN(n7988) );
  OAI211_X1 U9492 ( .C1(n7990), .C2(n7798), .A(n7986), .B(n7988), .ZN(n7806)
         );
  NAND2_X1 U9493 ( .A1(n8161), .A2(n7818), .ZN(n7801) );
  OR2_X1 U9494 ( .A1(n7820), .A2(n7799), .ZN(n7800) );
  INV_X1 U9495 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9357) );
  OR2_X1 U9496 ( .A1(n4979), .A2(n9357), .ZN(n7804) );
  INV_X1 U9497 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9576) );
  OR2_X1 U9498 ( .A1(n5790), .A2(n9576), .ZN(n7803) );
  INV_X1 U9499 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9651) );
  OR2_X1 U9500 ( .A1(n6072), .A2(n9651), .ZN(n7802) );
  INV_X1 U9501 ( .A(n9374), .ZN(n9206) );
  NOR2_X1 U9502 ( .A1(n9653), .A2(n9206), .ZN(n7981) );
  NOR2_X1 U9503 ( .A1(n7981), .A2(n7944), .ZN(n7995) );
  INV_X1 U9504 ( .A(n7995), .ZN(n7805) );
  AOI21_X1 U9505 ( .B1(n7991), .B2(n7806), .A(n7805), .ZN(n7826) );
  NAND2_X1 U9506 ( .A1(n7808), .A2(n7807), .ZN(n7812) );
  INV_X1 U9507 ( .A(SI_30_), .ZN(n7809) );
  NAND2_X1 U9508 ( .A1(n7810), .A2(n7809), .ZN(n7811) );
  INV_X1 U9509 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n7819) );
  INV_X1 U9510 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n7814) );
  MUX2_X1 U9511 ( .A(n7819), .B(n7814), .S(n7813), .Z(n7815) );
  XNOR2_X1 U9512 ( .A(n7815), .B(SI_31_), .ZN(n7816) );
  OR2_X1 U9513 ( .A1(n7820), .A2(n7819), .ZN(n7821) );
  INV_X1 U9514 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9926) );
  INV_X1 U9515 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n7822) );
  OR2_X1 U9516 ( .A1(n4979), .A2(n7822), .ZN(n7824) );
  INV_X1 U9517 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9572) );
  OR2_X1 U9518 ( .A1(n5790), .A2(n9572), .ZN(n7823) );
  OAI211_X1 U9519 ( .C1(n6072), .C2(n9926), .A(n7824), .B(n7823), .ZN(n9353)
         );
  INV_X1 U9520 ( .A(n8006), .ZN(n7825) );
  OAI21_X1 U9521 ( .B1(n9374), .B2(n9360), .A(n7825), .ZN(n7983) );
  OAI21_X1 U9522 ( .B1(n7826), .B2(n7983), .A(n4534), .ZN(n8011) );
  INV_X1 U9523 ( .A(n7829), .ZN(n7833) );
  AND3_X1 U9524 ( .A1(n7831), .A2(n7830), .A3(n7950), .ZN(n7832) );
  OAI21_X1 U9525 ( .B1(n7834), .B2(n7833), .A(n7832), .ZN(n7835) );
  AOI21_X1 U9526 ( .B1(n7847), .B2(n7838), .A(n7837), .ZN(n7843) );
  OR2_X1 U9527 ( .A1(n7840), .A2(n7839), .ZN(n7842) );
  OAI22_X1 U9528 ( .A1(n7843), .A2(n7842), .B1(n7841), .B2(n7950), .ZN(n7856)
         );
  INV_X1 U9529 ( .A(n7844), .ZN(n7846) );
  OAI21_X1 U9530 ( .B1(n7847), .B2(n7846), .A(n7845), .ZN(n7849) );
  NAND3_X1 U9531 ( .A1(n7849), .A2(n7848), .A3(n7947), .ZN(n7855) );
  NAND2_X1 U9532 ( .A1(n7851), .A2(n7850), .ZN(n7852) );
  MUX2_X1 U9533 ( .A(n7853), .B(n7852), .S(n7950), .Z(n7854) );
  AOI21_X1 U9534 ( .B1(n7856), .B2(n7855), .A(n7854), .ZN(n7861) );
  NAND2_X1 U9535 ( .A1(n7874), .A2(n7857), .ZN(n7858) );
  MUX2_X1 U9536 ( .A(n7859), .B(n7858), .S(n7950), .Z(n7860) );
  OR2_X1 U9537 ( .A1(n7861), .A2(n7860), .ZN(n7875) );
  NAND2_X1 U9538 ( .A1(n7875), .A2(n7862), .ZN(n7864) );
  NAND3_X1 U9539 ( .A1(n7869), .A2(n7868), .A3(n4810), .ZN(n7871) );
  NAND2_X1 U9540 ( .A1(n7871), .A2(n7870), .ZN(n7872) );
  AOI21_X1 U9541 ( .B1(n7875), .B2(n7874), .A(n7873), .ZN(n7877) );
  OAI211_X1 U9542 ( .C1(n7877), .C2(n7876), .A(n7947), .B(n7882), .ZN(n7889)
         );
  NAND2_X1 U9543 ( .A1(n7893), .A2(n7950), .ZN(n7878) );
  NAND2_X1 U9544 ( .A1(n7879), .A2(n7878), .ZN(n7888) );
  OR2_X1 U9545 ( .A1(n7880), .A2(n7950), .ZN(n7881) );
  OAI21_X1 U9546 ( .B1(n7882), .B2(n7947), .A(n7881), .ZN(n7886) );
  INV_X1 U9547 ( .A(n7883), .ZN(n7884) );
  NAND2_X1 U9548 ( .A1(n7884), .A2(n7950), .ZN(n7885) );
  OAI21_X1 U9549 ( .B1(n7886), .B2(n7971), .A(n7885), .ZN(n7887) );
  NAND3_X1 U9550 ( .A1(n7891), .A2(n7890), .A3(n7947), .ZN(n7892) );
  OAI21_X1 U9551 ( .B1(n7893), .B2(n7950), .A(n7892), .ZN(n7894) );
  INV_X1 U9552 ( .A(n7894), .ZN(n7896) );
  INV_X1 U9553 ( .A(n7974), .ZN(n7895) );
  INV_X1 U9554 ( .A(n7897), .ZN(n7900) );
  NAND2_X1 U9555 ( .A1(n7898), .A2(n9547), .ZN(n7899) );
  MUX2_X1 U9556 ( .A(n7900), .B(n7899), .S(n7950), .Z(n7901) );
  OR2_X1 U9557 ( .A1(n7902), .A2(n7901), .ZN(n7915) );
  INV_X1 U9558 ( .A(n7917), .ZN(n7905) );
  AOI211_X1 U9559 ( .C1(n7908), .C2(n7907), .A(n7906), .B(n7905), .ZN(n7912)
         );
  OAI211_X1 U9560 ( .C1(n7912), .C2(n7911), .A(n7910), .B(n7909), .ZN(n7913)
         );
  INV_X1 U9561 ( .A(n7915), .ZN(n7919) );
  OAI211_X1 U9562 ( .C1(n7919), .C2(n7918), .A(n7917), .B(n7916), .ZN(n7921)
         );
  AND3_X1 U9563 ( .A1(n7921), .A2(n7987), .A3(n7920), .ZN(n7924) );
  OAI21_X1 U9564 ( .B1(n7924), .B2(n7923), .A(n7922), .ZN(n7927) );
  INV_X1 U9565 ( .A(n7925), .ZN(n7926) );
  INV_X1 U9566 ( .A(n9436), .ZN(n7933) );
  INV_X1 U9567 ( .A(n7929), .ZN(n7930) );
  MUX2_X1 U9568 ( .A(n7931), .B(n7930), .S(n7950), .Z(n7932) );
  AOI21_X1 U9569 ( .B1(n7938), .B2(n7940), .A(n7939), .ZN(n7935) );
  AOI21_X1 U9570 ( .B1(n7941), .B2(n7940), .A(n7939), .ZN(n7943) );
  MUX2_X1 U9571 ( .A(n7945), .B(n7944), .S(n7950), .Z(n7946) );
  INV_X1 U9572 ( .A(n9353), .ZN(n7948) );
  NOR2_X1 U9573 ( .A1(n7948), .A2(n9374), .ZN(n7985) );
  INV_X1 U9574 ( .A(n9368), .ZN(n7980) );
  INV_X1 U9575 ( .A(n9060), .ZN(n9214) );
  XNOR2_X1 U9576 ( .A(n9946), .B(n9214), .ZN(n9501) );
  INV_X1 U9577 ( .A(n10076), .ZN(n7953) );
  NAND4_X1 U9578 ( .A1(n7955), .A2(n7954), .A3(n7953), .A4(n7952), .ZN(n7959)
         );
  INV_X1 U9579 ( .A(n7956), .ZN(n7958) );
  NOR3_X1 U9580 ( .A1(n7959), .A2(n7958), .A3(n7957), .ZN(n7963) );
  NAND4_X1 U9581 ( .A1(n7963), .A2(n7962), .A3(n7961), .A4(n7960), .ZN(n7966)
         );
  OR4_X1 U9582 ( .A1(n7967), .A2(n7966), .A3(n7965), .A4(n7964), .ZN(n7968) );
  NOR4_X1 U9583 ( .A1(n7971), .A2(n7970), .A3(n7969), .A4(n7968), .ZN(n7972)
         );
  NAND4_X1 U9584 ( .A1(n9549), .A2(n7974), .A3(n7973), .A4(n7972), .ZN(n7975)
         );
  NOR4_X1 U9585 ( .A1(n9501), .A2(n4502), .A3(n9516), .A4(n7975), .ZN(n7977)
         );
  INV_X1 U9586 ( .A(n9483), .ZN(n7976) );
  NAND4_X1 U9587 ( .A1(n9459), .A2(n9469), .A3(n7977), .A4(n7976), .ZN(n7978)
         );
  NOR4_X1 U9588 ( .A1(n4918), .A2(n9418), .A3(n9436), .A4(n7978), .ZN(n7979)
         );
  NAND4_X1 U9589 ( .A1(n9370), .A2(n7980), .A3(n7979), .A4(n9409), .ZN(n7984)
         );
  INV_X1 U9590 ( .A(n7985), .ZN(n7997) );
  INV_X1 U9591 ( .A(n7986), .ZN(n7993) );
  NAND2_X1 U9592 ( .A1(n9495), .A2(n7987), .ZN(n7989) );
  OAI21_X1 U9593 ( .B1(n7990), .B2(n7989), .A(n7988), .ZN(n7992) );
  OAI21_X1 U9594 ( .B1(n7993), .B2(n7992), .A(n7991), .ZN(n7994) );
  OAI211_X1 U9595 ( .C1(n9653), .C2(n9353), .A(n7995), .B(n7994), .ZN(n7996)
         );
  OAI21_X1 U9596 ( .B1(n9360), .B2(n7997), .A(n7996), .ZN(n7999) );
  AOI211_X1 U9597 ( .C1(n7999), .C2(n4534), .A(n8006), .B(n7998), .ZN(n8000)
         );
  NOR2_X1 U9598 ( .A1(n8011), .A2(n9342), .ZN(n8003) );
  NAND2_X1 U9599 ( .A1(n8003), .A2(n7108), .ZN(n8004) );
  NOR2_X1 U9600 ( .A1(n4534), .A2(n9342), .ZN(n8008) );
  NOR4_X1 U9601 ( .A1(n8009), .A2(n8015), .A3(n8008), .A4(n8007), .ZN(n8010)
         );
  NAND4_X1 U9602 ( .A1(n9173), .A2(n8013), .A3(n8012), .A4(n10031), .ZN(n8014)
         );
  OAI211_X1 U9603 ( .C1(n8015), .C2(n8017), .A(n8014), .B(P1_B_REG_SCAN_IN), 
        .ZN(n8016) );
  INV_X1 U9604 ( .A(n8018), .ZN(n8023) );
  AOI22_X1 U9605 ( .A1(n9076), .A2(n10091), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n10102), .ZN(n8019) );
  OAI21_X1 U9606 ( .B1(n9362), .B2(n10096), .A(n8019), .ZN(n8022) );
  NOR2_X1 U9607 ( .A1(n8020), .A2(n10102), .ZN(n8021) );
  AOI211_X1 U9608 ( .C1(n10081), .C2(n8023), .A(n8022), .B(n8021), .ZN(n8024)
         );
  OAI21_X1 U9609 ( .B1(n8025), .B2(n9557), .A(n8024), .ZN(P1_U3265) );
  NOR4_X1 U9610 ( .A1(n8028), .A2(n6488), .A3(n8027), .A4(n8026), .ZN(n8257)
         );
  OAI21_X1 U9611 ( .B1(n8243), .B2(n8029), .A(P2_B_REG_SCAN_IN), .ZN(n8256) );
  INV_X1 U9612 ( .A(n8030), .ZN(n8031) );
  AOI21_X1 U9613 ( .B1(n8033), .B2(n8032), .A(n8031), .ZN(n8089) );
  AOI211_X1 U9614 ( .C1(n8241), .C2(n8035), .A(n8171), .B(n8034), .ZN(n8038)
         );
  AOI22_X1 U9615 ( .A1(n8212), .A2(n8036), .B1(n8186), .B2(n8042), .ZN(n8037)
         );
  OAI21_X1 U9616 ( .B1(n8038), .B2(n8037), .A(n8757), .ZN(n8047) );
  INV_X1 U9617 ( .A(n8039), .ZN(n8069) );
  OAI21_X1 U9618 ( .B1(n8041), .B2(n8069), .A(n8186), .ZN(n8046) );
  NOR3_X1 U9619 ( .A1(n8041), .A2(n8069), .A3(n8040), .ZN(n8044) );
  INV_X1 U9620 ( .A(n8042), .ZN(n8043) );
  MUX2_X1 U9621 ( .A(n8044), .B(n8043), .S(n8171), .Z(n8045) );
  AOI21_X1 U9622 ( .B1(n8047), .B2(n8046), .A(n8045), .ZN(n8050) );
  AOI21_X1 U9623 ( .B1(n8051), .B2(n8048), .A(n8186), .ZN(n8049) );
  OAI21_X1 U9624 ( .B1(n8050), .B2(n8049), .A(n8213), .ZN(n8070) );
  INV_X1 U9625 ( .A(n8051), .ZN(n8053) );
  OAI211_X1 U9626 ( .C1(n8070), .C2(n8053), .A(n8071), .B(n8052), .ZN(n8054)
         );
  NAND3_X1 U9627 ( .A1(n8054), .A2(n8074), .A3(n8068), .ZN(n8057) );
  NAND2_X1 U9628 ( .A1(n8064), .A2(n8059), .ZN(n8055) );
  NAND2_X1 U9629 ( .A1(n8079), .A2(n8078), .ZN(n8058) );
  MUX2_X1 U9630 ( .A(n8055), .B(n8058), .S(n8186), .Z(n8082) );
  NOR2_X1 U9631 ( .A1(n8082), .A2(n8056), .ZN(n8075) );
  NAND3_X1 U9632 ( .A1(n8057), .A2(n8075), .A3(n8072), .ZN(n8065) );
  INV_X1 U9633 ( .A(n8058), .ZN(n8062) );
  NAND2_X1 U9634 ( .A1(n8060), .A2(n8059), .ZN(n8061) );
  NAND2_X1 U9635 ( .A1(n8062), .A2(n8061), .ZN(n8063) );
  NAND4_X1 U9636 ( .A1(n8065), .A2(n8083), .A3(n8064), .A4(n8063), .ZN(n8066)
         );
  OAI211_X1 U9637 ( .C1(n8070), .C2(n8069), .A(n8068), .B(n8067), .ZN(n8073)
         );
  NAND3_X1 U9638 ( .A1(n8073), .A2(n8072), .A3(n8071), .ZN(n8076) );
  AND3_X1 U9639 ( .A1(n8076), .A2(n8075), .A3(n8074), .ZN(n8085) );
  AND2_X1 U9640 ( .A1(n8078), .A2(n8077), .ZN(n8081) );
  OAI211_X1 U9641 ( .C1(n8082), .C2(n8081), .A(n8080), .B(n8079), .ZN(n8084)
         );
  NOR2_X1 U9642 ( .A1(n8087), .A2(n8086), .ZN(n8210) );
  INV_X1 U9643 ( .A(n8090), .ZN(n8091) );
  MUX2_X1 U9644 ( .A(n8092), .B(n8091), .S(n8171), .Z(n8094) );
  NOR3_X1 U9645 ( .A1(n8095), .A2(n8094), .A3(n8093), .ZN(n8103) );
  XNOR2_X1 U9646 ( .A(n8907), .B(n8730), .ZN(n8209) );
  MUX2_X1 U9647 ( .A(n8097), .B(n8096), .S(n8186), .Z(n8098) );
  NAND2_X1 U9648 ( .A1(n8209), .A2(n8098), .ZN(n8102) );
  INV_X1 U9649 ( .A(n8726), .ZN(n8728) );
  MUX2_X1 U9650 ( .A(n8100), .B(n8099), .S(n8171), .Z(n8101) );
  OAI211_X1 U9651 ( .C1(n8103), .C2(n8102), .A(n8728), .B(n8101), .ZN(n8107)
         );
  INV_X1 U9652 ( .A(n8721), .ZN(n8713) );
  MUX2_X1 U9653 ( .A(n8105), .B(n8104), .S(n8171), .Z(n8106) );
  NAND3_X1 U9654 ( .A1(n8107), .A2(n8713), .A3(n8106), .ZN(n8116) );
  NAND3_X1 U9655 ( .A1(n8116), .A2(n8683), .A3(n8108), .ZN(n8110) );
  NAND3_X1 U9656 ( .A1(n8110), .A2(n8117), .A3(n8109), .ZN(n8111) );
  NAND3_X1 U9657 ( .A1(n8111), .A2(n8119), .A3(n8670), .ZN(n8112) );
  NAND3_X1 U9658 ( .A1(n8112), .A2(n8123), .A3(n8118), .ZN(n8113) );
  NAND2_X1 U9659 ( .A1(n8113), .A2(n8120), .ZN(n8126) );
  INV_X1 U9660 ( .A(n8670), .ZN(n8115) );
  INV_X1 U9661 ( .A(n8683), .ZN(n8114) );
  AOI211_X1 U9662 ( .C1(n8116), .C2(n8682), .A(n8115), .B(n8114), .ZN(n8122)
         );
  NAND2_X1 U9663 ( .A1(n8118), .A2(n8117), .ZN(n8121) );
  OAI211_X1 U9664 ( .C1(n8122), .C2(n8121), .A(n8120), .B(n8119), .ZN(n8124)
         );
  NAND2_X1 U9665 ( .A1(n8124), .A2(n8123), .ZN(n8125) );
  INV_X1 U9666 ( .A(n8127), .ZN(n8648) );
  MUX2_X1 U9667 ( .A(n8129), .B(n8128), .S(n8171), .Z(n8131) );
  INV_X1 U9668 ( .A(n8623), .ZN(n8130) );
  INV_X1 U9669 ( .A(n8208), .ZN(n8132) );
  AOI21_X1 U9670 ( .B1(n8134), .B2(n8133), .A(n8132), .ZN(n8139) );
  OAI21_X1 U9671 ( .B1(n8136), .B2(n8135), .A(n8207), .ZN(n8137) );
  NAND2_X1 U9672 ( .A1(n8137), .A2(n8208), .ZN(n8138) );
  MUX2_X1 U9673 ( .A(n8139), .B(n8138), .S(n8186), .Z(n8146) );
  INV_X1 U9674 ( .A(n8144), .ZN(n8140) );
  INV_X1 U9675 ( .A(n8149), .ZN(n8141) );
  INV_X1 U9676 ( .A(n8142), .ZN(n8143) );
  MUX2_X1 U9677 ( .A(n8144), .B(n8143), .S(n8171), .Z(n8145) );
  OAI211_X1 U9678 ( .C1(n8146), .C2(n8618), .A(n8604), .B(n8145), .ZN(n8155)
         );
  INV_X1 U9679 ( .A(n8584), .ZN(n8591) );
  INV_X1 U9680 ( .A(n8147), .ZN(n8148) );
  MUX2_X1 U9681 ( .A(n8149), .B(n8148), .S(n8186), .Z(n8150) );
  NOR2_X1 U9682 ( .A1(n8591), .A2(n8150), .ZN(n8154) );
  NOR2_X1 U9683 ( .A1(n8843), .A2(n8400), .ZN(n8151) );
  MUX2_X1 U9684 ( .A(n8152), .B(n8151), .S(n8186), .Z(n8153) );
  AOI21_X1 U9685 ( .B1(n8155), .B2(n8154), .A(n8153), .ZN(n8167) );
  INV_X1 U9686 ( .A(n8167), .ZN(n8160) );
  MUX2_X1 U9687 ( .A(n8156), .B(n8782), .S(n8186), .Z(n8165) );
  INV_X1 U9688 ( .A(n8165), .ZN(n8159) );
  INV_X1 U9689 ( .A(n8286), .ZN(n8399) );
  MUX2_X1 U9690 ( .A(n8171), .B(n8399), .S(n8184), .Z(n8157) );
  AOI21_X1 U9691 ( .B1(n8286), .B2(n8186), .A(n8157), .ZN(n8166) );
  INV_X1 U9692 ( .A(n8166), .ZN(n8158) );
  OAI21_X1 U9693 ( .B1(n8160), .B2(n8159), .A(n8158), .ZN(n8183) );
  NAND2_X1 U9694 ( .A1(n8161), .A2(n5176), .ZN(n8163) );
  NAND2_X1 U9695 ( .A1(n5461), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8162) );
  NAND2_X1 U9696 ( .A1(n8835), .A2(n8169), .ZN(n8170) );
  NAND2_X1 U9697 ( .A1(n8184), .A2(n8286), .ZN(n8164) );
  AND2_X1 U9698 ( .A1(n8170), .A2(n8164), .ZN(n8194) );
  NOR3_X1 U9699 ( .A1(n8167), .A2(n8166), .A3(n8165), .ZN(n8187) );
  INV_X1 U9700 ( .A(n8187), .ZN(n8168) );
  OAI211_X1 U9701 ( .C1(n8183), .C2(n8588), .A(n8194), .B(n8168), .ZN(n8190)
         );
  OR2_X1 U9702 ( .A1(n8835), .A2(n8169), .ZN(n8198) );
  INV_X1 U9703 ( .A(n8198), .ZN(n8172) );
  OAI21_X1 U9704 ( .B1(n8172), .B2(n8171), .A(n8170), .ZN(n8189) );
  NAND2_X1 U9705 ( .A1(n8912), .A2(n5176), .ZN(n8175) );
  NAND2_X1 U9706 ( .A1(n5461), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8174) );
  INV_X1 U9707 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8178) );
  NAND2_X1 U9708 ( .A1(n5189), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8177) );
  INV_X1 U9709 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n9886) );
  OR2_X1 U9710 ( .A1(n4393), .A2(n9886), .ZN(n8176) );
  OAI211_X1 U9711 ( .C1(n8179), .C2(n8178), .A(n8177), .B(n8176), .ZN(n8180)
         );
  INV_X1 U9712 ( .A(n8180), .ZN(n8181) );
  OR2_X1 U9713 ( .A1(n8831), .A2(n8570), .ZN(n8195) );
  INV_X1 U9714 ( .A(n8195), .ZN(n8188) );
  NOR2_X1 U9715 ( .A1(n8184), .A2(n8286), .ZN(n8192) );
  INV_X1 U9716 ( .A(n8192), .ZN(n8185) );
  NAND2_X1 U9717 ( .A1(n8198), .A2(n8185), .ZN(n8237) );
  AND2_X1 U9718 ( .A1(n8831), .A2(n8570), .ZN(n8238) );
  XNOR2_X1 U9719 ( .A(n8191), .B(n8555), .ZN(n8253) );
  NOR2_X1 U9720 ( .A1(n8193), .A2(n8192), .ZN(n8202) );
  NAND2_X1 U9721 ( .A1(n8195), .A2(n8194), .ZN(n8239) );
  INV_X1 U9722 ( .A(n8239), .ZN(n8197) );
  INV_X1 U9723 ( .A(n8831), .ZN(n8573) );
  INV_X1 U9724 ( .A(n8570), .ZN(n8398) );
  NAND2_X1 U9725 ( .A1(n8198), .A2(n8398), .ZN(n8199) );
  NOR2_X1 U9726 ( .A1(n8203), .A2(n8555), .ZN(n8240) );
  NAND3_X1 U9727 ( .A1(n8205), .A2(n8204), .A3(n8240), .ZN(n8252) );
  AND2_X1 U9728 ( .A1(n8555), .A2(n8254), .ZN(n8242) );
  INV_X1 U9729 ( .A(n8242), .ZN(n8206) );
  NOR2_X1 U9730 ( .A1(n8206), .A2(n8241), .ZN(n8249) );
  NAND2_X1 U9731 ( .A1(n8208), .A2(n8207), .ZN(n8627) );
  INV_X1 U9732 ( .A(n8657), .ZN(n8661) );
  INV_X1 U9733 ( .A(n8674), .ZN(n8671) );
  INV_X1 U9734 ( .A(n8210), .ZN(n8224) );
  NAND4_X1 U9735 ( .A1(n8213), .A2(n8212), .A3(n8211), .A4(n8757), .ZN(n8218)
         );
  NAND2_X1 U9736 ( .A1(n8215), .A2(n8214), .ZN(n8217) );
  NOR3_X1 U9737 ( .A1(n8218), .A2(n8217), .A3(n8216), .ZN(n8221) );
  NAND4_X1 U9738 ( .A1(n8221), .A2(n4607), .A3(n8220), .A4(n8219), .ZN(n8222)
         );
  NOR3_X1 U9739 ( .A1(n8224), .A2(n8223), .A3(n8222), .ZN(n8226) );
  NAND3_X1 U9740 ( .A1(n8227), .A2(n8226), .A3(n8225), .ZN(n8228) );
  NOR3_X1 U9741 ( .A1(n8726), .A2(n8739), .A3(n8228), .ZN(n8229) );
  NAND3_X1 U9742 ( .A1(n8703), .A2(n8713), .A3(n8229), .ZN(n8230) );
  NOR2_X1 U9743 ( .A1(n8231), .A2(n8230), .ZN(n8232) );
  NAND4_X1 U9744 ( .A1(n8648), .A2(n8661), .A3(n8671), .A4(n8232), .ZN(n8233)
         );
  OR4_X1 U9745 ( .A1(n8618), .A2(n8627), .A3(n8233), .A4(n8638), .ZN(n8234) );
  NOR2_X1 U9746 ( .A1(n8599), .A2(n8234), .ZN(n8235) );
  NAND3_X1 U9747 ( .A1(n8279), .A2(n8235), .A3(n8584), .ZN(n8236) );
  NAND2_X1 U9748 ( .A1(n8240), .A2(n8241), .ZN(n8246) );
  NAND3_X1 U9749 ( .A1(n8247), .A2(n8242), .A3(n8241), .ZN(n8245) );
  INV_X1 U9750 ( .A(n8243), .ZN(n8244) );
  OAI211_X1 U9751 ( .C1(n8247), .C2(n8246), .A(n8245), .B(n8244), .ZN(n8248)
         );
  AOI21_X1 U9752 ( .B1(n8250), .B2(n8249), .A(n8248), .ZN(n8251) );
  OAI211_X1 U9753 ( .C1(n8254), .C2(n8253), .A(n8252), .B(n8251), .ZN(n8255)
         );
  OAI21_X1 U9754 ( .B1(n8257), .B2(n8256), .A(n8255), .ZN(P2_U3296) );
  OAI222_X1 U9755 ( .A1(n8260), .A2(P2_U3151), .B1(n8918), .B2(n8259), .C1(
        n9755), .C2(n8258), .ZN(P2_U3265) );
  AOI21_X1 U9756 ( .B1(n8651), .B2(n8261), .A(n8346), .ZN(n8267) );
  AOI22_X1 U9757 ( .A1(n8640), .A2(n8372), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8263) );
  NAND2_X1 U9758 ( .A1(n8394), .A2(n8642), .ZN(n8262) );
  OAI211_X1 U9759 ( .C1(n8264), .C2(n8376), .A(n8263), .B(n8262), .ZN(n8265)
         );
  AOI21_X1 U9760 ( .B1(n8865), .B2(n8379), .A(n8265), .ZN(n8266) );
  OAI21_X1 U9761 ( .B1(n8267), .B2(n8381), .A(n8266), .ZN(P2_U3156) );
  XNOR2_X1 U9762 ( .A(n8268), .B(n8357), .ZN(n8269) );
  XNOR2_X1 U9763 ( .A(n8270), .B(n8269), .ZN(n8275) );
  NAND2_X1 U9764 ( .A1(n8390), .A2(n8714), .ZN(n8271) );
  NAND2_X1 U9765 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8556) );
  OAI211_X1 U9766 ( .C1(n8693), .C2(n8392), .A(n8271), .B(n8556), .ZN(n8272)
         );
  AOI21_X1 U9767 ( .B1(n8698), .B2(n8394), .A(n8272), .ZN(n8274) );
  NAND2_X1 U9768 ( .A1(n8889), .A2(n8379), .ZN(n8273) );
  OAI211_X1 U9769 ( .C1(n8275), .C2(n8381), .A(n8274), .B(n8273), .ZN(P2_U3159) );
  INV_X1 U9770 ( .A(n8276), .ZN(n8278) );
  XOR2_X1 U9771 ( .A(n8280), .B(n8279), .Z(n8281) );
  XNOR2_X1 U9772 ( .A(n8282), .B(n8281), .ZN(n8290) );
  AOI22_X1 U9773 ( .A1(n8400), .A2(n8390), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8285) );
  NAND2_X1 U9774 ( .A1(n8283), .A2(n8394), .ZN(n8284) );
  OAI211_X1 U9775 ( .C1(n8286), .C2(n8392), .A(n8285), .B(n8284), .ZN(n8287)
         );
  AOI21_X1 U9776 ( .B1(n8288), .B2(n8379), .A(n8287), .ZN(n8289) );
  OAI21_X1 U9777 ( .B1(n8290), .B2(n8381), .A(n8289), .ZN(P2_U3160) );
  INV_X1 U9778 ( .A(n8877), .ZN(n8300) );
  NOR3_X1 U9779 ( .A1(n4420), .A2(n4782), .A3(n8292), .ZN(n8295) );
  INV_X1 U9780 ( .A(n8293), .ZN(n8294) );
  OAI21_X1 U9781 ( .B1(n8295), .B2(n8294), .A(n8387), .ZN(n8299) );
  AOI22_X1 U9782 ( .A1(n8372), .A2(n8664), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8296) );
  OAI21_X1 U9783 ( .B1(n8693), .B2(n8376), .A(n8296), .ZN(n8297) );
  AOI21_X1 U9784 ( .B1(n8667), .B2(n8394), .A(n8297), .ZN(n8298) );
  OAI211_X1 U9785 ( .C1(n8300), .C2(n8397), .A(n8299), .B(n8298), .ZN(P2_U3163) );
  OAI21_X1 U9786 ( .B1(n8303), .B2(n8302), .A(n8301), .ZN(n8305) );
  XNOR2_X1 U9787 ( .A(n8305), .B(n8304), .ZN(n8314) );
  NAND2_X1 U9788 ( .A1(n10282), .A2(n8379), .ZN(n8311) );
  NAND2_X1 U9789 ( .A1(n8390), .A2(n8404), .ZN(n8307) );
  OAI211_X1 U9790 ( .C1(n8308), .C2(n8392), .A(n8307), .B(n8306), .ZN(n8309)
         );
  INV_X1 U9791 ( .A(n8309), .ZN(n8310) );
  OAI211_X1 U9792 ( .C1(n8312), .C2(n8339), .A(n8311), .B(n8310), .ZN(n8313)
         );
  AOI21_X1 U9793 ( .B1(n8314), .B2(n8387), .A(n8313), .ZN(n8315) );
  INV_X1 U9794 ( .A(n8315), .ZN(P2_U3164) );
  INV_X1 U9795 ( .A(n8853), .ZN(n8793) );
  AND3_X1 U9796 ( .A1(n8316), .A2(n8318), .A3(n8317), .ZN(n8319) );
  OAI21_X1 U9797 ( .B1(n8386), .B2(n8319), .A(n8387), .ZN(n8323) );
  AOI22_X1 U9798 ( .A1(n8587), .A2(n8372), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8320) );
  OAI21_X1 U9799 ( .B1(n8614), .B2(n8376), .A(n8320), .ZN(n8321) );
  AOI21_X1 U9800 ( .B1(n8616), .B2(n8394), .A(n8321), .ZN(n8322) );
  OAI211_X1 U9801 ( .C1(n8793), .C2(n8397), .A(n8323), .B(n8322), .ZN(P2_U3165) );
  INV_X1 U9802 ( .A(n8324), .ZN(n8335) );
  AOI21_X1 U9803 ( .B1(n8326), .B2(n8325), .A(n8335), .ZN(n8331) );
  NAND2_X1 U9804 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8496) );
  OAI21_X1 U9805 ( .B1(n8392), .B2(n8377), .A(n8496), .ZN(n8327) );
  AOI21_X1 U9806 ( .B1(n8390), .B2(n8730), .A(n8327), .ZN(n8328) );
  OAI21_X1 U9807 ( .B1(n8734), .B2(n8339), .A(n8328), .ZN(n8329) );
  AOI21_X1 U9808 ( .B1(n8901), .B2(n8379), .A(n8329), .ZN(n8330) );
  OAI21_X1 U9809 ( .B1(n8331), .B2(n8381), .A(n8330), .ZN(P2_U3166) );
  INV_X1 U9810 ( .A(n8818), .ZN(n8344) );
  INV_X1 U9811 ( .A(n8332), .ZN(n8334) );
  NOR3_X1 U9812 ( .A1(n8335), .A2(n8334), .A3(n8333), .ZN(n8338) );
  INV_X1 U9813 ( .A(n8336), .ZN(n8337) );
  OAI21_X1 U9814 ( .B1(n8338), .B2(n8337), .A(n8387), .ZN(n8343) );
  OAI22_X1 U9815 ( .A1(n8392), .A2(n8692), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10234), .ZN(n8341) );
  NOR2_X1 U9816 ( .A1(n8339), .A2(n8716), .ZN(n8340) );
  AOI211_X1 U9817 ( .C1(n8390), .C2(n8743), .A(n8341), .B(n8340), .ZN(n8342)
         );
  OAI211_X1 U9818 ( .C1(n8344), .C2(n8397), .A(n8343), .B(n8342), .ZN(P2_U3168) );
  INV_X1 U9819 ( .A(n8859), .ZN(n8798) );
  INV_X1 U9820 ( .A(n8316), .ZN(n8348) );
  NOR3_X1 U9821 ( .A1(n8346), .A2(n4414), .A3(n8345), .ZN(n8347) );
  OAI21_X1 U9822 ( .B1(n8348), .B2(n8347), .A(n8387), .ZN(n8352) );
  AOI22_X1 U9823 ( .A1(n8401), .A2(n8372), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8349) );
  OAI21_X1 U9824 ( .B1(n8630), .B2(n8376), .A(n8349), .ZN(n8350) );
  AOI21_X1 U9825 ( .B1(n8634), .B2(n8394), .A(n8350), .ZN(n8351) );
  OAI211_X1 U9826 ( .C1(n8798), .C2(n8397), .A(n8352), .B(n8351), .ZN(P2_U3169) );
  AOI21_X1 U9827 ( .B1(n8354), .B2(n8353), .A(n4420), .ZN(n8360) );
  AOI22_X1 U9828 ( .A1(n8372), .A2(n8676), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8356) );
  NAND2_X1 U9829 ( .A1(n8394), .A2(n8679), .ZN(n8355) );
  OAI211_X1 U9830 ( .C1(n8357), .C2(n8376), .A(n8356), .B(n8355), .ZN(n8358)
         );
  AOI21_X1 U9831 ( .B1(n8883), .B2(n8379), .A(n8358), .ZN(n8359) );
  OAI21_X1 U9832 ( .B1(n8360), .B2(n8381), .A(n8359), .ZN(P2_U3173) );
  INV_X1 U9833 ( .A(n8871), .ZN(n8369) );
  AOI21_X1 U9834 ( .B1(n8362), .B2(n8361), .A(n8381), .ZN(n8364) );
  NAND2_X1 U9835 ( .A1(n8364), .A2(n8363), .ZN(n8368) );
  AOI22_X1 U9836 ( .A1(n8390), .A2(n8676), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8365) );
  OAI21_X1 U9837 ( .B1(n8630), .B2(n8392), .A(n8365), .ZN(n8366) );
  AOI21_X1 U9838 ( .B1(n8654), .B2(n8394), .A(n8366), .ZN(n8367) );
  OAI211_X1 U9839 ( .C1(n8369), .C2(n8397), .A(n8368), .B(n8367), .ZN(P2_U3175) );
  XOR2_X1 U9840 ( .A(n8371), .B(n8370), .Z(n8382) );
  AOI22_X1 U9841 ( .A1(n8372), .A2(n8706), .B1(P2_REG3_REG_18__SCAN_IN), .B2(
        P2_U3151), .ZN(n8375) );
  INV_X1 U9842 ( .A(n8373), .ZN(n8709) );
  NAND2_X1 U9843 ( .A1(n8394), .A2(n8709), .ZN(n8374) );
  OAI211_X1 U9844 ( .C1(n8377), .C2(n8376), .A(n8375), .B(n8374), .ZN(n8378)
         );
  AOI21_X1 U9845 ( .B1(n8894), .B2(n8379), .A(n8378), .ZN(n8380) );
  OAI21_X1 U9846 ( .B1(n8382), .B2(n8381), .A(n8380), .ZN(P2_U3178) );
  INV_X1 U9847 ( .A(n8846), .ZN(n8790) );
  INV_X1 U9848 ( .A(n8383), .ZN(n8389) );
  NOR3_X1 U9849 ( .A1(n8386), .A2(n8385), .A3(n8384), .ZN(n8388) );
  OAI21_X1 U9850 ( .B1(n8389), .B2(n8388), .A(n8387), .ZN(n8396) );
  AOI22_X1 U9851 ( .A1(n8401), .A2(n8390), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8391) );
  OAI21_X1 U9852 ( .B1(n8607), .B2(n8392), .A(n8391), .ZN(n8393) );
  AOI21_X1 U9853 ( .B1(n8609), .B2(n8394), .A(n8393), .ZN(n8395) );
  OAI211_X1 U9854 ( .C1(n8790), .C2(n8397), .A(n8396), .B(n8395), .ZN(P2_U3180) );
  MUX2_X1 U9855 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8398), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U9856 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8399), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U9857 ( .A(n8588), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8527), .Z(
        P2_U3519) );
  MUX2_X1 U9858 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8400), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9859 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8587), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U9860 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8401), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9861 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8640), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9862 ( .A(n8651), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8527), .Z(
        P2_U3514) );
  MUX2_X1 U9863 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8664), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9864 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8676), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9865 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8663), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9866 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8706), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9867 ( .A(n8714), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8527), .Z(
        P2_U3509) );
  MUX2_X1 U9868 ( .A(n8731), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8527), .Z(
        P2_U3508) );
  MUX2_X1 U9869 ( .A(n8743), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8527), .Z(
        P2_U3507) );
  MUX2_X1 U9870 ( .A(n8730), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8527), .Z(
        P2_U3506) );
  MUX2_X1 U9871 ( .A(n8742), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8527), .Z(
        P2_U3505) );
  MUX2_X1 U9872 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8402), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U9873 ( .A(n8403), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8527), .Z(
        P2_U3503) );
  MUX2_X1 U9874 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8404), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U9875 ( .A(n8405), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8527), .Z(
        P2_U3501) );
  MUX2_X1 U9876 ( .A(n8406), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8527), .Z(
        P2_U3500) );
  MUX2_X1 U9877 ( .A(n8407), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8527), .Z(
        P2_U3499) );
  MUX2_X1 U9878 ( .A(n8408), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8527), .Z(
        P2_U3498) );
  MUX2_X1 U9879 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8409), .S(P2_U3893), .Z(
        P2_U3497) );
  MUX2_X1 U9880 ( .A(n8410), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8527), .Z(
        P2_U3496) );
  MUX2_X1 U9881 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8411), .S(P2_U3893), .Z(
        P2_U3495) );
  MUX2_X1 U9882 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8412), .S(P2_U3893), .Z(
        P2_U3494) );
  MUX2_X1 U9883 ( .A(n8413), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8527), .Z(
        P2_U3493) );
  MUX2_X1 U9884 ( .A(n8414), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8527), .Z(
        P2_U3492) );
  MUX2_X1 U9885 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n8415), .S(P2_U3893), .Z(
        P2_U3491) );
  NAND2_X1 U9886 ( .A1(n8428), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n8416) );
  AOI21_X1 U9887 ( .B1(n8418), .B2(n8420), .A(n8453), .ZN(n8437) );
  NAND2_X1 U9888 ( .A1(n8551), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8419) );
  OAI21_X1 U9889 ( .B1(n8551), .B2(n8420), .A(n8419), .ZN(n8445) );
  XNOR2_X1 U9890 ( .A(n8445), .B(n8452), .ZN(n8425) );
  OR2_X1 U9891 ( .A1(n8428), .A2(n8421), .ZN(n8423) );
  NAND2_X1 U9892 ( .A1(n8423), .A2(n8422), .ZN(n8424) );
  NAND2_X1 U9893 ( .A1(n8425), .A2(n8424), .ZN(n8446) );
  OAI21_X1 U9894 ( .B1(n8425), .B2(n8424), .A(n8446), .ZN(n8435) );
  INV_X1 U9895 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n10008) );
  NAND2_X1 U9896 ( .A1(n10213), .A2(n8452), .ZN(n8427) );
  OAI211_X1 U9897 ( .C1(n10008), .C2(n10192), .A(n8427), .B(n8426), .ZN(n8434)
         );
  NAND2_X1 U9898 ( .A1(n8428), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n8429) );
  AOI21_X1 U9899 ( .B1(n9752), .B2(n8431), .A(n8439), .ZN(n8432) );
  NOR2_X1 U9900 ( .A1(n8432), .A2(n10229), .ZN(n8433) );
  AOI211_X1 U9901 ( .C1(n10225), .C2(n8435), .A(n8434), .B(n8433), .ZN(n8436)
         );
  OAI21_X1 U9902 ( .B1(n8437), .B2(n10220), .A(n8436), .ZN(P2_U3195) );
  AOI22_X1 U9903 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8455), .B1(n8475), .B2(
        n8440), .ZN(n8441) );
  NOR2_X1 U9904 ( .A1(n8442), .A2(n8441), .ZN(n8474) );
  AOI21_X1 U9905 ( .B1(n8442), .B2(n8441), .A(n8474), .ZN(n8463) );
  OR2_X1 U9906 ( .A1(n8551), .A2(n9911), .ZN(n8444) );
  NAND2_X1 U9907 ( .A1(n8551), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8443) );
  NAND2_X1 U9908 ( .A1(n8444), .A2(n8443), .ZN(n8467) );
  XNOR2_X1 U9909 ( .A(n8467), .B(n8455), .ZN(n8449) );
  OR2_X1 U9910 ( .A1(n4639), .A2(n8445), .ZN(n8447) );
  NAND2_X1 U9911 ( .A1(n8447), .A2(n8446), .ZN(n8448) );
  NAND2_X1 U9912 ( .A1(n8449), .A2(n8448), .ZN(n8468) );
  OAI21_X1 U9913 ( .B1(n8449), .B2(n8448), .A(n8468), .ZN(n8461) );
  NAND2_X1 U9914 ( .A1(n10212), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n8451) );
  OAI211_X1 U9915 ( .C1(n10204), .C2(n8475), .A(n8451), .B(n8450), .ZN(n8460)
         );
  NOR2_X1 U9916 ( .A1(n8452), .A2(n4438), .ZN(n8454) );
  AOI22_X1 U9917 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8455), .B1(n8475), .B2(
        n9911), .ZN(n8456) );
  NOR2_X1 U9918 ( .A1(n8457), .A2(n8456), .ZN(n8464) );
  AOI21_X1 U9919 ( .B1(n8457), .B2(n8456), .A(n8464), .ZN(n8458) );
  NOR2_X1 U9920 ( .A1(n8458), .A2(n10220), .ZN(n8459) );
  AOI211_X1 U9921 ( .C1(n10225), .C2(n8461), .A(n8460), .B(n8459), .ZN(n8462)
         );
  OAI21_X1 U9922 ( .B1(n8463), .B2(n10229), .A(n8462), .ZN(P2_U3196) );
  AOI21_X1 U9923 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8475), .A(n8464), .ZN(
        n8483) );
  XNOR2_X1 U9924 ( .A(n8483), .B(n8499), .ZN(n8465) );
  NOR2_X1 U9925 ( .A1(n8746), .A2(n8465), .ZN(n8484) );
  AOI21_X1 U9926 ( .B1(n8465), .B2(n8746), .A(n8484), .ZN(n8482) );
  NAND2_X1 U9927 ( .A1(n8551), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8466) );
  OAI21_X1 U9928 ( .B1(n8551), .B2(n8746), .A(n8466), .ZN(n8490) );
  XNOR2_X1 U9929 ( .A(n8490), .B(n8499), .ZN(n8471) );
  OR2_X1 U9930 ( .A1(n8475), .A2(n8467), .ZN(n8469) );
  NAND2_X1 U9931 ( .A1(n8469), .A2(n8468), .ZN(n8470) );
  NAND2_X1 U9932 ( .A1(n8471), .A2(n8470), .ZN(n8492) );
  OAI21_X1 U9933 ( .B1(n8471), .B2(n8470), .A(n8492), .ZN(n8480) );
  INV_X1 U9934 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n10014) );
  NAND2_X1 U9935 ( .A1(n10213), .A2(n8499), .ZN(n8473) );
  OAI211_X1 U9936 ( .C1(n10014), .C2(n10192), .A(n8473), .B(n8472), .ZN(n8479)
         );
  XNOR2_X1 U9937 ( .A(n8498), .B(n8499), .ZN(n8476) );
  NOR2_X1 U9938 ( .A1(n8825), .A2(n8476), .ZN(n8500) );
  AOI21_X1 U9939 ( .B1(n8825), .B2(n8476), .A(n8500), .ZN(n8477) );
  NOR2_X1 U9940 ( .A1(n8477), .A2(n10229), .ZN(n8478) );
  AOI211_X1 U9941 ( .C1(n10225), .C2(n8480), .A(n8479), .B(n8478), .ZN(n8481)
         );
  OAI21_X1 U9942 ( .B1(n8482), .B2(n10220), .A(n8481), .ZN(P2_U3197) );
  NOR2_X1 U9943 ( .A1(n8499), .A2(n8483), .ZN(n8485) );
  AOI22_X1 U9944 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8502), .B1(n8533), .B2(
        n8733), .ZN(n8486) );
  AOI21_X1 U9945 ( .B1(n8487), .B2(n8486), .A(n8511), .ZN(n8510) );
  OR2_X1 U9946 ( .A1(n8551), .A2(n8733), .ZN(n8489) );
  NAND2_X1 U9947 ( .A1(n8551), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8488) );
  NAND2_X1 U9948 ( .A1(n8489), .A2(n8488), .ZN(n8519) );
  XNOR2_X1 U9949 ( .A(n8519), .B(n8502), .ZN(n8495) );
  INV_X1 U9950 ( .A(n8490), .ZN(n8491) );
  NAND2_X1 U9951 ( .A1(n8499), .A2(n8491), .ZN(n8493) );
  NAND2_X1 U9952 ( .A1(n8493), .A2(n8492), .ZN(n8494) );
  NAND2_X1 U9953 ( .A1(n8495), .A2(n8494), .ZN(n8520) );
  OAI21_X1 U9954 ( .B1(n8495), .B2(n8494), .A(n8520), .ZN(n8508) );
  NAND2_X1 U9955 ( .A1(n10212), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n8497) );
  OAI211_X1 U9956 ( .C1(n10204), .C2(n8533), .A(n8497), .B(n8496), .ZN(n8507)
         );
  NOR2_X1 U9957 ( .A1(n8499), .A2(n8498), .ZN(n8501) );
  AOI22_X1 U9958 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8502), .B1(n8533), .B2(
        n8822), .ZN(n8503) );
  AOI21_X1 U9959 ( .B1(n8504), .B2(n8503), .A(n8532), .ZN(n8505) );
  NOR2_X1 U9960 ( .A1(n8505), .A2(n10229), .ZN(n8506) );
  AOI211_X1 U9961 ( .C1(n10225), .C2(n8508), .A(n8507), .B(n8506), .ZN(n8509)
         );
  OAI21_X1 U9962 ( .B1(n8510), .B2(n10220), .A(n8509), .ZN(P2_U3198) );
  NOR2_X1 U9963 ( .A1(n10214), .A2(n8512), .ZN(n8513) );
  NOR2_X1 U9964 ( .A1(n8717), .A2(n10219), .ZN(n10218) );
  NOR2_X1 U9965 ( .A1(n8513), .A2(n10218), .ZN(n8515) );
  NAND2_X1 U9966 ( .A1(n8536), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8543) );
  OAI21_X1 U9967 ( .B1(n8536), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8543), .ZN(
        n8514) );
  NOR2_X1 U9968 ( .A1(n8515), .A2(n8514), .ZN(n8545) );
  AOI21_X1 U9969 ( .B1(n8515), .B2(n8514), .A(n8545), .ZN(n8542) );
  NAND2_X1 U9970 ( .A1(n8551), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8516) );
  OAI21_X1 U9971 ( .B1(n8551), .B2(n8717), .A(n8516), .ZN(n8518) );
  OR2_X1 U9972 ( .A1(n8518), .A2(n8517), .ZN(n8522) );
  XNOR2_X1 U9973 ( .A(n8518), .B(n10214), .ZN(n10224) );
  OR2_X1 U9974 ( .A1(n8533), .A2(n8519), .ZN(n8521) );
  NAND2_X1 U9975 ( .A1(n8521), .A2(n8520), .ZN(n10223) );
  NAND2_X1 U9976 ( .A1(n10224), .A2(n10223), .ZN(n10222) );
  AND2_X1 U9977 ( .A1(n8522), .A2(n10222), .ZN(n8525) );
  INV_X1 U9978 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8708) );
  NAND2_X1 U9979 ( .A1(n8551), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8523) );
  OAI21_X1 U9980 ( .B1(n8551), .B2(n8708), .A(n8523), .ZN(n8524) );
  NOR2_X1 U9981 ( .A1(n8525), .A2(n8524), .ZN(n8549) );
  INV_X1 U9982 ( .A(n8549), .ZN(n8526) );
  NAND2_X1 U9983 ( .A1(n8525), .A2(n8524), .ZN(n8547) );
  NAND2_X1 U9984 ( .A1(n8526), .A2(n8547), .ZN(n8528) );
  OAI21_X1 U9985 ( .B1(n8528), .B2(n8527), .A(n10204), .ZN(n8541) );
  INV_X1 U9986 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10314) );
  NAND3_X1 U9987 ( .A1(n8528), .A2(n10225), .A3(n8536), .ZN(n8531) );
  INV_X1 U9988 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8529) );
  OR2_X1 U9989 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8529), .ZN(n8530) );
  OAI211_X1 U9990 ( .C1(n10314), .C2(n10192), .A(n8531), .B(n8530), .ZN(n8540)
         );
  NOR2_X1 U9991 ( .A1(n10214), .A2(n8534), .ZN(n8535) );
  NAND2_X1 U9992 ( .A1(n8536), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8560) );
  OAI21_X1 U9993 ( .B1(n8536), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8560), .ZN(
        n8537) );
  NOR2_X1 U9994 ( .A1(n8538), .A2(n8537), .ZN(n8562) );
  INV_X1 U9995 ( .A(n8543), .ZN(n8544) );
  NOR2_X1 U9996 ( .A1(n8545), .A2(n8544), .ZN(n8546) );
  XNOR2_X1 U9997 ( .A(n8555), .B(n8697), .ZN(n8550) );
  XNOR2_X1 U9998 ( .A(n8546), .B(n8550), .ZN(n8568) );
  OAI21_X1 U9999 ( .B1(n8549), .B2(n8548), .A(n8547), .ZN(n8554) );
  INV_X1 U10000 ( .A(n8550), .ZN(n8552) );
  XNOR2_X1 U10001 ( .A(n8555), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8563) );
  MUX2_X1 U10002 ( .A(n8552), .B(n8563), .S(n8551), .Z(n8553) );
  XNOR2_X1 U10003 ( .A(n8554), .B(n8553), .ZN(n8559) );
  NOR2_X1 U10004 ( .A1(n10204), .A2(n8555), .ZN(n8558) );
  INV_X1 U10005 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n9781) );
  OAI21_X1 U10006 ( .B1(n10192), .B2(n9781), .A(n8556), .ZN(n8557) );
  AOI211_X1 U10007 ( .C1(n8559), .C2(n10225), .A(n8558), .B(n8557), .ZN(n8567)
         );
  INV_X1 U10008 ( .A(n8560), .ZN(n8561) );
  NOR2_X1 U10009 ( .A1(n8562), .A2(n8561), .ZN(n8564) );
  XNOR2_X1 U10010 ( .A(n8564), .B(n8563), .ZN(n8565) );
  NAND2_X1 U10011 ( .A1(n8565), .A2(n10197), .ZN(n8566) );
  OAI211_X1 U10012 ( .C1(n8568), .C2(n10220), .A(n8567), .B(n8566), .ZN(
        P2_U3201) );
  NAND2_X1 U10013 ( .A1(n8571), .A2(n8748), .ZN(n8579) );
  OAI21_X1 U10014 ( .B1(n8725), .B2(n8776), .A(n8579), .ZN(n8574) );
  AOI21_X1 U10015 ( .B1(n8725), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8574), .ZN(
        n8572) );
  OAI21_X1 U10016 ( .B1(n8573), .B2(n8595), .A(n8572), .ZN(P2_U3202) );
  INV_X1 U10017 ( .A(n8835), .ZN(n8780) );
  AOI21_X1 U10018 ( .B1(n8725), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8574), .ZN(
        n8575) );
  OAI21_X1 U10019 ( .B1(n8780), .B2(n8595), .A(n8575), .ZN(P2_U3203) );
  INV_X1 U10020 ( .A(n8576), .ZN(n8583) );
  NAND2_X1 U10021 ( .A1(n8725), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8578) );
  OAI211_X1 U10022 ( .C1(n8580), .C2(n8595), .A(n8579), .B(n8578), .ZN(n8581)
         );
  AOI21_X1 U10023 ( .B1(n8577), .B2(n8745), .A(n8581), .ZN(n8582) );
  OAI21_X1 U10024 ( .B1(n8583), .B2(n8752), .A(n8582), .ZN(P2_U3204) );
  XNOR2_X1 U10025 ( .A(n8585), .B(n8584), .ZN(n8586) );
  NAND2_X1 U10026 ( .A1(n8586), .A2(n8765), .ZN(n8590) );
  AOI22_X1 U10027 ( .A1(n8588), .A2(n5047), .B1(n8741), .B2(n8587), .ZN(n8589)
         );
  NAND2_X1 U10028 ( .A1(n8590), .A2(n8589), .ZN(n8786) );
  INV_X1 U10029 ( .A(n8786), .ZN(n8598) );
  XNOR2_X1 U10030 ( .A(n8592), .B(n8591), .ZN(n8787) );
  AOI22_X1 U10031 ( .A1(n8593), .A2(n8748), .B1(n8725), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n8594) );
  OAI21_X1 U10032 ( .B1(n8843), .B2(n8595), .A(n8594), .ZN(n8596) );
  AOI21_X1 U10033 ( .B1(n8787), .B2(n8619), .A(n8596), .ZN(n8597) );
  OAI21_X1 U10034 ( .B1(n8725), .B2(n8598), .A(n8597), .ZN(P2_U3206) );
  XNOR2_X1 U10035 ( .A(n8600), .B(n8599), .ZN(n8849) );
  INV_X1 U10036 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8608) );
  NAND2_X1 U10037 ( .A1(n8603), .A2(n8602), .ZN(n8605) );
  XNOR2_X1 U10038 ( .A(n8605), .B(n8604), .ZN(n8606) );
  OAI222_X1 U10039 ( .A1(n8762), .A2(n8607), .B1(n8761), .B2(n8631), .C1(n8629), .C2(n8606), .ZN(n8789) );
  INV_X1 U10040 ( .A(n8789), .ZN(n8844) );
  MUX2_X1 U10041 ( .A(n8608), .B(n8844), .S(n8745), .Z(n8611) );
  AOI22_X1 U10042 ( .A1(n8846), .A2(n8749), .B1(n8748), .B2(n8609), .ZN(n8610)
         );
  OAI211_X1 U10043 ( .C1(n8849), .C2(n8752), .A(n8611), .B(n8610), .ZN(
        P2_U3207) );
  NOR2_X1 U10044 ( .A1(n8793), .A2(n8632), .ZN(n8615) );
  XNOR2_X1 U10045 ( .A(n8612), .B(n8618), .ZN(n8613) );
  OAI222_X1 U10046 ( .A1(n8762), .A2(n6273), .B1(n8761), .B2(n8614), .C1(n8613), .C2(n8629), .ZN(n8850) );
  AOI211_X1 U10047 ( .C1(n8748), .C2(n8616), .A(n8615), .B(n8850), .ZN(n8622)
         );
  XOR2_X1 U10048 ( .A(n8618), .B(n8617), .Z(n8856) );
  INV_X1 U10049 ( .A(n8856), .ZN(n8620) );
  AOI22_X1 U10050 ( .A1(n8620), .A2(n8619), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n8725), .ZN(n8621) );
  OAI21_X1 U10051 ( .B1(n8622), .B2(n8725), .A(n8621), .ZN(P2_U3208) );
  NAND2_X1 U10052 ( .A1(n8624), .A2(n8623), .ZN(n8625) );
  XNOR2_X1 U10053 ( .A(n8625), .B(n8627), .ZN(n8862) );
  XOR2_X1 U10054 ( .A(n8627), .B(n8626), .Z(n8628) );
  OAI222_X1 U10055 ( .A1(n8762), .A2(n8631), .B1(n8761), .B2(n8630), .C1(n8629), .C2(n8628), .ZN(n8796) );
  INV_X1 U10056 ( .A(n8796), .ZN(n8857) );
  OAI21_X1 U10057 ( .B1(n8798), .B2(n8632), .A(n8857), .ZN(n8633) );
  NAND2_X1 U10058 ( .A1(n8633), .A2(n8745), .ZN(n8636) );
  AOI22_X1 U10059 ( .A1(n8748), .A2(n8634), .B1(n8725), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n8635) );
  OAI211_X1 U10060 ( .C1(n8862), .C2(n8752), .A(n8636), .B(n8635), .ZN(
        P2_U3209) );
  XOR2_X1 U10061 ( .A(n8637), .B(n8638), .Z(n8868) );
  INV_X1 U10062 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n9881) );
  XNOR2_X1 U10063 ( .A(n8639), .B(n8638), .ZN(n8641) );
  AOI222_X1 U10064 ( .A1(n8765), .A2(n8641), .B1(n8640), .B2(n5047), .C1(n8664), .C2(n8741), .ZN(n8863) );
  MUX2_X1 U10065 ( .A(n9881), .B(n8863), .S(n8745), .Z(n8644) );
  AOI22_X1 U10066 ( .A1(n8865), .A2(n8749), .B1(n8748), .B2(n8642), .ZN(n8643)
         );
  OAI211_X1 U10067 ( .C1(n8868), .C2(n8752), .A(n8644), .B(n8643), .ZN(
        P2_U3210) );
  XNOR2_X1 U10068 ( .A(n8645), .B(n8648), .ZN(n8874) );
  INV_X1 U10069 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8653) );
  NAND3_X1 U10070 ( .A1(n8646), .A2(n8648), .A3(n8647), .ZN(n8649) );
  NAND2_X1 U10071 ( .A1(n8650), .A2(n8649), .ZN(n8652) );
  AOI222_X1 U10072 ( .A1(n8765), .A2(n8652), .B1(n8651), .B2(n5047), .C1(n8676), .C2(n8741), .ZN(n8869) );
  MUX2_X1 U10073 ( .A(n8653), .B(n8869), .S(n8745), .Z(n8656) );
  AOI22_X1 U10074 ( .A1(n8871), .A2(n8749), .B1(n8748), .B2(n8654), .ZN(n8655)
         );
  OAI211_X1 U10075 ( .C1(n8874), .C2(n8752), .A(n8656), .B(n8655), .ZN(
        P2_U3211) );
  XNOR2_X1 U10076 ( .A(n8658), .B(n8657), .ZN(n8880) );
  INV_X1 U10077 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8666) );
  NAND3_X1 U10078 ( .A1(n8659), .A2(n8661), .A3(n8660), .ZN(n8662) );
  NAND2_X1 U10079 ( .A1(n8646), .A2(n8662), .ZN(n8665) );
  AOI222_X1 U10080 ( .A1(n8765), .A2(n8665), .B1(n8664), .B2(n5047), .C1(n8663), .C2(n8741), .ZN(n8875) );
  MUX2_X1 U10081 ( .A(n8666), .B(n8875), .S(n8745), .Z(n8669) );
  AOI22_X1 U10082 ( .A1(n8877), .A2(n8749), .B1(n8748), .B2(n8667), .ZN(n8668)
         );
  OAI211_X1 U10083 ( .C1(n8880), .C2(n8752), .A(n8669), .B(n8668), .ZN(
        P2_U3212) );
  NAND2_X1 U10084 ( .A1(n8685), .A2(n8670), .ZN(n8672) );
  XNOR2_X1 U10085 ( .A(n8672), .B(n8671), .ZN(n8886) );
  AND2_X1 U10086 ( .A1(n8690), .A2(n8673), .ZN(n8675) );
  OAI21_X1 U10087 ( .B1(n8675), .B2(n8674), .A(n8659), .ZN(n8677) );
  AOI222_X1 U10088 ( .A1(n8765), .A2(n8677), .B1(n8676), .B2(n5047), .C1(n8706), .C2(n8741), .ZN(n8881) );
  MUX2_X1 U10089 ( .A(n8678), .B(n8881), .S(n8745), .Z(n8681) );
  AOI22_X1 U10090 ( .A1(n8883), .A2(n8749), .B1(n8748), .B2(n8679), .ZN(n8680)
         );
  OAI211_X1 U10091 ( .C1(n8886), .C2(n8752), .A(n8681), .B(n8680), .ZN(
        P2_U3213) );
  NAND2_X1 U10092 ( .A1(n8718), .A2(n8682), .ZN(n8684) );
  NAND2_X1 U10093 ( .A1(n8684), .A2(n8683), .ZN(n8686) );
  OAI21_X1 U10094 ( .B1(n8686), .B2(n8688), .A(n8685), .ZN(n8892) );
  NAND2_X1 U10095 ( .A1(n8704), .A2(n8687), .ZN(n8689) );
  NAND2_X1 U10096 ( .A1(n8689), .A2(n8688), .ZN(n8691) );
  NAND3_X1 U10097 ( .A1(n8691), .A2(n8765), .A3(n8690), .ZN(n8696) );
  OAI22_X1 U10098 ( .A1(n8693), .A2(n8762), .B1(n8692), .B2(n8761), .ZN(n8694)
         );
  INV_X1 U10099 ( .A(n8694), .ZN(n8695) );
  AND2_X1 U10100 ( .A1(n8696), .A2(n8695), .ZN(n8887) );
  MUX2_X1 U10101 ( .A(n8697), .B(n8887), .S(n8745), .Z(n8700) );
  AOI22_X1 U10102 ( .A1(n8889), .A2(n8749), .B1(n8748), .B2(n8698), .ZN(n8699)
         );
  OAI211_X1 U10103 ( .C1(n8892), .C2(n8752), .A(n8700), .B(n8699), .ZN(
        P2_U3214) );
  NAND2_X1 U10104 ( .A1(n8718), .A2(n8701), .ZN(n8702) );
  XOR2_X1 U10105 ( .A(n8703), .B(n8702), .Z(n8897) );
  OAI21_X1 U10106 ( .B1(n8705), .B2(n5453), .A(n8704), .ZN(n8707) );
  AOI222_X1 U10107 ( .A1(n8765), .A2(n8707), .B1(n8706), .B2(n5047), .C1(n8731), .C2(n8741), .ZN(n8893) );
  MUX2_X1 U10108 ( .A(n8708), .B(n8893), .S(n8745), .Z(n8711) );
  AOI22_X1 U10109 ( .A1(n8894), .A2(n8749), .B1(n8748), .B2(n8709), .ZN(n8710)
         );
  OAI211_X1 U10110 ( .C1(n8897), .C2(n8752), .A(n8711), .B(n8710), .ZN(
        P2_U3215) );
  XNOR2_X1 U10111 ( .A(n8712), .B(n8713), .ZN(n8715) );
  AOI222_X1 U10112 ( .A1(n8765), .A2(n8715), .B1(n8714), .B2(n5047), .C1(n8743), .C2(n8741), .ZN(n8820) );
  OAI22_X1 U10113 ( .A1(n8745), .A2(n8717), .B1(n8716), .B2(n8771), .ZN(n8723)
         );
  INV_X1 U10114 ( .A(n8718), .ZN(n8719) );
  AOI21_X1 U10115 ( .B1(n8721), .B2(n8720), .A(n8719), .ZN(n8821) );
  NOR2_X1 U10116 ( .A1(n8821), .A2(n8752), .ZN(n8722) );
  AOI211_X1 U10117 ( .C1(n8749), .C2(n8818), .A(n8723), .B(n8722), .ZN(n8724)
         );
  OAI21_X1 U10118 ( .B1(n8725), .B2(n8820), .A(n8724), .ZN(P2_U3216) );
  XNOR2_X1 U10119 ( .A(n8727), .B(n8726), .ZN(n8904) );
  XNOR2_X1 U10120 ( .A(n8729), .B(n8728), .ZN(n8732) );
  AOI222_X1 U10121 ( .A1(n8765), .A2(n8732), .B1(n8731), .B2(n5047), .C1(n8730), .C2(n8741), .ZN(n8899) );
  MUX2_X1 U10122 ( .A(n8733), .B(n8899), .S(n8745), .Z(n8737) );
  INV_X1 U10123 ( .A(n8734), .ZN(n8735) );
  AOI22_X1 U10124 ( .A1(n8901), .A2(n8749), .B1(n8748), .B2(n8735), .ZN(n8736)
         );
  OAI211_X1 U10125 ( .C1(n8904), .C2(n8752), .A(n8737), .B(n8736), .ZN(
        P2_U3217) );
  XNOR2_X1 U10126 ( .A(n8738), .B(n8739), .ZN(n8911) );
  XNOR2_X1 U10127 ( .A(n8740), .B(n8739), .ZN(n8744) );
  AOI222_X1 U10128 ( .A1(n8765), .A2(n8744), .B1(n8743), .B2(n5047), .C1(n8742), .C2(n8741), .ZN(n8905) );
  MUX2_X1 U10129 ( .A(n8746), .B(n8905), .S(n8745), .Z(n8751) );
  AOI22_X1 U10130 ( .A1(n8907), .A2(n8749), .B1(n8748), .B2(n8747), .ZN(n8750)
         );
  OAI211_X1 U10131 ( .C1(n8911), .C2(n8752), .A(n8751), .B(n8750), .ZN(
        P2_U3218) );
  OAI21_X1 U10132 ( .B1(n8754), .B2(n8757), .A(n8753), .ZN(n10242) );
  NAND2_X1 U10133 ( .A1(n10242), .A2(n8755), .ZN(n8768) );
  NAND3_X1 U10134 ( .A1(n8758), .A2(n8757), .A3(n8756), .ZN(n8759) );
  NAND2_X1 U10135 ( .A1(n8760), .A2(n8759), .ZN(n8766) );
  OAI22_X1 U10136 ( .A1(n8763), .A2(n8762), .B1(n6187), .B2(n8761), .ZN(n8764)
         );
  AOI21_X1 U10137 ( .B1(n8766), .B2(n8765), .A(n8764), .ZN(n8767) );
  AND2_X1 U10138 ( .A1(n8768), .A2(n8767), .ZN(n10244) );
  NAND2_X1 U10139 ( .A1(n10240), .A2(n8769), .ZN(n8770) );
  OAI21_X1 U10140 ( .B1(n6728), .B2(n8771), .A(n8770), .ZN(n8772) );
  AOI21_X1 U10141 ( .B1(n10242), .B2(n8773), .A(n8772), .ZN(n8774) );
  NAND2_X1 U10142 ( .A1(n10244), .A2(n8774), .ZN(n8775) );
  MUX2_X1 U10143 ( .A(n8775), .B(P2_REG2_REG_2__SCAN_IN), .S(n8725), .Z(
        P2_U3231) );
  NAND2_X1 U10144 ( .A1(n8831), .A2(n8826), .ZN(n8777) );
  INV_X1 U10145 ( .A(n8776), .ZN(n8832) );
  NAND2_X1 U10146 ( .A1(n8832), .A2(n10303), .ZN(n8779) );
  OAI211_X1 U10147 ( .C1(n10303), .C2(n8178), .A(n8777), .B(n8779), .ZN(
        P2_U3490) );
  NAND2_X1 U10148 ( .A1(n6312), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8778) );
  OAI211_X1 U10149 ( .C1(n8780), .C2(n8797), .A(n8779), .B(n8778), .ZN(
        P2_U3489) );
  MUX2_X1 U10150 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8781), .S(n10303), .Z(
        n8785) );
  OAI22_X1 U10151 ( .A1(n8783), .A2(n8829), .B1(n8782), .B2(n8797), .ZN(n8784)
         );
  OR2_X1 U10152 ( .A1(n8785), .A2(n8784), .ZN(P2_U3487) );
  AOI21_X1 U10153 ( .B1(n8787), .B2(n10279), .A(n8786), .ZN(n8839) );
  MUX2_X1 U10154 ( .A(n9900), .B(n8839), .S(n10303), .Z(n8788) );
  OAI21_X1 U10155 ( .B1(n8843), .B2(n8797), .A(n8788), .ZN(P2_U3486) );
  MUX2_X1 U10156 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8789), .S(n10303), .Z(
        n8792) );
  OAI22_X1 U10157 ( .A1(n8849), .A2(n8829), .B1(n8790), .B2(n8797), .ZN(n8791)
         );
  OR2_X1 U10158 ( .A1(n8792), .A2(n8791), .ZN(P2_U3485) );
  OAI22_X1 U10159 ( .A1(n8856), .A2(n8829), .B1(n8793), .B2(n8797), .ZN(n8795)
         );
  MUX2_X1 U10160 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8850), .S(n10303), .Z(
        n8794) );
  OR2_X1 U10161 ( .A1(n8795), .A2(n8794), .ZN(P2_U3484) );
  MUX2_X1 U10162 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8796), .S(n10303), .Z(
        n8800) );
  OAI22_X1 U10163 ( .A1(n8862), .A2(n8829), .B1(n8798), .B2(n8797), .ZN(n8799)
         );
  OR2_X1 U10164 ( .A1(n8800), .A2(n8799), .ZN(P2_U3483) );
  INV_X1 U10165 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8801) );
  MUX2_X1 U10166 ( .A(n8801), .B(n8863), .S(n10303), .Z(n8803) );
  NAND2_X1 U10167 ( .A1(n8865), .A2(n8826), .ZN(n8802) );
  OAI211_X1 U10168 ( .C1(n8868), .C2(n8829), .A(n8803), .B(n8802), .ZN(
        P2_U3482) );
  INV_X1 U10169 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8804) );
  MUX2_X1 U10170 ( .A(n8804), .B(n8869), .S(n10303), .Z(n8806) );
  NAND2_X1 U10171 ( .A1(n8871), .A2(n8826), .ZN(n8805) );
  OAI211_X1 U10172 ( .C1(n8874), .C2(n8829), .A(n8806), .B(n8805), .ZN(
        P2_U3481) );
  INV_X1 U10173 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8807) );
  MUX2_X1 U10174 ( .A(n8807), .B(n8875), .S(n10303), .Z(n8809) );
  NAND2_X1 U10175 ( .A1(n8877), .A2(n8826), .ZN(n8808) );
  OAI211_X1 U10176 ( .C1(n8829), .C2(n8880), .A(n8809), .B(n8808), .ZN(
        P2_U3480) );
  MUX2_X1 U10177 ( .A(n8810), .B(n8881), .S(n10303), .Z(n8812) );
  NAND2_X1 U10178 ( .A1(n8883), .A2(n8826), .ZN(n8811) );
  OAI211_X1 U10179 ( .C1(n8886), .C2(n8829), .A(n8812), .B(n8811), .ZN(
        P2_U3479) );
  MUX2_X1 U10180 ( .A(n9730), .B(n8887), .S(n10303), .Z(n8814) );
  NAND2_X1 U10181 ( .A1(n8889), .A2(n8826), .ZN(n8813) );
  OAI211_X1 U10182 ( .C1(n8829), .C2(n8892), .A(n8814), .B(n8813), .ZN(
        P2_U3478) );
  MUX2_X1 U10183 ( .A(n8815), .B(n8893), .S(n10303), .Z(n8817) );
  NAND2_X1 U10184 ( .A1(n8894), .A2(n8826), .ZN(n8816) );
  OAI211_X1 U10185 ( .C1(n8829), .C2(n8897), .A(n8817), .B(n8816), .ZN(
        P2_U3477) );
  NAND2_X1 U10186 ( .A1(n8818), .A2(n10281), .ZN(n8819) );
  OAI211_X1 U10187 ( .C1(n8821), .C2(n10247), .A(n8820), .B(n8819), .ZN(n8898)
         );
  MUX2_X1 U10188 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8898), .S(n10303), .Z(
        P2_U3476) );
  MUX2_X1 U10189 ( .A(n8822), .B(n8899), .S(n10303), .Z(n8824) );
  NAND2_X1 U10190 ( .A1(n8901), .A2(n8826), .ZN(n8823) );
  OAI211_X1 U10191 ( .C1(n8829), .C2(n8904), .A(n8824), .B(n8823), .ZN(
        P2_U3475) );
  MUX2_X1 U10192 ( .A(n8825), .B(n8905), .S(n10303), .Z(n8828) );
  NAND2_X1 U10193 ( .A1(n8907), .A2(n8826), .ZN(n8827) );
  OAI211_X1 U10194 ( .C1(n8911), .C2(n8829), .A(n8828), .B(n8827), .ZN(
        P2_U3474) );
  MUX2_X1 U10195 ( .A(n8830), .B(P2_REG1_REG_0__SCAN_IN), .S(n6312), .Z(
        P2_U3459) );
  INV_X1 U10196 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8834) );
  NAND2_X1 U10197 ( .A1(n8831), .A2(n5698), .ZN(n8833) );
  NAND2_X1 U10198 ( .A1(n8832), .A2(n10286), .ZN(n8836) );
  OAI211_X1 U10199 ( .C1(n8834), .C2(n10286), .A(n8833), .B(n8836), .ZN(
        P2_U3458) );
  INV_X1 U10200 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8838) );
  NAND2_X1 U10201 ( .A1(n8835), .A2(n5698), .ZN(n8837) );
  OAI211_X1 U10202 ( .C1(n8838), .C2(n10286), .A(n8837), .B(n8836), .ZN(
        P2_U3457) );
  INV_X1 U10203 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8840) );
  MUX2_X1 U10204 ( .A(n8840), .B(n8839), .S(n10286), .Z(n8841) );
  OAI21_X1 U10205 ( .B1(n8843), .B2(n8842), .A(n8841), .ZN(P2_U3454) );
  MUX2_X1 U10206 ( .A(n8845), .B(n8844), .S(n10286), .Z(n8848) );
  NAND2_X1 U10207 ( .A1(n8846), .A2(n5698), .ZN(n8847) );
  OAI211_X1 U10208 ( .C1(n8849), .C2(n8910), .A(n8848), .B(n8847), .ZN(
        P2_U3453) );
  INV_X1 U10209 ( .A(n8850), .ZN(n8851) );
  MUX2_X1 U10210 ( .A(n8852), .B(n8851), .S(n10286), .Z(n8855) );
  NAND2_X1 U10211 ( .A1(n8853), .A2(n5698), .ZN(n8854) );
  OAI211_X1 U10212 ( .C1(n8856), .C2(n8910), .A(n8855), .B(n8854), .ZN(
        P2_U3452) );
  MUX2_X1 U10213 ( .A(n8858), .B(n8857), .S(n10286), .Z(n8861) );
  NAND2_X1 U10214 ( .A1(n8859), .A2(n5698), .ZN(n8860) );
  OAI211_X1 U10215 ( .C1(n8862), .C2(n8910), .A(n8861), .B(n8860), .ZN(
        P2_U3451) );
  MUX2_X1 U10216 ( .A(n8864), .B(n8863), .S(n10286), .Z(n8867) );
  NAND2_X1 U10217 ( .A1(n8865), .A2(n5698), .ZN(n8866) );
  OAI211_X1 U10218 ( .C1(n8868), .C2(n8910), .A(n8867), .B(n8866), .ZN(
        P2_U3450) );
  MUX2_X1 U10219 ( .A(n8870), .B(n8869), .S(n10286), .Z(n8873) );
  NAND2_X1 U10220 ( .A1(n8871), .A2(n5698), .ZN(n8872) );
  OAI211_X1 U10221 ( .C1(n8874), .C2(n8910), .A(n8873), .B(n8872), .ZN(
        P2_U3449) );
  MUX2_X1 U10222 ( .A(n8876), .B(n8875), .S(n10286), .Z(n8879) );
  NAND2_X1 U10223 ( .A1(n8877), .A2(n5698), .ZN(n8878) );
  OAI211_X1 U10224 ( .C1(n8880), .C2(n8910), .A(n8879), .B(n8878), .ZN(
        P2_U3448) );
  INV_X1 U10225 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8882) );
  MUX2_X1 U10226 ( .A(n8882), .B(n8881), .S(n10286), .Z(n8885) );
  NAND2_X1 U10227 ( .A1(n8883), .A2(n5698), .ZN(n8884) );
  OAI211_X1 U10228 ( .C1(n8886), .C2(n8910), .A(n8885), .B(n8884), .ZN(
        P2_U3447) );
  MUX2_X1 U10229 ( .A(n8888), .B(n8887), .S(n10286), .Z(n8891) );
  NAND2_X1 U10230 ( .A1(n8889), .A2(n5698), .ZN(n8890) );
  OAI211_X1 U10231 ( .C1(n8892), .C2(n8910), .A(n8891), .B(n8890), .ZN(
        P2_U3446) );
  MUX2_X1 U10232 ( .A(n9796), .B(n8893), .S(n10286), .Z(n8896) );
  NAND2_X1 U10233 ( .A1(n8894), .A2(n5698), .ZN(n8895) );
  OAI211_X1 U10234 ( .C1(n8897), .C2(n8910), .A(n8896), .B(n8895), .ZN(
        P2_U3444) );
  MUX2_X1 U10235 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8898), .S(n10286), .Z(
        P2_U3441) );
  INV_X1 U10236 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8900) );
  MUX2_X1 U10237 ( .A(n8900), .B(n8899), .S(n10286), .Z(n8903) );
  NAND2_X1 U10238 ( .A1(n8901), .A2(n5698), .ZN(n8902) );
  OAI211_X1 U10239 ( .C1(n8904), .C2(n8910), .A(n8903), .B(n8902), .ZN(
        P2_U3438) );
  INV_X1 U10240 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8906) );
  MUX2_X1 U10241 ( .A(n8906), .B(n8905), .S(n10286), .Z(n8909) );
  NAND2_X1 U10242 ( .A1(n8907), .A2(n5698), .ZN(n8908) );
  OAI211_X1 U10243 ( .C1(n8911), .C2(n8910), .A(n8909), .B(n8908), .ZN(
        P2_U3435) );
  INV_X1 U10244 ( .A(n8912), .ZN(n9964) );
  NOR4_X1 U10245 ( .A1(n8914), .A2(P2_IR_REG_30__SCAN_IN), .A3(n8913), .A4(
        P2_U3151), .ZN(n8915) );
  AOI21_X1 U10246 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n8916), .A(n8915), .ZN(
        n8917) );
  OAI21_X1 U10247 ( .B1(n9964), .B2(n8918), .A(n8917), .ZN(P2_U3264) );
  MUX2_X1 U10248 ( .A(n8919), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  NOR2_X1 U10249 ( .A1(n8920), .A2(n9065), .ZN(n8921) );
  AOI21_X1 U10250 ( .B1(n9202), .B2(n7541), .A(n8921), .ZN(n9115) );
  NAND2_X1 U10251 ( .A1(n9202), .A2(n9070), .ZN(n8923) );
  NAND2_X1 U10252 ( .A1(n4655), .A2(n7541), .ZN(n8922) );
  NAND2_X1 U10253 ( .A1(n8923), .A2(n8922), .ZN(n8924) );
  XNOR2_X1 U10254 ( .A(n8924), .B(n9068), .ZN(n9117) );
  NOR2_X1 U10255 ( .A1(n8926), .A2(n8925), .ZN(n8930) );
  INV_X1 U10256 ( .A(n8926), .ZN(n8928) );
  OAI22_X2 U10257 ( .A1(n8930), .A2(n8929), .B1(n8928), .B2(n8927), .ZN(n9116)
         );
  NAND2_X1 U10258 ( .A1(n9126), .A2(n9070), .ZN(n8932) );
  NAND2_X1 U10259 ( .A1(n9218), .A2(n7541), .ZN(n8931) );
  NAND2_X1 U10260 ( .A1(n8932), .A2(n8931), .ZN(n8933) );
  XNOR2_X1 U10261 ( .A(n8933), .B(n8997), .ZN(n9118) );
  OAI22_X1 U10262 ( .A1(n9957), .A2(n4394), .B1(n9132), .B2(n9065), .ZN(n8935)
         );
  NAND2_X1 U10263 ( .A1(n9118), .A2(n8935), .ZN(n8934) );
  OAI211_X1 U10264 ( .C1(n9115), .C2(n9117), .A(n9116), .B(n8934), .ZN(n8940)
         );
  INV_X1 U10265 ( .A(n8935), .ZN(n9119) );
  AOI21_X1 U10266 ( .B1(n9117), .B2(n9115), .A(n9119), .ZN(n8936) );
  NAND3_X1 U10267 ( .A1(n9119), .A2(n9115), .A3(n9117), .ZN(n8937) );
  OAI22_X1 U10268 ( .A1(n9544), .A2(n4394), .B1(n8941), .B2(n9065), .ZN(n8946)
         );
  NAND2_X1 U10269 ( .A1(n9636), .A2(n9070), .ZN(n8943) );
  NAND2_X1 U10270 ( .A1(n9217), .A2(n7541), .ZN(n8942) );
  NAND2_X1 U10271 ( .A1(n8943), .A2(n8942), .ZN(n8944) );
  XNOR2_X1 U10272 ( .A(n8944), .B(n8997), .ZN(n8945) );
  XOR2_X1 U10273 ( .A(n8946), .B(n8945), .Z(n9130) );
  INV_X1 U10274 ( .A(n8945), .ZN(n8948) );
  INV_X1 U10275 ( .A(n8946), .ZN(n8947) );
  NAND2_X1 U10276 ( .A1(n8948), .A2(n8947), .ZN(n8949) );
  AOI22_X1 U10277 ( .A1(n9531), .A2(n9070), .B1(n7541), .B2(n9216), .ZN(n8950)
         );
  XNOR2_X1 U10278 ( .A(n8950), .B(n8997), .ZN(n8953) );
  AND2_X1 U10279 ( .A1(n9216), .A2(n9002), .ZN(n8952) );
  AOI21_X1 U10280 ( .B1(n9531), .B2(n7541), .A(n8952), .ZN(n9171) );
  NAND2_X1 U10281 ( .A1(n9167), .A2(n9171), .ZN(n8955) );
  NAND2_X1 U10282 ( .A1(n8955), .A2(n9168), .ZN(n9058) );
  NAND2_X1 U10283 ( .A1(n9625), .A2(n9070), .ZN(n8957) );
  INV_X1 U10284 ( .A(n9175), .ZN(n9215) );
  NAND2_X1 U10285 ( .A1(n9215), .A2(n7541), .ZN(n8956) );
  NAND2_X1 U10286 ( .A1(n8957), .A2(n8956), .ZN(n8958) );
  XNOR2_X1 U10287 ( .A(n8958), .B(n9068), .ZN(n8961) );
  NOR2_X1 U10288 ( .A1(n9175), .A2(n9065), .ZN(n8959) );
  AOI21_X1 U10289 ( .B1(n9625), .B2(n7541), .A(n8959), .ZN(n8960) );
  OR2_X1 U10290 ( .A1(n8961), .A2(n8960), .ZN(n9056) );
  NAND2_X1 U10291 ( .A1(n9058), .A2(n9056), .ZN(n8962) );
  NAND2_X1 U10292 ( .A1(n8961), .A2(n8960), .ZN(n9055) );
  OAI22_X1 U10293 ( .A1(n9946), .A2(n4394), .B1(n9060), .B2(n9065), .ZN(n8965)
         );
  OAI22_X1 U10294 ( .A1(n9946), .A2(n8996), .B1(n9060), .B2(n4394), .ZN(n8963)
         );
  XNOR2_X1 U10295 ( .A(n8963), .B(n8997), .ZN(n8964) );
  XOR2_X1 U10296 ( .A(n8965), .B(n8964), .Z(n9148) );
  INV_X1 U10297 ( .A(n8964), .ZN(n8967) );
  INV_X1 U10298 ( .A(n8965), .ZN(n8966) );
  NAND2_X1 U10299 ( .A1(n8967), .A2(n8966), .ZN(n8968) );
  OAI22_X1 U10300 ( .A1(n9942), .A2(n4394), .B1(n9160), .B2(n9065), .ZN(n8973)
         );
  NAND2_X1 U10301 ( .A1(n9486), .A2(n9070), .ZN(n8970) );
  NAND2_X1 U10302 ( .A1(n9213), .A2(n7541), .ZN(n8969) );
  NAND2_X1 U10303 ( .A1(n8970), .A2(n8969), .ZN(n8971) );
  XNOR2_X1 U10304 ( .A(n8971), .B(n8997), .ZN(n8972) );
  XOR2_X1 U10305 ( .A(n8973), .B(n8972), .Z(n9098) );
  INV_X1 U10306 ( .A(n8972), .ZN(n8975) );
  INV_X1 U10307 ( .A(n8973), .ZN(n8974) );
  NAND2_X1 U10308 ( .A1(n9474), .A2(n9070), .ZN(n8977) );
  NAND2_X1 U10309 ( .A1(n9212), .A2(n7541), .ZN(n8976) );
  NAND2_X1 U10310 ( .A1(n8977), .A2(n8976), .ZN(n8978) );
  XNOR2_X1 U10311 ( .A(n8978), .B(n8997), .ZN(n8980) );
  XNOR2_X1 U10312 ( .A(n8979), .B(n8980), .ZN(n9158) );
  AOI22_X1 U10313 ( .A1(n9474), .A2(n7541), .B1(n9002), .B2(n9212), .ZN(n9159)
         );
  INV_X1 U10314 ( .A(n8979), .ZN(n8981) );
  OAI22_X1 U10315 ( .A1(n9456), .A2(n8996), .B1(n9161), .B2(n4394), .ZN(n8983)
         );
  XNOR2_X1 U10316 ( .A(n8983), .B(n8997), .ZN(n8986) );
  OR2_X1 U10317 ( .A1(n9456), .A2(n4394), .ZN(n8985) );
  OR2_X1 U10318 ( .A1(n9161), .A2(n9065), .ZN(n8984) );
  NAND2_X1 U10319 ( .A1(n8985), .A2(n8984), .ZN(n8987) );
  NAND2_X1 U10320 ( .A1(n8986), .A2(n8987), .ZN(n9032) );
  NAND2_X1 U10321 ( .A1(n9035), .A2(n9032), .ZN(n8990) );
  INV_X1 U10322 ( .A(n8986), .ZN(n8989) );
  INV_X1 U10323 ( .A(n8987), .ZN(n8988) );
  NAND2_X1 U10324 ( .A1(n8989), .A2(n8988), .ZN(n9033) );
  AOI22_X1 U10325 ( .A1(n9443), .A2(n9070), .B1(n7541), .B2(n9211), .ZN(n8991)
         );
  XOR2_X1 U10326 ( .A(n8997), .B(n8991), .Z(n8993) );
  OAI22_X1 U10327 ( .A1(n4703), .A2(n4394), .B1(n9037), .B2(n9065), .ZN(n8992)
         );
  NOR2_X1 U10328 ( .A1(n8993), .A2(n8992), .ZN(n8994) );
  AOI21_X1 U10329 ( .B1(n8993), .B2(n8992), .A(n8994), .ZN(n9139) );
  INV_X1 U10330 ( .A(n8994), .ZN(n8995) );
  OAI22_X1 U10331 ( .A1(n9663), .A2(n4394), .B1(n9186), .B2(n9065), .ZN(n9004)
         );
  OAI22_X1 U10332 ( .A1(n9663), .A2(n8996), .B1(n9186), .B2(n4394), .ZN(n8998)
         );
  XNOR2_X1 U10333 ( .A(n8998), .B(n8997), .ZN(n9005) );
  XOR2_X1 U10334 ( .A(n9004), .B(n9005), .Z(n9107) );
  NAND2_X1 U10335 ( .A1(n9590), .A2(n9070), .ZN(n9000) );
  NAND2_X1 U10336 ( .A1(n9209), .A2(n7541), .ZN(n8999) );
  NAND2_X1 U10337 ( .A1(n9000), .A2(n8999), .ZN(n9001) );
  XNOR2_X1 U10338 ( .A(n9001), .B(n9068), .ZN(n9007) );
  AND2_X1 U10339 ( .A1(n9209), .A2(n9002), .ZN(n9003) );
  AOI21_X1 U10340 ( .B1(n9590), .B2(n7541), .A(n9003), .ZN(n9008) );
  XNOR2_X1 U10341 ( .A(n9007), .B(n9008), .ZN(n9180) );
  NOR2_X1 U10342 ( .A1(n9005), .A2(n9004), .ZN(n9181) );
  NOR2_X1 U10343 ( .A1(n9180), .A2(n9181), .ZN(n9006) );
  INV_X1 U10344 ( .A(n9007), .ZN(n9010) );
  INV_X1 U10345 ( .A(n9008), .ZN(n9009) );
  NAND2_X1 U10346 ( .A1(n9010), .A2(n9009), .ZN(n9020) );
  NAND2_X1 U10347 ( .A1(n9389), .A2(n9070), .ZN(n9012) );
  INV_X1 U10348 ( .A(n9187), .ZN(n9208) );
  NAND2_X1 U10349 ( .A1(n9208), .A2(n7541), .ZN(n9011) );
  NAND2_X1 U10350 ( .A1(n9012), .A2(n9011), .ZN(n9013) );
  XNOR2_X1 U10351 ( .A(n9013), .B(n9068), .ZN(n9016) );
  INV_X1 U10352 ( .A(n9016), .ZN(n9018) );
  NOR2_X1 U10353 ( .A1(n9187), .A2(n9065), .ZN(n9014) );
  AOI21_X1 U10354 ( .B1(n9389), .B2(n7541), .A(n9014), .ZN(n9015) );
  INV_X1 U10355 ( .A(n9015), .ZN(n9017) );
  AOI21_X1 U10356 ( .B1(n9018), .B2(n9017), .A(n9081), .ZN(n9019) );
  AOI21_X1 U10357 ( .B1(n9183), .B2(n9020), .A(n9019), .ZN(n9024) );
  INV_X1 U10358 ( .A(n9019), .ZN(n9022) );
  INV_X1 U10359 ( .A(n9020), .ZN(n9021) );
  NOR2_X1 U10360 ( .A1(n9022), .A2(n9021), .ZN(n9023) );
  OAI21_X1 U10361 ( .B1(n9024), .B2(n9075), .A(n9184), .ZN(n9031) );
  OR2_X1 U10362 ( .A1(n9372), .A2(n9350), .ZN(n9026) );
  NAND2_X1 U10363 ( .A1(n9209), .A2(n9173), .ZN(n9025) );
  AND2_X1 U10364 ( .A1(n9026), .A2(n9025), .ZN(n9397) );
  INV_X1 U10365 ( .A(n9391), .ZN(n9027) );
  AOI22_X1 U10366 ( .A1(n9027), .A2(n9145), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n9028) );
  OAI21_X1 U10367 ( .B1(n9397), .B2(n9143), .A(n9028), .ZN(n9029) );
  AOI21_X1 U10368 ( .B1(n9389), .B2(n9201), .A(n9029), .ZN(n9030) );
  NAND2_X1 U10369 ( .A1(n9031), .A2(n9030), .ZN(P1_U3214) );
  NAND2_X1 U10370 ( .A1(n9033), .A2(n9032), .ZN(n9034) );
  XNOR2_X1 U10371 ( .A(n9035), .B(n9034), .ZN(n9043) );
  OAI22_X1 U10372 ( .A1(n9037), .A2(n9350), .B1(n9036), .B2(n9373), .ZN(n9460)
         );
  INV_X1 U10373 ( .A(n9460), .ZN(n9040) );
  INV_X1 U10374 ( .A(n9038), .ZN(n9454) );
  AOI22_X1 U10375 ( .A1(n9454), .A2(n9145), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n9039) );
  OAI21_X1 U10376 ( .B1(n9040), .B2(n9143), .A(n9039), .ZN(n9041) );
  AOI21_X1 U10377 ( .B1(n6126), .B2(n9201), .A(n9041), .ZN(n9042) );
  OAI21_X1 U10378 ( .B1(n9043), .B2(n9204), .A(n9042), .ZN(P1_U3216) );
  OAI21_X1 U10379 ( .B1(n9046), .B2(n9045), .A(n9044), .ZN(n9047) );
  NAND2_X1 U10380 ( .A1(n9047), .A2(n9184), .ZN(n9054) );
  AOI22_X1 U10381 ( .A1(n9048), .A2(n9195), .B1(P1_REG3_REG_10__SCAN_IN), .B2(
        P1_U3086), .ZN(n9053) );
  NAND2_X1 U10382 ( .A1(n9049), .A2(n9201), .ZN(n9052) );
  NAND2_X1 U10383 ( .A1(n9145), .A2(n9050), .ZN(n9051) );
  NAND4_X1 U10384 ( .A1(n9054), .A2(n9053), .A3(n9052), .A4(n9051), .ZN(
        P1_U3217) );
  NAND2_X1 U10385 ( .A1(n9056), .A2(n9055), .ZN(n9057) );
  XNOR2_X1 U10386 ( .A(n9058), .B(n9057), .ZN(n9064) );
  NAND2_X1 U10387 ( .A1(n9216), .A2(n9173), .ZN(n9059) );
  OAI21_X1 U10388 ( .B1(n9060), .B2(n9350), .A(n9059), .ZN(n9514) );
  NAND2_X1 U10389 ( .A1(n9514), .A2(n9195), .ZN(n9061) );
  NAND2_X1 U10390 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9345) );
  OAI211_X1 U10391 ( .C1(n9198), .C2(n9519), .A(n9061), .B(n9345), .ZN(n9062)
         );
  AOI21_X1 U10392 ( .B1(n9625), .B2(n9201), .A(n9062), .ZN(n9063) );
  OAI21_X1 U10393 ( .B1(n9064), .B2(n9204), .A(n9063), .ZN(P1_U3219) );
  NAND2_X1 U10394 ( .A1(n9071), .A2(n7541), .ZN(n9067) );
  OR2_X1 U10395 ( .A1(n9372), .A2(n9065), .ZN(n9066) );
  NAND2_X1 U10396 ( .A1(n9067), .A2(n9066), .ZN(n9069) );
  XNOR2_X1 U10397 ( .A(n9069), .B(n9068), .ZN(n9074) );
  NAND2_X1 U10398 ( .A1(n9071), .A2(n9070), .ZN(n9072) );
  OAI21_X1 U10399 ( .B1(n9372), .B2(n4394), .A(n9072), .ZN(n9073) );
  XNOR2_X1 U10400 ( .A(n9074), .B(n9073), .ZN(n9082) );
  NAND3_X1 U10401 ( .A1(n9075), .A2(n9184), .A3(n9082), .ZN(n9085) );
  INV_X1 U10402 ( .A(n9076), .ZN(n9077) );
  OAI22_X1 U10403 ( .A1(n9077), .A2(n9198), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9378), .ZN(n9079) );
  NOR2_X1 U10404 ( .A1(n9362), .A2(n9191), .ZN(n9078) );
  AOI211_X1 U10405 ( .C1(n9195), .C2(n9080), .A(n9079), .B(n9078), .ZN(n9084)
         );
  NAND3_X1 U10406 ( .A1(n9082), .A2(n9184), .A3(n9081), .ZN(n9083) );
  NAND4_X1 U10407 ( .A1(n9086), .A2(n9085), .A3(n9084), .A4(n9083), .ZN(
        P1_U3220) );
  OAI21_X1 U10408 ( .B1(n9089), .B2(n9088), .A(n9087), .ZN(n9090) );
  NAND2_X1 U10409 ( .A1(n9090), .A2(n9184), .ZN(n9096) );
  AOI22_X1 U10410 ( .A1(n9091), .A2(n9195), .B1(P1_REG3_REG_8__SCAN_IN), .B2(
        P1_U3086), .ZN(n9095) );
  NAND2_X1 U10411 ( .A1(n9201), .A2(n9564), .ZN(n9094) );
  INV_X1 U10412 ( .A(n9560), .ZN(n9092) );
  NAND2_X1 U10413 ( .A1(n9145), .A2(n9092), .ZN(n9093) );
  NAND4_X1 U10414 ( .A1(n9096), .A2(n9095), .A3(n9094), .A4(n9093), .ZN(
        P1_U3221) );
  XOR2_X1 U10415 ( .A(n9098), .B(n9097), .Z(n9105) );
  NOR2_X1 U10416 ( .A1(n9198), .A2(n9487), .ZN(n9103) );
  NAND2_X1 U10417 ( .A1(n9214), .A2(n9173), .ZN(n9100) );
  NAND2_X1 U10418 ( .A1(n9212), .A2(n9150), .ZN(n9099) );
  AND2_X1 U10419 ( .A1(n9100), .A2(n9099), .ZN(n9481) );
  OAI22_X1 U10420 ( .A1(n9481), .A2(n9143), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9101), .ZN(n9102) );
  AOI211_X1 U10421 ( .C1(n9486), .C2(n9201), .A(n9103), .B(n9102), .ZN(n9104)
         );
  OAI21_X1 U10422 ( .B1(n9105), .B2(n9204), .A(n9104), .ZN(P1_U3223) );
  OAI21_X1 U10423 ( .B1(n9107), .B2(n9106), .A(n9179), .ZN(n9108) );
  NAND2_X1 U10424 ( .A1(n9108), .A2(n9184), .ZN(n9114) );
  AOI22_X1 U10425 ( .A1(n9209), .A2(n9150), .B1(n9173), .B2(n9211), .ZN(n9423)
         );
  INV_X1 U10426 ( .A(n9423), .ZN(n9112) );
  INV_X1 U10427 ( .A(n9428), .ZN(n9110) );
  OAI22_X1 U10428 ( .A1(n9110), .A2(n9198), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9109), .ZN(n9111) );
  AOI21_X1 U10429 ( .B1(n9112), .B2(n9195), .A(n9111), .ZN(n9113) );
  OAI211_X1 U10430 ( .C1(n9663), .C2(n9191), .A(n9114), .B(n9113), .ZN(
        P1_U3225) );
  XNOR2_X1 U10431 ( .A(n9116), .B(n9117), .ZN(n9194) );
  INV_X1 U10432 ( .A(n9115), .ZN(n9193) );
  NOR2_X1 U10433 ( .A1(n9194), .A2(n9193), .ZN(n9192) );
  AOI21_X1 U10434 ( .B1(n9117), .B2(n9116), .A(n9192), .ZN(n9121) );
  XNOR2_X1 U10435 ( .A(n9119), .B(n9118), .ZN(n9120) );
  XNOR2_X1 U10436 ( .A(n9121), .B(n9120), .ZN(n9128) );
  AOI22_X1 U10437 ( .A1(n9122), .A2(n9195), .B1(P1_REG3_REG_16__SCAN_IN), .B2(
        P1_U3086), .ZN(n9123) );
  OAI21_X1 U10438 ( .B1(n9124), .B2(n9198), .A(n9123), .ZN(n9125) );
  AOI21_X1 U10439 ( .B1(n9126), .B2(n9201), .A(n9125), .ZN(n9127) );
  OAI21_X1 U10440 ( .B1(n9128), .B2(n9204), .A(n9127), .ZN(P1_U3226) );
  XOR2_X1 U10441 ( .A(n9130), .B(n9129), .Z(n9136) );
  NAND2_X1 U10442 ( .A1(n9216), .A2(n9150), .ZN(n9131) );
  OAI21_X1 U10443 ( .B1(n9132), .B2(n9373), .A(n9131), .ZN(n9551) );
  NAND2_X1 U10444 ( .A1(n9551), .A2(n9195), .ZN(n9133) );
  NAND2_X1 U10445 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9301) );
  OAI211_X1 U10446 ( .C1(n9198), .C2(n9541), .A(n9133), .B(n9301), .ZN(n9134)
         );
  AOI21_X1 U10447 ( .B1(n9636), .B2(n9201), .A(n9134), .ZN(n9135) );
  OAI21_X1 U10448 ( .B1(n9136), .B2(n9204), .A(n9135), .ZN(P1_U3228) );
  OAI21_X1 U10449 ( .B1(n9139), .B2(n9138), .A(n9137), .ZN(n9140) );
  NAND2_X1 U10450 ( .A1(n9140), .A2(n9184), .ZN(n9147) );
  INV_X1 U10451 ( .A(n9186), .ZN(n9210) );
  NOR2_X1 U10452 ( .A1(n9161), .A2(n9373), .ZN(n9141) );
  AOI21_X1 U10453 ( .B1(n9210), .B2(n9150), .A(n9141), .ZN(n9440) );
  OAI22_X1 U10454 ( .A1(n9440), .A2(n9143), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9142), .ZN(n9144) );
  AOI21_X1 U10455 ( .B1(n9444), .B2(n9145), .A(n9144), .ZN(n9146) );
  OAI211_X1 U10456 ( .C1(n4703), .C2(n9191), .A(n9147), .B(n9146), .ZN(
        P1_U3229) );
  XOR2_X1 U10457 ( .A(n9149), .B(n9148), .Z(n9156) );
  OR2_X1 U10458 ( .A1(n9175), .A2(n9373), .ZN(n9152) );
  NAND2_X1 U10459 ( .A1(n9213), .A2(n9150), .ZN(n9151) );
  NAND2_X1 U10460 ( .A1(n9152), .A2(n9151), .ZN(n9498) );
  AOI22_X1 U10461 ( .A1(n9498), .A2(n9195), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n9153) );
  OAI21_X1 U10462 ( .B1(n9505), .B2(n9198), .A(n9153), .ZN(n9154) );
  AOI21_X1 U10463 ( .B1(n9504), .B2(n9201), .A(n9154), .ZN(n9155) );
  OAI21_X1 U10464 ( .B1(n9156), .B2(n9204), .A(n9155), .ZN(P1_U3233) );
  OAI21_X1 U10465 ( .B1(n9159), .B2(n9158), .A(n9157), .ZN(n9165) );
  NAND2_X1 U10466 ( .A1(n9474), .A2(n9201), .ZN(n9163) );
  OAI22_X1 U10467 ( .A1(n9161), .A2(n9350), .B1(n9160), .B2(n9373), .ZN(n9466)
         );
  AOI22_X1 U10468 ( .A1(n9466), .A2(n9195), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n9162) );
  OAI211_X1 U10469 ( .C1(n9198), .C2(n9471), .A(n9163), .B(n9162), .ZN(n9164)
         );
  AOI21_X1 U10470 ( .B1(n9165), .B2(n9184), .A(n9164), .ZN(n9166) );
  INV_X1 U10471 ( .A(n9166), .ZN(P1_U3235) );
  AND2_X1 U10472 ( .A1(n9168), .A2(n9167), .ZN(n9170) );
  NAND2_X1 U10473 ( .A1(n9170), .A2(n9171), .ZN(n9169) );
  OAI21_X1 U10474 ( .B1(n9171), .B2(n9170), .A(n9169), .ZN(n9172) );
  NAND2_X1 U10475 ( .A1(n9172), .A2(n9184), .ZN(n9178) );
  NAND2_X1 U10476 ( .A1(n9217), .A2(n9173), .ZN(n9174) );
  OAI21_X1 U10477 ( .B1(n9175), .B2(n9350), .A(n9174), .ZN(n9534) );
  AND2_X1 U10478 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9316) );
  NOR2_X1 U10479 ( .A1(n9198), .A2(n9526), .ZN(n9176) );
  AOI211_X1 U10480 ( .C1(n9195), .C2(n9534), .A(n9316), .B(n9176), .ZN(n9177)
         );
  OAI211_X1 U10481 ( .C1(n9951), .C2(n9191), .A(n9178), .B(n9177), .ZN(
        P1_U3238) );
  INV_X1 U10482 ( .A(n9179), .ZN(n9182) );
  OAI21_X1 U10483 ( .B1(n9182), .B2(n9181), .A(n9180), .ZN(n9185) );
  NAND3_X1 U10484 ( .A1(n9185), .A2(n9184), .A3(n9183), .ZN(n9190) );
  OAI22_X1 U10485 ( .A1(n9187), .A2(n9350), .B1(n9186), .B2(n9373), .ZN(n9411)
         );
  OAI22_X1 U10486 ( .A1(n9405), .A2(n9198), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9775), .ZN(n9188) );
  AOI21_X1 U10487 ( .B1(n9411), .B2(n9195), .A(n9188), .ZN(n9189) );
  OAI211_X1 U10488 ( .C1(n9408), .C2(n9191), .A(n9190), .B(n9189), .ZN(
        P1_U3240) );
  AOI21_X1 U10489 ( .B1(n9194), .B2(n9193), .A(n9192), .ZN(n9205) );
  AOI22_X1 U10490 ( .A1(n9196), .A2(n9195), .B1(P1_REG3_REG_15__SCAN_IN), .B2(
        P1_U3086), .ZN(n9197) );
  OAI21_X1 U10491 ( .B1(n9199), .B2(n9198), .A(n9197), .ZN(n9200) );
  AOI21_X1 U10492 ( .B1(n9202), .B2(n9201), .A(n9200), .ZN(n9203) );
  OAI21_X1 U10493 ( .B1(n9205), .B2(n9204), .A(n9203), .ZN(P1_U3241) );
  MUX2_X1 U10494 ( .A(n9353), .B(P1_DATAO_REG_31__SCAN_IN), .S(n9231), .Z(
        P1_U3585) );
  MUX2_X1 U10495 ( .A(n9206), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9231), .Z(
        P1_U3584) );
  MUX2_X1 U10496 ( .A(n9207), .B(P1_DATAO_REG_29__SCAN_IN), .S(n9231), .Z(
        P1_U3583) );
  MUX2_X1 U10497 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9208), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10498 ( .A(n9209), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9231), .Z(
        P1_U3580) );
  MUX2_X1 U10499 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9210), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10500 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9211), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10501 ( .A(n9212), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9231), .Z(
        P1_U3576) );
  MUX2_X1 U10502 ( .A(n9213), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9231), .Z(
        P1_U3575) );
  MUX2_X1 U10503 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9214), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10504 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9215), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10505 ( .A(n9216), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9231), .Z(
        P1_U3572) );
  MUX2_X1 U10506 ( .A(n9217), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9231), .Z(
        P1_U3571) );
  MUX2_X1 U10507 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9218), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10508 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n4655), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10509 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9219), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10510 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9220), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10511 ( .A(n9221), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9231), .Z(
        P1_U3565) );
  MUX2_X1 U10512 ( .A(n9222), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9231), .Z(
        P1_U3564) );
  MUX2_X1 U10513 ( .A(n9223), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9231), .Z(
        P1_U3563) );
  MUX2_X1 U10514 ( .A(n9224), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9231), .Z(
        P1_U3562) );
  MUX2_X1 U10515 ( .A(n9225), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9231), .Z(
        P1_U3561) );
  MUX2_X1 U10516 ( .A(n9226), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9231), .Z(
        P1_U3560) );
  MUX2_X1 U10517 ( .A(n9227), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9231), .Z(
        P1_U3559) );
  MUX2_X1 U10518 ( .A(n9228), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9231), .Z(
        P1_U3558) );
  MUX2_X1 U10519 ( .A(n9229), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9231), .Z(
        P1_U3557) );
  MUX2_X1 U10520 ( .A(n6805), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9231), .Z(
        P1_U3556) );
  MUX2_X1 U10521 ( .A(n9230), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9231), .Z(
        P1_U3555) );
  MUX2_X1 U10522 ( .A(n6109), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9231), .Z(
        P1_U3554) );
  AOI211_X1 U10523 ( .C1(n9243), .C2(n9233), .A(n9232), .B(n10044), .ZN(n9234)
         );
  INV_X1 U10524 ( .A(n9234), .ZN(n9242) );
  AOI22_X1 U10525 ( .A1(n10043), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9241) );
  NAND2_X1 U10526 ( .A1(n10052), .A2(n9235), .ZN(n9240) );
  OAI211_X1 U10527 ( .C1(n9238), .C2(n9237), .A(n10057), .B(n9236), .ZN(n9239)
         );
  NAND4_X1 U10528 ( .A1(n9242), .A2(n9241), .A3(n9240), .A4(n9239), .ZN(
        P1_U3244) );
  MUX2_X1 U10529 ( .A(n9244), .B(n9243), .S(n10031), .Z(n9247) );
  NOR2_X1 U10530 ( .A1(n6372), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9245) );
  OR2_X1 U10531 ( .A1(n9245), .A2(n9246), .ZN(n10032) );
  NAND2_X1 U10532 ( .A1(n10032), .A2(n10034), .ZN(n10037) );
  OAI211_X1 U10533 ( .C1(n9247), .C2(n9246), .A(P1_U3973), .B(n10037), .ZN(
        n10048) );
  AOI22_X1 U10534 ( .A1(P1_U3086), .A2(P1_REG3_REG_2__SCAN_IN), .B1(n10043), 
        .B2(P1_ADDR_REG_2__SCAN_IN), .ZN(n9259) );
  AOI211_X1 U10535 ( .C1(n9250), .C2(n9249), .A(n9248), .B(n10044), .ZN(n9257)
         );
  OAI21_X1 U10536 ( .B1(n9253), .B2(n9252), .A(n9251), .ZN(n9254) );
  OAI22_X1 U10537 ( .A1(n9255), .A2(n9335), .B1(n9336), .B2(n9254), .ZN(n9256)
         );
  NOR2_X1 U10538 ( .A1(n9257), .A2(n9256), .ZN(n9258) );
  NAND3_X1 U10539 ( .A1(n10048), .A2(n9259), .A3(n9258), .ZN(P1_U3245) );
  NOR2_X1 U10540 ( .A1(n7629), .A2(n9262), .ZN(n9280) );
  AOI211_X1 U10541 ( .C1(n7629), .C2(n9262), .A(n9280), .B(n10044), .ZN(n9271)
         );
  OAI21_X1 U10542 ( .B1(n9264), .B2(n7266), .A(n9263), .ZN(n9272) );
  XNOR2_X1 U10543 ( .A(n9278), .B(n9272), .ZN(n9265) );
  NAND2_X1 U10544 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n9265), .ZN(n9274) );
  OAI211_X1 U10545 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n9265), .A(n10057), .B(
        n9274), .ZN(n9269) );
  NOR2_X1 U10546 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9266), .ZN(n9267) );
  AOI21_X1 U10547 ( .B1(n10043), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n9267), .ZN(
        n9268) );
  OAI211_X1 U10548 ( .C1(n9335), .C2(n9278), .A(n9269), .B(n9268), .ZN(n9270)
         );
  OR2_X1 U10549 ( .A1(n9271), .A2(n9270), .ZN(P1_U3258) );
  NAND2_X1 U10550 ( .A1(n9273), .A2(n9272), .ZN(n9275) );
  NAND2_X1 U10551 ( .A1(n9275), .A2(n9274), .ZN(n9277) );
  XNOR2_X1 U10552 ( .A(n9294), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n9276) );
  NOR2_X1 U10553 ( .A1(n9276), .A2(n9277), .ZN(n9296) );
  AOI21_X1 U10554 ( .B1(n9277), .B2(n9276), .A(n9296), .ZN(n9291) );
  NOR2_X1 U10555 ( .A1(n9279), .A2(n9278), .ZN(n9281) );
  NOR2_X1 U10556 ( .A1(n9281), .A2(n9280), .ZN(n9284) );
  NAND2_X1 U10557 ( .A1(n9294), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9282) );
  OAI21_X1 U10558 ( .B1(n9294), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9282), .ZN(
        n9283) );
  NOR2_X1 U10559 ( .A1(n9284), .A2(n9283), .ZN(n9293) );
  AOI211_X1 U10560 ( .C1(n9284), .C2(n9283), .A(n9293), .B(n10044), .ZN(n9285)
         );
  INV_X1 U10561 ( .A(n9285), .ZN(n9290) );
  NOR2_X1 U10562 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9286), .ZN(n9288) );
  NOR2_X1 U10563 ( .A1(n9335), .A2(n9297), .ZN(n9287) );
  AOI211_X1 U10564 ( .C1(n10043), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n9288), .B(
        n9287), .ZN(n9289) );
  OAI211_X1 U10565 ( .C1(n9291), .C2(n9336), .A(n9290), .B(n9289), .ZN(
        P1_U3259) );
  XNOR2_X1 U10566 ( .A(n9317), .B(n9292), .ZN(n9308) );
  AOI21_X1 U10567 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n9294), .A(n9293), .ZN(
        n9309) );
  XOR2_X1 U10568 ( .A(n9308), .B(n9309), .Z(n9307) );
  XNOR2_X1 U10569 ( .A(n9317), .B(n9295), .ZN(n9300) );
  AOI21_X1 U10570 ( .B1(n9297), .B2(n9845), .A(n9296), .ZN(n9298) );
  INV_X1 U10571 ( .A(n9298), .ZN(n9299) );
  NAND2_X1 U10572 ( .A1(n9300), .A2(n9299), .ZN(n9319) );
  OAI21_X1 U10573 ( .B1(n9300), .B2(n9299), .A(n9319), .ZN(n9305) );
  NAND2_X1 U10574 ( .A1(n10043), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n9302) );
  OAI211_X1 U10575 ( .C1(n9335), .C2(n9303), .A(n9302), .B(n9301), .ZN(n9304)
         );
  AOI21_X1 U10576 ( .B1(n10057), .B2(n9305), .A(n9304), .ZN(n9306) );
  OAI21_X1 U10577 ( .B1(n9307), .B2(n10044), .A(n9306), .ZN(P1_U3260) );
  INV_X1 U10578 ( .A(n9330), .ZN(n9325) );
  NAND2_X1 U10579 ( .A1(n9309), .A2(n9308), .ZN(n9311) );
  OR2_X1 U10580 ( .A1(n9317), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9310) );
  NAND2_X1 U10581 ( .A1(n9311), .A2(n9310), .ZN(n9314) );
  NAND2_X1 U10582 ( .A1(n9330), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9326) );
  OR2_X1 U10583 ( .A1(n9330), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9312) );
  NAND2_X1 U10584 ( .A1(n9326), .A2(n9312), .ZN(n9313) );
  NOR2_X1 U10585 ( .A1(n9314), .A2(n9313), .ZN(n9328) );
  AOI211_X1 U10586 ( .C1(n9314), .C2(n9313), .A(n9328), .B(n10044), .ZN(n9315)
         );
  AOI211_X1 U10587 ( .C1(n10043), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n9316), .B(
        n9315), .ZN(n9324) );
  OR2_X1 U10588 ( .A1(n9317), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9318) );
  NAND2_X1 U10589 ( .A1(n9319), .A2(n9318), .ZN(n9321) );
  XNOR2_X1 U10590 ( .A(n9330), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9320) );
  NAND2_X1 U10591 ( .A1(n9321), .A2(n9320), .ZN(n9322) );
  NAND3_X1 U10592 ( .A1(n10057), .A2(n9332), .A3(n9322), .ZN(n9323) );
  OAI211_X1 U10593 ( .C1(n9335), .C2(n9325), .A(n9324), .B(n9323), .ZN(
        P1_U3261) );
  INV_X1 U10594 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9348) );
  INV_X1 U10595 ( .A(n9326), .ZN(n9327) );
  OR2_X1 U10596 ( .A1(n9328), .A2(n9327), .ZN(n9329) );
  XNOR2_X1 U10597 ( .A(n9329), .B(n9520), .ZN(n9341) );
  INV_X1 U10598 ( .A(n9341), .ZN(n9338) );
  NAND2_X1 U10599 ( .A1(n9330), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9331) );
  NAND2_X1 U10600 ( .A1(n9332), .A2(n9331), .ZN(n9334) );
  XNOR2_X1 U10601 ( .A(n9334), .B(n9333), .ZN(n9339) );
  OAI21_X1 U10602 ( .B1(n9336), .B2(n9339), .A(n9335), .ZN(n9337) );
  AOI21_X1 U10603 ( .B1(n9338), .B2(n9340), .A(n9337), .ZN(n9344) );
  AOI22_X1 U10604 ( .A1(n9341), .A2(n9340), .B1(n10057), .B2(n9339), .ZN(n9343) );
  MUX2_X1 U10605 ( .A(n9344), .B(n9343), .S(n9342), .Z(n9346) );
  OAI211_X1 U10606 ( .C1(n9348), .C2(n9347), .A(n9346), .B(n9345), .ZN(
        P1_U3262) );
  NAND2_X1 U10607 ( .A1(n9349), .A2(n10094), .ZN(n9571) );
  AND2_X1 U10608 ( .A1(n10031), .A2(P1_B_REG_SCAN_IN), .ZN(n9351) );
  OR2_X1 U10609 ( .A1(n9351), .A2(n9350), .ZN(n9375) );
  INV_X1 U10610 ( .A(n9375), .ZN(n9352) );
  NAND2_X1 U10611 ( .A1(n9353), .A2(n9352), .ZN(n9574) );
  NOR2_X1 U10612 ( .A1(n9574), .A2(n10102), .ZN(n9358) );
  NOR2_X1 U10613 ( .A1(n9649), .A2(n10096), .ZN(n9354) );
  AOI211_X1 U10614 ( .C1(n10102), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9358), .B(
        n9354), .ZN(n9355) );
  OAI21_X1 U10615 ( .B1(n10097), .B2(n9571), .A(n9355), .ZN(P1_U3263) );
  OAI211_X1 U10616 ( .C1(n9653), .C2(n9376), .A(n10094), .B(n9356), .ZN(n9575)
         );
  NOR2_X1 U10617 ( .A1(n9562), .A2(n9357), .ZN(n9359) );
  AOI211_X1 U10618 ( .C1(n9360), .C2(n10074), .A(n9359), .B(n9358), .ZN(n9361)
         );
  OAI21_X1 U10619 ( .B1(n9575), .B2(n10097), .A(n9361), .ZN(P1_U3264) );
  NAND2_X1 U10620 ( .A1(n9071), .A2(n9363), .ZN(n9364) );
  NAND2_X1 U10621 ( .A1(n9365), .A2(n9364), .ZN(n9366) );
  XNOR2_X1 U10622 ( .A(n9366), .B(n9370), .ZN(n9578) );
  INV_X1 U10623 ( .A(n9578), .ZN(n9386) );
  INV_X1 U10624 ( .A(n9370), .ZN(n9371) );
  AOI211_X1 U10625 ( .C1(n9581), .C2(n9377), .A(n9540), .B(n9376), .ZN(n9580)
         );
  NAND2_X1 U10626 ( .A1(n9580), .A2(n10081), .ZN(n9382) );
  NOR3_X1 U10627 ( .A1(n9379), .A2(n9378), .A3(n9559), .ZN(n9380) );
  AOI21_X1 U10628 ( .B1(n10102), .B2(P1_REG2_REG_29__SCAN_IN), .A(n9380), .ZN(
        n9381) );
  OAI211_X1 U10629 ( .C1(n9383), .C2(n10096), .A(n9382), .B(n9381), .ZN(n9384)
         );
  AOI21_X1 U10630 ( .B1(n9579), .B2(n9562), .A(n9384), .ZN(n9385) );
  OAI21_X1 U10631 ( .B1(n9386), .B2(n9557), .A(n9385), .ZN(P1_U3356) );
  XNOR2_X1 U10632 ( .A(n9387), .B(n9394), .ZN(n9586) );
  INV_X1 U10633 ( .A(n9586), .ZN(n9401) );
  AOI211_X1 U10634 ( .C1(n9389), .C2(n9403), .A(n9540), .B(n9388), .ZN(n9585)
         );
  NOR2_X1 U10635 ( .A1(n9658), .A2(n10096), .ZN(n9393) );
  OAI22_X1 U10636 ( .A1(n9391), .A2(n9559), .B1(n9390), .B2(n9562), .ZN(n9392)
         );
  AOI211_X1 U10637 ( .C1(n9585), .C2(n10081), .A(n9393), .B(n9392), .ZN(n9400)
         );
  XNOR2_X1 U10638 ( .A(n9395), .B(n9394), .ZN(n9396) );
  NAND2_X1 U10639 ( .A1(n9396), .A2(n10072), .ZN(n9398) );
  NAND2_X1 U10640 ( .A1(n9398), .A2(n9397), .ZN(n9584) );
  NAND2_X1 U10641 ( .A1(n9584), .A2(n9562), .ZN(n9399) );
  OAI211_X1 U10642 ( .C1(n9401), .C2(n9557), .A(n9400), .B(n9399), .ZN(
        P1_U3266) );
  XNOR2_X1 U10643 ( .A(n9402), .B(n9409), .ZN(n9593) );
  INV_X1 U10644 ( .A(n9425), .ZN(n9404) );
  AOI211_X1 U10645 ( .C1(n9590), .C2(n9404), .A(n9540), .B(n4699), .ZN(n9589)
         );
  INV_X1 U10646 ( .A(n9405), .ZN(n9406) );
  AOI22_X1 U10647 ( .A1(n9406), .A2(n10091), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n10102), .ZN(n9407) );
  OAI21_X1 U10648 ( .B1(n9408), .B2(n10096), .A(n9407), .ZN(n9414) );
  XNOR2_X1 U10649 ( .A(n9410), .B(n9409), .ZN(n9412) );
  AOI21_X1 U10650 ( .B1(n9412), .B2(n10072), .A(n9411), .ZN(n9592) );
  NOR2_X1 U10651 ( .A1(n9592), .A2(n10102), .ZN(n9413) );
  AOI211_X1 U10652 ( .C1(n9589), .C2(n10081), .A(n9414), .B(n9413), .ZN(n9415)
         );
  OAI21_X1 U10653 ( .B1(n9593), .B2(n9557), .A(n9415), .ZN(P1_U3267) );
  XOR2_X1 U10654 ( .A(n9418), .B(n9416), .Z(n9596) );
  INV_X1 U10655 ( .A(n9596), .ZN(n9433) );
  NAND2_X1 U10656 ( .A1(n9438), .A2(n9417), .ZN(n9419) );
  NAND2_X1 U10657 ( .A1(n9419), .A2(n9418), .ZN(n9421) );
  NAND2_X1 U10658 ( .A1(n9421), .A2(n9420), .ZN(n9422) );
  NAND2_X1 U10659 ( .A1(n9422), .A2(n10072), .ZN(n9424) );
  NAND2_X1 U10660 ( .A1(n9424), .A2(n9423), .ZN(n9594) );
  INV_X1 U10661 ( .A(n9442), .ZN(n9426) );
  AOI211_X1 U10662 ( .C1(n9427), .C2(n9426), .A(n9540), .B(n9425), .ZN(n9595)
         );
  NAND2_X1 U10663 ( .A1(n9595), .A2(n10081), .ZN(n9430) );
  AOI22_X1 U10664 ( .A1(n9428), .A2(n10091), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n10102), .ZN(n9429) );
  OAI211_X1 U10665 ( .C1(n9663), .C2(n10096), .A(n9430), .B(n9429), .ZN(n9431)
         );
  AOI21_X1 U10666 ( .B1(n9594), .B2(n9562), .A(n9431), .ZN(n9432) );
  OAI21_X1 U10667 ( .B1(n9433), .B2(n9557), .A(n9432), .ZN(P1_U3268) );
  XNOR2_X1 U10668 ( .A(n9434), .B(n9436), .ZN(n9601) );
  INV_X1 U10669 ( .A(n9601), .ZN(n9449) );
  NAND2_X1 U10670 ( .A1(n9457), .A2(n9435), .ZN(n9437) );
  NAND2_X1 U10671 ( .A1(n9437), .A2(n9436), .ZN(n9439) );
  NAND3_X1 U10672 ( .A1(n9439), .A2(n10072), .A3(n9438), .ZN(n9441) );
  NAND2_X1 U10673 ( .A1(n9441), .A2(n9440), .ZN(n9599) );
  AOI211_X1 U10674 ( .C1(n9443), .C2(n9452), .A(n9540), .B(n9442), .ZN(n9600)
         );
  NAND2_X1 U10675 ( .A1(n9600), .A2(n10081), .ZN(n9446) );
  AOI22_X1 U10676 ( .A1(n9444), .A2(n10091), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n10102), .ZN(n9445) );
  OAI211_X1 U10677 ( .C1(n4703), .C2(n10096), .A(n9446), .B(n9445), .ZN(n9447)
         );
  AOI21_X1 U10678 ( .B1(n9599), .B2(n9562), .A(n9447), .ZN(n9448) );
  OAI21_X1 U10679 ( .B1(n9449), .B2(n9557), .A(n9448), .ZN(P1_U3269) );
  XNOR2_X1 U10680 ( .A(n9450), .B(n4491), .ZN(n9607) );
  INV_X1 U10681 ( .A(n9452), .ZN(n9453) );
  AOI211_X1 U10682 ( .C1(n6126), .C2(n9451), .A(n9540), .B(n9453), .ZN(n9604)
         );
  AOI22_X1 U10683 ( .A1(n9454), .A2(n10091), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n10102), .ZN(n9455) );
  OAI21_X1 U10684 ( .B1(n9456), .B2(n10096), .A(n9455), .ZN(n9463) );
  OAI21_X1 U10685 ( .B1(n9459), .B2(n9458), .A(n9457), .ZN(n9461) );
  AOI21_X1 U10686 ( .B1(n9461), .B2(n10072), .A(n9460), .ZN(n9606) );
  NOR2_X1 U10687 ( .A1(n9606), .A2(n10102), .ZN(n9462) );
  AOI211_X1 U10688 ( .C1(n9604), .C2(n10081), .A(n9463), .B(n9462), .ZN(n9464)
         );
  OAI21_X1 U10689 ( .B1(n9607), .B2(n9557), .A(n9464), .ZN(P1_U3270) );
  XNOR2_X1 U10690 ( .A(n9465), .B(n9469), .ZN(n9467) );
  AOI21_X1 U10691 ( .B1(n9467), .B2(n10072), .A(n9466), .ZN(n9609) );
  XOR2_X1 U10692 ( .A(n9468), .B(n9469), .Z(n9612) );
  NAND2_X1 U10693 ( .A1(n9612), .A2(n10082), .ZN(n9476) );
  INV_X1 U10694 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9470) );
  OAI22_X1 U10695 ( .A1(n9471), .A2(n9559), .B1(n9562), .B2(n9470), .ZN(n9473)
         );
  OAI211_X1 U10696 ( .C1(n9485), .C2(n9610), .A(n10094), .B(n9451), .ZN(n9608)
         );
  NOR2_X1 U10697 ( .A1(n9608), .A2(n10097), .ZN(n9472) );
  AOI211_X1 U10698 ( .C1(n10074), .C2(n9474), .A(n9473), .B(n9472), .ZN(n9475)
         );
  OAI211_X1 U10699 ( .C1(n10102), .C2(n9609), .A(n9476), .B(n9475), .ZN(
        P1_U3271) );
  NAND2_X1 U10700 ( .A1(n9477), .A2(n9483), .ZN(n9478) );
  NAND2_X1 U10701 ( .A1(n9479), .A2(n9478), .ZN(n9480) );
  NAND2_X1 U10702 ( .A1(n9480), .A2(n10072), .ZN(n9482) );
  NAND2_X1 U10703 ( .A1(n9482), .A2(n9481), .ZN(n9614) );
  INV_X1 U10704 ( .A(n9614), .ZN(n9493) );
  XNOR2_X1 U10705 ( .A(n9484), .B(n9483), .ZN(n9616) );
  NAND2_X1 U10706 ( .A1(n9616), .A2(n10082), .ZN(n9492) );
  AOI211_X1 U10707 ( .C1(n9486), .C2(n4698), .A(n9540), .B(n9485), .ZN(n9615)
         );
  NOR2_X1 U10708 ( .A1(n9942), .A2(n10096), .ZN(n9490) );
  OAI22_X1 U10709 ( .A1(n9562), .A2(n9488), .B1(n9487), .B2(n9559), .ZN(n9489)
         );
  AOI211_X1 U10710 ( .C1(n9615), .C2(n10081), .A(n9490), .B(n9489), .ZN(n9491)
         );
  OAI211_X1 U10711 ( .C1(n10102), .C2(n9493), .A(n9492), .B(n9491), .ZN(
        P1_U3272) );
  AOI21_X1 U10712 ( .B1(n9495), .B2(n9501), .A(n10087), .ZN(n9496) );
  OAI21_X1 U10713 ( .B1(n9497), .B2(n4817), .A(n9496), .ZN(n9500) );
  INV_X1 U10714 ( .A(n9498), .ZN(n9499) );
  NAND2_X1 U10715 ( .A1(n9500), .A2(n9499), .ZN(n9618) );
  INV_X1 U10716 ( .A(n9618), .ZN(n9511) );
  XOR2_X1 U10717 ( .A(n9502), .B(n9501), .Z(n9620) );
  NAND2_X1 U10718 ( .A1(n9620), .A2(n10082), .ZN(n9510) );
  AOI211_X1 U10719 ( .C1(n9504), .C2(n4975), .A(n9540), .B(n9503), .ZN(n9619)
         );
  NOR2_X1 U10720 ( .A1(n9946), .A2(n10096), .ZN(n9508) );
  OAI22_X1 U10721 ( .A1(n9562), .A2(n9506), .B1(n9505), .B2(n9559), .ZN(n9507)
         );
  AOI211_X1 U10722 ( .C1(n9619), .C2(n10081), .A(n9508), .B(n9507), .ZN(n9509)
         );
  OAI211_X1 U10723 ( .C1(n10102), .C2(n9511), .A(n9510), .B(n9509), .ZN(
        P1_U3273) );
  XNOR2_X1 U10724 ( .A(n9513), .B(n9512), .ZN(n9515) );
  AOI21_X1 U10725 ( .B1(n9515), .B2(n10072), .A(n9514), .ZN(n9627) );
  OR2_X1 U10726 ( .A1(n4476), .A2(n9516), .ZN(n9623) );
  NAND3_X1 U10727 ( .A1(n9623), .A2(n9622), .A3(n10082), .ZN(n9524) );
  INV_X1 U10728 ( .A(n4975), .ZN(n9517) );
  AOI211_X1 U10729 ( .C1(n9625), .C2(n9528), .A(n9540), .B(n9517), .ZN(n9624)
         );
  NOR2_X1 U10730 ( .A1(n9518), .A2(n10096), .ZN(n9522) );
  OAI22_X1 U10731 ( .A1(n9562), .A2(n9520), .B1(n9519), .B2(n9559), .ZN(n9521)
         );
  AOI211_X1 U10732 ( .C1(n9624), .C2(n10081), .A(n9522), .B(n9521), .ZN(n9523)
         );
  OAI211_X1 U10733 ( .C1(n10102), .C2(n9627), .A(n9524), .B(n9523), .ZN(
        P1_U3274) );
  XNOR2_X1 U10734 ( .A(n9525), .B(n4502), .ZN(n9631) );
  OAI22_X1 U10735 ( .A1(n9562), .A2(n9527), .B1(n9526), .B2(n9559), .ZN(n9530)
         );
  OAI211_X1 U10736 ( .C1(n9539), .C2(n9951), .A(n9528), .B(n10094), .ZN(n9629)
         );
  NOR2_X1 U10737 ( .A1(n9629), .A2(n10097), .ZN(n9529) );
  AOI211_X1 U10738 ( .C1(n10074), .C2(n9531), .A(n9530), .B(n9529), .ZN(n9537)
         );
  XNOR2_X1 U10739 ( .A(n9533), .B(n9532), .ZN(n9535) );
  AOI21_X1 U10740 ( .B1(n9535), .B2(n10072), .A(n9534), .ZN(n9630) );
  OR2_X1 U10741 ( .A1(n9630), .A2(n10102), .ZN(n9536) );
  OAI211_X1 U10742 ( .C1(n9631), .C2(n9557), .A(n9537), .B(n9536), .ZN(
        P1_U3275) );
  XNOR2_X1 U10743 ( .A(n9538), .B(n9549), .ZN(n9640) );
  AOI211_X1 U10744 ( .C1(n9636), .C2(n4978), .A(n9540), .B(n9539), .ZN(n9635)
         );
  INV_X1 U10745 ( .A(n9541), .ZN(n9542) );
  AOI22_X1 U10746 ( .A1(n10102), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9542), 
        .B2(n10091), .ZN(n9543) );
  OAI21_X1 U10747 ( .B1(n9544), .B2(n10096), .A(n9543), .ZN(n9555) );
  INV_X1 U10748 ( .A(n9545), .ZN(n9546) );
  AOI21_X1 U10749 ( .B1(n9548), .B2(n9546), .A(n10087), .ZN(n9553) );
  INV_X1 U10750 ( .A(n9547), .ZN(n9550) );
  OAI21_X1 U10751 ( .B1(n9550), .B2(n9549), .A(n9548), .ZN(n9552) );
  AOI21_X1 U10752 ( .B1(n9553), .B2(n9552), .A(n9551), .ZN(n9638) );
  NOR2_X1 U10753 ( .A1(n9638), .A2(n10102), .ZN(n9554) );
  AOI211_X1 U10754 ( .C1(n9635), .C2(n10081), .A(n9555), .B(n9554), .ZN(n9556)
         );
  OAI21_X1 U10755 ( .B1(n9640), .B2(n9557), .A(n9556), .ZN(P1_U3276) );
  NAND2_X1 U10756 ( .A1(n9558), .A2(n9562), .ZN(n9570) );
  OAI22_X1 U10757 ( .A1(n9562), .A2(n9561), .B1(n9560), .B2(n9559), .ZN(n9563)
         );
  AOI21_X1 U10758 ( .B1(n10074), .B2(n9564), .A(n9563), .ZN(n9569) );
  NAND2_X1 U10759 ( .A1(n9565), .A2(n10082), .ZN(n9568) );
  NAND2_X1 U10760 ( .A1(n9566), .A2(n10081), .ZN(n9567) );
  NAND4_X1 U10761 ( .A1(n9570), .A2(n9569), .A3(n9568), .A4(n9567), .ZN(
        P1_U3285) );
  OAI21_X1 U10762 ( .B1(n9649), .B2(n9646), .A(n9573), .ZN(P1_U3553) );
  AND2_X1 U10763 ( .A1(n9575), .A2(n9574), .ZN(n9650) );
  MUX2_X1 U10764 ( .A(n9576), .B(n9650), .S(n10186), .Z(n9577) );
  OAI21_X1 U10765 ( .B1(n9653), .B2(n9646), .A(n9577), .ZN(P1_U3552) );
  NAND2_X1 U10766 ( .A1(n9578), .A2(n10161), .ZN(n9583) );
  NAND2_X1 U10767 ( .A1(n9583), .A2(n9582), .ZN(n9654) );
  MUX2_X1 U10768 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9654), .S(n10186), .Z(
        P1_U3551) );
  AOI211_X1 U10769 ( .C1(n9586), .C2(n10161), .A(n9585), .B(n9584), .ZN(n9655)
         );
  MUX2_X1 U10770 ( .A(n9587), .B(n9655), .S(n10186), .Z(n9588) );
  OAI21_X1 U10771 ( .B1(n9658), .B2(n9646), .A(n9588), .ZN(P1_U3549) );
  AOI21_X1 U10772 ( .B1(n10165), .B2(n9590), .A(n9589), .ZN(n9591) );
  OAI211_X1 U10773 ( .C1(n9593), .C2(n9639), .A(n9592), .B(n9591), .ZN(n9659)
         );
  MUX2_X1 U10774 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9659), .S(n10186), .Z(
        P1_U3548) );
  AOI211_X1 U10775 ( .C1(n9596), .C2(n10161), .A(n9595), .B(n9594), .ZN(n9660)
         );
  MUX2_X1 U10776 ( .A(n9597), .B(n9660), .S(n10186), .Z(n9598) );
  OAI21_X1 U10777 ( .B1(n9663), .B2(n9646), .A(n9598), .ZN(P1_U3547) );
  AOI211_X1 U10778 ( .C1(n9601), .C2(n10161), .A(n9600), .B(n9599), .ZN(n9664)
         );
  MUX2_X1 U10779 ( .A(n9602), .B(n9664), .S(n10186), .Z(n9603) );
  OAI21_X1 U10780 ( .B1(n4703), .B2(n9646), .A(n9603), .ZN(P1_U3546) );
  AOI21_X1 U10781 ( .B1(n10165), .B2(n6126), .A(n9604), .ZN(n9605) );
  OAI211_X1 U10782 ( .C1(n9607), .C2(n9639), .A(n9606), .B(n9605), .ZN(n9667)
         );
  MUX2_X1 U10783 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9667), .S(n10186), .Z(
        P1_U3545) );
  INV_X1 U10784 ( .A(n10165), .ZN(n10159) );
  OAI211_X1 U10785 ( .C1(n9610), .C2(n10159), .A(n9609), .B(n9608), .ZN(n9611)
         );
  AOI21_X1 U10786 ( .B1(n9612), .B2(n10161), .A(n9611), .ZN(n9669) );
  NAND2_X1 U10787 ( .A1(n10184), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n9613) );
  OAI21_X1 U10788 ( .B1(n9669), .B2(n10184), .A(n9613), .ZN(P1_U3544) );
  AOI211_X1 U10789 ( .C1(n9616), .C2(n10161), .A(n9615), .B(n9614), .ZN(n9939)
         );
  MUX2_X1 U10790 ( .A(n9786), .B(n9939), .S(n10186), .Z(n9617) );
  OAI21_X1 U10791 ( .B1(n9942), .B2(n9646), .A(n9617), .ZN(P1_U3543) );
  AOI211_X1 U10792 ( .C1(n9620), .C2(n10161), .A(n9619), .B(n9618), .ZN(n9943)
         );
  MUX2_X1 U10793 ( .A(n9840), .B(n9943), .S(n10186), .Z(n9621) );
  OAI21_X1 U10794 ( .B1(n9946), .B2(n9646), .A(n9621), .ZN(P1_U3542) );
  NAND3_X1 U10795 ( .A1(n9623), .A2(n9622), .A3(n10161), .ZN(n9628) );
  AOI21_X1 U10796 ( .B1(n10165), .B2(n9625), .A(n9624), .ZN(n9626) );
  NAND3_X1 U10797 ( .A1(n9628), .A2(n9627), .A3(n9626), .ZN(n9947) );
  MUX2_X1 U10798 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9947), .S(n10186), .Z(
        P1_U3541) );
  OAI211_X1 U10799 ( .C1(n9631), .C2(n9639), .A(n9630), .B(n9629), .ZN(n9632)
         );
  INV_X1 U10800 ( .A(n9632), .ZN(n9948) );
  MUX2_X1 U10801 ( .A(n9633), .B(n9948), .S(n10186), .Z(n9634) );
  OAI21_X1 U10802 ( .B1(n9951), .B2(n9646), .A(n9634), .ZN(P1_U3540) );
  AOI21_X1 U10803 ( .B1(n10165), .B2(n9636), .A(n9635), .ZN(n9637) );
  OAI211_X1 U10804 ( .C1(n9640), .C2(n9639), .A(n9638), .B(n9637), .ZN(n9952)
         );
  MUX2_X1 U10805 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9952), .S(n10186), .Z(
        P1_U3539) );
  NAND2_X1 U10806 ( .A1(n9642), .A2(n9641), .ZN(n9643) );
  AOI21_X1 U10807 ( .B1(n9644), .B2(n10161), .A(n9643), .ZN(n9953) );
  MUX2_X1 U10808 ( .A(n9845), .B(n9953), .S(n10186), .Z(n9645) );
  OAI21_X1 U10809 ( .B1(n9957), .B2(n9646), .A(n9645), .ZN(P1_U3538) );
  OAI21_X1 U10810 ( .B1(n9649), .B2(n9956), .A(n9648), .ZN(P1_U3521) );
  MUX2_X1 U10811 ( .A(n9651), .B(n9650), .S(n10174), .Z(n9652) );
  OAI21_X1 U10812 ( .B1(n9653), .B2(n9956), .A(n9652), .ZN(P1_U3520) );
  MUX2_X1 U10813 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9654), .S(n10174), .Z(
        P1_U3519) );
  MUX2_X1 U10814 ( .A(n9656), .B(n9655), .S(n10174), .Z(n9657) );
  OAI21_X1 U10815 ( .B1(n9658), .B2(n9956), .A(n9657), .ZN(P1_U3517) );
  MUX2_X1 U10816 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9659), .S(n10174), .Z(
        P1_U3516) );
  MUX2_X1 U10817 ( .A(n9661), .B(n9660), .S(n10174), .Z(n9662) );
  OAI21_X1 U10818 ( .B1(n9663), .B2(n9956), .A(n9662), .ZN(P1_U3515) );
  MUX2_X1 U10819 ( .A(n9665), .B(n9664), .S(n10174), .Z(n9666) );
  OAI21_X1 U10820 ( .B1(n4703), .B2(n9956), .A(n9666), .ZN(P1_U3514) );
  MUX2_X1 U10821 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9667), .S(n10174), .Z(
        P1_U3513) );
  NOR2_X1 U10822 ( .A1(n10174), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n9668) );
  AOI21_X1 U10823 ( .B1(n9669), .B2(n10174), .A(n9668), .ZN(n9938) );
  NAND4_X1 U10824 ( .A1(P1_REG0_REG_16__SCAN_IN), .A2(P1_REG2_REG_15__SCAN_IN), 
        .A3(n9845), .A4(n7266), .ZN(n9670) );
  NOR3_X1 U10825 ( .A1(P1_REG1_REG_21__SCAN_IN), .A2(P1_REG0_REG_20__SCAN_IN), 
        .A3(n9670), .ZN(n9681) );
  INV_X1 U10826 ( .A(SI_12_), .ZN(n9892) );
  NOR4_X1 U10827 ( .A1(n9892), .A2(n9893), .A3(n9733), .A4(SI_0_), .ZN(n9671)
         );
  NAND3_X1 U10828 ( .A1(n9671), .A2(P2_DATAO_REG_5__SCAN_IN), .A3(
        P2_DATAO_REG_4__SCAN_IN), .ZN(n9679) );
  NOR4_X1 U10829 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_REG0_REG_21__SCAN_IN), 
        .A3(n6876), .A4(n9763), .ZN(n9677) );
  NOR4_X1 U10830 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(SI_17_), .A3(
        P2_DATAO_REG_15__SCAN_IN), .A4(n9874), .ZN(n9673) );
  NOR4_X1 U10831 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(SI_20_), .A3(n9776), 
        .A4(n9924), .ZN(n9672) );
  AND4_X1 U10832 ( .A1(n9674), .A2(P1_REG3_REG_4__SCAN_IN), .A3(n9673), .A4(
        n9672), .ZN(n9676) );
  INV_X1 U10833 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9675) );
  NAND4_X1 U10834 ( .A1(n9677), .A2(P1_IR_REG_30__SCAN_IN), .A3(n9676), .A4(
        n9675), .ZN(n9678) );
  NOR4_X1 U10835 ( .A1(n9869), .A2(n9798), .A3(n9679), .A4(n9678), .ZN(n9680)
         );
  NAND4_X1 U10836 ( .A1(P1_REG1_REG_20__SCAN_IN), .A2(P1_REG0_REG_17__SCAN_IN), 
        .A3(n9681), .A4(n9680), .ZN(n9718) );
  NOR2_X1 U10837 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .ZN(
        n9687) );
  NOR2_X1 U10838 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n9973) );
  INV_X1 U10839 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9912) );
  NAND4_X1 U10840 ( .A1(P1_STATE_REG_SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(n9912), .ZN(n9685) );
  NAND4_X1 U10841 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .A3(P1_IR_REG_20__SCAN_IN), .A4(n9750), .ZN(n9684) );
  NAND4_X1 U10842 ( .A1(P2_RD_REG_SCAN_IN), .A2(P1_D_REG_28__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(n9781), .ZN(n9683) );
  NAND4_X1 U10843 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n9682) );
  NOR4_X1 U10844 ( .A1(n9685), .A2(n9684), .A3(n9683), .A4(n9682), .ZN(n9686)
         );
  NAND4_X1 U10845 ( .A1(n9688), .A2(n9687), .A3(n9973), .A4(n9686), .ZN(n9717)
         );
  NAND4_X1 U10846 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(P1_REG1_REG_10__SCAN_IN), 
        .A3(P1_REG0_REG_9__SCAN_IN), .A4(n5843), .ZN(n9689) );
  NOR3_X1 U10847 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(P1_REG1_REG_12__SCAN_IN), 
        .A3(n9689), .ZN(n9695) );
  NAND4_X1 U10848 ( .A1(P1_REG0_REG_28__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .A3(n10297), .A4(n5293), .ZN(n9693) );
  NAND4_X1 U10849 ( .A1(P1_REG2_REG_2__SCAN_IN), .A2(P2_REG2_REG_23__SCAN_IN), 
        .A3(n10175), .A4(n5774), .ZN(n9691) );
  NAND4_X1 U10850 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(P2_STATE_REG_SCAN_IN), 
        .A3(P2_REG2_REG_31__SCAN_IN), .A4(n9755), .ZN(n9690) );
  OR4_X1 U10851 ( .A1(P1_REG2_REG_28__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), 
        .A3(n9691), .A4(n9690), .ZN(n9692) );
  NOR4_X1 U10852 ( .A1(n9693), .A2(n9752), .A3(n9753), .A4(n9692), .ZN(n9694)
         );
  NAND4_X1 U10853 ( .A1(P1_REG0_REG_13__SCAN_IN), .A2(n9695), .A3(n9694), .A4(
        n7493), .ZN(n9714) );
  NOR4_X1 U10854 ( .A1(P2_REG0_REG_18__SCAN_IN), .A2(P2_REG1_REG_19__SCAN_IN), 
        .A3(P1_REG2_REG_30__SCAN_IN), .A4(n9721), .ZN(n9699) );
  NOR4_X1 U10855 ( .A1(P2_REG1_REG_30__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), 
        .A3(n9897), .A4(n9900), .ZN(n9698) );
  NOR4_X1 U10856 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(n9871), .A3(n9764), .A4(
        n9926), .ZN(n9697) );
  NOR4_X1 U10857 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(P2_REG0_REG_3__SCAN_IN), 
        .A3(P1_REG2_REG_27__SCAN_IN), .A4(P2_ADDR_REG_17__SCAN_IN), .ZN(n9696)
         );
  NAND4_X1 U10858 ( .A1(n9699), .A2(n9698), .A3(n9697), .A4(n9696), .ZN(n9713)
         );
  INV_X1 U10859 ( .A(n9700), .ZN(n9712) );
  NAND4_X1 U10860 ( .A1(n9815), .A2(n9915), .A3(P2_IR_REG_27__SCAN_IN), .A4(
        P2_REG2_REG_27__SCAN_IN), .ZN(n9704) );
  INV_X1 U10861 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10259) );
  NOR2_X1 U10862 ( .A1(n10259), .A2(n6047), .ZN(n9702) );
  NOR4_X1 U10863 ( .A1(P2_REG1_REG_7__SCAN_IN), .A2(P2_REG2_REG_9__SCAN_IN), 
        .A3(P2_REG2_REG_20__SCAN_IN), .A4(n9783), .ZN(n9701) );
  NAND4_X1 U10864 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(n9702), .A3(n9701), .A4(
        P1_REG2_REG_29__SCAN_IN), .ZN(n9703) );
  NOR4_X1 U10865 ( .A1(n9704), .A2(n9703), .A3(P2_IR_REG_14__SCAN_IN), .A4(
        P2_IR_REG_9__SCAN_IN), .ZN(n9710) );
  AND4_X1 U10866 ( .A1(n9911), .A2(P2_REG1_REG_11__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .A4(P2_REG1_REG_0__SCAN_IN), .ZN(n9709) );
  NOR4_X1 U10867 ( .A1(n9705), .A2(P1_REG3_REG_26__SCAN_IN), .A3(
        P2_REG3_REG_2__SCAN_IN), .A4(P2_REG3_REG_0__SCAN_IN), .ZN(n9708) );
  INV_X1 U10868 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9706) );
  NOR4_X1 U10869 ( .A1(n9706), .A2(P1_IR_REG_24__SCAN_IN), .A3(
        P1_ADDR_REG_14__SCAN_IN), .A4(P2_D_REG_1__SCAN_IN), .ZN(n9707) );
  NAND4_X1 U10870 ( .A1(n9710), .A2(n9709), .A3(n9708), .A4(n9707), .ZN(n9711)
         );
  OR4_X1 U10871 ( .A1(n9714), .A2(n9713), .A3(n9712), .A4(n9711), .ZN(n9716)
         );
  INV_X1 U10872 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9974) );
  OR4_X1 U10873 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .A3(n9987), .A4(n9974), .ZN(n9715) );
  NOR4_X1 U10874 ( .A1(n9718), .A2(n9717), .A3(n9716), .A4(n9715), .ZN(n9936)
         );
  INV_X1 U10875 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10110) );
  AOI22_X1 U10876 ( .A1(n5304), .A2(keyinput54), .B1(keyinput0), .B2(n10110), 
        .ZN(n9719) );
  OAI221_X1 U10877 ( .B1(n5304), .B2(keyinput54), .C1(n10110), .C2(keyinput0), 
        .A(n9719), .ZN(n9728) );
  INV_X1 U10878 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10108) );
  AOI22_X1 U10879 ( .A1(n9721), .A2(keyinput62), .B1(keyinput71), .B2(n10108), 
        .ZN(n9720) );
  OAI221_X1 U10880 ( .B1(n9721), .B2(keyinput62), .C1(n10108), .C2(keyinput71), 
        .A(n9720), .ZN(n9727) );
  INV_X1 U10881 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10107) );
  AOI22_X1 U10882 ( .A1(n9723), .A2(keyinput105), .B1(keyinput28), .B2(n10107), 
        .ZN(n9722) );
  OAI221_X1 U10883 ( .B1(n9723), .B2(keyinput105), .C1(n10107), .C2(keyinput28), .A(n9722), .ZN(n9726) );
  AOI22_X1 U10884 ( .A1(n6712), .A2(keyinput101), .B1(n6728), .B2(keyinput60), 
        .ZN(n9724) );
  OAI221_X1 U10885 ( .B1(n6712), .B2(keyinput101), .C1(n6728), .C2(keyinput60), 
        .A(n9724), .ZN(n9725) );
  NOR4_X1 U10886 ( .A1(n9728), .A2(n9727), .A3(n9726), .A4(n9725), .ZN(n9745)
         );
  AOI22_X1 U10887 ( .A1(n9730), .A2(keyinput53), .B1(keyinput127), .B2(n9357), 
        .ZN(n9729) );
  OAI221_X1 U10888 ( .B1(n9730), .B2(keyinput53), .C1(n9357), .C2(keyinput127), 
        .A(n9729), .ZN(n9737) );
  AOI22_X1 U10889 ( .A1(n9733), .A2(keyinput88), .B1(n9732), .B2(keyinput51), 
        .ZN(n9731) );
  OAI221_X1 U10890 ( .B1(n9733), .B2(keyinput88), .C1(n9732), .C2(keyinput51), 
        .A(n9731), .ZN(n9736) );
  XNOR2_X1 U10891 ( .A(keyinput81), .B(n10300), .ZN(n9735) );
  XNOR2_X1 U10892 ( .A(keyinput78), .B(n5941), .ZN(n9734) );
  NOR4_X1 U10893 ( .A1(n9737), .A2(n9736), .A3(n9735), .A4(n9734), .ZN(n9744)
         );
  INV_X1 U10894 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9976) );
  AOI22_X1 U10895 ( .A1(n9976), .A2(keyinput6), .B1(n5926), .B2(keyinput41), 
        .ZN(n9738) );
  OAI221_X1 U10896 ( .B1(n9976), .B2(keyinput6), .C1(n5926), .C2(keyinput41), 
        .A(n9738), .ZN(n9742) );
  AOI22_X1 U10897 ( .A1(n9740), .A2(keyinput103), .B1(n5293), .B2(keyinput85), 
        .ZN(n9739) );
  OAI221_X1 U10898 ( .B1(n9740), .B2(keyinput103), .C1(n5293), .C2(keyinput85), 
        .A(n9739), .ZN(n9741) );
  NOR2_X1 U10899 ( .A1(n9742), .A2(n9741), .ZN(n9743) );
  NAND3_X1 U10900 ( .A1(n9745), .A2(n9744), .A3(n9743), .ZN(n9867) );
  INV_X1 U10901 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n9748) );
  AOI22_X1 U10902 ( .A1(n9748), .A2(keyinput69), .B1(n9747), .B2(keyinput114), 
        .ZN(n9746) );
  OAI221_X1 U10903 ( .B1(n9748), .B2(keyinput69), .C1(n9747), .C2(keyinput114), 
        .A(n9746), .ZN(n9760) );
  AOI22_X1 U10904 ( .A1(n9390), .A2(keyinput34), .B1(n9750), .B2(keyinput106), 
        .ZN(n9749) );
  OAI221_X1 U10905 ( .B1(n9390), .B2(keyinput34), .C1(n9750), .C2(keyinput106), 
        .A(n9749), .ZN(n9759) );
  INV_X1 U10906 ( .A(SI_25_), .ZN(n9753) );
  AOI22_X1 U10907 ( .A1(n9753), .A2(keyinput39), .B1(keyinput20), .B2(n9752), 
        .ZN(n9751) );
  OAI221_X1 U10908 ( .B1(n9753), .B2(keyinput39), .C1(n9752), .C2(keyinput20), 
        .A(n9751), .ZN(n9758) );
  AOI22_X1 U10909 ( .A1(n9756), .A2(keyinput50), .B1(keyinput29), .B2(n9755), 
        .ZN(n9754) );
  OAI221_X1 U10910 ( .B1(n9756), .B2(keyinput50), .C1(n9755), .C2(keyinput29), 
        .A(n9754), .ZN(n9757) );
  NOR4_X1 U10911 ( .A1(n9760), .A2(n9759), .A3(n9758), .A4(n9757), .ZN(n9793)
         );
  AOI22_X1 U10912 ( .A1(n8678), .A2(keyinput125), .B1(keyinput118), .B2(n6047), 
        .ZN(n9761) );
  OAI221_X1 U10913 ( .B1(n8678), .B2(keyinput125), .C1(n6047), .C2(keyinput118), .A(n9761), .ZN(n9769) );
  AOI22_X1 U10914 ( .A1(n9764), .A2(keyinput97), .B1(keyinput46), .B2(n9763), 
        .ZN(n9762) );
  OAI221_X1 U10915 ( .B1(n9764), .B2(keyinput97), .C1(n9763), .C2(keyinput46), 
        .A(n9762), .ZN(n9768) );
  AOI22_X1 U10916 ( .A1(n9766), .A2(keyinput79), .B1(keyinput95), .B2(n9940), 
        .ZN(n9765) );
  OAI221_X1 U10917 ( .B1(n9766), .B2(keyinput79), .C1(n9940), .C2(keyinput95), 
        .A(n9765), .ZN(n9767) );
  NOR3_X1 U10918 ( .A1(n9769), .A2(n9768), .A3(n9767), .ZN(n9792) );
  INV_X1 U10919 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10022) );
  AOI22_X1 U10920 ( .A1(n9771), .A2(keyinput19), .B1(keyinput94), .B2(n10022), 
        .ZN(n9770) );
  OAI221_X1 U10921 ( .B1(n9771), .B2(keyinput19), .C1(n10022), .C2(keyinput94), 
        .A(n9770), .ZN(n9779) );
  AOI22_X1 U10922 ( .A1(n9773), .A2(keyinput119), .B1(keyinput84), .B2(n10175), 
        .ZN(n9772) );
  OAI221_X1 U10923 ( .B1(n9773), .B2(keyinput119), .C1(n10175), .C2(keyinput84), .A(n9772), .ZN(n9778) );
  AOI22_X1 U10924 ( .A1(n9776), .A2(keyinput45), .B1(keyinput44), .B2(n9775), 
        .ZN(n9774) );
  OAI221_X1 U10925 ( .B1(n9776), .B2(keyinput45), .C1(n9775), .C2(keyinput44), 
        .A(n9774), .ZN(n9777) );
  NOR3_X1 U10926 ( .A1(n9779), .A2(n9778), .A3(n9777), .ZN(n9791) );
  AOI22_X1 U10927 ( .A1(n9781), .A2(keyinput92), .B1(keyinput25), .B2(n6908), 
        .ZN(n9780) );
  OAI221_X1 U10928 ( .B1(n9781), .B2(keyinput92), .C1(n6908), .C2(keyinput25), 
        .A(n9780), .ZN(n9789) );
  INV_X1 U10929 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9784) );
  AOI22_X1 U10930 ( .A1(n9784), .A2(keyinput98), .B1(n9783), .B2(keyinput76), 
        .ZN(n9782) );
  OAI221_X1 U10931 ( .B1(n9784), .B2(keyinput98), .C1(n9783), .C2(keyinput76), 
        .A(n9782), .ZN(n9788) );
  INV_X1 U10932 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10111) );
  AOI22_X1 U10933 ( .A1(n10111), .A2(keyinput22), .B1(keyinput18), .B2(n9786), 
        .ZN(n9785) );
  OAI221_X1 U10934 ( .B1(n10111), .B2(keyinput22), .C1(n9786), .C2(keyinput18), 
        .A(n9785), .ZN(n9787) );
  NOR3_X1 U10935 ( .A1(n9789), .A2(n9788), .A3(n9787), .ZN(n9790) );
  NAND4_X1 U10936 ( .A1(n9793), .A2(n9792), .A3(n9791), .A4(n9790), .ZN(n9866)
         );
  AOI22_X1 U10937 ( .A1(n7493), .A2(keyinput117), .B1(keyinput121), .B2(n6676), 
        .ZN(n9794) );
  OAI221_X1 U10938 ( .B1(n7493), .B2(keyinput117), .C1(n6676), .C2(keyinput121), .A(n9794), .ZN(n9835) );
  XNOR2_X1 U10939 ( .A(n9795), .B(keyinput4), .ZN(n9802) );
  XNOR2_X1 U10940 ( .A(n9796), .B(keyinput11), .ZN(n9801) );
  XNOR2_X1 U10941 ( .A(n9797), .B(keyinput67), .ZN(n9800) );
  XNOR2_X1 U10942 ( .A(n9798), .B(keyinput47), .ZN(n9799) );
  NOR4_X1 U10943 ( .A1(n9802), .A2(n9801), .A3(n9800), .A4(n9799), .ZN(n9823)
         );
  XOR2_X1 U10944 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput70), .Z(n9807) );
  XOR2_X1 U10945 ( .A(SI_0_), .B(keyinput123), .Z(n9806) );
  XNOR2_X1 U10946 ( .A(P1_U3086), .B(keyinput14), .ZN(n9805) );
  XNOR2_X1 U10947 ( .A(n9803), .B(keyinput32), .ZN(n9804) );
  NOR4_X1 U10948 ( .A1(n9807), .A2(n9806), .A3(n9805), .A4(n9804), .ZN(n9822)
         );
  XNOR2_X1 U10949 ( .A(n9808), .B(keyinput13), .ZN(n9814) );
  XOR2_X1 U10950 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput48), .Z(n9813) );
  XNOR2_X1 U10951 ( .A(n9809), .B(keyinput83), .ZN(n9812) );
  XNOR2_X1 U10952 ( .A(n9810), .B(keyinput66), .ZN(n9811) );
  NOR4_X1 U10953 ( .A1(n9814), .A2(n9813), .A3(n9812), .A4(n9811), .ZN(n9821)
         );
  XOR2_X1 U10954 ( .A(P2_IR_REG_0__SCAN_IN), .B(keyinput59), .Z(n9819) );
  XOR2_X1 U10955 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput49), .Z(n9818) );
  XNOR2_X1 U10956 ( .A(n9815), .B(keyinput111), .ZN(n9817) );
  XNOR2_X1 U10957 ( .A(keyinput52), .B(n9974), .ZN(n9816) );
  NOR4_X1 U10958 ( .A1(n9819), .A2(n9818), .A3(n9817), .A4(n9816), .ZN(n9820)
         );
  NAND4_X1 U10959 ( .A1(n9823), .A2(n9822), .A3(n9821), .A4(n9820), .ZN(n9834)
         );
  XNOR2_X1 U10960 ( .A(P1_REG2_REG_28__SCAN_IN), .B(keyinput90), .ZN(n9827) );
  XNOR2_X1 U10961 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(keyinput24), .ZN(n9826) );
  XNOR2_X1 U10962 ( .A(P2_IR_REG_12__SCAN_IN), .B(keyinput36), .ZN(n9825) );
  XNOR2_X1 U10963 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput110), .ZN(n9824) );
  NAND4_X1 U10964 ( .A1(n9827), .A2(n9826), .A3(n9825), .A4(n9824), .ZN(n9833)
         );
  XNOR2_X1 U10965 ( .A(SI_17_), .B(keyinput96), .ZN(n9831) );
  XNOR2_X1 U10966 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput74), .ZN(n9830) );
  XNOR2_X1 U10967 ( .A(P2_REG1_REG_0__SCAN_IN), .B(keyinput122), .ZN(n9829) );
  XNOR2_X1 U10968 ( .A(P1_REG2_REG_2__SCAN_IN), .B(keyinput73), .ZN(n9828) );
  NAND4_X1 U10969 ( .A1(n9831), .A2(n9830), .A3(n9829), .A4(n9828), .ZN(n9832)
         );
  OR4_X1 U10970 ( .A1(n9835), .A2(n9834), .A3(n9833), .A4(n9832), .ZN(n9865)
         );
  INV_X1 U10971 ( .A(keyinput89), .ZN(n9837) );
  AOI22_X1 U10972 ( .A1(n5774), .A2(keyinput1), .B1(P1_ADDR_REG_14__SCAN_IN), 
        .B2(n9837), .ZN(n9836) );
  OAI221_X1 U10973 ( .B1(n5774), .B2(keyinput1), .C1(n9837), .C2(
        P1_ADDR_REG_14__SCAN_IN), .A(n9836), .ZN(n9842) );
  INV_X1 U10974 ( .A(keyinput37), .ZN(n9839) );
  AOI22_X1 U10975 ( .A1(n9840), .A2(keyinput9), .B1(P2_ADDR_REG_17__SCAN_IN), 
        .B2(n9839), .ZN(n9838) );
  OAI221_X1 U10976 ( .B1(n9840), .B2(keyinput9), .C1(n9839), .C2(
        P2_ADDR_REG_17__SCAN_IN), .A(n9838), .ZN(n9841) );
  NOR2_X1 U10977 ( .A1(n9842), .A2(n9841), .ZN(n9863) );
  INV_X1 U10978 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10113) );
  AOI22_X1 U10979 ( .A1(n7254), .A2(keyinput124), .B1(n10113), .B2(keyinput17), 
        .ZN(n9843) );
  OAI221_X1 U10980 ( .B1(n7254), .B2(keyinput124), .C1(n10113), .C2(keyinput17), .A(n9843), .ZN(n9847) );
  INV_X1 U10981 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10105) );
  AOI22_X1 U10982 ( .A1(n9845), .A2(keyinput61), .B1(n10105), .B2(keyinput126), 
        .ZN(n9844) );
  OAI221_X1 U10983 ( .B1(n9845), .B2(keyinput61), .C1(n10105), .C2(keyinput126), .A(n9844), .ZN(n9846) );
  NOR2_X1 U10984 ( .A1(n9847), .A2(n9846), .ZN(n9862) );
  INV_X1 U10985 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10114) );
  AOI22_X1 U10986 ( .A1(n9954), .A2(keyinput57), .B1(n10114), .B2(keyinput80), 
        .ZN(n9848) );
  OAI221_X1 U10987 ( .B1(n9954), .B2(keyinput57), .C1(n10114), .C2(keyinput80), 
        .A(n9848), .ZN(n9852) );
  INV_X1 U10988 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n9850) );
  AOI22_X1 U10989 ( .A1(n10297), .A2(keyinput58), .B1(keyinput55), .B2(n9850), 
        .ZN(n9849) );
  OAI221_X1 U10990 ( .B1(n10297), .B2(keyinput58), .C1(n9850), .C2(keyinput55), 
        .A(n9849), .ZN(n9851) );
  NOR2_X1 U10991 ( .A1(n9852), .A2(n9851), .ZN(n9861) );
  AOI22_X1 U10992 ( .A1(n7266), .A2(keyinput100), .B1(P2_U3151), .B2(
        keyinput42), .ZN(n9853) );
  OAI221_X1 U10993 ( .B1(n7266), .B2(keyinput100), .C1(P2_U3151), .C2(
        keyinput42), .A(n9853), .ZN(n9859) );
  XNOR2_X1 U10994 ( .A(keyinput115), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n9857)
         );
  XNOR2_X1 U10995 ( .A(keyinput102), .B(P2_REG0_REG_7__SCAN_IN), .ZN(n9856) );
  XNOR2_X1 U10996 ( .A(keyinput116), .B(P2_REG0_REG_3__SCAN_IN), .ZN(n9855) );
  XNOR2_X1 U10997 ( .A(keyinput77), .B(P2_D_REG_1__SCAN_IN), .ZN(n9854) );
  NAND4_X1 U10998 ( .A1(n9857), .A2(n9856), .A3(n9855), .A4(n9854), .ZN(n9858)
         );
  NOR2_X1 U10999 ( .A1(n9859), .A2(n9858), .ZN(n9860) );
  NAND4_X1 U11000 ( .A1(n9863), .A2(n9862), .A3(n9861), .A4(n9860), .ZN(n9864)
         );
  NOR4_X1 U11001 ( .A1(n9867), .A2(n9866), .A3(n9865), .A4(n9864), .ZN(n9908)
         );
  INV_X1 U11002 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10117) );
  AOI22_X1 U11003 ( .A1(n10117), .A2(keyinput7), .B1(n9869), .B2(keyinput109), 
        .ZN(n9868) );
  OAI221_X1 U11004 ( .B1(n10117), .B2(keyinput7), .C1(n9869), .C2(keyinput109), 
        .A(n9868), .ZN(n9879) );
  AOI22_X1 U11005 ( .A1(n6876), .A2(keyinput82), .B1(n9871), .B2(keyinput8), 
        .ZN(n9870) );
  OAI221_X1 U11006 ( .B1(n6876), .B2(keyinput82), .C1(n9871), .C2(keyinput8), 
        .A(n9870), .ZN(n9878) );
  INV_X1 U11007 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10112) );
  AOI22_X1 U11008 ( .A1(n7629), .A2(keyinput16), .B1(n10112), .B2(keyinput5), 
        .ZN(n9872) );
  OAI221_X1 U11009 ( .B1(n7629), .B2(keyinput16), .C1(n10112), .C2(keyinput5), 
        .A(n9872), .ZN(n9877) );
  AOI22_X1 U11010 ( .A1(n9875), .A2(keyinput99), .B1(keyinput21), .B2(n9874), 
        .ZN(n9873) );
  OAI221_X1 U11011 ( .B1(n9875), .B2(keyinput99), .C1(n9874), .C2(keyinput21), 
        .A(n9873), .ZN(n9876) );
  NOR4_X1 U11012 ( .A1(n9879), .A2(n9878), .A3(n9877), .A4(n9876), .ZN(n9907)
         );
  AOI22_X1 U11013 ( .A1(n9987), .A2(keyinput75), .B1(n9881), .B2(keyinput113), 
        .ZN(n9880) );
  OAI221_X1 U11014 ( .B1(n9987), .B2(keyinput75), .C1(n9881), .C2(keyinput113), 
        .A(n9880), .ZN(n9890) );
  INV_X1 U11015 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10104) );
  INV_X1 U11016 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n9985) );
  AOI22_X1 U11017 ( .A1(n10104), .A2(keyinput10), .B1(keyinput23), .B2(n9985), 
        .ZN(n9882) );
  OAI221_X1 U11018 ( .B1(n10104), .B2(keyinput10), .C1(n9985), .C2(keyinput23), 
        .A(n9882), .ZN(n9889) );
  AOI22_X1 U11019 ( .A1(n9706), .A2(keyinput120), .B1(n9884), .B2(keyinput68), 
        .ZN(n9883) );
  OAI221_X1 U11020 ( .B1(n9706), .B2(keyinput120), .C1(n9884), .C2(keyinput68), 
        .A(n9883), .ZN(n9888) );
  AOI22_X1 U11021 ( .A1(n9886), .A2(keyinput91), .B1(n5879), .B2(keyinput108), 
        .ZN(n9885) );
  OAI221_X1 U11022 ( .B1(n9886), .B2(keyinput91), .C1(n5879), .C2(keyinput108), 
        .A(n9885), .ZN(n9887) );
  NOR4_X1 U11023 ( .A1(n9890), .A2(n9889), .A3(n9888), .A4(n9887), .ZN(n9906)
         );
  AOI22_X1 U11024 ( .A1(n9893), .A2(keyinput26), .B1(keyinput104), .B2(n9892), 
        .ZN(n9891) );
  OAI221_X1 U11025 ( .B1(n9893), .B2(keyinput26), .C1(n9892), .C2(keyinput104), 
        .A(n9891), .ZN(n9904) );
  AOI22_X1 U11026 ( .A1(n9895), .A2(keyinput93), .B1(keyinput87), .B2(n5843), 
        .ZN(n9894) );
  OAI221_X1 U11027 ( .B1(n9895), .B2(keyinput93), .C1(n5843), .C2(keyinput87), 
        .A(n9894), .ZN(n9903) );
  AOI22_X1 U11028 ( .A1(n9944), .A2(keyinput27), .B1(n9897), .B2(keyinput72), 
        .ZN(n9896) );
  OAI221_X1 U11029 ( .B1(n9944), .B2(keyinput27), .C1(n9897), .C2(keyinput72), 
        .A(n9896), .ZN(n9902) );
  AOI22_X1 U11030 ( .A1(n9900), .A2(keyinput64), .B1(n9899), .B2(keyinput35), 
        .ZN(n9898) );
  OAI221_X1 U11031 ( .B1(n9900), .B2(keyinput64), .C1(n9899), .C2(keyinput35), 
        .A(n9898), .ZN(n9901) );
  NOR4_X1 U11032 ( .A1(n9904), .A2(n9903), .A3(n9902), .A4(n9901), .ZN(n9905)
         );
  AND4_X1 U11033 ( .A1(n9908), .A2(n9907), .A3(n9906), .A4(n9905), .ZN(n9934)
         );
  AOI22_X1 U11034 ( .A1(n10311), .A2(keyinput15), .B1(n9705), .B2(keyinput3), 
        .ZN(n9909) );
  OAI221_X1 U11035 ( .B1(n10311), .B2(keyinput15), .C1(n9705), .C2(keyinput3), 
        .A(n9909), .ZN(n9919) );
  AOI22_X1 U11036 ( .A1(n9912), .A2(keyinput31), .B1(n9911), .B2(keyinput30), 
        .ZN(n9910) );
  OAI221_X1 U11037 ( .B1(n9912), .B2(keyinput31), .C1(n9911), .C2(keyinput30), 
        .A(n9910), .ZN(n9918) );
  INV_X1 U11038 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10109) );
  INV_X1 U11039 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10106) );
  AOI22_X1 U11040 ( .A1(n10109), .A2(keyinput65), .B1(keyinput33), .B2(n10106), 
        .ZN(n9913) );
  OAI221_X1 U11041 ( .B1(n10109), .B2(keyinput65), .C1(n10106), .C2(keyinput33), .A(n9913), .ZN(n9917) );
  INV_X1 U11042 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10115) );
  AOI22_X1 U11043 ( .A1(n9915), .A2(keyinput56), .B1(keyinput63), .B2(n10115), 
        .ZN(n9914) );
  OAI221_X1 U11044 ( .B1(n9915), .B2(keyinput56), .C1(n10115), .C2(keyinput63), 
        .A(n9914), .ZN(n9916) );
  NOR4_X1 U11045 ( .A1(n9919), .A2(n9918), .A3(n9917), .A4(n9916), .ZN(n9933)
         );
  INV_X1 U11046 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9986) );
  AOI22_X1 U11047 ( .A1(n9986), .A2(keyinput40), .B1(n9921), .B2(keyinput2), 
        .ZN(n9920) );
  OAI221_X1 U11048 ( .B1(n9986), .B2(keyinput40), .C1(n9921), .C2(keyinput2), 
        .A(n9920), .ZN(n9931) );
  AOI22_X1 U11049 ( .A1(n9924), .A2(keyinput38), .B1(n9923), .B2(keyinput43), 
        .ZN(n9922) );
  OAI221_X1 U11050 ( .B1(n9924), .B2(keyinput38), .C1(n9923), .C2(keyinput43), 
        .A(n9922), .ZN(n9930) );
  INV_X1 U11051 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10103) );
  AOI22_X1 U11052 ( .A1(n10103), .A2(keyinput86), .B1(keyinput12), .B2(n9926), 
        .ZN(n9925) );
  OAI221_X1 U11053 ( .B1(n10103), .B2(keyinput86), .C1(n9926), .C2(keyinput12), 
        .A(n9925), .ZN(n9929) );
  AOI22_X1 U11054 ( .A1(n9674), .A2(keyinput107), .B1(n5867), .B2(keyinput112), 
        .ZN(n9927) );
  OAI221_X1 U11055 ( .B1(n9674), .B2(keyinput107), .C1(n5867), .C2(keyinput112), .A(n9927), .ZN(n9928) );
  NOR4_X1 U11056 ( .A1(n9931), .A2(n9930), .A3(n9929), .A4(n9928), .ZN(n9932)
         );
  NAND3_X1 U11057 ( .A1(n9934), .A2(n9933), .A3(n9932), .ZN(n9935) );
  XOR2_X1 U11058 ( .A(n9936), .B(n9935), .Z(n9937) );
  XNOR2_X1 U11059 ( .A(n9938), .B(n9937), .ZN(P1_U3512) );
  MUX2_X1 U11060 ( .A(n9940), .B(n9939), .S(n10174), .Z(n9941) );
  OAI21_X1 U11061 ( .B1(n9942), .B2(n9956), .A(n9941), .ZN(P1_U3511) );
  MUX2_X1 U11062 ( .A(n9944), .B(n9943), .S(n10174), .Z(n9945) );
  OAI21_X1 U11063 ( .B1(n9946), .B2(n9956), .A(n9945), .ZN(P1_U3510) );
  MUX2_X1 U11064 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9947), .S(n10174), .Z(
        P1_U3509) );
  MUX2_X1 U11065 ( .A(n9949), .B(n9948), .S(n10174), .Z(n9950) );
  OAI21_X1 U11066 ( .B1(n9951), .B2(n9956), .A(n9950), .ZN(P1_U3507) );
  MUX2_X1 U11067 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9952), .S(n10174), .Z(
        P1_U3504) );
  MUX2_X1 U11068 ( .A(n9954), .B(n9953), .S(n10174), .Z(n9955) );
  OAI21_X1 U11069 ( .B1(n9957), .B2(n9956), .A(n9955), .ZN(P1_U3501) );
  MUX2_X1 U11070 ( .A(n9958), .B(P1_D_REG_1__SCAN_IN), .S(n10116), .Z(P1_U3440) );
  MUX2_X1 U11071 ( .A(n9959), .B(P1_D_REG_0__SCAN_IN), .S(n10116), .Z(P1_U3439) );
  NOR3_X1 U11072 ( .A1(n9960), .A2(n4808), .A3(P1_U3086), .ZN(n9961) );
  AOI21_X1 U11073 ( .B1(n9962), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9961), .ZN(
        n9963) );
  OAI21_X1 U11074 ( .B1(n9964), .B2(n9969), .A(n9963), .ZN(P1_U3324) );
  OAI222_X1 U11075 ( .A1(n9969), .A2(n9968), .B1(P1_U3086), .B2(n9965), .C1(
        n9967), .C2(n9966), .ZN(P1_U3326) );
  MUX2_X1 U11076 ( .A(n9970), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  NOR2_X1 U11077 ( .A1(n9972), .A2(n9971), .ZN(n10025) );
  INV_X1 U11078 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n10021) );
  NOR2_X1 U11079 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10019) );
  NOR2_X1 U11080 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10017) );
  NOR2_X1 U11081 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(P2_ADDR_REG_14__SCAN_IN), 
        .ZN(n10013) );
  NOR2_X1 U11082 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10011) );
  NOR2_X1 U11083 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10007) );
  NOR2_X1 U11084 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n10005) );
  NOR2_X1 U11085 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n10001) );
  NOR2_X1 U11086 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n9997) );
  NOR2_X1 U11087 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(P2_ADDR_REG_8__SCAN_IN), 
        .ZN(n9994) );
  NOR2_X1 U11088 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n9991) );
  NOR2_X1 U11089 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n9989) );
  AOI21_X1 U11090 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n9973), .ZN(n10335) );
  NOR2_X1 U11091 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9983) );
  NAND2_X1 U11092 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9981) );
  AOI22_X1 U11093 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .B1(n9975), .B2(n9974), .ZN(n10345) );
  NAND2_X1 U11094 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n9979) );
  AOI21_X1 U11095 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10308) );
  INV_X1 U11096 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10310) );
  NOR2_X1 U11097 ( .A1(n10311), .A2(n10310), .ZN(n10309) );
  AOI21_X1 U11098 ( .B1(n10309), .B2(P1_ADDR_REG_1__SCAN_IN), .A(
        P2_ADDR_REG_1__SCAN_IN), .ZN(n10304) );
  NOR2_X1 U11099 ( .A1(n10308), .A2(n10304), .ZN(n10343) );
  INV_X1 U11100 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n9977) );
  AOI22_X1 U11101 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .B1(n9977), .B2(n9976), .ZN(n10342) );
  NAND2_X1 U11102 ( .A1(n10343), .A2(n10342), .ZN(n9978) );
  NAND2_X1 U11103 ( .A1(n9979), .A2(n9978), .ZN(n10344) );
  NAND2_X1 U11104 ( .A1(n10345), .A2(n10344), .ZN(n9980) );
  NAND2_X1 U11105 ( .A1(n9981), .A2(n9980), .ZN(n10347) );
  XNOR2_X1 U11106 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10346) );
  NOR2_X1 U11107 ( .A1(n10347), .A2(n10346), .ZN(n9982) );
  NOR2_X1 U11108 ( .A1(n9983), .A2(n9982), .ZN(n10334) );
  NAND2_X1 U11109 ( .A1(n10335), .A2(n10334), .ZN(n9984) );
  OAI21_X1 U11110 ( .B1(n9986), .B2(n9985), .A(n9984), .ZN(n10333) );
  AOI22_X1 U11111 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n6458), .B1(
        P1_ADDR_REG_6__SCAN_IN), .B2(n9987), .ZN(n10332) );
  NOR2_X1 U11112 ( .A1(n10333), .A2(n10332), .ZN(n9988) );
  NOR2_X1 U11113 ( .A1(n9989), .A2(n9988), .ZN(n10339) );
  XNOR2_X1 U11114 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10338) );
  NOR2_X1 U11115 ( .A1(n10339), .A2(n10338), .ZN(n9990) );
  NOR2_X1 U11116 ( .A1(n9991), .A2(n9990), .ZN(n10341) );
  INV_X1 U11117 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n9992) );
  AOI22_X1 U11118 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9992), .B1(
        P2_ADDR_REG_8__SCAN_IN), .B2(n9706), .ZN(n10340) );
  NOR2_X1 U11119 ( .A1(n10341), .A2(n10340), .ZN(n9993) );
  NOR2_X1 U11120 ( .A1(n9994), .A2(n9993), .ZN(n10337) );
  AOI22_X1 U11121 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n6476), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(n9995), .ZN(n10336) );
  NOR2_X1 U11122 ( .A1(n10337), .A2(n10336), .ZN(n9996) );
  NOR2_X1 U11123 ( .A1(n9997), .A2(n9996), .ZN(n10331) );
  INV_X1 U11124 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9999) );
  AOI22_X1 U11125 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n9999), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(n9998), .ZN(n10330) );
  NOR2_X1 U11126 ( .A1(n10331), .A2(n10330), .ZN(n10000) );
  NOR2_X1 U11127 ( .A1(n10001), .A2(n10000), .ZN(n10329) );
  INV_X1 U11128 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10003) );
  AOI22_X1 U11129 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n10003), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(n10002), .ZN(n10328) );
  NOR2_X1 U11130 ( .A1(n10329), .A2(n10328), .ZN(n10004) );
  NOR2_X1 U11131 ( .A1(n10005), .A2(n10004), .ZN(n10327) );
  XNOR2_X1 U11132 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10326) );
  NOR2_X1 U11133 ( .A1(n10327), .A2(n10326), .ZN(n10006) );
  NOR2_X1 U11134 ( .A1(n10007), .A2(n10006), .ZN(n10325) );
  INV_X1 U11135 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10009) );
  AOI22_X1 U11136 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(n10009), .B1(
        P1_ADDR_REG_13__SCAN_IN), .B2(n10008), .ZN(n10324) );
  NOR2_X1 U11137 ( .A1(n10325), .A2(n10324), .ZN(n10010) );
  NOR2_X1 U11138 ( .A1(n10011), .A2(n10010), .ZN(n10323) );
  XNOR2_X1 U11139 ( .A(P1_ADDR_REG_14__SCAN_IN), .B(P2_ADDR_REG_14__SCAN_IN), 
        .ZN(n10322) );
  NOR2_X1 U11140 ( .A1(n10323), .A2(n10322), .ZN(n10012) );
  NOR2_X1 U11141 ( .A1(n10013), .A2(n10012), .ZN(n10321) );
  INV_X1 U11142 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10015) );
  AOI22_X1 U11143 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n10015), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n10014), .ZN(n10320) );
  NOR2_X1 U11144 ( .A1(n10321), .A2(n10320), .ZN(n10016) );
  NOR2_X1 U11145 ( .A1(n10017), .A2(n10016), .ZN(n10319) );
  XNOR2_X1 U11146 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10318) );
  NOR2_X1 U11147 ( .A1(n10319), .A2(n10318), .ZN(n10018) );
  NOR2_X1 U11148 ( .A1(n10019), .A2(n10018), .ZN(n10317) );
  AOI22_X1 U11149 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n10021), .B1(
        P2_ADDR_REG_17__SCAN_IN), .B2(n10022), .ZN(n10316) );
  NOR2_X1 U11150 ( .A1(n10317), .A2(n10316), .ZN(n10020) );
  AOI21_X1 U11151 ( .B1(n10022), .B2(n10021), .A(n10020), .ZN(n10313) );
  NOR2_X1 U11152 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10313), .ZN(n10023) );
  NAND2_X1 U11153 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10313), .ZN(n10312) );
  OAI21_X1 U11154 ( .B1(n10023), .B2(n10314), .A(n10312), .ZN(n10024) );
  XOR2_X1 U11155 ( .A(n10025), .B(n10024), .Z(ADD_1068_U4) );
  OAI211_X1 U11156 ( .C1(n4656), .C2(n10159), .A(n10027), .B(n10026), .ZN(
        n10028) );
  AOI21_X1 U11157 ( .B1(n10029), .B2(n10161), .A(n10028), .ZN(n10030) );
  AOI22_X1 U11158 ( .A1(n10186), .A2(n10030), .B1(n5969), .B2(n10184), .ZN(
        P1_U3537) );
  AOI22_X1 U11159 ( .A1(n10174), .A2(n10030), .B1(n5968), .B2(n10173), .ZN(
        P1_U3498) );
  XNOR2_X1 U11160 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  NOR2_X1 U11161 ( .A1(n10031), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10033) );
  OR2_X1 U11162 ( .A1(n10032), .A2(n10033), .ZN(n10036) );
  INV_X1 U11163 ( .A(n10033), .ZN(n10035) );
  MUX2_X1 U11164 ( .A(n10036), .B(n10035), .S(n10034), .Z(n10038) );
  NAND2_X1 U11165 ( .A1(n10038), .A2(n10037), .ZN(n10040) );
  AOI22_X1 U11166 ( .A1(n10043), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n10039) );
  OAI21_X1 U11167 ( .B1(n10041), .B2(n10040), .A(n10039), .ZN(P1_U3243) );
  AOI22_X1 U11168 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(n10043), .B1(
        P1_REG3_REG_4__SCAN_IN), .B2(P1_U3086), .ZN(n10060) );
  AOI211_X1 U11169 ( .C1(n10047), .C2(n10046), .A(n10045), .B(n10044), .ZN(
        n10050) );
  INV_X1 U11170 ( .A(n10048), .ZN(n10049) );
  AOI211_X1 U11171 ( .C1(n10052), .C2(n10051), .A(n10050), .B(n10049), .ZN(
        n10059) );
  NAND2_X1 U11172 ( .A1(n10054), .A2(n10053), .ZN(n10055) );
  NAND3_X1 U11173 ( .A1(n10057), .A2(n10056), .A3(n10055), .ZN(n10058) );
  NAND3_X1 U11174 ( .A1(n10060), .A2(n10059), .A3(n10058), .ZN(P1_U3247) );
  NAND2_X1 U11175 ( .A1(n10061), .A2(n10081), .ZN(n10064) );
  AOI22_X1 U11176 ( .A1(n10102), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n10062), 
        .B2(n10091), .ZN(n10063) );
  OAI211_X1 U11177 ( .C1(n10065), .C2(n10096), .A(n10064), .B(n10063), .ZN(
        n10066) );
  AOI21_X1 U11178 ( .B1(n10082), .B2(n10067), .A(n10066), .ZN(n10068) );
  OAI21_X1 U11179 ( .B1(n10102), .B2(n10069), .A(n10068), .ZN(P1_U3288) );
  XNOR2_X1 U11180 ( .A(n10070), .B(n10076), .ZN(n10073) );
  AOI21_X1 U11181 ( .B1(n10073), .B2(n10072), .A(n10071), .ZN(n10125) );
  AOI222_X1 U11182 ( .A1(n5795), .A2(n10074), .B1(P1_REG2_REG_2__SCAN_IN), 
        .B2(n10102), .C1(n10091), .C2(P1_REG3_REG_2__SCAN_IN), .ZN(n10084) );
  XNOR2_X1 U11183 ( .A(n10075), .B(n10076), .ZN(n10128) );
  INV_X1 U11184 ( .A(n10093), .ZN(n10079) );
  INV_X1 U11185 ( .A(n10077), .ZN(n10078) );
  OAI211_X1 U11186 ( .C1(n5796), .C2(n10079), .A(n10078), .B(n10094), .ZN(
        n10124) );
  INV_X1 U11187 ( .A(n10124), .ZN(n10080) );
  AOI22_X1 U11188 ( .A1(n10128), .A2(n10082), .B1(n10081), .B2(n10080), .ZN(
        n10083) );
  OAI211_X1 U11189 ( .C1(n10102), .C2(n10125), .A(n10084), .B(n10083), .ZN(
        P1_U3291) );
  XNOR2_X1 U11190 ( .A(n10085), .B(n6108), .ZN(n10123) );
  XNOR2_X1 U11191 ( .A(n6108), .B(n10086), .ZN(n10088) );
  NOR2_X1 U11192 ( .A1(n10088), .A2(n10087), .ZN(n10089) );
  AOI211_X1 U11193 ( .C1(n10123), .C2(n10172), .A(n10090), .B(n10089), .ZN(
        n10120) );
  AOI22_X1 U11194 ( .A1(n10091), .A2(P1_REG3_REG_1__SCAN_IN), .B1(
        P1_REG2_REG_1__SCAN_IN), .B2(n10102), .ZN(n10101) );
  NOR2_X1 U11195 ( .A1(n10102), .A2(n10092), .ZN(n10099) );
  OAI211_X1 U11196 ( .C1(n10095), .C2(n6106), .A(n10094), .B(n10093), .ZN(
        n10119) );
  OAI22_X1 U11197 ( .A1(n10097), .A2(n10119), .B1(n6106), .B2(n10096), .ZN(
        n10098) );
  AOI21_X1 U11198 ( .B1(n10123), .B2(n10099), .A(n10098), .ZN(n10100) );
  OAI211_X1 U11199 ( .C1(n10102), .C2(n10120), .A(n10101), .B(n10100), .ZN(
        P1_U3292) );
  AND2_X1 U11200 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10116), .ZN(P1_U3294) );
  AND2_X1 U11201 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10116), .ZN(P1_U3295) );
  NOR2_X1 U11202 ( .A1(n10118), .A2(n10103), .ZN(P1_U3296) );
  NOR2_X1 U11203 ( .A1(n10118), .A2(n10104), .ZN(P1_U3297) );
  NOR2_X1 U11204 ( .A1(n10118), .A2(n10105), .ZN(P1_U3298) );
  AND2_X1 U11205 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10116), .ZN(P1_U3299) );
  AND2_X1 U11206 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10116), .ZN(P1_U3300) );
  NOR2_X1 U11207 ( .A1(n10118), .A2(n10106), .ZN(P1_U3301) );
  AND2_X1 U11208 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10116), .ZN(P1_U3302) );
  AND2_X1 U11209 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10116), .ZN(P1_U3303) );
  NOR2_X1 U11210 ( .A1(n10118), .A2(n10107), .ZN(P1_U3304) );
  NOR2_X1 U11211 ( .A1(n10118), .A2(n10108), .ZN(P1_U3305) );
  NOR2_X1 U11212 ( .A1(n10118), .A2(n10109), .ZN(P1_U3306) );
  NOR2_X1 U11213 ( .A1(n10118), .A2(n10110), .ZN(P1_U3307) );
  NOR2_X1 U11214 ( .A1(n10118), .A2(n10111), .ZN(P1_U3308) );
  NOR2_X1 U11215 ( .A1(n10118), .A2(n10112), .ZN(P1_U3309) );
  AND2_X1 U11216 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10116), .ZN(P1_U3310) );
  AND2_X1 U11217 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10116), .ZN(P1_U3311) );
  NOR2_X1 U11218 ( .A1(n10118), .A2(n10113), .ZN(P1_U3312) );
  AND2_X1 U11219 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10116), .ZN(P1_U3313) );
  NOR2_X1 U11220 ( .A1(n10118), .A2(n10114), .ZN(P1_U3314) );
  AND2_X1 U11221 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10116), .ZN(P1_U3315) );
  AND2_X1 U11222 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10116), .ZN(P1_U3316) );
  NOR2_X1 U11223 ( .A1(n10118), .A2(n10115), .ZN(P1_U3317) );
  AND2_X1 U11224 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10116), .ZN(P1_U3318) );
  AND2_X1 U11225 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10116), .ZN(P1_U3319) );
  AND2_X1 U11226 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10116), .ZN(P1_U3320) );
  AND2_X1 U11227 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10116), .ZN(P1_U3321) );
  AND2_X1 U11228 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10116), .ZN(P1_U3322) );
  NOR2_X1 U11229 ( .A1(n10118), .A2(n10117), .ZN(P1_U3323) );
  OAI21_X1 U11230 ( .B1(n6106), .B2(n10159), .A(n10119), .ZN(n10122) );
  INV_X1 U11231 ( .A(n10120), .ZN(n10121) );
  AOI211_X1 U11232 ( .C1(n10148), .C2(n10123), .A(n10122), .B(n10121), .ZN(
        n10176) );
  AOI22_X1 U11233 ( .A1(n10174), .A2(n10176), .B1(n5762), .B2(n10173), .ZN(
        P1_U3456) );
  OAI21_X1 U11234 ( .B1(n5796), .B2(n10159), .A(n10124), .ZN(n10127) );
  INV_X1 U11235 ( .A(n10125), .ZN(n10126) );
  AOI211_X1 U11236 ( .C1(n10161), .C2(n10128), .A(n10127), .B(n10126), .ZN(
        n10177) );
  AOI22_X1 U11237 ( .A1(n10174), .A2(n10177), .B1(n5791), .B2(n10173), .ZN(
        P1_U3459) );
  INV_X1 U11238 ( .A(n10129), .ZN(n10133) );
  OAI21_X1 U11239 ( .B1(n5810), .B2(n10159), .A(n10130), .ZN(n10132) );
  AOI211_X1 U11240 ( .C1(n10161), .C2(n10133), .A(n10132), .B(n10131), .ZN(
        n10178) );
  AOI22_X1 U11241 ( .A1(n10174), .A2(n10178), .B1(n5799), .B2(n10173), .ZN(
        P1_U3462) );
  OAI21_X1 U11242 ( .B1(n10135), .B2(n10159), .A(n10134), .ZN(n10138) );
  INV_X1 U11243 ( .A(n10136), .ZN(n10137) );
  AOI211_X1 U11244 ( .C1(n10161), .C2(n10139), .A(n10138), .B(n10137), .ZN(
        n10179) );
  AOI22_X1 U11245 ( .A1(n10174), .A2(n10179), .B1(n5814), .B2(n10173), .ZN(
        P1_U3465) );
  OAI211_X1 U11246 ( .C1(n10142), .C2(n10159), .A(n10141), .B(n10140), .ZN(
        n10143) );
  AOI21_X1 U11247 ( .B1(n10161), .B2(n10144), .A(n10143), .ZN(n10180) );
  AOI22_X1 U11248 ( .A1(n10174), .A2(n10180), .B1(n5879), .B2(n10173), .ZN(
        P1_U3480) );
  OAI21_X1 U11249 ( .B1(n10146), .B2(n10159), .A(n10145), .ZN(n10147) );
  AOI21_X1 U11250 ( .B1(n10149), .B2(n10148), .A(n10147), .ZN(n10150) );
  AOI22_X1 U11251 ( .A1(n10174), .A2(n10181), .B1(n5916), .B2(n10173), .ZN(
        P1_U3486) );
  OAI211_X1 U11252 ( .C1(n10154), .C2(n10159), .A(n10153), .B(n10152), .ZN(
        n10155) );
  AOI21_X1 U11253 ( .B1(n10156), .B2(n10161), .A(n10155), .ZN(n10182) );
  AOI22_X1 U11254 ( .A1(n10174), .A2(n10182), .B1(n5929), .B2(n10173), .ZN(
        P1_U3489) );
  OAI211_X1 U11255 ( .C1(n4692), .C2(n10159), .A(n10158), .B(n10157), .ZN(
        n10160) );
  AOI21_X1 U11256 ( .B1(n10162), .B2(n10161), .A(n10160), .ZN(n10183) );
  AOI22_X1 U11257 ( .A1(n10174), .A2(n10183), .B1(n5941), .B2(n10173), .ZN(
        P1_U3492) );
  AOI21_X1 U11258 ( .B1(n10165), .B2(n10164), .A(n10163), .ZN(n10166) );
  OAI211_X1 U11259 ( .C1(n10169), .C2(n10168), .A(n10167), .B(n10166), .ZN(
        n10170) );
  AOI21_X1 U11260 ( .B1(n10172), .B2(n10171), .A(n10170), .ZN(n10185) );
  AOI22_X1 U11261 ( .A1(n10174), .A2(n10185), .B1(n5957), .B2(n10173), .ZN(
        P1_U3495) );
  AOI22_X1 U11262 ( .A1(n10186), .A2(n10176), .B1(n10175), .B2(n10184), .ZN(
        P1_U3523) );
  AOI22_X1 U11263 ( .A1(n10186), .A2(n10177), .B1(n6380), .B2(n10184), .ZN(
        P1_U3524) );
  AOI22_X1 U11264 ( .A1(n10186), .A2(n10178), .B1(n6376), .B2(n10184), .ZN(
        P1_U3525) );
  AOI22_X1 U11265 ( .A1(n10186), .A2(n10179), .B1(n5812), .B2(n10184), .ZN(
        P1_U3526) );
  AOI22_X1 U11266 ( .A1(n10186), .A2(n10180), .B1(n6468), .B2(n10184), .ZN(
        P1_U3531) );
  AOI22_X1 U11267 ( .A1(n10186), .A2(n10181), .B1(n6794), .B2(n10184), .ZN(
        P1_U3533) );
  AOI22_X1 U11268 ( .A1(n10186), .A2(n10182), .B1(n5930), .B2(n10184), .ZN(
        P1_U3534) );
  AOI22_X1 U11269 ( .A1(n10186), .A2(n10183), .B1(n7082), .B2(n10184), .ZN(
        P1_U3535) );
  AOI22_X1 U11270 ( .A1(n10186), .A2(n10185), .B1(n7266), .B2(n10184), .ZN(
        P1_U3536) );
  AOI22_X1 U11271 ( .A1(n10213), .A2(P2_IR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .ZN(n10191) );
  XNOR2_X1 U11272 ( .A(n10187), .B(P2_IR_REG_0__SCAN_IN), .ZN(n10188) );
  OAI21_X1 U11273 ( .B1(n10189), .B2(n10225), .A(n10188), .ZN(n10190) );
  OAI211_X1 U11274 ( .C1(n10310), .C2(n10192), .A(n10191), .B(n10190), .ZN(
        P2_U3182) );
  INV_X1 U11275 ( .A(n10193), .ZN(n10195) );
  OAI21_X1 U11276 ( .B1(n10195), .B2(P2_REG1_REG_1__SCAN_IN), .A(n10194), .ZN(
        n10196) );
  AOI22_X1 U11277 ( .A1(n10212), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(n10197), 
        .B2(n10196), .ZN(n10202) );
  OAI211_X1 U11278 ( .C1(n10200), .C2(n10199), .A(n10198), .B(n10225), .ZN(
        n10201) );
  OAI211_X1 U11279 ( .C1(n10204), .C2(n10203), .A(n10202), .B(n10201), .ZN(
        n10205) );
  INV_X1 U11280 ( .A(n10205), .ZN(n10211) );
  INV_X1 U11281 ( .A(n10206), .ZN(n10207) );
  AOI21_X1 U11282 ( .B1(n6849), .B2(n10208), .A(n10207), .ZN(n10209) );
  OR2_X1 U11283 ( .A1(n10220), .A2(n10209), .ZN(n10210) );
  OAI211_X1 U11284 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n6734), .A(n10211), .B(
        n10210), .ZN(P2_U3183) );
  AOI22_X1 U11285 ( .A1(n10214), .A2(n10213), .B1(n10212), .B2(
        P2_ADDR_REG_17__SCAN_IN), .ZN(n10233) );
  AOI21_X1 U11286 ( .B1(n10217), .B2(n10216), .A(n10215), .ZN(n10230) );
  AOI21_X1 U11287 ( .B1(n8717), .B2(n10219), .A(n10218), .ZN(n10221) );
  OR2_X1 U11288 ( .A1(n10221), .A2(n10220), .ZN(n10228) );
  OAI21_X1 U11289 ( .B1(n10224), .B2(n10223), .A(n10222), .ZN(n10226) );
  NAND2_X1 U11290 ( .A1(n10226), .A2(n10225), .ZN(n10227) );
  OAI211_X1 U11291 ( .C1(n10230), .C2(n10229), .A(n10228), .B(n10227), .ZN(
        n10231) );
  INV_X1 U11292 ( .A(n10231), .ZN(n10232) );
  OAI211_X1 U11293 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10234), .A(n10233), .B(
        n10232), .ZN(P2_U3199) );
  INV_X1 U11294 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10239) );
  INV_X1 U11295 ( .A(n10235), .ZN(n10238) );
  OAI22_X1 U11296 ( .A1(n10236), .A2(n10268), .B1(n6186), .B2(n10274), .ZN(
        n10237) );
  NOR2_X1 U11297 ( .A1(n10238), .A2(n10237), .ZN(n10288) );
  AOI22_X1 U11298 ( .A1(n10287), .A2(n10239), .B1(n10288), .B2(n10286), .ZN(
        P2_U3393) );
  INV_X1 U11299 ( .A(n10268), .ZN(n10241) );
  AOI22_X1 U11300 ( .A1(n10242), .A2(n10241), .B1(n10281), .B2(n10240), .ZN(
        n10243) );
  AND2_X1 U11301 ( .A1(n10244), .A2(n10243), .ZN(n10290) );
  AOI22_X1 U11302 ( .A1(n10287), .A2(n9705), .B1(n10290), .B2(n10286), .ZN(
        P2_U3396) );
  INV_X1 U11303 ( .A(n10245), .ZN(n10250) );
  OAI22_X1 U11304 ( .A1(n10248), .A2(n10247), .B1(n10246), .B2(n10274), .ZN(
        n10249) );
  NOR2_X1 U11305 ( .A1(n10250), .A2(n10249), .ZN(n10292) );
  AOI22_X1 U11306 ( .A1(n10287), .A2(n5225), .B1(n10292), .B2(n10286), .ZN(
        P2_U3399) );
  OAI21_X1 U11307 ( .B1(n10252), .B2(n10274), .A(n10251), .ZN(n10253) );
  AOI21_X1 U11308 ( .B1(n10254), .B2(n10279), .A(n10253), .ZN(n10293) );
  AOI22_X1 U11309 ( .A1(n10287), .A2(n5265), .B1(n10293), .B2(n10286), .ZN(
        P2_U3408) );
  OAI22_X1 U11310 ( .A1(n10256), .A2(n10268), .B1(n10255), .B2(n10274), .ZN(
        n10257) );
  NOR2_X1 U11311 ( .A1(n10258), .A2(n10257), .ZN(n10294) );
  AOI22_X1 U11312 ( .A1(n10287), .A2(n10259), .B1(n10294), .B2(n10286), .ZN(
        P2_U3411) );
  OAI21_X1 U11313 ( .B1(n10261), .B2(n10274), .A(n10260), .ZN(n10262) );
  AOI21_X1 U11314 ( .B1(n10279), .B2(n10263), .A(n10262), .ZN(n10296) );
  AOI22_X1 U11315 ( .A1(n10287), .A2(n5293), .B1(n10296), .B2(n10286), .ZN(
        P2_U3414) );
  NOR2_X1 U11316 ( .A1(n10264), .A2(n10268), .ZN(n10266) );
  AOI211_X1 U11317 ( .C1(n10281), .C2(n10267), .A(n10266), .B(n10265), .ZN(
        n10298) );
  AOI22_X1 U11318 ( .A1(n10287), .A2(n5307), .B1(n10298), .B2(n10286), .ZN(
        P2_U3417) );
  INV_X1 U11319 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10273) );
  NOR2_X1 U11320 ( .A1(n10269), .A2(n10268), .ZN(n10271) );
  AOI211_X1 U11321 ( .C1(n10281), .C2(n10272), .A(n10271), .B(n10270), .ZN(
        n10299) );
  AOI22_X1 U11322 ( .A1(n10287), .A2(n10273), .B1(n10299), .B2(n10286), .ZN(
        P2_U3420) );
  NOR2_X1 U11323 ( .A1(n10275), .A2(n10274), .ZN(n10277) );
  AOI211_X1 U11324 ( .C1(n10279), .C2(n10278), .A(n10277), .B(n10276), .ZN(
        n10301) );
  AOI22_X1 U11325 ( .A1(n10287), .A2(n5348), .B1(n10301), .B2(n10286), .ZN(
        P2_U3423) );
  NAND2_X1 U11326 ( .A1(n10280), .A2(n10279), .ZN(n10285) );
  NAND2_X1 U11327 ( .A1(n10282), .A2(n10281), .ZN(n10283) );
  AND3_X1 U11328 ( .A1(n10285), .A2(n10284), .A3(n10283), .ZN(n10302) );
  AOI22_X1 U11329 ( .A1(n10287), .A2(n5364), .B1(n10302), .B2(n10286), .ZN(
        P2_U3426) );
  AOI22_X1 U11330 ( .A1(n10303), .A2(n10288), .B1(n6490), .B2(n6312), .ZN(
        P2_U3460) );
  AOI22_X1 U11331 ( .A1(n10303), .A2(n10290), .B1(n10289), .B2(n6312), .ZN(
        P2_U3461) );
  AOI22_X1 U11332 ( .A1(n10303), .A2(n10292), .B1(n10291), .B2(n6312), .ZN(
        P2_U3462) );
  AOI22_X1 U11333 ( .A1(n10303), .A2(n10293), .B1(n6754), .B2(n6312), .ZN(
        P2_U3465) );
  AOI22_X1 U11334 ( .A1(n10303), .A2(n10294), .B1(n6908), .B2(n6312), .ZN(
        P2_U3466) );
  INV_X1 U11335 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10295) );
  AOI22_X1 U11336 ( .A1(n10303), .A2(n10296), .B1(n10295), .B2(n6312), .ZN(
        P2_U3467) );
  AOI22_X1 U11337 ( .A1(n10303), .A2(n10298), .B1(n10297), .B2(n6312), .ZN(
        P2_U3468) );
  AOI22_X1 U11338 ( .A1(n10303), .A2(n10299), .B1(n5328), .B2(n6312), .ZN(
        P2_U3469) );
  AOI22_X1 U11339 ( .A1(n10303), .A2(n10301), .B1(n10300), .B2(n6312), .ZN(
        P2_U3470) );
  AOI22_X1 U11340 ( .A1(n10303), .A2(n10302), .B1(n7412), .B2(n6312), .ZN(
        P2_U3471) );
  INV_X1 U11341 ( .A(n10304), .ZN(n10307) );
  AOI21_X1 U11342 ( .B1(n10309), .B2(P1_ADDR_REG_1__SCAN_IN), .A(n10308), .ZN(
        n10306) );
  INV_X1 U11343 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10305) );
  OAI22_X1 U11344 ( .A1(n10308), .A2(n10307), .B1(n10306), .B2(n10305), .ZN(
        ADD_1068_U5) );
  AOI21_X1 U11345 ( .B1(n10311), .B2(n10310), .A(n10309), .ZN(ADD_1068_U46) );
  OAI21_X1 U11346 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n10313), .A(n10312), 
        .ZN(n10315) );
  XOR2_X1 U11347 ( .A(n10315), .B(n10314), .Z(ADD_1068_U55) );
  XNOR2_X1 U11348 ( .A(n10317), .B(n10316), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11349 ( .A(n10319), .B(n10318), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11350 ( .A(n10321), .B(n10320), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11351 ( .A(n10323), .B(n10322), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11352 ( .A(n10325), .B(n10324), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11353 ( .A(n10327), .B(n10326), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11354 ( .A(n10329), .B(n10328), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11355 ( .A(n10331), .B(n10330), .ZN(ADD_1068_U63) );
  XNOR2_X1 U11356 ( .A(n10333), .B(n10332), .ZN(ADD_1068_U50) );
  XOR2_X1 U11357 ( .A(n10335), .B(n10334), .Z(ADD_1068_U51) );
  XNOR2_X1 U11358 ( .A(n10337), .B(n10336), .ZN(ADD_1068_U47) );
  XNOR2_X1 U11359 ( .A(n10339), .B(n10338), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11360 ( .A(n10341), .B(n10340), .ZN(ADD_1068_U48) );
  XOR2_X1 U11361 ( .A(n10343), .B(n10342), .Z(ADD_1068_U54) );
  XOR2_X1 U11362 ( .A(n10345), .B(n10344), .Z(ADD_1068_U53) );
  XNOR2_X1 U11363 ( .A(n10347), .B(n10346), .ZN(ADD_1068_U52) );
  INV_X4 U4972 ( .A(n5188), .ZN(n5461) );
  CLKBUF_X1 U4899 ( .A(n5768), .Z(n7820) );
  CLKBUF_X1 U4914 ( .A(n6130), .Z(n9246) );
endmodule

