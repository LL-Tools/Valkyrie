

module b14_C_gen_AntiSAT_k_128_5 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, 
        U3344, U3343, U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, 
        U3334, U3333, U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, 
        U3324, U3323, U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, 
        U3316, U3315, U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, 
        U3306, U3305, U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, 
        U3296, U3295, U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, 
        U3475, U3477, U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, 
        U3495, U3497, U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, 
        U3510, U3511, U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, 
        U3520, U3521, U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, 
        U3530, U3531, U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, 
        U3540, U3541, U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, 
        U3290, U3289, U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, 
        U3280, U3279, U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, 
        U3270, U3269, U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, 
        U3261, U3260, U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, 
        U3251, U3250, U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, 
        U3241, U3240, U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, 
        U3558, U3559, U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, 
        U3568, U3569, U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, 
        U3578, U3579, U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, 
        U3233, U3232, U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, 
        U3223, U3222, U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, 
        U3213, U3212, U3211, U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761;

  INV_X2 U2290 ( .A(n3645), .ZN(n3641) );
  CLKBUF_X1 U2291 ( .A(n4300), .Z(n2048) );
  NOR2_X1 U2292 ( .A1(n2879), .A2(n2855), .ZN(n4300) );
  XNOR2_X1 U2293 ( .A(n4028), .B(n4050), .ZN(n4029) );
  OAI22_X1 U2294 ( .A1(n4029), .A2(n4502), .B1(n4028), .B2(n4050), .ZN(n4402)
         );
  AND3_X1 U2295 ( .A1(n2319), .A2(n2320), .A3(n2321), .ZN(n2542) );
  NAND2_X1 U2296 ( .A1(n3634), .A2(n3743), .ZN(n3712) );
  NOR2_X1 U2297 ( .A1(n4112), .A2(n4251), .ZN(n4094) );
  NOR2_X2 U2299 ( .A1(n3167), .A2(n3395), .ZN(n3316) );
  XNOR2_X1 U2300 ( .A(n2399), .B(IR_REG_2__SCAN_IN), .ZN(n4392) );
  NAND3_X2 U2301 ( .A1(n4383), .A2(n2714), .A3(n4382), .ZN(n2968) );
  OAI21_X1 U2302 ( .B1(n3712), .B2(n2278), .A(n2274), .ZN(n3670) );
  OR2_X1 U2303 ( .A1(n3702), .A2(n3697), .ZN(n2315) );
  NAND2_X1 U2304 ( .A1(n3763), .A2(n3623), .ZN(n3676) );
  NAND2_X1 U2305 ( .A1(n2315), .A2(n2313), .ZN(n3763) );
  NAND2_X1 U2306 ( .A1(n2618), .A2(n2157), .ZN(n4140) );
  NOR2_X1 U2307 ( .A1(n2058), .A2(n2233), .ZN(n4039) );
  OR2_X1 U2308 ( .A1(n3339), .A2(n2544), .ZN(n3360) );
  OAI22_X1 U2309 ( .A1(n4442), .A2(n4438), .B1(REG2_REG_13__SCAN_IN), .B2(
        n4046), .ZN(n4036) );
  NOR2_X1 U2310 ( .A1(n2050), .A2(n4190), .ZN(n4191) );
  NOR2_X1 U2311 ( .A1(n3124), .A2(n2061), .ZN(n3186) );
  NOR2_X1 U2312 ( .A1(n3428), .A2(n4323), .ZN(n3464) );
  AND3_X1 U2313 ( .A1(n2197), .A2(n2196), .A3(n2195), .ZN(n3108) );
  INV_X1 U2314 ( .A(n3167), .ZN(n3273) );
  INV_X1 U2315 ( .A(n2207), .ZN(n2206) );
  AOI21_X1 U2316 ( .B1(n2207), .B2(n2203), .A(n2053), .ZN(n2202) );
  INV_X2 U2317 ( .A(n4213), .ZN(n4519) );
  AND3_X1 U2318 ( .A1(n2236), .A2(n2234), .A3(n2089), .ZN(n4028) );
  AND2_X2 U2319 ( .A1(n2878), .A2(n4500), .ZN(n3779) );
  NAND2_X1 U2320 ( .A1(n3913), .A2(n2660), .ZN(n2659) );
  NAND2_X4 U2321 ( .A1(n2813), .A2(n2968), .ZN(n3645) );
  NAND2_X2 U2322 ( .A1(n2812), .A2(n2968), .ZN(n3657) );
  NAND2_X2 U2323 ( .A1(n2812), .A2(n2864), .ZN(n3658) );
  NAND2_X1 U2324 ( .A1(n2069), .A2(n2143), .ZN(n3149) );
  AND2_X2 U2325 ( .A1(n2343), .A2(n2755), .ZN(n2414) );
  AND2_X1 U2326 ( .A1(n2542), .A2(n2541), .ZN(n2575) );
  AND2_X1 U2327 ( .A1(n2574), .A2(n2302), .ZN(n2301) );
  NOR2_X1 U2328 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2398)
         );
  NAND2_X1 U2329 ( .A1(n2692), .A2(n2170), .ZN(n2351) );
  NAND2_X1 U2330 ( .A1(n2691), .A2(IR_REG_28__SCAN_IN), .ZN(n2352) );
  NAND2_X1 U2331 ( .A1(n2261), .A2(n2476), .ZN(n2260) );
  OR2_X1 U2332 ( .A1(n3070), .A2(n2456), .ZN(n2162) );
  OR2_X1 U2333 ( .A1(n2368), .A2(n4596), .ZN(n2620) );
  NAND2_X1 U2334 ( .A1(n2490), .A2(n2256), .ZN(n2255) );
  NOR2_X1 U2335 ( .A1(n2500), .A2(n2257), .ZN(n2256) );
  INV_X1 U2336 ( .A(n2489), .ZN(n2257) );
  AOI21_X1 U2337 ( .B1(n2221), .B2(n3212), .A(n3211), .ZN(n2219) );
  INV_X1 U2338 ( .A(n3014), .ZN(n2200) );
  INV_X1 U2339 ( .A(n2232), .ZN(n2230) );
  AND2_X1 U2340 ( .A1(n4044), .A2(REG2_REG_15__SCAN_IN), .ZN(n2233) );
  NAND2_X1 U2341 ( .A1(n3192), .A2(n3131), .ZN(n2164) );
  NAND2_X1 U2342 ( .A1(n3117), .A2(n3051), .ZN(n3921) );
  NAND2_X1 U2343 ( .A1(n2920), .A2(n2411), .ZN(n3058) );
  NOR2_X1 U2344 ( .A1(n4004), .A2(n2977), .ZN(n2410) );
  AND4_X1 U2345 ( .A1(n2331), .A2(n2318), .A3(n2317), .A4(n2316), .ZN(n2319)
         );
  NOR2_X1 U2346 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2317)
         );
  NOR2_X1 U2347 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2318)
         );
  INV_X1 U2348 ( .A(n2405), .ZN(n2320) );
  NAND2_X1 U2349 ( .A1(n3442), .A2(n3443), .ZN(n2216) );
  AOI21_X1 U2350 ( .B1(n3623), .B2(n2311), .A(n2310), .ZN(n2309) );
  AOI22_X1 U2351 ( .A1(n2387), .A2(n2960), .B1(n3189), .B2(n3149), .ZN(n2909)
         );
  OR2_X1 U2352 ( .A1(n2620), .A2(n2328), .ZN(n2622) );
  NOR2_X1 U2353 ( .A1(n2801), .A2(n2431), .ZN(n2122) );
  NAND2_X1 U2354 ( .A1(n4422), .A2(n4423), .ZN(n4421) );
  XNOR2_X1 U2355 ( .A(n4034), .B(n4531), .ZN(n4430) );
  NAND2_X1 U2356 ( .A1(n4470), .A2(n2560), .ZN(n4469) );
  NAND2_X1 U2357 ( .A1(n4478), .A2(n4480), .ZN(n4479) );
  AOI21_X1 U2358 ( .B1(n2248), .B2(n2055), .A(n2083), .ZN(n4160) );
  AOI21_X1 U2359 ( .B1(n2176), .B2(n2173), .A(n2171), .ZN(n4226) );
  OAI21_X1 U2360 ( .B1(n2596), .B2(n2172), .A(n2078), .ZN(n2171) );
  AND2_X1 U2361 ( .A1(n2174), .A2(n2605), .ZN(n2173) );
  NAND2_X1 U2362 ( .A1(n3996), .A2(n3282), .ZN(n2258) );
  NOR2_X1 U2363 ( .A1(n2259), .A2(n2488), .ZN(n2158) );
  OAI211_X1 U2364 ( .C1(IR_REG_31__SCAN_IN), .C2(IR_REG_29__SCAN_IN), .A(n2339), .B(n2095), .ZN(n2342) );
  NAND2_X1 U2365 ( .A1(n2051), .A2(n2084), .ZN(n2095) );
  NAND2_X1 U2366 ( .A1(n2181), .A2(n2180), .ZN(n2183) );
  NOR2_X1 U2367 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2316)
         );
  NOR2_X1 U2368 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2572)
         );
  AND2_X1 U2369 ( .A1(n2283), .A2(n2077), .ZN(n2231) );
  INV_X1 U2370 ( .A(n2280), .ZN(n2227) );
  AOI21_X1 U2371 ( .B1(n2283), .B2(n2286), .A(n2281), .ZN(n2280) );
  INV_X1 U2372 ( .A(n3606), .ZN(n2281) );
  INV_X1 U2373 ( .A(IR_REG_1__SCAN_IN), .ZN(n2133) );
  NAND2_X1 U2374 ( .A1(n4019), .A2(n2792), .ZN(n2793) );
  NOR2_X1 U2375 ( .A1(n3960), .A2(n2100), .ZN(n2099) );
  INV_X1 U2376 ( .A(n2099), .ZN(n2098) );
  AND2_X1 U2377 ( .A1(n4219), .A2(n2680), .ZN(n3951) );
  OR2_X1 U2378 ( .A1(n3476), .A2(n3829), .ZN(n4220) );
  NOR2_X1 U2379 ( .A1(n2264), .A2(n2175), .ZN(n2174) );
  NOR2_X1 U2380 ( .A1(n3435), .A2(n2267), .ZN(n2266) );
  INV_X1 U2381 ( .A(n2558), .ZN(n2267) );
  NAND2_X1 U2382 ( .A1(n3226), .A2(n3188), .ZN(n3930) );
  AND2_X1 U2383 ( .A1(n2091), .A2(n3923), .ZN(n2112) );
  INV_X1 U2384 ( .A(n3927), .ZN(n2115) );
  NAND2_X1 U2385 ( .A1(n3018), .A2(n2977), .ZN(n3920) );
  NAND2_X1 U2386 ( .A1(n4005), .A2(n2992), .ZN(n3918) );
  OR2_X1 U2387 ( .A1(n2393), .A2(n2936), .ZN(n2401) );
  NAND2_X1 U2388 ( .A1(n3688), .A2(n3703), .ZN(n2153) );
  AND2_X1 U2389 ( .A1(n2057), .A2(n3524), .ZN(n2150) );
  OR2_X1 U2390 ( .A1(n3168), .A2(n3282), .ZN(n3167) );
  NAND2_X1 U2391 ( .A1(n2162), .A2(n2164), .ZN(n3040) );
  INV_X1 U2392 ( .A(IR_REG_27__SCAN_IN), .ZN(n2338) );
  NOR2_X1 U2393 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2700)
         );
  NOR2_X1 U2394 ( .A1(IR_REG_21__SCAN_IN), .A2(IR_REG_22__SCAN_IN), .ZN(n2194)
         );
  AND4_X1 U2395 ( .A1(n2572), .A2(n2334), .A3(n2333), .A4(n2332), .ZN(n2335)
         );
  NOR2_X1 U2396 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_13__SCAN_IN), .ZN(n2334)
         );
  NOR2_X1 U2397 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2333)
         );
  NOR2_X1 U2398 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2332)
         );
  INV_X1 U2399 ( .A(IR_REG_6__SCAN_IN), .ZN(n2461) );
  NOR2_X1 U2400 ( .A1(IR_REG_3__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2321)
         );
  INV_X1 U2401 ( .A(IR_REG_2__SCAN_IN), .ZN(n2330) );
  INV_X1 U2402 ( .A(n3183), .ZN(n2223) );
  OR2_X1 U2403 ( .A1(n3514), .A2(n3513), .ZN(n2306) );
  NAND2_X1 U2404 ( .A1(n3514), .A2(n3513), .ZN(n2305) );
  NAND2_X1 U2405 ( .A1(n2289), .A2(n2288), .ZN(n2287) );
  AOI21_X1 U2406 ( .B1(n2284), .B2(n2285), .A(n3687), .ZN(n2283) );
  INV_X1 U2407 ( .A(n2287), .ZN(n2284) );
  AOI22_X1 U2408 ( .A1(n3189), .A2(n2817), .B1(n3649), .B2(n3150), .ZN(n2866)
         );
  OR2_X1 U2409 ( .A1(n2393), .A2(n2392), .ZN(n2395) );
  NOR2_X1 U2410 ( .A1(n3108), .A2(n3107), .ZN(n3112) );
  NOR2_X1 U2411 ( .A1(n3106), .A2(n3105), .ZN(n3107) );
  NOR2_X1 U2412 ( .A1(n3112), .A2(n3111), .ZN(n3124) );
  INV_X1 U2413 ( .A(REG3_REG_17__SCAN_IN), .ZN(n4573) );
  AOI21_X1 U2414 ( .B1(n2200), .B2(n2201), .A(n2070), .ZN(n2196) );
  INV_X1 U2415 ( .A(n3012), .ZN(n2198) );
  INV_X1 U2416 ( .A(n3013), .ZN(n2199) );
  NAND2_X1 U2417 ( .A1(n2960), .A2(n2817), .ZN(n2816) );
  NAND2_X1 U2418 ( .A1(n2213), .A2(n2215), .ZN(n2212) );
  NAND2_X1 U2419 ( .A1(n2290), .A2(n2291), .ZN(n3442) );
  AOI21_X1 U2420 ( .B1(n2293), .B2(n3280), .A(n2079), .ZN(n2291) );
  OAI22_X1 U2421 ( .A1(n3004), .A2(n3645), .B1(n3657), .B2(n3157), .ZN(n2865)
         );
  NAND2_X1 U2422 ( .A1(n2088), .A2(n3730), .ZN(n2232) );
  AND3_X1 U2423 ( .A1(n2925), .A2(n2853), .A3(n2923), .ZN(n2884) );
  OR2_X1 U2424 ( .A1(n3645), .A2(n2861), .ZN(n2882) );
  OAI22_X1 U2425 ( .A1(n2891), .A2(n2388), .B1(n2393), .B2(n2780), .ZN(n2323)
         );
  NAND2_X1 U2426 ( .A1(n2131), .A2(n2133), .ZN(n2180) );
  NAND2_X1 U2427 ( .A1(n2132), .A2(IR_REG_0__SCAN_IN), .ZN(n2181) );
  NAND2_X1 U2428 ( .A1(n2133), .A2(IR_REG_31__SCAN_IN), .ZN(n2132) );
  NAND2_X1 U2429 ( .A1(n4011), .A2(n2788), .ZN(n2838) );
  XNOR2_X1 U2430 ( .A(n2893), .B(n2185), .ZN(n2806) );
  NOR2_X1 U2431 ( .A1(n2899), .A2(n2238), .ZN(n2237) );
  OR2_X1 U2432 ( .A1(n2239), .A2(n2899), .ZN(n2236) );
  NOR2_X1 U2433 ( .A1(n2804), .A2(n2186), .ZN(n2893) );
  NOR2_X1 U2434 ( .A1(n2801), .A2(n2187), .ZN(n2186) );
  INV_X1 U2435 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2187) );
  NOR2_X1 U2436 ( .A1(n2806), .A2(n2805), .ZN(n2894) );
  NAND2_X1 U2437 ( .A1(n4418), .A2(n4058), .ZN(n4060) );
  NAND2_X1 U2438 ( .A1(n4421), .A2(n4033), .ZN(n4034) );
  NAND2_X1 U2439 ( .A1(n4430), .A2(REG2_REG_12__SCAN_IN), .ZN(n4429) );
  NAND2_X1 U2440 ( .A1(n4446), .A2(n4062), .ZN(n4064) );
  OR2_X1 U2441 ( .A1(n4451), .A2(n4037), .ZN(n2119) );
  NAND2_X1 U2442 ( .A1(n4469), .A2(n4040), .ZN(n4478) );
  AOI21_X1 U2443 ( .B1(n4128), .B2(n3861), .A(n3862), .ZN(n4111) );
  AOI21_X1 U2444 ( .B1(n2156), .B2(n2155), .A(n2154), .ZN(n4128) );
  AND2_X1 U2445 ( .A1(n3988), .A2(n4146), .ZN(n2154) );
  NAND2_X1 U2446 ( .A1(n4285), .A2(n4152), .ZN(n2155) );
  INV_X1 U2447 ( .A(n4140), .ZN(n2156) );
  NAND2_X1 U2448 ( .A1(n2685), .A2(n2684), .ZN(n2102) );
  NAND2_X1 U2449 ( .A1(n3551), .A2(n2081), .ZN(n2248) );
  INV_X1 U2450 ( .A(n4211), .ZN(n4201) );
  NOR2_X1 U2451 ( .A1(n4208), .A2(n2250), .ZN(n2249) );
  INV_X1 U2452 ( .A(n2252), .ZN(n2250) );
  NOR2_X1 U2453 ( .A1(n2577), .A2(n4573), .ZN(n2597) );
  INV_X1 U2454 ( .A(n3778), .ZN(n3597) );
  NAND2_X1 U2455 ( .A1(n2176), .A2(n2174), .ZN(n3472) );
  AND2_X1 U2456 ( .A1(n3950), .A2(n3822), .ZN(n3435) );
  OAI21_X1 U2457 ( .B1(n2674), .B2(n2105), .A(n2103), .ZN(n3434) );
  INV_X1 U2458 ( .A(n2104), .ZN(n2103) );
  OAI21_X1 U2459 ( .B1(n2056), .B2(n2105), .A(n3435), .ZN(n2104) );
  INV_X1 U2460 ( .A(n3827), .ZN(n2105) );
  NAND2_X1 U2461 ( .A1(n2559), .A2(n2266), .ZN(n2324) );
  NAND2_X1 U2462 ( .A1(n2674), .A2(n2056), .ZN(n3357) );
  AND2_X1 U2463 ( .A1(n2514), .A2(n2258), .ZN(n2254) );
  AND2_X1 U2464 ( .A1(n3299), .A2(n3301), .ZN(n3897) );
  NAND2_X1 U2465 ( .A1(n2116), .A2(n3931), .ZN(n3139) );
  NAND2_X1 U2466 ( .A1(n3232), .A2(n3935), .ZN(n2116) );
  OAI21_X1 U2467 ( .B1(n2260), .B2(n2466), .A(n2477), .ZN(n2259) );
  NAND2_X1 U2468 ( .A1(n2160), .A2(n2162), .ZN(n2159) );
  INV_X1 U2469 ( .A(n2164), .ZN(n2163) );
  AND2_X1 U2470 ( .A1(n2432), .A2(REG3_REG_6__SCAN_IN), .ZN(n2458) );
  AND2_X1 U2471 ( .A1(n3932), .A2(n3930), .ZN(n3896) );
  AOI21_X1 U2472 ( .B1(n3058), .B2(n2428), .A(n2430), .ZN(n3024) );
  NAND2_X1 U2473 ( .A1(n2298), .A2(IR_REG_31__SCAN_IN), .ZN(n2648) );
  AND2_X1 U2474 ( .A1(n2301), .A2(n2300), .ZN(n2299) );
  INV_X1 U2475 ( .A(IR_REG_18__SCAN_IN), .ZN(n2300) );
  INV_X1 U2476 ( .A(IR_REG_19__SCAN_IN), .ZN(n2647) );
  NAND2_X1 U2477 ( .A1(n3000), .A2(n3150), .ZN(n3912) );
  INV_X1 U2478 ( .A(n3150), .ZN(n3001) );
  AND2_X1 U2479 ( .A1(n2697), .A2(n2875), .ZN(n2998) );
  AND2_X1 U2480 ( .A1(n2658), .A2(n2998), .ZN(n2811) );
  AND3_X1 U2481 ( .A1(n2729), .A2(n2728), .A3(n2852), .ZN(n2743) );
  NAND2_X1 U2482 ( .A1(n2712), .A2(n4382), .ZN(n2761) );
  NOR2_X1 U2483 ( .A1(n2703), .A2(IR_REG_26__SCAN_IN), .ZN(n2140) );
  INV_X1 U2484 ( .A(IR_REG_23__SCAN_IN), .ZN(n2716) );
  NAND2_X1 U2485 ( .A1(n2575), .A2(n2301), .ZN(n2604) );
  NAND2_X1 U2486 ( .A1(n2575), .A2(n2574), .ZN(n2593) );
  AND2_X1 U2487 ( .A1(n2569), .A2(n2554), .ZN(n4044) );
  INV_X1 U2488 ( .A(IR_REG_7__SCAN_IN), .ZN(n2463) );
  INV_X1 U2489 ( .A(IR_REG_3__SCAN_IN), .ZN(n2406) );
  OR2_X1 U2490 ( .A1(n2329), .A2(n2630), .ZN(n4114) );
  NAND2_X1 U2491 ( .A1(n2295), .A2(n2292), .ZN(n3287) );
  INV_X1 U2492 ( .A(n2294), .ZN(n2292) );
  AOI21_X1 U2493 ( .B1(n2272), .B2(n2278), .A(n2086), .ZN(n2271) );
  NAND2_X1 U2494 ( .A1(n2427), .A2(n4393), .ZN(n2143) );
  INV_X1 U2495 ( .A(DATAI_1_), .ZN(n2144) );
  AND2_X1 U2496 ( .A1(n2622), .A2(n2621), .ZN(n4132) );
  OAI211_X1 U2497 ( .C1(n2402), .C2(n4376), .A(n2603), .B(n2602), .ZN(n4223)
         );
  NOR2_X1 U2498 ( .A1(n2785), .A2(n2784), .ZN(n2802) );
  AND2_X1 U2499 ( .A1(n2189), .A2(n2188), .ZN(n2804) );
  INV_X1 U2500 ( .A(n2794), .ZN(n2188) );
  XNOR2_X1 U2501 ( .A(n2121), .B(n2185), .ZN(n2898) );
  NAND2_X1 U2502 ( .A1(n4419), .A2(n4420), .ZN(n4418) );
  XNOR2_X1 U2503 ( .A(n4060), .B(n4531), .ZN(n4435) );
  NAND2_X1 U2504 ( .A1(n4447), .A2(n4448), .ZN(n4446) );
  XNOR2_X1 U2505 ( .A(n4064), .B(n2120), .ZN(n4456) );
  NOR2_X1 U2506 ( .A1(n4452), .A2(n2534), .ZN(n4451) );
  NOR2_X1 U2507 ( .A1(n4474), .A2(n4068), .ZN(n4484) );
  OAI21_X1 U2508 ( .B1(n4490), .B2(n2242), .A(n2241), .ZN(n2240) );
  AOI21_X1 U2509 ( .B1(n4493), .B2(ADDR_REG_18__SCAN_IN), .A(n4492), .ZN(n2241) );
  AND2_X1 U2510 ( .A1(n4479), .A2(n2136), .ZN(n4490) );
  NAND2_X1 U2511 ( .A1(n2243), .A2(n4440), .ZN(n2242) );
  AND2_X1 U2512 ( .A1(n2796), .A2(n2783), .ZN(n4495) );
  INV_X1 U2513 ( .A(n3997), .ZN(n3290) );
  INV_X1 U2514 ( .A(n4195), .ZN(n4513) );
  NAND3_X1 U2515 ( .A1(n2148), .A2(n2147), .A3(n2146), .ZN(n4395) );
  NAND2_X1 U2516 ( .A1(n3853), .A2(n2736), .ZN(n2146) );
  OR2_X1 U2517 ( .A1(n4094), .A2(n4245), .ZN(n2147) );
  NOR2_X1 U2518 ( .A1(n2169), .A2(IR_REG_29__SCAN_IN), .ZN(n2167) );
  INV_X1 U2519 ( .A(n4043), .ZN(n4522) );
  INV_X1 U2520 ( .A(n2325), .ZN(n2307) );
  INV_X1 U2521 ( .A(n2305), .ZN(n2303) );
  AND2_X1 U2522 ( .A1(n2306), .A2(n2215), .ZN(n2207) );
  NOR2_X1 U2523 ( .A1(n2211), .A2(n2208), .ZN(n2205) );
  INV_X1 U2524 ( .A(n3658), .ZN(n3652) );
  INV_X1 U2525 ( .A(n2313), .ZN(n2311) );
  INV_X1 U2526 ( .A(n3630), .ZN(n2310) );
  INV_X1 U2527 ( .A(n3623), .ZN(n2312) );
  NAND2_X1 U2528 ( .A1(n2216), .A2(n3490), .ZN(n2213) );
  INV_X1 U2529 ( .A(n3489), .ZN(n2215) );
  INV_X1 U2530 ( .A(n3391), .ZN(n3392) );
  NOR2_X1 U2531 ( .A1(n3865), .A2(n3834), .ZN(n2101) );
  INV_X1 U2532 ( .A(n2605), .ZN(n2172) );
  AND2_X1 U2533 ( .A1(n2419), .A2(REG3_REG_5__SCAN_IN), .ZN(n2432) );
  AND2_X1 U2534 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2419) );
  INV_X1 U2535 ( .A(n2761), .ZN(n2730) );
  NAND2_X1 U2536 ( .A1(n4090), .A2(n3846), .ZN(n2110) );
  NAND2_X1 U2537 ( .A1(n3157), .A2(n3001), .ZN(n2991) );
  INV_X1 U2538 ( .A(IR_REG_26__SCAN_IN), .ZN(n2269) );
  AND3_X1 U2539 ( .A1(n2700), .A2(n2336), .A3(n2655), .ZN(n2337) );
  NOR2_X1 U2540 ( .A1(IR_REG_22__SCAN_IN), .A2(IR_REG_25__SCAN_IN), .ZN(n2336)
         );
  INV_X1 U2541 ( .A(IR_REG_17__SCAN_IN), .ZN(n2302) );
  INV_X1 U2542 ( .A(IR_REG_15__SCAN_IN), .ZN(n2552) );
  INV_X1 U2543 ( .A(IR_REG_13__SCAN_IN), .ZN(n2541) );
  INV_X1 U2544 ( .A(IR_REG_11__SCAN_IN), .ZN(n2511) );
  OR3_X1 U2545 ( .A1(n2486), .A2(IR_REG_8__SCAN_IN), .A3(IR_REG_7__SCAN_IN), 
        .ZN(n2498) );
  NAND2_X1 U2546 ( .A1(n3711), .A2(n2277), .ZN(n2276) );
  INV_X1 U2547 ( .A(n3710), .ZN(n2277) );
  NOR2_X1 U2548 ( .A1(n3766), .A2(n2314), .ZN(n2313) );
  INV_X1 U2549 ( .A(n3698), .ZN(n2314) );
  NOR2_X1 U2550 ( .A1(n3279), .A2(n3278), .ZN(n2294) );
  NAND2_X1 U2551 ( .A1(n2297), .A2(n2296), .ZN(n2295) );
  INV_X1 U2552 ( .A(n3281), .ZN(n2297) );
  INV_X1 U2553 ( .A(n3789), .ZN(n2279) );
  INV_X1 U2554 ( .A(n2219), .ZN(n2217) );
  INV_X1 U2555 ( .A(REG3_REG_12__SCAN_IN), .ZN(n4724) );
  INV_X1 U2556 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4596) );
  NAND2_X1 U2557 ( .A1(n3676), .A2(n3628), .ZN(n3742) );
  INV_X1 U2558 ( .A(n3016), .ZN(n2195) );
  AOI21_X1 U2559 ( .B1(n3251), .B2(n3250), .A(n3249), .ZN(n3281) );
  NAND2_X1 U2560 ( .A1(n2819), .A2(n2818), .ZN(n2867) );
  NOR2_X1 U2561 ( .A1(n2229), .A2(n2227), .ZN(n2226) );
  AND2_X1 U2562 ( .A1(n2283), .A2(n2230), .ZN(n2229) );
  NOR2_X1 U2563 ( .A1(n2516), .A2(n4724), .ZN(n2527) );
  AND2_X1 U2564 ( .A1(n2527), .A2(REG3_REG_13__SCAN_IN), .ZN(n2535) );
  NAND2_X1 U2565 ( .A1(n2535), .A2(REG3_REG_14__SCAN_IN), .ZN(n2563) );
  INV_X1 U2566 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2562) );
  NAND2_X1 U2567 ( .A1(n2128), .A2(n2184), .ZN(n2127) );
  INV_X1 U2568 ( .A(n2180), .ZN(n2128) );
  NAND2_X1 U2569 ( .A1(n2183), .A2(n2126), .ZN(n2125) );
  AND2_X1 U2570 ( .A1(REG2_REG_1__SCAN_IN), .A2(n2184), .ZN(n2126) );
  NAND2_X1 U2571 ( .A1(n2837), .A2(n2789), .ZN(n2791) );
  AND2_X1 U2572 ( .A1(n2827), .A2(REG1_REG_4__SCAN_IN), .ZN(n2825) );
  OR2_X1 U2573 ( .A1(n2825), .A2(n2190), .ZN(n2189) );
  AND2_X1 U2574 ( .A1(n2793), .A2(n4390), .ZN(n2190) );
  NAND2_X1 U2575 ( .A1(n4409), .A2(n4032), .ZN(n4422) );
  NAND2_X1 U2576 ( .A1(n4463), .A2(n4066), .ZN(n4067) );
  XNOR2_X1 U2577 ( .A(n4039), .B(n4524), .ZN(n4470) );
  INV_X1 U2578 ( .A(n4483), .ZN(n2193) );
  NAND2_X1 U2579 ( .A1(n2244), .A2(n4491), .ZN(n2243) );
  NAND2_X1 U2580 ( .A1(n4479), .A2(n2245), .ZN(n2244) );
  INV_X1 U2581 ( .A(n4480), .ZN(n2135) );
  OR2_X1 U2582 ( .A1(n4108), .A2(n3837), .ZN(n4090) );
  NAND2_X1 U2583 ( .A1(n2097), .A2(n2065), .ZN(n4106) );
  OR2_X1 U2584 ( .A1(n2685), .A2(n2098), .ZN(n2097) );
  NAND2_X1 U2585 ( .A1(n2099), .A2(n3836), .ZN(n2096) );
  NAND2_X1 U2586 ( .A1(n2102), .A2(n2101), .ZN(n4142) );
  NAND2_X1 U2587 ( .A1(n4189), .A2(n4168), .ZN(n2157) );
  AND2_X1 U2588 ( .A1(n2374), .A2(n2373), .ZN(n4204) );
  NAND2_X1 U2589 ( .A1(n2253), .A2(n3703), .ZN(n2252) );
  AND2_X1 U2590 ( .A1(n4181), .A2(n2682), .ZN(n4208) );
  OR2_X1 U2591 ( .A1(n2617), .A2(n2616), .ZN(n2251) );
  INV_X1 U2592 ( .A(n3551), .ZN(n2617) );
  NAND2_X1 U2593 ( .A1(n2681), .A2(n3831), .ZN(n4178) );
  AND2_X1 U2594 ( .A1(REG3_REG_19__SCAN_IN), .A2(REG3_REG_18__SCAN_IN), .ZN(
        n2327) );
  INV_X1 U2595 ( .A(n2585), .ZN(n2265) );
  NAND2_X1 U2596 ( .A1(n3434), .A2(n3822), .ZN(n3476) );
  OR2_X1 U2597 ( .A1(n2502), .A2(n2501), .ZN(n2516) );
  OAI21_X1 U2598 ( .B1(n3139), .B2(n3138), .A(n3936), .ZN(n3165) );
  OR2_X1 U2599 ( .A1(n3034), .A2(n2666), .ZN(n2667) );
  OAI21_X1 U2600 ( .B1(n2113), .B2(n2114), .A(n2111), .ZN(n3071) );
  INV_X1 U2601 ( .A(n2091), .ZN(n2113) );
  NOR2_X1 U2602 ( .A1(n2115), .A2(n2066), .ZN(n2114) );
  NAND2_X1 U2603 ( .A1(n4003), .A2(n3056), .ZN(n3923) );
  INV_X1 U2604 ( .A(n2811), .ZN(n3481) );
  INV_X1 U2605 ( .A(n3894), .ZN(n2661) );
  AND2_X1 U2606 ( .A1(n3920), .A2(n3917), .ZN(n3893) );
  OAI21_X1 U2607 ( .B1(n2659), .B2(n3912), .A(n2660), .ZN(n2983) );
  NAND2_X1 U2608 ( .A1(n3894), .A2(n2983), .ZN(n2982) );
  AND2_X1 U2609 ( .A1(n3918), .A2(n2662), .ZN(n3894) );
  NOR2_X1 U2610 ( .A1(n2117), .A2(n2059), .ZN(n3018) );
  OR2_X1 U2611 ( .A1(n2388), .A2(REG3_REG_3__SCAN_IN), .ZN(n2404) );
  INV_X1 U2612 ( .A(n3149), .ZN(n3157) );
  NOR2_X1 U2613 ( .A1(n3853), .A2(n2736), .ZN(n2149) );
  AOI21_X1 U2614 ( .B1(n2108), .B2(n4231), .A(n2107), .ZN(n3562) );
  AND2_X1 U2615 ( .A1(n4084), .A2(n3986), .ZN(n2107) );
  XNOR2_X1 U2616 ( .A(n2109), .B(n3883), .ZN(n2108) );
  NAND2_X1 U2617 ( .A1(n2110), .A2(n2639), .ZN(n2109) );
  OR2_X1 U2618 ( .A1(n4130), .A2(n4260), .ZN(n4112) );
  NOR2_X1 U2619 ( .A1(n2427), .A2(n2353), .ZN(n4260) );
  OR2_X1 U2620 ( .A1(n4151), .A2(n4269), .ZN(n4130) );
  INV_X1 U2621 ( .A(n4134), .ZN(n4269) );
  NAND2_X1 U2622 ( .A1(n4162), .A2(n4152), .ZN(n4151) );
  AND2_X1 U2623 ( .A1(n4191), .A2(n4168), .ZN(n4162) );
  NOR2_X1 U2624 ( .A1(n2427), .A2(n4684), .ZN(n4190) );
  OR2_X1 U2625 ( .A1(n4235), .A2(n4201), .ZN(n2152) );
  NOR3_X1 U2626 ( .A1(n3543), .A2(n4235), .A3(n3599), .ZN(n4234) );
  OR2_X1 U2627 ( .A1(n3482), .A2(n3597), .ZN(n3543) );
  NAND2_X1 U2628 ( .A1(n3316), .A2(n2082), .ZN(n3428) );
  NAND2_X1 U2629 ( .A1(n3316), .A2(n2150), .ZN(n3362) );
  NAND2_X1 U2630 ( .A1(n3316), .A2(n2057), .ZN(n3346) );
  INV_X1 U2631 ( .A(n3492), .ZN(n3497) );
  AND2_X1 U2632 ( .A1(n3316), .A2(n3454), .ZN(n3318) );
  INV_X1 U2633 ( .A(n3395), .ZN(n3399) );
  NOR2_X1 U2634 ( .A1(n3075), .A2(n3188), .ZN(n3239) );
  AND2_X1 U2635 ( .A1(n3239), .A2(n3238), .ZN(n3241) );
  NAND2_X1 U2636 ( .A1(n2263), .A2(n2262), .ZN(n4555) );
  INV_X1 U2637 ( .A(n3896), .ZN(n2262) );
  AND2_X1 U2638 ( .A1(n4227), .A2(n4540), .ZN(n4551) );
  NAND2_X1 U2639 ( .A1(n2145), .A2(n3131), .ZN(n3075) );
  INV_X1 U2640 ( .A(n3077), .ZN(n2145) );
  NOR2_X1 U2641 ( .A1(n3050), .A2(n3051), .ZN(n3049) );
  NAND2_X1 U2642 ( .A1(n3049), .A2(n3114), .ZN(n3077) );
  AND2_X1 U2643 ( .A1(n2753), .A2(n2998), .ZN(n4324) );
  INV_X1 U2644 ( .A(n4304), .ZN(n4325) );
  NOR2_X1 U2645 ( .A1(n2984), .A2(n2991), .ZN(n2993) );
  INV_X1 U2646 ( .A(n2853), .ZN(n2926) );
  AND2_X1 U2647 ( .A1(n2321), .A2(n2170), .ZN(n2166) );
  NOR2_X1 U2648 ( .A1(n2140), .A2(n2087), .ZN(n2691) );
  NAND2_X1 U2649 ( .A1(n2349), .A2(n2350), .ZN(n2692) );
  NAND2_X1 U2650 ( .A1(n2704), .A2(n2703), .ZN(n2713) );
  MUX2_X1 U2651 ( .A(IR_REG_31__SCAN_IN), .B(n2702), .S(IR_REG_25__SCAN_IN), 
        .Z(n2704) );
  XNOR2_X1 U2652 ( .A(n2715), .B(n2716), .ZN(n2769) );
  INV_X1 U2653 ( .A(IR_REG_20__SCAN_IN), .ZN(n2650) );
  INV_X1 U2654 ( .A(n3998), .ZN(n3257) );
  OAI21_X1 U2655 ( .B1(n3186), .B2(n2224), .A(n2220), .ZN(n3213) );
  NAND2_X1 U2656 ( .A1(n2304), .A2(n2305), .ZN(n3570) );
  NAND2_X1 U2657 ( .A1(n2295), .A2(n2293), .ZN(n3393) );
  NAND2_X1 U2658 ( .A1(n3773), .A2(n2287), .ZN(n2282) );
  OAI21_X1 U2659 ( .B1(n3773), .B2(n2286), .A(n2283), .ZN(n3685) );
  AND4_X1 U2660 ( .A1(n2397), .A2(n2396), .A3(n2395), .A4(n2394), .ZN(n2967)
         );
  OR2_X1 U2661 ( .A1(n2388), .A2(n2836), .ZN(n2396) );
  INV_X1 U2662 ( .A(n3995), .ZN(n3455) );
  AND2_X1 U2663 ( .A1(n2214), .A2(n2216), .ZN(n3491) );
  NAND2_X1 U2664 ( .A1(n3445), .A2(n3444), .ZN(n2214) );
  AND2_X1 U2665 ( .A1(n2424), .A2(n2423), .ZN(n3117) );
  NOR2_X1 U2666 ( .A1(n2418), .A2(n2417), .ZN(n2424) );
  NAND2_X1 U2667 ( .A1(n2884), .A2(n2880), .ZN(n3808) );
  INV_X1 U2668 ( .A(n2387), .ZN(n3004) );
  NAND2_X1 U2669 ( .A1(n2068), .A2(n2141), .ZN(n3150) );
  NAND2_X1 U2670 ( .A1(n2427), .A2(IR_REG_0__SCAN_IN), .ZN(n2141) );
  INV_X1 U2671 ( .A(DATAI_0_), .ZN(n2142) );
  NAND2_X1 U2672 ( .A1(n2315), .A2(n3698), .ZN(n3765) );
  NAND2_X1 U2673 ( .A1(n2908), .A2(n2910), .ZN(n2911) );
  INV_X1 U2674 ( .A(n2909), .ZN(n2910) );
  INV_X1 U2675 ( .A(n2984), .ZN(n2992) );
  AND3_X1 U2676 ( .A1(n2459), .A2(n2460), .A3(n2165), .ZN(n3226) );
  NOR2_X1 U2677 ( .A1(n2054), .A2(n2060), .ZN(n2165) );
  NAND2_X1 U2678 ( .A1(n2884), .A2(n2871), .ZN(n3800) );
  NAND2_X1 U2679 ( .A1(n2973), .A2(n2972), .ZN(n3793) );
  NAND2_X1 U2680 ( .A1(n2273), .A2(n3711), .ZN(n3791) );
  INV_X1 U2681 ( .A(n3800), .ZN(n3806) );
  INV_X1 U2682 ( .A(n3793), .ZN(n3819) );
  OAI21_X1 U2683 ( .B1(n4114), .B2(n2388), .A(n2348), .ZN(n4270) );
  NAND2_X1 U2684 ( .A1(n2628), .A2(n2627), .ZN(n4261) );
  NAND2_X1 U2685 ( .A1(n2359), .A2(n2358), .ZN(n3988) );
  INV_X1 U2686 ( .A(n4204), .ZN(n4282) );
  OAI21_X1 U2687 ( .B1(n4212), .B2(n2388), .A(n2380), .ZN(n4186) );
  OAI211_X1 U2688 ( .C1(n4232), .C2(n2388), .A(n2609), .B(n2608), .ZN(n4301)
         );
  INV_X1 U2689 ( .A(n3226), .ZN(n3999) );
  CLKBUF_X1 U2690 ( .A(U4043), .Z(n4000) );
  INV_X1 U2691 ( .A(n3117), .ZN(n4003) );
  INV_X1 U2692 ( .A(n3018), .ZN(n4004) );
  INV_X1 U2693 ( .A(n2967), .ZN(n4005) );
  INV_X1 U2694 ( .A(n2323), .ZN(n2322) );
  NAND2_X1 U2695 ( .A1(n2247), .A2(n2246), .ZN(n4008) );
  NOR2_X1 U2696 ( .A1(n2131), .A2(n2780), .ZN(n2246) );
  NAND2_X1 U2697 ( .A1(n2130), .A2(n2125), .ZN(n2247) );
  OAI211_X1 U2698 ( .C1(n2181), .C2(n2129), .A(n2779), .B(n2127), .ZN(n2130)
         );
  NAND3_X1 U2699 ( .A1(n2179), .A2(n2182), .A3(n2178), .ZN(n4013) );
  NAND2_X1 U2700 ( .A1(n2129), .A2(n2787), .ZN(n2182) );
  NAND2_X1 U2701 ( .A1(n2183), .A2(n2062), .ZN(n2179) );
  NAND2_X1 U2702 ( .A1(n4013), .A2(n4012), .ZN(n4011) );
  XNOR2_X1 U2703 ( .A(n2791), .B(n2790), .ZN(n4020) );
  AND2_X1 U2704 ( .A1(n2124), .A2(n2123), .ZN(n2785) );
  NAND2_X1 U2705 ( .A1(n2824), .A2(REG2_REG_4__SCAN_IN), .ZN(n2124) );
  INV_X1 U2706 ( .A(n2189), .ZN(n2795) );
  AND2_X1 U2707 ( .A1(n2235), .A2(n2239), .ZN(n2900) );
  NAND2_X1 U2708 ( .A1(n2898), .A2(REG2_REG_6__SCAN_IN), .ZN(n2235) );
  AOI21_X1 U2709 ( .B1(n4388), .B2(n2895), .A(n2894), .ZN(n2949) );
  NAND2_X1 U2710 ( .A1(n4414), .A2(n4057), .ZN(n4419) );
  NAND2_X1 U2711 ( .A1(n4434), .A2(n4061), .ZN(n4447) );
  NAND2_X1 U2712 ( .A1(n4429), .A2(n4035), .ZN(n4442) );
  XNOR2_X1 U2713 ( .A(n4036), .B(n2120), .ZN(n4452) );
  NAND2_X1 U2714 ( .A1(n4455), .A2(n4065), .ZN(n4464) );
  NAND2_X1 U2715 ( .A1(n4464), .A2(n4465), .ZN(n4463) );
  INV_X1 U2716 ( .A(n4459), .ZN(n2118) );
  INV_X1 U2717 ( .A(n2119), .ZN(n4460) );
  XNOR2_X1 U2718 ( .A(n4067), .B(n4524), .ZN(n4473) );
  OAI21_X1 U2719 ( .B1(n4478), .B2(n2137), .A(n2134), .ZN(n2138) );
  AOI21_X1 U2720 ( .B1(n2136), .B2(n2135), .A(n2139), .ZN(n2134) );
  AND2_X1 U2721 ( .A1(n2637), .A2(n2636), .ZN(n4264) );
  NAND2_X1 U2722 ( .A1(n2102), .A2(n3867), .ZN(n4158) );
  NAND2_X1 U2723 ( .A1(n2248), .A2(n2052), .ZN(n4176) );
  NAND2_X1 U2724 ( .A1(n3472), .A2(n2596), .ZN(n3532) );
  NAND2_X1 U2725 ( .A1(n2324), .A2(n2571), .ZN(n3463) );
  NAND2_X1 U2726 ( .A1(n3357), .A2(n3827), .ZN(n3436) );
  INV_X1 U2727 ( .A(n3991), .ZN(n4329) );
  NAND2_X1 U2728 ( .A1(n2674), .A2(n3820), .ZN(n3356) );
  INV_X1 U2729 ( .A(n3992), .ZN(n3809) );
  NAND2_X1 U2730 ( .A1(n2255), .A2(n2258), .ZN(n3267) );
  NAND2_X1 U2731 ( .A1(n2490), .A2(n2489), .ZN(n3166) );
  INV_X1 U2732 ( .A(n2259), .ZN(n2161) );
  INV_X1 U2733 ( .A(n3561), .ZN(n4167) );
  INV_X1 U2734 ( .A(n4198), .ZN(n4209) );
  XNOR2_X1 U2735 ( .A(n2648), .B(n2647), .ZN(n4078) );
  INV_X1 U2736 ( .A(n4500), .ZN(n4511) );
  AND2_X2 U2737 ( .A1(n2743), .A2(n2853), .ZN(n4568) );
  NOR2_X1 U2738 ( .A1(n4244), .A2(n4245), .ZN(n4243) );
  AND2_X2 U2739 ( .A1(n2743), .A2(n2926), .ZN(n4559) );
  INV_X1 U2740 ( .A(n4521), .ZN(n2762) );
  NAND2_X1 U2741 ( .A1(n2761), .A2(n2876), .ZN(n4520) );
  NAND2_X1 U2742 ( .A1(n2339), .A2(IR_REG_31__SCAN_IN), .ZN(n2340) );
  INV_X1 U2743 ( .A(n2342), .ZN(n2755) );
  AND2_X1 U2744 ( .A1(n2711), .A2(n2710), .ZN(n4382) );
  INV_X1 U2745 ( .A(n2140), .ZN(n2710) );
  NAND2_X1 U2746 ( .A1(n2706), .A2(IR_REG_31__SCAN_IN), .ZN(n2707) );
  INV_X1 U2747 ( .A(DATAI_23_), .ZN(n4684) );
  AND2_X1 U2748 ( .A1(n2769), .A2(STATE_REG_SCAN_IN), .ZN(n4521) );
  XNOR2_X1 U2749 ( .A(n2656), .B(IR_REG_22__SCAN_IN), .ZN(n3981) );
  NAND2_X1 U2750 ( .A1(n2652), .A2(n2655), .ZN(n2699) );
  XNOR2_X1 U2751 ( .A(n2654), .B(IR_REG_21__SCAN_IN), .ZN(n4384) );
  INV_X1 U2752 ( .A(n4078), .ZN(n4385) );
  AND2_X1 U2753 ( .A1(n2472), .A2(n2465), .ZN(n4387) );
  AND2_X1 U2754 ( .A1(n2425), .A2(n2408), .ZN(n4391) );
  NAND2_X1 U2755 ( .A1(n2183), .A2(n2184), .ZN(n4393) );
  NOR2_X1 U2756 ( .A1(n4484), .A2(n4483), .ZN(n4485) );
  INV_X1 U2757 ( .A(n2240), .ZN(n4498) );
  AOI21_X1 U2758 ( .B1(n4395), .B2(n4513), .A(n2092), .ZN(n4396) );
  INV_X1 U2759 ( .A(n2427), .ZN(n2640) );
  NAND2_X2 U2760 ( .A1(n2755), .A2(n2341), .ZN(n2388) );
  INV_X2 U2761 ( .A(n3657), .ZN(n3649) );
  OR2_X2 U2762 ( .A1(n2811), .A2(n3657), .ZN(n2907) );
  INV_X2 U2763 ( .A(n2907), .ZN(n2960) );
  OR3_X1 U2764 ( .A1(n3543), .A2(n2153), .A3(n2152), .ZN(n2050) );
  NAND2_X1 U2765 ( .A1(n2542), .A2(n2064), .ZN(n2703) );
  OR2_X1 U2766 ( .A1(n2169), .A2(n2268), .ZN(n2051) );
  NAND2_X1 U2767 ( .A1(n2320), .A2(n2321), .ZN(n2440) );
  OAI21_X1 U2768 ( .B1(n2265), .B2(n2571), .A(n2067), .ZN(n2264) );
  OR2_X1 U2769 ( .A1(n2249), .A2(n2076), .ZN(n2052) );
  OR2_X1 U2770 ( .A1(n2303), .A2(n2307), .ZN(n2053) );
  AND2_X1 U2771 ( .A1(n2580), .A2(REG0_REG_7__SCAN_IN), .ZN(n2054) );
  AND2_X1 U2772 ( .A1(n2052), .A2(n2085), .ZN(n2055) );
  INV_X1 U2773 ( .A(IR_REG_21__SCAN_IN), .ZN(n2655) );
  AND2_X1 U2774 ( .A1(n2343), .A2(n2342), .ZN(n2413) );
  NAND2_X1 U2775 ( .A1(n2559), .A2(n2080), .ZN(n2176) );
  OAI211_X1 U2776 ( .C1(n3709), .C2(n2388), .A(n2615), .B(n2614), .ZN(n4202)
         );
  AND2_X1 U2777 ( .A1(n2106), .A2(n3820), .ZN(n2056) );
  AND2_X1 U2778 ( .A1(n3454), .A2(n3497), .ZN(n2057) );
  AND2_X1 U2779 ( .A1(n2176), .A2(n2177), .ZN(n3471) );
  INV_X1 U2780 ( .A(n3280), .ZN(n2296) );
  NAND2_X1 U2781 ( .A1(n2279), .A2(n3711), .ZN(n2278) );
  NAND2_X1 U2782 ( .A1(n2366), .A2(n2365), .ZN(n4147) );
  INV_X1 U2783 ( .A(n4147), .ZN(n4189) );
  NOR2_X1 U2784 ( .A1(n3183), .A2(n3184), .ZN(n2224) );
  XNOR2_X1 U2785 ( .A(n2340), .B(IR_REG_30__SCAN_IN), .ZN(n2341) );
  AND2_X1 U2786 ( .A1(n2542), .A2(n2335), .ZN(n2652) );
  AOI21_X1 U2787 ( .B1(n4068), .B2(n2193), .A(n4071), .ZN(n2192) );
  NAND2_X1 U2788 ( .A1(n2658), .A2(n4384), .ZN(n2812) );
  AND2_X1 U2789 ( .A1(n2119), .A2(n2118), .ZN(n2058) );
  NAND2_X1 U2790 ( .A1(n2168), .A2(n2167), .ZN(n2339) );
  AND2_X1 U2791 ( .A1(n2414), .A2(REG1_REG_3__SCAN_IN), .ZN(n2059) );
  AND2_X1 U2792 ( .A1(n2414), .A2(REG1_REG_7__SCAN_IN), .ZN(n2060) );
  NAND2_X1 U2793 ( .A1(IR_REG_1__SCAN_IN), .A2(n2758), .ZN(n2184) );
  INV_X1 U2794 ( .A(n2184), .ZN(n2129) );
  AND2_X1 U2795 ( .A1(n3125), .A2(n3126), .ZN(n2061) );
  AND2_X1 U2796 ( .A1(n2184), .A2(REG1_REG_1__SCAN_IN), .ZN(n2062) );
  AND2_X1 U2797 ( .A1(n2282), .A2(n2285), .ZN(n2063) );
  AND2_X1 U2798 ( .A1(n2335), .A2(n2337), .ZN(n2064) );
  AND2_X1 U2799 ( .A1(n2687), .A2(n2096), .ZN(n2065) );
  AND2_X1 U2800 ( .A1(n2664), .A2(n3923), .ZN(n2066) );
  NAND2_X1 U2801 ( .A1(n4326), .A2(n3590), .ZN(n2067) );
  OR2_X1 U2802 ( .A1(n2427), .A2(n2142), .ZN(n2068) );
  OR2_X1 U2803 ( .A1(n2427), .A2(n2144), .ZN(n2069) );
  OR2_X1 U2804 ( .A1(n2802), .A2(n2122), .ZN(n2121) );
  INV_X1 U2805 ( .A(n2221), .ZN(n2220) );
  NOR2_X1 U2806 ( .A1(n2223), .A2(n3185), .ZN(n2221) );
  AND2_X1 U2807 ( .A1(n2199), .A2(n2198), .ZN(n2070) );
  INV_X1 U2808 ( .A(IR_REG_0__SCAN_IN), .ZN(n2131) );
  INV_X1 U2809 ( .A(n2224), .ZN(n2222) );
  AND2_X1 U2810 ( .A1(n2222), .A2(n3212), .ZN(n2071) );
  NOR2_X1 U2811 ( .A1(n3286), .A2(n2294), .ZN(n2293) );
  AND2_X1 U2812 ( .A1(n2192), .A2(n2191), .ZN(n2072) );
  AND2_X1 U2813 ( .A1(n2338), .A2(n2269), .ZN(n2073) );
  INV_X1 U2814 ( .A(n4388), .ZN(n2185) );
  INV_X1 U2815 ( .A(n2413), .ZN(n2402) );
  INV_X1 U2816 ( .A(n3774), .ZN(n2288) );
  OR2_X1 U2817 ( .A1(n3543), .A2(n3599), .ZN(n2074) );
  INV_X1 U2818 ( .A(n2286), .ZN(n2285) );
  NOR2_X1 U2819 ( .A1(n2289), .A2(n2288), .ZN(n2286) );
  NAND2_X1 U2820 ( .A1(n2251), .A2(n2249), .ZN(n2075) );
  XNOR2_X1 U2821 ( .A(n2707), .B(IR_REG_24__SCAN_IN), .ZN(n2714) );
  AND2_X1 U2822 ( .A1(n4186), .A2(n4201), .ZN(n2076) );
  INV_X1 U2823 ( .A(n3574), .ZN(n3810) );
  AND2_X1 U2824 ( .A1(n3730), .A2(n3718), .ZN(n2077) );
  NAND2_X1 U2825 ( .A1(n2228), .A2(n2232), .ZN(n3773) );
  OR2_X1 U2826 ( .A1(n4223), .A2(n3599), .ZN(n2078) );
  INV_X1 U2827 ( .A(n3996), .ZN(n3398) );
  INV_X1 U2828 ( .A(n2101), .ZN(n2100) );
  OAI22_X1 U2829 ( .A1(n3192), .A2(n2907), .B1(n3645), .B2(n3131), .ZN(n3184)
         );
  AND2_X1 U2830 ( .A1(n3390), .A2(n3392), .ZN(n2079) );
  INV_X1 U2831 ( .A(n2151), .ZN(n4210) );
  NOR3_X1 U2832 ( .A1(n3543), .A2(n2153), .A3(n4235), .ZN(n2151) );
  NAND2_X1 U2833 ( .A1(n2251), .A2(n2252), .ZN(n4207) );
  AND2_X1 U2834 ( .A1(n2266), .A2(n2585), .ZN(n2080) );
  NOR2_X1 U2835 ( .A1(n2076), .A2(n2616), .ZN(n2081) );
  AND2_X1 U2836 ( .A1(n2150), .A2(n3810), .ZN(n2082) );
  AND2_X1 U2837 ( .A1(n4282), .A2(n4190), .ZN(n2083) );
  AND2_X1 U2838 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_29__SCAN_IN), .ZN(n2084)
         );
  INV_X1 U2839 ( .A(n2275), .ZN(n2274) );
  OAI21_X1 U2840 ( .B1(n3789), .B2(n2276), .A(n3787), .ZN(n2275) );
  INV_X1 U2841 ( .A(n2211), .ZN(n2210) );
  NAND2_X1 U2842 ( .A1(n2215), .A2(n3444), .ZN(n2211) );
  NAND2_X1 U2843 ( .A1(n4204), .A2(n3679), .ZN(n2085) );
  NOR2_X1 U2844 ( .A1(n3656), .A2(n3655), .ZN(n2086) );
  NAND2_X1 U2845 ( .A1(IR_REG_27__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2087) );
  NAND2_X1 U2846 ( .A1(n3727), .A2(n3729), .ZN(n2088) );
  NOR2_X1 U2847 ( .A1(n3669), .A2(n2275), .ZN(n2272) );
  INV_X1 U2848 ( .A(IR_REG_31__SCAN_IN), .ZN(n2758) );
  NAND2_X1 U2849 ( .A1(n4387), .A2(REG2_REG_7__SCAN_IN), .ZN(n2089) );
  INV_X1 U2850 ( .A(IR_REG_28__SCAN_IN), .ZN(n2170) );
  OR2_X1 U2851 ( .A1(n2312), .A2(n3697), .ZN(n2090) );
  INV_X1 U2852 ( .A(n4235), .ZN(n3757) );
  INV_X1 U2853 ( .A(n2817), .ZN(n3000) );
  INV_X1 U2854 ( .A(n3477), .ZN(n2175) );
  NAND2_X1 U2855 ( .A1(n2400), .A2(n2661), .ZN(n2920) );
  NAND2_X1 U2856 ( .A1(n4002), .A2(n3114), .ZN(n2091) );
  AND2_X1 U2857 ( .A1(n4519), .A2(REG2_REG_30__SCAN_IN), .ZN(n2092) );
  AND2_X1 U2858 ( .A1(n3921), .A2(n3923), .ZN(n3053) );
  NAND2_X1 U2859 ( .A1(n4555), .A2(n2466), .ZN(n3231) );
  AOI21_X1 U2860 ( .B1(n2218), .B2(n2071), .A(n2217), .ZN(n3251) );
  NOR2_X1 U2861 ( .A1(n2964), .A2(n2201), .ZN(n2093) );
  INV_X1 U2862 ( .A(n3490), .ZN(n2203) );
  INV_X1 U2863 ( .A(n3892), .ZN(n2106) );
  AND2_X1 U2864 ( .A1(n2559), .A2(n2558), .ZN(n2094) );
  NAND2_X1 U2865 ( .A1(n2640), .A2(DATAI_21_), .ZN(n3703) );
  NAND2_X1 U2866 ( .A1(n2705), .A2(IR_REG_31__SCAN_IN), .ZN(n2715) );
  INV_X1 U2867 ( .A(n3697), .ZN(n2308) );
  INV_X1 U2868 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2238) );
  INV_X1 U2869 ( .A(n2264), .ZN(n2177) );
  INV_X1 U2870 ( .A(n4063), .ZN(n2120) );
  NAND2_X1 U2871 ( .A1(n2168), .A2(n2542), .ZN(n2349) );
  INV_X1 U2872 ( .A(n4440), .ZN(n4489) );
  AND2_X1 U2873 ( .A1(n2796), .A2(n3978), .ZN(n4440) );
  NAND2_X1 U2874 ( .A1(n2640), .A2(DATAI_24_), .ZN(n4168) );
  INV_X1 U2875 ( .A(n2137), .ZN(n2136) );
  OR2_X1 U2876 ( .A1(n4491), .A2(n4027), .ZN(n2137) );
  OR2_X1 U2877 ( .A1(n4070), .A2(REG2_REG_17__SCAN_IN), .ZN(n2245) );
  NOR2_X2 U2878 ( .A1(n2968), .A2(n2762), .ZN(U4043) );
  NAND2_X1 U2879 ( .A1(n3054), .A2(n2112), .ZN(n2111) );
  NAND2_X1 U2880 ( .A1(n3071), .A2(n3925), .ZN(n2665) );
  OAI21_X1 U2881 ( .B1(n3054), .B2(n2664), .A(n3923), .ZN(n3025) );
  NAND3_X1 U2882 ( .A1(n2403), .A2(n2404), .A3(n2401), .ZN(n2117) );
  NAND2_X1 U2883 ( .A1(n2782), .A2(n4390), .ZN(n2123) );
  INV_X1 U2884 ( .A(n2138), .ZN(n4041) );
  AND2_X1 U2885 ( .A1(n4043), .A2(REG2_REG_18__SCAN_IN), .ZN(n2139) );
  NAND2_X1 U2886 ( .A1(n4094), .A2(n3844), .ZN(n4244) );
  NAND2_X1 U2887 ( .A1(n4094), .A2(n2149), .ZN(n2148) );
  NAND2_X1 U2888 ( .A1(n2158), .A2(n2159), .ZN(n2490) );
  NAND2_X1 U2889 ( .A1(n2159), .A2(n2161), .ZN(n3145) );
  NOR2_X1 U2890 ( .A1(n2260), .A2(n2163), .ZN(n2160) );
  NAND3_X1 U2891 ( .A1(n2319), .A2(n2320), .A3(n2166), .ZN(n2169) );
  INV_X1 U2892 ( .A(n2268), .ZN(n2168) );
  NAND3_X1 U2893 ( .A1(n2180), .A2(n2181), .A3(n2787), .ZN(n2178) );
  NAND3_X1 U2894 ( .A1(n2191), .A2(n4496), .A3(n2192), .ZN(n4494) );
  NAND2_X1 U2895 ( .A1(n4474), .A2(n2193), .ZN(n2191) );
  OAI22_X1 U2896 ( .A1(n2949), .A2(n2948), .B1(n4566), .B2(n2947), .ZN(n4051)
         );
  NOR2_X1 U2897 ( .A1(REG1_REG_16__SCAN_IN), .A2(n4473), .ZN(n4474) );
  NAND2_X1 U2898 ( .A1(n2652), .A2(n2194), .ZN(n2705) );
  NAND2_X1 U2899 ( .A1(n2197), .A2(n2196), .ZN(n3015) );
  NAND2_X1 U2900 ( .A1(n2964), .A2(n2200), .ZN(n2197) );
  AND2_X1 U2901 ( .A1(n2965), .A2(n2966), .ZN(n2201) );
  NAND2_X1 U2902 ( .A1(n3445), .A2(n2205), .ZN(n2204) );
  NAND2_X1 U2903 ( .A1(n3445), .A2(n2210), .ZN(n2209) );
  OAI211_X1 U2904 ( .C1(n2216), .C2(n2206), .A(n2204), .B(n2202), .ZN(n3572)
         );
  NAND2_X1 U2905 ( .A1(n3515), .A2(n2306), .ZN(n2304) );
  NAND2_X1 U2906 ( .A1(n2209), .A2(n2212), .ZN(n3515) );
  INV_X1 U2907 ( .A(n2306), .ZN(n2208) );
  INV_X1 U2908 ( .A(n3186), .ZN(n2218) );
  NAND2_X1 U2909 ( .A1(n2225), .A2(n2226), .ZN(n3699) );
  NAND3_X1 U2910 ( .A1(n3586), .A2(n3803), .A3(n2231), .ZN(n2225) );
  NAND3_X1 U2911 ( .A1(n3586), .A2(n3803), .A3(n2077), .ZN(n2228) );
  NAND3_X1 U2912 ( .A1(n3586), .A2(n3803), .A3(n3718), .ZN(n3728) );
  NAND2_X1 U2913 ( .A1(n2898), .A2(n2237), .ZN(n2234) );
  NAND2_X1 U2914 ( .A1(n2234), .A2(n2236), .ZN(n2951) );
  NAND2_X1 U2915 ( .A1(n2121), .A2(n4388), .ZN(n2239) );
  INV_X1 U2916 ( .A(n4202), .ZN(n2253) );
  NAND2_X1 U2917 ( .A1(n2255), .A2(n2254), .ZN(n3265) );
  NAND2_X1 U2918 ( .A1(n3896), .A2(n2466), .ZN(n2261) );
  INV_X1 U2919 ( .A(n3040), .ZN(n2263) );
  NAND3_X1 U2920 ( .A1(n2335), .A2(n2073), .A3(n2337), .ZN(n2268) );
  NAND2_X1 U2921 ( .A1(n2270), .A2(n2271), .ZN(n3663) );
  NAND2_X1 U2922 ( .A1(n3712), .A2(n2272), .ZN(n2270) );
  NAND2_X1 U2923 ( .A1(n3712), .A2(n3710), .ZN(n2273) );
  INV_X1 U2924 ( .A(n3775), .ZN(n2289) );
  NAND2_X1 U2925 ( .A1(n3281), .A2(n2293), .ZN(n2290) );
  INV_X1 U2926 ( .A(n3442), .ZN(n3441) );
  NAND2_X1 U2927 ( .A1(n2575), .A2(n2299), .ZN(n2298) );
  OAI21_X1 U2928 ( .B1(n3702), .B2(n2090), .A(n2309), .ZN(n3633) );
  NAND3_X1 U2929 ( .A1(n2390), .A2(n2322), .A3(n2389), .ZN(n2817) );
  INV_X1 U2930 ( .A(n2713), .ZN(n4383) );
  OAI21_X1 U2931 ( .B1(n2705), .B2(n2701), .A(IR_REG_31__SCAN_IN), .ZN(n2702)
         );
  AND2_X1 U2932 ( .A1(n2968), .A2(n4521), .ZN(n2876) );
  OR2_X1 U2933 ( .A1(n3485), .A2(n3481), .ZN(n4195) );
  NAND2_X1 U2934 ( .A1(n2649), .A2(IR_REG_31__SCAN_IN), .ZN(n2651) );
  NAND2_X2 U2935 ( .A1(n2927), .A2(n4500), .ZN(n4213) );
  INV_X1 U2936 ( .A(n4378), .ZN(n2739) );
  INV_X2 U2937 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U2938 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3704) );
  NAND2_X1 U2939 ( .A1(n2967), .A2(n2984), .ZN(n2662) );
  INV_X1 U2940 ( .A(n3564), .ZN(n2740) );
  OR2_X1 U2941 ( .A1(n3521), .A2(n3520), .ZN(n2325) );
  NOR2_X1 U2942 ( .A1(n2410), .A2(n2409), .ZN(n2411) );
  INV_X1 U2943 ( .A(n3104), .ZN(n3106) );
  INV_X1 U2944 ( .A(n2814), .ZN(n2815) );
  NOR2_X1 U2945 ( .A1(n2253), .A2(n3703), .ZN(n2616) );
  INV_X1 U2946 ( .A(n4324), .ZN(n3539) );
  AND2_X1 U2947 ( .A1(n3677), .A2(n3678), .ZN(n3623) );
  AND2_X1 U2948 ( .A1(n3630), .A2(n3631), .ZN(n3628) );
  INV_X1 U2949 ( .A(n3579), .ZN(n3803) );
  INV_X1 U2950 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4720) );
  NOR2_X1 U2951 ( .A1(n2393), .A2(n2412), .ZN(n2418) );
  INV_X1 U2952 ( .A(n3897), .ZN(n2514) );
  NOR2_X1 U2953 ( .A1(n2427), .A2(n2610), .ZN(n4235) );
  AND2_X1 U2954 ( .A1(n3981), .A2(n4384), .ZN(n2770) );
  AND2_X1 U2955 ( .A1(n2858), .A2(n2876), .ZN(n2924) );
  NAND2_X1 U2956 ( .A1(n2376), .A2(REG3_REG_23__SCAN_IN), .ZN(n2368) );
  INV_X1 U2957 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2561) );
  INV_X1 U2958 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4690) );
  INV_X1 U2959 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2501) );
  NOR2_X1 U2960 ( .A1(n2622), .A2(n4720), .ZN(n2630) );
  AND2_X1 U2961 ( .A1(n2612), .A2(REG3_REG_22__SCAN_IN), .ZN(n2376) );
  OAI21_X1 U2962 ( .B1(n4255), .B2(n4117), .A(n2629), .ZN(n4092) );
  INV_X1 U2963 ( .A(n3988), .ZN(n4285) );
  INV_X1 U2964 ( .A(n3252), .ZN(n3258) );
  NAND2_X1 U2965 ( .A1(n4548), .A2(n2877), .ZN(n4500) );
  NOR2_X1 U2966 ( .A1(n2427), .A2(n2638), .ZN(n4251) );
  INV_X1 U2967 ( .A(n3449), .ZN(n3454) );
  INV_X1 U2968 ( .A(n2048), .ZN(n4328) );
  NAND2_X1 U2969 ( .A1(n2657), .A2(n4078), .ZN(n4227) );
  NAND2_X1 U2970 ( .A1(n2879), .A2(n2770), .ZN(n4304) );
  AND2_X1 U2971 ( .A1(n2631), .A2(n3563), .ZN(n4096) );
  NOR2_X1 U2972 ( .A1(n2611), .A2(n3704), .ZN(n2612) );
  OR3_X1 U2973 ( .A1(n2563), .A2(n2561), .A3(n2562), .ZN(n2577) );
  OR2_X1 U2974 ( .A1(n2606), .A2(n4690), .ZN(n2611) );
  NOR2_X1 U2975 ( .A1(n2913), .A2(n2914), .ZN(n2964) );
  AND2_X1 U2976 ( .A1(n2870), .A2(n2876), .ZN(n2871) );
  AND3_X1 U2977 ( .A1(n3841), .A2(n3840), .A3(n3839), .ZN(n4086) );
  OR2_X1 U2978 ( .A1(n4164), .A2(n2388), .ZN(n2366) );
  NAND2_X1 U2979 ( .A1(n2690), .A2(n2051), .ZN(n2879) );
  AND2_X1 U2980 ( .A1(n4213), .A2(n2048), .ZN(n3561) );
  AND2_X1 U2981 ( .A1(n3929), .A2(n3925), .ZN(n3888) );
  INV_X1 U2982 ( .A(n4319), .ZN(n2746) );
  AND2_X1 U2983 ( .A1(n2734), .A2(n2733), .ZN(n2853) );
  INV_X1 U2984 ( .A(n3590), .ZN(n3733) );
  INV_X1 U2985 ( .A(n4551), .ZN(n4316) );
  INV_X1 U2986 ( .A(n4540), .ZN(n4548) );
  AND2_X1 U2987 ( .A1(n2522), .A2(n2513), .ZN(n4047) );
  AND2_X1 U2988 ( .A1(n2774), .A2(n2773), .ZN(n4493) );
  AND4_X1 U2989 ( .A1(n3798), .A2(n3797), .A3(n3796), .A4(n3795), .ZN(n3799)
         );
  INV_X1 U2990 ( .A(n4264), .ZN(n3987) );
  NAND2_X1 U2991 ( .A1(n2796), .A2(n2879), .ZN(n4499) );
  XNOR2_X1 U2992 ( .A(n2646), .B(n3883), .ZN(n3569) );
  NAND2_X1 U2993 ( .A1(n4213), .A2(n3042), .ZN(n4198) );
  NAND2_X1 U2994 ( .A1(n4568), .A2(n2811), .ZN(n4319) );
  INV_X1 U2995 ( .A(n4568), .ZN(n4565) );
  NAND2_X1 U2996 ( .A1(n2740), .A2(n2739), .ZN(n2741) );
  NAND2_X1 U2997 ( .A1(n4559), .A2(n2811), .ZN(n4378) );
  INV_X1 U2998 ( .A(n4559), .ZN(n4557) );
  INV_X1 U2999 ( .A(D_REG_1__SCAN_IN), .ZN(n2766) );
  INV_X1 U3000 ( .A(n4047), .ZN(n4532) );
  NAND2_X1 U3001 ( .A1(n2458), .A2(REG3_REG_7__SCAN_IN), .ZN(n2478) );
  NAND2_X1 U3002 ( .A1(REG3_REG_8__SCAN_IN), .A2(REG3_REG_9__SCAN_IN), .ZN(
        n2326) );
  NOR2_X1 U3003 ( .A1(n2478), .A2(n2326), .ZN(n2492) );
  NAND2_X1 U3004 ( .A1(n2492), .A2(REG3_REG_10__SCAN_IN), .ZN(n2502) );
  NAND2_X1 U3005 ( .A1(n2597), .A2(n2327), .ZN(n2606) );
  NAND2_X1 U3006 ( .A1(REG3_REG_25__SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .ZN(
        n2328) );
  AND2_X1 U3007 ( .A1(n2622), .A2(n4720), .ZN(n2329) );
  NAND2_X1 U3008 ( .A1(n2398), .A2(n2330), .ZN(n2405) );
  NOR2_X1 U3009 ( .A1(IR_REG_5__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2331)
         );
  INV_X1 U3010 ( .A(REG2_REG_27__SCAN_IN), .ZN(n2346) );
  NAND2_X2 U3011 ( .A1(n2342), .A2(n2341), .ZN(n2393) );
  INV_X1 U3012 ( .A(n2341), .ZN(n2343) );
  NAND2_X1 U3013 ( .A1(n2414), .A2(REG1_REG_27__SCAN_IN), .ZN(n2345) );
  NAND2_X1 U3014 ( .A1(n2413), .A2(REG0_REG_27__SCAN_IN), .ZN(n2344) );
  OAI211_X1 U3015 ( .C1(n2346), .C2(n2393), .A(n2345), .B(n2344), .ZN(n2347)
         );
  INV_X1 U3016 ( .A(n2347), .ZN(n2348) );
  INV_X1 U3017 ( .A(n4270), .ZN(n4255) );
  NAND2_X1 U3018 ( .A1(n2338), .A2(n2758), .ZN(n2350) );
  NAND2_X2 U3019 ( .A1(n2352), .A2(n2351), .ZN(n2427) );
  INV_X1 U3020 ( .A(DATAI_27_), .ZN(n2353) );
  INV_X1 U3021 ( .A(n4260), .ZN(n4117) );
  NAND2_X1 U3022 ( .A1(n2640), .A2(DATAI_25_), .ZN(n4152) );
  INV_X1 U3023 ( .A(n4152), .ZN(n4146) );
  XNOR2_X1 U3024 ( .A(n2620), .B(REG3_REG_25__SCAN_IN), .ZN(n4153) );
  NAND2_X1 U3025 ( .A1(n4153), .A2(n2382), .ZN(n2359) );
  INV_X1 U3026 ( .A(REG2_REG_25__SCAN_IN), .ZN(n2356) );
  NAND2_X1 U3027 ( .A1(n2414), .A2(REG1_REG_25__SCAN_IN), .ZN(n2355) );
  NAND2_X1 U3028 ( .A1(n2413), .A2(REG0_REG_25__SCAN_IN), .ZN(n2354) );
  OAI211_X1 U3029 ( .C1(n2356), .C2(n2393), .A(n2355), .B(n2354), .ZN(n2357)
         );
  INV_X1 U3030 ( .A(n2357), .ZN(n2358) );
  INV_X1 U3031 ( .A(n4168), .ZN(n4281) );
  NAND2_X1 U3032 ( .A1(n2368), .A2(n4596), .ZN(n2360) );
  NAND2_X1 U3033 ( .A1(n2620), .A2(n2360), .ZN(n4164) );
  INV_X1 U3034 ( .A(REG2_REG_24__SCAN_IN), .ZN(n2363) );
  NAND2_X1 U3035 ( .A1(n2414), .A2(REG1_REG_24__SCAN_IN), .ZN(n2362) );
  NAND2_X1 U3036 ( .A1(n2413), .A2(REG0_REG_24__SCAN_IN), .ZN(n2361) );
  OAI211_X1 U3037 ( .C1(n2363), .C2(n2393), .A(n2362), .B(n2361), .ZN(n2364)
         );
  INV_X1 U3038 ( .A(n2364), .ZN(n2365) );
  OR2_X1 U3039 ( .A1(n2376), .A2(REG3_REG_23__SCAN_IN), .ZN(n2367) );
  AND2_X1 U3040 ( .A1(n2368), .A2(n2367), .ZN(n4193) );
  NAND2_X1 U3041 ( .A1(n4193), .A2(n2382), .ZN(n2374) );
  INV_X1 U3042 ( .A(REG2_REG_23__SCAN_IN), .ZN(n2371) );
  NAND2_X1 U3043 ( .A1(n2414), .A2(REG1_REG_23__SCAN_IN), .ZN(n2370) );
  NAND2_X1 U3044 ( .A1(n2413), .A2(REG0_REG_23__SCAN_IN), .ZN(n2369) );
  OAI211_X1 U3045 ( .C1(n2371), .C2(n2393), .A(n2370), .B(n2369), .ZN(n2372)
         );
  INV_X1 U3046 ( .A(n2372), .ZN(n2373) );
  INV_X1 U3047 ( .A(n4190), .ZN(n3679) );
  NAND2_X1 U3048 ( .A1(n2640), .A2(DATAI_22_), .ZN(n4211) );
  NOR2_X1 U3049 ( .A1(n2612), .A2(REG3_REG_22__SCAN_IN), .ZN(n2375) );
  OR2_X1 U3050 ( .A1(n2376), .A2(n2375), .ZN(n4212) );
  INV_X1 U3051 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4214) );
  NAND2_X1 U3052 ( .A1(n2580), .A2(REG0_REG_22__SCAN_IN), .ZN(n2378) );
  NAND2_X1 U3053 ( .A1(n2414), .A2(REG1_REG_22__SCAN_IN), .ZN(n2377) );
  OAI211_X1 U3054 ( .C1(n2393), .C2(n4214), .A(n2378), .B(n2377), .ZN(n2379)
         );
  INV_X1 U3055 ( .A(n2379), .ZN(n2380) );
  INV_X1 U3056 ( .A(n2393), .ZN(n2381) );
  NAND2_X1 U3057 ( .A1(n2381), .A2(REG2_REG_1__SCAN_IN), .ZN(n2386) );
  INV_X1 U3058 ( .A(n2388), .ZN(n2382) );
  NAND2_X1 U3059 ( .A1(n2382), .A2(REG3_REG_1__SCAN_IN), .ZN(n2385) );
  NAND2_X1 U3060 ( .A1(n2414), .A2(REG1_REG_1__SCAN_IN), .ZN(n2384) );
  NAND2_X1 U3061 ( .A1(n2413), .A2(REG0_REG_1__SCAN_IN), .ZN(n2383) );
  NAND4_X1 U3062 ( .A1(n2386), .A2(n2385), .A3(n2384), .A4(n2383), .ZN(n2387)
         );
  NAND2_X1 U3063 ( .A1(n2387), .A2(n3157), .ZN(n3913) );
  NAND2_X1 U3064 ( .A1(n3004), .A2(n3149), .ZN(n2660) );
  NAND2_X1 U3065 ( .A1(n2414), .A2(REG1_REG_0__SCAN_IN), .ZN(n2390) );
  NAND2_X1 U3066 ( .A1(n2413), .A2(REG0_REG_0__SCAN_IN), .ZN(n2389) );
  INV_X1 U3067 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2891) );
  INV_X1 U3068 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2780) );
  AND2_X1 U3069 ( .A1(n2817), .A2(n3150), .ZN(n3151) );
  NAND2_X1 U3070 ( .A1(n2659), .A2(n3151), .ZN(n3153) );
  NAND2_X1 U3071 ( .A1(n2387), .A2(n3149), .ZN(n2391) );
  NAND2_X1 U3072 ( .A1(n3153), .A2(n2391), .ZN(n2981) );
  INV_X1 U3073 ( .A(n2981), .ZN(n2400) );
  NAND2_X1 U3074 ( .A1(n2414), .A2(REG1_REG_2__SCAN_IN), .ZN(n2397) );
  INV_X1 U3075 ( .A(REG3_REG_2__SCAN_IN), .ZN(n2836) );
  INV_X1 U3076 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2392) );
  NAND2_X1 U3077 ( .A1(n2413), .A2(REG0_REG_2__SCAN_IN), .ZN(n2394) );
  OR2_X1 U3078 ( .A1(n2398), .A2(n2758), .ZN(n2399) );
  MUX2_X1 U3079 ( .A(DATAI_2_), .B(n2049), .S(n2427), .Z(n2984) );
  INV_X1 U3080 ( .A(REG2_REG_3__SCAN_IN), .ZN(n2936) );
  INV_X2 U3081 ( .A(n2402), .ZN(n2580) );
  NAND2_X1 U3082 ( .A1(n2580), .A2(REG0_REG_3__SCAN_IN), .ZN(n2403) );
  NAND2_X1 U3083 ( .A1(n2405), .A2(IR_REG_31__SCAN_IN), .ZN(n2407) );
  NAND2_X1 U3084 ( .A1(n2407), .A2(n2406), .ZN(n2425) );
  OR2_X1 U3085 ( .A1(n2407), .A2(n2406), .ZN(n2408) );
  MUX2_X1 U3086 ( .A(DATAI_3_), .B(n4391), .S(n2427), .Z(n2977) );
  NAND2_X1 U3087 ( .A1(n2967), .A2(n2992), .ZN(n2921) );
  INV_X1 U3088 ( .A(n2921), .ZN(n2409) );
  NAND2_X1 U3089 ( .A1(n4004), .A2(n2977), .ZN(n3057) );
  INV_X1 U3090 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2412) );
  NAND2_X1 U3091 ( .A1(n2413), .A2(REG0_REG_4__SCAN_IN), .ZN(n2416) );
  NAND2_X1 U3092 ( .A1(n2414), .A2(REG1_REG_4__SCAN_IN), .ZN(n2415) );
  NAND2_X1 U3093 ( .A1(n2416), .A2(n2415), .ZN(n2417) );
  INV_X1 U3094 ( .A(n2419), .ZN(n2434) );
  INV_X1 U3095 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2421) );
  INV_X1 U3096 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2420) );
  NAND2_X1 U3097 ( .A1(n2421), .A2(n2420), .ZN(n2422) );
  NAND2_X1 U3098 ( .A1(n2434), .A2(n2422), .ZN(n3052) );
  OR2_X1 U3099 ( .A1(n2388), .A2(n3052), .ZN(n2423) );
  NAND2_X1 U3100 ( .A1(n2425), .A2(IR_REG_31__SCAN_IN), .ZN(n2426) );
  XNOR2_X1 U3101 ( .A(n2426), .B(IR_REG_4__SCAN_IN), .ZN(n4390) );
  MUX2_X1 U3102 ( .A(DATAI_4_), .B(n4390), .S(n2427), .Z(n3051) );
  NAND2_X1 U3103 ( .A1(n4003), .A2(n3051), .ZN(n2429) );
  AND2_X1 U3104 ( .A1(n3057), .A2(n2429), .ZN(n2428) );
  INV_X1 U3105 ( .A(n3051), .ZN(n3056) );
  AND2_X1 U3106 ( .A1(n2429), .A2(n3053), .ZN(n2430) );
  NAND2_X1 U3107 ( .A1(n2414), .A2(REG1_REG_5__SCAN_IN), .ZN(n2439) );
  NAND2_X1 U3108 ( .A1(n2580), .A2(REG0_REG_5__SCAN_IN), .ZN(n2438) );
  INV_X1 U3109 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2431) );
  OR2_X1 U3110 ( .A1(n2393), .A2(n2431), .ZN(n2437) );
  INV_X1 U3111 ( .A(n2432), .ZN(n2448) );
  INV_X1 U3112 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2433) );
  NAND2_X1 U3113 ( .A1(n2434), .A2(n2433), .ZN(n2435) );
  NAND2_X1 U3114 ( .A1(n2448), .A2(n2435), .ZN(n3122) );
  OR2_X1 U3115 ( .A1(n2388), .A2(n3122), .ZN(n2436) );
  NAND4_X1 U3116 ( .A1(n2439), .A2(n2438), .A3(n2437), .A4(n2436), .ZN(n4002)
         );
  INV_X1 U3117 ( .A(n4002), .ZN(n3130) );
  INV_X1 U3118 ( .A(DATAI_5_), .ZN(n4693) );
  NAND2_X1 U3119 ( .A1(n2440), .A2(IR_REG_31__SCAN_IN), .ZN(n2441) );
  MUX2_X1 U3120 ( .A(IR_REG_31__SCAN_IN), .B(n2441), .S(IR_REG_5__SCAN_IN), 
        .Z(n2443) );
  NOR2_X1 U3121 ( .A1(n2440), .A2(IR_REG_5__SCAN_IN), .ZN(n2462) );
  INV_X1 U3122 ( .A(n2462), .ZN(n2442) );
  NAND2_X1 U3123 ( .A1(n2443), .A2(n2442), .ZN(n2801) );
  MUX2_X1 U3124 ( .A(n4693), .B(n2801), .S(n2427), .Z(n3114) );
  NAND2_X1 U3125 ( .A1(n3130), .A2(n3114), .ZN(n2444) );
  NAND2_X1 U3126 ( .A1(n3024), .A2(n2444), .ZN(n2446) );
  INV_X1 U3127 ( .A(n3114), .ZN(n3027) );
  NAND2_X1 U3128 ( .A1(n4002), .A2(n3027), .ZN(n2445) );
  NAND2_X1 U3129 ( .A1(n2446), .A2(n2445), .ZN(n3070) );
  NAND2_X1 U3130 ( .A1(n2414), .A2(REG1_REG_6__SCAN_IN), .ZN(n2454) );
  NAND2_X1 U3131 ( .A1(n2580), .A2(REG0_REG_6__SCAN_IN), .ZN(n2453) );
  OR2_X1 U3132 ( .A1(n2393), .A2(n2238), .ZN(n2452) );
  INV_X1 U3133 ( .A(n2458), .ZN(n2450) );
  INV_X1 U3134 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2447) );
  NAND2_X1 U3135 ( .A1(n2448), .A2(n2447), .ZN(n2449) );
  NAND2_X1 U3136 ( .A1(n2450), .A2(n2449), .ZN(n3137) );
  OR2_X1 U3137 ( .A1(n2388), .A2(n3137), .ZN(n2451) );
  NAND4_X1 U3138 ( .A1(n2454), .A2(n2453), .A3(n2452), .A4(n2451), .ZN(n4001)
         );
  OR2_X1 U3139 ( .A1(n2462), .A2(n2758), .ZN(n2455) );
  XNOR2_X1 U3140 ( .A(n2455), .B(IR_REG_6__SCAN_IN), .ZN(n4388) );
  MUX2_X1 U3141 ( .A(DATAI_6_), .B(n4388), .S(n2427), .Z(n3083) );
  AND2_X1 U3142 ( .A1(n4001), .A2(n3083), .ZN(n2456) );
  INV_X1 U3143 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2457) );
  OR2_X1 U3144 ( .A1(n2393), .A2(n2457), .ZN(n2460) );
  OAI21_X1 U3145 ( .B1(n2458), .B2(REG3_REG_7__SCAN_IN), .A(n2478), .ZN(n3199)
         );
  OR2_X1 U3146 ( .A1(n2388), .A2(n3199), .ZN(n2459) );
  NAND2_X1 U3147 ( .A1(n2462), .A2(n2461), .ZN(n2486) );
  NAND2_X1 U31480 ( .A1(n2486), .A2(IR_REG_31__SCAN_IN), .ZN(n2464) );
  NAND2_X1 U31490 ( .A1(n2464), .A2(n2463), .ZN(n2472) );
  OR2_X1 U3150 ( .A1(n2464), .A2(n2463), .ZN(n2465) );
  MUX2_X1 U3151 ( .A(DATAI_7_), .B(n4387), .S(n2427), .Z(n3188) );
  INV_X1 U3152 ( .A(n3188), .ZN(n3193) );
  NAND2_X1 U3153 ( .A1(n3999), .A2(n3193), .ZN(n3932) );
  NAND2_X1 U3154 ( .A1(n3999), .A2(n3188), .ZN(n2466) );
  NAND2_X1 U3155 ( .A1(n2414), .A2(REG1_REG_8__SCAN_IN), .ZN(n2471) );
  NAND2_X1 U3156 ( .A1(n2580), .A2(REG0_REG_8__SCAN_IN), .ZN(n2470) );
  INV_X1 U3157 ( .A(REG2_REG_8__SCAN_IN), .ZN(n4502) );
  OR2_X1 U3158 ( .A1(n2393), .A2(n4502), .ZN(n2469) );
  INV_X1 U3159 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2467) );
  XNOR2_X1 U3160 ( .A(n2478), .B(n2467), .ZN(n4501) );
  OR2_X1 U3161 ( .A1(n2388), .A2(n4501), .ZN(n2468) );
  NAND4_X1 U3162 ( .A1(n2471), .A2(n2470), .A3(n2469), .A4(n2468), .ZN(n3998)
         );
  INV_X1 U3163 ( .A(DATAI_8_), .ZN(n2475) );
  NAND2_X1 U3164 ( .A1(n2472), .A2(IR_REG_31__SCAN_IN), .ZN(n2474) );
  INV_X1 U3165 ( .A(IR_REG_8__SCAN_IN), .ZN(n2473) );
  XNOR2_X1 U3166 ( .A(n2474), .B(n2473), .ZN(n4050) );
  MUX2_X1 U3167 ( .A(n2475), .B(n4050), .S(n2427), .Z(n3238) );
  NAND2_X1 U3168 ( .A1(n3257), .A2(n3238), .ZN(n2476) );
  INV_X1 U3169 ( .A(n3238), .ZN(n3233) );
  NAND2_X1 U3170 ( .A1(n3998), .A2(n3233), .ZN(n2477) );
  NAND2_X1 U3171 ( .A1(n2414), .A2(REG1_REG_9__SCAN_IN), .ZN(n2485) );
  NAND2_X1 U3172 ( .A1(n2580), .A2(REG0_REG_9__SCAN_IN), .ZN(n2484) );
  INV_X1 U3173 ( .A(n2478), .ZN(n2479) );
  AOI21_X1 U3174 ( .B1(n2479), .B2(REG3_REG_8__SCAN_IN), .A(
        REG3_REG_9__SCAN_IN), .ZN(n2480) );
  OR2_X1 U3175 ( .A1(n2480), .A2(n2492), .ZN(n3264) );
  OR2_X1 U3176 ( .A1(n2388), .A2(n3264), .ZN(n2483) );
  INV_X1 U3177 ( .A(REG2_REG_9__SCAN_IN), .ZN(n2481) );
  OR2_X1 U3178 ( .A1(n2393), .A2(n2481), .ZN(n2482) );
  NAND4_X1 U3179 ( .A1(n2485), .A2(n2484), .A3(n2483), .A4(n2482), .ZN(n3997)
         );
  NAND2_X1 U3180 ( .A1(n2498), .A2(IR_REG_31__SCAN_IN), .ZN(n2487) );
  XNOR2_X1 U3181 ( .A(n2487), .B(IR_REG_9__SCAN_IN), .ZN(n4049) );
  MUX2_X1 U3182 ( .A(DATAI_9_), .B(n4049), .S(n2427), .Z(n3252) );
  AND2_X1 U3183 ( .A1(n3997), .A2(n3252), .ZN(n2488) );
  NAND2_X1 U3184 ( .A1(n3290), .A2(n3258), .ZN(n2489) );
  NAND2_X1 U3185 ( .A1(n2414), .A2(REG1_REG_10__SCAN_IN), .ZN(n2497) );
  NAND2_X1 U3186 ( .A1(n2580), .A2(REG0_REG_10__SCAN_IN), .ZN(n2496) );
  INV_X1 U3187 ( .A(REG2_REG_10__SCAN_IN), .ZN(n2491) );
  OR2_X1 U3188 ( .A1(n2393), .A2(n2491), .ZN(n2495) );
  OR2_X1 U3189 ( .A1(n2492), .A2(REG3_REG_10__SCAN_IN), .ZN(n2493) );
  NAND2_X1 U3190 ( .A1(n2502), .A2(n2493), .ZN(n3295) );
  OR2_X1 U3191 ( .A1(n2388), .A2(n3295), .ZN(n2494) );
  NAND4_X1 U3192 ( .A1(n2497), .A2(n2496), .A3(n2495), .A4(n2494), .ZN(n3996)
         );
  NOR2_X1 U3193 ( .A1(n2498), .A2(IR_REG_9__SCAN_IN), .ZN(n2509) );
  OR2_X1 U3194 ( .A1(n2509), .A2(n2758), .ZN(n2499) );
  XNOR2_X1 U3195 ( .A(n2499), .B(IR_REG_10__SCAN_IN), .ZN(n4055) );
  MUX2_X1 U3196 ( .A(DATAI_10_), .B(n4055), .S(n2427), .Z(n3282) );
  NOR2_X1 U3197 ( .A1(n3996), .A2(n3282), .ZN(n2500) );
  INV_X1 U3198 ( .A(n3282), .ZN(n3289) );
  NAND2_X1 U3199 ( .A1(n2414), .A2(REG1_REG_11__SCAN_IN), .ZN(n2507) );
  NAND2_X1 U3200 ( .A1(n2580), .A2(REG0_REG_11__SCAN_IN), .ZN(n2506) );
  INV_X1 U3201 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3271) );
  OR2_X1 U3202 ( .A1(n2393), .A2(n3271), .ZN(n2505) );
  NAND2_X1 U3203 ( .A1(n2502), .A2(n2501), .ZN(n2503) );
  NAND2_X1 U3204 ( .A1(n2516), .A2(n2503), .ZN(n3405) );
  OR2_X1 U3205 ( .A1(n2388), .A2(n3405), .ZN(n2504) );
  NAND4_X1 U3206 ( .A1(n2507), .A2(n2506), .A3(n2505), .A4(n2504), .ZN(n3995)
         );
  INV_X1 U3207 ( .A(IR_REG_10__SCAN_IN), .ZN(n2508) );
  NAND2_X1 U3208 ( .A1(n2509), .A2(n2508), .ZN(n2510) );
  NAND2_X1 U3209 ( .A1(n2510), .A2(IR_REG_31__SCAN_IN), .ZN(n2512) );
  NAND2_X1 U32100 ( .A1(n2512), .A2(n2511), .ZN(n2522) );
  OR2_X1 U32110 ( .A1(n2512), .A2(n2511), .ZN(n2513) );
  MUX2_X1 U32120 ( .A(DATAI_11_), .B(n4047), .S(n2427), .Z(n3395) );
  NAND2_X1 U32130 ( .A1(n3455), .A2(n3395), .ZN(n3299) );
  NAND2_X1 U32140 ( .A1(n3995), .A2(n3399), .ZN(n3301) );
  NAND2_X1 U32150 ( .A1(n3455), .A2(n3399), .ZN(n2515) );
  NAND2_X1 U32160 ( .A1(n3265), .A2(n2515), .ZN(n3313) );
  NAND2_X1 U32170 ( .A1(n2414), .A2(REG1_REG_12__SCAN_IN), .ZN(n2521) );
  NAND2_X1 U32180 ( .A1(n2580), .A2(REG0_REG_12__SCAN_IN), .ZN(n2520) );
  INV_X1 U32190 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3319) );
  OR2_X1 U32200 ( .A1(n2393), .A2(n3319), .ZN(n2519) );
  AND2_X1 U32210 ( .A1(n2516), .A2(n4724), .ZN(n2517) );
  OR2_X1 U32220 ( .A1(n2517), .A2(n2527), .ZN(n3460) );
  OR2_X1 U32230 ( .A1(n2388), .A2(n3460), .ZN(n2518) );
  NAND4_X1 U32240 ( .A1(n2521), .A2(n2520), .A3(n2519), .A4(n2518), .ZN(n3994)
         );
  NAND2_X1 U32250 ( .A1(n2522), .A2(IR_REG_31__SCAN_IN), .ZN(n2523) );
  XNOR2_X1 U32260 ( .A(n2523), .B(IR_REG_12__SCAN_IN), .ZN(n4059) );
  MUX2_X1 U32270 ( .A(DATAI_12_), .B(n4059), .S(n2427), .Z(n3449) );
  NAND2_X1 U32280 ( .A1(n3994), .A2(n3449), .ZN(n2524) );
  NAND2_X1 U32290 ( .A1(n3313), .A2(n2524), .ZN(n2526) );
  INV_X1 U32300 ( .A(n3994), .ZN(n3496) );
  NAND2_X1 U32310 ( .A1(n3496), .A2(n3454), .ZN(n2525) );
  NAND2_X1 U32320 ( .A1(n2526), .A2(n2525), .ZN(n3339) );
  NAND2_X1 U32330 ( .A1(n2414), .A2(REG1_REG_13__SCAN_IN), .ZN(n2532) );
  NAND2_X1 U32340 ( .A1(n2580), .A2(REG0_REG_13__SCAN_IN), .ZN(n2531) );
  NOR2_X1 U32350 ( .A1(n2527), .A2(REG3_REG_13__SCAN_IN), .ZN(n2528) );
  OR2_X1 U32360 ( .A1(n2535), .A2(n2528), .ZN(n3503) );
  OR2_X1 U32370 ( .A1(n2388), .A2(n3503), .ZN(n2530) );
  INV_X1 U32380 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4439) );
  OR2_X1 U32390 ( .A1(n2393), .A2(n4439), .ZN(n2529) );
  NAND4_X1 U32400 ( .A1(n2532), .A2(n2531), .A3(n2530), .A4(n2529), .ZN(n3993)
         );
  OR2_X1 U32410 ( .A1(n2542), .A2(n2758), .ZN(n2533) );
  XNOR2_X1 U32420 ( .A(n2533), .B(IR_REG_13__SCAN_IN), .ZN(n4046) );
  MUX2_X1 U32430 ( .A(DATAI_13_), .B(n4046), .S(n2427), .Z(n3492) );
  NOR2_X1 U32440 ( .A1(n3993), .A2(n3492), .ZN(n3338) );
  NAND2_X1 U32450 ( .A1(n2414), .A2(REG1_REG_14__SCAN_IN), .ZN(n2540) );
  NAND2_X1 U32460 ( .A1(n2580), .A2(REG0_REG_14__SCAN_IN), .ZN(n2539) );
  INV_X1 U32470 ( .A(REG2_REG_14__SCAN_IN), .ZN(n2534) );
  OR2_X1 U32480 ( .A1(n2393), .A2(n2534), .ZN(n2538) );
  OR2_X1 U32490 ( .A1(n2535), .A2(REG3_REG_14__SCAN_IN), .ZN(n2536) );
  NAND2_X1 U32500 ( .A1(n2563), .A2(n2536), .ZN(n3531) );
  OR2_X1 U32510 ( .A1(n2388), .A2(n3531), .ZN(n2537) );
  NAND4_X1 U32520 ( .A1(n2540), .A2(n2539), .A3(n2538), .A4(n2537), .ZN(n3992)
         );
  OR2_X1 U32530 ( .A1(n2575), .A2(n2758), .ZN(n2543) );
  XNOR2_X1 U32540 ( .A(n2543), .B(IR_REG_14__SCAN_IN), .ZN(n4063) );
  MUX2_X1 U32550 ( .A(DATAI_14_), .B(n4063), .S(n2427), .Z(n3519) );
  INV_X1 U32560 ( .A(n3519), .ZN(n3524) );
  AND2_X1 U32570 ( .A1(n3809), .A2(n3524), .ZN(n2555) );
  OR2_X1 U32580 ( .A1(n3338), .A2(n2555), .ZN(n2544) );
  NAND2_X1 U32590 ( .A1(n2414), .A2(REG1_REG_15__SCAN_IN), .ZN(n2549) );
  NAND2_X1 U32600 ( .A1(n2580), .A2(REG0_REG_15__SCAN_IN), .ZN(n2548) );
  INV_X1 U32610 ( .A(REG2_REG_15__SCAN_IN), .ZN(n2545) );
  OR2_X1 U32620 ( .A1(n2393), .A2(n2545), .ZN(n2547) );
  XNOR2_X1 U32630 ( .A(n2563), .B(n2562), .ZN(n3818) );
  OR2_X1 U32640 ( .A1(n2388), .A2(n3818), .ZN(n2546) );
  NAND4_X1 U32650 ( .A1(n2549), .A2(n2548), .A3(n2547), .A4(n2546), .ZN(n3991)
         );
  INV_X1 U32660 ( .A(IR_REG_14__SCAN_IN), .ZN(n2550) );
  NAND2_X1 U32670 ( .A1(n2575), .A2(n2550), .ZN(n2551) );
  NAND2_X1 U32680 ( .A1(n2551), .A2(IR_REG_31__SCAN_IN), .ZN(n2553) );
  NAND2_X1 U32690 ( .A1(n2553), .A2(n2552), .ZN(n2569) );
  OR2_X1 U32700 ( .A1(n2553), .A2(n2552), .ZN(n2554) );
  MUX2_X1 U32710 ( .A(DATAI_15_), .B(n4044), .S(n2427), .Z(n3574) );
  NAND2_X1 U32720 ( .A1(n3991), .A2(n3574), .ZN(n2556) );
  NAND2_X1 U32730 ( .A1(n3809), .A2(n3519), .ZN(n3820) );
  NAND2_X1 U32740 ( .A1(n3992), .A2(n3524), .ZN(n3828) );
  NAND2_X1 U32750 ( .A1(n3820), .A2(n3828), .ZN(n3344) );
  NAND2_X1 U32760 ( .A1(n3993), .A2(n3492), .ZN(n3340) );
  AND2_X1 U32770 ( .A1(n3344), .A2(n3340), .ZN(n3341) );
  OR2_X1 U32780 ( .A1(n2555), .A2(n3341), .ZN(n3359) );
  AND2_X1 U32790 ( .A1(n2556), .A2(n3359), .ZN(n2557) );
  NAND2_X1 U32800 ( .A1(n3360), .A2(n2557), .ZN(n2559) );
  NAND2_X1 U32810 ( .A1(n4329), .A2(n3810), .ZN(n2558) );
  NAND2_X1 U32820 ( .A1(n2414), .A2(REG1_REG_16__SCAN_IN), .ZN(n2568) );
  NAND2_X1 U32830 ( .A1(n2580), .A2(REG0_REG_16__SCAN_IN), .ZN(n2567) );
  INV_X1 U32840 ( .A(REG2_REG_16__SCAN_IN), .ZN(n2560) );
  OR2_X1 U32850 ( .A1(n2393), .A2(n2560), .ZN(n2566) );
  OAI21_X1 U32860 ( .B1(n2563), .B2(n2562), .A(n2561), .ZN(n2564) );
  NAND2_X1 U32870 ( .A1(n2564), .A2(n2577), .ZN(n3726) );
  OR2_X1 U32880 ( .A1(n2388), .A2(n3726), .ZN(n2565) );
  NAND4_X1 U32890 ( .A1(n2568), .A2(n2567), .A3(n2566), .A4(n2565), .ZN(n3990)
         );
  INV_X1 U32900 ( .A(n3990), .ZN(n3812) );
  NAND2_X1 U32910 ( .A1(n2569), .A2(IR_REG_31__SCAN_IN), .ZN(n2570) );
  XNOR2_X1 U32920 ( .A(n2570), .B(IR_REG_16__SCAN_IN), .ZN(n4524) );
  MUX2_X1 U32930 ( .A(DATAI_16_), .B(n4524), .S(n2427), .Z(n4323) );
  NAND2_X1 U32940 ( .A1(n3812), .A2(n4323), .ZN(n3950) );
  INV_X1 U32950 ( .A(n4323), .ZN(n3721) );
  NAND2_X1 U32960 ( .A1(n3990), .A2(n3721), .ZN(n3822) );
  NAND2_X1 U32970 ( .A1(n3990), .A2(n4323), .ZN(n2571) );
  INV_X1 U32980 ( .A(n2572), .ZN(n2573) );
  NOR2_X1 U32990 ( .A1(n2573), .A2(IR_REG_16__SCAN_IN), .ZN(n2574) );
  NAND2_X1 U33000 ( .A1(n2593), .A2(IR_REG_31__SCAN_IN), .ZN(n2576) );
  XNOR2_X1 U33010 ( .A(n2576), .B(IR_REG_17__SCAN_IN), .ZN(n4070) );
  MUX2_X1 U33020 ( .A(DATAI_17_), .B(n4070), .S(n2427), .Z(n3590) );
  AND2_X1 U33030 ( .A1(n2577), .A2(n4573), .ZN(n2578) );
  NOR2_X1 U33040 ( .A1(n2597), .A2(n2578), .ZN(n3738) );
  NAND2_X1 U33050 ( .A1(n3738), .A2(n2382), .ZN(n2584) );
  INV_X1 U33060 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2579) );
  OR2_X1 U33070 ( .A1(n2393), .A2(n2579), .ZN(n2583) );
  NAND2_X1 U33080 ( .A1(n2414), .A2(REG1_REG_17__SCAN_IN), .ZN(n2582) );
  NAND2_X1 U33090 ( .A1(n2580), .A2(REG0_REG_17__SCAN_IN), .ZN(n2581) );
  NAND4_X1 U33100 ( .A1(n2584), .A2(n2583), .A3(n2582), .A4(n2581), .ZN(n4326)
         );
  OR2_X1 U33110 ( .A1(n3590), .A2(n4326), .ZN(n2585) );
  INV_X1 U33120 ( .A(REG0_REG_18__SCAN_IN), .ZN(n2592) );
  INV_X1 U33130 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2586) );
  XNOR2_X1 U33140 ( .A(n2597), .B(n2586), .ZN(n3783) );
  NAND2_X1 U33150 ( .A1(n3783), .A2(n2382), .ZN(n2591) );
  NAND2_X1 U33160 ( .A1(n2414), .A2(REG1_REG_18__SCAN_IN), .ZN(n2589) );
  INV_X1 U33170 ( .A(REG2_REG_18__SCAN_IN), .ZN(n2587) );
  OR2_X1 U33180 ( .A1(n2393), .A2(n2587), .ZN(n2588) );
  AND2_X1 U33190 ( .A1(n2589), .A2(n2588), .ZN(n2590) );
  OAI211_X1 U33200 ( .C1(n2402), .C2(n2592), .A(n2591), .B(n2590), .ZN(n3989)
         );
  INV_X1 U33210 ( .A(DATAI_18_), .ZN(n2595) );
  NAND2_X1 U33220 ( .A1(n2604), .A2(IR_REG_31__SCAN_IN), .ZN(n2594) );
  XNOR2_X1 U33230 ( .A(n2594), .B(IR_REG_18__SCAN_IN), .ZN(n4043) );
  MUX2_X1 U33240 ( .A(n2595), .B(n4522), .S(n2427), .Z(n3778) );
  OR2_X1 U33250 ( .A1(n3989), .A2(n3778), .ZN(n3533) );
  NAND2_X1 U33260 ( .A1(n3989), .A2(n3778), .ZN(n3534) );
  NAND2_X1 U33270 ( .A1(n3533), .A2(n3534), .ZN(n3477) );
  INV_X1 U33280 ( .A(n3989), .ZN(n3735) );
  NAND2_X1 U33290 ( .A1(n3735), .A2(n3778), .ZN(n2596) );
  INV_X1 U33300 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4376) );
  NAND2_X1 U33310 ( .A1(n2597), .A2(REG3_REG_18__SCAN_IN), .ZN(n2598) );
  INV_X1 U33320 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4598) );
  NAND2_X1 U33330 ( .A1(n2598), .A2(n4598), .ZN(n2599) );
  NAND2_X1 U33340 ( .A1(n2599), .A2(n2606), .ZN(n3692) );
  OR2_X1 U33350 ( .A1(n3692), .A2(n2388), .ZN(n2603) );
  NAND2_X1 U33360 ( .A1(n2414), .A2(REG1_REG_19__SCAN_IN), .ZN(n2601) );
  INV_X1 U33370 ( .A(REG2_REG_19__SCAN_IN), .ZN(n3545) );
  OR2_X1 U33380 ( .A1(n2393), .A2(n3545), .ZN(n2600) );
  AND2_X1 U33390 ( .A1(n2601), .A2(n2600), .ZN(n2602) );
  MUX2_X1 U33400 ( .A(DATAI_19_), .B(n4385), .S(n2427), .Z(n3599) );
  NAND2_X1 U33410 ( .A1(n4223), .A2(n3599), .ZN(n2605) );
  NAND2_X1 U33420 ( .A1(n2606), .A2(n4690), .ZN(n2607) );
  NAND2_X1 U33430 ( .A1(n2611), .A2(n2607), .ZN(n4232) );
  AOI22_X1 U33440 ( .A1(n2381), .A2(REG2_REG_20__SCAN_IN), .B1(n2414), .B2(
        REG1_REG_20__SCAN_IN), .ZN(n2609) );
  NAND2_X1 U33450 ( .A1(n2413), .A2(REG0_REG_20__SCAN_IN), .ZN(n2608) );
  INV_X1 U33460 ( .A(DATAI_20_), .ZN(n2610) );
  AND2_X1 U33470 ( .A1(n4301), .A2(n4235), .ZN(n3877) );
  OR2_X1 U33480 ( .A1(n4301), .A2(n4235), .ZN(n3878) );
  OAI21_X1 U33490 ( .B1(n4226), .B2(n3877), .A(n3878), .ZN(n3551) );
  AND2_X1 U33500 ( .A1(n2611), .A2(n3704), .ZN(n2613) );
  OR2_X1 U33510 ( .A1(n2613), .A2(n2612), .ZN(n3709) );
  AOI22_X1 U33520 ( .A1(n2381), .A2(REG2_REG_21__SCAN_IN), .B1(n2414), .B2(
        REG1_REG_21__SCAN_IN), .ZN(n2615) );
  NAND2_X1 U3353 ( .A1(n2413), .A2(REG0_REG_21__SCAN_IN), .ZN(n2614) );
  INV_X1 U33540 ( .A(n3703), .ZN(n4299) );
  OR2_X1 U3355 ( .A1(n4186), .A2(n4211), .ZN(n4181) );
  NAND2_X1 U3356 ( .A1(n4186), .A2(n4211), .ZN(n2682) );
  OAI21_X1 U3357 ( .B1(n4189), .B2(n4168), .A(n4160), .ZN(n2618) );
  INV_X1 U3358 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4726) );
  INV_X1 U3359 ( .A(REG3_REG_26__SCAN_IN), .ZN(n2619) );
  OAI21_X1 U3360 ( .B1(n2620), .B2(n4726), .A(n2619), .ZN(n2621) );
  NAND2_X1 U3361 ( .A1(n4132), .A2(n2382), .ZN(n2628) );
  INV_X1 U3362 ( .A(REG2_REG_26__SCAN_IN), .ZN(n2625) );
  NAND2_X1 U3363 ( .A1(n2414), .A2(REG1_REG_26__SCAN_IN), .ZN(n2624) );
  NAND2_X1 U3364 ( .A1(n2413), .A2(REG0_REG_26__SCAN_IN), .ZN(n2623) );
  OAI211_X1 U3365 ( .C1(n2625), .C2(n2393), .A(n2624), .B(n2623), .ZN(n2626)
         );
  INV_X1 U3366 ( .A(n2626), .ZN(n2627) );
  NAND2_X1 U3367 ( .A1(n2640), .A2(DATAI_26_), .ZN(n4134) );
  NAND2_X1 U3368 ( .A1(n4261), .A2(n4269), .ZN(n3861) );
  NOR2_X1 U3369 ( .A1(n4261), .A2(n4269), .ZN(n3862) );
  OAI21_X1 U3370 ( .B1(n4260), .B2(n4270), .A(n4111), .ZN(n2629) );
  OR2_X1 U3371 ( .A1(n2630), .A2(REG3_REG_28__SCAN_IN), .ZN(n2631) );
  NAND2_X1 U3372 ( .A1(n2630), .A2(REG3_REG_28__SCAN_IN), .ZN(n3563) );
  NAND2_X1 U3373 ( .A1(n4096), .A2(n2382), .ZN(n2637) );
  INV_X1 U3374 ( .A(REG2_REG_28__SCAN_IN), .ZN(n2634) );
  NAND2_X1 U3375 ( .A1(n2413), .A2(REG0_REG_28__SCAN_IN), .ZN(n2633) );
  NAND2_X1 U3376 ( .A1(n2414), .A2(REG1_REG_28__SCAN_IN), .ZN(n2632) );
  OAI211_X1 U3377 ( .C1(n2393), .C2(n2634), .A(n2633), .B(n2632), .ZN(n2635)
         );
  INV_X1 U3378 ( .A(n2635), .ZN(n2636) );
  INV_X1 U3379 ( .A(DATAI_28_), .ZN(n2638) );
  AND2_X1 U3380 ( .A1(n4264), .A2(n4251), .ZN(n3838) );
  INV_X1 U3381 ( .A(n3838), .ZN(n2639) );
  INV_X1 U3382 ( .A(n4251), .ZN(n4098) );
  NAND2_X1 U3383 ( .A1(n3987), .A2(n4098), .ZN(n3846) );
  NAND2_X1 U3384 ( .A1(n2639), .A2(n3846), .ZN(n4093) );
  AOI22_X1 U3385 ( .A1(n4092), .A2(n4093), .B1(n4251), .B2(n3987), .ZN(n2646)
         );
  NAND2_X1 U3386 ( .A1(n2640), .A2(DATAI_29_), .ZN(n3844) );
  OR2_X1 U3387 ( .A1(n3563), .A2(n2388), .ZN(n2645) );
  INV_X1 U3388 ( .A(REG2_REG_29__SCAN_IN), .ZN(n3559) );
  NAND2_X1 U3389 ( .A1(n2413), .A2(REG0_REG_29__SCAN_IN), .ZN(n2642) );
  NAND2_X1 U3390 ( .A1(n2414), .A2(REG1_REG_29__SCAN_IN), .ZN(n2641) );
  OAI211_X1 U3391 ( .C1(n2393), .C2(n3559), .A(n2642), .B(n2641), .ZN(n2643)
         );
  INV_X1 U3392 ( .A(n2643), .ZN(n2644) );
  NAND2_X1 U3393 ( .A1(n2645), .A2(n2644), .ZN(n4252) );
  XOR2_X1 U3394 ( .A(n3844), .B(n4252), .Z(n3883) );
  NAND2_X1 U3395 ( .A1(n2648), .A2(n2647), .ZN(n2649) );
  XNOR2_X1 U3396 ( .A(n2651), .B(n2650), .ZN(n2658) );
  INV_X1 U3397 ( .A(n2652), .ZN(n2653) );
  NAND2_X1 U3398 ( .A1(n2653), .A2(IR_REG_31__SCAN_IN), .ZN(n2654) );
  NAND2_X1 U3399 ( .A1(n2699), .A2(IR_REG_31__SCAN_IN), .ZN(n2656) );
  XNOR2_X1 U3400 ( .A(n2812), .B(n3981), .ZN(n2657) );
  NAND2_X1 U3401 ( .A1(n2658), .A2(n4385), .ZN(n3005) );
  OR2_X1 U3402 ( .A1(n3005), .A2(n3981), .ZN(n4540) );
  NAND2_X1 U3403 ( .A1(n2982), .A2(n2662), .ZN(n2929) );
  INV_X1 U3404 ( .A(n2977), .ZN(n2961) );
  NAND2_X1 U3405 ( .A1(n4004), .A2(n2961), .ZN(n3917) );
  NAND2_X1 U3406 ( .A1(n2929), .A2(n3893), .ZN(n2663) );
  NAND2_X1 U3407 ( .A1(n2663), .A2(n3920), .ZN(n3054) );
  INV_X1 U3408 ( .A(n3921), .ZN(n2664) );
  NAND2_X1 U3409 ( .A1(n3130), .A2(n3027), .ZN(n3927) );
  INV_X1 U3410 ( .A(n3083), .ZN(n3131) );
  NAND2_X1 U3411 ( .A1(n4001), .A2(n3131), .ZN(n3925) );
  INV_X1 U3412 ( .A(n4001), .ZN(n3192) );
  NAND2_X1 U3413 ( .A1(n3192), .A2(n3083), .ZN(n3929) );
  NAND2_X1 U3414 ( .A1(n2665), .A2(n3929), .ZN(n3034) );
  INV_X1 U3415 ( .A(n3930), .ZN(n2666) );
  NAND2_X1 U3416 ( .A1(n2667), .A2(n3932), .ZN(n3232) );
  NAND2_X1 U3417 ( .A1(n3257), .A2(n3233), .ZN(n3935) );
  NAND2_X1 U3418 ( .A1(n3998), .A2(n3238), .ZN(n3931) );
  AND2_X1 U3419 ( .A1(n3997), .A2(n3258), .ZN(n3138) );
  NAND2_X1 U3420 ( .A1(n3290), .A2(n3252), .ZN(n3936) );
  NAND2_X1 U3421 ( .A1(n3996), .A2(n3289), .ZN(n3940) );
  NAND2_X1 U3422 ( .A1(n3165), .A2(n3940), .ZN(n2668) );
  NAND2_X1 U3423 ( .A1(n3398), .A2(n3282), .ZN(n3944) );
  NAND2_X1 U3424 ( .A1(n2668), .A2(n3944), .ZN(n3302) );
  NAND2_X1 U3425 ( .A1(n3994), .A2(n3454), .ZN(n3314) );
  NAND2_X1 U3426 ( .A1(n3993), .A2(n3497), .ZN(n3296) );
  NAND2_X1 U3427 ( .A1(n3314), .A2(n3296), .ZN(n2670) );
  INV_X1 U3428 ( .A(n3301), .ZN(n2669) );
  NOR2_X1 U3429 ( .A1(n2670), .A2(n2669), .ZN(n3941) );
  NAND2_X1 U3430 ( .A1(n3302), .A2(n3941), .ZN(n2673) );
  NAND2_X1 U3431 ( .A1(n3496), .A2(n3449), .ZN(n3315) );
  NAND2_X1 U3432 ( .A1(n3299), .A2(n3315), .ZN(n2672) );
  INV_X1 U3433 ( .A(n2670), .ZN(n2671) );
  NOR2_X1 U3434 ( .A1(n3993), .A2(n3497), .ZN(n3297) );
  AOI21_X1 U3435 ( .B1(n2672), .B2(n2671), .A(n3297), .ZN(n3946) );
  NAND2_X1 U3436 ( .A1(n2673), .A2(n3946), .ZN(n3821) );
  INV_X1 U3437 ( .A(n3344), .ZN(n3898) );
  NAND2_X1 U3438 ( .A1(n3821), .A2(n3898), .ZN(n2674) );
  NAND2_X1 U3439 ( .A1(n4329), .A2(n3574), .ZN(n3824) );
  NAND2_X1 U3440 ( .A1(n3991), .A2(n3810), .ZN(n3827) );
  NAND2_X1 U3441 ( .A1(n3824), .A2(n3827), .ZN(n3892) );
  INV_X1 U3442 ( .A(n3599), .ZN(n3688) );
  NAND2_X1 U3443 ( .A1(n4223), .A2(n3688), .ZN(n2675) );
  NAND2_X1 U3444 ( .A1(n3534), .A2(n2675), .ZN(n2676) );
  AND2_X1 U3445 ( .A1(n4326), .A2(n3733), .ZN(n3475) );
  OR2_X1 U3446 ( .A1(n2676), .A2(n3475), .ZN(n3829) );
  INV_X1 U3447 ( .A(n2676), .ZN(n2679) );
  OR2_X1 U3448 ( .A1(n3733), .A2(n4326), .ZN(n3474) );
  NAND2_X1 U3449 ( .A1(n3533), .A2(n3474), .ZN(n2678) );
  NOR2_X1 U3450 ( .A1(n4223), .A2(n3688), .ZN(n2677) );
  AOI21_X1 U3451 ( .B1(n2679), .B2(n2678), .A(n2677), .ZN(n4219) );
  OR2_X1 U3452 ( .A1(n4301), .A2(n3757), .ZN(n2680) );
  NAND2_X1 U3453 ( .A1(n4220), .A2(n3951), .ZN(n2681) );
  NAND2_X1 U3454 ( .A1(n4301), .A2(n3757), .ZN(n3831) );
  OR2_X1 U3455 ( .A1(n4202), .A2(n3703), .ZN(n4179) );
  AND2_X1 U3456 ( .A1(n4181), .A2(n4179), .ZN(n3958) );
  NAND2_X1 U3457 ( .A1(n4178), .A2(n3958), .ZN(n2685) );
  OR2_X1 U34580 ( .A1(n4204), .A2(n4190), .ZN(n3866) );
  AND2_X1 U34590 ( .A1(n3866), .A2(n2682), .ZN(n3962) );
  AND2_X1 U3460 ( .A1(n4202), .A2(n3703), .ZN(n4177) );
  NAND2_X1 U3461 ( .A1(n4181), .A2(n4177), .ZN(n2683) );
  NAND2_X1 U3462 ( .A1(n3962), .A2(n2683), .ZN(n3836) );
  INV_X1 U3463 ( .A(n3836), .ZN(n2684) );
  AND2_X1 U3464 ( .A1(n4204), .A2(n4190), .ZN(n3834) );
  INV_X1 U3465 ( .A(n3834), .ZN(n3867) );
  NOR2_X1 U3466 ( .A1(n4147), .A2(n4168), .ZN(n3865) );
  OR2_X1 U34670 ( .A1(n3988), .A2(n4152), .ZN(n4124) );
  OAI21_X1 U3468 ( .B1(n4261), .B2(n4134), .A(n4124), .ZN(n3960) );
  NAND2_X1 U34690 ( .A1(n3988), .A2(n4152), .ZN(n3860) );
  NAND2_X1 U3470 ( .A1(n4147), .A2(n4168), .ZN(n4141) );
  AND2_X1 U34710 ( .A1(n3860), .A2(n4141), .ZN(n4123) );
  OR2_X1 U3472 ( .A1(n3960), .A2(n4123), .ZN(n2686) );
  NAND2_X1 U34730 ( .A1(n4261), .A2(n4134), .ZN(n3847) );
  NAND2_X1 U3474 ( .A1(n2686), .A2(n3847), .ZN(n3965) );
  INV_X1 U34750 ( .A(n3965), .ZN(n2687) );
  XNOR2_X1 U3476 ( .A(n4270), .B(n4260), .ZN(n4110) );
  INV_X1 U34770 ( .A(n4110), .ZN(n4105) );
  NOR2_X1 U3478 ( .A1(n4106), .A2(n4105), .ZN(n4108) );
  NOR2_X1 U34790 ( .A1(n4270), .A2(n4117), .ZN(n3837) );
  INV_X1 U3480 ( .A(n2658), .ZN(n2753) );
  NAND2_X1 U34810 ( .A1(n2753), .A2(n4384), .ZN(n3854) );
  NAND2_X1 U3482 ( .A1(n4385), .A2(n3981), .ZN(n2688) );
  NAND2_X2 U34830 ( .A1(n3854), .A2(n2688), .ZN(n4231) );
  NAND2_X1 U3484 ( .A1(n2349), .A2(IR_REG_31__SCAN_IN), .ZN(n2689) );
  MUX2_X1 U34850 ( .A(IR_REG_31__SCAN_IN), .B(n2689), .S(IR_REG_28__SCAN_IN), 
        .Z(n2690) );
  NOR2_X1 U3486 ( .A1(n2692), .A2(n2691), .ZN(n2821) );
  AND2_X1 U34870 ( .A1(n2821), .A2(B_REG_SCAN_IN), .ZN(n2693) );
  NOR2_X1 U3488 ( .A1(n4304), .A2(n2693), .ZN(n4084) );
  INV_X1 U34890 ( .A(REG2_REG_30__SCAN_IN), .ZN(n2696) );
  NAND2_X1 U3490 ( .A1(n2414), .A2(REG1_REG_30__SCAN_IN), .ZN(n2695) );
  NAND2_X1 U34910 ( .A1(n2413), .A2(REG0_REG_30__SCAN_IN), .ZN(n2694) );
  OAI211_X1 U3492 ( .C1(n2393), .C2(n2696), .A(n2695), .B(n2694), .ZN(n3986)
         );
  INV_X1 U34930 ( .A(n2770), .ZN(n2855) );
  INV_X1 U3494 ( .A(n3844), .ZN(n2736) );
  INV_X1 U34950 ( .A(n3981), .ZN(n2697) );
  INV_X1 U3496 ( .A(n4384), .ZN(n2875) );
  AOI22_X1 U34970 ( .A1(n3987), .A2(n2048), .B1(n2736), .B2(n4324), .ZN(n2698)
         );
  OAI211_X1 U3498 ( .C1(n3569), .C2(n4551), .A(n3562), .B(n2698), .ZN(n2744)
         );
  INV_X1 U34990 ( .A(n2700), .ZN(n2701) );
  NAND2_X1 U3500 ( .A1(n2713), .A2(B_REG_SCAN_IN), .ZN(n2708) );
  NAND2_X1 U35010 ( .A1(n2715), .A2(n2716), .ZN(n2706) );
  MUX2_X1 U3502 ( .A(n2708), .B(B_REG_SCAN_IN), .S(n2714), .Z(n2712) );
  NAND2_X1 U35030 ( .A1(n2703), .A2(IR_REG_31__SCAN_IN), .ZN(n2709) );
  MUX2_X1 U3504 ( .A(IR_REG_31__SCAN_IN), .B(n2709), .S(IR_REG_26__SCAN_IN), 
        .Z(n2711) );
  NAND2_X1 U35050 ( .A1(n2730), .A2(n2766), .ZN(n2923) );
  INV_X1 U35060 ( .A(n4382), .ZN(n2731) );
  NAND2_X1 U35070 ( .A1(n2713), .A2(n2731), .ZN(n2851) );
  NAND2_X1 U35080 ( .A1(n2923), .A2(n2851), .ZN(n2729) );
  NAND2_X1 U35090 ( .A1(n2658), .A2(n4078), .ZN(n2854) );
  NAND2_X1 U35100 ( .A1(n2854), .A2(n2770), .ZN(n2858) );
  OR2_X1 U35110 ( .A1(n4540), .A2(n4384), .ZN(n2717) );
  AND2_X1 U35120 ( .A1(n2924), .A2(n2717), .ZN(n2728) );
  NOR4_X1 U35130 ( .A1(D_REG_18__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_20__SCAN_IN), .A4(D_REG_21__SCAN_IN), .ZN(n2721) );
  NOR4_X1 U35140 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_15__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n2720) );
  NOR4_X1 U35150 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2719) );
  NOR4_X1 U35160 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_23__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_25__SCAN_IN), .ZN(n2718) );
  NAND4_X1 U35170 ( .A1(n2721), .A2(n2720), .A3(n2719), .A4(n2718), .ZN(n2727)
         );
  NOR2_X1 U35180 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_3__SCAN_IN), .ZN(n2725) );
  NOR4_X1 U35190 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_4__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2724) );
  NOR4_X1 U35200 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(
        D_REG_12__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2723) );
  NOR4_X1 U35210 ( .A1(D_REG_6__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_8__SCAN_IN), .A4(D_REG_9__SCAN_IN), .ZN(n2722) );
  NAND4_X1 U35220 ( .A1(n2725), .A2(n2724), .A3(n2723), .A4(n2722), .ZN(n2726)
         );
  OAI21_X1 U35230 ( .B1(n2727), .B2(n2726), .A(n2730), .ZN(n2852) );
  INV_X1 U35240 ( .A(D_REG_0__SCAN_IN), .ZN(n2764) );
  NAND2_X1 U35250 ( .A1(n2730), .A2(n2764), .ZN(n2734) );
  INV_X1 U35260 ( .A(n2714), .ZN(n2732) );
  NAND2_X1 U35270 ( .A1(n2732), .A2(n2731), .ZN(n2733) );
  MUX2_X1 U35280 ( .A(REG0_REG_29__SCAN_IN), .B(n2744), .S(n4559), .Z(n2735)
         );
  INV_X1 U35290 ( .A(n2735), .ZN(n2742) );
  NAND2_X1 U35300 ( .A1(n2993), .A2(n2961), .ZN(n3050) );
  NAND2_X1 U35310 ( .A1(n3241), .A2(n3258), .ZN(n3168) );
  NAND2_X1 U35320 ( .A1(n3464), .A2(n3733), .ZN(n3482) );
  INV_X1 U35330 ( .A(n4094), .ZN(n2737) );
  NAND2_X1 U35340 ( .A1(n2737), .A2(n2736), .ZN(n2738) );
  NAND2_X1 U35350 ( .A1(n4244), .A2(n2738), .ZN(n3564) );
  NAND2_X1 U35360 ( .A1(n2742), .A2(n2741), .ZN(U3515) );
  MUX2_X1 U35370 ( .A(REG1_REG_29__SCAN_IN), .B(n2744), .S(n4568), .Z(n2745)
         );
  INV_X1 U35380 ( .A(n2745), .ZN(n2748) );
  NAND2_X1 U35390 ( .A1(n2740), .A2(n2746), .ZN(n2747) );
  NAND2_X1 U35400 ( .A1(n2748), .A2(n2747), .ZN(U3547) );
  INV_X1 U35410 ( .A(DATAI_22_), .ZN(n4571) );
  NAND2_X1 U35420 ( .A1(n3981), .A2(STATE_REG_SCAN_IN), .ZN(n2749) );
  OAI21_X1 U35430 ( .B1(STATE_REG_SCAN_IN), .B2(n4571), .A(n2749), .ZN(U3330)
         );
  NAND2_X1 U35440 ( .A1(n2821), .A2(STATE_REG_SCAN_IN), .ZN(n2750) );
  OAI21_X1 U35450 ( .B1(STATE_REG_SCAN_IN), .B2(n2353), .A(n2750), .ZN(U3325)
         );
  INV_X1 U35460 ( .A(DATAI_24_), .ZN(n2752) );
  NAND2_X1 U35470 ( .A1(n2714), .A2(STATE_REG_SCAN_IN), .ZN(n2751) );
  OAI21_X1 U35480 ( .B1(STATE_REG_SCAN_IN), .B2(n2752), .A(n2751), .ZN(U3328)
         );
  NAND2_X1 U35490 ( .A1(n2753), .A2(STATE_REG_SCAN_IN), .ZN(n2754) );
  OAI21_X1 U35500 ( .B1(STATE_REG_SCAN_IN), .B2(n2610), .A(n2754), .ZN(U3332)
         );
  INV_X1 U35510 ( .A(DATAI_29_), .ZN(n4584) );
  NAND2_X1 U35520 ( .A1(n2755), .A2(STATE_REG_SCAN_IN), .ZN(n2756) );
  OAI21_X1 U35530 ( .B1(STATE_REG_SCAN_IN), .B2(n4584), .A(n2756), .ZN(U3323)
         );
  INV_X1 U35540 ( .A(DATAI_30_), .ZN(n4718) );
  NAND2_X1 U35550 ( .A1(n2341), .A2(STATE_REG_SCAN_IN), .ZN(n2757) );
  OAI21_X1 U35560 ( .B1(STATE_REG_SCAN_IN), .B2(n4718), .A(n2757), .ZN(U3322)
         );
  INV_X1 U35570 ( .A(DATAI_31_), .ZN(n4637) );
  OR4_X1 U35580 ( .A1(n2339), .A2(IR_REG_30__SCAN_IN), .A3(n2758), .A4(U3149), 
        .ZN(n2759) );
  OAI21_X1 U35590 ( .B1(STATE_REG_SCAN_IN), .B2(n4637), .A(n2759), .ZN(U3321)
         );
  INV_X1 U35600 ( .A(n2879), .ZN(n2881) );
  NAND2_X1 U35610 ( .A1(n2881), .A2(STATE_REG_SCAN_IN), .ZN(n2760) );
  OAI21_X1 U35620 ( .B1(STATE_REG_SCAN_IN), .B2(n2638), .A(n2760), .ZN(U3324)
         );
  NOR3_X1 U35630 ( .A1(n2762), .A2(n2714), .A3(n4382), .ZN(n2763) );
  AOI21_X1 U35640 ( .B1(n4520), .B2(n2764), .A(n2763), .ZN(U3458) );
  INV_X1 U35650 ( .A(n2851), .ZN(n2765) );
  AOI22_X1 U35660 ( .A1(n4520), .A2(n2766), .B1(n2765), .B2(n4521), .ZN(U3459)
         );
  INV_X1 U35670 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4560) );
  AOI21_X1 U35680 ( .B1(n2821), .B2(n2780), .A(n2879), .ZN(n2823) );
  OAI21_X1 U35690 ( .B1(n2821), .B2(REG1_REG_0__SCAN_IN), .A(n2823), .ZN(n2767) );
  MUX2_X1 U35700 ( .A(n2767), .B(n2823), .S(IR_REG_0__SCAN_IN), .Z(n2778) );
  INV_X1 U35710 ( .A(n2876), .ZN(n2768) );
  OR2_X1 U35720 ( .A1(n2769), .A2(U3149), .ZN(n3983) );
  NAND2_X1 U35730 ( .A1(n2768), .A2(n3983), .ZN(n2774) );
  AND2_X1 U35740 ( .A1(n2770), .A2(n2769), .ZN(n2771) );
  NOR2_X1 U35750 ( .A1(n2771), .A2(n2427), .ZN(n2772) );
  AND2_X1 U35760 ( .A1(n2774), .A2(n2772), .ZN(n2796) );
  INV_X1 U35770 ( .A(n2796), .ZN(n2777) );
  INV_X1 U35780 ( .A(n2821), .ZN(n2783) );
  NAND3_X1 U35790 ( .A1(n4495), .A2(IR_REG_0__SCAN_IN), .A3(n4560), .ZN(n2776)
         );
  INV_X1 U35800 ( .A(n2772), .ZN(n2773) );
  AOI22_X1 U35810 ( .A1(n4493), .A2(ADDR_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n2775) );
  OAI211_X1 U3582 ( .C1(n2778), .C2(n2777), .A(n2776), .B(n2775), .ZN(U3240)
         );
  INV_X1 U3583 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2779) );
  NAND2_X1 U3584 ( .A1(n4393), .A2(REG2_REG_1__SCAN_IN), .ZN(n2842) );
  MUX2_X1 U3585 ( .A(n2392), .B(REG2_REG_2__SCAN_IN), .S(n4392), .Z(n2841) );
  AOI21_X1 U3586 ( .B1(n4008), .B2(n2842), .A(n2841), .ZN(n2840) );
  AOI21_X1 U3587 ( .B1(n2049), .B2(REG2_REG_2__SCAN_IN), .A(n2840), .ZN(n2781)
         );
  INV_X1 U3588 ( .A(n4391), .ZN(n2790) );
  XNOR2_X1 U3589 ( .A(n2781), .B(n2790), .ZN(n4021) );
  OAI22_X1 U3590 ( .A1(n4021), .A2(n2936), .B1(n2781), .B2(n2790), .ZN(n2782)
         );
  INV_X1 U3591 ( .A(n4390), .ZN(n2831) );
  XNOR2_X1 U3592 ( .A(n2782), .B(n2831), .ZN(n2824) );
  MUX2_X1 U3593 ( .A(REG2_REG_5__SCAN_IN), .B(n2431), .S(n2801), .Z(n2784) );
  NOR2_X1 U3594 ( .A1(n2879), .A2(n2783), .ZN(n3978) );
  AOI211_X1 U3595 ( .C1(n2785), .C2(n2784), .A(n4489), .B(n2802), .ZN(n2800)
         );
  INV_X1 U3596 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2786) );
  XNOR2_X1 U3597 ( .A(n2049), .B(n2786), .ZN(n2839) );
  INV_X1 U3598 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2787) );
  AND2_X1 U3599 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n4012)
         );
  NAND2_X1 U3600 ( .A1(n4393), .A2(REG1_REG_1__SCAN_IN), .ZN(n2788) );
  NAND2_X1 U3601 ( .A1(n2839), .A2(n2838), .ZN(n2837) );
  NAND2_X1 U3602 ( .A1(n2049), .A2(REG1_REG_2__SCAN_IN), .ZN(n2789) );
  NAND2_X1 U3603 ( .A1(n4020), .A2(REG1_REG_3__SCAN_IN), .ZN(n4019) );
  NAND2_X1 U3604 ( .A1(n2791), .A2(n4391), .ZN(n2792) );
  XNOR2_X1 U3605 ( .A(n2793), .B(n2831), .ZN(n2827) );
  XOR2_X1 U3606 ( .A(REG1_REG_5__SCAN_IN), .B(n2801), .Z(n2794) );
  INV_X1 U3607 ( .A(n4495), .ZN(n2904) );
  AOI211_X1 U3608 ( .C1(n2795), .C2(n2794), .A(n2804), .B(n2904), .ZN(n2799)
         );
  NOR2_X1 U3609 ( .A1(STATE_REG_SCAN_IN), .A2(n2433), .ZN(n3115) );
  AOI21_X1 U3610 ( .B1(n4493), .B2(ADDR_REG_5__SCAN_IN), .A(n3115), .ZN(n2797)
         );
  OAI21_X1 U3611 ( .B1(n4499), .B2(n2801), .A(n2797), .ZN(n2798) );
  OR3_X1 U3612 ( .A1(n2800), .A2(n2799), .A3(n2798), .ZN(U3245) );
  NOR2_X1 U3613 ( .A1(n4493), .A2(n4000), .ZN(U3148) );
  INV_X1 U3614 ( .A(n2801), .ZN(n4389) );
  XNOR2_X1 U3615 ( .A(n2898), .B(REG2_REG_6__SCAN_IN), .ZN(n2810) );
  INV_X1 U3616 ( .A(n4499), .ZN(n4018) );
  NAND2_X1 U3617 ( .A1(n4493), .A2(ADDR_REG_6__SCAN_IN), .ZN(n2803) );
  NAND2_X1 U3618 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3132) );
  NAND2_X1 U3619 ( .A1(n2803), .A2(n3132), .ZN(n2808) );
  INV_X1 U3620 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2805) );
  AOI211_X1 U3621 ( .C1(n2806), .C2(n2805), .A(n2904), .B(n2894), .ZN(n2807)
         );
  AOI211_X1 U3622 ( .C1(n4018), .C2(n4388), .A(n2808), .B(n2807), .ZN(n2809)
         );
  OAI21_X1 U3623 ( .B1(n2810), .B2(n4489), .A(n2809), .ZN(U3246) );
  INV_X1 U3624 ( .A(n2812), .ZN(n2813) );
  OAI22_X1 U3625 ( .A1(n3645), .A2(n3001), .B1(n2968), .B2(n2131), .ZN(n2814)
         );
  NAND2_X1 U3626 ( .A1(n2816), .A2(n2815), .ZN(n2819) );
  INV_X1 U3627 ( .A(n3645), .ZN(n3189) );
  OAI21_X1 U3628 ( .B1(n2968), .B2(n4560), .A(n2866), .ZN(n2818) );
  OAI21_X1 U3629 ( .B1(n2819), .B2(n2818), .A(n2867), .ZN(n2888) );
  NAND2_X1 U3630 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n4007) );
  AOI21_X1 U3631 ( .B1(n2821), .B2(n4007), .A(n2879), .ZN(n2820) );
  OAI21_X1 U3632 ( .B1(n2888), .B2(n2821), .A(n2820), .ZN(n2822) );
  OAI211_X1 U3633 ( .C1(IR_REG_0__SCAN_IN), .C2(n2823), .A(n2822), .B(U4043), 
        .ZN(n2850) );
  XOR2_X1 U3634 ( .A(REG2_REG_4__SCAN_IN), .B(n2824), .Z(n2833) );
  INV_X1 U3635 ( .A(n2825), .ZN(n2826) );
  OAI211_X1 U3636 ( .C1(REG1_REG_4__SCAN_IN), .C2(n2827), .A(n4495), .B(n2826), 
        .ZN(n2830) );
  NAND2_X1 U3637 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n3019) );
  INV_X1 U3638 ( .A(n3019), .ZN(n2828) );
  AOI21_X1 U3639 ( .B1(n4493), .B2(ADDR_REG_4__SCAN_IN), .A(n2828), .ZN(n2829)
         );
  OAI211_X1 U3640 ( .C1(n4499), .C2(n2831), .A(n2830), .B(n2829), .ZN(n2832)
         );
  AOI21_X1 U3641 ( .B1(n4440), .B2(n2833), .A(n2832), .ZN(n2834) );
  NAND2_X1 U3642 ( .A1(n2850), .A2(n2834), .ZN(U3244) );
  NAND2_X1 U3643 ( .A1(n4493), .A2(ADDR_REG_2__SCAN_IN), .ZN(n2835) );
  OAI21_X1 U3644 ( .B1(STATE_REG_SCAN_IN), .B2(n2836), .A(n2835), .ZN(n2848)
         );
  OAI211_X1 U3645 ( .C1(n2839), .C2(n2838), .A(n4495), .B(n2837), .ZN(n2846)
         );
  INV_X1 U3646 ( .A(n2840), .ZN(n2844) );
  NAND3_X1 U3647 ( .A1(n4008), .A2(n2842), .A3(n2841), .ZN(n2843) );
  NAND3_X1 U3648 ( .A1(n4440), .A2(n2844), .A3(n2843), .ZN(n2845) );
  NAND2_X1 U3649 ( .A1(n2846), .A2(n2845), .ZN(n2847) );
  AOI211_X1 U3650 ( .C1(n2049), .C2(n4018), .A(n2848), .B(n2847), .ZN(n2849)
         );
  NAND2_X1 U3651 ( .A1(n2850), .A2(n2849), .ZN(U3242) );
  AND2_X1 U3652 ( .A1(n2852), .A2(n2851), .ZN(n2925) );
  INV_X1 U3653 ( .A(n2884), .ZN(n2862) );
  NAND2_X1 U3654 ( .A1(n2854), .A2(n2998), .ZN(n2856) );
  NAND2_X1 U3655 ( .A1(n2856), .A2(n2855), .ZN(n2869) );
  NAND2_X1 U3656 ( .A1(n2869), .A2(n3539), .ZN(n2857) );
  NAND2_X1 U3657 ( .A1(n2862), .A2(n2857), .ZN(n2859) );
  NAND2_X1 U3658 ( .A1(n2859), .A2(n2858), .ZN(n2970) );
  INV_X1 U3659 ( .A(n2970), .ZN(n2863) );
  NAND2_X1 U3660 ( .A1(n4078), .A2(n3981), .ZN(n2864) );
  INV_X1 U3661 ( .A(n2864), .ZN(n2860) );
  NAND2_X1 U3662 ( .A1(n2860), .A2(n4521), .ZN(n2861) );
  INV_X1 U3663 ( .A(n2882), .ZN(n3979) );
  NAND2_X1 U3664 ( .A1(n2862), .A2(n3979), .ZN(n2971) );
  NAND3_X1 U3665 ( .A1(n2863), .A2(n2876), .A3(n2971), .ZN(n2917) );
  INV_X1 U3666 ( .A(n2917), .ZN(n2892) );
  INV_X1 U3667 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3154) );
  XNOR2_X1 U3668 ( .A(n2865), .B(n3658), .ZN(n2908) );
  XNOR2_X1 U3669 ( .A(n2908), .B(n2909), .ZN(n2873) );
  INV_X1 U3670 ( .A(n2866), .ZN(n2868) );
  OAI21_X1 U3671 ( .B1(n2868), .B2(n3658), .A(n2867), .ZN(n2872) );
  NAND2_X1 U3672 ( .A1(n2873), .A2(n2872), .ZN(n2912) );
  INV_X1 U3673 ( .A(n2869), .ZN(n2870) );
  OAI211_X1 U3674 ( .C1(n2873), .C2(n2872), .A(n2912), .B(n3806), .ZN(n2887)
         );
  AND2_X1 U3675 ( .A1(n2876), .A2(n4324), .ZN(n2874) );
  NAND2_X1 U3676 ( .A1(n2884), .A2(n2874), .ZN(n2878) );
  AND2_X1 U3677 ( .A1(n2876), .A2(n2875), .ZN(n2877) );
  INV_X1 U3678 ( .A(n3779), .ZN(n2976) );
  NOR2_X1 U3679 ( .A1(n2882), .A2(n2879), .ZN(n2880) );
  NOR2_X1 U3680 ( .A1(n2882), .A2(n2881), .ZN(n2883) );
  NAND2_X2 U3681 ( .A1(n2884), .A2(n2883), .ZN(n3813) );
  OAI22_X1 U3682 ( .A1(n3000), .A2(n3808), .B1(n3813), .B2(n2967), .ZN(n2885)
         );
  AOI21_X1 U3683 ( .B1(n3149), .B2(n2976), .A(n2885), .ZN(n2886) );
  OAI211_X1 U3684 ( .C1(n2892), .C2(n3154), .A(n2887), .B(n2886), .ZN(U3219)
         );
  OAI22_X1 U3685 ( .A1(n2888), .A2(n3800), .B1(n3004), .B2(n3813), .ZN(n2889)
         );
  AOI21_X1 U3686 ( .B1(n3150), .B2(n2976), .A(n2889), .ZN(n2890) );
  OAI21_X1 U3687 ( .B1(n2892), .B2(n2891), .A(n2890), .ZN(U3229) );
  INV_X1 U3688 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4566) );
  MUX2_X1 U3689 ( .A(REG1_REG_7__SCAN_IN), .B(n4566), .S(n4387), .Z(n2896) );
  INV_X1 U3690 ( .A(n2893), .ZN(n2895) );
  XOR2_X1 U3691 ( .A(n2896), .B(n2949), .Z(n2905) );
  NAND2_X1 U3692 ( .A1(n4493), .A2(ADDR_REG_7__SCAN_IN), .ZN(n2897) );
  NAND2_X1 U3693 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3194) );
  NAND2_X1 U3694 ( .A1(n2897), .A2(n3194), .ZN(n2902) );
  MUX2_X1 U3695 ( .A(n2457), .B(REG2_REG_7__SCAN_IN), .S(n4387), .Z(n2899) );
  AOI211_X1 U3696 ( .C1(n2900), .C2(n2899), .A(n4489), .B(n2951), .ZN(n2901)
         );
  AOI211_X1 U3697 ( .C1(n4018), .C2(n4387), .A(n2902), .B(n2901), .ZN(n2903)
         );
  OAI21_X1 U3698 ( .B1(n2905), .B2(n2904), .A(n2903), .ZN(U3247) );
  OAI22_X1 U3699 ( .A1(n2967), .A2(n3645), .B1(n3657), .B2(n2992), .ZN(n2906)
         );
  XNOR2_X1 U3700 ( .A(n2906), .B(n3658), .ZN(n2963) );
  OAI22_X1 U3701 ( .A1(n2967), .A2(n2907), .B1(n3645), .B2(n2992), .ZN(n2962)
         );
  XNOR2_X1 U3702 ( .A(n2963), .B(n2962), .ZN(n2914) );
  NAND2_X1 U3703 ( .A1(n2912), .A2(n2911), .ZN(n2913) );
  AOI21_X1 U3704 ( .B1(n2914), .B2(n2913), .A(n2964), .ZN(n2919) );
  INV_X1 U3705 ( .A(n3813), .ZN(n3792) );
  INV_X1 U3706 ( .A(n3808), .ZN(n3794) );
  AOI22_X1 U3707 ( .A1(n3792), .A2(n4004), .B1(n3794), .B2(n2387), .ZN(n2915)
         );
  OAI21_X1 U3708 ( .B1(n3779), .B2(n2992), .A(n2915), .ZN(n2916) );
  AOI21_X1 U3709 ( .B1(REG3_REG_2__SCAN_IN), .B2(n2917), .A(n2916), .ZN(n2918)
         );
  OAI21_X1 U3710 ( .B1(n2919), .B2(n3800), .A(n2918), .ZN(U3234) );
  NAND2_X1 U3711 ( .A1(n2920), .A2(n2921), .ZN(n2922) );
  XNOR2_X1 U3712 ( .A(n2922), .B(n3893), .ZN(n2940) );
  NAND4_X1 U3713 ( .A1(n2926), .A2(n2925), .A3(n2924), .A4(n2923), .ZN(n2927)
         );
  OR2_X1 U3714 ( .A1(n2812), .A2(n4078), .ZN(n3041) );
  INV_X1 U3715 ( .A(n3041), .ZN(n2928) );
  NAND2_X1 U3716 ( .A1(n4213), .A2(n2928), .ZN(n4238) );
  XNOR2_X1 U3717 ( .A(n2929), .B(n3893), .ZN(n2932) );
  AOI22_X1 U3718 ( .A1(n4005), .A2(n2048), .B1(n4324), .B2(n2977), .ZN(n2930)
         );
  OAI21_X1 U3719 ( .B1(n3117), .B2(n4304), .A(n2930), .ZN(n2931) );
  AOI21_X1 U3720 ( .B1(n2932), .B2(n4231), .A(n2931), .ZN(n2933) );
  OAI21_X1 U3721 ( .B1(n2940), .B2(n4227), .A(n2933), .ZN(n2941) );
  NAND2_X1 U3722 ( .A1(n2941), .A2(n4213), .ZN(n2939) );
  NAND2_X1 U3723 ( .A1(n4213), .A2(n4078), .ZN(n3485) );
  INV_X1 U3724 ( .A(n2993), .ZN(n2934) );
  NAND2_X1 U3725 ( .A1(n2934), .A2(n2977), .ZN(n2935) );
  AND2_X1 U3726 ( .A1(n2935), .A2(n3050), .ZN(n2944) );
  OAI22_X1 U3727 ( .A1(n4213), .A2(n2936), .B1(REG3_REG_3__SCAN_IN), .B2(n4500), .ZN(n2937) );
  AOI21_X1 U3728 ( .B1(n4513), .B2(n2944), .A(n2937), .ZN(n2938) );
  OAI211_X1 U3729 ( .C1(n2940), .C2(n4238), .A(n2939), .B(n2938), .ZN(U3287)
         );
  INV_X1 U3730 ( .A(n2940), .ZN(n2942) );
  AOI21_X1 U3731 ( .B1(n4548), .B2(n2942), .A(n2941), .ZN(n2946) );
  AOI22_X1 U3732 ( .A1(n2739), .A2(n2944), .B1(REG0_REG_3__SCAN_IN), .B2(n4557), .ZN(n2943) );
  OAI21_X1 U3733 ( .B1(n2946), .B2(n4557), .A(n2943), .ZN(U3473) );
  AOI22_X1 U3734 ( .A1(n2746), .A2(n2944), .B1(REG1_REG_3__SCAN_IN), .B2(n4565), .ZN(n2945) );
  OAI21_X1 U3735 ( .B1(n2946), .B2(n4565), .A(n2945), .ZN(U3521) );
  NOR2_X1 U3736 ( .A1(n4387), .A2(REG1_REG_7__SCAN_IN), .ZN(n2948) );
  INV_X1 U3737 ( .A(n4387), .ZN(n2947) );
  XNOR2_X1 U3738 ( .A(n4051), .B(n4050), .ZN(n4052) );
  XOR2_X1 U3739 ( .A(REG1_REG_8__SCAN_IN), .B(n4052), .Z(n2950) );
  NAND2_X1 U3740 ( .A1(n2950), .A2(n4495), .ZN(n2956) );
  XNOR2_X1 U3741 ( .A(REG2_REG_8__SCAN_IN), .B(n4029), .ZN(n2952) );
  NAND2_X1 U3742 ( .A1(n4440), .A2(n2952), .ZN(n2953) );
  NAND2_X1 U3743 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3225) );
  NAND2_X1 U3744 ( .A1(n2953), .A2(n3225), .ZN(n2954) );
  AOI21_X1 U3745 ( .B1(n4493), .B2(ADDR_REG_8__SCAN_IN), .A(n2954), .ZN(n2955)
         );
  OAI211_X1 U3746 ( .C1(n4499), .C2(n4050), .A(n2956), .B(n2955), .ZN(U3248)
         );
  NAND2_X1 U3747 ( .A1(n4004), .A2(n3189), .ZN(n2958) );
  NAND2_X1 U3748 ( .A1(n2977), .A2(n3649), .ZN(n2957) );
  NAND2_X1 U3749 ( .A1(n2958), .A2(n2957), .ZN(n2959) );
  XNOR2_X1 U3750 ( .A(n2959), .B(n3658), .ZN(n3013) );
  OAI22_X1 U3751 ( .A1(n3018), .A2(n2907), .B1(n3645), .B2(n2961), .ZN(n3012)
         );
  XNOR2_X1 U3752 ( .A(n3013), .B(n3012), .ZN(n3014) );
  INV_X1 U3753 ( .A(n2962), .ZN(n2966) );
  INV_X1 U3754 ( .A(n2963), .ZN(n2965) );
  XOR2_X1 U3755 ( .A(n3014), .B(n2093), .Z(n2979) );
  OAI22_X1 U3756 ( .A1(n2967), .A2(n3808), .B1(n3813), .B2(n3117), .ZN(n2975)
         );
  INV_X1 U3757 ( .A(n2968), .ZN(n2969) );
  OAI21_X1 U3758 ( .B1(n2970), .B2(n2969), .A(STATE_REG_SCAN_IN), .ZN(n2973)
         );
  AND2_X1 U3759 ( .A1(n2971), .A2(n3983), .ZN(n2972) );
  MUX2_X1 U3760 ( .A(n3793), .B(U3149), .S(REG3_REG_3__SCAN_IN), .Z(n2974) );
  AOI211_X1 U3761 ( .C1(n2977), .C2(n2976), .A(n2975), .B(n2974), .ZN(n2978)
         );
  OAI21_X1 U3762 ( .B1(n2979), .B2(n3800), .A(n2978), .ZN(U3215) );
  INV_X1 U3763 ( .A(n2920), .ZN(n2980) );
  AOI21_X1 U3764 ( .B1(n3894), .B2(n2981), .A(n2980), .ZN(n2986) );
  INV_X1 U3765 ( .A(n2986), .ZN(n4515) );
  OAI21_X1 U3766 ( .B1(n3894), .B2(n2983), .A(n2982), .ZN(n2989) );
  AOI22_X1 U3767 ( .A1(n2387), .A2(n2048), .B1(n2984), .B2(n4324), .ZN(n2985)
         );
  OAI21_X1 U3768 ( .B1(n3018), .B2(n4304), .A(n2985), .ZN(n2988) );
  NOR2_X1 U3769 ( .A1(n2986), .A2(n4227), .ZN(n2987) );
  AOI211_X1 U3770 ( .C1(n4231), .C2(n2989), .A(n2988), .B(n2987), .ZN(n4518)
         );
  INV_X1 U3771 ( .A(n4518), .ZN(n2990) );
  AOI21_X1 U3772 ( .B1(n4548), .B2(n4515), .A(n2990), .ZN(n2997) );
  INV_X1 U3773 ( .A(n2991), .ZN(n3148) );
  NOR2_X1 U3774 ( .A1(n3148), .A2(n2992), .ZN(n2994) );
  NOR2_X1 U3775 ( .A1(n2994), .A2(n2993), .ZN(n4512) );
  AOI22_X1 U3776 ( .A1(n2746), .A2(n4512), .B1(REG1_REG_2__SCAN_IN), .B2(n4565), .ZN(n2995) );
  OAI21_X1 U3777 ( .B1(n2997), .B2(n4565), .A(n2995), .ZN(U3520) );
  AOI22_X1 U3778 ( .A1(n2739), .A2(n4512), .B1(REG0_REG_2__SCAN_IN), .B2(n4557), .ZN(n2996) );
  OAI21_X1 U3779 ( .B1(n2997), .B2(n4557), .A(n2996), .ZN(U3471) );
  INV_X1 U3780 ( .A(n2998), .ZN(n2999) );
  NOR2_X1 U3781 ( .A1(n3001), .A2(n2999), .ZN(n4537) );
  INV_X1 U3782 ( .A(n4227), .ZN(n3002) );
  NAND2_X1 U3783 ( .A1(n2817), .A2(n3001), .ZN(n3914) );
  NAND2_X1 U3784 ( .A1(n3912), .A2(n3914), .ZN(n4538) );
  OAI21_X1 U3785 ( .B1(n3002), .B2(n4231), .A(n4538), .ZN(n3003) );
  OAI21_X1 U3786 ( .B1(n3004), .B2(n4304), .A(n3003), .ZN(n4536) );
  AOI21_X1 U3787 ( .B1(n4537), .B2(n3005), .A(n4536), .ZN(n3008) );
  AOI22_X1 U3788 ( .A1(n4519), .A2(REG2_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(n4511), .ZN(n3007) );
  INV_X1 U3789 ( .A(n4238), .ZN(n4514) );
  NAND2_X1 U3790 ( .A1(n4514), .A2(n4538), .ZN(n3006) );
  OAI211_X1 U3791 ( .C1(n3008), .C2(n4519), .A(n3007), .B(n3006), .ZN(U3290)
         );
  AOI22_X1 U3792 ( .A1(n4003), .A2(n2960), .B1(n3189), .B2(n3051), .ZN(n3105)
         );
  NAND2_X1 U3793 ( .A1(n4003), .A2(n3641), .ZN(n3010) );
  NAND2_X1 U3794 ( .A1(n3051), .A2(n3649), .ZN(n3009) );
  NAND2_X1 U3795 ( .A1(n3010), .A2(n3009), .ZN(n3011) );
  XNOR2_X1 U3796 ( .A(n3011), .B(n3658), .ZN(n3104) );
  XOR2_X1 U3797 ( .A(n3105), .B(n3104), .Z(n3016) );
  AOI211_X1 U3798 ( .C1(n3016), .C2(n3015), .A(n3800), .B(n3108), .ZN(n3017)
         );
  INV_X1 U3799 ( .A(n3017), .ZN(n3023) );
  OAI22_X1 U3800 ( .A1(n3779), .A2(n3056), .B1(n3018), .B2(n3808), .ZN(n3021)
         );
  OAI21_X1 U3801 ( .B1(n3813), .B2(n3130), .A(n3019), .ZN(n3020) );
  NOR2_X1 U3802 ( .A1(n3021), .A2(n3020), .ZN(n3022) );
  OAI211_X1 U3803 ( .C1(n3819), .C2(n3052), .A(n3023), .B(n3022), .ZN(U3227)
         );
  AND2_X1 U3804 ( .A1(n2091), .A2(n3927), .ZN(n3890) );
  XNOR2_X1 U3805 ( .A(n3024), .B(n3890), .ZN(n3102) );
  XOR2_X1 U3806 ( .A(n3890), .B(n3025), .Z(n3026) );
  NAND2_X1 U3807 ( .A1(n3026), .A2(n4231), .ZN(n3099) );
  AOI22_X1 U3808 ( .A1(n4001), .A2(n4325), .B1(n4324), .B2(n3027), .ZN(n3028)
         );
  OAI211_X1 U3809 ( .C1(n3117), .C2(n4328), .A(n3099), .B(n3028), .ZN(n3029)
         );
  AOI21_X1 U3810 ( .B1(n3102), .B2(n4316), .A(n3029), .ZN(n3033) );
  OR2_X1 U3811 ( .A1(n3049), .A2(n3114), .ZN(n3030) );
  AND2_X1 U3812 ( .A1(n3077), .A2(n3030), .ZN(n3093) );
  AOI22_X1 U3813 ( .A1(n3093), .A2(n2746), .B1(REG1_REG_5__SCAN_IN), .B2(n4565), .ZN(n3031) );
  OAI21_X1 U3814 ( .B1(n3033), .B2(n4565), .A(n3031), .ZN(U3523) );
  AOI22_X1 U3815 ( .A1(n3093), .A2(n2739), .B1(REG0_REG_5__SCAN_IN), .B2(n4557), .ZN(n3032) );
  OAI21_X1 U3816 ( .B1(n3033), .B2(n4557), .A(n3032), .ZN(U3477) );
  XOR2_X1 U3817 ( .A(n3896), .B(n3034), .Z(n3037) );
  INV_X1 U3818 ( .A(n4231), .ZN(n3408) );
  OAI22_X1 U3819 ( .A1(n3257), .A2(n4304), .B1(n3539), .B2(n3193), .ZN(n3035)
         );
  AOI21_X1 U3820 ( .B1(n2048), .B2(n4001), .A(n3035), .ZN(n3036) );
  OAI21_X1 U3821 ( .B1(n3037), .B2(n3408), .A(n3036), .ZN(n4553) );
  INV_X1 U3822 ( .A(n4553), .ZN(n3048) );
  INV_X1 U3823 ( .A(n3485), .ZN(n3046) );
  NAND2_X1 U3824 ( .A1(n3075), .A2(n3188), .ZN(n3038) );
  NAND2_X1 U3825 ( .A1(n3038), .A2(n2811), .ZN(n3039) );
  NOR2_X1 U3826 ( .A1(n3239), .A2(n3039), .ZN(n4554) );
  OAI22_X1 U3827 ( .A1(n4213), .A2(n2457), .B1(n3199), .B2(n4500), .ZN(n3045)
         );
  INV_X1 U3828 ( .A(n4555), .ZN(n3043) );
  AND2_X1 U3829 ( .A1(n3040), .A2(n3896), .ZN(n4552) );
  NAND2_X1 U3830 ( .A1(n4227), .A2(n3041), .ZN(n3042) );
  NOR3_X1 U3831 ( .A1(n3043), .A2(n4552), .A3(n4198), .ZN(n3044) );
  AOI211_X1 U3832 ( .C1(n3046), .C2(n4554), .A(n3045), .B(n3044), .ZN(n3047)
         );
  OAI21_X1 U3833 ( .B1(n4519), .B2(n3048), .A(n3047), .ZN(U3283) );
  AOI211_X1 U3834 ( .C1(n3051), .C2(n3050), .A(n3481), .B(n3049), .ZN(n4547)
         );
  NOR2_X1 U3835 ( .A1(n4500), .A2(n3052), .ZN(n3066) );
  XOR2_X1 U3836 ( .A(n3053), .B(n3054), .Z(n3065) );
  NAND2_X1 U3837 ( .A1(n4004), .A2(n2048), .ZN(n3055) );
  OAI21_X1 U3838 ( .B1(n3539), .B2(n3056), .A(n3055), .ZN(n3063) );
  AND2_X1 U3839 ( .A1(n3058), .A2(n3057), .ZN(n3059) );
  OR2_X1 U3840 ( .A1(n3059), .A2(n3053), .ZN(n3061) );
  NAND2_X1 U3841 ( .A1(n3059), .A2(n3053), .ZN(n3060) );
  NAND2_X1 U3842 ( .A1(n3061), .A2(n3060), .ZN(n3067) );
  NOR2_X1 U3843 ( .A1(n3067), .A2(n4227), .ZN(n3062) );
  AOI211_X1 U3844 ( .C1(n4325), .C2(n4002), .A(n3063), .B(n3062), .ZN(n3064)
         );
  OAI21_X1 U3845 ( .B1(n3408), .B2(n3065), .A(n3064), .ZN(n4546) );
  AOI211_X1 U3846 ( .C1(n4547), .C2(n4078), .A(n3066), .B(n4546), .ZN(n3069)
         );
  INV_X1 U3847 ( .A(n3067), .ZN(n4549) );
  AOI22_X1 U3848 ( .A1(n4549), .A2(n4514), .B1(REG2_REG_4__SCAN_IN), .B2(n4519), .ZN(n3068) );
  OAI21_X1 U3849 ( .B1(n3069), .B2(n4519), .A(n3068), .ZN(U3286) );
  XNOR2_X1 U3850 ( .A(n3070), .B(n3888), .ZN(n3089) );
  XOR2_X1 U3851 ( .A(n3888), .B(n3071), .Z(n3092) );
  OAI22_X1 U3852 ( .A1(n3226), .A2(n4304), .B1(n3131), .B2(n3539), .ZN(n3072)
         );
  AOI21_X1 U3853 ( .B1(n2048), .B2(n4002), .A(n3072), .ZN(n3073) );
  OAI21_X1 U3854 ( .B1(n3092), .B2(n3408), .A(n3073), .ZN(n3074) );
  AOI21_X1 U3855 ( .B1(n3089), .B2(n4316), .A(n3074), .ZN(n3082) );
  INV_X1 U3856 ( .A(n3075), .ZN(n3076) );
  AOI21_X1 U3857 ( .B1(n3083), .B2(n3077), .A(n3076), .ZN(n3088) );
  AOI22_X1 U3858 ( .A1(n3088), .A2(n2746), .B1(n4565), .B2(REG1_REG_6__SCAN_IN), .ZN(n3078) );
  OAI21_X1 U3859 ( .B1(n3082), .B2(n4565), .A(n3078), .ZN(U3524) );
  INV_X1 U3860 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3079) );
  NOR2_X1 U3861 ( .A1(n4559), .A2(n3079), .ZN(n3080) );
  AOI21_X1 U3862 ( .B1(n3088), .B2(n2739), .A(n3080), .ZN(n3081) );
  OAI21_X1 U3863 ( .B1(n3082), .B2(n4557), .A(n3081), .ZN(U3479) );
  NAND2_X1 U3864 ( .A1(n4213), .A2(n4231), .ZN(n3355) );
  NAND2_X1 U3865 ( .A1(n4213), .A2(n4324), .ZN(n4169) );
  INV_X1 U3866 ( .A(n4169), .ZN(n3430) );
  NAND2_X1 U3867 ( .A1(n4213), .A2(n4325), .ZN(n4170) );
  INV_X1 U3868 ( .A(n4170), .ZN(n3429) );
  AOI22_X1 U3869 ( .A1(n3083), .A2(n3430), .B1(n3429), .B2(n3999), .ZN(n3086)
         );
  INV_X1 U3870 ( .A(n3137), .ZN(n3084) );
  AOI22_X1 U3871 ( .A1(n4519), .A2(REG2_REG_6__SCAN_IN), .B1(n3084), .B2(n4511), .ZN(n3085) );
  OAI211_X1 U3872 ( .C1(n3130), .C2(n4167), .A(n3086), .B(n3085), .ZN(n3087)
         );
  AOI21_X1 U3873 ( .B1(n4513), .B2(n3088), .A(n3087), .ZN(n3091) );
  NAND2_X1 U3874 ( .A1(n3089), .A2(n4209), .ZN(n3090) );
  OAI211_X1 U3875 ( .C1(n3092), .C2(n3355), .A(n3091), .B(n3090), .ZN(U3284)
         );
  INV_X1 U3876 ( .A(n3093), .ZN(n3098) );
  OAI22_X1 U3877 ( .A1(n4213), .A2(n2431), .B1(n3122), .B2(n4500), .ZN(n3094)
         );
  AOI21_X1 U3878 ( .B1(n3561), .B2(n4003), .A(n3094), .ZN(n3097) );
  OAI22_X1 U3879 ( .A1(n3192), .A2(n4170), .B1(n4169), .B2(n3114), .ZN(n3095)
         );
  INV_X1 U3880 ( .A(n3095), .ZN(n3096) );
  OAI211_X1 U3881 ( .C1(n4195), .C2(n3098), .A(n3097), .B(n3096), .ZN(n3101)
         );
  NOR2_X1 U3882 ( .A1(n3099), .A2(n4519), .ZN(n3100) );
  AOI211_X1 U3883 ( .C1(n3102), .C2(n4209), .A(n3101), .B(n3100), .ZN(n3103)
         );
  INV_X1 U3884 ( .A(n3103), .ZN(U3285) );
  NOR2_X1 U3885 ( .A1(n3645), .A2(n3114), .ZN(n3109) );
  AOI21_X1 U3886 ( .B1(n4002), .B2(n2960), .A(n3109), .ZN(n3123) );
  OAI22_X1 U3887 ( .A1(n3130), .A2(n3645), .B1(n3657), .B2(n3114), .ZN(n3110)
         );
  XNOR2_X1 U3888 ( .A(n3110), .B(n3658), .ZN(n3125) );
  XOR2_X1 U3889 ( .A(n3123), .B(n3125), .Z(n3111) );
  AOI211_X1 U3890 ( .C1(n3112), .C2(n3111), .A(n3800), .B(n3124), .ZN(n3113)
         );
  INV_X1 U3891 ( .A(n3113), .ZN(n3121) );
  OAI22_X1 U3892 ( .A1(n3779), .A2(n3114), .B1(n3192), .B2(n3813), .ZN(n3119)
         );
  INV_X1 U3893 ( .A(n3115), .ZN(n3116) );
  OAI21_X1 U3894 ( .B1(n3808), .B2(n3117), .A(n3116), .ZN(n3118) );
  NOR2_X1 U3895 ( .A1(n3119), .A2(n3118), .ZN(n3120) );
  OAI211_X1 U3896 ( .C1(n3819), .C2(n3122), .A(n3121), .B(n3120), .ZN(U3224)
         );
  INV_X1 U3897 ( .A(n3123), .ZN(n3126) );
  OAI22_X1 U3898 ( .A1(n3192), .A2(n3645), .B1(n3657), .B2(n3131), .ZN(n3127)
         );
  XNOR2_X1 U3899 ( .A(n3127), .B(n3658), .ZN(n3183) );
  INV_X1 U3900 ( .A(n3184), .ZN(n3185) );
  XNOR2_X1 U3901 ( .A(n3183), .B(n3185), .ZN(n3128) );
  XNOR2_X1 U3902 ( .A(n3186), .B(n3128), .ZN(n3129) );
  NAND2_X1 U3903 ( .A1(n3129), .A2(n3806), .ZN(n3136) );
  OAI22_X1 U3904 ( .A1(n3779), .A2(n3131), .B1(n3130), .B2(n3808), .ZN(n3134)
         );
  OAI21_X1 U3905 ( .B1(n3813), .B2(n3226), .A(n3132), .ZN(n3133) );
  NOR2_X1 U3906 ( .A1(n3134), .A2(n3133), .ZN(n3135) );
  OAI211_X1 U3907 ( .C1(n3819), .C2(n3137), .A(n3136), .B(n3135), .ZN(U3236)
         );
  INV_X1 U3908 ( .A(n3138), .ZN(n3938) );
  AND2_X1 U3909 ( .A1(n3938), .A2(n3936), .ZN(n3891) );
  XOR2_X1 U3910 ( .A(n3891), .B(n3139), .Z(n3140) );
  NAND2_X1 U3911 ( .A1(n3140), .A2(n4231), .ZN(n3176) );
  OR2_X1 U3912 ( .A1(n3241), .A2(n3258), .ZN(n3141) );
  AND2_X1 U3913 ( .A1(n3168), .A2(n3141), .ZN(n3180) );
  AOI22_X1 U3914 ( .A1(n3429), .A2(n3996), .B1(n3561), .B2(n3998), .ZN(n3142)
         );
  OAI21_X1 U3915 ( .B1(n3258), .B2(n4169), .A(n3142), .ZN(n3144) );
  OAI22_X1 U3916 ( .A1(n3264), .A2(n4500), .B1(n2481), .B2(n4213), .ZN(n3143)
         );
  AOI211_X1 U3917 ( .C1(n3180), .C2(n4513), .A(n3144), .B(n3143), .ZN(n3147)
         );
  XNOR2_X1 U3918 ( .A(n3145), .B(n3891), .ZN(n3178) );
  NAND2_X1 U3919 ( .A1(n3178), .A2(n4209), .ZN(n3146) );
  OAI211_X1 U3920 ( .C1(n3176), .C2(n4519), .A(n3147), .B(n3146), .ZN(U3281)
         );
  AOI21_X1 U3921 ( .B1(n3150), .B2(n3149), .A(n3148), .ZN(n4544) );
  OR2_X1 U3922 ( .A1(n2659), .A2(n3151), .ZN(n3152) );
  NAND2_X1 U3923 ( .A1(n3153), .A2(n3152), .ZN(n4541) );
  OAI22_X1 U3924 ( .A1(n4541), .A2(n4238), .B1(n3154), .B2(n4500), .ZN(n3163)
         );
  NAND2_X1 U3925 ( .A1(n2817), .A2(n2048), .ZN(n3156) );
  NAND2_X1 U3926 ( .A1(n4005), .A2(n4325), .ZN(n3155) );
  OAI211_X1 U3927 ( .C1(n3539), .C2(n3157), .A(n3156), .B(n3155), .ZN(n3158)
         );
  INV_X1 U3928 ( .A(n3158), .ZN(n3161) );
  XNOR2_X1 U3929 ( .A(n2659), .B(n3912), .ZN(n3159) );
  NAND2_X1 U3930 ( .A1(n3159), .A2(n4231), .ZN(n3160) );
  OAI211_X1 U3931 ( .C1(n4541), .C2(n4227), .A(n3161), .B(n3160), .ZN(n4542)
         );
  MUX2_X1 U3932 ( .A(n4542), .B(REG2_REG_1__SCAN_IN), .S(n4519), .Z(n3162) );
  AOI211_X1 U3933 ( .C1(n4513), .C2(n4544), .A(n3163), .B(n3162), .ZN(n3164)
         );
  INV_X1 U3934 ( .A(n3164), .ZN(U3289) );
  NAND2_X1 U3935 ( .A1(n3944), .A2(n3940), .ZN(n3886) );
  XNOR2_X1 U3936 ( .A(n3165), .B(n3886), .ZN(n3202) );
  XNOR2_X1 U3937 ( .A(n3166), .B(n3886), .ZN(n3204) );
  NAND2_X1 U3938 ( .A1(n3204), .A2(n4209), .ZN(n3174) );
  AOI21_X1 U3939 ( .B1(n3282), .B2(n3168), .A(n3273), .ZN(n3206) );
  AOI22_X1 U3940 ( .A1(n3430), .A2(n3282), .B1(n3429), .B2(n3995), .ZN(n3171)
         );
  INV_X1 U3941 ( .A(n3295), .ZN(n3169) );
  AOI22_X1 U3942 ( .A1(n4519), .A2(REG2_REG_10__SCAN_IN), .B1(n3169), .B2(
        n4511), .ZN(n3170) );
  OAI211_X1 U3943 ( .C1(n3290), .C2(n4167), .A(n3171), .B(n3170), .ZN(n3172)
         );
  AOI21_X1 U3944 ( .B1(n3206), .B2(n4513), .A(n3172), .ZN(n3173) );
  OAI211_X1 U3945 ( .C1(n3202), .C2(n3355), .A(n3174), .B(n3173), .ZN(U3280)
         );
  AOI22_X1 U3946 ( .A1(n3996), .A2(n4325), .B1(n4324), .B2(n3252), .ZN(n3175)
         );
  OAI211_X1 U3947 ( .C1(n3257), .C2(n4328), .A(n3176), .B(n3175), .ZN(n3177)
         );
  AOI21_X1 U3948 ( .B1(n3178), .B2(n4316), .A(n3177), .ZN(n3182) );
  AOI22_X1 U3949 ( .A1(n3180), .A2(n2746), .B1(REG1_REG_9__SCAN_IN), .B2(n4565), .ZN(n3179) );
  OAI21_X1 U3950 ( .B1(n3182), .B2(n4565), .A(n3179), .ZN(U3527) );
  AOI22_X1 U3951 ( .A1(n3180), .A2(n2739), .B1(REG0_REG_9__SCAN_IN), .B2(n4557), .ZN(n3181) );
  OAI21_X1 U3952 ( .B1(n3182), .B2(n4557), .A(n3181), .ZN(U3485) );
  OAI22_X1 U3953 ( .A1(n3226), .A2(n3645), .B1(n3657), .B2(n3193), .ZN(n3187)
         );
  XOR2_X1 U3954 ( .A(n3658), .B(n3187), .Z(n3210) );
  INV_X1 U3955 ( .A(n3210), .ZN(n3190) );
  AOI22_X1 U3956 ( .A1(n3999), .A2(n2960), .B1(n3189), .B2(n3188), .ZN(n3209)
         );
  XNOR2_X1 U3957 ( .A(n3190), .B(n3209), .ZN(n3212) );
  XOR2_X1 U3958 ( .A(n3213), .B(n3212), .Z(n3191) );
  NAND2_X1 U3959 ( .A1(n3191), .A2(n3806), .ZN(n3198) );
  OAI22_X1 U3960 ( .A1(n3779), .A2(n3193), .B1(n3192), .B2(n3808), .ZN(n3196)
         );
  OAI21_X1 U3961 ( .B1(n3813), .B2(n3257), .A(n3194), .ZN(n3195) );
  NOR2_X1 U3962 ( .A1(n3196), .A2(n3195), .ZN(n3197) );
  OAI211_X1 U3963 ( .C1(n3819), .C2(n3199), .A(n3198), .B(n3197), .ZN(U3210)
         );
  OAI22_X1 U3964 ( .A1(n3455), .A2(n4304), .B1(n3539), .B2(n3289), .ZN(n3200)
         );
  AOI21_X1 U3965 ( .B1(n2048), .B2(n3997), .A(n3200), .ZN(n3201) );
  OAI21_X1 U3966 ( .B1(n3202), .B2(n3408), .A(n3201), .ZN(n3203) );
  AOI21_X1 U3967 ( .B1(n4316), .B2(n3204), .A(n3203), .ZN(n3208) );
  AOI22_X1 U3968 ( .A1(n3206), .A2(n2739), .B1(REG0_REG_10__SCAN_IN), .B2(
        n4557), .ZN(n3205) );
  OAI21_X1 U3969 ( .B1(n3208), .B2(n4557), .A(n3205), .ZN(U3487) );
  AOI22_X1 U3970 ( .A1(n3206), .A2(n2746), .B1(REG1_REG_10__SCAN_IN), .B2(
        n4565), .ZN(n3207) );
  OAI21_X1 U3971 ( .B1(n3208), .B2(n4565), .A(n3207), .ZN(U3528) );
  NOR2_X1 U3972 ( .A1(n3210), .A2(n3209), .ZN(n3211) );
  NAND2_X1 U3973 ( .A1(n3998), .A2(n3641), .ZN(n3215) );
  NAND2_X1 U3974 ( .A1(n3233), .A2(n3649), .ZN(n3214) );
  NAND2_X1 U3975 ( .A1(n3215), .A2(n3214), .ZN(n3216) );
  XNOR2_X1 U3976 ( .A(n3216), .B(n3652), .ZN(n3221) );
  INV_X1 U3977 ( .A(n3221), .ZN(n3219) );
  NOR2_X1 U3978 ( .A1(n3645), .A2(n3238), .ZN(n3217) );
  AOI21_X1 U3979 ( .B1(n3998), .B2(n2960), .A(n3217), .ZN(n3220) );
  INV_X1 U3980 ( .A(n3220), .ZN(n3218) );
  NAND2_X1 U3981 ( .A1(n3219), .A2(n3218), .ZN(n3250) );
  INV_X1 U3982 ( .A(n3250), .ZN(n3222) );
  AND2_X1 U3983 ( .A1(n3221), .A2(n3220), .ZN(n3249) );
  NOR2_X1 U3984 ( .A1(n3222), .A2(n3249), .ZN(n3223) );
  XNOR2_X1 U3985 ( .A(n3251), .B(n3223), .ZN(n3224) );
  NAND2_X1 U3986 ( .A1(n3224), .A2(n3806), .ZN(n3230) );
  OAI22_X1 U3987 ( .A1(n3779), .A2(n3238), .B1(n3290), .B2(n3813), .ZN(n3228)
         );
  OAI21_X1 U3988 ( .B1(n3808), .B2(n3226), .A(n3225), .ZN(n3227) );
  NOR2_X1 U3989 ( .A1(n3228), .A2(n3227), .ZN(n3229) );
  OAI211_X1 U3990 ( .C1(n3819), .C2(n4501), .A(n3230), .B(n3229), .ZN(U3218)
         );
  AND2_X1 U3991 ( .A1(n3935), .A2(n3931), .ZN(n3889) );
  XOR2_X1 U3992 ( .A(n3889), .B(n3231), .Z(n4504) );
  XOR2_X1 U3993 ( .A(n3889), .B(n3232), .Z(n3237) );
  AOI22_X1 U3994 ( .A1(n3999), .A2(n2048), .B1(n3233), .B2(n4324), .ZN(n3234)
         );
  OAI21_X1 U3995 ( .B1(n3290), .B2(n4304), .A(n3234), .ZN(n3236) );
  NOR2_X1 U3996 ( .A1(n4504), .A2(n4227), .ZN(n3235) );
  AOI211_X1 U3997 ( .C1(n4231), .C2(n3237), .A(n3236), .B(n3235), .ZN(n4510)
         );
  OAI21_X1 U3998 ( .B1(n4540), .B2(n4504), .A(n4510), .ZN(n3247) );
  NOR2_X1 U3999 ( .A1(n3239), .A2(n3238), .ZN(n3240) );
  OR2_X1 U4000 ( .A1(n3241), .A2(n3240), .ZN(n4505) );
  INV_X1 U4001 ( .A(REG1_REG_8__SCAN_IN), .ZN(n3242) );
  OAI22_X1 U4002 ( .A1(n4505), .A2(n4319), .B1(n4568), .B2(n3242), .ZN(n3243)
         );
  AOI21_X1 U4003 ( .B1(n3247), .B2(n4568), .A(n3243), .ZN(n3244) );
  INV_X1 U4004 ( .A(n3244), .ZN(U3526) );
  INV_X1 U4005 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3245) );
  OAI22_X1 U4006 ( .A1(n4505), .A2(n4378), .B1(n4559), .B2(n3245), .ZN(n3246)
         );
  AOI21_X1 U4007 ( .B1(n3247), .B2(n4559), .A(n3246), .ZN(n3248) );
  INV_X1 U4008 ( .A(n3248), .ZN(U3483) );
  NAND2_X1 U4009 ( .A1(n3997), .A2(n3189), .ZN(n3254) );
  NAND2_X1 U4010 ( .A1(n3252), .A2(n3649), .ZN(n3253) );
  NAND2_X1 U4011 ( .A1(n3254), .A2(n3253), .ZN(n3255) );
  XNOR2_X1 U4012 ( .A(n3255), .B(n3658), .ZN(n3279) );
  OAI22_X1 U4013 ( .A1(n3290), .A2(n2907), .B1(n3645), .B2(n3258), .ZN(n3278)
         );
  XNOR2_X1 U4014 ( .A(n3279), .B(n3278), .ZN(n3280) );
  XNOR2_X1 U4015 ( .A(n3281), .B(n3280), .ZN(n3256) );
  NAND2_X1 U4016 ( .A1(n3256), .A2(n3806), .ZN(n3263) );
  OAI22_X1 U4017 ( .A1(n3779), .A2(n3258), .B1(n3257), .B2(n3808), .ZN(n3261)
         );
  INV_X1 U4018 ( .A(REG3_REG_9__SCAN_IN), .ZN(n4677) );
  NOR2_X1 U4019 ( .A1(STATE_REG_SCAN_IN), .A2(n4677), .ZN(n4407) );
  INV_X1 U4020 ( .A(n4407), .ZN(n3259) );
  OAI21_X1 U4021 ( .B1(n3813), .B2(n3398), .A(n3259), .ZN(n3260) );
  NOR2_X1 U4022 ( .A1(n3261), .A2(n3260), .ZN(n3262) );
  OAI211_X1 U4023 ( .C1(n3819), .C2(n3264), .A(n3263), .B(n3262), .ZN(U3228)
         );
  INV_X1 U4024 ( .A(n3265), .ZN(n3266) );
  AOI21_X1 U4025 ( .B1(n3897), .B2(n3267), .A(n3266), .ZN(n3329) );
  AOI22_X1 U4026 ( .A1(n3994), .A2(n4325), .B1(n4324), .B2(n3395), .ZN(n3270)
         );
  XNOR2_X1 U4027 ( .A(n3302), .B(n3897), .ZN(n3268) );
  NAND2_X1 U4028 ( .A1(n3268), .A2(n4231), .ZN(n3269) );
  OAI211_X1 U4029 ( .C1(n3329), .C2(n4227), .A(n3270), .B(n3269), .ZN(n3331)
         );
  NAND2_X1 U4030 ( .A1(n3331), .A2(n4213), .ZN(n3277) );
  OAI22_X1 U4031 ( .A1(n4213), .A2(n3271), .B1(n3405), .B2(n4500), .ZN(n3275)
         );
  INV_X1 U4032 ( .A(n3316), .ZN(n3272) );
  OAI21_X1 U4033 ( .B1(n3273), .B2(n3399), .A(n3272), .ZN(n3337) );
  NOR2_X1 U4034 ( .A1(n3337), .A2(n4195), .ZN(n3274) );
  AOI211_X1 U4035 ( .C1(n3561), .C2(n3996), .A(n3275), .B(n3274), .ZN(n3276)
         );
  OAI211_X1 U4036 ( .C1(n3329), .C2(n4238), .A(n3277), .B(n3276), .ZN(U3279)
         );
  AOI22_X1 U4037 ( .A1(n3996), .A2(n2960), .B1(n3641), .B2(n3282), .ZN(n3391)
         );
  NAND2_X1 U4038 ( .A1(n3996), .A2(n3641), .ZN(n3284) );
  NAND2_X1 U4039 ( .A1(n3282), .A2(n3649), .ZN(n3283) );
  NAND2_X1 U4040 ( .A1(n3284), .A2(n3283), .ZN(n3285) );
  XNOR2_X1 U4041 ( .A(n3285), .B(n3658), .ZN(n3390) );
  XOR2_X1 U4042 ( .A(n3391), .B(n3390), .Z(n3286) );
  AOI21_X1 U40430 ( .B1(n3287), .B2(n3286), .A(n3800), .ZN(n3288) );
  NAND2_X1 U4044 ( .A1(n3288), .A2(n3393), .ZN(n3294) );
  OAI22_X1 U4045 ( .A1(n3779), .A2(n3289), .B1(n3455), .B2(n3813), .ZN(n3292)
         );
  NAND2_X1 U4046 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4411) );
  OAI21_X1 U4047 ( .B1(n3808), .B2(n3290), .A(n4411), .ZN(n3291) );
  NOR2_X1 U4048 ( .A1(n3292), .A2(n3291), .ZN(n3293) );
  OAI211_X1 U4049 ( .C1(n3819), .C2(n3295), .A(n3294), .B(n3293), .ZN(U3214)
         );
  INV_X1 U4050 ( .A(n3296), .ZN(n3298) );
  OR2_X1 U4051 ( .A1(n3298), .A2(n3297), .ZN(n3887) );
  XNOR2_X1 U4052 ( .A(n3339), .B(n3887), .ZN(n3372) );
  INV_X1 U4053 ( .A(n3372), .ZN(n3312) );
  INV_X1 U4054 ( .A(n3299), .ZN(n3300) );
  AOI21_X1 U4055 ( .B1(n3302), .B2(n3301), .A(n3300), .ZN(n3324) );
  INV_X1 U4056 ( .A(n3314), .ZN(n3303) );
  AOI21_X1 U4057 ( .B1(n3324), .B2(n3315), .A(n3303), .ZN(n3304) );
  XNOR2_X1 U4058 ( .A(n3304), .B(n3887), .ZN(n3307) );
  OAI22_X1 U4059 ( .A1(n3809), .A2(n4304), .B1(n3539), .B2(n3497), .ZN(n3305)
         );
  AOI21_X1 U4060 ( .B1(n2048), .B2(n3994), .A(n3305), .ZN(n3306) );
  OAI21_X1 U4061 ( .B1(n3307), .B2(n3408), .A(n3306), .ZN(n3371) );
  OAI21_X1 U4062 ( .B1(n3318), .B2(n3497), .A(n3346), .ZN(n3377) );
  INV_X1 U4063 ( .A(n3503), .ZN(n3308) );
  AOI22_X1 U4064 ( .A1(n4519), .A2(REG2_REG_13__SCAN_IN), .B1(n3308), .B2(
        n4511), .ZN(n3309) );
  OAI21_X1 U4065 ( .B1(n3377), .B2(n4195), .A(n3309), .ZN(n3310) );
  AOI21_X1 U4066 ( .B1(n3371), .B2(n4213), .A(n3310), .ZN(n3311) );
  OAI21_X1 U4067 ( .B1(n3312), .B2(n4198), .A(n3311), .ZN(U3277) );
  NAND2_X1 U4068 ( .A1(n3315), .A2(n3314), .ZN(n3873) );
  XNOR2_X1 U4069 ( .A(n3313), .B(n3873), .ZN(n3381) );
  NOR2_X1 U4070 ( .A1(n3316), .A2(n3454), .ZN(n3317) );
  OR2_X1 U4071 ( .A1(n3318), .A2(n3317), .ZN(n3389) );
  OAI22_X1 U4072 ( .A1(n4213), .A2(n3319), .B1(n3460), .B2(n4500), .ZN(n3320)
         );
  AOI21_X1 U4073 ( .B1(n3561), .B2(n3995), .A(n3320), .ZN(n3323) );
  INV_X1 U4074 ( .A(n3993), .ZN(n3526) );
  OAI22_X1 U4075 ( .A1(n3526), .A2(n4170), .B1(n4169), .B2(n3454), .ZN(n3321)
         );
  INV_X1 U4076 ( .A(n3321), .ZN(n3322) );
  OAI211_X1 U4077 ( .C1(n3389), .C2(n4195), .A(n3323), .B(n3322), .ZN(n3327)
         );
  XNOR2_X1 U4078 ( .A(n3324), .B(n3873), .ZN(n3325) );
  NAND2_X1 U4079 ( .A1(n3325), .A2(n4231), .ZN(n3379) );
  NOR2_X1 U4080 ( .A1(n3379), .A2(n4519), .ZN(n3326) );
  AOI211_X1 U4081 ( .C1(n4209), .C2(n3381), .A(n3327), .B(n3326), .ZN(n3328)
         );
  INV_X1 U4082 ( .A(n3328), .ZN(U3278) );
  INV_X1 U4083 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3332) );
  OAI22_X1 U4084 ( .A1(n3329), .A2(n4540), .B1(n3398), .B2(n4328), .ZN(n3330)
         );
  NOR2_X1 U4085 ( .A1(n3331), .A2(n3330), .ZN(n3334) );
  MUX2_X1 U4086 ( .A(n3332), .B(n3334), .S(n4568), .Z(n3333) );
  OAI21_X1 U4087 ( .B1(n4319), .B2(n3337), .A(n3333), .ZN(U3529) );
  INV_X1 U4088 ( .A(REG0_REG_11__SCAN_IN), .ZN(n3335) );
  MUX2_X1 U4089 ( .A(n3335), .B(n3334), .S(n4559), .Z(n3336) );
  OAI21_X1 U4090 ( .B1(n3337), .B2(n4378), .A(n3336), .ZN(U3489) );
  XNOR2_X1 U4091 ( .A(n3821), .B(n3344), .ZN(n3409) );
  OR2_X1 U4092 ( .A1(n3339), .A2(n3338), .ZN(n3342) );
  AND2_X1 U4093 ( .A1(n3342), .A2(n3340), .ZN(n3345) );
  NAND2_X1 U4094 ( .A1(n3342), .A2(n3341), .ZN(n3343) );
  OAI21_X1 U4095 ( .B1(n3345), .B2(n3344), .A(n3343), .ZN(n3411) );
  NAND2_X1 U4096 ( .A1(n3411), .A2(n4209), .ZN(n3354) );
  INV_X1 U4097 ( .A(n3346), .ZN(n3347) );
  OAI21_X1 U4098 ( .B1(n3347), .B2(n3524), .A(n3362), .ZN(n3417) );
  INV_X1 U4099 ( .A(n3417), .ZN(n3352) );
  AOI22_X1 U4100 ( .A1(n3430), .A2(n3519), .B1(n3429), .B2(n3991), .ZN(n3350)
         );
  INV_X1 U4101 ( .A(n3531), .ZN(n3348) );
  AOI22_X1 U4102 ( .A1(n4519), .A2(REG2_REG_14__SCAN_IN), .B1(n3348), .B2(
        n4511), .ZN(n3349) );
  OAI211_X1 U4103 ( .C1(n3526), .C2(n4167), .A(n3350), .B(n3349), .ZN(n3351)
         );
  AOI21_X1 U4104 ( .B1(n3352), .B2(n4513), .A(n3351), .ZN(n3353) );
  OAI211_X1 U4105 ( .C1(n3409), .C2(n3355), .A(n3354), .B(n3353), .ZN(U3276)
         );
  AOI21_X1 U4106 ( .B1(n3356), .B2(n3892), .A(n3408), .ZN(n3358) );
  NAND2_X1 U4107 ( .A1(n3358), .A2(n3357), .ZN(n3419) );
  AND2_X1 U4108 ( .A1(n3360), .A2(n3359), .ZN(n3361) );
  XNOR2_X1 U4109 ( .A(n3361), .B(n3892), .ZN(n3421) );
  NAND2_X1 U4110 ( .A1(n3421), .A2(n4209), .ZN(n3370) );
  INV_X1 U4111 ( .A(n3362), .ZN(n3363) );
  OAI21_X1 U4112 ( .B1(n3363), .B2(n3810), .A(n3428), .ZN(n3427) );
  INV_X1 U4113 ( .A(n3427), .ZN(n3368) );
  AOI22_X1 U4114 ( .A1(n3430), .A2(n3574), .B1(n3429), .B2(n3990), .ZN(n3366)
         );
  INV_X1 U4115 ( .A(n3818), .ZN(n3364) );
  AOI22_X1 U4116 ( .A1(n4519), .A2(REG2_REG_15__SCAN_IN), .B1(n3364), .B2(
        n4511), .ZN(n3365) );
  OAI211_X1 U4117 ( .C1(n3809), .C2(n4167), .A(n3366), .B(n3365), .ZN(n3367)
         );
  AOI21_X1 U4118 ( .B1(n3368), .B2(n4513), .A(n3367), .ZN(n3369) );
  OAI211_X1 U4119 ( .C1(n4519), .C2(n3419), .A(n3370), .B(n3369), .ZN(U3275)
         );
  AOI21_X1 U4120 ( .B1(n4316), .B2(n3372), .A(n3371), .ZN(n3374) );
  MUX2_X1 U4121 ( .A(n4045), .B(n3374), .S(n4568), .Z(n3373) );
  OAI21_X1 U4122 ( .B1(n4319), .B2(n3377), .A(n3373), .ZN(U3531) );
  INV_X1 U4123 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3375) );
  MUX2_X1 U4124 ( .A(n3375), .B(n3374), .S(n4559), .Z(n3376) );
  OAI21_X1 U4125 ( .B1(n3377), .B2(n4378), .A(n3376), .ZN(U3493) );
  INV_X1 U4126 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3384) );
  AOI22_X1 U4127 ( .A1(n2048), .A2(n3995), .B1(n3993), .B2(n4325), .ZN(n3378)
         );
  OAI211_X1 U4128 ( .C1(n3539), .C2(n3454), .A(n3379), .B(n3378), .ZN(n3380)
         );
  INV_X1 U4129 ( .A(n3380), .ZN(n3383) );
  NAND2_X1 U4130 ( .A1(n3381), .A2(n4316), .ZN(n3382) );
  AND2_X1 U4131 ( .A1(n3383), .A2(n3382), .ZN(n3386) );
  MUX2_X1 U4132 ( .A(n3384), .B(n3386), .S(n4559), .Z(n3385) );
  OAI21_X1 U4133 ( .B1(n3389), .B2(n4378), .A(n3385), .ZN(U3491) );
  INV_X1 U4134 ( .A(REG1_REG_12__SCAN_IN), .ZN(n3387) );
  MUX2_X1 U4135 ( .A(n3387), .B(n3386), .S(n4568), .Z(n3388) );
  OAI21_X1 U4136 ( .B1(n4319), .B2(n3389), .A(n3388), .ZN(U3530) );
  OAI22_X1 U4137 ( .A1(n3455), .A2(n3645), .B1(n3657), .B2(n3399), .ZN(n3394)
         );
  XNOR2_X1 U4138 ( .A(n3394), .B(n3658), .ZN(n3444) );
  AOI22_X1 U4139 ( .A1(n3995), .A2(n2960), .B1(n3641), .B2(n3395), .ZN(n3440)
         );
  INV_X1 U4140 ( .A(n3440), .ZN(n3443) );
  XNOR2_X1 U4141 ( .A(n3444), .B(n3443), .ZN(n3396) );
  XNOR2_X1 U4142 ( .A(n3442), .B(n3396), .ZN(n3397) );
  NAND2_X1 U4143 ( .A1(n3397), .A2(n3806), .ZN(n3404) );
  OAI22_X1 U4144 ( .A1(n3779), .A2(n3399), .B1(n3398), .B2(n3808), .ZN(n3402)
         );
  AND2_X1 U4145 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4427) );
  INV_X1 U4146 ( .A(n4427), .ZN(n3400) );
  OAI21_X1 U4147 ( .B1(n3813), .B2(n3496), .A(n3400), .ZN(n3401) );
  NOR2_X1 U4148 ( .A1(n3402), .A2(n3401), .ZN(n3403) );
  OAI211_X1 U4149 ( .C1(n3819), .C2(n3405), .A(n3404), .B(n3403), .ZN(U3233)
         );
  OAI22_X1 U4150 ( .A1(n4329), .A2(n4304), .B1(n3539), .B2(n3524), .ZN(n3406)
         );
  AOI21_X1 U4151 ( .B1(n2048), .B2(n3993), .A(n3406), .ZN(n3407) );
  OAI21_X1 U4152 ( .B1(n3409), .B2(n3408), .A(n3407), .ZN(n3410) );
  AOI21_X1 U4153 ( .B1(n3411), .B2(n4316), .A(n3410), .ZN(n3415) );
  INV_X1 U4154 ( .A(REG1_REG_14__SCAN_IN), .ZN(n3412) );
  MUX2_X1 U4155 ( .A(n3415), .B(n3412), .S(n4565), .Z(n3413) );
  OAI21_X1 U4156 ( .B1(n4319), .B2(n3417), .A(n3413), .ZN(U3532) );
  INV_X1 U4157 ( .A(REG0_REG_14__SCAN_IN), .ZN(n3414) );
  MUX2_X1 U4158 ( .A(n3415), .B(n3414), .S(n4557), .Z(n3416) );
  OAI21_X1 U4159 ( .B1(n3417), .B2(n4378), .A(n3416), .ZN(U3495) );
  AOI22_X1 U4160 ( .A1(n3990), .A2(n4325), .B1(n4324), .B2(n3574), .ZN(n3418)
         );
  OAI211_X1 U4161 ( .C1(n3809), .C2(n4328), .A(n3419), .B(n3418), .ZN(n3420)
         );
  AOI21_X1 U4162 ( .B1(n3421), .B2(n4316), .A(n3420), .ZN(n3425) );
  INV_X1 U4163 ( .A(REG0_REG_15__SCAN_IN), .ZN(n3422) );
  MUX2_X1 U4164 ( .A(n3425), .B(n3422), .S(n4557), .Z(n3423) );
  OAI21_X1 U4165 ( .B1(n3427), .B2(n4378), .A(n3423), .ZN(U3497) );
  INV_X1 U4166 ( .A(REG1_REG_15__SCAN_IN), .ZN(n3424) );
  MUX2_X1 U4167 ( .A(n3425), .B(n3424), .S(n4565), .Z(n3426) );
  OAI21_X1 U4168 ( .B1(n4319), .B2(n3427), .A(n3426), .ZN(U3533) );
  INV_X1 U4169 ( .A(n3435), .ZN(n3869) );
  OAI21_X1 U4170 ( .B1(n2094), .B2(n3869), .A(n2324), .ZN(n4334) );
  AOI21_X1 U4171 ( .B1(n4323), .B2(n3428), .A(n3464), .ZN(n4331) );
  AOI22_X1 U4172 ( .A1(n3430), .A2(n4323), .B1(n3429), .B2(n4326), .ZN(n3433)
         );
  INV_X1 U4173 ( .A(n3726), .ZN(n3431) );
  AOI22_X1 U4174 ( .A1(n4519), .A2(REG2_REG_16__SCAN_IN), .B1(n3431), .B2(
        n4511), .ZN(n3432) );
  OAI211_X1 U4175 ( .C1(n4329), .C2(n4167), .A(n3433), .B(n3432), .ZN(n3438)
         );
  OAI211_X1 U4176 ( .C1(n3436), .C2(n3435), .A(n3434), .B(n4231), .ZN(n4332)
         );
  NOR2_X1 U4177 ( .A1(n4332), .A2(n4519), .ZN(n3437) );
  AOI211_X1 U4178 ( .C1(n4331), .C2(n4513), .A(n3438), .B(n3437), .ZN(n3439)
         );
  OAI21_X1 U4179 ( .B1(n4334), .B2(n4198), .A(n3439), .ZN(U3274) );
  NAND2_X1 U4180 ( .A1(n3441), .A2(n3440), .ZN(n3445) );
  NAND2_X1 U4181 ( .A1(n3994), .A2(n3641), .ZN(n3447) );
  NAND2_X1 U4182 ( .A1(n3449), .A2(n3649), .ZN(n3446) );
  NAND2_X1 U4183 ( .A1(n3447), .A2(n3446), .ZN(n3448) );
  XNOR2_X1 U4184 ( .A(n3448), .B(n3652), .ZN(n3451) );
  AOI22_X1 U4185 ( .A1(n3994), .A2(n2960), .B1(n3641), .B2(n3449), .ZN(n3450)
         );
  OR2_X1 U4186 ( .A1(n3451), .A2(n3450), .ZN(n3490) );
  AND2_X1 U4187 ( .A1(n3451), .A2(n3450), .ZN(n3489) );
  NOR2_X1 U4188 ( .A1(n2203), .A2(n3489), .ZN(n3452) );
  XNOR2_X1 U4189 ( .A(n3491), .B(n3452), .ZN(n3453) );
  NAND2_X1 U4190 ( .A1(n3453), .A2(n3806), .ZN(n3459) );
  OAI22_X1 U4191 ( .A1(n3779), .A2(n3454), .B1(n3526), .B2(n3813), .ZN(n3457)
         );
  NAND2_X1 U4192 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4431) );
  OAI21_X1 U4193 ( .B1(n3808), .B2(n3455), .A(n4431), .ZN(n3456) );
  NOR2_X1 U4194 ( .A1(n3457), .A2(n3456), .ZN(n3458) );
  OAI211_X1 U4195 ( .C1(n3819), .C2(n3460), .A(n3459), .B(n3458), .ZN(U3221)
         );
  INV_X1 U4196 ( .A(n3475), .ZN(n3461) );
  NAND2_X1 U4197 ( .A1(n3461), .A2(n3474), .ZN(n3868) );
  XNOR2_X1 U4198 ( .A(n3476), .B(n3868), .ZN(n3462) );
  NAND2_X1 U4199 ( .A1(n3462), .A2(n4231), .ZN(n3505) );
  XOR2_X1 U4200 ( .A(n3868), .B(n3463), .Z(n3507) );
  NAND2_X1 U4201 ( .A1(n3507), .A2(n4209), .ZN(n3470) );
  OAI21_X1 U4202 ( .B1(n3464), .B2(n3733), .A(n3482), .ZN(n3512) );
  INV_X1 U4203 ( .A(n3512), .ZN(n3468) );
  AOI22_X1 U4204 ( .A1(n4519), .A2(REG2_REG_17__SCAN_IN), .B1(n3738), .B2(
        n4511), .ZN(n3465) );
  OAI21_X1 U4205 ( .B1(n4167), .B2(n3812), .A(n3465), .ZN(n3467) );
  OAI22_X1 U4206 ( .A1(n3735), .A2(n4170), .B1(n4169), .B2(n3733), .ZN(n3466)
         );
  AOI211_X1 U4207 ( .C1(n3468), .C2(n4513), .A(n3467), .B(n3466), .ZN(n3469)
         );
  OAI211_X1 U4208 ( .C1(n4519), .C2(n3505), .A(n3470), .B(n3469), .ZN(U3273)
         );
  OAI21_X1 U4209 ( .B1(n3471), .B2(n3477), .A(n3472), .ZN(n3473) );
  INV_X1 U4210 ( .A(n3473), .ZN(n4322) );
  OAI21_X1 U4211 ( .B1(n3476), .B2(n3475), .A(n3474), .ZN(n3536) );
  XNOR2_X1 U4212 ( .A(n3536), .B(n2175), .ZN(n3480) );
  INV_X1 U4213 ( .A(n4326), .ZN(n3777) );
  AOI22_X1 U4214 ( .A1(n4223), .A2(n4325), .B1(n4324), .B2(n3597), .ZN(n3478)
         );
  OAI21_X1 U4215 ( .B1(n3777), .B2(n4328), .A(n3478), .ZN(n3479) );
  AOI21_X1 U4216 ( .B1(n3480), .B2(n4231), .A(n3479), .ZN(n4321) );
  INV_X1 U4217 ( .A(n4321), .ZN(n3487) );
  AOI21_X1 U4218 ( .B1(n3482), .B2(n3597), .A(n3481), .ZN(n3483) );
  NAND2_X1 U4219 ( .A1(n3483), .A2(n3543), .ZN(n4320) );
  AOI22_X1 U4220 ( .A1(n4519), .A2(REG2_REG_18__SCAN_IN), .B1(n3783), .B2(
        n4511), .ZN(n3484) );
  OAI21_X1 U4221 ( .B1(n4320), .B2(n3485), .A(n3484), .ZN(n3486) );
  AOI21_X1 U4222 ( .B1(n3487), .B2(n4213), .A(n3486), .ZN(n3488) );
  OAI21_X1 U4223 ( .B1(n4322), .B2(n4198), .A(n3488), .ZN(U3272) );
  AOI22_X1 U4224 ( .A1(n3993), .A2(n3641), .B1(n3649), .B2(n3492), .ZN(n3493)
         );
  XOR2_X1 U4225 ( .A(n3658), .B(n3493), .Z(n3514) );
  OAI22_X1 U4226 ( .A1(n3526), .A2(n2907), .B1(n3645), .B2(n3497), .ZN(n3513)
         );
  XNOR2_X1 U4227 ( .A(n3514), .B(n3513), .ZN(n3494) );
  XNOR2_X1 U4228 ( .A(n3515), .B(n3494), .ZN(n3495) );
  NAND2_X1 U4229 ( .A1(n3495), .A2(n3806), .ZN(n3502) );
  OAI22_X1 U4230 ( .A1(n3779), .A2(n3497), .B1(n3496), .B2(n3808), .ZN(n3500)
         );
  INV_X1 U4231 ( .A(REG3_REG_13__SCAN_IN), .ZN(n4574) );
  NOR2_X1 U4232 ( .A1(STATE_REG_SCAN_IN), .A2(n4574), .ZN(n4444) );
  INV_X1 U4233 ( .A(n4444), .ZN(n3498) );
  OAI21_X1 U4234 ( .B1(n3813), .B2(n3809), .A(n3498), .ZN(n3499) );
  NOR2_X1 U4235 ( .A1(n3500), .A2(n3499), .ZN(n3501) );
  OAI211_X1 U4236 ( .C1(n3819), .C2(n3503), .A(n3502), .B(n3501), .ZN(U3231)
         );
  AOI22_X1 U4237 ( .A1(n3990), .A2(n2048), .B1(n3590), .B2(n4324), .ZN(n3504)
         );
  OAI211_X1 U4238 ( .C1(n3735), .C2(n4304), .A(n3505), .B(n3504), .ZN(n3506)
         );
  AOI21_X1 U4239 ( .B1(n3507), .B2(n4316), .A(n3506), .ZN(n3510) );
  MUX2_X1 U4240 ( .A(n3510), .B(n4069), .S(n4565), .Z(n3508) );
  OAI21_X1 U4241 ( .B1(n4319), .B2(n3512), .A(n3508), .ZN(U3535) );
  INV_X1 U4242 ( .A(REG0_REG_17__SCAN_IN), .ZN(n3509) );
  MUX2_X1 U4243 ( .A(n3510), .B(n3509), .S(n4557), .Z(n3511) );
  OAI21_X1 U4244 ( .B1(n3512), .B2(n4378), .A(n3511), .ZN(U3501) );
  NAND2_X1 U4245 ( .A1(n3992), .A2(n3189), .ZN(n3517) );
  NAND2_X1 U4246 ( .A1(n3519), .A2(n3649), .ZN(n3516) );
  NAND2_X1 U4247 ( .A1(n3517), .A2(n3516), .ZN(n3518) );
  XNOR2_X1 U4248 ( .A(n3518), .B(n3652), .ZN(n3521) );
  AOI22_X1 U4249 ( .A1(n3992), .A2(n2960), .B1(n3641), .B2(n3519), .ZN(n3520)
         );
  NAND2_X1 U4250 ( .A1(n3521), .A2(n3520), .ZN(n3571) );
  NAND2_X1 U4251 ( .A1(n2325), .A2(n3571), .ZN(n3522) );
  XNOR2_X1 U4252 ( .A(n3570), .B(n3522), .ZN(n3523) );
  NAND2_X1 U4253 ( .A1(n3523), .A2(n3806), .ZN(n3530) );
  OAI22_X1 U4254 ( .A1(n3779), .A2(n3524), .B1(n4329), .B2(n3813), .ZN(n3528)
         );
  INV_X1 U4255 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4694) );
  NOR2_X1 U4256 ( .A1(n4694), .A2(STATE_REG_SCAN_IN), .ZN(n4454) );
  INV_X1 U4257 ( .A(n4454), .ZN(n3525) );
  OAI21_X1 U4258 ( .B1(n3808), .B2(n3526), .A(n3525), .ZN(n3527) );
  NOR2_X1 U4259 ( .A1(n3528), .A2(n3527), .ZN(n3529) );
  OAI211_X1 U4260 ( .C1(n3819), .C2(n3531), .A(n3530), .B(n3529), .ZN(U3212)
         );
  XNOR2_X1 U4261 ( .A(n4223), .B(n3599), .ZN(n3875) );
  XOR2_X1 U4262 ( .A(n3875), .B(n3532), .Z(n4317) );
  INV_X1 U4263 ( .A(n4317), .ZN(n3549) );
  INV_X1 U4264 ( .A(n3533), .ZN(n3535) );
  OAI21_X1 U4265 ( .B1(n3536), .B2(n3535), .A(n3534), .ZN(n3537) );
  XOR2_X1 U4266 ( .A(n3875), .B(n3537), .Z(n3538) );
  NAND2_X1 U4267 ( .A1(n3538), .A2(n4231), .ZN(n3542) );
  NOR2_X1 U4268 ( .A1(n3688), .A2(n3539), .ZN(n3540) );
  AOI21_X1 U4269 ( .B1(n4301), .B2(n4325), .A(n3540), .ZN(n3541) );
  OAI211_X1 U4270 ( .C1(n3735), .C2(n4328), .A(n3542), .B(n3541), .ZN(n4315)
         );
  INV_X1 U4271 ( .A(n3543), .ZN(n3544) );
  OAI21_X1 U4272 ( .B1(n3544), .B2(n3688), .A(n2074), .ZN(n4379) );
  NOR2_X1 U4273 ( .A1(n4379), .A2(n4195), .ZN(n3547) );
  OAI22_X1 U4274 ( .A1(n4213), .A2(n3545), .B1(n3692), .B2(n4500), .ZN(n3546)
         );
  AOI211_X1 U4275 ( .C1(n4315), .C2(n4213), .A(n3547), .B(n3546), .ZN(n3548)
         );
  OAI21_X1 U4276 ( .B1(n3549), .B2(n4198), .A(n3548), .ZN(U3271) );
  INV_X1 U4277 ( .A(n4177), .ZN(n3954) );
  NAND2_X1 U4278 ( .A1(n3954), .A2(n4179), .ZN(n3872) );
  XNOR2_X1 U4279 ( .A(n4178), .B(n3872), .ZN(n3550) );
  NAND2_X1 U4280 ( .A1(n3550), .A2(n4231), .ZN(n4303) );
  XNOR2_X1 U4281 ( .A(n3551), .B(n3872), .ZN(n4307) );
  NAND2_X1 U4282 ( .A1(n4307), .A2(n4209), .ZN(n3558) );
  OAI21_X1 U4283 ( .B1(n4234), .B2(n3703), .A(n4210), .ZN(n4373) );
  INV_X1 U4284 ( .A(n4373), .ZN(n3556) );
  INV_X1 U4285 ( .A(n4301), .ZN(n3689) );
  INV_X1 U4286 ( .A(n3709), .ZN(n3552) );
  AOI22_X1 U4287 ( .A1(n4519), .A2(REG2_REG_21__SCAN_IN), .B1(n3552), .B2(
        n4511), .ZN(n3553) );
  OAI21_X1 U4288 ( .B1(n4167), .B2(n3689), .A(n3553), .ZN(n3555) );
  INV_X1 U4289 ( .A(n4186), .ZN(n4305) );
  OAI22_X1 U4290 ( .A1(n4305), .A2(n4170), .B1(n4169), .B2(n3703), .ZN(n3554)
         );
  AOI211_X1 U4291 ( .C1(n3556), .C2(n4513), .A(n3555), .B(n3554), .ZN(n3557)
         );
  OAI211_X1 U4292 ( .C1(n4519), .C2(n4303), .A(n3558), .B(n3557), .ZN(U3269)
         );
  OAI22_X1 U4293 ( .A1(n4169), .A2(n3844), .B1(n3559), .B2(n4213), .ZN(n3560)
         );
  AOI21_X1 U4294 ( .B1(n3987), .B2(n3561), .A(n3560), .ZN(n3568) );
  INV_X1 U4295 ( .A(n3562), .ZN(n3566) );
  OAI22_X1 U4296 ( .A1(n3564), .A2(n4195), .B1(n3563), .B2(n4500), .ZN(n3565)
         );
  OAI21_X1 U4297 ( .B1(n3566), .B2(n3565), .A(n4213), .ZN(n3567) );
  OAI211_X1 U4298 ( .C1(n3569), .C2(n4198), .A(n3568), .B(n3567), .ZN(U3354)
         );
  NAND2_X1 U4299 ( .A1(n3572), .A2(n3571), .ZN(n3578) );
  OAI22_X1 U4300 ( .A1(n4329), .A2(n3645), .B1(n3657), .B2(n3810), .ZN(n3573)
         );
  XOR2_X1 U4301 ( .A(n3658), .B(n3573), .Z(n3577) );
  NAND2_X1 U4302 ( .A1(n3578), .A2(n3577), .ZN(n3802) );
  NAND2_X1 U4303 ( .A1(n3991), .A2(n2960), .ZN(n3576) );
  NAND2_X1 U4304 ( .A1(n3574), .A2(n3641), .ZN(n3575) );
  NAND2_X1 U4305 ( .A1(n3576), .A2(n3575), .ZN(n3804) );
  NAND2_X1 U4306 ( .A1(n3802), .A2(n3804), .ZN(n3586) );
  NOR2_X1 U4307 ( .A1(n3578), .A2(n3577), .ZN(n3579) );
  NAND2_X1 U4308 ( .A1(n3990), .A2(n3641), .ZN(n3581) );
  NAND2_X1 U4309 ( .A1(n4323), .A2(n3649), .ZN(n3580) );
  NAND2_X1 U4310 ( .A1(n3581), .A2(n3580), .ZN(n3582) );
  XNOR2_X1 U4311 ( .A(n3582), .B(n3652), .ZN(n3584) );
  AOI22_X1 U4312 ( .A1(n3990), .A2(n2960), .B1(n3641), .B2(n4323), .ZN(n3583)
         );
  NAND2_X1 U4313 ( .A1(n3584), .A2(n3583), .ZN(n3727) );
  OAI21_X1 U4314 ( .B1(n3584), .B2(n3583), .A(n3727), .ZN(n3585) );
  INV_X1 U4315 ( .A(n3585), .ZN(n3718) );
  NAND2_X1 U4316 ( .A1(n4326), .A2(n3641), .ZN(n3588) );
  NAND2_X1 U4317 ( .A1(n3590), .A2(n3649), .ZN(n3587) );
  NAND2_X1 U4318 ( .A1(n3588), .A2(n3587), .ZN(n3589) );
  XNOR2_X1 U4319 ( .A(n3589), .B(n3658), .ZN(n3596) );
  INV_X1 U4320 ( .A(n3596), .ZN(n3594) );
  NAND2_X1 U4321 ( .A1(n4326), .A2(n2960), .ZN(n3592) );
  NAND2_X1 U4322 ( .A1(n3590), .A2(n3641), .ZN(n3591) );
  NAND2_X1 U4323 ( .A1(n3592), .A2(n3591), .ZN(n3595) );
  INV_X1 U4324 ( .A(n3595), .ZN(n3593) );
  NAND2_X1 U4325 ( .A1(n3594), .A2(n3593), .ZN(n3729) );
  NAND2_X1 U4326 ( .A1(n3596), .A2(n3595), .ZN(n3730) );
  AOI22_X1 U4327 ( .A1(n3989), .A2(n2960), .B1(n3641), .B2(n3597), .ZN(n3774)
         );
  OAI22_X1 U4328 ( .A1(n3735), .A2(n3645), .B1(n3657), .B2(n3778), .ZN(n3598)
         );
  XOR2_X1 U4329 ( .A(n3658), .B(n3598), .Z(n3775) );
  NAND2_X1 U4330 ( .A1(n4223), .A2(n3641), .ZN(n3601) );
  NAND2_X1 U4331 ( .A1(n3599), .A2(n3649), .ZN(n3600) );
  NAND2_X1 U4332 ( .A1(n3601), .A2(n3600), .ZN(n3602) );
  XNOR2_X1 U4333 ( .A(n3602), .B(n3652), .ZN(n3605) );
  NOR2_X1 U4334 ( .A1(n3688), .A2(n3645), .ZN(n3603) );
  AOI21_X1 U4335 ( .B1(n4223), .B2(n2960), .A(n3603), .ZN(n3604) );
  NAND2_X1 U4336 ( .A1(n3605), .A2(n3604), .ZN(n3606) );
  OAI21_X1 U4337 ( .B1(n3605), .B2(n3604), .A(n3606), .ZN(n3687) );
  NAND2_X1 U4338 ( .A1(n4301), .A2(n3641), .ZN(n3608) );
  NAND2_X1 U4339 ( .A1(n3649), .A2(n4235), .ZN(n3607) );
  NAND2_X1 U4340 ( .A1(n3608), .A2(n3607), .ZN(n3609) );
  XNOR2_X1 U4341 ( .A(n3609), .B(n3652), .ZN(n3612) );
  NOR2_X1 U4342 ( .A1(n3645), .A2(n3757), .ZN(n3610) );
  AOI21_X1 U4343 ( .B1(n4301), .B2(n2960), .A(n3610), .ZN(n3611) );
  OR2_X1 U4344 ( .A1(n3612), .A2(n3611), .ZN(n3754) );
  NAND2_X1 U4345 ( .A1(n3699), .A2(n3754), .ZN(n3751) );
  NAND2_X1 U4346 ( .A1(n3612), .A2(n3611), .ZN(n3753) );
  NAND2_X1 U4347 ( .A1(n3751), .A2(n3753), .ZN(n3702) );
  NAND2_X1 U4348 ( .A1(n4202), .A2(n3641), .ZN(n3614) );
  NAND2_X1 U4349 ( .A1(n3649), .A2(n4299), .ZN(n3613) );
  NAND2_X1 U4350 ( .A1(n3614), .A2(n3613), .ZN(n3615) );
  XNOR2_X1 U4351 ( .A(n3615), .B(n3652), .ZN(n3618) );
  NOR2_X1 U4352 ( .A1(n3645), .A2(n3703), .ZN(n3616) );
  AOI21_X1 U4353 ( .B1(n4202), .B2(n2960), .A(n3616), .ZN(n3617) );
  AND2_X1 U4354 ( .A1(n3618), .A2(n3617), .ZN(n3697) );
  OR2_X1 U4355 ( .A1(n3618), .A2(n3617), .ZN(n3698) );
  AOI22_X1 U4356 ( .A1(n4186), .A2(n3641), .B1(n3649), .B2(n4201), .ZN(n3619)
         );
  XNOR2_X1 U4357 ( .A(n3619), .B(n3658), .ZN(n3622) );
  AOI22_X1 U4358 ( .A1(n4186), .A2(n2960), .B1(n3641), .B2(n4201), .ZN(n3621)
         );
  XNOR2_X1 U4359 ( .A(n3622), .B(n3621), .ZN(n3766) );
  OAI22_X1 U4360 ( .A1(n4204), .A2(n3645), .B1(n3657), .B2(n3679), .ZN(n3620)
         );
  XNOR2_X1 U4361 ( .A(n3620), .B(n3652), .ZN(n3624) );
  OAI22_X1 U4362 ( .A1(n4204), .A2(n2907), .B1(n3645), .B2(n3679), .ZN(n3625)
         );
  XNOR2_X1 U4363 ( .A(n3624), .B(n3625), .ZN(n3677) );
  NAND2_X1 U4364 ( .A1(n3622), .A2(n3621), .ZN(n3678) );
  INV_X1 U4365 ( .A(n3624), .ZN(n3626) );
  NAND2_X1 U4366 ( .A1(n3626), .A2(n3625), .ZN(n3630) );
  NOR2_X1 U4367 ( .A1(n3645), .A2(n4168), .ZN(n3627) );
  AOI21_X1 U4368 ( .B1(n4147), .B2(n2960), .A(n3627), .ZN(n3631) );
  OAI22_X1 U4369 ( .A1(n4189), .A2(n3645), .B1(n3657), .B2(n4168), .ZN(n3629)
         );
  XNOR2_X1 U4370 ( .A(n3629), .B(n3658), .ZN(n3745) );
  NAND2_X1 U4371 ( .A1(n3742), .A2(n3745), .ZN(n3634) );
  INV_X1 U4372 ( .A(n3631), .ZN(n3632) );
  NAND2_X1 U4373 ( .A1(n3633), .A2(n3632), .ZN(n3743) );
  NAND2_X1 U4374 ( .A1(n3988), .A2(n3641), .ZN(n3636) );
  NAND2_X1 U4375 ( .A1(n3649), .A2(n4146), .ZN(n3635) );
  NAND2_X1 U4376 ( .A1(n3636), .A2(n3635), .ZN(n3637) );
  XNOR2_X1 U4377 ( .A(n3637), .B(n3652), .ZN(n3640) );
  NOR2_X1 U4378 ( .A1(n3645), .A2(n4152), .ZN(n3638) );
  AOI21_X1 U4379 ( .B1(n3988), .B2(n2960), .A(n3638), .ZN(n3639) );
  NAND2_X1 U4380 ( .A1(n3640), .A2(n3639), .ZN(n3710) );
  OR2_X1 U4381 ( .A1(n3640), .A2(n3639), .ZN(n3711) );
  NAND2_X1 U4382 ( .A1(n4261), .A2(n3641), .ZN(n3643) );
  NAND2_X1 U4383 ( .A1(n3649), .A2(n4269), .ZN(n3642) );
  NAND2_X1 U4384 ( .A1(n3643), .A2(n3642), .ZN(n3644) );
  XNOR2_X1 U4385 ( .A(n3644), .B(n3652), .ZN(n3648) );
  NOR2_X1 U4386 ( .A1(n3645), .A2(n4134), .ZN(n3646) );
  AOI21_X1 U4387 ( .B1(n4261), .B2(n2960), .A(n3646), .ZN(n3647) );
  NOR2_X1 U4388 ( .A1(n3648), .A2(n3647), .ZN(n3789) );
  NAND2_X1 U4389 ( .A1(n3648), .A2(n3647), .ZN(n3787) );
  NAND2_X1 U4390 ( .A1(n4270), .A2(n3641), .ZN(n3651) );
  NAND2_X1 U4391 ( .A1(n3649), .A2(n4260), .ZN(n3650) );
  NAND2_X1 U4392 ( .A1(n3651), .A2(n3650), .ZN(n3653) );
  XNOR2_X1 U4393 ( .A(n3653), .B(n3652), .ZN(n3656) );
  NOR2_X1 U4394 ( .A1(n3645), .A2(n4117), .ZN(n3654) );
  AOI21_X1 U4395 ( .B1(n4270), .B2(n2960), .A(n3654), .ZN(n3655) );
  XNOR2_X1 U4396 ( .A(n3656), .B(n3655), .ZN(n3669) );
  OAI22_X1 U4397 ( .A1(n4264), .A2(n2907), .B1(n3645), .B2(n4098), .ZN(n3661)
         );
  OAI22_X1 U4398 ( .A1(n4264), .A2(n3645), .B1(n3657), .B2(n4098), .ZN(n3659)
         );
  XNOR2_X1 U4399 ( .A(n3659), .B(n3658), .ZN(n3660) );
  XOR2_X1 U4400 ( .A(n3661), .B(n3660), .Z(n3662) );
  XNOR2_X1 U4401 ( .A(n3663), .B(n3662), .ZN(n3668) );
  INV_X1 U4402 ( .A(n4252), .ZN(n4099) );
  INV_X1 U4403 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3664) );
  OAI22_X1 U4404 ( .A1(n4099), .A2(n3813), .B1(STATE_REG_SCAN_IN), .B2(n3664), 
        .ZN(n3666) );
  OAI22_X1 U4405 ( .A1(n4255), .A2(n3808), .B1(n3779), .B2(n4098), .ZN(n3665)
         );
  AOI211_X1 U4406 ( .C1(n4096), .C2(n3793), .A(n3666), .B(n3665), .ZN(n3667)
         );
  OAI21_X1 U4407 ( .B1(n3668), .B2(n3800), .A(n3667), .ZN(U3217) );
  XNOR2_X1 U4408 ( .A(n3670), .B(n3669), .ZN(n3675) );
  NOR2_X1 U4409 ( .A1(n4114), .A2(n3819), .ZN(n3673) );
  AOI22_X1 U4410 ( .A1(n4261), .A2(n3794), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3671) );
  OAI21_X1 U4411 ( .B1(n3779), .B2(n4117), .A(n3671), .ZN(n3672) );
  AOI211_X1 U4412 ( .C1(n3987), .C2(n3792), .A(n3673), .B(n3672), .ZN(n3674)
         );
  OAI21_X1 U4413 ( .B1(n3675), .B2(n3800), .A(n3674), .ZN(U3211) );
  NAND2_X1 U4414 ( .A1(n3676), .A2(n3806), .ZN(n3684) );
  AOI21_X1 U4415 ( .B1(n3763), .B2(n3678), .A(n3677), .ZN(n3683) );
  OAI22_X1 U4416 ( .A1(n4305), .A2(n3808), .B1(n3779), .B2(n3679), .ZN(n3681)
         );
  INV_X1 U4417 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4691) );
  OAI22_X1 U4418 ( .A1(n4189), .A2(n3813), .B1(STATE_REG_SCAN_IN), .B2(n4691), 
        .ZN(n3680) );
  AOI211_X1 U4419 ( .C1(n4193), .C2(n3793), .A(n3681), .B(n3680), .ZN(n3682)
         );
  OAI21_X1 U4420 ( .B1(n3684), .B2(n3683), .A(n3682), .ZN(U3213) );
  INV_X1 U4421 ( .A(n3685), .ZN(n3686) );
  AOI21_X1 U4422 ( .B1(n3687), .B2(n2063), .A(n3686), .ZN(n3696) );
  OAI22_X1 U4423 ( .A1(n3779), .A2(n3688), .B1(n3735), .B2(n3808), .ZN(n3691)
         );
  NAND2_X1 U4424 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4077) );
  OAI21_X1 U4425 ( .B1(n3813), .B2(n3689), .A(n4077), .ZN(n3690) );
  NOR2_X1 U4426 ( .A1(n3691), .A2(n3690), .ZN(n3695) );
  INV_X1 U4427 ( .A(n3692), .ZN(n3693) );
  NAND2_X1 U4428 ( .A1(n3793), .A2(n3693), .ZN(n3694) );
  OAI211_X1 U4429 ( .C1(n3696), .C2(n3800), .A(n3695), .B(n3694), .ZN(U3216)
         );
  NAND2_X1 U4430 ( .A1(n2308), .A2(n3698), .ZN(n3701) );
  INV_X1 U4431 ( .A(n3753), .ZN(n3752) );
  OAI211_X1 U4432 ( .C1(n3699), .C2(n3752), .A(n3754), .B(n3701), .ZN(n3700)
         );
  OAI211_X1 U4433 ( .C1(n3702), .C2(n3701), .A(n3806), .B(n3700), .ZN(n3708)
         );
  NOR2_X1 U4434 ( .A1(n3779), .A2(n3703), .ZN(n3706) );
  OAI22_X1 U4435 ( .A1(n4305), .A2(n3813), .B1(STATE_REG_SCAN_IN), .B2(n3704), 
        .ZN(n3705) );
  AOI211_X1 U4436 ( .C1(n3794), .C2(n4301), .A(n3706), .B(n3705), .ZN(n3707)
         );
  OAI211_X1 U4437 ( .C1(n3819), .C2(n3709), .A(n3708), .B(n3707), .ZN(U3220)
         );
  NAND2_X1 U4438 ( .A1(n3711), .A2(n3710), .ZN(n3713) );
  XOR2_X1 U4439 ( .A(n3713), .B(n3712), .Z(n3717) );
  OAI22_X1 U4440 ( .A1(n4189), .A2(n3808), .B1(n3779), .B2(n4152), .ZN(n3715)
         );
  INV_X1 U4441 ( .A(n4261), .ZN(n4150) );
  OAI22_X1 U4442 ( .A1(n4150), .A2(n3813), .B1(STATE_REG_SCAN_IN), .B2(n4726), 
        .ZN(n3714) );
  AOI211_X1 U4443 ( .C1(n4153), .C2(n3793), .A(n3715), .B(n3714), .ZN(n3716)
         );
  OAI21_X1 U4444 ( .B1(n3717), .B2(n3800), .A(n3716), .ZN(U3222) );
  OAI21_X1 U4445 ( .B1(n3579), .B2(n3804), .A(n3802), .ZN(n3719) );
  XNOR2_X1 U4446 ( .A(n3719), .B(n3718), .ZN(n3720) );
  NAND2_X1 U4447 ( .A1(n3720), .A2(n3806), .ZN(n3725) );
  OAI22_X1 U4448 ( .A1(n3779), .A2(n3721), .B1(n4329), .B2(n3808), .ZN(n3723)
         );
  NAND2_X1 U4449 ( .A1(U3149), .A2(REG3_REG_16__SCAN_IN), .ZN(n4468) );
  OAI21_X1 U4450 ( .B1(n3813), .B2(n3777), .A(n4468), .ZN(n3722) );
  NOR2_X1 U4451 ( .A1(n3723), .A2(n3722), .ZN(n3724) );
  OAI211_X1 U4452 ( .C1(n3819), .C2(n3726), .A(n3725), .B(n3724), .ZN(U3223)
         );
  NAND2_X1 U4453 ( .A1(n3728), .A2(n3727), .ZN(n3732) );
  NAND2_X1 U4454 ( .A1(n3730), .A2(n3729), .ZN(n3731) );
  XNOR2_X1 U4455 ( .A(n3732), .B(n3731), .ZN(n3741) );
  OAI22_X1 U4456 ( .A1(n3779), .A2(n3733), .B1(n3812), .B2(n3808), .ZN(n3737)
         );
  AND2_X1 U4457 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4482) );
  INV_X1 U4458 ( .A(n4482), .ZN(n3734) );
  OAI21_X1 U4459 ( .B1(n3813), .B2(n3735), .A(n3734), .ZN(n3736) );
  NOR2_X1 U4460 ( .A1(n3737), .A2(n3736), .ZN(n3740) );
  NAND2_X1 U4461 ( .A1(n3793), .A2(n3738), .ZN(n3739) );
  OAI211_X1 U4462 ( .C1(n3741), .C2(n3800), .A(n3740), .B(n3739), .ZN(U3225)
         );
  NAND2_X1 U4463 ( .A1(n3743), .A2(n3742), .ZN(n3744) );
  XOR2_X1 U4464 ( .A(n3745), .B(n3744), .Z(n3750) );
  NOR2_X1 U4465 ( .A1(n3819), .A2(n4164), .ZN(n3748) );
  AOI22_X1 U4466 ( .A1(n4282), .A2(n3794), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n3746) );
  OAI21_X1 U4467 ( .B1(n3779), .B2(n4168), .A(n3746), .ZN(n3747) );
  AOI211_X1 U4468 ( .C1(n3792), .C2(n3988), .A(n3748), .B(n3747), .ZN(n3749)
         );
  OAI21_X1 U4469 ( .B1(n3750), .B2(n3800), .A(n3749), .ZN(U3226) );
  NOR2_X1 U4470 ( .A1(n3751), .A2(n3752), .ZN(n3756) );
  AOI21_X1 U4471 ( .B1(n3754), .B2(n3753), .A(n3699), .ZN(n3755) );
  OAI21_X1 U4472 ( .B1(n3756), .B2(n3755), .A(n3806), .ZN(n3762) );
  INV_X1 U4473 ( .A(n4223), .ZN(n3780) );
  OAI22_X1 U4474 ( .A1(n3779), .A2(n3757), .B1(n3780), .B2(n3808), .ZN(n3760)
         );
  NAND2_X1 U4475 ( .A1(n3792), .A2(n4202), .ZN(n3758) );
  OAI21_X1 U4476 ( .B1(STATE_REG_SCAN_IN), .B2(n4690), .A(n3758), .ZN(n3759)
         );
  NOR2_X1 U4477 ( .A1(n3760), .A2(n3759), .ZN(n3761) );
  OAI211_X1 U4478 ( .C1(n3819), .C2(n4232), .A(n3762), .B(n3761), .ZN(U3230)
         );
  INV_X1 U4479 ( .A(n3763), .ZN(n3764) );
  AOI21_X1 U4480 ( .B1(n3766), .B2(n3765), .A(n3764), .ZN(n3772) );
  INV_X1 U4481 ( .A(n4212), .ZN(n3770) );
  OAI22_X1 U4482 ( .A1(n2253), .A2(n3808), .B1(n3779), .B2(n4211), .ZN(n3769)
         );
  INV_X1 U4483 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3767) );
  OAI22_X1 U4484 ( .A1(n4204), .A2(n3813), .B1(STATE_REG_SCAN_IN), .B2(n3767), 
        .ZN(n3768) );
  AOI211_X1 U4485 ( .C1(n3770), .C2(n3793), .A(n3769), .B(n3768), .ZN(n3771)
         );
  OAI21_X1 U4486 ( .B1(n3772), .B2(n3800), .A(n3771), .ZN(U3232) );
  XNOR2_X1 U4487 ( .A(n3775), .B(n3774), .ZN(n3776) );
  XNOR2_X1 U4488 ( .A(n3773), .B(n3776), .ZN(n3786) );
  OAI22_X1 U4489 ( .A1(n3779), .A2(n3778), .B1(n3777), .B2(n3808), .ZN(n3782)
         );
  NAND2_X1 U4490 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4488) );
  OAI21_X1 U4491 ( .B1(n3813), .B2(n3780), .A(n4488), .ZN(n3781) );
  NOR2_X1 U4492 ( .A1(n3782), .A2(n3781), .ZN(n3785) );
  NAND2_X1 U4493 ( .A1(n3793), .A2(n3783), .ZN(n3784) );
  OAI211_X1 U4494 ( .C1(n3786), .C2(n3800), .A(n3785), .B(n3784), .ZN(U3235)
         );
  INV_X1 U4495 ( .A(n3787), .ZN(n3788) );
  NOR2_X1 U4496 ( .A1(n3789), .A2(n3788), .ZN(n3790) );
  XNOR2_X1 U4497 ( .A(n3791), .B(n3790), .ZN(n3801) );
  AOI22_X1 U4498 ( .A1(n4270), .A2(n3792), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n3798) );
  NAND2_X1 U4499 ( .A1(n4132), .A2(n3793), .ZN(n3797) );
  NAND2_X1 U4500 ( .A1(n3988), .A2(n3794), .ZN(n3796) );
  OR2_X1 U4501 ( .A1(n3779), .A2(n4134), .ZN(n3795) );
  OAI21_X1 U4502 ( .B1(n3801), .B2(n3800), .A(n3799), .ZN(U3237) );
  NAND2_X1 U4503 ( .A1(n3803), .A2(n3802), .ZN(n3805) );
  XNOR2_X1 U4504 ( .A(n3805), .B(n3804), .ZN(n3807) );
  NAND2_X1 U4505 ( .A1(n3807), .A2(n3806), .ZN(n3817) );
  OAI22_X1 U4506 ( .A1(n3779), .A2(n3810), .B1(n3809), .B2(n3808), .ZN(n3815)
         );
  AND2_X1 U4507 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4462) );
  INV_X1 U4508 ( .A(n4462), .ZN(n3811) );
  OAI21_X1 U4509 ( .B1(n3813), .B2(n3812), .A(n3811), .ZN(n3814) );
  NOR2_X1 U4510 ( .A1(n3815), .A2(n3814), .ZN(n3816) );
  OAI211_X1 U4511 ( .C1(n3819), .C2(n3818), .A(n3817), .B(n3816), .ZN(U3238)
         );
  INV_X1 U4512 ( .A(n3950), .ZN(n3825) );
  NAND2_X1 U4513 ( .A1(n3820), .A2(n3824), .ZN(n3948) );
  NOR3_X1 U4514 ( .A1(n3821), .A2(n3825), .A3(n3948), .ZN(n3823) );
  INV_X1 U4515 ( .A(n3822), .ZN(n3952) );
  OAI21_X1 U4516 ( .B1(n3823), .B2(n3952), .A(n3951), .ZN(n3833) );
  INV_X1 U4517 ( .A(n3824), .ZN(n3826) );
  AOI211_X1 U4518 ( .C1(n3828), .C2(n3827), .A(n3826), .B(n3825), .ZN(n3830)
         );
  OAI21_X1 U4519 ( .B1(n3830), .B2(n3829), .A(n3951), .ZN(n3832) );
  AND2_X1 U4520 ( .A1(n3832), .A2(n3831), .ZN(n3955) );
  NAND2_X1 U4521 ( .A1(n3833), .A2(n3955), .ZN(n3835) );
  NOR2_X1 U4522 ( .A1(n3865), .A2(n3834), .ZN(n3959) );
  OAI221_X1 U4523 ( .B1(n3836), .B2(n3958), .C1(n3836), .C2(n3835), .A(n3959), 
        .ZN(n3843) );
  OR2_X1 U4524 ( .A1(n3838), .A2(n3837), .ZN(n3849) );
  NAND2_X1 U4525 ( .A1(n2414), .A2(REG1_REG_31__SCAN_IN), .ZN(n3841) );
  NAND2_X1 U4526 ( .A1(n2413), .A2(REG0_REG_31__SCAN_IN), .ZN(n3840) );
  INV_X1 U4527 ( .A(REG2_REG_31__SCAN_IN), .ZN(n4088) );
  OR2_X1 U4528 ( .A1(n2393), .A2(n4088), .ZN(n3839) );
  INV_X1 U4529 ( .A(n4086), .ZN(n3985) );
  NOR2_X1 U4530 ( .A1(n2427), .A2(n4637), .ZN(n4087) );
  INV_X1 U4531 ( .A(n4087), .ZN(n4083) );
  AND2_X1 U4532 ( .A1(n3985), .A2(n4083), .ZN(n3969) );
  NOR2_X1 U4533 ( .A1(n2427), .A2(n4718), .ZN(n4245) );
  INV_X1 U4534 ( .A(n4245), .ZN(n3853) );
  NOR2_X1 U4535 ( .A1(n3986), .A2(n3853), .ZN(n3842) );
  NOR2_X1 U4536 ( .A1(n3969), .A2(n3842), .ZN(n3882) );
  OAI21_X1 U4537 ( .B1(n4252), .B2(n3844), .A(n3882), .ZN(n3848) );
  AOI211_X1 U4538 ( .C1(n4123), .C2(n3843), .A(n3849), .B(n3848), .ZN(n3852)
         );
  INV_X1 U4539 ( .A(n3960), .ZN(n3851) );
  NAND2_X1 U4540 ( .A1(n4252), .A2(n3844), .ZN(n3845) );
  AND2_X1 U4541 ( .A1(n3846), .A2(n3845), .ZN(n3963) );
  NAND3_X1 U4542 ( .A1(n4110), .A2(n3963), .A3(n3847), .ZN(n3850) );
  AOI21_X1 U4543 ( .B1(n3963), .B2(n3849), .A(n3848), .ZN(n3968) );
  AOI22_X1 U4544 ( .A1(n3852), .A2(n3851), .B1(n3850), .B2(n3968), .ZN(n3859)
         );
  NOR2_X1 U4545 ( .A1(n3985), .A2(n3853), .ZN(n3858) );
  INV_X1 U4546 ( .A(n3854), .ZN(n3857) );
  INV_X1 U4547 ( .A(n3986), .ZN(n3855) );
  NOR2_X1 U4548 ( .A1(n3855), .A2(n4245), .ZN(n3881) );
  OAI21_X1 U4549 ( .B1(n3881), .B2(n4086), .A(n4087), .ZN(n3856) );
  OAI211_X1 U4550 ( .C1(n3859), .C2(n3858), .A(n3857), .B(n3856), .ZN(n3976)
         );
  INV_X1 U4551 ( .A(n4093), .ZN(n3911) );
  NAND2_X1 U4552 ( .A1(n4124), .A2(n3860), .ZN(n4143) );
  INV_X1 U4553 ( .A(n4143), .ZN(n3910) );
  INV_X1 U4554 ( .A(n3861), .ZN(n3863) );
  OR2_X1 U4555 ( .A1(n3863), .A2(n3862), .ZN(n4129) );
  INV_X1 U4556 ( .A(n4129), .ZN(n3908) );
  INV_X1 U4557 ( .A(n4141), .ZN(n3864) );
  NOR2_X1 U4558 ( .A1(n3865), .A2(n3864), .ZN(n4161) );
  NAND2_X1 U4559 ( .A1(n3867), .A2(n3866), .ZN(n4183) );
  INV_X1 U4560 ( .A(n4183), .ZN(n3871) );
  NOR2_X1 U4561 ( .A1(n3869), .A2(n3868), .ZN(n3870) );
  NAND4_X1 U4562 ( .A1(n4161), .A2(n3871), .A3(n4208), .A4(n3870), .ZN(n3907)
         );
  INV_X1 U4563 ( .A(n3872), .ZN(n3876) );
  NOR2_X1 U4564 ( .A1(n4538), .A2(n3873), .ZN(n3874) );
  NAND4_X1 U4565 ( .A1(n3876), .A2(n2175), .A3(n3875), .A4(n3874), .ZN(n3906)
         );
  INV_X1 U4566 ( .A(n3877), .ZN(n3879) );
  AND2_X1 U4567 ( .A1(n3879), .A2(n3878), .ZN(n4225) );
  NOR2_X1 U4568 ( .A1(n3985), .A2(n4083), .ZN(n3880) );
  NOR2_X1 U4569 ( .A1(n3881), .A2(n3880), .ZN(n3970) );
  NAND4_X1 U4570 ( .A1(n3883), .A2(n4110), .A3(n3882), .A4(n3970), .ZN(n3884)
         );
  OR2_X1 U4571 ( .A1(n4384), .A2(n3884), .ZN(n3885) );
  NOR2_X1 U4572 ( .A1(n4225), .A2(n3885), .ZN(n3904) );
  NOR2_X1 U4573 ( .A1(n3887), .A2(n3886), .ZN(n3903) );
  AND4_X1 U4574 ( .A1(n3891), .A2(n3890), .A3(n3889), .A4(n3888), .ZN(n3902)
         );
  INV_X1 U4575 ( .A(n2659), .ZN(n3895) );
  NAND4_X1 U4576 ( .A1(n3895), .A2(n2106), .A3(n3894), .A4(n3893), .ZN(n3900)
         );
  NAND4_X1 U4577 ( .A1(n3898), .A2(n3897), .A3(n3896), .A4(n3053), .ZN(n3899)
         );
  NOR2_X1 U4578 ( .A1(n3900), .A2(n3899), .ZN(n3901) );
  NAND4_X1 U4579 ( .A1(n3904), .A2(n3903), .A3(n3902), .A4(n3901), .ZN(n3905)
         );
  NOR4_X1 U4580 ( .A1(n3908), .A2(n3907), .A3(n3906), .A4(n3905), .ZN(n3909)
         );
  NAND3_X1 U4581 ( .A1(n3911), .A2(n3910), .A3(n3909), .ZN(n3974) );
  NOR2_X1 U4582 ( .A1(n4255), .A2(n4260), .ZN(n3967) );
  INV_X1 U4583 ( .A(n3912), .ZN(n3915) );
  OAI211_X1 U4584 ( .C1(n3915), .C2(n4384), .A(n3914), .B(n3913), .ZN(n3916)
         );
  NAND3_X1 U4585 ( .A1(n3916), .A2(n2662), .A3(n2660), .ZN(n3919) );
  NAND3_X1 U4586 ( .A1(n3919), .A2(n3918), .A3(n3917), .ZN(n3922) );
  NAND3_X1 U4587 ( .A1(n3922), .A2(n3921), .A3(n3920), .ZN(n3924) );
  NAND3_X1 U4588 ( .A1(n3924), .A2(n3923), .A3(n2091), .ZN(n3928) );
  INV_X1 U4589 ( .A(n3925), .ZN(n3926) );
  AOI21_X1 U4590 ( .B1(n3928), .B2(n3927), .A(n3926), .ZN(n3934) );
  NAND2_X1 U4591 ( .A1(n3930), .A2(n3929), .ZN(n3933) );
  OAI211_X1 U4592 ( .C1(n3934), .C2(n3933), .A(n3932), .B(n3931), .ZN(n3937)
         );
  NAND3_X1 U4593 ( .A1(n3937), .A2(n3936), .A3(n3935), .ZN(n3939) );
  NAND2_X1 U4594 ( .A1(n3939), .A2(n3938), .ZN(n3945) );
  INV_X1 U4595 ( .A(n3940), .ZN(n3943) );
  INV_X1 U4596 ( .A(n3941), .ZN(n3942) );
  AOI211_X1 U4597 ( .C1(n3945), .C2(n3944), .A(n3943), .B(n3942), .ZN(n3949)
         );
  INV_X1 U4598 ( .A(n3946), .ZN(n3947) );
  NOR3_X1 U4599 ( .A1(n3949), .A2(n3948), .A3(n3947), .ZN(n3953) );
  OAI211_X1 U4600 ( .C1(n3953), .C2(n3952), .A(n3951), .B(n3950), .ZN(n3956)
         );
  NAND3_X1 U4601 ( .A1(n3956), .A2(n3955), .A3(n3954), .ZN(n3957) );
  NAND2_X1 U4602 ( .A1(n3958), .A2(n3957), .ZN(n3961) );
  AOI211_X1 U4603 ( .C1(n3962), .C2(n3961), .A(n3960), .B(n2100), .ZN(n3966)
         );
  INV_X1 U4604 ( .A(n3963), .ZN(n3964) );
  NOR4_X1 U4605 ( .A1(n3967), .A2(n3966), .A3(n3965), .A4(n3964), .ZN(n3972)
         );
  INV_X1 U4606 ( .A(n3968), .ZN(n3971) );
  OAI22_X1 U4607 ( .A1(n3972), .A2(n3971), .B1(n3970), .B2(n3969), .ZN(n3973)
         );
  MUX2_X1 U4608 ( .A(n3974), .B(n3973), .S(n2658), .Z(n3975) );
  NAND2_X1 U4609 ( .A1(n3976), .A2(n3975), .ZN(n3977) );
  XNOR2_X1 U4610 ( .A(n3977), .B(n4385), .ZN(n3984) );
  NAND2_X1 U4611 ( .A1(n3979), .A2(n3978), .ZN(n3980) );
  OAI211_X1 U4612 ( .C1(n3981), .C2(n3983), .A(n3980), .B(B_REG_SCAN_IN), .ZN(
        n3982) );
  OAI21_X1 U4613 ( .B1(n3984), .B2(n3983), .A(n3982), .ZN(U3239) );
  MUX2_X1 U4614 ( .A(DATAO_REG_31__SCAN_IN), .B(n3985), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4615 ( .A(DATAO_REG_30__SCAN_IN), .B(n3986), .S(U4043), .Z(U3580)
         );
  MUX2_X1 U4616 ( .A(DATAO_REG_29__SCAN_IN), .B(n4252), .S(U4043), .Z(U3579)
         );
  MUX2_X1 U4617 ( .A(DATAO_REG_28__SCAN_IN), .B(n3987), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4618 ( .A(DATAO_REG_27__SCAN_IN), .B(n4270), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4619 ( .A(DATAO_REG_26__SCAN_IN), .B(n4261), .S(U4043), .Z(U3576)
         );
  MUX2_X1 U4620 ( .A(DATAO_REG_25__SCAN_IN), .B(n3988), .S(U4043), .Z(U3575)
         );
  MUX2_X1 U4621 ( .A(DATAO_REG_24__SCAN_IN), .B(n4147), .S(U4043), .Z(U3574)
         );
  MUX2_X1 U4622 ( .A(DATAO_REG_23__SCAN_IN), .B(n4282), .S(n4000), .Z(U3573)
         );
  MUX2_X1 U4623 ( .A(DATAO_REG_22__SCAN_IN), .B(n4186), .S(n4000), .Z(U3572)
         );
  MUX2_X1 U4624 ( .A(DATAO_REG_21__SCAN_IN), .B(n4202), .S(n4000), .Z(U3571)
         );
  MUX2_X1 U4625 ( .A(DATAO_REG_20__SCAN_IN), .B(n4301), .S(n4000), .Z(U3570)
         );
  MUX2_X1 U4626 ( .A(DATAO_REG_19__SCAN_IN), .B(n4223), .S(n4000), .Z(U3569)
         );
  MUX2_X1 U4627 ( .A(DATAO_REG_18__SCAN_IN), .B(n3989), .S(n4000), .Z(U3568)
         );
  MUX2_X1 U4628 ( .A(DATAO_REG_17__SCAN_IN), .B(n4326), .S(n4000), .Z(U3567)
         );
  MUX2_X1 U4629 ( .A(DATAO_REG_16__SCAN_IN), .B(n3990), .S(n4000), .Z(U3566)
         );
  MUX2_X1 U4630 ( .A(DATAO_REG_15__SCAN_IN), .B(n3991), .S(n4000), .Z(U3565)
         );
  MUX2_X1 U4631 ( .A(DATAO_REG_14__SCAN_IN), .B(n3992), .S(n4000), .Z(U3564)
         );
  MUX2_X1 U4632 ( .A(DATAO_REG_13__SCAN_IN), .B(n3993), .S(n4000), .Z(U3563)
         );
  MUX2_X1 U4633 ( .A(DATAO_REG_12__SCAN_IN), .B(n3994), .S(n4000), .Z(U3562)
         );
  MUX2_X1 U4634 ( .A(DATAO_REG_11__SCAN_IN), .B(n3995), .S(n4000), .Z(U3561)
         );
  MUX2_X1 U4635 ( .A(DATAO_REG_10__SCAN_IN), .B(n3996), .S(n4000), .Z(U3560)
         );
  MUX2_X1 U4636 ( .A(DATAO_REG_9__SCAN_IN), .B(n3997), .S(U4043), .Z(U3559) );
  MUX2_X1 U4637 ( .A(DATAO_REG_8__SCAN_IN), .B(n3998), .S(n4000), .Z(U3558) );
  MUX2_X1 U4638 ( .A(DATAO_REG_7__SCAN_IN), .B(n3999), .S(n4000), .Z(U3557) );
  MUX2_X1 U4639 ( .A(DATAO_REG_6__SCAN_IN), .B(n4001), .S(n4000), .Z(U3556) );
  MUX2_X1 U4640 ( .A(DATAO_REG_5__SCAN_IN), .B(n4002), .S(U4043), .Z(U3555) );
  MUX2_X1 U4641 ( .A(DATAO_REG_4__SCAN_IN), .B(n4003), .S(U4043), .Z(U3554) );
  MUX2_X1 U4642 ( .A(DATAO_REG_3__SCAN_IN), .B(n4004), .S(U4043), .Z(U3553) );
  MUX2_X1 U4643 ( .A(DATAO_REG_2__SCAN_IN), .B(n4005), .S(U4043), .Z(U3552) );
  MUX2_X1 U4644 ( .A(DATAO_REG_1__SCAN_IN), .B(n2387), .S(U4043), .Z(U3551) );
  MUX2_X1 U4645 ( .A(DATAO_REG_0__SCAN_IN), .B(n2817), .S(U4043), .Z(U3550) );
  NAND2_X1 U4646 ( .A1(n4018), .A2(n4393), .ZN(n4017) );
  INV_X1 U4647 ( .A(n4007), .ZN(n4010) );
  MUX2_X1 U4648 ( .A(REG2_REG_1__SCAN_IN), .B(n2779), .S(n4393), .Z(n4009) );
  OAI211_X1 U4649 ( .C1(n4010), .C2(n4009), .A(n4440), .B(n4008), .ZN(n4016)
         );
  OAI211_X1 U4650 ( .C1(n4013), .C2(n4012), .A(n4495), .B(n4011), .ZN(n4015)
         );
  AOI22_X1 U4651 ( .A1(n4493), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4014) );
  NAND4_X1 U4652 ( .A1(n4017), .A2(n4016), .A3(n4015), .A4(n4014), .ZN(U3241)
         );
  NAND2_X1 U4653 ( .A1(n4018), .A2(n4391), .ZN(n4026) );
  OAI211_X1 U4654 ( .C1(REG1_REG_3__SCAN_IN), .C2(n4020), .A(n4495), .B(n4019), 
        .ZN(n4025) );
  AOI22_X1 U4655 ( .A1(n4493), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n4024) );
  XNOR2_X1 U4656 ( .A(n4021), .B(REG2_REG_3__SCAN_IN), .ZN(n4022) );
  NAND2_X1 U4657 ( .A1(n4440), .A2(n4022), .ZN(n4023) );
  NAND4_X1 U4658 ( .A1(n4026), .A2(n4025), .A3(n4024), .A4(n4023), .ZN(U3243)
         );
  MUX2_X1 U4659 ( .A(n3545), .B(REG2_REG_19__SCAN_IN), .S(n4078), .Z(n4042) );
  AOI22_X1 U4660 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4522), .B1(n4043), .B2(
        n2587), .ZN(n4491) );
  NOR2_X1 U4661 ( .A1(n4070), .A2(REG2_REG_17__SCAN_IN), .ZN(n4027) );
  AOI21_X1 U4662 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4070), .A(n4027), .ZN(n4480) );
  INV_X1 U4663 ( .A(n4046), .ZN(n4529) );
  NOR2_X1 U4664 ( .A1(n4439), .A2(n4529), .ZN(n4438) );
  NAND2_X1 U4665 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4047), .ZN(n4033) );
  AOI22_X1 U4666 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4047), .B1(n4532), .B2(
        n3271), .ZN(n4423) );
  NAND2_X1 U4667 ( .A1(n4049), .A2(REG2_REG_9__SCAN_IN), .ZN(n4030) );
  INV_X1 U4668 ( .A(n4049), .ZN(n4535) );
  AOI22_X1 U4669 ( .A1(n4049), .A2(REG2_REG_9__SCAN_IN), .B1(n2481), .B2(n4535), .ZN(n4403) );
  NAND2_X1 U4670 ( .A1(n4403), .A2(n4402), .ZN(n4401) );
  NAND2_X1 U4671 ( .A1(n4030), .A2(n4401), .ZN(n4031) );
  NAND2_X1 U4672 ( .A1(n4055), .A2(n4031), .ZN(n4032) );
  INV_X1 U4673 ( .A(n4055), .ZN(n4534) );
  XNOR2_X1 U4674 ( .A(n4031), .B(n4534), .ZN(n4410) );
  NAND2_X1 U4675 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4410), .ZN(n4409) );
  NAND2_X1 U4676 ( .A1(n4059), .A2(n4034), .ZN(n4035) );
  INV_X1 U4677 ( .A(n4059), .ZN(n4531) );
  NOR2_X1 U4678 ( .A1(n2120), .A2(n4036), .ZN(n4037) );
  NAND2_X1 U4679 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4044), .ZN(n4038) );
  OAI21_X1 U4680 ( .B1(REG2_REG_15__SCAN_IN), .B2(n4044), .A(n4038), .ZN(n4459) );
  INV_X1 U4681 ( .A(n4524), .ZN(n4477) );
  NAND2_X1 U4682 ( .A1(n4039), .A2(n4477), .ZN(n4040) );
  XOR2_X1 U4683 ( .A(n4042), .B(n4041), .Z(n4082) );
  INV_X1 U4684 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4072) );
  AOI22_X1 U4685 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4043), .B1(n4522), .B2(
        n4072), .ZN(n4496) );
  NOR2_X1 U4686 ( .A1(n4070), .A2(REG1_REG_17__SCAN_IN), .ZN(n4071) );
  NAND2_X1 U4687 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4044), .ZN(n4066) );
  INV_X1 U4688 ( .A(n4044), .ZN(n4526) );
  AOI22_X1 U4689 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4044), .B1(n4526), .B2(
        n3424), .ZN(n4465) );
  NAND2_X1 U4690 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4046), .ZN(n4062) );
  INV_X1 U4691 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4045) );
  AOI22_X1 U4692 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4046), .B1(n4529), .B2(
        n4045), .ZN(n4448) );
  NAND2_X1 U4693 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4047), .ZN(n4058) );
  AOI22_X1 U4694 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4047), .B1(n4532), .B2(
        n3332), .ZN(n4420) );
  NAND2_X1 U4695 ( .A1(n4049), .A2(REG1_REG_9__SCAN_IN), .ZN(n4054) );
  INV_X1 U4696 ( .A(REG1_REG_9__SCAN_IN), .ZN(n4048) );
  AOI22_X1 U4697 ( .A1(n4049), .A2(REG1_REG_9__SCAN_IN), .B1(n4048), .B2(n4535), .ZN(n4400) );
  INV_X1 U4698 ( .A(n4050), .ZN(n4386) );
  AOI22_X1 U4699 ( .A1(n4052), .A2(REG1_REG_8__SCAN_IN), .B1(n4386), .B2(n4051), .ZN(n4053) );
  INV_X1 U4700 ( .A(n4053), .ZN(n4399) );
  NAND2_X1 U4701 ( .A1(n4400), .A2(n4399), .ZN(n4398) );
  NAND2_X1 U4702 ( .A1(n4054), .A2(n4398), .ZN(n4056) );
  NAND2_X1 U4703 ( .A1(n4055), .A2(n4056), .ZN(n4057) );
  XNOR2_X1 U4704 ( .A(n4056), .B(n4534), .ZN(n4415) );
  NAND2_X1 U4705 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4415), .ZN(n4414) );
  NAND2_X1 U4706 ( .A1(n4059), .A2(n4060), .ZN(n4061) );
  NAND2_X1 U4707 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4435), .ZN(n4434) );
  NAND2_X1 U4708 ( .A1(n4063), .A2(n4064), .ZN(n4065) );
  NAND2_X1 U4709 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4456), .ZN(n4455) );
  NOR2_X1 U4710 ( .A1(n4524), .A2(n4067), .ZN(n4068) );
  INV_X1 U4711 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4069) );
  INV_X1 U4712 ( .A(n4070), .ZN(n4523) );
  AOI22_X1 U4713 ( .A1(n4070), .A2(n4069), .B1(REG1_REG_17__SCAN_IN), .B2(
        n4523), .ZN(n4483) );
  OAI21_X1 U4714 ( .B1(n4072), .B2(n4522), .A(n4494), .ZN(n4075) );
  INV_X1 U4715 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4073) );
  MUX2_X1 U4716 ( .A(REG1_REG_19__SCAN_IN), .B(n4073), .S(n4078), .Z(n4074) );
  XNOR2_X1 U4717 ( .A(n4075), .B(n4074), .ZN(n4080) );
  NAND2_X1 U4718 ( .A1(n4493), .A2(ADDR_REG_19__SCAN_IN), .ZN(n4076) );
  OAI211_X1 U4719 ( .C1(n4499), .C2(n4078), .A(n4077), .B(n4076), .ZN(n4079)
         );
  AOI21_X1 U4720 ( .B1(n4080), .B2(n4495), .A(n4079), .ZN(n4081) );
  OAI21_X1 U4721 ( .B1(n4082), .B2(n4489), .A(n4081), .ZN(U3259) );
  XNOR2_X1 U4722 ( .A(n4243), .B(n4083), .ZN(n4338) );
  INV_X1 U4723 ( .A(n4084), .ZN(n4085) );
  NOR2_X1 U4724 ( .A1(n4086), .A2(n4085), .ZN(n4247) );
  AOI21_X1 U4725 ( .B1(n4087), .B2(n4324), .A(n4247), .ZN(n4335) );
  MUX2_X1 U4726 ( .A(n4088), .B(n4335), .S(n4213), .Z(n4089) );
  OAI21_X1 U4727 ( .B1(n4338), .B2(n4195), .A(n4089), .ZN(U3260) );
  XOR2_X1 U4728 ( .A(n4093), .B(n4090), .Z(n4091) );
  NAND2_X1 U4729 ( .A1(n4091), .A2(n4231), .ZN(n4254) );
  XOR2_X1 U4730 ( .A(n4093), .B(n4092), .Z(n4257) );
  NAND2_X1 U4731 ( .A1(n4257), .A2(n4209), .ZN(n4104) );
  AND2_X1 U4732 ( .A1(n4112), .A2(n4251), .ZN(n4095) );
  OR2_X1 U4733 ( .A1(n4095), .A2(n4094), .ZN(n4345) );
  INV_X1 U4734 ( .A(n4345), .ZN(n4102) );
  AOI22_X1 U4735 ( .A1(n4096), .A2(n4511), .B1(REG2_REG_28__SCAN_IN), .B2(
        n4519), .ZN(n4097) );
  OAI21_X1 U4736 ( .B1(n4255), .B2(n4167), .A(n4097), .ZN(n4101) );
  OAI22_X1 U4737 ( .A1(n4099), .A2(n4170), .B1(n4098), .B2(n4169), .ZN(n4100)
         );
  AOI211_X1 U4738 ( .C1(n4102), .C2(n4513), .A(n4101), .B(n4100), .ZN(n4103)
         );
  OAI211_X1 U4739 ( .C1(n4519), .C2(n4254), .A(n4104), .B(n4103), .ZN(U3262)
         );
  AND2_X1 U4740 ( .A1(n4106), .A2(n4105), .ZN(n4107) );
  OR2_X1 U4741 ( .A1(n4108), .A2(n4107), .ZN(n4109) );
  NAND2_X1 U4742 ( .A1(n4109), .A2(n4231), .ZN(n4263) );
  XNOR2_X1 U4743 ( .A(n4111), .B(n4110), .ZN(n4266) );
  NAND2_X1 U4744 ( .A1(n4266), .A2(n4209), .ZN(n4122) );
  INV_X1 U4745 ( .A(n4130), .ZN(n4113) );
  OAI21_X1 U4746 ( .B1(n4113), .B2(n4117), .A(n4112), .ZN(n4349) );
  INV_X1 U4747 ( .A(n4349), .ZN(n4120) );
  INV_X1 U4748 ( .A(n4114), .ZN(n4115) );
  AOI22_X1 U4749 ( .A1(n4115), .A2(n4511), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4519), .ZN(n4116) );
  OAI21_X1 U4750 ( .B1(n4150), .B2(n4167), .A(n4116), .ZN(n4119) );
  OAI22_X1 U4751 ( .A1(n4264), .A2(n4170), .B1(n4117), .B2(n4169), .ZN(n4118)
         );
  AOI211_X1 U4752 ( .C1(n4120), .C2(n4513), .A(n4119), .B(n4118), .ZN(n4121)
         );
  OAI211_X1 U4753 ( .C1(n4519), .C2(n4263), .A(n4122), .B(n4121), .ZN(U3263)
         );
  NAND2_X1 U4754 ( .A1(n4142), .A2(n4123), .ZN(n4125) );
  NAND2_X1 U4755 ( .A1(n4125), .A2(n4124), .ZN(n4126) );
  XNOR2_X1 U4756 ( .A(n4126), .B(n4129), .ZN(n4127) );
  NAND2_X1 U4757 ( .A1(n4127), .A2(n4231), .ZN(n4272) );
  XOR2_X1 U4758 ( .A(n4129), .B(n4128), .Z(n4274) );
  NAND2_X1 U4759 ( .A1(n4274), .A2(n4209), .ZN(n4139) );
  INV_X1 U4760 ( .A(n4151), .ZN(n4131) );
  OAI21_X1 U4761 ( .B1(n4131), .B2(n4134), .A(n4130), .ZN(n4353) );
  INV_X1 U4762 ( .A(n4353), .ZN(n4137) );
  AOI22_X1 U4763 ( .A1(n4132), .A2(n4511), .B1(REG2_REG_26__SCAN_IN), .B2(
        n4519), .ZN(n4133) );
  OAI21_X1 U4764 ( .B1(n4255), .B2(n4170), .A(n4133), .ZN(n4136) );
  OAI22_X1 U4765 ( .A1(n4285), .A2(n4167), .B1(n4134), .B2(n4169), .ZN(n4135)
         );
  AOI211_X1 U4766 ( .C1(n4137), .C2(n4513), .A(n4136), .B(n4135), .ZN(n4138)
         );
  OAI211_X1 U4767 ( .C1(n4519), .C2(n4272), .A(n4139), .B(n4138), .ZN(U3264)
         );
  XNOR2_X1 U4768 ( .A(n4140), .B(n4143), .ZN(n4278) );
  INV_X1 U4769 ( .A(n4278), .ZN(n4157) );
  NAND2_X1 U4770 ( .A1(n4142), .A2(n4141), .ZN(n4144) );
  XNOR2_X1 U4771 ( .A(n4144), .B(n4143), .ZN(n4145) );
  NAND2_X1 U4772 ( .A1(n4145), .A2(n4231), .ZN(n4149) );
  AOI22_X1 U4773 ( .A1(n4147), .A2(n2048), .B1(n4146), .B2(n4324), .ZN(n4148)
         );
  OAI211_X1 U4774 ( .C1(n4150), .C2(n4304), .A(n4149), .B(n4148), .ZN(n4277)
         );
  OAI21_X1 U4775 ( .B1(n4162), .B2(n4152), .A(n4151), .ZN(n4357) );
  AOI22_X1 U4776 ( .A1(n4153), .A2(n4511), .B1(REG2_REG_25__SCAN_IN), .B2(
        n4519), .ZN(n4154) );
  OAI21_X1 U4777 ( .B1(n4357), .B2(n4195), .A(n4154), .ZN(n4155) );
  AOI21_X1 U4778 ( .B1(n4277), .B2(n4213), .A(n4155), .ZN(n4156) );
  OAI21_X1 U4779 ( .B1(n4157), .B2(n4198), .A(n4156), .ZN(U3265) );
  XNOR2_X1 U4780 ( .A(n4158), .B(n4161), .ZN(n4159) );
  NAND2_X1 U4781 ( .A1(n4159), .A2(n4231), .ZN(n4284) );
  XOR2_X1 U4782 ( .A(n4161), .B(n4160), .Z(n4287) );
  NAND2_X1 U4783 ( .A1(n4287), .A2(n4209), .ZN(n4175) );
  INV_X1 U4784 ( .A(n4162), .ZN(n4163) );
  OAI21_X1 U4785 ( .B1(n4191), .B2(n4168), .A(n4163), .ZN(n4361) );
  INV_X1 U4786 ( .A(n4361), .ZN(n4173) );
  INV_X1 U4787 ( .A(n4164), .ZN(n4165) );
  AOI22_X1 U4788 ( .A1(n4165), .A2(n4511), .B1(REG2_REG_24__SCAN_IN), .B2(
        n4519), .ZN(n4166) );
  OAI21_X1 U4789 ( .B1(n4204), .B2(n4167), .A(n4166), .ZN(n4172) );
  OAI22_X1 U4790 ( .A1(n4285), .A2(n4170), .B1(n4169), .B2(n4168), .ZN(n4171)
         );
  AOI211_X1 U4791 ( .C1(n4173), .C2(n4513), .A(n4172), .B(n4171), .ZN(n4174)
         );
  OAI211_X1 U4792 ( .C1(n4519), .C2(n4284), .A(n4175), .B(n4174), .ZN(U3266)
         );
  XNOR2_X1 U4793 ( .A(n4176), .B(n4183), .ZN(n4291) );
  INV_X1 U4794 ( .A(n4291), .ZN(n4199) );
  OR2_X1 U4795 ( .A1(n4178), .A2(n4177), .ZN(n4180) );
  NAND2_X1 U4796 ( .A1(n4180), .A2(n4179), .ZN(n4200) );
  INV_X1 U4797 ( .A(n4181), .ZN(n4182) );
  AOI21_X1 U4798 ( .B1(n4200), .B2(n4208), .A(n4182), .ZN(n4184) );
  XNOR2_X1 U4799 ( .A(n4184), .B(n4183), .ZN(n4185) );
  NAND2_X1 U4800 ( .A1(n4185), .A2(n4231), .ZN(n4188) );
  AOI22_X1 U4801 ( .A1(n4186), .A2(n2048), .B1(n4324), .B2(n4190), .ZN(n4187)
         );
  OAI211_X1 U4802 ( .C1(n4189), .C2(n4304), .A(n4188), .B(n4187), .ZN(n4290)
         );
  AND2_X1 U4803 ( .A1(n2050), .A2(n4190), .ZN(n4192) );
  OR2_X1 U4804 ( .A1(n4192), .A2(n4191), .ZN(n4365) );
  AOI22_X1 U4805 ( .A1(n4193), .A2(n4511), .B1(n4519), .B2(
        REG2_REG_23__SCAN_IN), .ZN(n4194) );
  OAI21_X1 U4806 ( .B1(n4365), .B2(n4195), .A(n4194), .ZN(n4196) );
  AOI21_X1 U4807 ( .B1(n4290), .B2(n4213), .A(n4196), .ZN(n4197) );
  OAI21_X1 U4808 ( .B1(n4199), .B2(n4198), .A(n4197), .ZN(U3267) );
  XNOR2_X1 U4809 ( .A(n4200), .B(n4208), .ZN(n4206) );
  AOI22_X1 U4810 ( .A1(n4202), .A2(n2048), .B1(n4201), .B2(n4324), .ZN(n4203)
         );
  OAI21_X1 U4811 ( .B1(n4204), .B2(n4304), .A(n4203), .ZN(n4205) );
  AOI21_X1 U4812 ( .B1(n4206), .B2(n4231), .A(n4205), .ZN(n4295) );
  NAND2_X1 U4813 ( .A1(n4207), .A2(n4208), .ZN(n4294) );
  NAND3_X1 U4814 ( .A1(n2075), .A2(n4209), .A3(n4294), .ZN(n4218) );
  OAI21_X1 U4815 ( .B1(n2151), .B2(n4211), .A(n2050), .ZN(n4369) );
  INV_X1 U4816 ( .A(n4369), .ZN(n4216) );
  OAI22_X1 U4817 ( .A1(n4214), .A2(n4213), .B1(n4212), .B2(n4500), .ZN(n4215)
         );
  AOI21_X1 U4818 ( .B1(n4216), .B2(n4513), .A(n4215), .ZN(n4217) );
  OAI211_X1 U4819 ( .C1(n4519), .C2(n4295), .A(n4218), .B(n4217), .ZN(U3268)
         );
  NAND2_X1 U4820 ( .A1(n4220), .A2(n4219), .ZN(n4222) );
  INV_X1 U4821 ( .A(n4225), .ZN(n4221) );
  XNOR2_X1 U4822 ( .A(n4222), .B(n4221), .ZN(n4230) );
  AOI22_X1 U4823 ( .A1(n4223), .A2(n2048), .B1(n4235), .B2(n4324), .ZN(n4224)
         );
  OAI21_X1 U4824 ( .B1(n2253), .B2(n4304), .A(n4224), .ZN(n4229) );
  XNOR2_X1 U4825 ( .A(n4226), .B(n4225), .ZN(n4314) );
  NOR2_X1 U4826 ( .A1(n4314), .A2(n4227), .ZN(n4228) );
  AOI211_X1 U4827 ( .C1(n4231), .C2(n4230), .A(n4229), .B(n4228), .ZN(n4313)
         );
  INV_X1 U4828 ( .A(n4232), .ZN(n4233) );
  AOI22_X1 U4829 ( .A1(n4519), .A2(REG2_REG_20__SCAN_IN), .B1(n4233), .B2(
        n4511), .ZN(n4237) );
  INV_X1 U4830 ( .A(n4234), .ZN(n4311) );
  NAND2_X1 U4831 ( .A1(n2074), .A2(n4235), .ZN(n4310) );
  NAND3_X1 U4832 ( .A1(n4311), .A2(n4513), .A3(n4310), .ZN(n4236) );
  OAI211_X1 U4833 ( .C1(n4314), .C2(n4238), .A(n4237), .B(n4236), .ZN(n4239)
         );
  INV_X1 U4834 ( .A(n4239), .ZN(n4240) );
  OAI21_X1 U4835 ( .B1(n4313), .B2(n4519), .A(n4240), .ZN(U3270) );
  NOR2_X1 U4836 ( .A1(n4335), .A2(n4565), .ZN(n4241) );
  AOI21_X1 U4837 ( .B1(REG1_REG_31__SCAN_IN), .B2(n4565), .A(n4241), .ZN(n4242) );
  OAI21_X1 U4838 ( .B1(n4338), .B2(n4319), .A(n4242), .ZN(U3549) );
  INV_X1 U4839 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4250) );
  NAND2_X1 U4840 ( .A1(n4395), .A2(n2746), .ZN(n4249) );
  AND2_X1 U4841 ( .A1(n4324), .A2(n4245), .ZN(n4246) );
  OR2_X1 U4842 ( .A1(n4247), .A2(n4246), .ZN(n4394) );
  NAND2_X1 U4843 ( .A1(n4394), .A2(n4568), .ZN(n4248) );
  OAI211_X1 U4844 ( .C1(n4568), .C2(n4250), .A(n4249), .B(n4248), .ZN(U3548)
         );
  INV_X1 U4845 ( .A(REG1_REG_28__SCAN_IN), .ZN(n4258) );
  AOI22_X1 U4846 ( .A1(n4252), .A2(n4325), .B1(n4251), .B2(n4324), .ZN(n4253)
         );
  OAI211_X1 U4847 ( .C1(n4255), .C2(n4328), .A(n4254), .B(n4253), .ZN(n4256)
         );
  AOI21_X1 U4848 ( .B1(n4257), .B2(n4316), .A(n4256), .ZN(n4342) );
  MUX2_X1 U4849 ( .A(n4258), .B(n4342), .S(n4568), .Z(n4259) );
  OAI21_X1 U4850 ( .B1(n4319), .B2(n4345), .A(n4259), .ZN(U3546) );
  INV_X1 U4851 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4267) );
  AOI22_X1 U4852 ( .A1(n4261), .A2(n2048), .B1(n4260), .B2(n4324), .ZN(n4262)
         );
  OAI211_X1 U4853 ( .C1(n4264), .C2(n4304), .A(n4263), .B(n4262), .ZN(n4265)
         );
  AOI21_X1 U4854 ( .B1(n4266), .B2(n4316), .A(n4265), .ZN(n4346) );
  MUX2_X1 U4855 ( .A(n4267), .B(n4346), .S(n4568), .Z(n4268) );
  OAI21_X1 U4856 ( .B1(n4319), .B2(n4349), .A(n4268), .ZN(U3545) );
  INV_X1 U4857 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4275) );
  AOI22_X1 U4858 ( .A1(n4270), .A2(n4325), .B1(n4324), .B2(n4269), .ZN(n4271)
         );
  OAI211_X1 U4859 ( .C1(n4285), .C2(n4328), .A(n4272), .B(n4271), .ZN(n4273)
         );
  AOI21_X1 U4860 ( .B1(n4274), .B2(n4316), .A(n4273), .ZN(n4350) );
  MUX2_X1 U4861 ( .A(n4275), .B(n4350), .S(n4568), .Z(n4276) );
  OAI21_X1 U4862 ( .B1(n4319), .B2(n4353), .A(n4276), .ZN(U3544) );
  INV_X1 U4863 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4279) );
  AOI21_X1 U4864 ( .B1(n4278), .B2(n4316), .A(n4277), .ZN(n4354) );
  MUX2_X1 U4865 ( .A(n4279), .B(n4354), .S(n4568), .Z(n4280) );
  OAI21_X1 U4866 ( .B1(n4319), .B2(n4357), .A(n4280), .ZN(U3543) );
  INV_X1 U4867 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4288) );
  AOI22_X1 U4868 ( .A1(n4282), .A2(n2048), .B1(n4324), .B2(n4281), .ZN(n4283)
         );
  OAI211_X1 U4869 ( .C1(n4285), .C2(n4304), .A(n4284), .B(n4283), .ZN(n4286)
         );
  AOI21_X1 U4870 ( .B1(n4287), .B2(n4316), .A(n4286), .ZN(n4358) );
  MUX2_X1 U4871 ( .A(n4288), .B(n4358), .S(n4568), .Z(n4289) );
  OAI21_X1 U4872 ( .B1(n4319), .B2(n4361), .A(n4289), .ZN(U3542) );
  INV_X1 U4873 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4292) );
  AOI21_X1 U4874 ( .B1(n4291), .B2(n4316), .A(n4290), .ZN(n4362) );
  MUX2_X1 U4875 ( .A(n4292), .B(n4362), .S(n4568), .Z(n4293) );
  OAI21_X1 U4876 ( .B1(n4319), .B2(n4365), .A(n4293), .ZN(U3541) );
  INV_X1 U4877 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4297) );
  NAND3_X1 U4878 ( .A1(n2075), .A2(n4316), .A3(n4294), .ZN(n4296) );
  AND2_X1 U4879 ( .A1(n4296), .A2(n4295), .ZN(n4366) );
  MUX2_X1 U4880 ( .A(n4297), .B(n4366), .S(n4568), .Z(n4298) );
  OAI21_X1 U4881 ( .B1(n4319), .B2(n4369), .A(n4298), .ZN(U3540) );
  INV_X1 U4882 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4308) );
  AOI22_X1 U4883 ( .A1(n4301), .A2(n2048), .B1(n4299), .B2(n4324), .ZN(n4302)
         );
  OAI211_X1 U4884 ( .C1(n4305), .C2(n4304), .A(n4303), .B(n4302), .ZN(n4306)
         );
  AOI21_X1 U4885 ( .B1(n4307), .B2(n4316), .A(n4306), .ZN(n4370) );
  MUX2_X1 U4886 ( .A(n4308), .B(n4370), .S(n4568), .Z(n4309) );
  OAI21_X1 U4887 ( .B1(n4319), .B2(n4373), .A(n4309), .ZN(U3539) );
  NAND3_X1 U4888 ( .A1(n4311), .A2(n2811), .A3(n4310), .ZN(n4312) );
  OAI211_X1 U4889 ( .C1(n4314), .C2(n4540), .A(n4313), .B(n4312), .ZN(n4374)
         );
  MUX2_X1 U4890 ( .A(REG1_REG_20__SCAN_IN), .B(n4374), .S(n4568), .Z(U3538) );
  AOI21_X1 U4891 ( .B1(n4317), .B2(n4316), .A(n4315), .ZN(n4375) );
  MUX2_X1 U4892 ( .A(n4073), .B(n4375), .S(n4568), .Z(n4318) );
  OAI21_X1 U4893 ( .B1(n4319), .B2(n4379), .A(n4318), .ZN(U3537) );
  OAI211_X1 U4894 ( .C1(n4322), .C2(n4551), .A(n4321), .B(n4320), .ZN(n4380)
         );
  MUX2_X1 U4895 ( .A(REG1_REG_18__SCAN_IN), .B(n4380), .S(n4568), .Z(U3536) );
  AOI22_X1 U4896 ( .A1(n4326), .A2(n4325), .B1(n4324), .B2(n4323), .ZN(n4327)
         );
  OAI21_X1 U4897 ( .B1(n4329), .B2(n4328), .A(n4327), .ZN(n4330) );
  AOI21_X1 U4898 ( .B1(n4331), .B2(n2811), .A(n4330), .ZN(n4333) );
  OAI211_X1 U4899 ( .C1(n4334), .C2(n4551), .A(n4333), .B(n4332), .ZN(n4381)
         );
  MUX2_X1 U4900 ( .A(REG1_REG_16__SCAN_IN), .B(n4381), .S(n4568), .Z(U3534) );
  NOR2_X1 U4901 ( .A1(n4335), .A2(n4557), .ZN(n4336) );
  AOI21_X1 U4902 ( .B1(REG0_REG_31__SCAN_IN), .B2(n4557), .A(n4336), .ZN(n4337) );
  OAI21_X1 U4903 ( .B1(n4338), .B2(n4378), .A(n4337), .ZN(U3517) );
  INV_X1 U4904 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4341) );
  NAND2_X1 U4905 ( .A1(n4395), .A2(n2739), .ZN(n4340) );
  NAND2_X1 U4906 ( .A1(n4394), .A2(n4559), .ZN(n4339) );
  OAI211_X1 U4907 ( .C1(n4559), .C2(n4341), .A(n4340), .B(n4339), .ZN(U3516)
         );
  INV_X1 U4908 ( .A(REG0_REG_28__SCAN_IN), .ZN(n4343) );
  MUX2_X1 U4909 ( .A(n4343), .B(n4342), .S(n4559), .Z(n4344) );
  OAI21_X1 U4910 ( .B1(n4345), .B2(n4378), .A(n4344), .ZN(U3514) );
  INV_X1 U4911 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4347) );
  MUX2_X1 U4912 ( .A(n4347), .B(n4346), .S(n4559), .Z(n4348) );
  OAI21_X1 U4913 ( .B1(n4349), .B2(n4378), .A(n4348), .ZN(U3513) );
  INV_X1 U4914 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4351) );
  MUX2_X1 U4915 ( .A(n4351), .B(n4350), .S(n4559), .Z(n4352) );
  OAI21_X1 U4916 ( .B1(n4353), .B2(n4378), .A(n4352), .ZN(U3512) );
  INV_X1 U4917 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4355) );
  MUX2_X1 U4918 ( .A(n4355), .B(n4354), .S(n4559), .Z(n4356) );
  OAI21_X1 U4919 ( .B1(n4357), .B2(n4378), .A(n4356), .ZN(U3511) );
  INV_X1 U4920 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4359) );
  MUX2_X1 U4921 ( .A(n4359), .B(n4358), .S(n4559), .Z(n4360) );
  OAI21_X1 U4922 ( .B1(n4361), .B2(n4378), .A(n4360), .ZN(U3510) );
  INV_X1 U4923 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4363) );
  MUX2_X1 U4924 ( .A(n4363), .B(n4362), .S(n4559), .Z(n4364) );
  OAI21_X1 U4925 ( .B1(n4365), .B2(n4378), .A(n4364), .ZN(U3509) );
  INV_X1 U4926 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4367) );
  MUX2_X1 U4927 ( .A(n4367), .B(n4366), .S(n4559), .Z(n4368) );
  OAI21_X1 U4928 ( .B1(n4369), .B2(n4378), .A(n4368), .ZN(U3508) );
  INV_X1 U4929 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4371) );
  MUX2_X1 U4930 ( .A(n4371), .B(n4370), .S(n4559), .Z(n4372) );
  OAI21_X1 U4931 ( .B1(n4373), .B2(n4378), .A(n4372), .ZN(U3507) );
  MUX2_X1 U4932 ( .A(REG0_REG_20__SCAN_IN), .B(n4374), .S(n4559), .Z(U3506) );
  MUX2_X1 U4933 ( .A(n4376), .B(n4375), .S(n4559), .Z(n4377) );
  OAI21_X1 U4934 ( .B1(n4379), .B2(n4378), .A(n4377), .ZN(U3505) );
  MUX2_X1 U4935 ( .A(REG0_REG_18__SCAN_IN), .B(n4380), .S(n4559), .Z(U3503) );
  MUX2_X1 U4936 ( .A(REG0_REG_16__SCAN_IN), .B(n4381), .S(n4559), .Z(U3499) );
  MUX2_X1 U4937 ( .A(n4382), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U4938 ( .A(n4383), .B(DATAI_25_), .S(U3149), .Z(U3327) );
  MUX2_X1 U4939 ( .A(n4384), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U4940 ( .A(DATAI_19_), .B(n4385), .S(STATE_REG_SCAN_IN), .Z(U3333)
         );
  MUX2_X1 U4941 ( .A(DATAI_8_), .B(n4386), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U4942 ( .A(n4387), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U4943 ( .A(n4388), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U4944 ( .A(n4389), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U4945 ( .A(DATAI_4_), .B(n4390), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4946 ( .A(n4391), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U4947 ( .A(n2049), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U4948 ( .A(n4393), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  INV_X1 U4949 ( .A(n4394), .ZN(n4397) );
  OAI21_X1 U4950 ( .B1(n4519), .B2(n4397), .A(n4396), .ZN(U3261) );
  OAI211_X1 U4951 ( .C1(n4400), .C2(n4399), .A(n4495), .B(n4398), .ZN(n4405)
         );
  OAI211_X1 U4952 ( .C1(n4403), .C2(n4402), .A(n4440), .B(n4401), .ZN(n4404)
         );
  OAI211_X1 U4953 ( .C1(n4499), .C2(n4535), .A(n4405), .B(n4404), .ZN(n4406)
         );
  AOI211_X1 U4954 ( .C1(n4493), .C2(ADDR_REG_9__SCAN_IN), .A(n4407), .B(n4406), 
        .ZN(n4408) );
  INV_X1 U4955 ( .A(n4408), .ZN(U3249) );
  OAI211_X1 U4956 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4410), .A(n4440), .B(n4409), .ZN(n4412) );
  NAND2_X1 U4957 ( .A1(n4412), .A2(n4411), .ZN(n4413) );
  AOI21_X1 U4958 ( .B1(n4493), .B2(ADDR_REG_10__SCAN_IN), .A(n4413), .ZN(n4417) );
  OAI211_X1 U4959 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4415), .A(n4495), .B(n4414), .ZN(n4416) );
  OAI211_X1 U4960 ( .C1(n4499), .C2(n4534), .A(n4417), .B(n4416), .ZN(U3250)
         );
  OAI211_X1 U4961 ( .C1(n4420), .C2(n4419), .A(n4495), .B(n4418), .ZN(n4425)
         );
  OAI211_X1 U4962 ( .C1(n4423), .C2(n4422), .A(n4440), .B(n4421), .ZN(n4424)
         );
  OAI211_X1 U4963 ( .C1(n4499), .C2(n4532), .A(n4425), .B(n4424), .ZN(n4426)
         );
  AOI211_X1 U4964 ( .C1(n4493), .C2(ADDR_REG_11__SCAN_IN), .A(n4427), .B(n4426), .ZN(n4428) );
  INV_X1 U4965 ( .A(n4428), .ZN(U3251) );
  OAI211_X1 U4966 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4430), .A(n4440), .B(n4429), .ZN(n4432) );
  NAND2_X1 U4967 ( .A1(n4432), .A2(n4431), .ZN(n4433) );
  AOI21_X1 U4968 ( .B1(n4493), .B2(ADDR_REG_12__SCAN_IN), .A(n4433), .ZN(n4437) );
  OAI211_X1 U4969 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4435), .A(n4495), .B(n4434), .ZN(n4436) );
  OAI211_X1 U4970 ( .C1(n4499), .C2(n4531), .A(n4437), .B(n4436), .ZN(U3252)
         );
  AOI21_X1 U4971 ( .B1(n4439), .B2(n4529), .A(n4438), .ZN(n4443) );
  OAI21_X1 U4972 ( .B1(n4443), .B2(n4442), .A(n4440), .ZN(n4441) );
  AOI21_X1 U4973 ( .B1(n4443), .B2(n4442), .A(n4441), .ZN(n4445) );
  AOI211_X1 U4974 ( .C1(n4493), .C2(ADDR_REG_13__SCAN_IN), .A(n4445), .B(n4444), .ZN(n4450) );
  OAI211_X1 U4975 ( .C1(n4448), .C2(n4447), .A(n4495), .B(n4446), .ZN(n4449)
         );
  OAI211_X1 U4976 ( .C1(n4499), .C2(n4529), .A(n4450), .B(n4449), .ZN(U3253)
         );
  AOI211_X1 U4977 ( .C1(n2534), .C2(n4452), .A(n4451), .B(n4489), .ZN(n4453)
         );
  AOI211_X1 U4978 ( .C1(n4493), .C2(ADDR_REG_14__SCAN_IN), .A(n4454), .B(n4453), .ZN(n4458) );
  OAI211_X1 U4979 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4456), .A(n4495), .B(n4455), .ZN(n4457) );
  OAI211_X1 U4980 ( .C1(n4499), .C2(n2120), .A(n4458), .B(n4457), .ZN(U3254)
         );
  AOI211_X1 U4981 ( .C1(n4460), .C2(n4459), .A(n2058), .B(n4489), .ZN(n4461)
         );
  AOI211_X1 U4982 ( .C1(n4493), .C2(ADDR_REG_15__SCAN_IN), .A(n4462), .B(n4461), .ZN(n4467) );
  OAI211_X1 U4983 ( .C1(n4465), .C2(n4464), .A(n4495), .B(n4463), .ZN(n4466)
         );
  OAI211_X1 U4984 ( .C1(n4499), .C2(n4526), .A(n4467), .B(n4466), .ZN(U3255)
         );
  INV_X1 U4985 ( .A(n4468), .ZN(n4472) );
  AOI221_X1 U4986 ( .B1(n4470), .B2(n4469), .C1(n2560), .C2(n4469), .A(n4489), 
        .ZN(n4471) );
  AOI211_X1 U4987 ( .C1(n4493), .C2(ADDR_REG_16__SCAN_IN), .A(n4472), .B(n4471), .ZN(n4476) );
  OAI221_X1 U4988 ( .B1(n4474), .B2(REG1_REG_16__SCAN_IN), .C1(n4474), .C2(
        n4473), .A(n4495), .ZN(n4475) );
  OAI211_X1 U4989 ( .C1(n4499), .C2(n4477), .A(n4476), .B(n4475), .ZN(U3256)
         );
  AOI221_X1 U4990 ( .B1(n4480), .B2(n4479), .C1(n4478), .C2(n4479), .A(n4489), 
        .ZN(n4481) );
  AOI211_X1 U4991 ( .C1(n4493), .C2(ADDR_REG_17__SCAN_IN), .A(n4482), .B(n4481), .ZN(n4487) );
  OAI221_X1 U4992 ( .B1(n4485), .B2(n4484), .C1(n4485), .C2(n4483), .A(n4495), 
        .ZN(n4486) );
  OAI211_X1 U4993 ( .C1(n4499), .C2(n4523), .A(n4487), .B(n4486), .ZN(U3257)
         );
  INV_X1 U4994 ( .A(n4488), .ZN(n4492) );
  OAI211_X1 U4995 ( .C1(n4496), .C2(n2072), .A(n4495), .B(n4494), .ZN(n4497)
         );
  OAI211_X1 U4996 ( .C1(n4499), .C2(n4522), .A(n4498), .B(n4497), .ZN(U3258)
         );
  OAI22_X1 U4997 ( .A1(n4213), .A2(n4502), .B1(n4501), .B2(n4500), .ZN(n4503)
         );
  INV_X1 U4998 ( .A(n4503), .ZN(n4509) );
  INV_X1 U4999 ( .A(n4504), .ZN(n4507) );
  INV_X1 U5000 ( .A(n4505), .ZN(n4506) );
  AOI22_X1 U5001 ( .A1(n4507), .A2(n4514), .B1(n4513), .B2(n4506), .ZN(n4508)
         );
  OAI211_X1 U5002 ( .C1(n4519), .C2(n4510), .A(n4509), .B(n4508), .ZN(U3282)
         );
  AOI22_X1 U5003 ( .A1(REG2_REG_2__SCAN_IN), .A2(n4519), .B1(
        REG3_REG_2__SCAN_IN), .B2(n4511), .ZN(n4517) );
  AOI22_X1 U5004 ( .A1(n4515), .A2(n4514), .B1(n4513), .B2(n4512), .ZN(n4516)
         );
  OAI211_X1 U5005 ( .C1(n4519), .C2(n4518), .A(n4517), .B(n4516), .ZN(U3288)
         );
  AND2_X1 U5006 ( .A1(D_REG_31__SCAN_IN), .A2(n4520), .ZN(U3291) );
  AND2_X1 U5007 ( .A1(D_REG_30__SCAN_IN), .A2(n4520), .ZN(U3292) );
  AND2_X1 U5008 ( .A1(D_REG_29__SCAN_IN), .A2(n4520), .ZN(U3293) );
  AND2_X1 U5009 ( .A1(D_REG_28__SCAN_IN), .A2(n4520), .ZN(U3294) );
  AND2_X1 U5010 ( .A1(D_REG_27__SCAN_IN), .A2(n4520), .ZN(U3295) );
  AND2_X1 U5011 ( .A1(D_REG_26__SCAN_IN), .A2(n4520), .ZN(U3296) );
  AND2_X1 U5012 ( .A1(D_REG_25__SCAN_IN), .A2(n4520), .ZN(U3297) );
  AND2_X1 U5013 ( .A1(D_REG_24__SCAN_IN), .A2(n4520), .ZN(U3298) );
  AND2_X1 U5014 ( .A1(D_REG_23__SCAN_IN), .A2(n4520), .ZN(U3299) );
  AND2_X1 U5015 ( .A1(D_REG_22__SCAN_IN), .A2(n4520), .ZN(U3300) );
  AND2_X1 U5016 ( .A1(D_REG_21__SCAN_IN), .A2(n4520), .ZN(U3301) );
  AND2_X1 U5017 ( .A1(D_REG_20__SCAN_IN), .A2(n4520), .ZN(U3302) );
  AND2_X1 U5018 ( .A1(D_REG_19__SCAN_IN), .A2(n4520), .ZN(U3303) );
  AND2_X1 U5019 ( .A1(D_REG_18__SCAN_IN), .A2(n4520), .ZN(U3304) );
  AND2_X1 U5020 ( .A1(D_REG_17__SCAN_IN), .A2(n4520), .ZN(U3305) );
  AND2_X1 U5021 ( .A1(D_REG_16__SCAN_IN), .A2(n4520), .ZN(U3306) );
  AND2_X1 U5022 ( .A1(D_REG_15__SCAN_IN), .A2(n4520), .ZN(U3307) );
  AND2_X1 U5023 ( .A1(D_REG_14__SCAN_IN), .A2(n4520), .ZN(U3308) );
  AND2_X1 U5024 ( .A1(D_REG_13__SCAN_IN), .A2(n4520), .ZN(U3309) );
  AND2_X1 U5025 ( .A1(D_REG_12__SCAN_IN), .A2(n4520), .ZN(U3310) );
  AND2_X1 U5026 ( .A1(D_REG_11__SCAN_IN), .A2(n4520), .ZN(U3311) );
  AND2_X1 U5027 ( .A1(D_REG_10__SCAN_IN), .A2(n4520), .ZN(U3312) );
  AND2_X1 U5028 ( .A1(D_REG_9__SCAN_IN), .A2(n4520), .ZN(U3313) );
  AND2_X1 U5029 ( .A1(D_REG_8__SCAN_IN), .A2(n4520), .ZN(U3314) );
  AND2_X1 U5030 ( .A1(D_REG_7__SCAN_IN), .A2(n4520), .ZN(U3315) );
  AND2_X1 U5031 ( .A1(D_REG_6__SCAN_IN), .A2(n4520), .ZN(U3316) );
  AND2_X1 U5032 ( .A1(D_REG_5__SCAN_IN), .A2(n4520), .ZN(U3317) );
  AND2_X1 U5033 ( .A1(D_REG_4__SCAN_IN), .A2(n4520), .ZN(U3318) );
  AND2_X1 U5034 ( .A1(D_REG_3__SCAN_IN), .A2(n4520), .ZN(U3319) );
  AND2_X1 U5035 ( .A1(D_REG_2__SCAN_IN), .A2(n4520), .ZN(U3320) );
  AOI21_X1 U5036 ( .B1(U3149), .B2(n4684), .A(n4521), .ZN(U3329) );
  AOI22_X1 U5037 ( .A1(STATE_REG_SCAN_IN), .A2(n4522), .B1(n2595), .B2(U3149), 
        .ZN(U3334) );
  INV_X1 U5038 ( .A(DATAI_17_), .ZN(n4723) );
  AOI22_X1 U5039 ( .A1(STATE_REG_SCAN_IN), .A2(n4523), .B1(n4723), .B2(U3149), 
        .ZN(U3335) );
  OAI22_X1 U5040 ( .A1(U3149), .A2(n4524), .B1(DATAI_16_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4525) );
  INV_X1 U5041 ( .A(n4525), .ZN(U3336) );
  INV_X1 U5042 ( .A(DATAI_15_), .ZN(n4676) );
  AOI22_X1 U5043 ( .A1(STATE_REG_SCAN_IN), .A2(n4526), .B1(n4676), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U5044 ( .A(DATAI_14_), .ZN(n4527) );
  AOI22_X1 U5045 ( .A1(STATE_REG_SCAN_IN), .A2(n2120), .B1(n4527), .B2(U3149), 
        .ZN(U3338) );
  INV_X1 U5046 ( .A(DATAI_13_), .ZN(n4528) );
  AOI22_X1 U5047 ( .A1(STATE_REG_SCAN_IN), .A2(n4529), .B1(n4528), .B2(U3149), 
        .ZN(U3339) );
  INV_X1 U5048 ( .A(DATAI_12_), .ZN(n4530) );
  AOI22_X1 U5049 ( .A1(STATE_REG_SCAN_IN), .A2(n4531), .B1(n4530), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U5050 ( .A(DATAI_11_), .ZN(n4609) );
  AOI22_X1 U5051 ( .A1(STATE_REG_SCAN_IN), .A2(n4532), .B1(n4609), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5052 ( .A(DATAI_10_), .ZN(n4533) );
  AOI22_X1 U5053 ( .A1(STATE_REG_SCAN_IN), .A2(n4534), .B1(n4533), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5054 ( .A(DATAI_9_), .ZN(n4588) );
  AOI22_X1 U5055 ( .A1(STATE_REG_SCAN_IN), .A2(n4535), .B1(n4588), .B2(U3149), 
        .ZN(U3343) );
  AOI211_X1 U5056 ( .C1(n4548), .C2(n4538), .A(n4537), .B(n4536), .ZN(n4561)
         );
  INV_X1 U5057 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4539) );
  AOI22_X1 U5058 ( .A1(n4559), .A2(n4561), .B1(n4539), .B2(n4557), .ZN(U3467)
         );
  NOR2_X1 U5059 ( .A1(n4541), .A2(n4540), .ZN(n4543) );
  AOI211_X1 U5060 ( .C1(n2811), .C2(n4544), .A(n4543), .B(n4542), .ZN(n4562)
         );
  INV_X1 U5061 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4545) );
  AOI22_X1 U5062 ( .A1(n4559), .A2(n4562), .B1(n4545), .B2(n4557), .ZN(U3469)
         );
  AOI211_X1 U5063 ( .C1(n4549), .C2(n4548), .A(n4547), .B(n4546), .ZN(n4564)
         );
  INV_X1 U5064 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4550) );
  AOI22_X1 U5065 ( .A1(n4559), .A2(n4564), .B1(n4550), .B2(n4557), .ZN(U3475)
         );
  NOR2_X1 U5066 ( .A1(n4552), .A2(n4551), .ZN(n4556) );
  AOI211_X1 U5067 ( .C1(n4556), .C2(n4555), .A(n4554), .B(n4553), .ZN(n4567)
         );
  INV_X1 U5068 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4558) );
  AOI22_X1 U5069 ( .A1(n4559), .A2(n4567), .B1(n4558), .B2(n4557), .ZN(U3481)
         );
  AOI22_X1 U5070 ( .A1(n4568), .A2(n4561), .B1(n4560), .B2(n4565), .ZN(U3518)
         );
  AOI22_X1 U5071 ( .A1(n4568), .A2(n4562), .B1(n2787), .B2(n4565), .ZN(U3519)
         );
  INV_X1 U5072 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4563) );
  AOI22_X1 U5073 ( .A1(n4568), .A2(n4564), .B1(n4563), .B2(n4565), .ZN(U3522)
         );
  AOI22_X1 U5074 ( .A1(n4568), .A2(n4567), .B1(n4566), .B2(n4565), .ZN(U3525)
         );
  AOI22_X1 U5075 ( .A1(STATE_REG_SCAN_IN), .A2(IR_REG_0__SCAN_IN), .B1(
        DATAI_0_), .B2(U3149), .ZN(n4761) );
  AOI22_X1 U5076 ( .A1(n2433), .A2(keyinput_g47), .B1(keyinput_g9), .B2(n4571), 
        .ZN(n4570) );
  OAI221_X1 U5077 ( .B1(n2433), .B2(keyinput_g47), .C1(n4571), .C2(keyinput_g9), .A(n4570), .ZN(n4581) );
  AOI22_X1 U5078 ( .A1(n4574), .A2(keyinput_g54), .B1(n4573), .B2(keyinput_g48), .ZN(n4572) );
  OAI221_X1 U5079 ( .B1(n4574), .B2(keyinput_g54), .C1(n4573), .C2(
        keyinput_g48), .A(n4572), .ZN(n4580) );
  XNOR2_X1 U5080 ( .A(DATAI_25_), .B(keyinput_g6), .ZN(n4578) );
  XNOR2_X1 U5081 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_g50), .ZN(n4577) );
  XNOR2_X1 U5082 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_g52), .ZN(n4576) );
  XNOR2_X1 U5083 ( .A(DATAI_0_), .B(keyinput_g31), .ZN(n4575) );
  NAND4_X1 U5084 ( .A1(n4578), .A2(n4577), .A3(n4576), .A4(n4575), .ZN(n4579)
         );
  NOR3_X1 U5085 ( .A1(n4581), .A2(n4580), .A3(n4579), .ZN(n4619) );
  INV_X1 U5086 ( .A(DATAI_6_), .ZN(n4583) );
  AOI22_X1 U5087 ( .A1(n4584), .A2(keyinput_g2), .B1(keyinput_g25), .B2(n4583), 
        .ZN(n4582) );
  OAI221_X1 U5088 ( .B1(n4584), .B2(keyinput_g2), .C1(n4583), .C2(keyinput_g25), .A(n4582), .ZN(n4594) );
  AOI22_X1 U5089 ( .A1(n4677), .A2(keyinput_g51), .B1(keyinput_g4), .B2(n2353), 
        .ZN(n4585) );
  OAI221_X1 U5090 ( .B1(n4677), .B2(keyinput_g51), .C1(n2353), .C2(keyinput_g4), .A(n4585), .ZN(n4593) );
  INV_X1 U5091 ( .A(DATAI_26_), .ZN(n4587) );
  AOI22_X1 U5092 ( .A1(n4588), .A2(keyinput_g22), .B1(n4587), .B2(keyinput_g5), 
        .ZN(n4586) );
  OAI221_X1 U5093 ( .B1(n4588), .B2(keyinput_g22), .C1(n4587), .C2(keyinput_g5), .A(n4586), .ZN(n4592) );
  XNOR2_X1 U5094 ( .A(IR_REG_0__SCAN_IN), .B(keyinput_g55), .ZN(n4590) );
  XNOR2_X1 U5095 ( .A(DATAI_15_), .B(keyinput_g16), .ZN(n4589) );
  NAND2_X1 U5096 ( .A1(n4590), .A2(n4589), .ZN(n4591) );
  NOR4_X1 U5097 ( .A1(n4594), .A2(n4593), .A3(n4592), .A4(n4591), .ZN(n4618)
         );
  AOI22_X1 U5098 ( .A1(n4724), .A2(keyinput_g44), .B1(n4596), .B2(keyinput_g49), .ZN(n4595) );
  OAI221_X1 U5099 ( .B1(n4724), .B2(keyinput_g44), .C1(n4596), .C2(
        keyinput_g49), .A(n4595), .ZN(n4605) );
  AOI22_X1 U5100 ( .A1(n2610), .A2(keyinput_g11), .B1(n4598), .B2(keyinput_g39), .ZN(n4597) );
  OAI221_X1 U5101 ( .B1(n2610), .B2(keyinput_g11), .C1(n4598), .C2(
        keyinput_g39), .A(n4597), .ZN(n4604) );
  AOI22_X1 U5102 ( .A1(n4693), .A2(keyinput_g26), .B1(n4690), .B2(keyinput_g53), .ZN(n4599) );
  OAI221_X1 U5103 ( .B1(n4693), .B2(keyinput_g26), .C1(n4690), .C2(
        keyinput_g53), .A(n4599), .ZN(n4603) );
  XNOR2_X1 U5104 ( .A(IR_REG_3__SCAN_IN), .B(keyinput_g58), .ZN(n4601) );
  XNOR2_X1 U5105 ( .A(REG3_REG_23__SCAN_IN), .B(keyinput_g36), .ZN(n4600) );
  NAND2_X1 U5106 ( .A1(n4601), .A2(n4600), .ZN(n4602) );
  NOR4_X1 U5107 ( .A1(n4605), .A2(n4604), .A3(n4603), .A4(n4602), .ZN(n4617)
         );
  AOI22_X1 U5108 ( .A1(n3704), .A2(keyinput_g43), .B1(keyinput_g35), .B2(n4694), .ZN(n4606) );
  OAI221_X1 U5109 ( .B1(n3704), .B2(keyinput_g43), .C1(n4694), .C2(
        keyinput_g35), .A(n4606), .ZN(n4615) );
  AOI22_X1 U5110 ( .A1(n4718), .A2(keyinput_g1), .B1(n2595), .B2(keyinput_g13), 
        .ZN(n4607) );
  OAI221_X1 U5111 ( .B1(n4718), .B2(keyinput_g1), .C1(n2595), .C2(keyinput_g13), .A(n4607), .ZN(n4614) );
  AOI22_X1 U5112 ( .A1(n4609), .A2(keyinput_g20), .B1(n4723), .B2(keyinput_g14), .ZN(n4608) );
  OAI221_X1 U5113 ( .B1(n4609), .B2(keyinput_g20), .C1(n4723), .C2(
        keyinput_g14), .A(n4608), .ZN(n4613) );
  XNOR2_X1 U5114 ( .A(IR_REG_1__SCAN_IN), .B(keyinput_g56), .ZN(n4611) );
  XNOR2_X1 U5115 ( .A(REG3_REG_25__SCAN_IN), .B(keyinput_g45), .ZN(n4610) );
  NAND2_X1 U5116 ( .A1(n4611), .A2(n4610), .ZN(n4612) );
  NOR4_X1 U5117 ( .A1(n4615), .A2(n4614), .A3(n4613), .A4(n4612), .ZN(n4616)
         );
  NAND4_X1 U5118 ( .A1(n4619), .A2(n4618), .A3(n4617), .A4(n4616), .ZN(n4759)
         );
  AOI22_X1 U5119 ( .A1(DATAI_14_), .A2(keyinput_g17), .B1(DATAI_16_), .B2(
        keyinput_g15), .ZN(n4620) );
  OAI221_X1 U5120 ( .B1(DATAI_14_), .B2(keyinput_g17), .C1(DATAI_16_), .C2(
        keyinput_g15), .A(n4620), .ZN(n4627) );
  AOI22_X1 U5121 ( .A1(REG3_REG_1__SCAN_IN), .A2(keyinput_g42), .B1(DATAI_19_), 
        .B2(keyinput_g12), .ZN(n4621) );
  OAI221_X1 U5122 ( .B1(REG3_REG_1__SCAN_IN), .B2(keyinput_g42), .C1(DATAI_19_), .C2(keyinput_g12), .A(n4621), .ZN(n4626) );
  AOI22_X1 U5123 ( .A1(DATAI_7_), .A2(keyinput_g24), .B1(DATAI_13_), .B2(
        keyinput_g18), .ZN(n4622) );
  OAI221_X1 U5124 ( .B1(DATAI_7_), .B2(keyinput_g24), .C1(DATAI_13_), .C2(
        keyinput_g18), .A(n4622), .ZN(n4625) );
  AOI22_X1 U5125 ( .A1(DATAI_10_), .A2(keyinput_g21), .B1(DATAI_12_), .B2(
        keyinput_g19), .ZN(n4623) );
  OAI221_X1 U5126 ( .B1(DATAI_10_), .B2(keyinput_g21), .C1(DATAI_12_), .C2(
        keyinput_g19), .A(n4623), .ZN(n4624) );
  NOR4_X1 U5127 ( .A1(n4627), .A2(n4626), .A3(n4625), .A4(n4624), .ZN(n4656)
         );
  XOR2_X1 U5128 ( .A(REG3_REG_28__SCAN_IN), .B(keyinput_g40), .Z(n4634) );
  AOI22_X1 U5129 ( .A1(DATAI_1_), .A2(keyinput_g30), .B1(STATE_REG_SCAN_IN), 
        .B2(keyinput_g32), .ZN(n4628) );
  OAI221_X1 U5130 ( .B1(DATAI_1_), .B2(keyinput_g30), .C1(STATE_REG_SCAN_IN), 
        .C2(keyinput_g32), .A(n4628), .ZN(n4633) );
  AOI22_X1 U5131 ( .A1(DATAI_21_), .A2(keyinput_g10), .B1(DATAI_28_), .B2(
        keyinput_g3), .ZN(n4629) );
  OAI221_X1 U5132 ( .B1(DATAI_21_), .B2(keyinput_g10), .C1(DATAI_28_), .C2(
        keyinput_g3), .A(n4629), .ZN(n4632) );
  AOI22_X1 U5133 ( .A1(DATAI_24_), .A2(keyinput_g7), .B1(DATAI_2_), .B2(
        keyinput_g29), .ZN(n4630) );
  OAI221_X1 U5134 ( .B1(DATAI_24_), .B2(keyinput_g7), .C1(DATAI_2_), .C2(
        keyinput_g29), .A(n4630), .ZN(n4631) );
  NOR4_X1 U5135 ( .A1(n4634), .A2(n4633), .A3(n4632), .A4(n4631), .ZN(n4655)
         );
  AOI22_X1 U5136 ( .A1(REG3_REG_8__SCAN_IN), .A2(keyinput_g41), .B1(
        REG3_REG_16__SCAN_IN), .B2(keyinput_g46), .ZN(n4635) );
  OAI221_X1 U5137 ( .B1(REG3_REG_8__SCAN_IN), .B2(keyinput_g41), .C1(
        REG3_REG_16__SCAN_IN), .C2(keyinput_g46), .A(n4635), .ZN(n4644) );
  AOI22_X1 U5138 ( .A1(n4637), .A2(keyinput_g0), .B1(n4684), .B2(keyinput_g8), 
        .ZN(n4636) );
  OAI221_X1 U5139 ( .B1(n4637), .B2(keyinput_g0), .C1(n4684), .C2(keyinput_g8), 
        .A(n4636), .ZN(n4643) );
  AOI22_X1 U5140 ( .A1(REG3_REG_10__SCAN_IN), .A2(keyinput_g37), .B1(
        REG3_REG_27__SCAN_IN), .B2(keyinput_g34), .ZN(n4638) );
  OAI221_X1 U5141 ( .B1(REG3_REG_10__SCAN_IN), .B2(keyinput_g37), .C1(
        REG3_REG_27__SCAN_IN), .C2(keyinput_g34), .A(n4638), .ZN(n4642) );
  XNOR2_X1 U5142 ( .A(IR_REG_6__SCAN_IN), .B(keyinput_g61), .ZN(n4640) );
  XNOR2_X1 U5143 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput_g38), .ZN(n4639) );
  NAND2_X1 U5144 ( .A1(n4640), .A2(n4639), .ZN(n4641) );
  NOR4_X1 U5145 ( .A1(n4644), .A2(n4643), .A3(n4642), .A4(n4641), .ZN(n4654)
         );
  AOI22_X1 U5146 ( .A1(DATAI_3_), .A2(keyinput_g28), .B1(IR_REG_2__SCAN_IN), 
        .B2(keyinput_g57), .ZN(n4645) );
  OAI221_X1 U5147 ( .B1(DATAI_3_), .B2(keyinput_g28), .C1(IR_REG_2__SCAN_IN), 
        .C2(keyinput_g57), .A(n4645), .ZN(n4652) );
  AOI22_X1 U5148 ( .A1(REG3_REG_7__SCAN_IN), .A2(keyinput_g33), .B1(
        IR_REG_7__SCAN_IN), .B2(keyinput_g62), .ZN(n4646) );
  OAI221_X1 U5149 ( .B1(REG3_REG_7__SCAN_IN), .B2(keyinput_g33), .C1(
        IR_REG_7__SCAN_IN), .C2(keyinput_g62), .A(n4646), .ZN(n4651) );
  AOI22_X1 U5150 ( .A1(DATAI_8_), .A2(keyinput_g23), .B1(IR_REG_8__SCAN_IN), 
        .B2(keyinput_g63), .ZN(n4647) );
  OAI221_X1 U5151 ( .B1(DATAI_8_), .B2(keyinput_g23), .C1(IR_REG_8__SCAN_IN), 
        .C2(keyinput_g63), .A(n4647), .ZN(n4650) );
  AOI22_X1 U5152 ( .A1(DATAI_4_), .A2(keyinput_g27), .B1(IR_REG_4__SCAN_IN), 
        .B2(keyinput_g59), .ZN(n4648) );
  OAI221_X1 U5153 ( .B1(DATAI_4_), .B2(keyinput_g27), .C1(IR_REG_4__SCAN_IN), 
        .C2(keyinput_g59), .A(n4648), .ZN(n4649) );
  NOR4_X1 U5154 ( .A1(n4652), .A2(n4651), .A3(n4650), .A4(n4649), .ZN(n4653)
         );
  NAND4_X1 U5155 ( .A1(n4656), .A2(n4655), .A3(n4654), .A4(n4653), .ZN(n4758)
         );
  INV_X1 U5156 ( .A(IR_REG_5__SCAN_IN), .ZN(n4752) );
  AOI22_X1 U5157 ( .A1(DATAI_21_), .A2(keyinput_f10), .B1(DATAI_22_), .B2(
        keyinput_f9), .ZN(n4657) );
  OAI221_X1 U5158 ( .B1(DATAI_21_), .B2(keyinput_f10), .C1(DATAI_22_), .C2(
        keyinput_f9), .A(n4657), .ZN(n4664) );
  AOI22_X1 U5159 ( .A1(DATAI_25_), .A2(keyinput_f6), .B1(DATAI_27_), .B2(
        keyinput_f4), .ZN(n4658) );
  OAI221_X1 U5160 ( .B1(DATAI_25_), .B2(keyinput_f6), .C1(DATAI_27_), .C2(
        keyinput_f4), .A(n4658), .ZN(n4663) );
  AOI22_X1 U5161 ( .A1(DATAI_16_), .A2(keyinput_f15), .B1(REG3_REG_13__SCAN_IN), .B2(keyinput_f54), .ZN(n4659) );
  OAI221_X1 U5162 ( .B1(DATAI_16_), .B2(keyinput_f15), .C1(
        REG3_REG_13__SCAN_IN), .C2(keyinput_f54), .A(n4659), .ZN(n4662) );
  AOI22_X1 U5163 ( .A1(REG3_REG_1__SCAN_IN), .A2(keyinput_f42), .B1(
        IR_REG_0__SCAN_IN), .B2(keyinput_f55), .ZN(n4660) );
  OAI221_X1 U5164 ( .B1(REG3_REG_1__SCAN_IN), .B2(keyinput_f42), .C1(
        IR_REG_0__SCAN_IN), .C2(keyinput_f55), .A(n4660), .ZN(n4661) );
  NOR4_X1 U5165 ( .A1(n4664), .A2(n4663), .A3(n4662), .A4(n4661), .ZN(n4716)
         );
  XNOR2_X1 U5166 ( .A(DATAI_3_), .B(keyinput_f28), .ZN(n4668) );
  XNOR2_X1 U5167 ( .A(IR_REG_1__SCAN_IN), .B(keyinput_f56), .ZN(n4667) );
  XNOR2_X1 U5168 ( .A(REG3_REG_17__SCAN_IN), .B(keyinput_f48), .ZN(n4666) );
  XNOR2_X1 U5169 ( .A(IR_REG_6__SCAN_IN), .B(keyinput_f61), .ZN(n4665) );
  NAND4_X1 U5170 ( .A1(n4668), .A2(n4667), .A3(n4666), .A4(n4665), .ZN(n4674)
         );
  XNOR2_X1 U5171 ( .A(keyinput_f19), .B(DATAI_12_), .ZN(n4672) );
  XNOR2_X1 U5172 ( .A(IR_REG_3__SCAN_IN), .B(keyinput_f58), .ZN(n4671) );
  XNOR2_X1 U5173 ( .A(keyinput_f5), .B(DATAI_26_), .ZN(n4670) );
  XNOR2_X1 U5174 ( .A(keyinput_f25), .B(DATAI_6_), .ZN(n4669) );
  NAND4_X1 U5175 ( .A1(n4672), .A2(n4671), .A3(n4670), .A4(n4669), .ZN(n4673)
         );
  NOR2_X1 U5176 ( .A1(n4674), .A2(n4673), .ZN(n4715) );
  AOI22_X1 U5177 ( .A1(n4677), .A2(keyinput_f51), .B1(keyinput_f16), .B2(n4676), .ZN(n4675) );
  OAI221_X1 U5178 ( .B1(n4677), .B2(keyinput_f51), .C1(n4676), .C2(
        keyinput_f16), .A(n4675), .ZN(n4682) );
  AOI22_X1 U5179 ( .A1(REG3_REG_16__SCAN_IN), .A2(keyinput_f46), .B1(
        REG3_REG_19__SCAN_IN), .B2(keyinput_f39), .ZN(n4678) );
  OAI221_X1 U5180 ( .B1(REG3_REG_16__SCAN_IN), .B2(keyinput_f46), .C1(
        REG3_REG_19__SCAN_IN), .C2(keyinput_f39), .A(n4678), .ZN(n4681) );
  AOI22_X1 U5181 ( .A1(DATAI_29_), .A2(keyinput_f2), .B1(REG3_REG_8__SCAN_IN), 
        .B2(keyinput_f41), .ZN(n4679) );
  OAI221_X1 U5182 ( .B1(DATAI_29_), .B2(keyinput_f2), .C1(REG3_REG_8__SCAN_IN), 
        .C2(keyinput_f41), .A(n4679), .ZN(n4680) );
  NOR3_X1 U5183 ( .A1(n4682), .A2(n4681), .A3(n4680), .ZN(n4714) );
  AOI22_X1 U5184 ( .A1(n2638), .A2(keyinput_f3), .B1(keyinput_f8), .B2(n4684), 
        .ZN(n4683) );
  OAI221_X1 U5185 ( .B1(n2638), .B2(keyinput_f3), .C1(n4684), .C2(keyinput_f8), 
        .A(n4683), .ZN(n4688) );
  INV_X1 U5186 ( .A(DATAI_19_), .ZN(n4686) );
  AOI22_X1 U5187 ( .A1(n4686), .A2(keyinput_f12), .B1(U3149), .B2(keyinput_f32), .ZN(n4685) );
  OAI221_X1 U5188 ( .B1(n4686), .B2(keyinput_f12), .C1(U3149), .C2(
        keyinput_f32), .A(n4685), .ZN(n4687) );
  NOR2_X1 U5189 ( .A1(n4688), .A2(n4687), .ZN(n4712) );
  AOI22_X1 U5190 ( .A1(n4691), .A2(keyinput_f36), .B1(keyinput_f53), .B2(n4690), .ZN(n4689) );
  OAI221_X1 U5191 ( .B1(n4691), .B2(keyinput_f36), .C1(n4690), .C2(
        keyinput_f53), .A(n4689), .ZN(n4696) );
  AOI22_X1 U5192 ( .A1(n4694), .A2(keyinput_f35), .B1(keyinput_f26), .B2(n4693), .ZN(n4692) );
  OAI221_X1 U5193 ( .B1(n4694), .B2(keyinput_f35), .C1(n4693), .C2(
        keyinput_f26), .A(n4692), .ZN(n4695) );
  NOR2_X1 U5194 ( .A1(n4696), .A2(n4695), .ZN(n4711) );
  XNOR2_X1 U5195 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput_f38), .ZN(n4700) );
  XNOR2_X1 U5196 ( .A(DATAI_9_), .B(keyinput_f22), .ZN(n4699) );
  XNOR2_X1 U5197 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_f50), .ZN(n4698) );
  XNOR2_X1 U5198 ( .A(DATAI_0_), .B(keyinput_f31), .ZN(n4697) );
  NAND4_X1 U5199 ( .A1(n4700), .A2(n4699), .A3(n4698), .A4(n4697), .ZN(n4706)
         );
  XNOR2_X1 U5200 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_f52), .ZN(n4704) );
  XNOR2_X1 U5201 ( .A(REG3_REG_10__SCAN_IN), .B(keyinput_f37), .ZN(n4703) );
  XNOR2_X1 U5202 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_f59), .ZN(n4702) );
  XNOR2_X1 U5203 ( .A(REG3_REG_7__SCAN_IN), .B(keyinput_f33), .ZN(n4701) );
  NAND4_X1 U5204 ( .A1(n4704), .A2(n4703), .A3(n4702), .A4(n4701), .ZN(n4705)
         );
  NOR2_X1 U5205 ( .A1(n4706), .A2(n4705), .ZN(n4710) );
  AOI22_X1 U5206 ( .A1(n2475), .A2(keyinput_f23), .B1(n3704), .B2(keyinput_f43), .ZN(n4707) );
  OAI221_X1 U5207 ( .B1(n2475), .B2(keyinput_f23), .C1(n3704), .C2(
        keyinput_f43), .A(n4707), .ZN(n4708) );
  INV_X1 U5208 ( .A(n4708), .ZN(n4709) );
  AND4_X1 U5209 ( .A1(n4712), .A2(n4711), .A3(n4710), .A4(n4709), .ZN(n4713)
         );
  AND4_X1 U5210 ( .A1(n4716), .A2(n4715), .A3(n4714), .A4(n4713), .ZN(n4750)
         );
  AOI22_X1 U5211 ( .A1(n4718), .A2(keyinput_f1), .B1(n2595), .B2(keyinput_f13), 
        .ZN(n4717) );
  OAI221_X1 U5212 ( .B1(n4718), .B2(keyinput_f1), .C1(n2595), .C2(keyinput_f13), .A(n4717), .ZN(n4731) );
  INV_X1 U5213 ( .A(DATAI_4_), .ZN(n4721) );
  AOI22_X1 U5214 ( .A1(n4721), .A2(keyinput_f27), .B1(n4720), .B2(keyinput_f34), .ZN(n4719) );
  OAI221_X1 U5215 ( .B1(n4721), .B2(keyinput_f27), .C1(n4720), .C2(
        keyinput_f34), .A(n4719), .ZN(n4730) );
  AOI22_X1 U5216 ( .A1(n4724), .A2(keyinput_f44), .B1(keyinput_f14), .B2(n4723), .ZN(n4722) );
  OAI221_X1 U5217 ( .B1(n4724), .B2(keyinput_f44), .C1(n4723), .C2(
        keyinput_f14), .A(n4722), .ZN(n4729) );
  INV_X1 U5218 ( .A(DATAI_7_), .ZN(n4727) );
  AOI22_X1 U5219 ( .A1(n4727), .A2(keyinput_f24), .B1(n4726), .B2(keyinput_f45), .ZN(n4725) );
  OAI221_X1 U5220 ( .B1(n4727), .B2(keyinput_f24), .C1(n4726), .C2(
        keyinput_f45), .A(n4725), .ZN(n4728) );
  NOR4_X1 U5221 ( .A1(n4731), .A2(n4730), .A3(n4729), .A4(n4728), .ZN(n4749)
         );
  AOI22_X1 U5222 ( .A1(DATAI_13_), .A2(keyinput_f18), .B1(IR_REG_7__SCAN_IN), 
        .B2(keyinput_f62), .ZN(n4732) );
  OAI221_X1 U5223 ( .B1(DATAI_13_), .B2(keyinput_f18), .C1(IR_REG_7__SCAN_IN), 
        .C2(keyinput_f62), .A(n4732), .ZN(n4739) );
  AOI22_X1 U5224 ( .A1(DATAI_10_), .A2(keyinput_f21), .B1(DATAI_14_), .B2(
        keyinput_f17), .ZN(n4733) );
  OAI221_X1 U5225 ( .B1(DATAI_10_), .B2(keyinput_f21), .C1(DATAI_14_), .C2(
        keyinput_f17), .A(n4733), .ZN(n4738) );
  AOI22_X1 U5226 ( .A1(DATAI_11_), .A2(keyinput_f20), .B1(IR_REG_8__SCAN_IN), 
        .B2(keyinput_f63), .ZN(n4734) );
  OAI221_X1 U5227 ( .B1(DATAI_11_), .B2(keyinput_f20), .C1(IR_REG_8__SCAN_IN), 
        .C2(keyinput_f63), .A(n4734), .ZN(n4737) );
  AOI22_X1 U5228 ( .A1(REG3_REG_5__SCAN_IN), .A2(keyinput_f47), .B1(
        IR_REG_2__SCAN_IN), .B2(keyinput_f57), .ZN(n4735) );
  OAI221_X1 U5229 ( .B1(REG3_REG_5__SCAN_IN), .B2(keyinput_f47), .C1(
        IR_REG_2__SCAN_IN), .C2(keyinput_f57), .A(n4735), .ZN(n4736) );
  NOR4_X1 U5230 ( .A1(n4739), .A2(n4738), .A3(n4737), .A4(n4736), .ZN(n4748)
         );
  XNOR2_X1 U5231 ( .A(DATAI_1_), .B(keyinput_f30), .ZN(n4746) );
  AOI22_X1 U5232 ( .A1(DATAI_2_), .A2(keyinput_f29), .B1(n2610), .B2(
        keyinput_f11), .ZN(n4740) );
  OAI221_X1 U5233 ( .B1(DATAI_2_), .B2(keyinput_f29), .C1(n2610), .C2(
        keyinput_f11), .A(n4740), .ZN(n4745) );
  AOI22_X1 U5234 ( .A1(DATAI_31_), .A2(keyinput_f0), .B1(REG3_REG_24__SCAN_IN), 
        .B2(keyinput_f49), .ZN(n4741) );
  OAI221_X1 U5235 ( .B1(DATAI_31_), .B2(keyinput_f0), .C1(REG3_REG_24__SCAN_IN), .C2(keyinput_f49), .A(n4741), .ZN(n4744) );
  AOI22_X1 U5236 ( .A1(DATAI_24_), .A2(keyinput_f7), .B1(REG3_REG_28__SCAN_IN), 
        .B2(keyinput_f40), .ZN(n4742) );
  OAI221_X1 U5237 ( .B1(DATAI_24_), .B2(keyinput_f7), .C1(REG3_REG_28__SCAN_IN), .C2(keyinput_f40), .A(n4742), .ZN(n4743) );
  NOR4_X1 U5238 ( .A1(n4746), .A2(n4745), .A3(n4744), .A4(n4743), .ZN(n4747)
         );
  NAND4_X1 U5239 ( .A1(n4750), .A2(n4749), .A3(n4748), .A4(n4747), .ZN(n4751)
         );
  OAI21_X1 U5240 ( .B1(keyinput_f60), .B2(n4752), .A(n4751), .ZN(n4754) );
  OAI211_X1 U5241 ( .C1(n4754), .C2(keyinput_f60), .A(keyinput_g60), .B(n4752), 
        .ZN(n4756) );
  INV_X1 U5242 ( .A(keyinput_g60), .ZN(n4753) );
  NAND3_X1 U5243 ( .A1(n4754), .A2(IR_REG_5__SCAN_IN), .A3(n4753), .ZN(n4755)
         );
  NAND2_X1 U5244 ( .A1(n4756), .A2(n4755), .ZN(n4757) );
  OAI21_X1 U5245 ( .B1(n4759), .B2(n4758), .A(n4757), .ZN(n4760) );
  XOR2_X1 U5246 ( .A(n4761), .B(n4760), .Z(U3352) );
  CLKBUF_X1 U2298 ( .A(n4392), .Z(n2049) );
endmodule

