

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593;

  NOR4_X1 U4898 ( .A1(n8329), .A2(n8411), .A3(n8328), .A4(n8327), .ZN(n8330)
         );
  NAND2_X1 U4899 ( .A1(n7174), .A2(n7173), .ZN(n9590) );
  CLKBUF_X1 U4900 ( .A(n5640), .Z(n6182) );
  AND3_X1 U4901 ( .A1(n6383), .A2(n6385), .A3(n6384), .ZN(n10447) );
  AND4_X1 U4902 ( .A1(n4441), .A2(n5548), .A3(n5547), .A4(n5546), .ZN(n7108)
         );
  CLKBUF_X2 U4903 ( .A(n6468), .Z(n9570) );
  CLKBUF_X2 U4904 ( .A(n5545), .Z(n5900) );
  INV_X1 U4905 ( .A(n6468), .ZN(n6788) );
  INV_X2 U4906 ( .A(n5641), .ZN(n7743) );
  NAND2_X2 U4907 ( .A1(n6282), .A2(n6279), .ZN(n6593) );
  BUF_X1 U4908 ( .A(n6281), .Z(n7720) );
  XNOR2_X1 U4909 ( .A(n6278), .B(n6277), .ZN(n6281) );
  INV_X2 U4910 ( .A(n4393), .ZN(n4394) );
  NOR4_X1 U4911 ( .A1(n8875), .A2(n8882), .A3(n8907), .A4(n8331), .ZN(n8332)
         );
  INV_X1 U4912 ( .A(n8494), .ZN(n8481) );
  INV_X2 U4913 ( .A(n5167), .ZN(n4396) );
  INV_X1 U4914 ( .A(n7291), .ZN(n7543) );
  OR2_X1 U4915 ( .A1(n8978), .A2(n8710), .ZN(n8479) );
  NAND2_X1 U4916 ( .A1(n5416), .A2(n5415), .ZN(n5697) );
  INV_X1 U4917 ( .A(n6861), .ZN(n6173) );
  NAND2_X1 U4918 ( .A1(n6861), .A2(n5167), .ZN(n5560) );
  NAND2_X2 U4919 ( .A1(n8687), .A2(n6034), .ZN(n6861) );
  AND2_X1 U4920 ( .A1(n5247), .A2(n5619), .ZN(n7291) );
  NAND2_X1 U4921 ( .A1(n5357), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5358) );
  INV_X1 U4922 ( .A(n6281), .ZN(n6279) );
  NAND2_X1 U4923 ( .A1(n7720), .A2(n6282), .ZN(n6468) );
  NAND2_X1 U4924 ( .A1(n7220), .A2(n9739), .ZN(n7239) );
  AND3_X1 U4925 ( .A1(n5587), .A2(n5586), .A3(n5585), .ZN(n7258) );
  INV_X1 U4926 ( .A(n8453), .ZN(n8841) );
  INV_X1 U4927 ( .A(n8850), .ZN(n8513) );
  INV_X1 U4928 ( .A(n10170), .ZN(n10118) );
  AND2_X2 U4929 ( .A1(n4521), .A2(n4520), .ZN(n5167) );
  OR2_X1 U4930 ( .A1(n6654), .A2(n6705), .ZN(n6697) );
  NAND4_X2 U4931 ( .A1(n6287), .A2(n6286), .A3(n6285), .A4(n6284), .ZN(n6654)
         );
  AND2_X1 U4932 ( .A1(n4521), .A2(n4520), .ZN(n4393) );
  INV_X2 U4933 ( .A(n4393), .ZN(n4395) );
  INV_X2 U4934 ( .A(n5167), .ZN(n4397) );
  BUF_X1 U4935 ( .A(n9008), .Z(n4398) );
  XNOR2_X2 U4936 ( .A(n5358), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5359) );
  XNOR2_X2 U4937 ( .A(n4766), .B(n5493), .ZN(n6034) );
  NAND2_X1 U4938 ( .A1(n7727), .A2(n7726), .ZN(n8978) );
  NAND2_X1 U4939 ( .A1(n4523), .A2(n9577), .ZN(n10004) );
  OR2_X1 U4940 ( .A1(n7475), .A2(n4905), .ZN(n4988) );
  NAND2_X1 U4941 ( .A1(n4779), .A2(n4778), .ZN(n5322) );
  AND2_X1 U4942 ( .A1(n9606), .A2(n9739), .ZN(n9603) );
  INV_X2 U4943 ( .A(n6504), .ZN(n8096) );
  NAND2_X1 U4944 ( .A1(n4527), .A2(n5177), .ZN(n5616) );
  NAND2_X1 U4945 ( .A1(n6663), .A2(n10447), .ZN(n9799) );
  INV_X2 U4946 ( .A(n8123), .ZN(n8084) );
  INV_X4 U4947 ( .A(n8127), .ZN(n8133) );
  CLKBUF_X1 U4948 ( .A(n6105), .Z(n10530) );
  INV_X1 U4949 ( .A(n7104), .ZN(n10518) );
  OR2_X2 U4950 ( .A1(n6329), .A2(n9829), .ZN(n10458) );
  INV_X2 U4951 ( .A(n5941), .ZN(n8308) );
  CLKBUF_X2 U4952 ( .A(n5526), .Z(n5641) );
  INV_X1 U4953 ( .A(n9680), .ZN(n7859) );
  OR2_X1 U4954 ( .A1(n9690), .A2(n9829), .ZN(n6696) );
  INV_X1 U4955 ( .A(n9829), .ZN(n7007) );
  NAND2_X2 U4956 ( .A1(n6197), .A2(n6533), .ZN(n6380) );
  MUX2_X1 U4957 ( .A(n8496), .B(n8495), .S(n8494), .Z(n8499) );
  NAND2_X1 U4958 ( .A1(n4731), .A2(n4729), .ZN(n8259) );
  NAND2_X1 U4959 ( .A1(n5016), .A2(n8484), .ZN(n8490) );
  NAND2_X1 U4960 ( .A1(n10217), .A2(n4415), .ZN(n10323) );
  OR2_X1 U4961 ( .A1(n4935), .A2(n9079), .ZN(n4931) );
  AOI21_X1 U4962 ( .B1(n8982), .B2(n9079), .A(n10537), .ZN(n4933) );
  NOR2_X1 U4963 ( .A1(n7774), .A2(n8476), .ZN(n8976) );
  AND2_X1 U4964 ( .A1(n8981), .A2(n8980), .ZN(n8982) );
  NOR2_X1 U4965 ( .A1(n5928), .A2(n8220), .ZN(n5929) );
  AOI21_X1 U4966 ( .B1(n4820), .B2(n10192), .A(n4817), .ZN(n10234) );
  AND2_X1 U4967 ( .A1(n4794), .A2(n4793), .ZN(n8220) );
  NAND2_X1 U4968 ( .A1(n5094), .A2(n5092), .ZN(n4794) );
  NAND2_X1 U4969 ( .A1(n4918), .A2(n4917), .ZN(n8120) );
  OAI21_X1 U4970 ( .B1(n10225), .B2(n10299), .A(n4799), .ZN(n4798) );
  NAND2_X1 U4971 ( .A1(n7994), .A2(n9820), .ZN(n9968) );
  AOI21_X1 U4972 ( .B1(n9426), .B2(n8069), .A(n8068), .ZN(n9496) );
  NAND2_X1 U4973 ( .A1(n8172), .A2(n5867), .ZN(n8233) );
  NAND2_X1 U4974 ( .A1(n9413), .A2(n8091), .ZN(n9488) );
  NAND2_X1 U4975 ( .A1(n5091), .A2(n5090), .ZN(n8172) );
  NAND2_X1 U4976 ( .A1(n8310), .A2(n8309), .ZN(n8963) );
  AND2_X1 U4977 ( .A1(n8476), .A2(n8475), .ZN(n5020) );
  INV_X1 U4978 ( .A(n8975), .ZN(n5018) );
  NAND2_X1 U4979 ( .A1(n4982), .A2(n8053), .ZN(n4981) );
  NAND2_X1 U4980 ( .A1(n5813), .A2(n5812), .ZN(n8204) );
  NAND2_X1 U4981 ( .A1(n4936), .A2(n4939), .ZN(n8840) );
  XNOR2_X1 U4982 ( .A(n8984), .B(n8742), .ZN(n8717) );
  AND2_X1 U4983 ( .A1(n6038), .A2(n7742), .ZN(n7777) );
  NAND2_X1 U4984 ( .A1(n4847), .A2(n4846), .ZN(n10046) );
  AND2_X1 U4985 ( .A1(n5367), .A2(n5366), .ZN(n8192) );
  NAND2_X1 U4986 ( .A1(n9407), .A2(n8036), .ZN(n8047) );
  NAND2_X1 U4987 ( .A1(n7515), .A2(n7516), .ZN(n4724) );
  NAND2_X1 U4988 ( .A1(n5962), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6037) );
  AND2_X1 U4989 ( .A1(n5903), .A2(n5902), .ZN(n8453) );
  NAND2_X1 U4990 ( .A1(n4767), .A2(n5033), .ZN(n4926) );
  NAND2_X1 U4991 ( .A1(n4838), .A2(n4836), .ZN(n10307) );
  NAND2_X1 U4992 ( .A1(n5498), .A2(n5497), .ZN(n9000) );
  NAND2_X1 U4993 ( .A1(n5882), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5919) );
  NAND2_X1 U4994 ( .A1(n7178), .A2(n7177), .ZN(n7457) );
  OAI21_X1 U4995 ( .B1(n5954), .B2(n5953), .A(n5955), .ZN(n5976) );
  NAND2_X1 U4996 ( .A1(n5146), .A2(n5145), .ZN(n7584) );
  NAND2_X1 U4997 ( .A1(n7556), .A2(n8391), .ZN(n5146) );
  NAND2_X1 U4998 ( .A1(n5492), .A2(n5491), .ZN(n5936) );
  NAND2_X1 U4999 ( .A1(n7843), .A2(n7842), .ZN(n10275) );
  NAND2_X1 U5000 ( .A1(n4644), .A2(n7833), .ZN(n10282) );
  NAND2_X1 U5001 ( .A1(n5823), .A2(n5822), .ZN(n9037) );
  NAND2_X1 U5002 ( .A1(n5799), .A2(n5798), .ZN(n8942) );
  NAND2_X1 U5003 ( .A1(n4844), .A2(n4418), .ZN(n4843) );
  NAND2_X1 U5004 ( .A1(n5339), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5840) );
  NAND2_X1 U5005 ( .A1(n4607), .A2(n5739), .ZN(n8407) );
  INV_X1 U5006 ( .A(n5824), .ZN(n5339) );
  NAND2_X1 U5007 ( .A1(n5760), .A2(n5759), .ZN(n9054) );
  NAND2_X1 U5008 ( .A1(n5721), .A2(n5720), .ZN(n9067) );
  NAND2_X1 U5009 ( .A1(n7388), .A2(n7387), .ZN(n10303) );
  NAND2_X1 U5010 ( .A1(n7033), .A2(n8356), .ZN(n4509) );
  INV_X1 U5011 ( .A(n9610), .ZN(n4399) );
  NAND2_X1 U5012 ( .A1(n8376), .A2(n8372), .ZN(n8320) );
  NAND2_X1 U5013 ( .A1(n4710), .A2(n4709), .ZN(n9739) );
  NAND2_X1 U5014 ( .A1(n7098), .A2(n8363), .ZN(n7033) );
  NAND2_X1 U5015 ( .A1(n4825), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5804) );
  XNOR2_X1 U5016 ( .A(n4770), .B(n5716), .ZN(n7385) );
  NAND2_X1 U5017 ( .A1(n5639), .A2(n5638), .ZN(n7483) );
  XNOR2_X1 U5018 ( .A(n5673), .B(n5319), .ZN(n9389) );
  INV_X1 U5019 ( .A(n7272), .ZN(n10529) );
  INV_X1 U5020 ( .A(n5781), .ZN(n4825) );
  NAND2_X2 U5021 ( .A1(n8352), .A2(n8363), .ZN(n7030) );
  NAND2_X1 U5022 ( .A1(n5616), .A2(n5414), .ZN(n5635) );
  INV_X1 U5023 ( .A(n7126), .ZN(n5060) );
  INV_X1 U5024 ( .A(n9848), .ZN(n7242) );
  NAND2_X1 U5025 ( .A1(n4822), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5762) );
  BUF_X2 U5026 ( .A(n7728), .Z(n4796) );
  XNOR2_X1 U5027 ( .A(n5616), .B(n5615), .ZN(n4780) );
  NAND2_X1 U5028 ( .A1(n5329), .A2(n6474), .ZN(n6659) );
  NAND4_X2 U5029 ( .A1(n6597), .A2(n6596), .A3(n6595), .A4(n6594), .ZN(n9851)
         );
  INV_X1 U5030 ( .A(n5741), .ZN(n4822) );
  INV_X2 U5031 ( .A(n5575), .ZN(n7728) );
  AND2_X2 U5032 ( .A1(n6199), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  NAND4_X1 U5033 ( .A1(n5595), .A2(n5594), .A3(n5593), .A4(n5592), .ZN(n8526)
         );
  NAND2_X1 U5034 ( .A1(n4435), .A2(n5271), .ZN(n9853) );
  INV_X1 U5035 ( .A(n5512), .ZN(n7729) );
  NAND2_X1 U5036 ( .A1(n4823), .A2(n4464), .ZN(n5741) );
  NAND2_X1 U5037 ( .A1(n4593), .A2(n5408), .ZN(n5581) );
  INV_X1 U5038 ( .A(n5725), .ZN(n4823) );
  AND4_X1 U5039 ( .A1(n5521), .A2(n5520), .A3(n5519), .A4(n5518), .ZN(n6617)
         );
  NAND2_X1 U5040 ( .A1(n6025), .A2(n6490), .ZN(n6105) );
  AND3_X1 U5041 ( .A1(n5553), .A2(n5552), .A3(n4448), .ZN(n6094) );
  CLKBUF_X1 U5042 ( .A(n5896), .Z(n5965) );
  AND3_X1 U5043 ( .A1(n6499), .A2(n6498), .A3(n6497), .ZN(n6660) );
  NAND3_X1 U5044 ( .A1(n6452), .A2(n6451), .A3(n6450), .ZN(n6945) );
  NAND2_X1 U5045 ( .A1(n4828), .A2(n5404), .ZN(n5559) );
  NOR2_X1 U5046 ( .A1(n5155), .A2(n5716), .ZN(n5154) );
  NAND2_X1 U5047 ( .A1(n5385), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5380) );
  BUF_X1 U5048 ( .A(n6280), .Z(n4749) );
  XNOR2_X1 U5049 ( .A(n6069), .B(n6068), .ZN(n7721) );
  NAND2_X1 U5050 ( .A1(n6861), .A2(n4395), .ZN(n5941) );
  INV_X1 U5051 ( .A(n6280), .ZN(n6282) );
  AND2_X1 U5052 ( .A1(n5360), .A2(n5361), .ZN(n5640) );
  NAND2_X2 U5053 ( .A1(n6380), .A2(n5167), .ZN(n9680) );
  XNOR2_X1 U5054 ( .A(n5383), .B(n5382), .ZN(n8337) );
  XNOR2_X1 U5055 ( .A(n6276), .B(n6275), .ZN(n6280) );
  NAND2_X1 U5056 ( .A1(n6055), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6057) );
  NAND2_X1 U5057 ( .A1(n4879), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6278) );
  XNOR2_X1 U5058 ( .A(n4904), .B(P1_IR_REG_20__SCAN_IN), .ZN(n9829) );
  XNOR2_X1 U5059 ( .A(n4694), .B(n6078), .ZN(n6533) );
  NAND2_X1 U5060 ( .A1(n5210), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6071) );
  NAND2_X1 U5061 ( .A1(n5335), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5643) );
  INV_X1 U5062 ( .A(n5621), .ZN(n5335) );
  NAND2_X1 U5063 ( .A1(n5353), .A2(n5258), .ZN(n5257) );
  NAND4_X1 U5064 ( .A1(n5347), .A2(n5345), .A3(n5346), .A4(n5368), .ZN(n5348)
         );
  NAND2_X1 U5065 ( .A1(n9137), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5606) );
  INV_X1 U5066 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n6160) );
  NOR2_X1 U5067 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n4867) );
  NOR2_X1 U5068 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n6065) );
  NOR2_X1 U5069 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n6053) );
  NOR2_X1 U5070 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n6052) );
  NOR2_X1 U5071 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n6051) );
  NOR2_X1 U5072 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5790) );
  NOR2_X1 U5073 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5345) );
  NOR2_X1 U5074 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5346) );
  INV_X1 U5075 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5379) );
  NOR2_X1 U5076 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5351) );
  NOR2_X1 U5077 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5350) );
  NOR2_X1 U5078 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n5349) );
  INV_X1 U5079 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5701) );
  INV_X1 U5080 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4592) );
  NAND2_X2 U5081 ( .A1(n8884), .A2(n8431), .ZN(n8863) );
  NOR2_X2 U5082 ( .A1(n5322), .A2(n4775), .ZN(n4582) );
  XNOR2_X1 U5083 ( .A(n5559), .B(n5558), .ZN(n6580) );
  NAND2_X2 U5084 ( .A1(n4806), .A2(n8915), .ZN(n5575) );
  NAND2_X1 U5085 ( .A1(n8286), .A2(n8285), .ZN(n8971) );
  NAND2_X1 U5086 ( .A1(n4604), .A2(n4404), .ZN(n8284) );
  AND2_X1 U5087 ( .A1(n8485), .A2(n8312), .ZN(n8489) );
  NAND2_X1 U5088 ( .A1(n5132), .A2(n5131), .ZN(n8881) );
  NOR2_X1 U5089 ( .A1(n7782), .A2(n8907), .ZN(n5131) );
  OR2_X1 U5090 ( .A1(n9049), .A2(n8925), .ZN(n7780) );
  INV_X1 U5091 ( .A(n6696), .ZN(n5179) );
  INV_X1 U5092 ( .A(n4852), .ZN(n4851) );
  NAND2_X1 U5093 ( .A1(n6380), .A2(n4396), .ZN(n6744) );
  NAND2_X1 U5094 ( .A1(n5439), .A2(n5438), .ZN(n5442) );
  INV_X1 U5095 ( .A(SI_12_), .ZN(n5438) );
  AND2_X1 U5096 ( .A1(n4455), .A2(n5093), .ZN(n5092) );
  NAND2_X1 U5097 ( .A1(n8233), .A2(n5097), .ZN(n5094) );
  INV_X1 U5098 ( .A(n5917), .ZN(n5093) );
  AND2_X1 U5099 ( .A1(n8701), .A2(n8702), .ZN(n8972) );
  AND2_X1 U5100 ( .A1(n8483), .A2(n8482), .ZN(n8975) );
  NAND2_X1 U5101 ( .A1(n4692), .A2(n4691), .ZN(n8832) );
  AOI21_X1 U5102 ( .B1(n4402), .B2(n5225), .A(n4465), .ZN(n4691) );
  NAND2_X1 U5103 ( .A1(n8900), .A2(n4402), .ZN(n4692) );
  INV_X1 U5104 ( .A(n4859), .ZN(n4858) );
  OAI21_X1 U5105 ( .B1(n9820), .B2(n4860), .A(n7961), .ZN(n4859) );
  NAND2_X1 U5106 ( .A1(n4862), .A2(n7951), .ZN(n4860) );
  INV_X1 U5107 ( .A(n6073), .ZN(n6075) );
  NAND2_X1 U5108 ( .A1(n4897), .A2(n4895), .ZN(n9617) );
  NAND2_X1 U5109 ( .A1(n4658), .A2(n4656), .ZN(n8465) );
  OR2_X1 U5110 ( .A1(n8435), .A2(n4657), .ZN(n4656) );
  AND2_X1 U5111 ( .A1(n4659), .A2(n4426), .ZN(n4658) );
  NAND2_X1 U5112 ( .A1(n4742), .A2(n6102), .ZN(n5512) );
  NAND2_X1 U5113 ( .A1(n4469), .A2(n4741), .ZN(n4742) );
  AND3_X1 U5114 ( .A1(n8340), .A2(n8350), .A3(n8339), .ZN(n8494) );
  NOR2_X1 U5115 ( .A1(n5840), .A2(n5839), .ZN(n4826) );
  NAND2_X1 U5116 ( .A1(n7291), .A2(n8524), .ZN(n8380) );
  AND2_X1 U5117 ( .A1(n10209), .A2(n4889), .ZN(n4888) );
  OR2_X1 U5118 ( .A1(n10208), .A2(n9688), .ZN(n4889) );
  AOI21_X1 U5119 ( .B1(n5157), .B2(n10208), .A(n10209), .ZN(n4886) );
  NAND2_X1 U5120 ( .A1(n5918), .A2(n5917), .ZN(n8162) );
  NAND2_X1 U5121 ( .A1(n4733), .A2(n4736), .ZN(n5918) );
  AND2_X1 U5122 ( .A1(n4455), .A2(n4737), .ZN(n4736) );
  INV_X1 U5123 ( .A(n6105), .ZN(n4806) );
  AND3_X1 U5124 ( .A1(n8489), .A2(n4975), .A3(n4974), .ZN(n8336) );
  INV_X1 U5125 ( .A(n8486), .ZN(n4975) );
  INV_X1 U5126 ( .A(n5963), .ZN(n5962) );
  OR2_X1 U5127 ( .A1(n8746), .A2(n8193), .ZN(n8470) );
  AND2_X1 U5128 ( .A1(n4517), .A2(n4515), .ZN(n5144) );
  NAND2_X1 U5129 ( .A1(n4586), .A2(n8467), .ZN(n4517) );
  OR2_X1 U5130 ( .A1(n9000), .A2(n8192), .ZN(n8466) );
  OR2_X1 U5131 ( .A1(n9005), .A2(n8824), .ZN(n8459) );
  AND2_X1 U5132 ( .A1(n8794), .A2(n8444), .ZN(n8792) );
  NAND2_X1 U5133 ( .A1(n4826), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5881) );
  AND2_X1 U5134 ( .A1(n7780), .A2(n7695), .ZN(n8420) );
  XNOR2_X1 U5135 ( .A(n8407), .B(n8156), .ZN(n7680) );
  NAND2_X1 U5136 ( .A1(n6025), .A2(n8350), .ZN(n6102) );
  NAND2_X1 U5137 ( .A1(n8975), .A2(n5240), .ZN(n5239) );
  NOR2_X1 U5138 ( .A1(n8973), .A2(n9079), .ZN(n5240) );
  NAND2_X1 U5139 ( .A1(n8881), .A2(n7785), .ZN(n8884) );
  NOR2_X1 U5140 ( .A1(n5257), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n5256) );
  NAND2_X1 U5141 ( .A1(n7457), .A2(n7179), .ZN(n7475) );
  NAND2_X1 U5142 ( .A1(n5198), .A2(n5197), .ZN(n5196) );
  OR2_X1 U5143 ( .A1(n8074), .A2(n8073), .ZN(n5197) );
  OR2_X1 U5144 ( .A1(n9497), .A2(n5200), .ZN(n5198) );
  NAND2_X1 U5145 ( .A1(n8082), .A2(n8081), .ZN(n9413) );
  OAI21_X1 U5146 ( .B1(n4981), .B2(n4408), .A(n4910), .ZN(n8082) );
  OR2_X1 U5147 ( .A1(n6401), .A2(n6628), .ZN(n6407) );
  OR2_X1 U5148 ( .A1(n9943), .A2(n9966), .ZN(n9724) );
  NAND2_X1 U5149 ( .A1(n9876), .A2(n9875), .ZN(n6425) );
  AND2_X1 U5150 ( .A1(n4446), .A2(n6424), .ZN(n5009) );
  OR2_X1 U5151 ( .A1(n7942), .A2(n7941), .ZN(n7967) );
  AOI21_X1 U5152 ( .B1(n4406), .B2(n4652), .A(n4651), .ZN(n4650) );
  INV_X1 U5153 ( .A(n9996), .ZN(n4651) );
  NAND2_X1 U5154 ( .A1(n10030), .A2(n4406), .ZN(n4649) );
  OR2_X1 U5155 ( .A1(n10238), .A2(n10013), .ZN(n9985) );
  INV_X1 U5156 ( .A(n4850), .ZN(n4849) );
  OAI21_X1 U5157 ( .B1(n4437), .B2(n4851), .A(n7879), .ZN(n4850) );
  OR2_X1 U5158 ( .A1(n10270), .A2(n9482), .ZN(n9643) );
  NOR2_X1 U5159 ( .A1(n10139), .A2(n4643), .ZN(n4642) );
  INV_X1 U5160 ( .A(n7833), .ZN(n4643) );
  NOR2_X1 U5161 ( .A1(n10292), .A2(n10190), .ZN(n5293) );
  OR2_X1 U5162 ( .A1(n10292), .A2(n10138), .ZN(n9633) );
  NAND2_X1 U5163 ( .A1(n4702), .A2(n4701), .ZN(n9611) );
  AOI21_X1 U5164 ( .B1(n9733), .B2(n4699), .A(n4399), .ZN(n4698) );
  INV_X1 U5165 ( .A(n9607), .ZN(n4699) );
  OR2_X1 U5166 ( .A1(n9852), .A2(n10457), .ZN(n9807) );
  AND2_X1 U5167 ( .A1(n9611), .A2(n9618), .ZN(n9710) );
  NAND2_X1 U5168 ( .A1(n7718), .A2(n7717), .ZN(n8011) );
  NAND2_X1 U5169 ( .A1(n7725), .A2(n7724), .ZN(n7718) );
  NAND2_X1 U5170 ( .A1(n5978), .A2(n5977), .ZN(n7711) );
  NAND2_X1 U5171 ( .A1(n5486), .A2(n5485), .ZN(n5890) );
  NAND2_X1 U5172 ( .A1(n5471), .A2(n9249), .ZN(n5474) );
  NOR2_X1 U5173 ( .A1(n5849), .A2(n5166), .ZN(n5165) );
  INV_X1 U5174 ( .A(n5469), .ZN(n5166) );
  AND2_X1 U5175 ( .A1(n5479), .A2(n5478), .ZN(n5868) );
  AND2_X1 U5176 ( .A1(n5170), .A2(n5466), .ZN(n5169) );
  NAND2_X1 U5177 ( .A1(n4970), .A2(n5451), .ZN(n5775) );
  NAND2_X1 U5178 ( .A1(n5442), .A2(n5441), .ZN(n5716) );
  NAND2_X1 U5179 ( .A1(n4596), .A2(n4594), .ZN(n5436) );
  AOI21_X1 U5180 ( .B1(n5695), .B2(n5692), .A(n4595), .ZN(n4594) );
  NAND2_X1 U5181 ( .A1(n5635), .A2(n4450), .ZN(n4596) );
  NAND2_X1 U5182 ( .A1(n5699), .A2(n5697), .ZN(n4595) );
  AND2_X1 U5183 ( .A1(n5429), .A2(n5634), .ZN(n4672) );
  AOI21_X1 U5184 ( .B1(n5178), .B2(n5412), .A(n4440), .ZN(n5177) );
  NAND2_X1 U5185 ( .A1(n5581), .A2(n4813), .ZN(n4527) );
  INV_X1 U5186 ( .A(n5411), .ZN(n5178) );
  INV_X1 U5187 ( .A(n8164), .ZN(n4793) );
  NOR2_X1 U5188 ( .A1(n8287), .A2(n4759), .ZN(n5138) );
  NAND2_X1 U5189 ( .A1(n5137), .A2(n8482), .ZN(n5136) );
  INV_X1 U5190 ( .A(n5139), .ZN(n5137) );
  INV_X1 U5191 ( .A(n5965), .ZN(n7747) );
  OR3_X1 U5192 ( .A1(n7528), .A2(n9122), .A3(n7653), .ZN(n6815) );
  OR2_X1 U5193 ( .A1(n8559), .A2(n6842), .ZN(n4563) );
  INV_X1 U5194 ( .A(n8638), .ZN(n4559) );
  NAND2_X1 U5195 ( .A1(n8832), .A2(n7766), .ZN(n7768) );
  NAND2_X1 U5196 ( .A1(n7764), .A2(n5228), .ZN(n5227) );
  INV_X1 U5197 ( .A(n7763), .ZN(n5228) );
  NOR2_X1 U5198 ( .A1(n7765), .A2(n5231), .ZN(n5229) );
  INV_X1 U5199 ( .A(n7764), .ZN(n5226) );
  NAND2_X1 U5200 ( .A1(n4582), .A2(n4581), .ZN(n8852) );
  NAND2_X1 U5201 ( .A1(n8900), .A2(n7762), .ZN(n8880) );
  NOR2_X1 U5202 ( .A1(n8328), .A2(n4947), .ZN(n5145) );
  INV_X1 U5203 ( .A(n8389), .ZN(n4947) );
  OAI21_X1 U5204 ( .B1(n8707), .B2(n4439), .A(n8935), .ZN(n8713) );
  AND2_X1 U5205 ( .A1(n5140), .A2(n8479), .ZN(n8706) );
  OAI21_X1 U5206 ( .B1(n8733), .B2(n4683), .A(n4681), .ZN(n7774) );
  NAND2_X1 U5207 ( .A1(n7772), .A2(n7773), .ZN(n4683) );
  OR2_X1 U5208 ( .A1(n4684), .A2(n4682), .ZN(n4681) );
  INV_X1 U5209 ( .A(n7773), .ZN(n4682) );
  INV_X1 U5210 ( .A(n9074), .ZN(n10528) );
  OR2_X1 U5211 ( .A1(n6484), .A2(n6483), .ZN(n6731) );
  NAND2_X1 U5212 ( .A1(n5533), .A2(n5531), .ZN(n5561) );
  NAND2_X1 U5213 ( .A1(n4403), .A2(n4613), .ZN(n4612) );
  AND2_X1 U5214 ( .A1(n5180), .A2(n4615), .ZN(n4614) );
  INV_X1 U5215 ( .A(n4987), .ZN(n4613) );
  NAND2_X1 U5216 ( .A1(n7169), .A2(n7168), .ZN(n7184) );
  INV_X1 U5217 ( .A(n6330), .ZN(n6667) );
  OR2_X1 U5218 ( .A1(n10226), .A2(n8138), .ZN(n9781) );
  NOR2_X1 U5219 ( .A1(n4552), .A2(n4470), .ZN(n9883) );
  XNOR2_X1 U5220 ( .A(n10209), .B(n10208), .ZN(n10205) );
  AOI22_X1 U5221 ( .A1(n4719), .A2(n10010), .B1(n5070), .B2(n9727), .ZN(n9965)
         );
  NOR3_X1 U5222 ( .A1(n5069), .A2(n5073), .A3(n4720), .ZN(n4719) );
  NAND2_X1 U5223 ( .A1(n9819), .A2(n5071), .ZN(n5070) );
  INV_X1 U5224 ( .A(n9665), .ZN(n5073) );
  INV_X1 U5225 ( .A(n7937), .ZN(n4863) );
  NAND2_X1 U5226 ( .A1(n4544), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n7903) );
  INV_X1 U5227 ( .A(n10114), .ZN(n7987) );
  NAND2_X1 U5228 ( .A1(n4645), .A2(n4459), .ZN(n10091) );
  OAI21_X1 U5229 ( .B1(n10154), .B2(n4647), .A(n4646), .ZN(n4645) );
  INV_X1 U5230 ( .A(n5289), .ZN(n4647) );
  NOR2_X1 U5231 ( .A1(n5299), .A2(n5293), .ZN(n5292) );
  NAND2_X1 U5232 ( .A1(n10131), .A2(n5300), .ZN(n5299) );
  INV_X1 U5233 ( .A(n7831), .ZN(n5300) );
  INV_X2 U5234 ( .A(n6744), .ZN(n9677) );
  AND2_X1 U5235 ( .A1(n6667), .A2(n9786), .ZN(n10187) );
  NOR2_X1 U5236 ( .A1(n7654), .A2(n7525), .ZN(n6060) );
  INV_X1 U5237 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n6275) );
  NAND2_X1 U5238 ( .A1(n10344), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6276) );
  AND2_X1 U5239 ( .A1(n5491), .A2(n5490), .ZN(n5912) );
  NAND2_X1 U5240 ( .A1(n5160), .A2(n5158), .ZN(n5878) );
  XNOR2_X1 U5241 ( .A(n6309), .B(n6308), .ZN(n6386) );
  INV_X1 U5242 ( .A(n4618), .ZN(n6307) );
  AOI21_X1 U5243 ( .B1(n6375), .B2(P1_IR_REG_31__SCAN_IN), .A(n4619), .ZN(
        n4618) );
  NAND2_X1 U5244 ( .A1(n5274), .A2(n6064), .ZN(n6375) );
  OAI21_X1 U5245 ( .B1(n8546), .B2(P2_REG2_REG_2__SCAN_IN), .A(n4763), .ZN(
        n8543) );
  NAND2_X1 U5246 ( .A1(n8546), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4763) );
  AOI21_X1 U5247 ( .B1(n8972), .B2(n8957), .A(n8714), .ZN(n4950) );
  NAND2_X1 U5248 ( .A1(n8367), .A2(n8372), .ZN(n5025) );
  NAND2_X1 U5249 ( .A1(n4673), .A2(n8481), .ZN(n8393) );
  NAND2_X1 U5250 ( .A1(n8390), .A2(n8389), .ZN(n4673) );
  NAND2_X1 U5251 ( .A1(n4478), .A2(n8494), .ZN(n4773) );
  NAND2_X1 U5252 ( .A1(n5022), .A2(n5021), .ZN(n8388) );
  NOR2_X1 U5253 ( .A1(n8383), .A2(n8384), .ZN(n5021) );
  NAND2_X1 U5254 ( .A1(n8447), .A2(n8444), .ZN(n5029) );
  AND2_X1 U5255 ( .A1(n8430), .A2(n8428), .ZN(n4774) );
  AND2_X1 U5256 ( .A1(n9642), .A2(n4876), .ZN(n4873) );
  NOR2_X1 U5257 ( .A1(n4878), .A2(n4877), .ZN(n4876) );
  NAND2_X1 U5258 ( .A1(n9753), .A2(n9688), .ZN(n4877) );
  INV_X1 U5259 ( .A(n9736), .ZN(n4878) );
  NOR2_X1 U5260 ( .A1(n4874), .A2(n4410), .ZN(n4870) );
  INV_X1 U5261 ( .A(n9642), .ZN(n4874) );
  AND2_X1 U5262 ( .A1(n9621), .A2(n9623), .ZN(n4875) );
  AOI21_X1 U5263 ( .B1(n8738), .B2(n8470), .A(n8494), .ZN(n4664) );
  NAND2_X1 U5264 ( .A1(n4893), .A2(n9746), .ZN(n4892) );
  NAND2_X1 U5265 ( .A1(n9660), .A2(n4894), .ZN(n4893) );
  INV_X1 U5266 ( .A(n9775), .ZN(n4894) );
  INV_X1 U5267 ( .A(n8480), .ZN(n5019) );
  NOR2_X1 U5268 ( .A1(n4739), .A2(n4735), .ZN(n4734) );
  INV_X1 U5269 ( .A(n5090), .ZN(n4735) );
  INV_X1 U5270 ( .A(n5097), .ZN(n4739) );
  INV_X1 U5271 ( .A(n9447), .ZN(n5181) );
  INV_X1 U5272 ( .A(n5185), .ZN(n5184) );
  OAI21_X1 U5273 ( .B1(n5328), .B2(n5186), .A(n9504), .ZN(n5185) );
  NAND2_X1 U5274 ( .A1(n9446), .A2(n9447), .ZN(n5186) );
  OR2_X1 U5275 ( .A1(n10243), .A2(n10025), .ZN(n9774) );
  INV_X1 U5276 ( .A(n9603), .ZN(n9702) );
  AND2_X1 U5277 ( .A1(n4416), .A2(n5486), .ZN(n4956) );
  INV_X1 U5278 ( .A(n5912), .ZN(n4959) );
  INV_X1 U5279 ( .A(n5163), .ZN(n5162) );
  OAI21_X1 U5280 ( .B1(n5165), .B2(n5164), .A(n5868), .ZN(n5163) );
  AND2_X1 U5281 ( .A1(n5176), .A2(n5326), .ZN(n5175) );
  NAND2_X1 U5282 ( .A1(n5774), .A2(n5457), .ZN(n5176) );
  INV_X1 U5283 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5458) );
  INV_X1 U5284 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n5452) );
  INV_X1 U5285 ( .A(n5152), .ZN(n5151) );
  OAI21_X1 U5286 ( .B1(n5154), .B2(n5153), .A(n5325), .ZN(n5152) );
  NAND2_X1 U5287 ( .A1(n4816), .A2(n4758), .ZN(n5413) );
  INV_X1 U5288 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4591) );
  INV_X1 U5289 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4590) );
  INV_X1 U5290 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5387) );
  NOR2_X1 U5291 ( .A1(n4436), .A2(n5098), .ZN(n5097) );
  INV_X1 U5292 ( .A(n5100), .ZN(n5098) );
  NOR2_X1 U5293 ( .A1(n5919), .A2(n8166), .ZN(n4827) );
  AND2_X1 U5294 ( .A1(n5341), .A2(n5340), .ZN(n5882) );
  INV_X1 U5295 ( .A(n8492), .ZN(n8315) );
  NAND2_X1 U5296 ( .A1(n5037), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5530) );
  OR3_X1 U5297 ( .A1(n6037), .A2(n6042), .A3(n6036), .ZN(n7742) );
  OR2_X1 U5298 ( .A1(n8996), .A2(n8741), .ZN(n8463) );
  OR2_X1 U5299 ( .A1(n5945), .A2(n5944), .ZN(n5963) );
  NOR2_X1 U5300 ( .A1(n8996), .A2(n9000), .ZN(n5270) );
  AND2_X1 U5301 ( .A1(n8463), .A2(n8468), .ZN(n8467) );
  AND2_X1 U5302 ( .A1(n8441), .A2(n8864), .ZN(n4940) );
  OR2_X1 U5303 ( .A1(n5261), .A2(n9032), .ZN(n5260) );
  INV_X1 U5304 ( .A(n8399), .ZN(n4943) );
  AND2_X1 U5305 ( .A1(n5129), .A2(n4946), .ZN(n4945) );
  NAND2_X1 U5306 ( .A1(n8399), .A2(n7629), .ZN(n4946) );
  NOR2_X1 U5307 ( .A1(n7680), .A2(n5130), .ZN(n5129) );
  INV_X1 U5308 ( .A(n8402), .ZN(n5130) );
  OAI22_X1 U5309 ( .A1(n5128), .A2(n7680), .B1(n9059), .B2(n8518), .ZN(n5127)
         );
  NAND2_X1 U5310 ( .A1(n7631), .A2(n8402), .ZN(n5128) );
  OR2_X1 U5311 ( .A1(n9054), .A2(n7700), .ZN(n8413) );
  NAND2_X1 U5312 ( .A1(n9059), .A2(n4574), .ZN(n4573) );
  INV_X1 U5313 ( .A(n9067), .ZN(n4574) );
  NAND2_X1 U5314 ( .A1(n9073), .A2(n7551), .ZN(n8399) );
  OR2_X1 U5315 ( .A1(n7645), .A2(n7554), .ZN(n8394) );
  NAND2_X1 U5316 ( .A1(n5337), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5681) );
  INV_X1 U5317 ( .A(n5656), .ZN(n5337) );
  AND2_X1 U5318 ( .A1(n8385), .A2(n8386), .ZN(n8325) );
  NOR2_X1 U5319 ( .A1(n7543), .A2(n7483), .ZN(n5264) );
  NAND2_X1 U5320 ( .A1(n5336), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5656) );
  INV_X1 U5321 ( .A(n5643), .ZN(n5336) );
  NAND2_X1 U5322 ( .A1(n8526), .A2(n7258), .ZN(n8370) );
  NAND2_X1 U5323 ( .A1(n8525), .A2(n10529), .ZN(n8372) );
  INV_X1 U5324 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5036) );
  INV_X1 U5325 ( .A(n8337), .ZN(n8350) );
  INV_X1 U5326 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5493) );
  NOR2_X1 U5327 ( .A1(n5354), .A2(n9103), .ZN(n5494) );
  INV_X1 U5328 ( .A(n4678), .ZN(n4577) );
  NOR2_X1 U5329 ( .A1(n4679), .A2(n4677), .ZN(n4575) );
  OR2_X1 U5330 ( .A1(n5738), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5792) );
  NAND2_X1 U5331 ( .A1(n5190), .A2(n4989), .ZN(n7465) );
  AND2_X1 U5332 ( .A1(n5188), .A2(n7170), .ZN(n4989) );
  INV_X1 U5333 ( .A(n9687), .ZN(n4538) );
  NAND2_X1 U5334 ( .A1(n4885), .A2(n4884), .ZN(n4883) );
  INV_X1 U5335 ( .A(n4886), .ZN(n4885) );
  INV_X1 U5336 ( .A(n4888), .ZN(n4884) );
  AOI22_X1 U5337 ( .A1(n4886), .A2(n4887), .B1(n4888), .B2(n9688), .ZN(n4881)
         );
  INV_X1 U5338 ( .A(n5157), .ZN(n4887) );
  AND2_X1 U5339 ( .A1(n6282), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4899) );
  INV_X1 U5340 ( .A(n6442), .ZN(n5010) );
  NAND2_X1 U5341 ( .A1(n10221), .A2(n9973), .ZN(n5053) );
  INV_X1 U5342 ( .A(n10238), .ZN(n8111) );
  OR2_X1 U5343 ( .A1(n10248), .A2(n10012), .ZN(n9747) );
  NOR2_X1 U5344 ( .A1(n10260), .A2(n10256), .ZN(n5047) );
  NOR2_X1 U5345 ( .A1(n5046), .A2(n5048), .ZN(n5045) );
  INV_X1 U5346 ( .A(n5047), .ZN(n5046) );
  OR2_X1 U5347 ( .A1(n10256), .A2(n9521), .ZN(n9768) );
  OR2_X1 U5348 ( .A1(n9761), .A2(n5068), .ZN(n5067) );
  NAND2_X1 U5349 ( .A1(n4704), .A2(n4706), .ZN(n4703) );
  INV_X1 U5350 ( .A(n9601), .ZN(n4706) );
  AND2_X1 U5351 ( .A1(n6950), .A2(n4705), .ZN(n4704) );
  AND2_X1 U5352 ( .A1(n9808), .A2(n6662), .ZN(n4705) );
  OR2_X1 U5353 ( .A1(n9851), .A2(n6990), .ZN(n9808) );
  OR2_X1 U5354 ( .A1(n6659), .A2(n6660), .ZN(n9803) );
  NAND2_X1 U5355 ( .A1(n4880), .A2(n9801), .ZN(n6950) );
  AND3_X1 U5356 ( .A1(n6662), .A2(n9800), .A3(n9799), .ZN(n4880) );
  OR2_X1 U5357 ( .A1(n6663), .A2(n10447), .ZN(n6694) );
  NAND2_X1 U5358 ( .A1(n7858), .A2(n6382), .ZN(n6383) );
  NAND2_X1 U5359 ( .A1(n4965), .A2(SI_29_), .ZN(n8299) );
  INV_X1 U5360 ( .A(n8011), .ZN(n4965) );
  NAND2_X1 U5361 ( .A1(n7713), .A2(n7712), .ZN(n7725) );
  OAI21_X1 U5362 ( .B1(n5936), .B2(n5935), .A(n5934), .ZN(n5954) );
  INV_X1 U5363 ( .A(n5931), .ZN(n5935) );
  AND2_X1 U5364 ( .A1(n5213), .A2(n5209), .ZN(n5208) );
  INV_X1 U5365 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5209) );
  NAND2_X1 U5366 ( .A1(n5474), .A2(n5473), .ZN(n5849) );
  INV_X1 U5367 ( .A(n5834), .ZN(n5467) );
  INV_X1 U5368 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6305) );
  AOI21_X1 U5369 ( .B1(n5175), .B2(n5173), .A(n5172), .ZN(n5171) );
  INV_X1 U5370 ( .A(n5463), .ZN(n5172) );
  INV_X1 U5371 ( .A(n5457), .ZN(n5173) );
  INV_X1 U5372 ( .A(n5175), .ZN(n5174) );
  NAND2_X1 U5373 ( .A1(n5454), .A2(n5453), .ZN(n5457) );
  INV_X1 U5374 ( .A(SI_15_), .ZN(n5453) );
  NOR2_X1 U5375 ( .A1(n6193), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n6187) );
  XNOR2_X1 U5376 ( .A(n5413), .B(n4641), .ZN(n5412) );
  INV_X1 U5377 ( .A(SI_6_), .ZN(n4641) );
  INV_X1 U5378 ( .A(n5582), .ZN(n5409) );
  NAND2_X1 U5379 ( .A1(n10343), .A2(n4550), .ZN(n4549) );
  INV_X1 U5380 ( .A(n6979), .ZN(n4804) );
  INV_X1 U5381 ( .A(n7084), .ZN(n4805) );
  XNOR2_X1 U5382 ( .A(n4746), .B(n7645), .ZN(n5688) );
  NAND2_X1 U5383 ( .A1(n8251), .A2(n8250), .ZN(n5091) );
  NAND2_X1 U5384 ( .A1(n8259), .A2(n5974), .ZN(n5995) );
  AOI21_X1 U5385 ( .B1(n5994), .B2(n5993), .A(n7741), .ZN(n5996) );
  AOI22_X1 U5386 ( .A1(n5523), .A2(n7050), .B1(n7729), .B2(n6487), .ZN(n6612)
         );
  NAND2_X1 U5387 ( .A1(n4827), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5945) );
  INV_X1 U5388 ( .A(n4827), .ZN(n5921) );
  AND2_X1 U5389 ( .A1(n5691), .A2(n5715), .ZN(n5085) );
  INV_X1 U5390 ( .A(n5817), .ZN(n4726) );
  NAND2_X1 U5391 ( .A1(n5334), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5621) );
  INV_X1 U5392 ( .A(n5606), .ZN(n5334) );
  NAND2_X1 U5393 ( .A1(n8188), .A2(n8189), .ZN(n4732) );
  NAND2_X1 U5394 ( .A1(n5952), .A2(n5951), .ZN(n4730) );
  NAND2_X1 U5395 ( .A1(n5135), .A2(n4425), .ZN(n5141) );
  NOR2_X1 U5396 ( .A1(n8315), .A2(n8340), .ZN(n5120) );
  AOI21_X1 U5397 ( .B1(n5118), .B2(n5120), .A(n5117), .ZN(n5116) );
  AND2_X1 U5398 ( .A1(n8315), .A2(n8340), .ZN(n5117) );
  INV_X1 U5399 ( .A(n8489), .ZN(n5118) );
  OAI211_X1 U5400 ( .C1(n8499), .C2(n4660), .A(n4815), .B(n4661), .ZN(n5122)
         );
  NAND2_X1 U5401 ( .A1(n8500), .A2(n8497), .ZN(n4661) );
  NAND2_X1 U5402 ( .A1(n8500), .A2(n4741), .ZN(n4660) );
  AND2_X1 U5403 ( .A1(n5970), .A2(n5969), .ZN(n8193) );
  OR2_X1 U5404 ( .A1(n8262), .A2(n5965), .ZN(n5970) );
  AND3_X1 U5405 ( .A1(n5844), .A2(n5843), .A3(n5842), .ZN(n8214) );
  INV_X1 U5406 ( .A(n6921), .ZN(n4555) );
  INV_X1 U5407 ( .A(n4558), .ZN(n4557) );
  OAI21_X1 U5408 ( .B1(n4559), .B2(n6854), .A(n6857), .ZN(n4558) );
  NOR2_X1 U5409 ( .A1(n6933), .A2(n4811), .ZN(n8652) );
  AND2_X1 U5410 ( .A1(n6858), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4811) );
  AND2_X1 U5411 ( .A1(n8504), .A2(n8350), .ZN(n6814) );
  NAND2_X1 U5412 ( .A1(n7606), .A2(n4560), .ZN(n7611) );
  NAND2_X1 U5413 ( .A1(n7603), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4560) );
  NAND2_X1 U5414 ( .A1(n7611), .A2(n7610), .ZN(n7668) );
  NAND2_X1 U5415 ( .A1(n8292), .A2(n8291), .ZN(n8694) );
  NOR2_X1 U5416 ( .A1(n8978), .A2(n8728), .ZN(n8973) );
  INV_X1 U5417 ( .A(n4685), .ZN(n4684) );
  OAI21_X1 U5418 ( .B1(n8738), .B2(n4686), .A(n8717), .ZN(n4685) );
  NAND2_X1 U5419 ( .A1(n8470), .A2(n8472), .ZN(n8738) );
  NAND2_X1 U5420 ( .A1(n8733), .A2(n8738), .ZN(n8735) );
  NAND2_X1 U5421 ( .A1(n4518), .A2(n8466), .ZN(n4586) );
  NAND2_X1 U5422 ( .A1(n4516), .A2(n4460), .ZN(n4584) );
  INV_X1 U5423 ( .A(n8467), .ZN(n8765) );
  NAND2_X1 U5424 ( .A1(n4589), .A2(n4588), .ZN(n8783) );
  NAND2_X1 U5425 ( .A1(n7788), .A2(n4413), .ZN(n4588) );
  NAND2_X1 U5426 ( .A1(n4516), .A2(n4400), .ZN(n4589) );
  NOR2_X1 U5427 ( .A1(n8775), .A2(n4921), .ZN(n4920) );
  INV_X1 U5428 ( .A(n7769), .ZN(n4921) );
  NOR2_X1 U5429 ( .A1(n8792), .A2(n5246), .ZN(n5245) );
  INV_X1 U5430 ( .A(n7767), .ZN(n5246) );
  NAND2_X1 U5431 ( .A1(n5244), .A2(n5243), .ZN(n8802) );
  AND2_X1 U5432 ( .A1(n8803), .A2(n4417), .ZN(n5243) );
  NOR2_X1 U5433 ( .A1(n8895), .A2(n8214), .ZN(n5231) );
  AND2_X1 U5434 ( .A1(n8440), .A2(n8846), .ZN(n8864) );
  NAND2_X1 U5435 ( .A1(n4824), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5824) );
  INV_X1 U5436 ( .A(n5804), .ZN(n4824) );
  NAND2_X1 U5437 ( .A1(n7781), .A2(n5133), .ZN(n5132) );
  NOR2_X1 U5438 ( .A1(n7783), .A2(n5134), .ZN(n5133) );
  INV_X1 U5439 ( .A(n7780), .ZN(n5134) );
  INV_X1 U5440 ( .A(n7704), .ZN(n4779) );
  NOR2_X1 U5441 ( .A1(n8928), .A2(n5242), .ZN(n5241) );
  INV_X1 U5442 ( .A(n7759), .ZN(n5242) );
  AND3_X1 U5443 ( .A1(n5829), .A2(n5828), .A3(n5827), .ZN(n8927) );
  NAND2_X1 U5444 ( .A1(n5338), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5781) );
  INV_X1 U5445 ( .A(n5762), .ZN(n5338) );
  OR2_X1 U5446 ( .A1(n9054), .A2(n8517), .ZN(n4928) );
  NOR2_X1 U5447 ( .A1(n7683), .A2(n4925), .ZN(n4924) );
  NAND2_X1 U5448 ( .A1(n7697), .A2(n8420), .ZN(n7781) );
  NAND2_X1 U5449 ( .A1(n7694), .A2(n8413), .ZN(n7697) );
  INV_X1 U5450 ( .A(n8420), .ZN(n7702) );
  AND4_X1 U5451 ( .A1(n5746), .A2(n5745), .A3(n5744), .A4(n5743), .ZN(n8156)
         );
  NAND2_X1 U5452 ( .A1(n4927), .A2(n5216), .ZN(n7623) );
  INV_X1 U5453 ( .A(n4930), .ZN(n4927) );
  AOI22_X1 U5454 ( .A1(n8327), .A2(n7619), .B1(n9073), .B2(n8520), .ZN(n7620)
         );
  NAND2_X1 U5455 ( .A1(n8398), .A2(n8399), .ZN(n8327) );
  NAND2_X1 U5456 ( .A1(n8390), .A2(n8394), .ZN(n8328) );
  NAND2_X1 U5457 ( .A1(n4689), .A2(n4688), .ZN(n7486) );
  NAND2_X1 U5458 ( .A1(n4690), .A2(n7484), .ZN(n4689) );
  NAND2_X1 U5459 ( .A1(n7486), .A2(n7492), .ZN(n7553) );
  INV_X1 U5460 ( .A(n8525), .ZN(n7451) );
  NAND2_X1 U5461 ( .A1(n7294), .A2(n5214), .ZN(n7446) );
  NAND2_X1 U5462 ( .A1(n8316), .A2(n10523), .ZN(n6097) );
  NAND2_X1 U5463 ( .A1(n8337), .A2(n8339), .ZN(n6107) );
  OR2_X1 U5464 ( .A1(n6379), .A2(n5560), .ZN(n4514) );
  INV_X1 U5465 ( .A(n4513), .ZN(n4512) );
  OAI22_X1 U5466 ( .A1(n5941), .A2(n6121), .B1(n6838), .B2(n6861), .ZN(n4513)
         );
  INV_X1 U5467 ( .A(n8926), .ZN(n8888) );
  NAND2_X1 U5468 ( .A1(n5984), .A2(n5983), .ZN(n8984) );
  INV_X1 U5469 ( .A(n8407), .ZN(n9059) );
  NAND2_X1 U5470 ( .A1(n4780), .A2(n8307), .ZN(n5247) );
  NAND2_X1 U5471 ( .A1(n5040), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5356) );
  AND2_X1 U5472 ( .A1(n5256), .A2(n5493), .ZN(n5039) );
  AND2_X2 U5473 ( .A1(n4511), .A2(n4510), .ZN(n5999) );
  NOR2_X1 U5474 ( .A1(n4678), .A2(n5348), .ZN(n4511) );
  NOR2_X1 U5475 ( .A1(n4679), .A2(n4677), .ZN(n4510) );
  NAND2_X1 U5476 ( .A1(n6006), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6024) );
  AND2_X1 U5477 ( .A1(n5352), .A2(n5351), .ZN(n4680) );
  INV_X1 U5478 ( .A(n4679), .ZN(n4676) );
  NAND2_X1 U5479 ( .A1(n5636), .A2(n5369), .ZN(n5381) );
  NOR2_X2 U5480 ( .A1(n5617), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5636) );
  NOR2_X2 U5481 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n4792) );
  NAND2_X1 U5482 ( .A1(n5190), .A2(n5188), .ZN(n7178) );
  AND2_X1 U5483 ( .A1(n4474), .A2(n9456), .ZN(n4917) );
  NOR2_X1 U5484 ( .A1(n5205), .A2(n4914), .ZN(n4913) );
  INV_X1 U5485 ( .A(n8110), .ZN(n4914) );
  NAND2_X1 U5486 ( .A1(n7465), .A2(n7202), .ZN(n7458) );
  NAND2_X1 U5487 ( .A1(n4907), .A2(n4906), .ZN(n4905) );
  INV_X1 U5488 ( .A(n8069), .ZN(n5199) );
  INV_X1 U5489 ( .A(n5196), .ZN(n5195) );
  NAND2_X1 U5490 ( .A1(n9488), .A2(n8110), .ZN(n4918) );
  NAND2_X1 U5491 ( .A1(n8045), .A2(n4983), .ZN(n4982) );
  NOR2_X1 U5492 ( .A1(n4985), .A2(n4984), .ZN(n4983) );
  AND2_X1 U5493 ( .A1(n6501), .A2(n6500), .ZN(n6577) );
  INV_X1 U5494 ( .A(n6390), .ZN(n6391) );
  NAND2_X1 U5495 ( .A1(n8084), .A2(n6654), .ZN(n6392) );
  OR2_X1 U5496 ( .A1(n8123), .A2(n6655), .ZN(n6397) );
  NOR2_X1 U5497 ( .A1(n6407), .A2(n6627), .ZN(n6408) );
  NAND2_X1 U5498 ( .A1(n6466), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6471) );
  NAND2_X1 U5499 ( .A1(n6466), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6286) );
  AND2_X1 U5500 ( .A1(n6241), .A2(n6240), .ZN(n6289) );
  NAND2_X1 U5501 ( .A1(n4505), .A2(n4546), .ZN(n9876) );
  INV_X1 U5502 ( .A(n6423), .ZN(n4546) );
  NOR2_X1 U5503 ( .A1(n6441), .A2(n5013), .ZN(n5012) );
  INV_X1 U5504 ( .A(n6426), .ZN(n5013) );
  XNOR2_X1 U5505 ( .A(n7592), .B(n7806), .ZN(n7155) );
  NAND2_X1 U5506 ( .A1(n5004), .A2(n5003), .ZN(n5002) );
  NAND2_X1 U5507 ( .A1(n9885), .A2(n9891), .ZN(n5003) );
  OR2_X1 U5508 ( .A1(n9915), .A2(n4503), .ZN(n5000) );
  OAI21_X1 U5509 ( .B1(n4996), .B2(n9917), .A(n4992), .ZN(n4991) );
  NAND2_X1 U5510 ( .A1(n9915), .A2(n4432), .ZN(n4995) );
  NAND2_X1 U5511 ( .A1(n4998), .A2(n4431), .ZN(n4994) );
  NOR2_X1 U5512 ( .A1(n5074), .A2(n7858), .ZN(n9689) );
  INV_X1 U5513 ( .A(n9561), .ZN(n5074) );
  NAND2_X1 U5514 ( .A1(n9566), .A2(n9565), .ZN(n9939) );
  AND2_X1 U5515 ( .A1(n9978), .A2(n5050), .ZN(n9947) );
  NOR2_X1 U5516 ( .A1(n5053), .A2(n5051), .ZN(n5050) );
  NAND2_X1 U5517 ( .A1(n5156), .A2(n9984), .ZN(n5051) );
  NAND2_X1 U5518 ( .A1(n9948), .A2(n4540), .ZN(n8139) );
  OAI21_X1 U5519 ( .B1(n7967), .B2(n9398), .A(n7966), .ZN(n4540) );
  NAND2_X1 U5520 ( .A1(n4716), .A2(n9952), .ZN(n4715) );
  NAND2_X1 U5521 ( .A1(n7996), .A2(n9576), .ZN(n4716) );
  INV_X1 U5522 ( .A(n9988), .ZN(n4821) );
  NAND2_X1 U5523 ( .A1(n9990), .A2(n10189), .ZN(n4819) );
  NAND2_X1 U5524 ( .A1(n4649), .A2(n4650), .ZN(n7938) );
  INV_X1 U5525 ( .A(n5304), .ZN(n4652) );
  NAND2_X1 U5526 ( .A1(n9577), .A2(n10025), .ZN(n5310) );
  NAND2_X1 U5527 ( .A1(n5304), .A2(n5302), .ZN(n5301) );
  INV_X1 U5528 ( .A(n5308), .ZN(n5302) );
  NAND2_X1 U5529 ( .A1(n9985), .A2(n9665), .ZN(n9996) );
  INV_X1 U5530 ( .A(n4541), .ZN(n7915) );
  NOR2_X1 U5531 ( .A1(n7910), .A2(n5309), .ZN(n5308) );
  INV_X1 U5532 ( .A(n7897), .ZN(n5309) );
  OAI21_X1 U5533 ( .B1(n7910), .B2(n5307), .A(n9578), .ZN(n5306) );
  NAND2_X1 U5534 ( .A1(n7898), .A2(n7897), .ZN(n5307) );
  NAND2_X1 U5535 ( .A1(n4484), .A2(n4412), .ZN(n4852) );
  AND2_X1 U5536 ( .A1(n10050), .A2(n9692), .ZN(n10072) );
  INV_X1 U5537 ( .A(n4405), .ZN(n5077) );
  AOI21_X1 U5538 ( .B1(n4405), .B2(n5076), .A(n9637), .ZN(n5075) );
  AND2_X1 U5539 ( .A1(n4648), .A2(n5297), .ZN(n5289) );
  NAND2_X1 U5540 ( .A1(n5292), .A2(n7818), .ZN(n4648) );
  AND2_X1 U5541 ( .A1(n7986), .A2(n10098), .ZN(n10113) );
  NAND2_X1 U5542 ( .A1(n6351), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7844) );
  INV_X1 U5543 ( .A(n7836), .ZN(n6351) );
  NAND2_X1 U5544 ( .A1(n9756), .A2(n9636), .ZN(n10131) );
  NAND2_X1 U5545 ( .A1(n5294), .A2(n5291), .ZN(n10141) );
  INV_X1 U5546 ( .A(n5293), .ZN(n5291) );
  NAND2_X1 U5547 ( .A1(n5296), .A2(n5295), .ZN(n5294) );
  NAND2_X1 U5548 ( .A1(n7984), .A2(n4401), .ZN(n5080) );
  AOI21_X1 U5549 ( .B1(n4401), .B2(n7983), .A(n9628), .ZN(n5079) );
  AND2_X1 U5550 ( .A1(n7809), .A2(n7808), .ZN(n10156) );
  OAI22_X1 U5551 ( .A1(n7806), .A2(n6380), .B1(n9680), .B2(n7805), .ZN(n7807)
         );
  OAI22_X1 U5552 ( .A1(n10173), .A2(n7803), .B1(n10183), .B2(n10166), .ZN(
        n10154) );
  OR2_X1 U5553 ( .A1(n7984), .A2(n7983), .ZN(n5081) );
  AOI21_X1 U5554 ( .B1(n10303), .B2(n10188), .A(n10307), .ZN(n10173) );
  NAND2_X1 U5555 ( .A1(n4840), .A2(n7347), .ZN(n7424) );
  NOR2_X1 U5556 ( .A1(n5285), .A2(n5284), .ZN(n5283) );
  INV_X1 U5557 ( .A(n7353), .ZN(n5285) );
  INV_X1 U5558 ( .A(n7409), .ZN(n5284) );
  NAND2_X1 U5559 ( .A1(n4845), .A2(n5282), .ZN(n4837) );
  NAND2_X1 U5560 ( .A1(n4483), .A2(n7409), .ZN(n5282) );
  AND2_X1 U5561 ( .A1(n9625), .A2(n9623), .ZN(n9707) );
  OAI211_X1 U5562 ( .C1(n7239), .C2(n4700), .A(n4697), .B(n9611), .ZN(n4696)
         );
  INV_X1 U5563 ( .A(n9733), .ZN(n4700) );
  AND2_X1 U5564 ( .A1(n9612), .A2(n4698), .ZN(n4697) );
  AND4_X1 U5565 ( .A1(n7376), .A2(n7375), .A3(n7374), .A4(n7373), .ZN(n8030)
         );
  OR2_X1 U5566 ( .A1(n7186), .A2(n7185), .ZN(n7210) );
  INV_X1 U5567 ( .A(n6713), .ZN(n5281) );
  AND2_X1 U5568 ( .A1(n9808), .A2(n9810), .ZN(n9699) );
  NAND2_X1 U5569 ( .A1(n6712), .A2(n9695), .ZN(n6714) );
  AND2_X1 U5570 ( .A1(n4623), .A2(n6386), .ZN(n4622) );
  NAND2_X1 U5571 ( .A1(n6696), .A2(n7721), .ZN(n4623) );
  INV_X1 U5572 ( .A(n10187), .ZN(n10167) );
  NOR2_X1 U5573 ( .A1(n10458), .A2(n10007), .ZN(n6632) );
  AND2_X1 U5574 ( .A1(n4492), .A2(n4856), .ZN(n10207) );
  AOI21_X1 U5575 ( .B1(n9959), .B2(n10192), .A(n9958), .ZN(n10217) );
  INV_X1 U5576 ( .A(n10223), .ZN(n4799) );
  NAND2_X1 U5577 ( .A1(n7940), .A2(n7939), .ZN(n10231) );
  NAND2_X1 U5578 ( .A1(n9117), .A2(n9677), .ZN(n7940) );
  INV_X1 U5579 ( .A(n10480), .ZN(n10463) );
  AND3_X1 U5580 ( .A1(n6585), .A2(n6584), .A3(n6583), .ZN(n10457) );
  OR2_X1 U5581 ( .A1(n6329), .A2(n9832), .ZN(n10480) );
  AND2_X1 U5582 ( .A1(n6311), .A2(n6310), .ZN(n6676) );
  AND2_X1 U5583 ( .A1(n5313), .A2(n6076), .ZN(n5312) );
  INV_X1 U5584 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n6277) );
  AND2_X1 U5585 ( .A1(n6074), .A2(n6078), .ZN(n5313) );
  INV_X1 U5586 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6056) );
  NAND2_X1 U5587 ( .A1(n4961), .A2(n5481), .ZN(n4960) );
  INV_X1 U5588 ( .A(n5890), .ZN(n4961) );
  NAND2_X1 U5589 ( .A1(n6305), .A2(n5213), .ZN(n4621) );
  INV_X1 U5590 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6050) );
  OAI21_X1 U5591 ( .B1(n6191), .B2(P1_IR_REG_12__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6270) );
  NAND2_X1 U5592 ( .A1(n5436), .A2(n5154), .ZN(n5150) );
  XNOR2_X1 U5593 ( .A(n5700), .B(n5699), .ZN(n7354) );
  XNOR2_X1 U5594 ( .A(n5678), .B(n5677), .ZN(n7349) );
  NAND2_X1 U5595 ( .A1(n5675), .A2(n5674), .ZN(n5678) );
  OAI21_X1 U5596 ( .B1(n5635), .B2(n4671), .A(n4669), .ZN(n5675) );
  NAND2_X1 U5597 ( .A1(n5635), .A2(n4672), .ZN(n5694) );
  INV_X1 U5598 ( .A(n4629), .ZN(n10382) );
  OAI21_X1 U5599 ( .B1(n10592), .B2(n10593), .A(n4481), .ZN(n4629) );
  NAND2_X1 U5600 ( .A1(n10577), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n10384) );
  NAND2_X1 U5601 ( .A1(n6115), .A2(n5614), .ZN(n5106) );
  NAND2_X1 U5602 ( .A1(n5915), .A2(n5914), .ZN(n9005) );
  AND2_X1 U5603 ( .A1(n5992), .A2(n5991), .ZN(n7741) );
  NAND2_X1 U5604 ( .A1(n5995), .A2(n5996), .ZN(n7758) );
  NAND2_X1 U5605 ( .A1(n5880), .A2(n5879), .ZN(n9015) );
  NOR2_X1 U5606 ( .A1(n5929), .A2(n4795), .ZN(n8191) );
  AND2_X1 U5607 ( .A1(n8221), .A2(n5930), .ZN(n4795) );
  NAND2_X1 U5608 ( .A1(n4740), .A2(n5654), .ZN(n7567) );
  NAND2_X1 U5609 ( .A1(n9389), .A2(n8307), .ZN(n4740) );
  NAND2_X1 U5610 ( .A1(n5871), .A2(n5870), .ZN(n9022) );
  AND2_X1 U5611 ( .A1(n5889), .A2(n5888), .ZN(n8850) );
  NAND2_X1 U5612 ( .A1(n5893), .A2(n5892), .ZN(n9010) );
  INV_X1 U5613 ( .A(n7561), .ZN(n9073) );
  AND2_X1 U5614 ( .A1(n5860), .A2(n5859), .ZN(n8848) );
  AND2_X1 U5615 ( .A1(n6604), .A2(n6028), .ZN(n8280) );
  NAND2_X1 U5616 ( .A1(n6841), .A2(n4561), .ZN(n8570) );
  AND2_X1 U5617 ( .A1(n4563), .A2(n4562), .ZN(n4561) );
  NAND2_X1 U5618 ( .A1(n8559), .A2(n6842), .ZN(n4562) );
  NAND2_X1 U5619 ( .A1(n8713), .A2(n8712), .ZN(n4951) );
  OR2_X1 U5620 ( .A1(n8880), .A2(n5227), .ZN(n5221) );
  NAND2_X1 U5621 ( .A1(n5604), .A2(n5603), .ZN(n7272) );
  NAND2_X1 U5622 ( .A1(n6861), .A2(n4419), .ZN(n4580) );
  AND2_X1 U5623 ( .A1(n7049), .A2(n4796), .ZN(n8957) );
  NAND2_X1 U5624 ( .A1(n8940), .A2(n6103), .ZN(n8899) );
  AND2_X2 U5625 ( .A1(n6486), .A2(n6485), .ZN(n10544) );
  AND2_X1 U5626 ( .A1(n4771), .A2(n8974), .ZN(n4519) );
  INV_X1 U5627 ( .A(n8982), .ZN(n4611) );
  INV_X1 U5628 ( .A(n7232), .ZN(n10473) );
  INV_X1 U5629 ( .A(n9845), .ZN(n10166) );
  INV_X1 U5630 ( .A(n8035), .ZN(n9407) );
  INV_X1 U5631 ( .A(n10156), .ZN(n10292) );
  INV_X1 U5632 ( .A(n9844), .ZN(n10168) );
  AND3_X1 U5633 ( .A1(n7856), .A2(n7855), .A3(n7854), .ZN(n9482) );
  INV_X1 U5634 ( .A(n6663), .ZN(n6655) );
  NAND2_X1 U5635 ( .A1(n7850), .A2(n7849), .ZN(n10270) );
  INV_X1 U5636 ( .A(n9558), .ZN(n9507) );
  AND2_X1 U5637 ( .A1(n7936), .A2(n7935), .ZN(n10013) );
  OR2_X1 U5638 ( .A1(n9998), .A2(n6593), .ZN(n7936) );
  AND4_X1 U5639 ( .A1(n7817), .A2(n7816), .A3(n7815), .A4(n7814), .ZN(n10138)
         );
  NAND2_X1 U5640 ( .A1(n7821), .A2(n7820), .ZN(n10285) );
  INV_X1 U5641 ( .A(n8138), .ZN(n9990) );
  INV_X1 U5642 ( .A(n10013), .ZN(n9989) );
  AND2_X1 U5643 ( .A1(n6358), .A2(n6357), .ZN(n10055) );
  NAND2_X1 U5644 ( .A1(n7878), .A2(n7877), .ZN(n10086) );
  INV_X1 U5645 ( .A(n10138), .ZN(n10190) );
  INV_X1 U5646 ( .A(n8030), .ZN(n10188) );
  NAND4_X2 U5647 ( .A1(n6517), .A2(n6516), .A3(n6515), .A4(n6514), .ZN(n9852)
         );
  NAND2_X1 U5648 ( .A1(n6222), .A2(n6258), .ZN(n6262) );
  OAI21_X1 U5649 ( .B1(n10411), .B2(n4592), .A(n9933), .ZN(n4789) );
  NAND2_X1 U5650 ( .A1(n4714), .A2(n4711), .ZN(n10224) );
  NOR2_X1 U5651 ( .A1(n4713), .A2(n4712), .ZN(n4711) );
  NAND2_X1 U5652 ( .A1(n4715), .A2(n10192), .ZN(n4714) );
  NOR2_X1 U5653 ( .A1(n8138), .A2(n10167), .ZN(n4712) );
  OR2_X1 U5654 ( .A1(n10458), .A2(n6404), .ZN(n10157) );
  AND3_X2 U5655 ( .A1(n6630), .A2(n10443), .A3(n6679), .ZN(n10488) );
  CLKBUF_X1 U5656 ( .A(n6386), .Z(n10059) );
  NOR2_X1 U5657 ( .A1(n10571), .A2(n4508), .ZN(n10570) );
  OR2_X1 U5658 ( .A1(n10570), .A2(n10569), .ZN(n4635) );
  OAI21_X1 U5659 ( .B1(n5026), .B2(n5024), .A(n5023), .ZN(n5022) );
  INV_X1 U5660 ( .A(n8377), .ZN(n5023) );
  INV_X1 U5661 ( .A(n8378), .ZN(n5026) );
  NOR2_X1 U5662 ( .A1(n4814), .A2(n8405), .ZN(n5031) );
  NAND2_X1 U5663 ( .A1(n8406), .A2(n4456), .ZN(n4814) );
  OAI21_X1 U5664 ( .B1(n8396), .B2(n8494), .A(n4773), .ZN(n5035) );
  AND2_X1 U5665 ( .A1(n8420), .A2(n8414), .ZN(n4769) );
  INV_X1 U5666 ( .A(n9589), .ZN(n4897) );
  NOR2_X1 U5667 ( .A1(n9588), .A2(n4896), .ZN(n4895) );
  OR2_X1 U5668 ( .A1(n9587), .A2(n9688), .ZN(n4896) );
  OAI21_X1 U5669 ( .B1(n8446), .B2(n8445), .A(n5028), .ZN(n4659) );
  NOR2_X1 U5670 ( .A1(n5029), .A2(n4471), .ZN(n5028) );
  NAND2_X1 U5671 ( .A1(n8465), .A2(n5027), .ZN(n8469) );
  AND2_X1 U5672 ( .A1(n8467), .A2(n8466), .ZN(n5027) );
  AND2_X1 U5673 ( .A1(n4871), .A2(n4869), .ZN(n9656) );
  INV_X1 U5674 ( .A(n9661), .ZN(n4745) );
  NAND2_X1 U5675 ( .A1(n4892), .A2(n4890), .ZN(n9662) );
  NOR2_X1 U5676 ( .A1(n9661), .A2(n4891), .ZN(n4890) );
  AND2_X1 U5677 ( .A1(n9611), .A2(n7428), .ZN(n9750) );
  NAND2_X1 U5678 ( .A1(n5097), .A2(n4738), .ZN(n4737) );
  NAND2_X1 U5679 ( .A1(n4665), .A2(n5017), .ZN(n5016) );
  NOR2_X1 U5680 ( .A1(n5019), .A2(n5018), .ZN(n5017) );
  NAND2_X1 U5681 ( .A1(n8963), .A2(n8689), .ZN(n8492) );
  NAND2_X1 U5682 ( .A1(n4976), .A2(n8311), .ZN(n8485) );
  INV_X1 U5683 ( .A(n8963), .ZN(n4976) );
  NOR2_X1 U5684 ( .A1(n5018), .A2(n8335), .ZN(n4974) );
  NAND2_X1 U5685 ( .A1(n8487), .A2(n8492), .ZN(n8486) );
  INV_X1 U5686 ( .A(n5348), .ZN(n4576) );
  NOR2_X1 U5687 ( .A1(n4911), .A2(n5193), .ZN(n4910) );
  OAI21_X1 U5688 ( .B1(n4408), .B2(n4980), .A(n9440), .ZN(n4911) );
  NAND2_X1 U5689 ( .A1(n10208), .A2(n9683), .ZN(n5157) );
  NOR2_X1 U5690 ( .A1(n7844), .A2(n9481), .ZN(n4545) );
  AND2_X1 U5691 ( .A1(n9612), .A2(n9610), .ZN(n7428) );
  NAND2_X1 U5692 ( .A1(n7239), .A2(n9607), .ZN(n7280) );
  NAND2_X1 U5693 ( .A1(n7280), .A2(n7279), .ZN(n9589) );
  INV_X1 U5694 ( .A(n5474), .ZN(n5164) );
  INV_X1 U5695 ( .A(n5451), .ZN(n4973) );
  INV_X1 U5696 ( .A(SI_16_), .ZN(n5459) );
  INV_X1 U5697 ( .A(n5442), .ZN(n5153) );
  INV_X1 U5698 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5443) );
  OAI21_X1 U5699 ( .B1(n4395), .B2(P1_DATAO_REG_12__SCAN_IN), .A(n4801), .ZN(
        n5439) );
  NAND2_X1 U5700 ( .A1(n4397), .A2(n5437), .ZN(n4801) );
  INV_X1 U5701 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5437) );
  AND2_X1 U5702 ( .A1(n5412), .A2(n4954), .ZN(n4813) );
  NAND2_X1 U5703 ( .A1(n5388), .A2(n5387), .ZN(n5252) );
  NAND2_X1 U5704 ( .A1(n5389), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5168) );
  NAND2_X1 U5705 ( .A1(n4592), .A2(n4591), .ZN(n5388) );
  NAND2_X1 U5706 ( .A1(n4590), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n5389) );
  OR2_X1 U5707 ( .A1(n4436), .A2(n5099), .ZN(n5096) );
  NAND2_X1 U5708 ( .A1(n5097), .A2(n8232), .ZN(n5095) );
  AND2_X1 U5709 ( .A1(n8179), .A2(n5911), .ZN(n5099) );
  AND2_X1 U5710 ( .A1(n5866), .A2(n5848), .ZN(n5090) );
  NOR2_X1 U5711 ( .A1(n4433), .A2(n5103), .ZN(n5102) );
  INV_X1 U5712 ( .A(n5773), .ZN(n5103) );
  OR2_X1 U5713 ( .A1(n8971), .A2(n8508), .ZN(n8483) );
  AND2_X1 U5714 ( .A1(n5269), .A2(n5270), .ZN(n5268) );
  NAND2_X1 U5715 ( .A1(n4939), .A2(n4938), .ZN(n4937) );
  INV_X1 U5716 ( .A(n4940), .ZN(n4938) );
  INV_X1 U5717 ( .A(n4826), .ZN(n5854) );
  INV_X1 U5718 ( .A(n7678), .ZN(n4925) );
  INV_X1 U5719 ( .A(n5220), .ZN(n5219) );
  INV_X1 U5720 ( .A(n7629), .ZN(n8398) );
  INV_X1 U5721 ( .A(n8328), .ZN(n7575) );
  AND2_X1 U5722 ( .A1(n8380), .A2(n8325), .ZN(n7302) );
  AND2_X1 U5723 ( .A1(n8391), .A2(n8389), .ZN(n8324) );
  NAND2_X1 U5724 ( .A1(n8380), .A2(n8379), .ZN(n8321) );
  NAND2_X1 U5725 ( .A1(n7451), .A2(n7272), .ZN(n8376) );
  NAND2_X1 U5726 ( .A1(n4509), .A2(n5142), .ZN(n7298) );
  NOR2_X1 U5727 ( .A1(n7110), .A2(n5143), .ZN(n5142) );
  AND2_X1 U5728 ( .A1(n10518), .A2(n6487), .ZN(n5253) );
  INV_X1 U5729 ( .A(n4807), .ZN(n4760) );
  AOI21_X1 U5730 ( .B1(n8510), .B2(n8886), .A(n4808), .ZN(n4807) );
  NOR2_X1 U5731 ( .A1(n8508), .A2(n8926), .ZN(n4808) );
  NOR2_X1 U5732 ( .A1(n4404), .A2(n7790), .ZN(n4599) );
  NAND2_X1 U5733 ( .A1(n8736), .A2(n4605), .ZN(n4604) );
  NOR2_X1 U5734 ( .A1(n8717), .A2(n4606), .ZN(n4605) );
  INV_X1 U5735 ( .A(n8472), .ZN(n4606) );
  NAND2_X1 U5736 ( .A1(n4604), .A2(n4601), .ZN(n4600) );
  NOR2_X1 U5737 ( .A1(n4759), .A2(n4602), .ZN(n4601) );
  NAND2_X1 U5738 ( .A1(n4404), .A2(n8935), .ZN(n4602) );
  NAND2_X1 U5739 ( .A1(n8284), .A2(n8476), .ZN(n5140) );
  AND2_X1 U5740 ( .A1(n7113), .A2(n7258), .ZN(n7269) );
  NOR2_X1 U5741 ( .A1(n7112), .A2(n6099), .ZN(n7113) );
  INV_X1 U5742 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5258) );
  NAND2_X1 U5743 ( .A1(n5352), .A2(n5531), .ZN(n4677) );
  INV_X1 U5744 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5353) );
  INV_X1 U5745 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n10377) );
  AND2_X1 U5746 ( .A1(n6787), .A2(n5189), .ZN(n5188) );
  NAND2_X1 U5747 ( .A1(n4403), .A2(n4986), .ZN(n4615) );
  NAND2_X1 U5748 ( .A1(n5187), .A2(n9447), .ZN(n5182) );
  INV_X1 U5749 ( .A(n5328), .ZN(n5187) );
  INV_X1 U5750 ( .A(n8044), .ZN(n4985) );
  NOR2_X1 U5751 ( .A1(n8046), .A2(n9548), .ZN(n4984) );
  NAND2_X1 U5752 ( .A1(n8089), .A2(n8088), .ZN(n9414) );
  NOR2_X1 U5753 ( .A1(n7153), .A2(n5005), .ZN(n7592) );
  AND2_X1 U5754 ( .A1(n7800), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5005) );
  INV_X1 U5755 ( .A(n9915), .ZN(n4998) );
  AOI21_X1 U5756 ( .B1(n4999), .B2(n4503), .A(n4997), .ZN(n4996) );
  INV_X1 U5757 ( .A(n9916), .ZN(n4997) );
  NAND2_X1 U5758 ( .A1(n4996), .A2(n4993), .ZN(n4992) );
  NAND2_X1 U5759 ( .A1(n10413), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n4993) );
  NAND2_X1 U5760 ( .A1(n5072), .A2(n9665), .ZN(n5071) );
  INV_X1 U5761 ( .A(n9774), .ZN(n5072) );
  NOR3_X1 U5762 ( .A1(n7903), .A2(n9519), .A3(n9420), .ZN(n4541) );
  OR2_X1 U5763 ( .A1(n5048), .A2(n10055), .ZN(n9746) );
  NAND2_X1 U5764 ( .A1(n4545), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n7871) );
  AOI21_X1 U5765 ( .B1(n5289), .B2(n5290), .A(n4480), .ZN(n4646) );
  NAND2_X1 U5766 ( .A1(n9581), .A2(n9737), .ZN(n5078) );
  INV_X1 U5767 ( .A(n9737), .ZN(n5076) );
  INV_X1 U5768 ( .A(n4545), .ZN(n7852) );
  INV_X1 U5769 ( .A(n4438), .ZN(n5298) );
  INV_X1 U5770 ( .A(n10154), .ZN(n5296) );
  NOR2_X1 U5771 ( .A1(n7812), .A2(n7811), .ZN(n4543) );
  NOR2_X1 U5772 ( .A1(n7348), .A2(n4842), .ZN(n4841) );
  INV_X1 U5773 ( .A(n7235), .ZN(n4842) );
  NOR2_X1 U5774 ( .A1(n5056), .A2(n10303), .ZN(n5055) );
  OR2_X1 U5775 ( .A1(n7366), .A2(n9624), .ZN(n9620) );
  INV_X1 U5776 ( .A(n7236), .ZN(n4844) );
  NAND2_X1 U5777 ( .A1(n10473), .A2(n5061), .ZN(n5059) );
  NOR2_X1 U5778 ( .A1(n5281), .A2(n4434), .ZN(n5280) );
  INV_X1 U5779 ( .A(n9699), .ZN(n5278) );
  NOR2_X1 U5780 ( .A1(n6998), .A2(n4434), .ZN(n5276) );
  INV_X1 U5781 ( .A(n7721), .ZN(n9789) );
  OR2_X1 U5782 ( .A1(n6402), .A2(n6330), .ZN(n6387) );
  NAND2_X1 U5783 ( .A1(n6386), .A2(n7007), .ZN(n6402) );
  NAND2_X1 U5784 ( .A1(n5043), .A2(n4525), .ZN(n4524) );
  AND2_X1 U5785 ( .A1(n5045), .A2(n5044), .ZN(n5043) );
  NAND2_X1 U5786 ( .A1(n7832), .A2(n9677), .ZN(n4644) );
  NAND2_X1 U5787 ( .A1(n5058), .A2(n5060), .ZN(n5316) );
  NOR2_X1 U5788 ( .A1(n9590), .A2(n5059), .ZN(n5058) );
  INV_X1 U5789 ( .A(n6721), .ZN(n6720) );
  NAND2_X1 U5790 ( .A1(n10447), .A2(n6705), .ZN(n6946) );
  INV_X1 U5791 ( .A(n6054), .ZN(n5062) );
  AND2_X1 U5792 ( .A1(n7712), .A2(n5982), .ZN(n7710) );
  AND2_X1 U5793 ( .A1(n5977), .A2(n5959), .ZN(n5975) );
  NAND2_X1 U5794 ( .A1(n4955), .A2(n4958), .ZN(n5492) );
  AOI21_X1 U5795 ( .B1(n4960), .B2(n5486), .A(n4959), .ZN(n4958) );
  AOI21_X1 U5796 ( .B1(n5162), .B2(n5164), .A(n5159), .ZN(n5158) );
  INV_X1 U5797 ( .A(n5479), .ZN(n5159) );
  NAND2_X1 U5798 ( .A1(n4620), .A2(n6306), .ZN(n4619) );
  NAND2_X1 U5799 ( .A1(n4621), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4620) );
  INV_X1 U5800 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n4902) );
  INV_X1 U5801 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n6049) );
  NAND2_X1 U5802 ( .A1(n5457), .A2(n5456), .ZN(n5774) );
  AOI21_X1 U5803 ( .B1(n5151), .B2(n5153), .A(n5148), .ZN(n5147) );
  INV_X1 U5804 ( .A(n5448), .ZN(n5148) );
  NAND2_X1 U5805 ( .A1(n5436), .A2(n5151), .ZN(n5149) );
  INV_X1 U5806 ( .A(n5435), .ZN(n5155) );
  INV_X1 U5807 ( .A(n4670), .ZN(n4669) );
  OAI21_X1 U5808 ( .B1(n4672), .B2(n4671), .A(n5319), .ZN(n4670) );
  INV_X1 U5809 ( .A(n5651), .ZN(n4671) );
  NOR2_X1 U5810 ( .A1(n6163), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n4744) );
  NOR2_X1 U5811 ( .A1(n6155), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n6161) );
  OR2_X1 U5812 ( .A1(n6150), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n6155) );
  OAI21_X1 U5813 ( .B1(n4394), .B2(P1_DATAO_REG_2__SCAN_IN), .A(SI_2_), .ZN(
        n4748) );
  NAND2_X1 U5814 ( .A1(n4724), .A2(n4424), .ZN(n8151) );
  INV_X1 U5815 ( .A(n8154), .ZN(n4783) );
  AND2_X1 U5816 ( .A1(n5524), .A2(n5517), .ZN(n6613) );
  NAND2_X1 U5817 ( .A1(n5876), .A2(n5877), .ZN(n5100) );
  OR2_X1 U5818 ( .A1(n6114), .A2(n6115), .ZN(n6900) );
  XNOR2_X1 U5819 ( .A(n7272), .B(n5985), .ZN(n6898) );
  NAND2_X1 U5820 ( .A1(n8151), .A2(n5773), .ZN(n8200) );
  INV_X1 U5821 ( .A(n5900), .ZN(n8288) );
  AND4_X2 U5822 ( .A1(n5530), .A2(n5529), .A3(n5528), .A4(n5527), .ZN(n6081)
         );
  NAND2_X1 U5823 ( .A1(n5640), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5527) );
  OR2_X1 U5824 ( .A1(n5545), .A2(n6837), .ZN(n5528) );
  NAND2_X1 U5825 ( .A1(n8652), .A2(n8653), .ZN(n8651) );
  NAND2_X1 U5826 ( .A1(n8651), .A2(n4762), .ZN(n6915) );
  OR2_X1 U5827 ( .A1(n8660), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4762) );
  NOR2_X1 U5828 ( .A1(n6913), .A2(n4812), .ZN(n6859) );
  AND2_X1 U5829 ( .A1(n6918), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4812) );
  NAND2_X1 U5830 ( .A1(n4566), .A2(n5784), .ZN(n4565) );
  NAND2_X1 U5831 ( .A1(n7010), .A2(n7503), .ZN(n4566) );
  NAND2_X1 U5832 ( .A1(n7668), .A2(n7669), .ZN(n8666) );
  NOR2_X1 U5833 ( .A1(n8702), .A2(n8694), .ZN(n8693) );
  NAND2_X1 U5834 ( .A1(n8720), .A2(n4583), .ZN(n8702) );
  NOR2_X1 U5835 ( .A1(n8978), .A2(n8971), .ZN(n4583) );
  NAND2_X1 U5836 ( .A1(n8720), .A2(n7779), .ZN(n8700) );
  AND2_X1 U5837 ( .A1(n8806), .A2(n5266), .ZN(n8720) );
  NOR2_X1 U5838 ( .A1(n8984), .A2(n5267), .ZN(n5266) );
  INV_X1 U5839 ( .A(n5268), .ZN(n5267) );
  AND2_X1 U5840 ( .A1(n8806), .A2(n5268), .ZN(n8748) );
  NAND2_X1 U5841 ( .A1(n5144), .A2(n8463), .ZN(n8737) );
  AND2_X1 U5842 ( .A1(n5963), .A2(n5946), .ZN(n8762) );
  NAND2_X1 U5843 ( .A1(n8806), .A2(n5270), .ZN(n8760) );
  AND2_X1 U5844 ( .A1(n8804), .A2(n8811), .ZN(n8806) );
  NAND2_X1 U5845 ( .A1(n8806), .A2(n8782), .ZN(n8776) );
  OR2_X1 U5846 ( .A1(n9010), .A2(n8453), .ZN(n8794) );
  AND2_X1 U5847 ( .A1(n9015), .A2(n8850), .ZN(n8823) );
  AND2_X1 U5848 ( .A1(n5927), .A2(n5926), .ZN(n8824) );
  AND2_X1 U5849 ( .A1(n8833), .A2(n8820), .ZN(n8804) );
  AND2_X1 U5850 ( .A1(n8434), .A2(n8443), .ZN(n8839) );
  NAND2_X1 U5851 ( .A1(n8863), .A2(n4940), .ZN(n4936) );
  AND2_X1 U5852 ( .A1(n5883), .A2(n5894), .ZN(n8834) );
  INV_X1 U5853 ( .A(n8839), .ZN(n8831) );
  NAND2_X1 U5854 ( .A1(n5224), .A2(n4784), .ZN(n4922) );
  AOI21_X1 U5855 ( .B1(n5224), .B2(n5227), .A(n5223), .ZN(n5222) );
  INV_X1 U5856 ( .A(n7762), .ZN(n4784) );
  NAND2_X1 U5857 ( .A1(n4777), .A2(n4776), .ZN(n4775) );
  INV_X1 U5858 ( .A(n5260), .ZN(n4777) );
  NAND2_X1 U5859 ( .A1(n8863), .A2(n8864), .ZN(n8862) );
  OR2_X1 U5860 ( .A1(n9037), .A2(n8942), .ZN(n5261) );
  NOR2_X1 U5861 ( .A1(n5322), .A2(n8942), .ZN(n8936) );
  NAND2_X1 U5862 ( .A1(n7781), .A2(n7780), .ZN(n8923) );
  NOR2_X1 U5863 ( .A1(n4573), .A2(n9054), .ZN(n4571) );
  NAND2_X1 U5864 ( .A1(n4945), .A2(n4943), .ZN(n4942) );
  NOR2_X1 U5865 ( .A1(n5127), .A2(n8411), .ZN(n5123) );
  INV_X1 U5866 ( .A(n4945), .ZN(n4944) );
  NAND2_X1 U5867 ( .A1(n4941), .A2(n4945), .ZN(n5124) );
  NAND2_X1 U5868 ( .A1(n7630), .A2(n8399), .ZN(n4941) );
  INV_X1 U5869 ( .A(n5127), .ZN(n5126) );
  INV_X1 U5870 ( .A(n5216), .ZN(n4767) );
  NOR2_X1 U5871 ( .A1(n5327), .A2(n4573), .ZN(n7686) );
  AND4_X1 U5872 ( .A1(n5767), .A2(n5766), .A3(n5765), .A4(n5764), .ZN(n7700)
         );
  NAND2_X1 U5873 ( .A1(n5125), .A2(n8402), .ZN(n7681) );
  OR2_X1 U5874 ( .A1(n7661), .A2(n7631), .ZN(n5125) );
  NOR2_X1 U5875 ( .A1(n5327), .A2(n9067), .ZN(n7635) );
  NAND2_X1 U5876 ( .A1(n5146), .A2(n8389), .ZN(n7580) );
  INV_X1 U5877 ( .A(n8324), .ZN(n7492) );
  AND2_X1 U5878 ( .A1(n5262), .A2(n5265), .ZN(n7578) );
  NOR2_X1 U5879 ( .A1(n5263), .A2(n7567), .ZN(n5262) );
  NAND2_X1 U5880 ( .A1(n5265), .A2(n5264), .ZN(n7487) );
  AND4_X1 U5881 ( .A1(n5648), .A2(n5647), .A3(n5646), .A4(n5645), .ZN(n7493)
         );
  NAND2_X1 U5882 ( .A1(n5265), .A2(n7291), .ZN(n7448) );
  NAND2_X1 U5883 ( .A1(n8527), .A2(n6099), .ZN(n6100) );
  INV_X1 U5884 ( .A(n9137), .ZN(n5589) );
  NAND3_X1 U5885 ( .A1(n5253), .A2(n5254), .A3(n6094), .ZN(n7112) );
  NAND2_X1 U5886 ( .A1(n5640), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5547) );
  NAND2_X1 U5887 ( .A1(n5037), .A2(n5036), .ZN(n5548) );
  NAND2_X1 U5888 ( .A1(n5254), .A2(n5253), .ZN(n7092) );
  NAND2_X1 U5889 ( .A1(n6733), .A2(n6089), .ZN(n6732) );
  NOR2_X1 U5890 ( .A1(n8950), .A2(n7050), .ZN(n7093) );
  INV_X1 U5891 ( .A(n4597), .ZN(n8981) );
  OAI211_X1 U5892 ( .C1(n4604), .C2(n4603), .A(n4600), .B(n4598), .ZN(n4597)
         );
  AOI21_X1 U5893 ( .B1(n4759), .B2(n4599), .A(n4760), .ZN(n4598) );
  NAND2_X1 U5894 ( .A1(n4759), .A2(n8935), .ZN(n4603) );
  INV_X1 U5895 ( .A(n5239), .ZN(n5235) );
  AND2_X1 U5896 ( .A1(n5233), .A2(n4772), .ZN(n4771) );
  OR2_X1 U5897 ( .A1(n5239), .A2(n4759), .ZN(n5233) );
  NOR2_X1 U5898 ( .A1(n4420), .A2(n8711), .ZN(n4772) );
  INV_X1 U5899 ( .A(n6094), .ZN(n7038) );
  INV_X1 U5900 ( .A(n10530), .ZN(n9075) );
  INV_X1 U5901 ( .A(n6107), .ZN(n6490) );
  NAND2_X1 U5902 ( .A1(n6815), .A2(n10514), .ZN(n10501) );
  NAND2_X1 U5903 ( .A1(n4723), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4766) );
  NAND2_X1 U5904 ( .A1(n5496), .A2(n5495), .ZN(n8687) );
  AND2_X1 U5905 ( .A1(n4723), .A2(n4494), .ZN(n5495) );
  NAND2_X1 U5906 ( .A1(n6011), .A2(n5494), .ZN(n5496) );
  NAND2_X1 U5907 ( .A1(n5999), .A2(n5255), .ZN(n6011) );
  INV_X1 U5908 ( .A(n5257), .ZN(n5255) );
  NAND2_X1 U5909 ( .A1(n5107), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6005) );
  AND2_X1 U5910 ( .A1(n5369), .A2(n5382), .ZN(n5108) );
  INV_X1 U5911 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6004) );
  OR3_X1 U5912 ( .A1(n5792), .A2(P2_IR_REG_13__SCAN_IN), .A3(n5791), .ZN(n5794) );
  INV_X1 U5913 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7185) );
  NAND2_X1 U5914 ( .A1(n6350), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7394) );
  INV_X1 U5915 ( .A(n7370), .ZN(n6350) );
  INV_X1 U5916 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7393) );
  AND2_X1 U5917 ( .A1(n8087), .A2(n8086), .ZN(n8095) );
  OR2_X1 U5918 ( .A1(n7533), .A2(n7534), .ZN(n4987) );
  OAI22_X1 U5919 ( .A1(n6655), .A2(n8127), .B1(n10447), .B2(n8121), .ZN(n6388)
         );
  OR2_X1 U5920 ( .A1(n6380), .A2(n6546), .ZN(n6450) );
  OR2_X1 U5921 ( .A1(n9680), .A2(n6448), .ZN(n6452) );
  NAND2_X1 U5922 ( .A1(n6749), .A2(n6748), .ZN(n5192) );
  OAI21_X1 U5923 ( .B1(n4535), .B2(n9687), .A(n9784), .ZN(n4534) );
  NAND2_X1 U5924 ( .A1(n9675), .A2(n10208), .ZN(n4535) );
  INV_X1 U5925 ( .A(n9826), .ZN(n4532) );
  NOR2_X1 U5926 ( .A1(n9789), .A2(n9690), .ZN(n4531) );
  AND2_X1 U5927 ( .A1(n9651), .A2(n9985), .ZN(n9819) );
  NAND2_X1 U5928 ( .A1(n4537), .A2(n9686), .ZN(n9793) );
  AND4_X1 U5929 ( .A1(n7365), .A2(n7364), .A3(n7363), .A4(n7362), .ZN(n7532)
         );
  OR2_X1 U5930 ( .A1(n9570), .A2(n6512), .ZN(n6516) );
  INV_X1 U5931 ( .A(n5272), .ZN(n5271) );
  OAI22_X1 U5932 ( .A1(n6593), .A2(n6411), .B1(n6472), .B2(n6410), .ZN(n5272)
         );
  NAND2_X1 U5933 ( .A1(n6279), .A2(n4898), .ZN(n4900) );
  NAND2_X1 U5934 ( .A1(n7720), .A2(n4899), .ZN(n4901) );
  AND2_X1 U5935 ( .A1(n4749), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n4898) );
  AND2_X1 U5936 ( .A1(n6253), .A2(n6206), .ZN(n6207) );
  NAND2_X1 U5937 ( .A1(n6247), .A2(n6246), .ZN(n6422) );
  NAND2_X1 U5938 ( .A1(n4744), .A2(n4743), .ZN(n6193) );
  INV_X1 U5939 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n4743) );
  NAND2_X1 U5940 ( .A1(n6425), .A2(n6424), .ZN(n9878) );
  NAND2_X1 U5941 ( .A1(n4446), .A2(n5008), .ZN(n5007) );
  INV_X1 U5942 ( .A(n5012), .ZN(n5008) );
  OR2_X1 U5943 ( .A1(n7594), .A2(n7593), .ZN(n5004) );
  NOR2_X1 U5944 ( .A1(n9900), .A2(n4502), .ZN(n9903) );
  AND2_X1 U5945 ( .A1(n7960), .A2(n7959), .ZN(n8138) );
  NOR2_X1 U5946 ( .A1(n10211), .A2(n10169), .ZN(n4713) );
  INV_X1 U5947 ( .A(n9965), .ZN(n7994) );
  AND2_X1 U5948 ( .A1(n7967), .A2(n7943), .ZN(n9982) );
  NAND2_X1 U5949 ( .A1(n7928), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n7942) );
  INV_X1 U5950 ( .A(n7930), .ZN(n7928) );
  OR2_X1 U5951 ( .A1(n10006), .A2(n6593), .ZN(n7922) );
  XNOR2_X1 U5952 ( .A(n9995), .B(n9996), .ZN(n4753) );
  NAND2_X1 U5953 ( .A1(n4541), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n7930) );
  NAND2_X1 U5954 ( .A1(n10081), .A2(n5045), .ZN(n10031) );
  NAND2_X1 U5955 ( .A1(n9768), .A2(n9655), .ZN(n10047) );
  AOI21_X1 U5956 ( .B1(n4849), .B2(n4851), .A(n4468), .ZN(n4846) );
  AOI21_X1 U5957 ( .B1(n4445), .B2(n5068), .A(n5065), .ZN(n5064) );
  INV_X1 U5958 ( .A(n9766), .ZN(n5065) );
  NAND2_X1 U5959 ( .A1(n10081), .A2(n10071), .ZN(n10066) );
  NOR2_X1 U5960 ( .A1(n10080), .A2(n10265), .ZN(n10081) );
  NOR2_X1 U5961 ( .A1(n10124), .A2(n10275), .ZN(n10108) );
  NAND2_X1 U5962 ( .A1(n4543), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n7836) );
  OR2_X1 U5963 ( .A1(n10123), .A2(n10282), .ZN(n10124) );
  NAND2_X1 U5964 ( .A1(n4717), .A2(n9633), .ZN(n10137) );
  INV_X1 U5965 ( .A(n10162), .ZN(n4718) );
  AND3_X1 U5966 ( .A1(n7840), .A2(n7839), .A3(n7838), .ZN(n10139) );
  OR2_X1 U5967 ( .A1(n7394), .A2(n7393), .ZN(n7812) );
  INV_X1 U5968 ( .A(n4543), .ZN(n7823) );
  AND2_X1 U5969 ( .A1(n4411), .A2(n4761), .ZN(n10155) );
  AND2_X1 U5970 ( .A1(n7439), .A2(n10156), .ZN(n4761) );
  NAND2_X1 U5971 ( .A1(n7439), .A2(n4411), .ZN(n10174) );
  NAND2_X1 U5972 ( .A1(n7439), .A2(n5055), .ZN(n10176) );
  OR2_X1 U5973 ( .A1(n5056), .A2(n7532), .ZN(n7981) );
  NAND2_X1 U5974 ( .A1(n5287), .A2(n5286), .ZN(n7426) );
  INV_X1 U5975 ( .A(n9710), .ZN(n5286) );
  NAND2_X1 U5976 ( .A1(n4528), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7370) );
  INV_X1 U5977 ( .A(n7359), .ZN(n4528) );
  INV_X1 U5978 ( .A(n9620), .ZN(n9711) );
  NAND2_X1 U5979 ( .A1(n4529), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7359) );
  INV_X1 U5980 ( .A(n7210), .ZN(n4529) );
  NOR2_X1 U5981 ( .A1(n5316), .A2(n7184), .ZN(n7438) );
  AND2_X1 U5982 ( .A1(n9612), .A2(n7427), .ZN(n9708) );
  NAND2_X1 U5983 ( .A1(n6349), .A2(n4473), .ZN(n6804) );
  NAND2_X1 U5984 ( .A1(n4542), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7186) );
  INV_X1 U5985 ( .A(n6804), .ZN(n4542) );
  NAND2_X1 U5986 ( .A1(n5060), .A2(n5057), .ZN(n7278) );
  INV_X1 U5987 ( .A(n5059), .ZN(n5057) );
  NAND2_X1 U5988 ( .A1(n5060), .A2(n6990), .ZN(n7226) );
  NOR2_X1 U5989 ( .A1(n7126), .A2(n4522), .ZN(n7225) );
  NAND3_X1 U5990 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n6766) );
  AND4_X1 U5991 ( .A1(n5042), .A2(n6383), .A3(n6705), .A4(n5041), .ZN(n6948)
         );
  AND2_X1 U5992 ( .A1(n6452), .A2(n6451), .ZN(n5041) );
  AND3_X1 U5993 ( .A1(n6384), .A2(n6385), .A3(n6450), .ZN(n5042) );
  NAND2_X1 U5994 ( .A1(n6948), .A2(n6660), .ZN(n6721) );
  INV_X1 U5995 ( .A(n9697), .ZN(n6952) );
  AND2_X1 U5996 ( .A1(n9801), .A2(n9799), .ZN(n6951) );
  AND2_X1 U5997 ( .A1(n10205), .A2(n10476), .ZN(n10206) );
  NAND2_X1 U5998 ( .A1(n10220), .A2(n5320), .ZN(n4833) );
  NAND2_X1 U5999 ( .A1(n7802), .A2(n7801), .ZN(n10295) );
  NAND2_X1 U6000 ( .A1(n4837), .A2(n4839), .ZN(n4836) );
  INV_X1 U6001 ( .A(n9707), .ZN(n4839) );
  INV_X1 U6002 ( .A(n10458), .ZN(n10464) );
  INV_X1 U6003 ( .A(n7796), .ZN(n6705) );
  NOR2_X1 U6004 ( .A1(n6677), .A2(n6676), .ZN(n6630) );
  OR2_X1 U6005 ( .A1(n10458), .A2(n10059), .ZN(n6324) );
  XNOR2_X1 U6006 ( .A(n4963), .B(n8306), .ZN(n9560) );
  XNOR2_X1 U6007 ( .A(n8013), .B(n8012), .ZN(n9563) );
  NAND2_X1 U6008 ( .A1(n8300), .A2(n8299), .ZN(n8013) );
  NAND2_X1 U6009 ( .A1(n6075), .A2(n5312), .ZN(n4879) );
  XNOR2_X1 U6010 ( .A(n8011), .B(n7719), .ZN(n9678) );
  XNOR2_X1 U6011 ( .A(n7725), .B(n7724), .ZN(n8006) );
  NAND2_X1 U6012 ( .A1(n4695), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4694) );
  XNOR2_X1 U6013 ( .A(n7711), .B(n7710), .ZN(n9114) );
  XNOR2_X1 U6014 ( .A(n5976), .B(n5975), .ZN(n9117) );
  NAND2_X1 U6015 ( .A1(n6073), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6058) );
  INV_X1 U6016 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6059) );
  NAND2_X1 U6017 ( .A1(n4962), .A2(n5481), .ZN(n5891) );
  NAND2_X1 U6018 ( .A1(n5274), .A2(n5207), .ZN(n5210) );
  AND2_X1 U6019 ( .A1(n5211), .A2(n6064), .ZN(n5207) );
  AND2_X1 U6020 ( .A1(n6066), .A2(n5208), .ZN(n5211) );
  NAND2_X1 U6021 ( .A1(n5161), .A2(n5474), .ZN(n5869) );
  NAND2_X1 U6022 ( .A1(n5470), .A2(n5165), .ZN(n5161) );
  OAI21_X1 U6023 ( .B1(n5775), .B2(n5174), .A(n5171), .ZN(n5819) );
  XNOR2_X1 U6024 ( .A(n5752), .B(n5751), .ZN(n7804) );
  NAND2_X1 U6025 ( .A1(n5149), .A2(n5147), .ZN(n5752) );
  NAND2_X1 U6026 ( .A1(n5436), .A2(n5435), .ZN(n4770) );
  INV_X1 U6027 ( .A(n4744), .ZN(n6178) );
  NAND2_X1 U6028 ( .A1(n5635), .A2(n5634), .ZN(n5650) );
  XNOR2_X1 U6029 ( .A(n5602), .B(n4640), .ZN(n6773) );
  INV_X1 U6030 ( .A(n5412), .ZN(n4640) );
  NAND2_X1 U6031 ( .A1(n5215), .A2(n5411), .ZN(n5602) );
  XNOR2_X1 U6032 ( .A(n5406), .B(SI_4_), .ZN(n5558) );
  OAI21_X1 U6033 ( .B1(n6127), .B2(n4551), .A(n4549), .ZN(n6129) );
  NAND2_X1 U6034 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n4551) );
  XNOR2_X1 U6035 ( .A(n5402), .B(SI_3_), .ZN(n5551) );
  OR2_X1 U6036 ( .A1(n6124), .A2(n10343), .ZN(n6149) );
  AND2_X1 U6037 ( .A1(n4638), .A2(n4637), .ZN(n10383) );
  INV_X1 U6038 ( .A(n10578), .ZN(n4637) );
  OR2_X1 U6039 ( .A1(n10579), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n4638) );
  NAND2_X1 U6040 ( .A1(n4632), .A2(n10387), .ZN(n10388) );
  NAND2_X1 U6041 ( .A1(n10575), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n4632) );
  NAND2_X1 U6042 ( .A1(n4724), .A2(n5750), .ZN(n8153) );
  INV_X1 U6043 ( .A(n4794), .ZN(n8163) );
  NOR2_X1 U6044 ( .A1(n5665), .A2(n5317), .ZN(n5666) );
  NAND2_X1 U6045 ( .A1(n4757), .A2(n5680), .ZN(n7645) );
  NAND2_X1 U6046 ( .A1(n7349), .A2(n8307), .ZN(n4757) );
  OAI21_X1 U6047 ( .B1(n6621), .B2(n6620), .A(n5543), .ZN(n6639) );
  NAND2_X1 U6048 ( .A1(n5091), .A2(n5848), .ZN(n8171) );
  AND4_X1 U6049 ( .A1(n5662), .A2(n5661), .A3(n5660), .A4(n5659), .ZN(n7582)
         );
  OR2_X1 U6050 ( .A1(n5896), .A2(n7045), .ZN(n5519) );
  NAND2_X1 U6051 ( .A1(n6613), .A2(n6612), .ZN(n5083) );
  NAND2_X1 U6052 ( .A1(n5101), .A2(n5100), .ZN(n8180) );
  OR2_X1 U6053 ( .A1(n8233), .A2(n8232), .ZN(n5101) );
  INV_X1 U6054 ( .A(n5086), .ZN(n7331) );
  AOI21_X1 U6055 ( .B1(n7138), .B2(n7139), .A(n5089), .ZN(n5086) );
  NAND2_X1 U6056 ( .A1(n5943), .A2(n5942), .ZN(n8996) );
  AND4_X1 U6057 ( .A1(n5788), .A2(n5787), .A3(n5786), .A4(n5785), .ZN(n8925)
         );
  NAND2_X1 U6058 ( .A1(n8204), .A2(n5817), .ZN(n8213) );
  CLKBUF_X1 U6059 ( .A(n6644), .Z(n6648) );
  AND4_X1 U6060 ( .A1(n5687), .A2(n5686), .A3(n5685), .A4(n5684), .ZN(n7554)
         );
  AND4_X1 U6061 ( .A1(n5731), .A2(n5730), .A3(n5729), .A4(n5728), .ZN(n7626)
         );
  NAND2_X1 U6062 ( .A1(n5833), .A2(n5832), .ZN(n8251) );
  NOR2_X1 U6063 ( .A1(n8212), .A2(n4726), .ZN(n4725) );
  AND2_X1 U6064 ( .A1(n8260), .A2(n4730), .ZN(n4729) );
  NAND2_X1 U6065 ( .A1(n4727), .A2(n4732), .ZN(n8261) );
  OR2_X1 U6066 ( .A1(n8191), .A2(n4728), .ZN(n4727) );
  INV_X1 U6067 ( .A(n4730), .ZN(n4728) );
  AND3_X1 U6068 ( .A1(n5808), .A2(n5807), .A3(n5806), .ZN(n8278) );
  NAND2_X1 U6069 ( .A1(n8227), .A2(n8888), .ZN(n8277) );
  INV_X1 U6070 ( .A(n8501), .ZN(n5113) );
  NAND2_X1 U6071 ( .A1(n5141), .A2(n8293), .ZN(n8297) );
  NAND2_X1 U6072 ( .A1(n5115), .A2(n8501), .ZN(n5114) );
  NAND2_X1 U6073 ( .A1(n5116), .A2(n5119), .ZN(n5115) );
  INV_X1 U6074 ( .A(n5120), .ZN(n5119) );
  NOR2_X1 U6075 ( .A1(n8313), .A2(n8506), .ZN(n4967) );
  INV_X1 U6076 ( .A(n8156), .ZN(n8518) );
  NAND4_X1 U6077 ( .A1(n5612), .A2(n5611), .A3(n5610), .A4(n5609), .ZN(n8525)
         );
  INV_X1 U6078 ( .A(n8316), .ZN(n8527) );
  INV_X1 U6079 ( .A(n6090), .ZN(n8528) );
  NAND2_X1 U6080 ( .A1(n8570), .A2(n8569), .ZN(n6845) );
  NAND2_X1 U6081 ( .A1(n6855), .A2(n6854), .ZN(n8639) );
  OAI21_X1 U6082 ( .B1(n6855), .B2(n4559), .A(n4557), .ZN(n8641) );
  OAI21_X1 U6083 ( .B1(n4557), .B2(n4556), .A(n4555), .ZN(n4554) );
  NOR3_X1 U6084 ( .A1(n6855), .A2(n4559), .A3(n4556), .ZN(n4553) );
  INV_X1 U6085 ( .A(n6922), .ZN(n4556) );
  OR2_X1 U6086 ( .A1(n6910), .A2(n6911), .ZN(n6908) );
  NOR2_X1 U6087 ( .A1(n4565), .A2(n7508), .ZN(n7507) );
  XNOR2_X1 U6088 ( .A(n8666), .B(n4764), .ZN(n7670) );
  INV_X1 U6089 ( .A(n8681), .ZN(n8654) );
  NAND2_X1 U6090 ( .A1(n8685), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4570) );
  INV_X1 U6091 ( .A(n8684), .ZN(n4569) );
  NAND2_X1 U6092 ( .A1(n8736), .A2(n8472), .ZN(n8726) );
  NAND2_X1 U6093 ( .A1(n8735), .A2(n7772), .ZN(n8718) );
  OAI21_X1 U6094 ( .B1(n8733), .B2(n4686), .A(n4684), .ZN(n8716) );
  NAND2_X1 U6095 ( .A1(n4585), .A2(n4584), .ZN(n8766) );
  INV_X1 U6096 ( .A(n4586), .ZN(n4585) );
  NAND2_X1 U6097 ( .A1(n8783), .A2(n8775), .ZN(n8786) );
  NAND2_X1 U6098 ( .A1(n8802), .A2(n7769), .ZN(n8774) );
  AND2_X1 U6099 ( .A1(n5244), .A2(n4417), .ZN(n8801) );
  NAND2_X1 U6100 ( .A1(n7768), .A2(n7767), .ZN(n8815) );
  NAND2_X1 U6101 ( .A1(n5232), .A2(n5230), .ZN(n8874) );
  INV_X1 U6102 ( .A(n5231), .ZN(n5230) );
  OR2_X1 U6103 ( .A1(n8880), .A2(n7763), .ZN(n5232) );
  NAND2_X1 U6104 ( .A1(n7760), .A2(n7759), .ZN(n8929) );
  NAND2_X1 U6105 ( .A1(n7623), .A2(n5033), .ZN(n7679) );
  INV_X1 U6106 ( .A(n7623), .ZN(n7624) );
  NAND2_X1 U6107 ( .A1(n7799), .A2(n8307), .ZN(n4607) );
  OAI21_X1 U6108 ( .B1(n7622), .B2(n7621), .A(n7620), .ZN(n7656) );
  AOI21_X2 U6109 ( .B1(n7354), .B2(n8307), .A(n5706), .ZN(n7561) );
  NAND2_X1 U6110 ( .A1(n4687), .A2(n7446), .ZN(n7485) );
  AND2_X1 U6111 ( .A1(n7446), .A2(n7295), .ZN(n7296) );
  INV_X1 U6112 ( .A(n4690), .ZN(n4687) );
  INV_X1 U6113 ( .A(n8954), .ZN(n8871) );
  NAND2_X1 U6114 ( .A1(n8940), .A2(n6108), .ZN(n8894) );
  INV_X1 U6115 ( .A(n8899), .ZN(n8953) );
  CLKBUF_X1 U6116 ( .A(n6104), .Z(n8950) );
  INV_X1 U6117 ( .A(n8894), .ZN(n8951) );
  INV_X1 U6118 ( .A(n10544), .ZN(n10542) );
  OR3_X1 U6119 ( .A1(n9026), .A2(n9025), .A3(n9024), .ZN(n9093) );
  AND2_X1 U6120 ( .A1(n6172), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10514) );
  INV_X1 U6121 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5038) );
  XNOR2_X1 U6122 ( .A(n6009), .B(n6008), .ZN(n7528) );
  INV_X1 U6123 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7722) );
  NAND2_X1 U6124 ( .A1(n4791), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5383) );
  INV_X1 U6125 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n9374) );
  INV_X1 U6126 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6743) );
  INV_X1 U6127 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6417) );
  INV_X1 U6128 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6268) );
  INV_X1 U6129 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n9294) );
  AND3_X1 U6130 ( .A1(n5531), .A2(n4792), .A3(n5344), .ZN(n4721) );
  XNOR2_X1 U6131 ( .A(n5550), .B(n5549), .ZN(n8559) );
  NAND2_X1 U6132 ( .A1(n5534), .A2(n5561), .ZN(n8546) );
  OAI22_X1 U6133 ( .A1(n4765), .A2(n5531), .B1(P2_IR_REG_2__SCAN_IN), .B2(
        P2_IR_REG_31__SCAN_IN), .ZN(n5532) );
  NAND2_X1 U6134 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4765) );
  XNOR2_X1 U6135 ( .A(n5505), .B(n5504), .ZN(n6838) );
  NOR2_X1 U6136 ( .A1(n4539), .A2(n7970), .ZN(n9966) );
  NOR2_X1 U6137 ( .A1(n8139), .A2(n6593), .ZN(n4539) );
  AOI21_X1 U6138 ( .B1(n5204), .B2(n4916), .A(n4452), .ZN(n4915) );
  INV_X1 U6139 ( .A(n4917), .ZN(n4916) );
  AND4_X1 U6140 ( .A1(n7192), .A2(n7191), .A3(n7190), .A4(n7189), .ZN(n9591)
         );
  INV_X1 U6141 ( .A(n7476), .ZN(n7471) );
  INV_X1 U6142 ( .A(n10086), .ZN(n10054) );
  OAI21_X1 U6143 ( .B1(n8120), .B2(n4452), .A(n5202), .ZN(n8149) );
  INV_X1 U6144 ( .A(n5203), .ZN(n5202) );
  OAI21_X1 U6145 ( .B1(n5204), .B2(n4452), .A(n8135), .ZN(n5203) );
  AND4_X1 U6146 ( .A1(n6796), .A2(n6795), .A3(n6794), .A4(n6793), .ZN(n7253)
         );
  INV_X1 U6147 ( .A(n4908), .ZN(n9439) );
  AOI22_X1 U6148 ( .A1(n4981), .A2(n4909), .B1(n4408), .B2(n4979), .ZN(n4908)
         );
  NOR2_X1 U6149 ( .A1(n5193), .A2(n9477), .ZN(n4909) );
  OAI21_X1 U6150 ( .B1(n4442), .B2(n9446), .A(n9447), .ZN(n9506) );
  AND2_X1 U6151 ( .A1(n7890), .A2(n7889), .ZN(n9521) );
  AND2_X1 U6152 ( .A1(n6413), .A2(n9786), .ZN(n9511) );
  INV_X1 U6153 ( .A(n9529), .ZN(n9551) );
  INV_X1 U6154 ( .A(n9511), .ZN(n9554) );
  NAND2_X1 U6155 ( .A1(n6405), .A2(n10157), .ZN(n9556) );
  OR3_X1 U6156 ( .A1(n6403), .A2(n6667), .A3(n10463), .ZN(n9558) );
  AOI21_X1 U6157 ( .B1(n4536), .B2(n4533), .A(n4530), .ZN(n9792) );
  NAND2_X1 U6158 ( .A1(n4532), .A2(n4531), .ZN(n4530) );
  NAND2_X1 U6159 ( .A1(n4534), .A2(n9688), .ZN(n4533) );
  INV_X1 U6160 ( .A(n9793), .ZN(n4536) );
  OAI21_X1 U6161 ( .B1(n6375), .B2(n5212), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n4904) );
  NAND2_X1 U6162 ( .A1(n6066), .A2(n5213), .ZN(n5212) );
  INV_X1 U6163 ( .A(n9966), .ZN(n9956) );
  NAND2_X1 U6164 ( .A1(n7909), .A2(n7908), .ZN(n10041) );
  INV_X1 U6165 ( .A(n9521), .ZN(n10074) );
  INV_X1 U6166 ( .A(n7532), .ZN(n9846) );
  OR2_X1 U6167 ( .A1(n6472), .A2(n6473), .ZN(n6474) );
  OR2_X1 U6168 ( .A1(n6472), .A2(n6332), .ZN(n6336) );
  OR2_X1 U6169 ( .A1(n7944), .A2(n6333), .ZN(n6335) );
  OR2_X1 U6170 ( .A1(n6593), .A2(n10406), .ZN(n6287) );
  AND2_X1 U6171 ( .A1(n10361), .A2(n6204), .ZN(n6552) );
  NAND2_X1 U6172 ( .A1(n6262), .A2(n6223), .ZN(n6226) );
  NAND2_X1 U6173 ( .A1(n4548), .A2(n4547), .ZN(n6241) );
  INV_X1 U6174 ( .A(n6225), .ZN(n4547) );
  INV_X1 U6175 ( .A(n6226), .ZN(n4548) );
  NAND2_X1 U6176 ( .A1(n5011), .A2(n6442), .ZN(n6568) );
  NAND2_X1 U6177 ( .A1(n9878), .A2(n5012), .ZN(n5011) );
  NAND2_X1 U6178 ( .A1(n9878), .A2(n6426), .ZN(n6443) );
  INV_X1 U6179 ( .A(n5004), .ZN(n9884) );
  AND2_X1 U6180 ( .A1(n5002), .A2(n5001), .ZN(n9900) );
  INV_X1 U6181 ( .A(n9887), .ZN(n5001) );
  INV_X1 U6182 ( .A(n5002), .ZN(n9888) );
  AOI21_X1 U6183 ( .B1(n9892), .B2(n9891), .A(n9890), .ZN(n9894) );
  AOI21_X1 U6184 ( .B1(n9920), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9919), .ZN(
        n10422) );
  NAND2_X1 U6185 ( .A1(n5000), .A2(n4999), .ZN(n10415) );
  INV_X1 U6186 ( .A(n5000), .ZN(n10412) );
  INV_X1 U6187 ( .A(n9689), .ZN(n10200) );
  INV_X1 U6188 ( .A(n9939), .ZN(n10204) );
  AOI21_X1 U6189 ( .B1(n10215), .B2(n10195), .A(n9960), .ZN(n4786) );
  INV_X1 U6190 ( .A(n5052), .ZN(n9945) );
  NAND2_X1 U6191 ( .A1(n4857), .A2(n7951), .ZN(n9963) );
  NAND2_X1 U6192 ( .A1(n7938), .A2(n4861), .ZN(n4857) );
  NAND2_X1 U6193 ( .A1(n4819), .A2(n4818), .ZN(n4817) );
  XNOR2_X1 U6194 ( .A(n9987), .B(n4821), .ZN(n4820) );
  NAND2_X1 U6195 ( .A1(n9989), .A2(n10187), .ZN(n4818) );
  INV_X1 U6196 ( .A(n10231), .ZN(n9984) );
  NAND2_X1 U6197 ( .A1(n7938), .A2(n7937), .ZN(n9977) );
  OAI21_X1 U6198 ( .B1(n10030), .B2(n4652), .A(n4406), .ZN(n9994) );
  NAND2_X1 U6199 ( .A1(n7927), .A2(n7926), .ZN(n10238) );
  NAND2_X1 U6200 ( .A1(n4752), .A2(n4750), .ZN(n10236) );
  AOI21_X1 U6201 ( .B1(n9841), .B2(n10189), .A(n4751), .ZN(n4750) );
  NAND2_X1 U6202 ( .A1(n4753), .A2(n10192), .ZN(n4752) );
  NOR2_X1 U6203 ( .A1(n10025), .A2(n10167), .ZN(n4751) );
  NAND2_X1 U6204 ( .A1(n5305), .A2(n5303), .ZN(n10003) );
  INV_X1 U6205 ( .A(n5306), .ZN(n5303) );
  NAND2_X1 U6206 ( .A1(n10030), .A2(n5308), .ZN(n5305) );
  OAI21_X1 U6207 ( .B1(n10030), .B2(n7898), .A(n7897), .ZN(n10017) );
  NAND2_X1 U6208 ( .A1(n7883), .A2(n7882), .ZN(n10256) );
  NAND2_X1 U6209 ( .A1(n4848), .A2(n4852), .ZN(n10065) );
  NAND2_X1 U6210 ( .A1(n10091), .A2(n4437), .ZN(n4848) );
  NAND2_X1 U6211 ( .A1(n5066), .A2(n9760), .ZN(n10085) );
  NAND2_X1 U6212 ( .A1(n10099), .A2(n9761), .ZN(n5066) );
  AND2_X1 U6213 ( .A1(n4853), .A2(n4855), .ZN(n10079) );
  NAND2_X1 U6214 ( .A1(n10091), .A2(n10100), .ZN(n4853) );
  NAND2_X1 U6215 ( .A1(n10154), .A2(n5292), .ZN(n5288) );
  OAI21_X1 U6216 ( .B1(n10141), .B2(n7831), .A(n4438), .ZN(n10122) );
  INV_X1 U6217 ( .A(n10285), .ZN(n10149) );
  NAND2_X1 U6218 ( .A1(n5080), .A2(n5079), .ZN(n10163) );
  NAND2_X1 U6219 ( .A1(n4401), .A2(n5081), .ZN(n10185) );
  AND2_X1 U6220 ( .A1(n5081), .A2(n9749), .ZN(n10186) );
  INV_X1 U6221 ( .A(n10295), .ZN(n10183) );
  AND2_X1 U6222 ( .A1(n4835), .A2(n4834), .ZN(n7410) );
  INV_X1 U6223 ( .A(n4837), .ZN(n4835) );
  NAND2_X1 U6224 ( .A1(n7424), .A2(n5283), .ZN(n4834) );
  NAND2_X1 U6225 ( .A1(n6747), .A2(n6746), .ZN(n7232) );
  AOI21_X1 U6226 ( .B1(n6998), .B2(n5281), .A(n4434), .ZN(n5279) );
  INV_X1 U6227 ( .A(n10457), .ZN(n7000) );
  INV_X1 U6228 ( .A(n6945), .ZN(n10452) );
  NAND2_X1 U6229 ( .A1(n10170), .A2(n6631), .ZN(n10182) );
  AND2_X1 U6230 ( .A1(n10170), .A2(n6632), .ZN(n10195) );
  INV_X1 U6231 ( .A(n10182), .ZN(n10048) );
  INV_X1 U6232 ( .A(n4798), .ZN(n4797) );
  INV_X1 U6233 ( .A(n10224), .ZN(n4800) );
  INV_X1 U6234 ( .A(n10439), .ZN(n10440) );
  AND2_X1 U6235 ( .A1(n6520), .A2(n6131), .ZN(n10443) );
  AND2_X1 U6236 ( .A1(n5312), .A2(n6277), .ZN(n5311) );
  AOI21_X1 U6237 ( .B1(n6057), .B2(n6056), .A(n10343), .ZN(n4990) );
  INV_X1 U6238 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7912) );
  INV_X1 U6239 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7900) );
  OAI21_X1 U6240 ( .B1(n4957), .B2(n4960), .A(n5486), .ZN(n5913) );
  INV_X1 U6241 ( .A(n4962), .ZN(n4957) );
  INV_X1 U6242 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7894) );
  XNOR2_X1 U6243 ( .A(n6071), .B(n6070), .ZN(n9690) );
  INV_X1 U6244 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7868) );
  INV_X1 U6245 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8005) );
  OAI21_X1 U6246 ( .B1(n6375), .B2(n4621), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6618) );
  INV_X1 U6247 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7805) );
  XNOR2_X1 U6248 ( .A(n6273), .B(n6272), .ZN(n7806) );
  XNOR2_X1 U6249 ( .A(n6270), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7800) );
  XNOR2_X1 U6250 ( .A(n6168), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7386) );
  INV_X1 U6251 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6190) );
  INV_X1 U6252 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9207) );
  NAND2_X1 U6253 ( .A1(n5694), .A2(n5651), .ZN(n5673) );
  NAND2_X1 U6254 ( .A1(n6147), .A2(n5014), .ZN(n6546) );
  NAND2_X1 U6255 ( .A1(n5015), .A2(P1_IR_REG_2__SCAN_IN), .ZN(n5014) );
  INV_X1 U6256 ( .A(n6149), .ZN(n5015) );
  XNOR2_X1 U6257 ( .A(n5511), .B(n5510), .ZN(n6379) );
  NAND2_X1 U6258 ( .A1(n4630), .A2(n10381), .ZN(n10592) );
  NAND2_X1 U6259 ( .A1(n10590), .A2(n10591), .ZN(n4630) );
  AND2_X1 U6260 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10382), .ZN(n10579) );
  XNOR2_X1 U6261 ( .A(n10383), .B(n4636), .ZN(n10577) );
  INV_X1 U6262 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n4636) );
  XNOR2_X1 U6263 ( .A(n10386), .B(n4633), .ZN(n10575) );
  INV_X1 U6264 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n4633) );
  XNOR2_X1 U6265 ( .A(n10388), .B(n4631), .ZN(n10581) );
  NOR2_X1 U6266 ( .A1(n10392), .A2(n10586), .ZN(n10573) );
  AND2_X1 U6267 ( .A1(n4635), .A2(n4634), .ZN(n10567) );
  NAND2_X1 U6268 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n4634) );
  NAND2_X1 U6269 ( .A1(n10567), .A2(n10566), .ZN(n10565) );
  OAI21_X1 U6270 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10565), .ZN(n10563) );
  OAI21_X1 U6271 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10562), .ZN(n10560) );
  OAI21_X1 U6272 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10559), .ZN(n10557) );
  NAND2_X1 U6273 ( .A1(n10557), .A2(n10558), .ZN(n10556) );
  NAND2_X1 U6274 ( .A1(n10556), .A2(n4627), .ZN(n10554) );
  NAND2_X1 U6275 ( .A1(n7013), .A2(n4628), .ZN(n4627) );
  NAND2_X1 U6276 ( .A1(n10554), .A2(n10555), .ZN(n10553) );
  NAND2_X1 U6277 ( .A1(n10553), .A2(n4626), .ZN(n10551) );
  NAND2_X1 U6278 ( .A1(n9221), .A2(n9173), .ZN(n4626) );
  OAI21_X1 U6279 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n10550), .ZN(n10583) );
  OAI21_X1 U6280 ( .B1(n8724), .B2(n8268), .A(n6045), .ZN(n6046) );
  OR2_X1 U6281 ( .A1(n7758), .A2(n7757), .ZN(n4782) );
  NAND2_X1 U6282 ( .A1(n4810), .A2(n4567), .ZN(P2_U3264) );
  AOI21_X1 U6283 ( .B1(n4809), .B2(n8915), .A(n4568), .ZN(n4567) );
  NAND2_X1 U6284 ( .A1(n8683), .A2(n8340), .ZN(n4810) );
  NAND2_X1 U6285 ( .A1(n4570), .A2(n4569), .ZN(n4568) );
  AOI21_X1 U6286 ( .B1(n4951), .B2(n8940), .A(n4949), .ZN(n4948) );
  INV_X1 U6287 ( .A(n4950), .ZN(n4949) );
  INV_X1 U6288 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n5237) );
  NAND2_X1 U6289 ( .A1(n4579), .A2(n4578), .ZN(P2_U3517) );
  NAND2_X1 U6290 ( .A1(n10537), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n4578) );
  NAND2_X1 U6291 ( .A1(n9084), .A2(n10538), .ZN(n4579) );
  NAND2_X1 U6292 ( .A1(n10537), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n4934) );
  NAND2_X1 U6293 ( .A1(n4933), .A2(n4609), .ZN(n4608) );
  OAI21_X1 U6294 ( .B1(n8976), .B2(n4611), .A(n4933), .ZN(n4610) );
  INV_X1 U6295 ( .A(n4789), .ZN(n4788) );
  NAND2_X1 U6296 ( .A1(n9932), .A2(n10059), .ZN(n4790) );
  NAND2_X1 U6297 ( .A1(n9931), .A2(n10007), .ZN(n4787) );
  NAND2_X1 U6298 ( .A1(n4655), .A2(n4653), .ZN(P1_U3552) );
  OR2_X1 U6299 ( .A1(n10499), .A2(n4654), .ZN(n4653) );
  NAND2_X1 U6300 ( .A1(n10323), .A2(n10499), .ZN(n4655) );
  INV_X1 U6301 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n4654) );
  NAND2_X1 U6302 ( .A1(n4756), .A2(n4754), .ZN(P1_U3548) );
  OR2_X1 U6303 ( .A1(n10499), .A2(n4755), .ZN(n4754) );
  INV_X1 U6304 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n4755) );
  OR2_X1 U6305 ( .A1(n10488), .A2(n4831), .ZN(n4830) );
  NAND2_X1 U6306 ( .A1(n10323), .A2(n10488), .ZN(n4832) );
  INV_X1 U6307 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n4831) );
  INV_X1 U6308 ( .A(n4635), .ZN(n10568) );
  AND2_X1 U6309 ( .A1(n7788), .A2(n4939), .ZN(n4400) );
  AND2_X1 U6310 ( .A1(n9749), .A2(n7985), .ZN(n4401) );
  AND2_X1 U6311 ( .A1(n4922), .A2(n5222), .ZN(n4402) );
  OR2_X1 U6312 ( .A1(n5184), .A2(n4414), .ZN(n4403) );
  OR2_X1 U6313 ( .A1(n8742), .A2(n8984), .ZN(n4404) );
  XNOR2_X1 U6314 ( .A(n5356), .B(n5355), .ZN(n5360) );
  NOR2_X1 U6315 ( .A1(n4461), .A2(n5196), .ZN(n5193) );
  AND2_X1 U6316 ( .A1(n9715), .A2(n5078), .ZN(n4405) );
  OR2_X1 U6317 ( .A1(n9022), .A2(n8182), .ZN(n8441) );
  NOR2_X1 U6318 ( .A1(n5229), .A2(n5226), .ZN(n5225) );
  AND2_X1 U6319 ( .A1(n5301), .A2(n5310), .ZN(n4406) );
  AND2_X1 U6320 ( .A1(n9635), .A2(n10140), .ZN(n4407) );
  NAND2_X1 U6321 ( .A1(n5195), .A2(n8056), .ZN(n4408) );
  AND2_X1 U6322 ( .A1(n5147), .A2(n5751), .ZN(n4409) );
  INV_X1 U6323 ( .A(n9760), .ZN(n5068) );
  AND2_X1 U6324 ( .A1(n4407), .A2(n4463), .ZN(n4410) );
  AND2_X1 U6325 ( .A1(n5055), .A2(n10183), .ZN(n4411) );
  OR2_X1 U6326 ( .A1(n10265), .A2(n10103), .ZN(n4412) );
  NAND2_X1 U6327 ( .A1(n4937), .A2(n5323), .ZN(n4413) );
  NAND2_X1 U6328 ( .A1(n7351), .A2(n7350), .ZN(n7352) );
  INV_X1 U6329 ( .A(n7352), .ZN(n4702) );
  INV_X1 U6330 ( .A(n5259), .ZN(n8868) );
  AND2_X1 U6331 ( .A1(n5328), .A2(n5183), .ZN(n4414) );
  AND3_X1 U6332 ( .A1(n10216), .A2(n4496), .A3(n4833), .ZN(n4415) );
  NAND2_X1 U6333 ( .A1(n7950), .A2(n7949), .ZN(n9841) );
  AND2_X1 U6334 ( .A1(n5158), .A2(n4500), .ZN(n4416) );
  OR2_X1 U6335 ( .A1(n9010), .A2(n8841), .ZN(n4417) );
  AND2_X1 U6336 ( .A1(n9703), .A2(n9702), .ZN(n4418) );
  NAND2_X1 U6337 ( .A1(n7954), .A2(n7953), .ZN(n10226) );
  AND2_X1 U6338 ( .A1(n4397), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n4419) );
  INV_X1 U6339 ( .A(n10025), .ZN(n9842) );
  AND2_X1 U6340 ( .A1(n7922), .A2(n7921), .ZN(n10025) );
  AND2_X1 U6341 ( .A1(n5018), .A2(n5315), .ZN(n4420) );
  AND2_X1 U6342 ( .A1(n4482), .A2(n4680), .ZN(n4421) );
  AND2_X1 U6343 ( .A1(n4565), .A2(n4564), .ZN(n4422) );
  NAND2_X1 U6344 ( .A1(n5132), .A2(n8421), .ZN(n4423) );
  AND2_X1 U6345 ( .A1(n4783), .A2(n5750), .ZN(n4424) );
  AND2_X1 U6346 ( .A1(n5136), .A2(n4504), .ZN(n4425) );
  NAND2_X1 U6347 ( .A1(n4479), .A2(n8441), .ZN(n4939) );
  AND2_X1 U6348 ( .A1(n7199), .A2(n7198), .ZN(n7474) );
  INV_X1 U6349 ( .A(n7474), .ZN(n4907) );
  INV_X1 U6350 ( .A(n7680), .ZN(n8406) );
  INV_X1 U6351 ( .A(n8406), .ZN(n5033) );
  AND3_X1 U6352 ( .A1(n8775), .A2(n8461), .A3(n4493), .ZN(n4426) );
  AND2_X1 U6353 ( .A1(n4650), .A2(n7951), .ZN(n4427) );
  AND2_X1 U6354 ( .A1(n5039), .A2(n5038), .ZN(n4428) );
  AND2_X1 U6355 ( .A1(n4485), .A2(n5116), .ZN(n4429) );
  NAND2_X1 U6356 ( .A1(n4572), .A2(n4571), .ZN(n7704) );
  OAI21_X1 U6357 ( .B1(n6714), .B2(n9698), .A(n5279), .ZN(n7121) );
  OR2_X1 U6358 ( .A1(n5322), .A2(n5261), .ZN(n4430) );
  NAND2_X1 U6359 ( .A1(n6720), .A2(n10457), .ZN(n7126) );
  AND2_X1 U6360 ( .A1(n4996), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n4431) );
  AND2_X1 U6361 ( .A1(n4999), .A2(n9917), .ZN(n4432) );
  NAND2_X1 U6362 ( .A1(n8901), .A2(n7761), .ZN(n8900) );
  INV_X2 U6363 ( .A(n7944), .ZN(n6466) );
  AND2_X1 U6364 ( .A1(n8199), .A2(n5809), .ZN(n4433) );
  NOR2_X1 U6365 ( .A1(n9852), .A2(n7000), .ZN(n4434) );
  INV_X1 U6366 ( .A(n5056), .ZN(n10309) );
  NAND2_X1 U6367 ( .A1(n7357), .A2(n7356), .ZN(n5056) );
  AND2_X1 U6368 ( .A1(n4901), .A2(n4900), .ZN(n4435) );
  NAND2_X1 U6369 ( .A1(n4514), .A2(n4512), .ZN(n6104) );
  AND3_X1 U6370 ( .A1(n5569), .A2(n5568), .A3(n5567), .ZN(n10523) );
  NAND2_X1 U6371 ( .A1(n5910), .A2(n5909), .ZN(n4436) );
  NAND2_X1 U6372 ( .A1(n6611), .A2(n10518), .ZN(n8352) );
  NAND2_X1 U6373 ( .A1(n5999), .A2(n5353), .ZN(n6002) );
  NOR2_X1 U6374 ( .A1(n5306), .A2(n7923), .ZN(n5304) );
  AND2_X1 U6375 ( .A1(n8466), .A2(n8462), .ZN(n8775) );
  INV_X1 U6376 ( .A(n8775), .ZN(n4587) );
  AND2_X1 U6377 ( .A1(n4412), .A2(n10100), .ZN(n4437) );
  OR2_X1 U6378 ( .A1(n10149), .A2(n10168), .ZN(n4438) );
  INV_X1 U6379 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9103) );
  AND2_X1 U6380 ( .A1(n5140), .A2(n5139), .ZN(n4439) );
  AND4_X1 U6381 ( .A1(n5503), .A2(n5502), .A3(n5501), .A4(n4693), .ZN(n6090)
         );
  AND2_X1 U6382 ( .A1(n5413), .A2(SI_6_), .ZN(n4440) );
  OR2_X1 U6383 ( .A1(n5641), .A2(n5544), .ZN(n4441) );
  AND2_X1 U6384 ( .A1(n4617), .A2(n4616), .ZN(n4442) );
  INV_X1 U6385 ( .A(n5359), .ZN(n5361) );
  AND2_X1 U6386 ( .A1(n5328), .A2(n5181), .ZN(n4443) );
  XNOR2_X1 U6387 ( .A(n5465), .B(n5464), .ZN(n5818) );
  AND2_X1 U6388 ( .A1(n4981), .A2(n4980), .ZN(n4444) );
  AND2_X1 U6389 ( .A1(n10084), .A2(n5067), .ZN(n4445) );
  NOR2_X1 U6390 ( .A1(n6569), .A2(n5010), .ZN(n4446) );
  OR2_X1 U6391 ( .A1(n8447), .A2(n8494), .ZN(n4447) );
  OR2_X1 U6392 ( .A1(n6861), .A2(n8559), .ZN(n4448) );
  INV_X1 U6393 ( .A(n8857), .ZN(n5223) );
  AND3_X1 U6394 ( .A1(n8434), .A2(n8441), .A3(n8481), .ZN(n4449) );
  INV_X1 U6395 ( .A(n9773), .ZN(n4891) );
  AND3_X1 U6396 ( .A1(n5429), .A2(n5695), .A3(n5634), .ZN(n4450) );
  NAND4_X1 U6397 ( .A1(n6772), .A2(n6771), .A3(n6770), .A4(n6769), .ZN(n9850)
         );
  INV_X1 U6398 ( .A(n9850), .ZN(n4709) );
  XOR2_X1 U6399 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n4451) );
  AND2_X1 U6400 ( .A1(n8125), .A2(n8124), .ZN(n4452) );
  NAND2_X1 U6401 ( .A1(n5221), .A2(n5224), .ZN(n8856) );
  OR2_X1 U6402 ( .A1(n10207), .A2(n7973), .ZN(n10225) );
  NAND2_X1 U6403 ( .A1(n7902), .A2(n7901), .ZN(n10248) );
  INV_X1 U6404 ( .A(n10248), .ZN(n5044) );
  AND2_X1 U6405 ( .A1(n10265), .A2(n10103), .ZN(n4453) );
  OAI21_X1 U6406 ( .B1(n8900), .B2(n5225), .A(n4402), .ZN(n8858) );
  AND4_X1 U6407 ( .A1(n6050), .A2(n6160), .A3(n6049), .A4(n6048), .ZN(n4454)
         );
  AND2_X1 U6408 ( .A1(n5095), .A2(n5096), .ZN(n4455) );
  AND3_X1 U6409 ( .A1(n8393), .A2(n8394), .A3(n8391), .ZN(n4456) );
  AND4_X1 U6410 ( .A1(n7215), .A2(n7214), .A3(n7213), .A4(n7212), .ZN(n9596)
         );
  INV_X1 U6411 ( .A(n9596), .ZN(n4701) );
  OR2_X1 U6412 ( .A1(n10240), .A2(n10299), .ZN(n4457) );
  NOR2_X1 U6413 ( .A1(n9979), .A2(n10226), .ZN(n4458) );
  OR2_X1 U6414 ( .A1(n10112), .A2(n10134), .ZN(n4459) );
  INV_X1 U6415 ( .A(n10260), .ZN(n10071) );
  NAND2_X1 U6416 ( .A1(n7870), .A2(n7869), .ZN(n10260) );
  AND2_X1 U6417 ( .A1(n4400), .A2(n8775), .ZN(n4460) );
  INV_X1 U6418 ( .A(n5194), .ZN(n9426) );
  NOR2_X1 U6419 ( .A1(n4444), .A2(n5201), .ZN(n5194) );
  AOI21_X1 U6420 ( .B1(n5184), .B2(n5182), .A(n4443), .ZN(n5180) );
  INV_X1 U6421 ( .A(n7818), .ZN(n5295) );
  NOR2_X1 U6422 ( .A1(n9497), .A2(n5199), .ZN(n4461) );
  INV_X1 U6423 ( .A(n4523), .ZN(n4526) );
  AND2_X1 U6424 ( .A1(n7289), .A2(n7444), .ZN(n4462) );
  INV_X1 U6425 ( .A(n8476), .ZN(n4759) );
  XNOR2_X1 U6426 ( .A(n5747), .B(n5748), .ZN(n7516) );
  NAND2_X1 U6427 ( .A1(n7038), .A2(n7108), .ZN(n8344) );
  INV_X1 U6428 ( .A(n8344), .ZN(n5143) );
  NAND2_X1 U6429 ( .A1(n10081), .A2(n5047), .ZN(n5049) );
  NAND3_X1 U6430 ( .A1(n9633), .A2(n9632), .A3(n9749), .ZN(n4463) );
  INV_X1 U6431 ( .A(n8984), .ZN(n8724) );
  NAND2_X1 U6432 ( .A1(n5838), .A2(n5837), .ZN(n9032) );
  AND2_X1 U6433 ( .A1(n7896), .A2(n7895), .ZN(n10035) );
  INV_X1 U6434 ( .A(n10035), .ZN(n5048) );
  AND2_X1 U6435 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_REG3_REG_11__SCAN_IN), 
        .ZN(n4464) );
  AND2_X1 U6436 ( .A1(n9022), .A2(n8866), .ZN(n4465) );
  AND2_X1 U6437 ( .A1(n6093), .A2(n7026), .ZN(n4466) );
  NAND2_X1 U6438 ( .A1(n8222), .A2(n5916), .ZN(n4467) );
  INV_X1 U6439 ( .A(n9727), .ZN(n5069) );
  INV_X1 U6440 ( .A(n5193), .ZN(n4979) );
  AND2_X1 U6441 ( .A1(n10260), .A2(n10086), .ZN(n4468) );
  INV_X1 U6442 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5213) );
  INV_X1 U6443 ( .A(n5205), .ZN(n5204) );
  NAND2_X1 U6444 ( .A1(n5206), .A2(n8119), .ZN(n5205) );
  AND2_X1 U6445 ( .A1(n6107), .A2(n8337), .ZN(n4469) );
  NOR2_X1 U6446 ( .A1(n7592), .A2(n7806), .ZN(n4470) );
  NAND3_X1 U6447 ( .A1(n8443), .A2(n8494), .A3(n8442), .ZN(n4471) );
  OR2_X1 U6448 ( .A1(n6861), .A2(n8546), .ZN(n4472) );
  AND2_X1 U6449 ( .A1(n7784), .A2(n8422), .ZN(n8903) );
  AND2_X1 U6450 ( .A1(n5331), .A2(n8421), .ZN(n8928) );
  AND2_X1 U6451 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n4473) );
  OR2_X1 U6452 ( .A1(n8109), .A2(n9490), .ZN(n4474) );
  AND2_X1 U6453 ( .A1(n4576), .A2(n5256), .ZN(n4475) );
  INV_X1 U6454 ( .A(n8056), .ZN(n5201) );
  OR2_X1 U6455 ( .A1(n8055), .A2(n8054), .ZN(n8056) );
  INV_X1 U6456 ( .A(n4986), .ZN(n4616) );
  AND2_X1 U6457 ( .A1(n8025), .A2(n8026), .ZN(n4986) );
  OR2_X1 U6458 ( .A1(n6375), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n4476) );
  INV_X1 U6459 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7209) );
  AND2_X1 U6460 ( .A1(n10282), .A2(n10115), .ZN(n4477) );
  AND2_X1 U6461 ( .A1(n8390), .A2(n8399), .ZN(n4478) );
  OR2_X1 U6462 ( .A1(n8857), .A2(n8437), .ZN(n4479) );
  NAND2_X1 U6463 ( .A1(n9682), .A2(n9681), .ZN(n10209) );
  INV_X1 U6464 ( .A(n10209), .ZN(n5156) );
  INV_X1 U6465 ( .A(n9577), .ZN(n10243) );
  AND2_X1 U6466 ( .A1(n7914), .A2(n7913), .ZN(n9577) );
  INV_X1 U6467 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6062) );
  INV_X1 U6468 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5354) );
  NOR2_X1 U6469 ( .A1(n10275), .A2(n10102), .ZN(n4480) );
  INV_X1 U6470 ( .A(n7772), .ZN(n4686) );
  OR2_X1 U6471 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n4481) );
  AND2_X1 U6472 ( .A1(n4676), .A2(n5790), .ZN(n4482) );
  INV_X1 U6473 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n10343) );
  AND2_X1 U6474 ( .A1(n5056), .A2(n9846), .ZN(n4483) );
  INV_X1 U6475 ( .A(n4544), .ZN(n7884) );
  NOR2_X1 U6476 ( .A1(n7871), .A2(n6352), .ZN(n4544) );
  OR2_X1 U6477 ( .A1(n4453), .A2(n4854), .ZN(n4484) );
  INV_X1 U6478 ( .A(n9943), .ZN(n10221) );
  NAND2_X1 U6479 ( .A1(n7963), .A2(n7962), .ZN(n9943) );
  INV_X1 U6480 ( .A(n4862), .ZN(n4861) );
  OR2_X1 U6481 ( .A1(n7952), .A2(n4863), .ZN(n4862) );
  NAND2_X1 U6482 ( .A1(n8489), .A2(n8340), .ZN(n4485) );
  NAND2_X1 U6483 ( .A1(n5651), .A2(n5427), .ZN(n5649) );
  INV_X1 U6484 ( .A(n8863), .ZN(n4516) );
  NAND2_X1 U6485 ( .A1(n5961), .A2(n5960), .ZN(n8746) );
  INV_X1 U6486 ( .A(n8746), .ZN(n5269) );
  AND2_X1 U6487 ( .A1(n8180), .A2(n8179), .ZN(n4486) );
  AND2_X1 U6488 ( .A1(n5171), .A2(n5818), .ZN(n4487) );
  NAND2_X1 U6489 ( .A1(n5410), .A2(SI_5_), .ZN(n5411) );
  AND2_X1 U6490 ( .A1(n5288), .A2(n5289), .ZN(n4488) );
  NAND2_X1 U6491 ( .A1(n7774), .A2(n8476), .ZN(n4935) );
  INV_X1 U6492 ( .A(n4935), .ZN(n4609) );
  AND2_X1 U6493 ( .A1(n7353), .A2(n7409), .ZN(n4489) );
  NOR3_X1 U6494 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .A3(
        P1_IR_REG_25__SCAN_IN), .ZN(n6074) );
  AND2_X1 U6495 ( .A1(n9781), .A2(n9726), .ZN(n9820) );
  INV_X1 U6496 ( .A(n9820), .ZN(n9964) );
  XNOR2_X1 U6497 ( .A(n5449), .B(SI_14_), .ZN(n5751) );
  AND2_X1 U6498 ( .A1(n7552), .A2(n5220), .ZN(n4490) );
  AOI21_X1 U6499 ( .B1(n10131), .B2(n5298), .A(n4477), .ZN(n5297) );
  NAND2_X1 U6500 ( .A1(n5483), .A2(n5482), .ZN(n5486) );
  INV_X1 U6501 ( .A(n5715), .ZN(n5089) );
  AND2_X1 U6502 ( .A1(n7789), .A2(n8463), .ZN(n4491) );
  NAND2_X1 U6503 ( .A1(n8120), .A2(n5204), .ZN(n9538) );
  AND2_X1 U6504 ( .A1(n4858), .A2(n9576), .ZN(n4492) );
  AND2_X1 U6505 ( .A1(n4447), .A2(n8436), .ZN(n4493) );
  INV_X1 U6506 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n6078) );
  OR2_X1 U6507 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4494) );
  AND2_X1 U6508 ( .A1(n8402), .A2(n8403), .ZN(n8323) );
  NAND2_X1 U6509 ( .A1(n9641), .A2(n9640), .ZN(n4495) );
  INV_X1 U6510 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4550) );
  NAND2_X1 U6511 ( .A1(n10207), .A2(n10206), .ZN(n4496) );
  OR2_X1 U6512 ( .A1(n4429), .A2(n5113), .ZN(n4497) );
  NAND2_X1 U6513 ( .A1(n7721), .A2(n9690), .ZN(n6329) );
  INV_X1 U6514 ( .A(n7473), .ZN(n4906) );
  NAND2_X1 U6515 ( .A1(n4674), .A2(n4466), .ZN(n6098) );
  NAND2_X1 U6516 ( .A1(n10309), .A2(n7439), .ZN(n7402) );
  INV_X2 U6517 ( .A(n10537), .ZN(n10538) );
  AND2_X1 U6518 ( .A1(n4843), .A2(n7235), .ZN(n4498) );
  XNOR2_X1 U6519 ( .A(n8996), .B(n5985), .ZN(n8189) );
  NAND2_X1 U6520 ( .A1(n6349), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n4499) );
  INV_X1 U6521 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5249) );
  NAND2_X1 U6522 ( .A1(n7280), .A2(n9733), .ZN(n7429) );
  INV_X1 U6523 ( .A(n7312), .ZN(n5265) );
  NOR2_X1 U6524 ( .A1(n7010), .A2(n7503), .ZN(n7508) );
  INV_X1 U6525 ( .A(n7508), .ZN(n4564) );
  NAND2_X1 U6526 ( .A1(n7861), .A2(n7860), .ZN(n10265) );
  INV_X1 U6527 ( .A(n10265), .ZN(n4525) );
  NAND2_X1 U6528 ( .A1(n4977), .A2(n6579), .ZN(n6749) );
  NAND2_X1 U6529 ( .A1(n7426), .A2(n7353), .ZN(n7408) );
  NAND2_X1 U6530 ( .A1(n6714), .A2(n6713), .ZN(n6999) );
  XOR2_X1 U6531 ( .A(n5480), .B(SI_21_), .Z(n4500) );
  INV_X1 U6532 ( .A(n9022), .ZN(n4581) );
  NAND2_X1 U6533 ( .A1(n5124), .A2(n5126), .ZN(n7682) );
  OR2_X1 U6534 ( .A1(n7559), .A2(n9073), .ZN(n5327) );
  INV_X1 U6535 ( .A(n5327), .ZN(n4572) );
  INV_X1 U6536 ( .A(n9477), .ZN(n4980) );
  INV_X1 U6537 ( .A(n4582), .ZN(n8869) );
  INV_X1 U6538 ( .A(n5292), .ZN(n5290) );
  NOR2_X1 U6539 ( .A1(n5322), .A2(n5260), .ZN(n5259) );
  INV_X1 U6540 ( .A(n8068), .ZN(n5200) );
  NAND2_X1 U6541 ( .A1(n5274), .A2(n5062), .ZN(n4501) );
  OR2_X1 U6542 ( .A1(n7535), .A2(n4987), .ZN(n4617) );
  NOR2_X1 U6543 ( .A1(n7155), .A2(n7154), .ZN(n4552) );
  INV_X1 U6544 ( .A(n4855), .ZN(n4854) );
  NAND2_X1 U6545 ( .A1(n10116), .A2(n10270), .ZN(n4855) );
  INV_X1 U6546 ( .A(n8340), .ZN(n8915) );
  NAND2_X1 U6547 ( .A1(n6666), .A2(n6665), .ZN(n10192) );
  AND2_X1 U6548 ( .A1(n8931), .A2(n9047), .ZN(n9079) );
  OR2_X1 U6549 ( .A1(n6330), .A2(n9786), .ZN(n10169) );
  INV_X1 U6550 ( .A(n10169), .ZN(n10189) );
  AND2_X1 U6551 ( .A1(n9906), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4502) );
  AND2_X1 U6552 ( .A1(n9920), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4503) );
  NAND2_X1 U6553 ( .A1(n5779), .A2(n5778), .ZN(n9049) );
  INV_X1 U6554 ( .A(n9049), .ZN(n4778) );
  NAND2_X1 U6555 ( .A1(n5852), .A2(n5851), .ZN(n9028) );
  INV_X1 U6556 ( .A(n9028), .ZN(n4776) );
  NAND2_X1 U6557 ( .A1(n8294), .A2(n8507), .ZN(n4504) );
  AND2_X1 U6558 ( .A1(n8033), .A2(n8032), .ZN(n9446) );
  INV_X1 U6559 ( .A(n9446), .ZN(n5183) );
  AND2_X1 U6560 ( .A1(n6422), .A2(n6421), .ZN(n4505) );
  INV_X1 U6561 ( .A(n4522), .ZN(n5061) );
  NAND2_X1 U6562 ( .A1(n7228), .A2(n6990), .ZN(n4522) );
  INV_X1 U6563 ( .A(n10413), .ZN(n4999) );
  INV_X1 U6564 ( .A(n6990), .ZN(n7134) );
  AND3_X1 U6565 ( .A1(n6759), .A2(n6758), .A3(n6757), .ZN(n6990) );
  AND2_X1 U6566 ( .A1(n6380), .A2(P1_STATE_REG_SCAN_IN), .ZN(n4506) );
  AND2_X1 U6567 ( .A1(n4703), .A2(n4707), .ZN(n4507) );
  INV_X1 U6568 ( .A(n8670), .ZN(n4764) );
  INV_X1 U6569 ( .A(n6386), .ZN(n10007) );
  INV_X1 U6570 ( .A(n8506), .ZN(n5121) );
  NAND2_X1 U6571 ( .A1(n8340), .A2(n8504), .ZN(n4741) );
  AND2_X1 U6572 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n4508) );
  INV_X1 U6573 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n4631) );
  INV_X1 U6574 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10376) );
  INV_X1 U6575 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n4628) );
  NAND2_X1 U6576 ( .A1(n4509), .A2(n8344), .ZN(n7106) );
  OAI21_X1 U6577 ( .B1(n7033), .B2(n8356), .A(n4509), .ZN(n7036) );
  NAND2_X2 U6578 ( .A1(n7584), .A2(n8394), .ZN(n7630) );
  NAND2_X1 U6579 ( .A1(n7491), .A2(n8386), .ZN(n7556) );
  NAND4_X1 U6580 ( .A1(n5790), .A2(n5344), .A3(n4792), .A4(n5351), .ZN(n4678)
         );
  NAND4_X1 U6581 ( .A1(n5349), .A2(n5350), .A3(n5379), .A4(n5701), .ZN(n4679)
         );
  NAND4_X1 U6582 ( .A1(n4400), .A2(n4516), .A3(n8467), .A4(n8775), .ZN(n4515)
         );
  NAND3_X1 U6583 ( .A1(n7788), .A2(n4413), .A3(n8775), .ZN(n4518) );
  NAND4_X1 U6584 ( .A1(n8977), .A2(n5234), .A3(n4519), .A4(n8713), .ZN(n9084)
         );
  NAND3_X1 U6585 ( .A1(n4592), .A2(n5387), .A3(n4591), .ZN(n4521) );
  NAND3_X1 U6586 ( .A1(n4590), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4520) );
  NOR2_X2 U6587 ( .A1(n10080), .A2(n4524), .ZN(n4523) );
  NOR2_X4 U6588 ( .A1(n10004), .A2(n10238), .ZN(n9978) );
  AND2_X2 U6589 ( .A1(n7438), .A2(n4702), .ZN(n7439) );
  NAND3_X1 U6590 ( .A1(n4538), .A2(n4881), .A3(n4882), .ZN(n4537) );
  AND2_X2 U6591 ( .A1(n4903), .A2(n6124), .ZN(n6127) );
  NOR2_X1 U6592 ( .A1(n4553), .A2(n4554), .ZN(n6933) );
  NAND2_X1 U6593 ( .A1(n6859), .A2(n6860), .ZN(n6890) );
  NOR2_X1 U6594 ( .A1(n6915), .A2(n6914), .ZN(n6913) );
  NAND2_X1 U6595 ( .A1(n4564), .A2(n4566), .ZN(n7012) );
  NAND3_X1 U6596 ( .A1(n4577), .A2(n4475), .A3(n4575), .ZN(n4723) );
  OAI211_X2 U6597 ( .C1(n6449), .C2(n5560), .A(n4580), .B(n4472), .ZN(n7104)
         );
  NOR2_X2 U6598 ( .A1(n8852), .A2(n9015), .ZN(n8833) );
  NAND2_X1 U6599 ( .A1(n5559), .A2(n5558), .ZN(n4593) );
  NAND3_X1 U6600 ( .A1(n4610), .A2(n4608), .A3(n4934), .ZN(P2_U3516) );
  OAI21_X2 U6601 ( .B1(n7535), .B2(n4612), .A(n4614), .ZN(n8035) );
  NAND2_X2 U6602 ( .A1(n6387), .A2(n4622), .ZN(n6661) );
  NAND2_X1 U6603 ( .A1(n6460), .A2(n6461), .ZN(n6465) );
  NAND2_X1 U6604 ( .A1(n6529), .A2(n4624), .ZN(n6461) );
  NAND2_X1 U6605 ( .A1(n4625), .A2(n6504), .ZN(n4624) );
  INV_X1 U6606 ( .A(n6530), .ZN(n4625) );
  NAND2_X1 U6607 ( .A1(n4639), .A2(n5551), .ZN(n4828) );
  XNOR2_X1 U6608 ( .A(n4639), .B(n5551), .ZN(n6495) );
  NAND2_X1 U6609 ( .A1(n5401), .A2(n5400), .ZN(n4639) );
  NAND2_X1 U6610 ( .A1(n5167), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n4758) );
  XNOR2_X1 U6611 ( .A(n5789), .B(n5326), .ZN(n7832) );
  NAND2_X1 U6612 ( .A1(n4644), .A2(n4642), .ZN(n9756) );
  NAND3_X1 U6613 ( .A1(n4427), .A2(n4649), .A3(n9964), .ZN(n4856) );
  NAND3_X1 U6614 ( .A1(n8459), .A2(n4449), .A3(n8794), .ZN(n4657) );
  NAND2_X1 U6615 ( .A1(n5122), .A2(n5114), .ZN(n5112) );
  NAND3_X1 U6616 ( .A1(n4662), .A2(n4668), .A3(n4667), .ZN(n4666) );
  NAND2_X1 U6617 ( .A1(n4663), .A2(n4664), .ZN(n4662) );
  NAND2_X1 U6618 ( .A1(n8471), .A2(n8470), .ZN(n4663) );
  NAND2_X1 U6619 ( .A1(n4666), .A2(n5020), .ZN(n4665) );
  INV_X1 U6620 ( .A(n8477), .ZN(n4667) );
  NAND4_X1 U6621 ( .A1(n8464), .A2(n8470), .A3(n8463), .A4(n8494), .ZN(n4668)
         );
  NAND2_X1 U6622 ( .A1(n6098), .A2(n5332), .ZN(n4919) );
  OAI21_X1 U6623 ( .B1(n6734), .B2(n4675), .A(n6091), .ZN(n4674) );
  INV_X1 U6624 ( .A(n6733), .ZN(n4675) );
  INV_X1 U6625 ( .A(n7026), .ZN(n8356) );
  NAND3_X1 U6626 ( .A1(n7294), .A2(n5214), .A3(n7484), .ZN(n4688) );
  NAND2_X1 U6627 ( .A1(n8383), .A2(n7295), .ZN(n4690) );
  NAND2_X2 U6628 ( .A1(n9106), .A2(n5359), .ZN(n5896) );
  NAND3_X1 U6629 ( .A1(n9106), .A2(P2_REG3_REG_1__SCAN_IN), .A3(n5359), .ZN(
        n4693) );
  INV_X1 U6630 ( .A(n5360), .ZN(n9106) );
  NAND3_X1 U6631 ( .A1(n5274), .A2(n6074), .A3(n5273), .ZN(n4695) );
  NAND2_X1 U6632 ( .A1(n9734), .A2(n4696), .ZN(n7389) );
  NAND2_X1 U6633 ( .A1(n6989), .A2(n9602), .ZN(n4708) );
  NAND3_X1 U6634 ( .A1(n4703), .A2(n4707), .A3(n9603), .ZN(n7220) );
  NAND2_X1 U6635 ( .A1(n6950), .A2(n6662), .ZN(n9743) );
  NAND2_X1 U6636 ( .A1(n4708), .A2(n9808), .ZN(n4707) );
  INV_X1 U6637 ( .A(n7228), .ZN(n4710) );
  NAND3_X1 U6638 ( .A1(n5080), .A2(n4718), .A3(n5079), .ZN(n4717) );
  OAI21_X2 U6639 ( .B1(n10137), .B2(n5077), .A(n5075), .ZN(n10114) );
  NAND2_X1 U6640 ( .A1(n10010), .A2(n10009), .ZN(n7993) );
  INV_X1 U6641 ( .A(n10009), .ZN(n4720) );
  NAND4_X1 U6642 ( .A1(n5531), .A2(n4792), .A3(n5344), .A4(n5368), .ZN(n5617)
         );
  OR2_X1 U6643 ( .A1(n4721), .A2(n9103), .ZN(n5601) );
  NAND2_X1 U6644 ( .A1(n4722), .A2(n5085), .ZN(n5084) );
  NAND2_X1 U6645 ( .A1(n4722), .A2(n5691), .ZN(n7138) );
  NAND2_X1 U6646 ( .A1(n7053), .A2(n7054), .ZN(n4722) );
  NAND2_X1 U6647 ( .A1(n8204), .A2(n4725), .ZN(n5833) );
  NAND2_X1 U6648 ( .A1(n8191), .A2(n4732), .ZN(n4731) );
  NAND2_X1 U6649 ( .A1(n5091), .A2(n4734), .ZN(n4733) );
  INV_X1 U6650 ( .A(n5867), .ZN(n4738) );
  NAND2_X1 U6651 ( .A1(n10036), .A2(n7989), .ZN(n10039) );
  NAND2_X2 U6652 ( .A1(n7987), .A2(n7986), .ZN(n10099) );
  XNOR2_X1 U6653 ( .A(n6104), .B(n5512), .ZN(n5515) );
  INV_X1 U6654 ( .A(n7083), .ZN(n5665) );
  OAI21_X2 U6655 ( .B1(n5381), .B2(n5321), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5836) );
  NAND2_X1 U6656 ( .A1(n9674), .A2(n9673), .ZN(n9676) );
  AOI21_X1 U6657 ( .B1(n4870), .B2(n4872), .A(n4495), .ZN(n4869) );
  NAND3_X1 U6658 ( .A1(n9649), .A2(n9747), .A3(n4745), .ZN(n9650) );
  INV_X1 U6659 ( .A(n5515), .ZN(n5513) );
  INV_X1 U6660 ( .A(n5088), .ZN(n5087) );
  BUF_X1 U6661 ( .A(n7729), .Z(n4746) );
  NAND2_X1 U6662 ( .A1(n4800), .A2(n4797), .ZN(n10324) );
  NAND2_X1 U6663 ( .A1(n5399), .A2(n4747), .ZN(n5400) );
  INV_X1 U6664 ( .A(n4748), .ZN(n4747) );
  NAND2_X1 U6665 ( .A1(n10073), .A2(n9692), .ZN(n10051) );
  NAND2_X1 U6666 ( .A1(n5063), .A2(n5064), .ZN(n10073) );
  NAND2_X1 U6667 ( .A1(n10327), .A2(n10499), .ZN(n4756) );
  NAND2_X1 U6668 ( .A1(n10239), .A2(n4457), .ZN(n10327) );
  AND4_X2 U6669 ( .A1(n4867), .A2(n4866), .A3(n4865), .A4(n4902), .ZN(n4864)
         );
  NAND4_X1 U6670 ( .A1(n6337), .A2(n6334), .A3(n6335), .A4(n6336), .ZN(n6663)
         );
  NAND2_X1 U6671 ( .A1(n5274), .A2(n5273), .ZN(n6073) );
  NAND2_X1 U6672 ( .A1(n5513), .A2(n5514), .ZN(n5524) );
  NAND2_X1 U6673 ( .A1(n4930), .A2(n5033), .ZN(n4923) );
  NAND2_X1 U6674 ( .A1(n7703), .A2(n7702), .ZN(n7760) );
  NAND2_X1 U6675 ( .A1(n8757), .A2(n8765), .ZN(n8756) );
  OAI21_X1 U6676 ( .B1(n7139), .B2(n5089), .A(n7332), .ZN(n5088) );
  NAND2_X1 U6677 ( .A1(n4832), .A2(n4830), .ZN(P1_U3520) );
  AOI22_X1 U6678 ( .A1(n10215), .A2(n10464), .B1(n10214), .B2(n10213), .ZN(
        n10216) );
  NAND2_X1 U6679 ( .A1(n6853), .A2(n6852), .ZN(n8625) );
  NAND2_X1 U6680 ( .A1(n6848), .A2(n6847), .ZN(n8598) );
  OAI22_X1 U6681 ( .A1(n8682), .A2(n8681), .B1(n8680), .B2(n8679), .ZN(n4809)
         );
  NAND2_X1 U6682 ( .A1(n4929), .A2(n4928), .ZN(n7703) );
  NAND3_X1 U6683 ( .A1(n5110), .A2(n4966), .A3(n8505), .ZN(P2_U3244) );
  NAND3_X1 U6684 ( .A1(n8429), .A2(n4774), .A3(n4768), .ZN(n8439) );
  NAND3_X1 U6685 ( .A1(n8424), .A2(n8417), .A3(n4769), .ZN(n4768) );
  NAND2_X1 U6686 ( .A1(n8397), .A2(n5031), .ZN(n5030) );
  OR2_X2 U6687 ( .A1(n9067), .A2(n7626), .ZN(n8402) );
  NAND2_X1 U6688 ( .A1(n4781), .A2(n6979), .ZN(n6934) );
  NAND2_X1 U6689 ( .A1(n5630), .A2(n5629), .ZN(n4781) );
  NAND2_X1 U6690 ( .A1(n7756), .A2(n4782), .ZN(P2_U3222) );
  NAND2_X1 U6691 ( .A1(n5238), .A2(n5236), .ZN(P2_U3549) );
  OAI21_X1 U6692 ( .B1(n4409), .B2(n4973), .A(n4487), .ZN(n4972) );
  OAI21_X1 U6693 ( .B1(n5775), .B2(n5774), .A(n5457), .ZN(n5789) );
  INV_X1 U6694 ( .A(n4785), .ZN(n9961) );
  OAI21_X1 U6695 ( .B1(n10217), .B2(n10118), .A(n4786), .ZN(n4785) );
  NAND2_X1 U6696 ( .A1(n7992), .A2(n9747), .ZN(n10010) );
  NAND2_X1 U6697 ( .A1(n4396), .A2(n5394), .ZN(n4953) );
  NAND3_X1 U6698 ( .A1(n4790), .A2(n4788), .A3(n4787), .ZN(P1_U3260) );
  XNOR2_X2 U6699 ( .A(n6125), .B(P1_IR_REG_3__SCAN_IN), .ZN(n10355) );
  NOR2_X2 U6700 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6124) );
  NAND2_X1 U6701 ( .A1(n5109), .A2(n4421), .ZN(n4791) );
  NAND2_X1 U6702 ( .A1(n8162), .A2(n4467), .ZN(n5928) );
  NAND2_X1 U6703 ( .A1(n5580), .A2(n6645), .ZN(n6114) );
  AND2_X1 U6704 ( .A1(n5633), .A2(n5106), .ZN(n5104) );
  NOR2_X1 U6705 ( .A1(n4805), .A2(n4804), .ZN(n4803) );
  INV_X1 U6706 ( .A(n5381), .ZN(n5109) );
  NAND2_X2 U6707 ( .A1(n7391), .A2(n7390), .ZN(n7984) );
  NAND2_X1 U6708 ( .A1(n5150), .A2(n5442), .ZN(n5737) );
  AND2_X1 U6709 ( .A1(n9810), .A2(n9742), .ZN(n9602) );
  INV_X1 U6710 ( .A(n5225), .ZN(n5224) );
  NAND2_X1 U6711 ( .A1(n5470), .A2(n5469), .ZN(n5850) );
  INV_X1 U6712 ( .A(n4972), .ZN(n4971) );
  NAND2_X1 U6713 ( .A1(n4971), .A2(n4973), .ZN(n4968) );
  OAI21_X1 U6714 ( .B1(n8715), .B2(n8899), .A(n4948), .ZN(P2_U3267) );
  NAND2_X1 U6715 ( .A1(n4802), .A2(n6047), .ZN(P2_U3216) );
  NAND3_X1 U6716 ( .A1(n6026), .A2(n7758), .A3(n7733), .ZN(n4802) );
  NAND2_X1 U6717 ( .A1(n6937), .A2(n4803), .ZN(n5667) );
  NAND2_X1 U6718 ( .A1(n5105), .A2(n5104), .ZN(n6937) );
  NAND2_X1 U6719 ( .A1(n5144), .A2(n4491), .ZN(n8736) );
  NAND2_X1 U6720 ( .A1(n4394), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n4816) );
  OAI211_X2 U6721 ( .C1(n7630), .C2(n4944), .A(n4942), .B(n5123), .ZN(n7694)
         );
  NAND2_X1 U6722 ( .A1(n9995), .A2(n9665), .ZN(n9986) );
  OAI21_X1 U6723 ( .B1(n5035), .B2(n8405), .A(n8404), .ZN(n5034) );
  NAND2_X1 U6724 ( .A1(n5034), .A2(n8406), .ZN(n5032) );
  INV_X1 U6725 ( .A(n8490), .ZN(n8488) );
  NAND2_X1 U6726 ( .A1(n5122), .A2(n4497), .ZN(n5111) );
  NAND2_X1 U6727 ( .A1(n8499), .A2(n8498), .ZN(n4815) );
  AND2_X2 U6728 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n9137) );
  NAND2_X1 U6729 ( .A1(n5112), .A2(n4967), .ZN(n4966) );
  AOI21_X4 U6730 ( .B1(n7777), .B2(n7747), .A(n6041), .ZN(n8710) );
  INV_X1 U6731 ( .A(n5264), .ZN(n5263) );
  NAND2_X1 U6732 ( .A1(n9697), .A2(n6944), .ZN(n4829) );
  NAND2_X1 U6733 ( .A1(n4829), .A2(n6658), .ZN(n6712) );
  NAND3_X1 U6734 ( .A1(n6714), .A2(n5280), .A3(n5278), .ZN(n5277) );
  NAND3_X1 U6735 ( .A1(n6945), .A2(n4435), .A3(n5271), .ZN(n6662) );
  AND3_X2 U6736 ( .A1(n4864), .A2(n4454), .A3(n6127), .ZN(n5274) );
  INV_X1 U6737 ( .A(n5274), .ZN(n6371) );
  NAND3_X1 U6738 ( .A1(n7424), .A2(n5283), .A3(n4839), .ZN(n4838) );
  NAND2_X1 U6739 ( .A1(n4841), .A2(n4843), .ZN(n4840) );
  NAND2_X1 U6740 ( .A1(n4489), .A2(n9710), .ZN(n4845) );
  NAND2_X1 U6741 ( .A1(n10091), .A2(n4849), .ZN(n4847) );
  NAND2_X1 U6742 ( .A1(n4856), .A2(n4858), .ZN(n7972) );
  NOR2_X2 U6743 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n4865) );
  NOR2_X2 U6744 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n4866) );
  NAND2_X1 U6745 ( .A1(n4868), .A2(n4873), .ZN(n4871) );
  NAND2_X1 U6746 ( .A1(n9626), .A2(n9625), .ZN(n4868) );
  NAND2_X1 U6747 ( .A1(n9622), .A2(n9621), .ZN(n9634) );
  NAND3_X1 U6748 ( .A1(n9622), .A2(n4875), .A3(n4407), .ZN(n4872) );
  NAND2_X1 U6749 ( .A1(n6662), .A2(n9800), .ZN(n9697) );
  NAND2_X1 U6750 ( .A1(n6694), .A2(n6697), .ZN(n9801) );
  NAND2_X1 U6751 ( .A1(n9676), .A2(n4883), .ZN(n4882) );
  NAND2_X2 U6752 ( .A1(n6280), .A2(n6279), .ZN(n7944) );
  NOR2_X1 U6753 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n4903) );
  NAND2_X1 U6754 ( .A1(n4912), .A2(n4915), .ZN(n9396) );
  NAND2_X1 U6755 ( .A1(n9488), .A2(n4913), .ZN(n4912) );
  AND2_X1 U6756 ( .A1(n4918), .A2(n4474), .ZN(n9455) );
  NAND2_X1 U6757 ( .A1(n4919), .A2(n5324), .ZN(n7290) );
  NAND2_X1 U6758 ( .A1(n8802), .A2(n4920), .ZN(n8772) );
  NAND2_X1 U6759 ( .A1(n8368), .A2(n8344), .ZN(n7026) );
  NAND2_X1 U6760 ( .A1(n6622), .A2(n6094), .ZN(n8368) );
  NAND3_X1 U6761 ( .A1(n4926), .A2(n7678), .A3(n4923), .ZN(n7701) );
  NAND3_X1 U6762 ( .A1(n4926), .A2(n4924), .A3(n4923), .ZN(n4929) );
  OAI21_X1 U6763 ( .B1(n7620), .B2(n5219), .A(n5218), .ZN(n4930) );
  NAND2_X1 U6764 ( .A1(n8976), .A2(n10536), .ZN(n4932) );
  NOR2_X1 U6765 ( .A1(n8976), .A2(n4609), .ZN(n8983) );
  NAND3_X1 U6766 ( .A1(n4932), .A2(n8982), .A3(n4931), .ZN(n9085) );
  OAI21_X1 U6767 ( .B1(n7630), .B2(n7629), .A(n8399), .ZN(n7661) );
  MUX2_X1 U6768 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n4393), .Z(n5410) );
  NAND2_X1 U6769 ( .A1(n5398), .A2(n5536), .ZN(n5401) );
  NAND2_X1 U6770 ( .A1(n4953), .A2(n4952), .ZN(n5536) );
  NAND2_X1 U6771 ( .A1(n4393), .A2(n5397), .ZN(n4952) );
  NAND2_X1 U6772 ( .A1(n5411), .A2(n5582), .ZN(n4954) );
  NAND2_X1 U6773 ( .A1(n5160), .A2(n4416), .ZN(n4962) );
  NAND2_X1 U6774 ( .A1(n5160), .A2(n4956), .ZN(n4955) );
  NAND2_X1 U6775 ( .A1(n8010), .A2(n8009), .ZN(n8300) );
  NAND3_X1 U6776 ( .A1(n8300), .A2(n8299), .A3(n8298), .ZN(n4964) );
  NAND2_X1 U6777 ( .A1(n4964), .A2(n8304), .ZN(n4963) );
  NAND2_X1 U6778 ( .A1(n5149), .A2(n4971), .ZN(n4969) );
  NAND2_X1 U6779 ( .A1(n5149), .A2(n4409), .ZN(n4970) );
  NAND3_X1 U6780 ( .A1(n4969), .A2(n5169), .A3(n4968), .ZN(n5835) );
  NAND2_X1 U6781 ( .A1(n6575), .A2(n6574), .ZN(n4977) );
  NAND2_X1 U6782 ( .A1(n4978), .A2(n6511), .ZN(n6575) );
  NAND2_X1 U6783 ( .A1(n6506), .A2(n6507), .ZN(n4978) );
  AND4_X2 U6784 ( .A1(n4988), .A2(n7472), .A3(n7470), .A4(n7471), .ZN(n7535)
         );
  XNOR2_X2 U6785 ( .A(n4990), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6132) );
  NOR2_X2 U6786 ( .A1(n6054), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n5273) );
  NAND3_X1 U6787 ( .A1(n4995), .A2(n4994), .A3(n4991), .ZN(n9929) );
  NAND2_X1 U6788 ( .A1(n6425), .A2(n5009), .ZN(n5006) );
  NAND2_X1 U6789 ( .A1(n5006), .A2(n5007), .ZN(n6686) );
  AOI21_X1 U6790 ( .B1(n8359), .B2(n8358), .A(n5025), .ZN(n5024) );
  NAND3_X1 U6791 ( .A1(n5032), .A2(n5030), .A3(n8412), .ZN(n8424) );
  INV_X1 U6792 ( .A(n5896), .ZN(n5037) );
  NAND2_X1 U6793 ( .A1(n5999), .A2(n5039), .ZN(n5357) );
  NAND2_X1 U6794 ( .A1(n4428), .A2(n5999), .ZN(n5040) );
  INV_X1 U6795 ( .A(n5049), .ZN(n10058) );
  NAND2_X1 U6796 ( .A1(n9978), .A2(n9984), .ZN(n9979) );
  NOR2_X2 U6797 ( .A1(n9979), .A2(n5053), .ZN(n5052) );
  NAND2_X1 U6798 ( .A1(n5054), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6077) );
  NAND3_X1 U6799 ( .A1(n5274), .A2(n5313), .A3(n5273), .ZN(n5054) );
  NAND2_X1 U6800 ( .A1(n10099), .A2(n4445), .ZN(n5063) );
  NAND2_X1 U6801 ( .A1(n7993), .A2(n9774), .ZN(n9995) );
  NAND2_X1 U6802 ( .A1(n6211), .A2(n6380), .ZN(n6079) );
  INV_X2 U6803 ( .A(n6380), .ZN(n7858) );
  OAI21_X1 U6804 ( .B1(n10137), .B2(n9581), .A(n9737), .ZN(n10132) );
  NAND2_X1 U6805 ( .A1(n9968), .A2(n7995), .ZN(n9952) );
  NAND2_X1 U6806 ( .A1(n5083), .A2(n5524), .ZN(n6621) );
  NAND2_X1 U6807 ( .A1(n5083), .A2(n5082), .ZN(n6614) );
  OR2_X1 U6808 ( .A1(n6612), .A2(n6613), .ZN(n5082) );
  NAND2_X1 U6809 ( .A1(n5084), .A2(n5087), .ZN(n5736) );
  NAND2_X1 U6810 ( .A1(n8151), .A2(n5102), .ZN(n5813) );
  NAND2_X1 U6811 ( .A1(n6114), .A2(n5614), .ZN(n5105) );
  NAND3_X1 U6812 ( .A1(n4421), .A2(n5108), .A3(n5636), .ZN(n5107) );
  NAND3_X1 U6813 ( .A1(n5111), .A2(n8313), .A3(n5121), .ZN(n5110) );
  NAND2_X1 U6814 ( .A1(n5135), .A2(n5136), .ZN(n8295) );
  NAND2_X1 U6815 ( .A1(n8284), .A2(n5138), .ZN(n5135) );
  AND2_X1 U6816 ( .A1(n8975), .A2(n8479), .ZN(n5139) );
  XNOR2_X1 U6817 ( .A(n8316), .B(n6099), .ZN(n7110) );
  NAND2_X1 U6818 ( .A1(n5470), .A2(n5162), .ZN(n5160) );
  NAND3_X1 U6819 ( .A1(n5252), .A2(n6496), .A3(n5168), .ZN(n5250) );
  NAND3_X1 U6820 ( .A1(n5171), .A2(n5174), .A3(n5818), .ZN(n5170) );
  INV_X1 U6821 ( .A(n9690), .ZN(n6378) );
  NAND2_X4 U6822 ( .A1(n5179), .A2(n6520), .ZN(n8127) );
  NAND2_X1 U6823 ( .A1(n6782), .A2(n5191), .ZN(n5189) );
  NAND3_X1 U6824 ( .A1(n6749), .A2(n6748), .A3(n6782), .ZN(n5190) );
  NAND2_X1 U6825 ( .A1(n5192), .A2(n6753), .ZN(n6872) );
  INV_X1 U6826 ( .A(n6753), .ZN(n5191) );
  NAND2_X1 U6827 ( .A1(n8120), .A2(n8119), .ZN(n9537) );
  INV_X1 U6828 ( .A(n9536), .ZN(n5206) );
  INV_X1 U6829 ( .A(n7293), .ZN(n5214) );
  NAND2_X1 U6830 ( .A1(n5581), .A2(n5409), .ZN(n5215) );
  INV_X1 U6831 ( .A(n7621), .ZN(n5217) );
  NAND3_X1 U6832 ( .A1(n5217), .A2(n4490), .A3(n7553), .ZN(n5216) );
  NAND2_X1 U6833 ( .A1(n7553), .A2(n7552), .ZN(n7622) );
  NAND2_X1 U6834 ( .A1(n8323), .A2(n5220), .ZN(n5218) );
  OR2_X1 U6835 ( .A1(n9067), .A2(n8519), .ZN(n5220) );
  NAND2_X1 U6836 ( .A1(n7774), .A2(n5235), .ZN(n5234) );
  NAND2_X1 U6837 ( .A1(n9084), .A2(n10544), .ZN(n5238) );
  OR2_X1 U6838 ( .A1(n10544), .A2(n5237), .ZN(n5236) );
  NAND2_X1 U6839 ( .A1(n7760), .A2(n5241), .ZN(n8901) );
  NAND2_X1 U6840 ( .A1(n7768), .A2(n5245), .ZN(n5244) );
  NAND3_X1 U6841 ( .A1(n5250), .A2(n5251), .A3(n5248), .ZN(n5402) );
  NAND3_X1 U6842 ( .A1(n5388), .A2(n5387), .A3(n5249), .ZN(n5248) );
  NAND3_X1 U6843 ( .A1(n5389), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(n5249), .ZN(
        n5251) );
  INV_X1 U6844 ( .A(n6104), .ZN(n5254) );
  NAND2_X1 U6845 ( .A1(n7578), .A2(n7579), .ZN(n7559) );
  NAND3_X1 U6846 ( .A1(n5277), .A2(n7001), .A3(n5275), .ZN(n7236) );
  NAND2_X1 U6847 ( .A1(n5278), .A2(n5276), .ZN(n5275) );
  INV_X1 U6848 ( .A(n7424), .ZN(n5287) );
  NAND2_X1 U6849 ( .A1(n5311), .A2(n6075), .ZN(n10344) );
  NAND2_X1 U6850 ( .A1(n5976), .A2(n5975), .ZN(n5978) );
  NAND2_X1 U6851 ( .A1(n7711), .A2(n7710), .ZN(n7713) );
  NAND2_X1 U6852 ( .A1(n9724), .A2(n9951), .ZN(n9576) );
  NAND2_X1 U6853 ( .A1(n5835), .A2(n5467), .ZN(n5470) );
  NAND2_X1 U6854 ( .A1(n6617), .A2(n7050), .ZN(n6605) );
  NAND2_X1 U6855 ( .A1(n8361), .A2(n8362), .ZN(n6733) );
  XNOR2_X1 U6856 ( .A(n5954), .B(n5953), .ZN(n7924) );
  INV_X1 U6857 ( .A(n8840), .ZN(n8791) );
  OR2_X1 U6858 ( .A1(n5526), .A2(n5525), .ZN(n5529) );
  OR2_X1 U6859 ( .A1(n5526), .A2(n5499), .ZN(n5503) );
  XOR2_X1 U6860 ( .A(n8963), .B(n8693), .Z(n8965) );
  AND2_X1 U6861 ( .A1(n7972), .A2(n7971), .ZN(n7973) );
  INV_X1 U6862 ( .A(n8958), .ZN(n8940) );
  AND2_X1 U6863 ( .A1(n10218), .A2(n10476), .ZN(n5314) );
  AND2_X1 U6864 ( .A1(n8973), .A2(n10536), .ZN(n5315) );
  AND2_X1 U6865 ( .A1(n5664), .A2(n6980), .ZN(n5317) );
  AND3_X1 U6866 ( .A1(n8375), .A2(n7300), .A3(n8376), .ZN(n5318) );
  AND2_X1 U6867 ( .A1(n5674), .A2(n5652), .ZN(n5319) );
  INV_X1 U6868 ( .A(SI_17_), .ZN(n5464) );
  AND2_X1 U6869 ( .A1(n10219), .A2(n5314), .ZN(n5320) );
  OR2_X1 U6870 ( .A1(n5375), .A2(n5374), .ZN(n5321) );
  INV_X1 U6871 ( .A(n8742), .ZN(n8510) );
  INV_X1 U6872 ( .A(n8193), .ZN(n8727) );
  AND3_X1 U6873 ( .A1(n8459), .A2(n8434), .A3(n8794), .ZN(n5323) );
  AND2_X1 U6874 ( .A1(n7261), .A2(n6100), .ZN(n5324) );
  INV_X1 U6875 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n6076) );
  AND2_X1 U6876 ( .A1(n5448), .A2(n5447), .ZN(n5325) );
  INV_X1 U6877 ( .A(n8886), .ZN(n8924) );
  AND2_X1 U6878 ( .A1(n5463), .A2(n5462), .ZN(n5326) );
  XNOR2_X1 U6879 ( .A(n6504), .B(n8034), .ZN(n5328) );
  AND3_X1 U6880 ( .A1(n6471), .A2(n6470), .A3(n6469), .ZN(n5329) );
  AND2_X1 U6881 ( .A1(n9517), .A2(n9414), .ZN(n5330) );
  INV_X1 U6882 ( .A(n8694), .ZN(n8293) );
  INV_X1 U6883 ( .A(n8738), .ZN(n7789) );
  OR2_X1 U6884 ( .A1(n8942), .A2(n8278), .ZN(n5331) );
  AND2_X1 U6885 ( .A1(n6097), .A2(n6096), .ZN(n5332) );
  INV_X1 U6886 ( .A(n8411), .ZN(n7683) );
  AND2_X1 U6887 ( .A1(n8143), .A2(n9507), .ZN(n5333) );
  INV_X1 U6888 ( .A(n10523), .ZN(n6099) );
  INV_X1 U6889 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n6048) );
  INV_X1 U6890 ( .A(n8421), .ZN(n7782) );
  INV_X1 U6891 ( .A(n5331), .ZN(n7783) );
  INV_X1 U6892 ( .A(P2_RD_REG_SCAN_IN), .ZN(n9227) );
  NAND2_X1 U6893 ( .A1(n6090), .A2(n6104), .ZN(n8362) );
  INV_X1 U6894 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5369) );
  NAND2_X1 U6895 ( .A1(n6393), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n6389) );
  OR2_X1 U6896 ( .A1(n10260), .A2(n10086), .ZN(n7879) );
  INV_X1 U6897 ( .A(n9638), .ZN(n7986) );
  OAI21_X1 U6898 ( .B1(n6695), .B2(n6655), .A(n10447), .ZN(n6657) );
  INV_X1 U6899 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6064) );
  INV_X1 U6900 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5368) );
  AOI21_X1 U6901 ( .B1(n7467), .B2(n7473), .A(n7474), .ZN(n7468) );
  INV_X1 U6902 ( .A(n7177), .ZN(n7170) );
  AOI21_X1 U6903 ( .B1(n8038), .B2(n9462), .A(n8037), .ZN(n9466) );
  OR2_X1 U6904 ( .A1(n6593), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6469) );
  INV_X1 U6905 ( .A(n9624), .ZN(n7390) );
  INV_X1 U6906 ( .A(n10184), .ZN(n7985) );
  INV_X1 U6907 ( .A(SI_19_), .ZN(n9249) );
  NOR2_X1 U6908 ( .A1(n5676), .A2(n5422), .ZN(n5695) );
  NAND2_X1 U6909 ( .A1(n5269), .A2(n8193), .ZN(n7772) );
  AOI21_X1 U6910 ( .B1(n5836), .B2(n5376), .A(n9103), .ZN(n5384) );
  INV_X1 U6911 ( .A(n6520), .ZN(n6393) );
  NAND2_X1 U6912 ( .A1(n7469), .A2(n7468), .ZN(n7470) );
  NOR2_X1 U6913 ( .A1(n8090), .A2(n5330), .ZN(n8091) );
  INV_X1 U6914 ( .A(n10443), .ZN(n6627) );
  NAND2_X1 U6915 ( .A1(n9789), .A2(n6378), .ZN(n6330) );
  INV_X1 U6916 ( .A(n9957), .ZN(n9958) );
  NAND2_X1 U6917 ( .A1(n10309), .A2(n7532), .ZN(n7409) );
  NAND2_X1 U6918 ( .A1(n5476), .A2(n5475), .ZN(n5479) );
  NAND2_X1 U6919 ( .A1(n5460), .A2(n5459), .ZN(n5463) );
  NAND2_X1 U6920 ( .A1(n5445), .A2(n5444), .ZN(n5448) );
  INV_X1 U6921 ( .A(n5996), .ZN(n5997) );
  INV_X1 U6922 ( .A(n8162), .ZN(n8219) );
  INV_X1 U6923 ( .A(n8188), .ZN(n5952) );
  INV_X1 U6924 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9163) );
  OR2_X1 U6925 ( .A1(n6817), .A2(n6816), .ZN(n6862) );
  INV_X1 U6926 ( .A(n8978), .ZN(n7779) );
  OR2_X1 U6927 ( .A1(n9047), .A2(n8350), .ZN(n6482) );
  AND2_X1 U6928 ( .A1(n6490), .A2(n6032), .ZN(n9074) );
  INV_X1 U6929 ( .A(n9550), .ZN(n9531) );
  INV_X1 U6930 ( .A(n6593), .ZN(n7955) );
  CLKBUF_X3 U6931 ( .A(n6341), .Z(n7974) );
  NOR2_X1 U6932 ( .A1(n5052), .A2(n5156), .ZN(n9946) );
  INV_X1 U6933 ( .A(n9841), .ZN(n9997) );
  INV_X1 U6934 ( .A(n10192), .ZN(n10165) );
  AND2_X1 U6935 ( .A1(n6667), .A2(n6402), .ZN(n6677) );
  XNOR2_X1 U6936 ( .A(n5468), .B(SI_18_), .ZN(n5834) );
  OAI21_X1 U6937 ( .B1(n4397), .B2(P1_DATAO_REG_4__SCAN_IN), .A(n5405), .ZN(
        n5406) );
  AND2_X1 U6938 ( .A1(n6033), .A2(n8502), .ZN(n8227) );
  INV_X1 U6939 ( .A(n8273), .ZN(n8254) );
  AND2_X1 U6940 ( .A1(n6031), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8273) );
  INV_X1 U6941 ( .A(n8339), .ZN(n8504) );
  INV_X1 U6942 ( .A(n8677), .ZN(n8661) );
  AND2_X1 U6943 ( .A1(n6862), .A2(n6818), .ZN(n8675) );
  INV_X1 U6944 ( .A(n8792), .ZN(n8822) );
  AND2_X1 U6945 ( .A1(n6814), .A2(n6035), .ZN(n8886) );
  AND2_X1 U6946 ( .A1(n7679), .A2(n7625), .ZN(n9063) );
  INV_X1 U6947 ( .A(n8325), .ZN(n8383) );
  OR2_X1 U6948 ( .A1(n6482), .A2(n10501), .ZN(n8954) );
  NAND2_X1 U6949 ( .A1(n4741), .A2(n8314), .ZN(n8935) );
  INV_X1 U6950 ( .A(n6731), .ZN(n6486) );
  INV_X1 U6951 ( .A(n9079), .ZN(n10536) );
  AOI21_X1 U6952 ( .B1(n7653), .B2(n6013), .A(n9122), .ZN(n10500) );
  AND2_X1 U6953 ( .A1(n5776), .A2(n5758), .ZN(n7015) );
  INV_X1 U6954 ( .A(n9924), .ZN(n10416) );
  INV_X1 U6955 ( .A(n9923), .ZN(n10425) );
  INV_X1 U6956 ( .A(n10205), .ZN(n10219) );
  AND2_X1 U6957 ( .A1(n9657), .A2(n9766), .ZN(n10084) );
  AND2_X1 U6958 ( .A1(n6994), .A2(n10157), .ZN(n10180) );
  INV_X1 U6959 ( .A(n10476), .ZN(n10299) );
  AND2_X1 U6960 ( .A1(n6324), .A2(n6323), .ZN(n6679) );
  OR3_X1 U6961 ( .A1(n6132), .A2(n6136), .A3(n6135), .ZN(n10429) );
  XNOR2_X1 U6962 ( .A(n6077), .B(n6076), .ZN(n6197) );
  INV_X1 U6963 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6070) );
  XNOR2_X1 U6964 ( .A(n5650), .B(n5649), .ZN(n7171) );
  NAND2_X1 U6965 ( .A1(n6177), .A2(n6176), .ZN(n8685) );
  NAND2_X1 U6966 ( .A1(n8227), .A2(n8886), .ZN(n8263) );
  INV_X1 U6967 ( .A(n8280), .ZN(n8268) );
  OR2_X1 U6968 ( .A1(n7732), .A2(n7731), .ZN(n8282) );
  INV_X1 U6969 ( .A(n8848), .ZN(n8889) );
  INV_X1 U6970 ( .A(n8957), .ZN(n8944) );
  AND2_X1 U6971 ( .A1(n7048), .A2(n8954), .ZN(n8958) );
  AND2_X1 U6972 ( .A1(n7634), .A2(n7633), .ZN(n9065) );
  INV_X1 U6973 ( .A(n8940), .ZN(n8949) );
  OR2_X1 U6974 ( .A1(n6731), .A2(n6730), .ZN(n10537) );
  NOR2_X1 U6975 ( .A1(n10501), .A2(n10500), .ZN(n10508) );
  INV_X1 U6976 ( .A(n10508), .ZN(n10511) );
  INV_X1 U6977 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n9253) );
  INV_X1 U6978 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6419) );
  INV_X1 U6979 ( .A(n9386), .ZN(n9118) );
  OR2_X1 U6980 ( .A1(n6409), .A2(n9786), .ZN(n9529) );
  INV_X1 U6981 ( .A(n9556), .ZN(n9544) );
  NAND2_X1 U6982 ( .A1(n7980), .A2(n7979), .ZN(n10208) );
  INV_X1 U6983 ( .A(n10139), .ZN(n10115) );
  OR2_X1 U6984 ( .A1(n10408), .A2(n10403), .ZN(n9923) );
  NAND2_X1 U6985 ( .A1(n10170), .A2(n7004), .ZN(n10197) );
  OR3_X1 U6986 ( .A1(n10118), .A2(n6696), .A3(n10059), .ZN(n10150) );
  AND2_X2 U6987 ( .A1(n6679), .A2(n6678), .ZN(n10499) );
  INV_X1 U6988 ( .A(n10499), .ZN(n10496) );
  INV_X1 U6989 ( .A(n10488), .ZN(n10486) );
  AND2_X1 U6990 ( .A1(n10443), .A2(n10429), .ZN(n10439) );
  NOR2_X1 U6991 ( .A1(n10588), .A2(n10587), .ZN(n10586) );
  NOR2_X1 U6992 ( .A1(n10573), .A2(n10572), .ZN(n10571) );
  INV_X1 U6993 ( .A(n8514), .ZN(P2_U3966) );
  OR2_X2 U6994 ( .A1(n5681), .A2(n9163), .ZN(n5725) );
  INV_X1 U6995 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5780) );
  INV_X1 U6996 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5839) );
  INV_X1 U6997 ( .A(n5881), .ZN(n5341) );
  AND2_X1 U6998 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(P2_REG3_REG_20__SCAN_IN), 
        .ZN(n5340) );
  INV_X1 U6999 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8166) );
  INV_X1 U7000 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5342) );
  NAND2_X1 U7001 ( .A1(n5921), .A2(n5342), .ZN(n5343) );
  NAND2_X1 U7002 ( .A1(n5945), .A2(n5343), .ZN(n8779) );
  NOR2_X4 U7003 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5531) );
  NOR2_X2 U7004 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5344) );
  NOR2_X1 U7005 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5347) );
  NOR2_X1 U7006 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5352) );
  INV_X1 U7007 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5355) );
  OR2_X1 U7008 ( .A1(n8779), .A2(n5896), .ZN(n5367) );
  INV_X1 U7009 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n5364) );
  NAND2_X1 U7010 ( .A1(n5360), .A2(n5359), .ZN(n5526) );
  NAND2_X1 U7011 ( .A1(n7743), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5363) );
  NAND2_X2 U7012 ( .A1(n9106), .A2(n5361), .ZN(n5545) );
  NAND2_X1 U7013 ( .A1(n8288), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5362) );
  OAI211_X1 U7014 ( .C1(n5364), .C2(n5826), .A(n5363), .B(n5362), .ZN(n5365)
         );
  INV_X1 U7015 ( .A(n5365), .ZN(n5366) );
  NOR2_X1 U7016 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n5371) );
  INV_X1 U7017 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5756) );
  INV_X1 U7018 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5370) );
  NAND4_X1 U7019 ( .A1(n5371), .A2(n5756), .A3(n5701), .A4(n5370), .ZN(n5375)
         );
  INV_X1 U7020 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n9162) );
  INV_X1 U7021 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5373) );
  INV_X1 U7022 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5795) );
  INV_X1 U7023 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5372) );
  NAND4_X1 U7024 ( .A1(n9162), .A2(n5373), .A3(n5795), .A4(n5372), .ZN(n5374)
         );
  INV_X1 U7025 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5376) );
  INV_X1 U7026 ( .A(n5384), .ZN(n5378) );
  INV_X1 U7027 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5377) );
  NAND2_X1 U7028 ( .A1(n5378), .A2(n5377), .ZN(n5385) );
  XNOR2_X2 U7029 ( .A(n5380), .B(n5379), .ZN(n6025) );
  XNOR2_X1 U7030 ( .A(n6005), .B(n6004), .ZN(n8339) );
  INV_X1 U7031 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5382) );
  NAND2_X1 U7032 ( .A1(n5384), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n5386) );
  AND2_X2 U7033 ( .A1(n5386), .A2(n5385), .ZN(n8340) );
  OR2_X1 U7034 ( .A1(n8192), .A2(n4796), .ZN(n5916) );
  INV_X1 U7035 ( .A(n5916), .ZN(n8221) );
  INV_X1 U7036 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6496) );
  INV_X1 U7037 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6122) );
  NAND2_X1 U7038 ( .A1(n4397), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5390) );
  INV_X1 U7039 ( .A(SI_2_), .ZN(n5535) );
  OAI211_X1 U7040 ( .C1(n4395), .C2(n6122), .A(n5390), .B(n5535), .ZN(n5398)
         );
  NOR2_X1 U7041 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(SI_1_), .ZN(n5393) );
  AND2_X1 U7042 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5506) );
  INV_X1 U7043 ( .A(n5506), .ZN(n5392) );
  NAND2_X1 U7044 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(SI_1_), .ZN(n5391) );
  OAI21_X1 U7045 ( .B1(n5393), .B2(n5392), .A(n5391), .ZN(n5394) );
  NOR2_X1 U7046 ( .A1(SI_1_), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5396) );
  NAND2_X1 U7047 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5507) );
  NAND2_X1 U7048 ( .A1(SI_1_), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5395) );
  OAI21_X1 U7049 ( .B1(n5396), .B2(n5507), .A(n5395), .ZN(n5397) );
  INV_X1 U7050 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6448) );
  NAND2_X1 U7051 ( .A1(n4396), .A2(n6448), .ZN(n5399) );
  INV_X1 U7052 ( .A(n5402), .ZN(n5403) );
  NAND2_X1 U7053 ( .A1(n5403), .A2(SI_3_), .ZN(n5404) );
  INV_X1 U7054 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6123) );
  INV_X1 U7055 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6581) );
  NAND2_X1 U7056 ( .A1(n4396), .A2(n6581), .ZN(n5405) );
  INV_X1 U7057 ( .A(n5406), .ZN(n5407) );
  NAND2_X1 U7058 ( .A1(n5407), .A2(SI_4_), .ZN(n5408) );
  XNOR2_X1 U7059 ( .A(n5410), .B(SI_5_), .ZN(n5582) );
  MUX2_X1 U7060 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n4397), .Z(n5428) );
  XNOR2_X1 U7061 ( .A(n5428), .B(SI_7_), .ZN(n5615) );
  INV_X1 U7062 ( .A(n5615), .ZN(n5414) );
  INV_X1 U7063 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6195) );
  MUX2_X1 U7064 ( .A(n6195), .B(n9207), .S(n4394), .Z(n5416) );
  INV_X1 U7065 ( .A(SI_10_), .ZN(n5415) );
  INV_X1 U7066 ( .A(n5416), .ZN(n5417) );
  NAND2_X1 U7067 ( .A1(n5417), .A2(SI_10_), .ZN(n5418) );
  NAND2_X1 U7068 ( .A1(n5697), .A2(n5418), .ZN(n5676) );
  INV_X1 U7069 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5420) );
  INV_X1 U7070 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5419) );
  MUX2_X1 U7071 ( .A(n5420), .B(n5419), .S(n4394), .Z(n5431) );
  INV_X1 U7072 ( .A(n5431), .ZN(n5421) );
  NAND2_X1 U7073 ( .A1(n5421), .A2(SI_9_), .ZN(n5652) );
  INV_X1 U7074 ( .A(n5652), .ZN(n5422) );
  INV_X1 U7075 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n5423) );
  INV_X1 U7076 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6166) );
  MUX2_X1 U7077 ( .A(n5423), .B(n6166), .S(n4396), .Z(n5425) );
  INV_X1 U7078 ( .A(SI_8_), .ZN(n5424) );
  NAND2_X1 U7079 ( .A1(n5425), .A2(n5424), .ZN(n5651) );
  INV_X1 U7080 ( .A(n5425), .ZN(n5426) );
  NAND2_X1 U7081 ( .A1(n5426), .A2(SI_8_), .ZN(n5427) );
  INV_X1 U7082 ( .A(n5649), .ZN(n5429) );
  NAND2_X1 U7083 ( .A1(n5428), .A2(SI_7_), .ZN(n5634) );
  INV_X1 U7084 ( .A(SI_9_), .ZN(n5430) );
  NAND2_X1 U7085 ( .A1(n5431), .A2(n5430), .ZN(n5674) );
  NAND2_X1 U7086 ( .A1(n5651), .A2(n5674), .ZN(n5692) );
  INV_X1 U7087 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5432) );
  MUX2_X1 U7088 ( .A(n5432), .B(n6190), .S(n4394), .Z(n5433) );
  XNOR2_X1 U7089 ( .A(n5433), .B(SI_11_), .ZN(n5699) );
  INV_X1 U7090 ( .A(n5433), .ZN(n5434) );
  NAND2_X1 U7091 ( .A1(n5434), .A2(SI_11_), .ZN(n5435) );
  INV_X1 U7092 ( .A(n5439), .ZN(n5440) );
  NAND2_X1 U7093 ( .A1(n5440), .A2(SI_12_), .ZN(n5441) );
  MUX2_X1 U7094 ( .A(n9294), .B(n5443), .S(n4396), .Z(n5445) );
  INV_X1 U7095 ( .A(SI_13_), .ZN(n5444) );
  INV_X1 U7096 ( .A(n5445), .ZN(n5446) );
  NAND2_X1 U7097 ( .A1(n5446), .A2(SI_13_), .ZN(n5447) );
  MUX2_X1 U7098 ( .A(n6268), .B(n7805), .S(n4396), .Z(n5449) );
  INV_X1 U7099 ( .A(n5449), .ZN(n5450) );
  NAND2_X1 U7100 ( .A1(n5450), .A2(SI_14_), .ZN(n5451) );
  MUX2_X1 U7101 ( .A(n6417), .B(n5452), .S(n4395), .Z(n5454) );
  INV_X1 U7102 ( .A(n5454), .ZN(n5455) );
  NAND2_X1 U7103 ( .A1(n5455), .A2(SI_15_), .ZN(n5456) );
  MUX2_X1 U7104 ( .A(n6419), .B(n5458), .S(n4397), .Z(n5460) );
  INV_X1 U7105 ( .A(n5460), .ZN(n5461) );
  NAND2_X1 U7106 ( .A1(n5461), .A2(SI_16_), .ZN(n5462) );
  MUX2_X1 U7107 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n4397), .Z(n5465) );
  NAND2_X1 U7108 ( .A1(n5465), .A2(SI_17_), .ZN(n5466) );
  MUX2_X1 U7109 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4394), .Z(n5468) );
  NAND2_X1 U7110 ( .A1(n5468), .A2(SI_18_), .ZN(n5469) );
  MUX2_X1 U7111 ( .A(n6743), .B(n8005), .S(n4394), .Z(n5471) );
  INV_X1 U7112 ( .A(n5471), .ZN(n5472) );
  NAND2_X1 U7113 ( .A1(n5472), .A2(SI_19_), .ZN(n5473) );
  MUX2_X1 U7114 ( .A(n9374), .B(n7868), .S(n4395), .Z(n5476) );
  INV_X1 U7115 ( .A(SI_20_), .ZN(n5475) );
  INV_X1 U7116 ( .A(n5476), .ZN(n5477) );
  NAND2_X1 U7117 ( .A1(n5477), .A2(SI_20_), .ZN(n5478) );
  MUX2_X1 U7118 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n4396), .Z(n5480) );
  NAND2_X1 U7119 ( .A1(n5480), .A2(SI_21_), .ZN(n5481) );
  MUX2_X1 U7120 ( .A(n7722), .B(n7894), .S(n4397), .Z(n5483) );
  INV_X1 U7121 ( .A(SI_22_), .ZN(n5482) );
  INV_X1 U7122 ( .A(n5483), .ZN(n5484) );
  NAND2_X1 U7123 ( .A1(n5484), .A2(SI_22_), .ZN(n5485) );
  INV_X1 U7124 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5487) );
  MUX2_X1 U7125 ( .A(n5487), .B(n7900), .S(n4394), .Z(n5488) );
  INV_X1 U7126 ( .A(SI_23_), .ZN(n9335) );
  NAND2_X1 U7127 ( .A1(n5488), .A2(n9335), .ZN(n5491) );
  INV_X1 U7128 ( .A(n5488), .ZN(n5489) );
  NAND2_X1 U7129 ( .A1(n5489), .A2(SI_23_), .ZN(n5490) );
  INV_X1 U7130 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7526) );
  MUX2_X1 U7131 ( .A(n7526), .B(n7912), .S(n4395), .Z(n5932) );
  XNOR2_X1 U7132 ( .A(n5932), .B(SI_24_), .ZN(n5931) );
  XNOR2_X1 U7133 ( .A(n5936), .B(n5931), .ZN(n7911) );
  INV_X4 U7134 ( .A(n5560), .ZN(n8307) );
  NAND2_X1 U7135 ( .A1(n7911), .A2(n8307), .ZN(n5498) );
  NAND2_X1 U7136 ( .A1(n8308), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5497) );
  XNOR2_X1 U7137 ( .A(n4746), .B(n9000), .ZN(n8222) );
  INV_X1 U7138 ( .A(n8222), .ZN(n5930) );
  INV_X1 U7139 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n5499) );
  INV_X1 U7140 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n5500) );
  INV_X1 U7141 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6839) );
  OR2_X1 U7142 ( .A1(n5545), .A2(n6839), .ZN(n5502) );
  NAND2_X1 U7143 ( .A1(n5640), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5501) );
  NOR2_X1 U7144 ( .A1(n6090), .A2(n7728), .ZN(n5516) );
  INV_X1 U7145 ( .A(n5516), .ZN(n5514) );
  INV_X1 U7146 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5505) );
  NAND2_X1 U7147 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5504) );
  INV_X1 U7148 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6121) );
  NAND2_X1 U7149 ( .A1(n4395), .A2(n5506), .ZN(n6327) );
  OAI21_X1 U7150 ( .B1(n4394), .B2(n5507), .A(n6327), .ZN(n5509) );
  INV_X1 U7151 ( .A(SI_1_), .ZN(n5508) );
  XNOR2_X1 U7152 ( .A(n5509), .B(n5508), .ZN(n5511) );
  MUX2_X1 U7153 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n4395), .Z(n5510) );
  NAND2_X1 U7154 ( .A1(n5516), .A2(n5515), .ZN(n5517) );
  NAND2_X1 U7155 ( .A1(n5640), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5521) );
  INV_X1 U7156 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6972) );
  OR2_X1 U7157 ( .A1(n5526), .A2(n6972), .ZN(n5520) );
  INV_X1 U7158 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7045) );
  INV_X1 U7159 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6971) );
  OR2_X1 U7160 ( .A1(n5545), .A2(n6971), .ZN(n5518) );
  NOR2_X1 U7161 ( .A1(n6617), .A2(n7728), .ZN(n5523) );
  NAND2_X1 U7162 ( .A1(n5167), .A2(SI_0_), .ZN(n5522) );
  XNOR2_X1 U7163 ( .A(n5522), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9392) );
  MUX2_X1 U7164 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9392), .S(n6861), .Z(n7050) );
  INV_X1 U7165 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n8544) );
  INV_X1 U7166 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n5525) );
  INV_X1 U7167 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6837) );
  OR2_X1 U7168 ( .A1(n6081), .A2(n7728), .ZN(n5539) );
  INV_X1 U7169 ( .A(n5532), .ZN(n5534) );
  INV_X1 U7170 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5533) );
  XNOR2_X1 U7171 ( .A(n5536), .B(n5535), .ZN(n5538) );
  MUX2_X1 U7172 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n4395), .Z(n5537) );
  XNOR2_X1 U7173 ( .A(n5538), .B(n5537), .ZN(n6449) );
  XNOR2_X1 U7174 ( .A(n7729), .B(n7104), .ZN(n5540) );
  XNOR2_X1 U7175 ( .A(n5540), .B(n5539), .ZN(n6620) );
  INV_X1 U7176 ( .A(n5539), .ZN(n5542) );
  INV_X1 U7177 ( .A(n5540), .ZN(n5541) );
  NAND2_X1 U7178 ( .A1(n5542), .A2(n5541), .ZN(n5543) );
  INV_X1 U7179 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5544) );
  INV_X1 U7180 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6842) );
  OR2_X1 U7181 ( .A1(n5545), .A2(n6842), .ZN(n5546) );
  OR2_X1 U7182 ( .A1(n7108), .A2(n4796), .ZN(n5556) );
  NAND2_X1 U7183 ( .A1(n5561), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5550) );
  INV_X1 U7184 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5549) );
  OR2_X1 U7185 ( .A1(n5560), .A2(n6495), .ZN(n5553) );
  OR2_X1 U7186 ( .A1(n5941), .A2(n5249), .ZN(n5552) );
  XNOR2_X1 U7187 ( .A(n5985), .B(n7038), .ZN(n5554) );
  XNOR2_X1 U7188 ( .A(n5556), .B(n5554), .ZN(n6638) );
  INV_X1 U7189 ( .A(n5554), .ZN(n5555) );
  NOR2_X1 U7190 ( .A1(n5556), .A2(n5555), .ZN(n5557) );
  AOI21_X1 U7191 ( .B1(n6639), .B2(n6638), .A(n5557), .ZN(n6644) );
  OR2_X1 U7192 ( .A1(n5560), .A2(n6580), .ZN(n5569) );
  OR2_X1 U7193 ( .A1(n5941), .A2(n6123), .ZN(n5568) );
  OR2_X1 U7194 ( .A1(n5561), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n5563) );
  NAND2_X1 U7195 ( .A1(n5563), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5562) );
  MUX2_X1 U7196 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5562), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n5566) );
  INV_X1 U7197 ( .A(n5563), .ZN(n5565) );
  INV_X1 U7198 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5564) );
  NAND2_X1 U7199 ( .A1(n5565), .A2(n5564), .ZN(n5583) );
  NAND2_X1 U7200 ( .A1(n5566), .A2(n5583), .ZN(n8568) );
  INV_X1 U7201 ( .A(n8568), .ZN(n8573) );
  NAND2_X1 U7202 ( .A1(n6173), .A2(n8573), .ZN(n5567) );
  XNOR2_X1 U7203 ( .A(n7729), .B(n10523), .ZN(n5576) );
  NAND2_X1 U7204 ( .A1(n7743), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5574) );
  INV_X2 U7205 ( .A(n5640), .ZN(n5826) );
  INV_X1 U7206 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5570) );
  OR2_X1 U7207 ( .A1(n5826), .A2(n5570), .ZN(n5573) );
  OAI21_X1 U7208 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n5589), .ZN(n6649) );
  OR2_X1 U7209 ( .A1(n5896), .A2(n6649), .ZN(n5572) );
  INV_X1 U7210 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6843) );
  OR2_X1 U7211 ( .A1(n5900), .A2(n6843), .ZN(n5571) );
  AND4_X2 U7212 ( .A1(n5574), .A2(n5573), .A3(n5572), .A4(n5571), .ZN(n8316)
         );
  AND2_X1 U7213 ( .A1(n8527), .A2(n5575), .ZN(n5577) );
  NAND2_X1 U7214 ( .A1(n5576), .A2(n5577), .ZN(n6646) );
  NAND2_X1 U7215 ( .A1(n6644), .A2(n6646), .ZN(n5580) );
  INV_X1 U7216 ( .A(n5576), .ZN(n5579) );
  INV_X1 U7217 ( .A(n5577), .ZN(n5578) );
  NAND2_X1 U7218 ( .A1(n5579), .A2(n5578), .ZN(n6645) );
  XNOR2_X1 U7219 ( .A(n5581), .B(n5582), .ZN(n6754) );
  NAND2_X1 U7220 ( .A1(n8307), .A2(n6754), .ZN(n5587) );
  NAND2_X1 U7221 ( .A1(n5583), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5584) );
  XNOR2_X1 U7222 ( .A(n5584), .B(P2_IR_REG_5__SCAN_IN), .ZN(n8587) );
  NAND2_X1 U7223 ( .A1(n6173), .A2(n8587), .ZN(n5586) );
  INV_X1 U7224 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6141) );
  OR2_X1 U7225 ( .A1(n5941), .A2(n6141), .ZN(n5585) );
  XNOR2_X1 U7226 ( .A(n7729), .B(n7258), .ZN(n5596) );
  NAND2_X1 U7227 ( .A1(n7743), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5595) );
  INV_X1 U7228 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6846) );
  OR2_X1 U7229 ( .A1(n5900), .A2(n6846), .ZN(n5594) );
  INV_X1 U7230 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U7231 ( .A1(n5589), .A2(n5588), .ZN(n5590) );
  NAND2_X1 U7232 ( .A1(n5606), .A2(n5590), .ZN(n6116) );
  OR2_X1 U7233 ( .A1(n5896), .A2(n6116), .ZN(n5593) );
  INV_X1 U7234 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5591) );
  OR2_X1 U7235 ( .A1(n5826), .A2(n5591), .ZN(n5592) );
  AND2_X1 U7236 ( .A1(n8526), .A2(n5575), .ZN(n5597) );
  NAND2_X1 U7237 ( .A1(n5596), .A2(n5597), .ZN(n6899) );
  INV_X1 U7238 ( .A(n5596), .ZN(n5599) );
  INV_X1 U7239 ( .A(n5597), .ZN(n5598) );
  NAND2_X1 U7240 ( .A1(n5599), .A2(n5598), .ZN(n5600) );
  NAND2_X1 U7241 ( .A1(n6899), .A2(n5600), .ZN(n6115) );
  XNOR2_X1 U7242 ( .A(n5601), .B(P2_IR_REG_6__SCAN_IN), .ZN(n8600) );
  AOI22_X1 U7243 ( .A1(n8308), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6173), .B2(
        n8600), .ZN(n5604) );
  NAND2_X1 U7244 ( .A1(n6773), .A2(n8307), .ZN(n5603) );
  NAND2_X1 U7245 ( .A1(n7743), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5612) );
  INV_X1 U7246 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7268) );
  OR2_X1 U7247 ( .A1(n5900), .A2(n7268), .ZN(n5611) );
  INV_X1 U7248 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5605) );
  NAND2_X1 U7249 ( .A1(n5606), .A2(n5605), .ZN(n5607) );
  NAND2_X1 U7250 ( .A1(n5621), .A2(n5607), .ZN(n7270) );
  OR2_X1 U7251 ( .A1(n5896), .A2(n7270), .ZN(n5610) );
  INV_X1 U7252 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5608) );
  OR2_X1 U7253 ( .A1(n5826), .A2(n5608), .ZN(n5609) );
  AND2_X1 U7254 ( .A1(n8525), .A2(n5575), .ZN(n6897) );
  NAND2_X1 U7255 ( .A1(n6898), .A2(n6897), .ZN(n5613) );
  AND2_X1 U7256 ( .A1(n5613), .A2(n6899), .ZN(n5614) );
  NAND2_X1 U7257 ( .A1(n5617), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5618) );
  XNOR2_X1 U7258 ( .A(n5618), .B(P2_IR_REG_7__SCAN_IN), .ZN(n8614) );
  AOI22_X1 U7259 ( .A1(n8308), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6173), .B2(
        n8614), .ZN(n5619) );
  INV_X2 U7260 ( .A(n7729), .ZN(n5985) );
  XNOR2_X1 U7261 ( .A(n7543), .B(n5985), .ZN(n5627) );
  NAND2_X1 U7262 ( .A1(n7743), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5626) );
  INV_X1 U7263 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6851) );
  OR2_X1 U7264 ( .A1(n5900), .A2(n6851), .ZN(n5625) );
  INV_X1 U7265 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5620) );
  NAND2_X1 U7266 ( .A1(n5621), .A2(n5620), .ZN(n5622) );
  NAND2_X1 U7267 ( .A1(n5643), .A2(n5622), .ZN(n6939) );
  OR2_X1 U7268 ( .A1(n5896), .A2(n6939), .ZN(n5624) );
  INV_X1 U7269 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9248) );
  OR2_X1 U7270 ( .A1(n5826), .A2(n9248), .ZN(n5623) );
  AND4_X2 U7271 ( .A1(n5626), .A2(n5625), .A3(n5624), .A4(n5623), .ZN(n7305)
         );
  NOR2_X1 U7272 ( .A1(n7305), .A2(n4796), .ZN(n5628) );
  NAND2_X1 U7273 ( .A1(n5627), .A2(n5628), .ZN(n6979) );
  INV_X1 U7274 ( .A(n5627), .ZN(n5630) );
  INV_X1 U7275 ( .A(n5628), .ZN(n5629) );
  INV_X1 U7276 ( .A(n6898), .ZN(n5632) );
  INV_X1 U7277 ( .A(n6897), .ZN(n5631) );
  AND2_X1 U7278 ( .A1(n5632), .A2(n5631), .ZN(n6935) );
  NOR2_X1 U7279 ( .A1(n6934), .A2(n6935), .ZN(n5633) );
  NAND2_X1 U7280 ( .A1(n7171), .A2(n8307), .ZN(n5639) );
  OR2_X1 U7281 ( .A1(n5636), .A2(n9103), .ZN(n5637) );
  XNOR2_X1 U7282 ( .A(n5637), .B(P2_IR_REG_8__SCAN_IN), .ZN(n8627) );
  AOI22_X1 U7283 ( .A1(n8308), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6173), .B2(
        n8627), .ZN(n5638) );
  XNOR2_X1 U7284 ( .A(n7483), .B(n5985), .ZN(n6981) );
  NAND2_X1 U7285 ( .A1(n6182), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5648) );
  INV_X1 U7286 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7310) );
  OR2_X1 U7287 ( .A1(n5900), .A2(n7310), .ZN(n5647) );
  INV_X1 U7288 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9238) );
  OR2_X1 U7289 ( .A1(n5641), .A2(n9238), .ZN(n5646) );
  INV_X1 U7290 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5642) );
  NAND2_X1 U7291 ( .A1(n5643), .A2(n5642), .ZN(n5644) );
  NAND2_X1 U7292 ( .A1(n5656), .A2(n5644), .ZN(n7314) );
  OR2_X1 U7293 ( .A1(n5965), .A2(n7314), .ZN(n5645) );
  NOR2_X1 U7294 ( .A1(n7493), .A2(n4796), .ZN(n5663) );
  NAND2_X1 U7295 ( .A1(n6981), .A2(n5663), .ZN(n7084) );
  NAND2_X1 U7296 ( .A1(n5381), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5653) );
  XNOR2_X1 U7297 ( .A(n5653), .B(P2_IR_REG_9__SCAN_IN), .ZN(n9387) );
  AOI22_X1 U7298 ( .A1(n8308), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6173), .B2(
        n9387), .ZN(n5654) );
  XNOR2_X1 U7299 ( .A(n4746), .B(n7567), .ZN(n5668) );
  NAND2_X1 U7300 ( .A1(n7743), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5662) );
  INV_X1 U7301 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6856) );
  OR2_X1 U7302 ( .A1(n5900), .A2(n6856), .ZN(n5661) );
  INV_X1 U7303 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5655) );
  NAND2_X1 U7304 ( .A1(n5656), .A2(n5655), .ZN(n5657) );
  NAND2_X1 U7305 ( .A1(n5681), .A2(n5657), .ZN(n7565) );
  OR2_X1 U7306 ( .A1(n5965), .A2(n7565), .ZN(n5660) );
  INV_X1 U7307 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5658) );
  OR2_X1 U7308 ( .A1(n5826), .A2(n5658), .ZN(n5659) );
  OR2_X1 U7309 ( .A1(n7582), .A2(n4796), .ZN(n5669) );
  NAND2_X1 U7310 ( .A1(n5668), .A2(n5669), .ZN(n7083) );
  INV_X1 U7311 ( .A(n6981), .ZN(n5664) );
  INV_X1 U7312 ( .A(n5663), .ZN(n6980) );
  NAND2_X1 U7313 ( .A1(n5667), .A2(n5666), .ZN(n5672) );
  INV_X1 U7314 ( .A(n5668), .ZN(n5671) );
  INV_X1 U7315 ( .A(n5669), .ZN(n5670) );
  NAND2_X1 U7316 ( .A1(n5671), .A2(n5670), .ZN(n7082) );
  NAND2_X1 U7317 ( .A1(n5672), .A2(n7082), .ZN(n7053) );
  INV_X1 U7318 ( .A(n5676), .ZN(n5677) );
  NOR2_X1 U7319 ( .A1(n5381), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5718) );
  INV_X1 U7320 ( .A(n5718), .ZN(n5679) );
  NAND2_X1 U7321 ( .A1(n5679), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5702) );
  XNOR2_X1 U7322 ( .A(n5702), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6858) );
  AOI22_X1 U7323 ( .A1(n8308), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6173), .B2(
        n6858), .ZN(n5680) );
  NAND2_X1 U7324 ( .A1(n6182), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5687) );
  INV_X1 U7325 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9224) );
  OR2_X1 U7326 ( .A1(n5641), .A2(n9224), .ZN(n5686) );
  NAND2_X1 U7327 ( .A1(n5681), .A2(n9163), .ZN(n5682) );
  NAND2_X1 U7328 ( .A1(n5725), .A2(n5682), .ZN(n7643) );
  OR2_X1 U7329 ( .A1(n5896), .A2(n7643), .ZN(n5685) );
  INV_X1 U7330 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n5683) );
  OR2_X1 U7331 ( .A1(n5545), .A2(n5683), .ZN(n5684) );
  NOR2_X1 U7332 ( .A1(n7554), .A2(n4796), .ZN(n5689) );
  XNOR2_X1 U7333 ( .A(n5688), .B(n5689), .ZN(n7054) );
  INV_X1 U7334 ( .A(n5688), .ZN(n5690) );
  NAND2_X1 U7335 ( .A1(n5690), .A2(n5689), .ZN(n5691) );
  INV_X1 U7336 ( .A(n5692), .ZN(n5693) );
  NAND2_X1 U7337 ( .A1(n5694), .A2(n5693), .ZN(n5696) );
  NAND2_X1 U7338 ( .A1(n5696), .A2(n5695), .ZN(n5698) );
  NAND2_X1 U7339 ( .A1(n5698), .A2(n5697), .ZN(n5700) );
  NAND2_X1 U7340 ( .A1(n5702), .A2(n5701), .ZN(n5703) );
  NAND2_X1 U7341 ( .A1(n5703), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5704) );
  XNOR2_X1 U7342 ( .A(n5704), .B(P2_IR_REG_11__SCAN_IN), .ZN(n8660) );
  AOI22_X1 U7343 ( .A1(n8308), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6173), .B2(
        n8660), .ZN(n5705) );
  INV_X1 U7344 ( .A(n5705), .ZN(n5706) );
  XNOR2_X1 U7345 ( .A(n4746), .B(n7561), .ZN(n5714) );
  NAND2_X1 U7346 ( .A1(n7743), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5711) );
  INV_X1 U7347 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7558) );
  OR2_X1 U7348 ( .A1(n5900), .A2(n7558), .ZN(n5710) );
  INV_X1 U7349 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5724) );
  XNOR2_X1 U7350 ( .A(n5725), .B(n5724), .ZN(n7560) );
  OR2_X1 U7351 ( .A1(n5896), .A2(n7560), .ZN(n5709) );
  INV_X1 U7352 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n5707) );
  OR2_X1 U7353 ( .A1(n5826), .A2(n5707), .ZN(n5708) );
  NAND4_X1 U7354 ( .A1(n5711), .A2(n5710), .A3(n5709), .A4(n5708), .ZN(n8520)
         );
  NAND2_X1 U7355 ( .A1(n8520), .A2(n5575), .ZN(n5712) );
  XNOR2_X1 U7356 ( .A(n5714), .B(n5712), .ZN(n7139) );
  INV_X1 U7357 ( .A(n5712), .ZN(n5713) );
  NAND2_X1 U7358 ( .A1(n5714), .A2(n5713), .ZN(n5715) );
  NAND2_X1 U7359 ( .A1(n7385), .A2(n8307), .ZN(n5721) );
  NOR2_X1 U7360 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5717) );
  NAND2_X1 U7361 ( .A1(n5718), .A2(n5717), .ZN(n5738) );
  NAND2_X1 U7362 ( .A1(n5738), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5719) );
  XNOR2_X1 U7363 ( .A(n5719), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6918) );
  AOI22_X1 U7364 ( .A1(n8308), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6173), .B2(
        n6918), .ZN(n5720) );
  XNOR2_X1 U7365 ( .A(n4746), .B(n9067), .ZN(n5732) );
  NAND2_X1 U7366 ( .A1(n6182), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5731) );
  INV_X1 U7367 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n5722) );
  OR2_X1 U7368 ( .A1(n5641), .A2(n5722), .ZN(n5730) );
  INV_X1 U7369 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5723) );
  OAI21_X1 U7370 ( .B1(n5725), .B2(n5724), .A(n5723), .ZN(n5726) );
  NAND2_X1 U7371 ( .A1(n5726), .A2(n5741), .ZN(n7333) );
  OR2_X1 U7372 ( .A1(n5965), .A2(n7333), .ZN(n5729) );
  INV_X1 U7373 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n5727) );
  OR2_X1 U7374 ( .A1(n5545), .A2(n5727), .ZN(n5728) );
  NOR2_X1 U7375 ( .A1(n7626), .A2(n4796), .ZN(n5733) );
  XNOR2_X1 U7376 ( .A(n5732), .B(n5733), .ZN(n7332) );
  INV_X1 U7377 ( .A(n5732), .ZN(n5734) );
  NAND2_X1 U7378 ( .A1(n5734), .A2(n5733), .ZN(n5735) );
  NAND2_X1 U7379 ( .A1(n5736), .A2(n5735), .ZN(n7515) );
  XNOR2_X1 U7380 ( .A(n5737), .B(n5325), .ZN(n7799) );
  NAND2_X1 U7381 ( .A1(n5792), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5754) );
  XNOR2_X1 U7382 ( .A(n5754), .B(P2_IR_REG_13__SCAN_IN), .ZN(n6883) );
  AOI22_X1 U7383 ( .A1(n8308), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6173), .B2(
        n6883), .ZN(n5739) );
  XNOR2_X1 U7384 ( .A(n4746), .B(n8407), .ZN(n5747) );
  NAND2_X1 U7385 ( .A1(n8288), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5746) );
  INV_X1 U7386 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6819) );
  OR2_X1 U7387 ( .A1(n5641), .A2(n6819), .ZN(n5745) );
  INV_X1 U7388 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5740) );
  NAND2_X1 U7389 ( .A1(n5741), .A2(n5740), .ZN(n5742) );
  NAND2_X1 U7390 ( .A1(n5762), .A2(n5742), .ZN(n7637) );
  OR2_X1 U7391 ( .A1(n5896), .A2(n7637), .ZN(n5744) );
  INV_X1 U7392 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9293) );
  OR2_X1 U7393 ( .A1(n5826), .A2(n9293), .ZN(n5743) );
  NOR2_X1 U7394 ( .A1(n8156), .A2(n4796), .ZN(n5748) );
  INV_X1 U7395 ( .A(n5747), .ZN(n5749) );
  NAND2_X1 U7396 ( .A1(n5749), .A2(n5748), .ZN(n5750) );
  NAND2_X1 U7397 ( .A1(n7804), .A2(n8307), .ZN(n5760) );
  INV_X1 U7398 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5753) );
  NAND2_X1 U7399 ( .A1(n5754), .A2(n5753), .ZN(n5755) );
  NAND2_X1 U7400 ( .A1(n5755), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5757) );
  NAND2_X1 U7401 ( .A1(n5757), .A2(n5756), .ZN(n5776) );
  OR2_X1 U7402 ( .A1(n5757), .A2(n5756), .ZN(n5758) );
  AOI22_X1 U7403 ( .A1(n7015), .A2(n6173), .B1(n8308), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n5759) );
  XNOR2_X1 U7404 ( .A(n4746), .B(n9054), .ZN(n5768) );
  NAND2_X1 U7405 ( .A1(n6182), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5767) );
  INV_X1 U7406 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n6880) );
  OR2_X1 U7407 ( .A1(n5641), .A2(n6880), .ZN(n5766) );
  INV_X1 U7408 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6887) );
  OR2_X1 U7409 ( .A1(n5900), .A2(n6887), .ZN(n5765) );
  INV_X1 U7410 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5761) );
  NAND2_X1 U7411 ( .A1(n5762), .A2(n5761), .ZN(n5763) );
  NAND2_X1 U7412 ( .A1(n5781), .A2(n5763), .ZN(n8157) );
  OR2_X1 U7413 ( .A1(n5965), .A2(n8157), .ZN(n5764) );
  OR2_X1 U7414 ( .A1(n7700), .A2(n4796), .ZN(n5769) );
  NAND2_X1 U7415 ( .A1(n5768), .A2(n5769), .ZN(n5773) );
  INV_X1 U7416 ( .A(n5768), .ZN(n5771) );
  INV_X1 U7417 ( .A(n5769), .ZN(n5770) );
  NAND2_X1 U7418 ( .A1(n5771), .A2(n5770), .ZN(n5772) );
  NAND2_X1 U7419 ( .A1(n5773), .A2(n5772), .ZN(n8154) );
  XNOR2_X1 U7420 ( .A(n5775), .B(n5774), .ZN(n7819) );
  NAND2_X1 U7421 ( .A1(n7819), .A2(n8307), .ZN(n5779) );
  NAND2_X1 U7422 ( .A1(n5776), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5777) );
  XNOR2_X1 U7423 ( .A(n5777), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7503) );
  AOI22_X1 U7424 ( .A1(n7503), .A2(n6173), .B1(n8308), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5778) );
  XNOR2_X1 U7425 ( .A(n4746), .B(n9049), .ZN(n8199) );
  NAND2_X1 U7426 ( .A1(n5781), .A2(n5780), .ZN(n5782) );
  AND2_X1 U7427 ( .A1(n5804), .A2(n5782), .ZN(n8272) );
  NAND2_X1 U7428 ( .A1(n7747), .A2(n8272), .ZN(n5788) );
  INV_X1 U7429 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7019) );
  OR2_X1 U7430 ( .A1(n5641), .A2(n7019), .ZN(n5787) );
  INV_X1 U7431 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n5783) );
  OR2_X1 U7432 ( .A1(n5826), .A2(n5783), .ZN(n5786) );
  INV_X1 U7433 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n5784) );
  OR2_X1 U7434 ( .A1(n5545), .A2(n5784), .ZN(n5785) );
  OR2_X1 U7435 ( .A1(n8925), .A2(n4796), .ZN(n5809) );
  NAND2_X1 U7436 ( .A1(n7832), .A2(n8307), .ZN(n5799) );
  INV_X1 U7437 ( .A(n5790), .ZN(n5791) );
  NAND2_X1 U7438 ( .A1(n5794), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5793) );
  MUX2_X1 U7439 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5793), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n5797) );
  INV_X1 U7440 ( .A(n5794), .ZN(n5796) );
  NAND2_X1 U7441 ( .A1(n5796), .A2(n5795), .ZN(n5820) );
  NAND2_X1 U7442 ( .A1(n5797), .A2(n5820), .ZN(n7607) );
  INV_X1 U7443 ( .A(n7607), .ZN(n7603) );
  AOI22_X1 U7444 ( .A1(n7603), .A2(n6173), .B1(n8308), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n5798) );
  XNOR2_X1 U7445 ( .A(n8942), .B(n5985), .ZN(n5814) );
  INV_X1 U7446 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n5800) );
  OR2_X1 U7447 ( .A1(n5641), .A2(n5800), .ZN(n5802) );
  INV_X1 U7448 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8939) );
  OR2_X1 U7449 ( .A1(n5900), .A2(n8939), .ZN(n5801) );
  AND2_X1 U7450 ( .A1(n5802), .A2(n5801), .ZN(n5808) );
  INV_X1 U7451 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5803) );
  NAND2_X1 U7452 ( .A1(n5804), .A2(n5803), .ZN(n5805) );
  NAND2_X1 U7453 ( .A1(n5824), .A2(n5805), .ZN(n8938) );
  OR2_X1 U7454 ( .A1(n8938), .A2(n5896), .ZN(n5807) );
  NAND2_X1 U7455 ( .A1(n6182), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5806) );
  INV_X1 U7456 ( .A(n8278), .ZN(n8515) );
  NAND2_X1 U7457 ( .A1(n8515), .A2(n5575), .ZN(n5815) );
  XNOR2_X1 U7458 ( .A(n5814), .B(n5815), .ZN(n8202) );
  INV_X1 U7459 ( .A(n8199), .ZN(n5810) );
  INV_X1 U7460 ( .A(n5809), .ZN(n8271) );
  NAND2_X1 U7461 ( .A1(n5810), .A2(n8271), .ZN(n5811) );
  AND2_X1 U7462 ( .A1(n8202), .A2(n5811), .ZN(n5812) );
  INV_X1 U7463 ( .A(n5814), .ZN(n5816) );
  NAND2_X1 U7464 ( .A1(n5816), .A2(n5815), .ZN(n5817) );
  XNOR2_X1 U7465 ( .A(n5819), .B(n5818), .ZN(n7841) );
  NAND2_X1 U7466 ( .A1(n7841), .A2(n8307), .ZN(n5823) );
  NAND2_X1 U7467 ( .A1(n5820), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5821) );
  XNOR2_X1 U7468 ( .A(n5821), .B(P2_IR_REG_17__SCAN_IN), .ZN(n7672) );
  AOI22_X1 U7469 ( .A1(n7672), .A2(n6173), .B1(n8308), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n5822) );
  XNOR2_X1 U7470 ( .A(n9037), .B(n5985), .ZN(n5831) );
  INV_X1 U7471 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n7612) );
  NAND2_X1 U7472 ( .A1(n5824), .A2(n7612), .ZN(n5825) );
  NAND2_X1 U7473 ( .A1(n5840), .A2(n5825), .ZN(n8916) );
  OR2_X1 U7474 ( .A1(n8916), .A2(n5896), .ZN(n5829) );
  AOI22_X1 U7475 ( .A1(n8288), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n7743), .B2(
        P2_REG1_REG_17__SCAN_IN), .ZN(n5828) );
  INV_X1 U7476 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9175) );
  OR2_X1 U7477 ( .A1(n5826), .A2(n9175), .ZN(n5827) );
  NOR2_X1 U7478 ( .A1(n8927), .A2(n4796), .ZN(n5830) );
  XNOR2_X1 U7479 ( .A(n5831), .B(n5830), .ZN(n8212) );
  NAND2_X1 U7480 ( .A1(n5831), .A2(n5830), .ZN(n5832) );
  XNOR2_X1 U7481 ( .A(n5835), .B(n5834), .ZN(n7848) );
  NAND2_X1 U7482 ( .A1(n7848), .A2(n8307), .ZN(n5838) );
  XNOR2_X1 U7483 ( .A(n5836), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8670) );
  AOI22_X1 U7484 ( .A1(n8308), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6173), .B2(
        n8670), .ZN(n5837) );
  XNOR2_X1 U7485 ( .A(n4746), .B(n9032), .ZN(n5845) );
  NAND2_X1 U7486 ( .A1(n5840), .A2(n5839), .ZN(n5841) );
  AND2_X1 U7487 ( .A1(n5854), .A2(n5841), .ZN(n8253) );
  NAND2_X1 U7488 ( .A1(n8253), .A2(n7747), .ZN(n5844) );
  AOI22_X1 U7489 ( .A1(n7743), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n6182), .B2(
        P2_REG0_REG_18__SCAN_IN), .ZN(n5843) );
  NAND2_X1 U7490 ( .A1(n8288), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5842) );
  NOR2_X1 U7491 ( .A1(n8214), .A2(n4796), .ZN(n5846) );
  XNOR2_X1 U7492 ( .A(n5845), .B(n5846), .ZN(n8250) );
  INV_X1 U7493 ( .A(n5845), .ZN(n5847) );
  NAND2_X1 U7494 ( .A1(n5847), .A2(n5846), .ZN(n5848) );
  XNOR2_X1 U7495 ( .A(n5850), .B(n5849), .ZN(n7857) );
  NAND2_X1 U7496 ( .A1(n7857), .A2(n8307), .ZN(n5852) );
  AOI22_X1 U7497 ( .A1(n8308), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8340), .B2(
        n6173), .ZN(n5851) );
  XNOR2_X1 U7498 ( .A(n4746), .B(n9028), .ZN(n5861) );
  INV_X1 U7499 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5853) );
  NAND2_X1 U7500 ( .A1(n5854), .A2(n5853), .ZN(n5855) );
  NAND2_X1 U7501 ( .A1(n5881), .A2(n5855), .ZN(n8870) );
  OR2_X1 U7502 ( .A1(n8870), .A2(n5965), .ZN(n5860) );
  INV_X1 U7503 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9185) );
  NAND2_X1 U7504 ( .A1(n8288), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5857) );
  NAND2_X1 U7505 ( .A1(n6182), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5856) );
  OAI211_X1 U7506 ( .C1(n5641), .C2(n9185), .A(n5857), .B(n5856), .ZN(n5858)
         );
  INV_X1 U7507 ( .A(n5858), .ZN(n5859) );
  NAND2_X1 U7508 ( .A1(n8889), .A2(n5575), .ZN(n5862) );
  NAND2_X1 U7509 ( .A1(n5861), .A2(n5862), .ZN(n5867) );
  INV_X1 U7510 ( .A(n5861), .ZN(n5864) );
  INV_X1 U7511 ( .A(n5862), .ZN(n5863) );
  NAND2_X1 U7512 ( .A1(n5864), .A2(n5863), .ZN(n5865) );
  NAND2_X1 U7513 ( .A1(n5867), .A2(n5865), .ZN(n8174) );
  INV_X1 U7514 ( .A(n8174), .ZN(n5866) );
  XNOR2_X1 U7515 ( .A(n5869), .B(n5868), .ZN(n7867) );
  NAND2_X1 U7516 ( .A1(n7867), .A2(n8307), .ZN(n5871) );
  OR2_X1 U7517 ( .A1(n5941), .A2(n9374), .ZN(n5870) );
  XNOR2_X1 U7518 ( .A(n9022), .B(n5985), .ZN(n5876) );
  XNOR2_X1 U7519 ( .A(n5881), .B(P2_REG3_REG_20__SCAN_IN), .ZN(n8853) );
  INV_X1 U7520 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n5874) );
  NAND2_X1 U7521 ( .A1(n7743), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5873) );
  NAND2_X1 U7522 ( .A1(n6182), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5872) );
  OAI211_X1 U7523 ( .C1(n5545), .C2(n5874), .A(n5873), .B(n5872), .ZN(n5875)
         );
  AOI21_X1 U7524 ( .B1(n8853), .B2(n7747), .A(n5875), .ZN(n8182) );
  NOR2_X1 U7525 ( .A1(n8182), .A2(n4796), .ZN(n5877) );
  XNOR2_X1 U7526 ( .A(n5876), .B(n5877), .ZN(n8232) );
  XNOR2_X1 U7527 ( .A(n5878), .B(n4500), .ZN(n7880) );
  NAND2_X1 U7528 ( .A1(n7880), .A2(n8307), .ZN(n5880) );
  NAND2_X1 U7529 ( .A1(n8308), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5879) );
  XNOR2_X1 U7530 ( .A(n9015), .B(n5985), .ZN(n5908) );
  INV_X1 U7531 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8234) );
  INV_X1 U7532 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8181) );
  OAI21_X1 U7533 ( .B1(n5881), .B2(n8234), .A(n8181), .ZN(n5883) );
  INV_X1 U7534 ( .A(n5882), .ZN(n5894) );
  NAND2_X1 U7535 ( .A1(n8834), .A2(n7747), .ZN(n5889) );
  INV_X1 U7536 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n5886) );
  NAND2_X1 U7537 ( .A1(n7743), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5885) );
  NAND2_X1 U7538 ( .A1(n6182), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5884) );
  OAI211_X1 U7539 ( .C1(n5900), .C2(n5886), .A(n5885), .B(n5884), .ZN(n5887)
         );
  INV_X1 U7540 ( .A(n5887), .ZN(n5888) );
  NAND2_X1 U7541 ( .A1(n8513), .A2(n5575), .ZN(n5904) );
  XNOR2_X1 U7542 ( .A(n5908), .B(n5904), .ZN(n8179) );
  XNOR2_X1 U7543 ( .A(n5891), .B(n5890), .ZN(n7893) );
  NAND2_X1 U7544 ( .A1(n7893), .A2(n8307), .ZN(n5893) );
  NAND2_X1 U7545 ( .A1(n8308), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5892) );
  XNOR2_X1 U7546 ( .A(n9010), .B(n5985), .ZN(n5906) );
  INV_X1 U7547 ( .A(n5906), .ZN(n8243) );
  INV_X1 U7548 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9325) );
  NAND2_X1 U7549 ( .A1(n5894), .A2(n9325), .ZN(n5895) );
  NAND2_X1 U7550 ( .A1(n5919), .A2(n5895), .ZN(n8817) );
  OR2_X1 U7551 ( .A1(n8817), .A2(n5896), .ZN(n5903) );
  INV_X1 U7552 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n5899) );
  NAND2_X1 U7553 ( .A1(n6182), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5898) );
  NAND2_X1 U7554 ( .A1(n7743), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5897) );
  OAI211_X1 U7555 ( .C1(n5900), .C2(n5899), .A(n5898), .B(n5897), .ZN(n5901)
         );
  INV_X1 U7556 ( .A(n5901), .ZN(n5902) );
  NAND2_X1 U7557 ( .A1(n8841), .A2(n5575), .ZN(n8242) );
  NAND2_X1 U7558 ( .A1(n8243), .A2(n8242), .ZN(n5911) );
  INV_X1 U7559 ( .A(n5904), .ZN(n5907) );
  NAND2_X1 U7560 ( .A1(n5908), .A2(n5907), .ZN(n8240) );
  NAND2_X1 U7561 ( .A1(n8240), .A2(n8242), .ZN(n5905) );
  NAND2_X1 U7562 ( .A1(n5906), .A2(n5905), .ZN(n5910) );
  NAND3_X1 U7563 ( .A1(n5908), .A2(n5907), .A3(n8841), .ZN(n5909) );
  XNOR2_X1 U7564 ( .A(n5913), .B(n5912), .ZN(n7899) );
  NAND2_X1 U7565 ( .A1(n7899), .A2(n8307), .ZN(n5915) );
  NAND2_X1 U7566 ( .A1(n8308), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5914) );
  XNOR2_X1 U7567 ( .A(n4746), .B(n9005), .ZN(n5917) );
  NAND2_X1 U7568 ( .A1(n5919), .A2(n8166), .ZN(n5920) );
  NAND2_X1 U7569 ( .A1(n5921), .A2(n5920), .ZN(n8807) );
  OR2_X1 U7570 ( .A1(n8807), .A2(n5965), .ZN(n5927) );
  INV_X1 U7571 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n5924) );
  NAND2_X1 U7572 ( .A1(n6182), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5923) );
  NAND2_X1 U7573 ( .A1(n7743), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5922) );
  OAI211_X1 U7574 ( .C1(n5545), .C2(n5924), .A(n5923), .B(n5922), .ZN(n5925)
         );
  INV_X1 U7575 ( .A(n5925), .ZN(n5926) );
  NOR2_X1 U7576 ( .A1(n8824), .A2(n4796), .ZN(n8164) );
  INV_X1 U7577 ( .A(n5932), .ZN(n5933) );
  NAND2_X1 U7578 ( .A1(n5933), .A2(SI_24_), .ZN(n5934) );
  INV_X1 U7579 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7925) );
  MUX2_X1 U7580 ( .A(n9253), .B(n7925), .S(n4396), .Z(n5938) );
  INV_X1 U7581 ( .A(SI_25_), .ZN(n5937) );
  NAND2_X1 U7582 ( .A1(n5938), .A2(n5937), .ZN(n5955) );
  INV_X1 U7583 ( .A(n5938), .ZN(n5939) );
  NAND2_X1 U7584 ( .A1(n5939), .A2(SI_25_), .ZN(n5940) );
  NAND2_X1 U7585 ( .A1(n5955), .A2(n5940), .ZN(n5953) );
  NAND2_X1 U7586 ( .A1(n7924), .A2(n8307), .ZN(n5943) );
  OR2_X1 U7587 ( .A1(n5941), .A2(n9253), .ZN(n5942) );
  INV_X1 U7588 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5944) );
  NAND2_X1 U7589 ( .A1(n5945), .A2(n5944), .ZN(n5946) );
  INV_X1 U7590 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n5949) );
  NAND2_X1 U7591 ( .A1(n6182), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5948) );
  NAND2_X1 U7592 ( .A1(n7743), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5947) );
  OAI211_X1 U7593 ( .C1(n5545), .C2(n5949), .A(n5948), .B(n5947), .ZN(n5950)
         );
  AOI21_X2 U7594 ( .B1(n8762), .B2(n7747), .A(n5950), .ZN(n8741) );
  NOR2_X1 U7595 ( .A1(n8741), .A2(n4796), .ZN(n8188) );
  INV_X1 U7596 ( .A(n8189), .ZN(n5951) );
  INV_X1 U7597 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9119) );
  INV_X1 U7598 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n10352) );
  MUX2_X1 U7599 ( .A(n9119), .B(n10352), .S(n4397), .Z(n5957) );
  INV_X1 U7600 ( .A(SI_26_), .ZN(n5956) );
  NAND2_X1 U7601 ( .A1(n5957), .A2(n5956), .ZN(n5977) );
  INV_X1 U7602 ( .A(n5957), .ZN(n5958) );
  NAND2_X1 U7603 ( .A1(n5958), .A2(SI_26_), .ZN(n5959) );
  NAND2_X1 U7604 ( .A1(n9117), .A2(n8307), .ZN(n5961) );
  NAND2_X1 U7605 ( .A1(n8308), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5960) );
  XNOR2_X1 U7606 ( .A(n4746), .B(n8746), .ZN(n5972) );
  INV_X1 U7607 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9254) );
  NAND2_X1 U7608 ( .A1(n5963), .A2(n9254), .ZN(n5964) );
  NAND2_X1 U7609 ( .A1(n6037), .A2(n5964), .ZN(n8262) );
  INV_X1 U7610 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9327) );
  NAND2_X1 U7611 ( .A1(n8288), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5967) );
  INV_X1 U7612 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9240) );
  OR2_X1 U7613 ( .A1(n5826), .A2(n9240), .ZN(n5966) );
  OAI211_X1 U7614 ( .C1(n5641), .C2(n9327), .A(n5967), .B(n5966), .ZN(n5968)
         );
  INV_X1 U7615 ( .A(n5968), .ZN(n5969) );
  NAND2_X1 U7616 ( .A1(n8727), .A2(n5575), .ZN(n5971) );
  NOR2_X1 U7617 ( .A1(n5972), .A2(n5971), .ZN(n5973) );
  AOI21_X1 U7618 ( .B1(n5972), .B2(n5971), .A(n5973), .ZN(n8260) );
  INV_X1 U7619 ( .A(n5973), .ZN(n5974) );
  INV_X1 U7620 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5979) );
  INV_X1 U7621 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9351) );
  MUX2_X1 U7622 ( .A(n5979), .B(n9351), .S(n4394), .Z(n5980) );
  INV_X1 U7623 ( .A(SI_27_), .ZN(n9297) );
  NAND2_X1 U7624 ( .A1(n5980), .A2(n9297), .ZN(n7712) );
  INV_X1 U7625 ( .A(n5980), .ZN(n5981) );
  NAND2_X1 U7626 ( .A1(n5981), .A2(SI_27_), .ZN(n5982) );
  NAND2_X1 U7627 ( .A1(n9114), .A2(n8307), .ZN(n5984) );
  NAND2_X1 U7628 ( .A1(n8308), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5983) );
  XNOR2_X1 U7629 ( .A(n8984), .B(n5985), .ZN(n5992) );
  INV_X1 U7630 ( .A(n5992), .ZN(n5994) );
  XNOR2_X1 U7631 ( .A(n6037), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8722) );
  NAND2_X1 U7632 ( .A1(n8722), .A2(n7747), .ZN(n5990) );
  INV_X1 U7633 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9356) );
  NAND2_X1 U7634 ( .A1(n6182), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5987) );
  NAND2_X1 U7635 ( .A1(n8288), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5986) );
  OAI211_X1 U7636 ( .C1(n5641), .C2(n9356), .A(n5987), .B(n5986), .ZN(n5988)
         );
  INV_X1 U7637 ( .A(n5988), .ZN(n5989) );
  AND2_X2 U7638 ( .A1(n5990), .A2(n5989), .ZN(n8742) );
  NOR2_X1 U7639 ( .A1(n8742), .A2(n4796), .ZN(n5991) );
  INV_X1 U7640 ( .A(n5991), .ZN(n5993) );
  INV_X1 U7641 ( .A(n5995), .ZN(n5998) );
  NAND2_X1 U7642 ( .A1(n5998), .A2(n5997), .ZN(n6026) );
  NOR2_X1 U7643 ( .A1(n5999), .A2(n9103), .ZN(n6000) );
  MUX2_X1 U7644 ( .A(n9103), .B(n6000), .S(P2_IR_REG_25__SCAN_IN), .Z(n6001)
         );
  INV_X1 U7645 ( .A(n6001), .ZN(n6003) );
  NAND2_X1 U7646 ( .A1(n6003), .A2(n6002), .ZN(n7653) );
  NAND2_X1 U7647 ( .A1(n6005), .A2(n6004), .ZN(n6006) );
  INV_X1 U7648 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U7649 ( .A1(n6024), .A2(n6023), .ZN(n6007) );
  NAND2_X1 U7650 ( .A1(n6007), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6009) );
  INV_X1 U7651 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6008) );
  XNOR2_X1 U7652 ( .A(n7528), .B(P2_B_REG_SCAN_IN), .ZN(n6013) );
  NAND2_X1 U7653 ( .A1(n6002), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6010) );
  MUX2_X1 U7654 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6010), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6012) );
  NAND2_X1 U7655 ( .A1(n6012), .A2(n6011), .ZN(n9122) );
  INV_X1 U7656 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10509) );
  AND2_X1 U7657 ( .A1(n7528), .A2(n9122), .ZN(n10510) );
  AOI21_X1 U7658 ( .B1(n10500), .B2(n10509), .A(n10510), .ZN(n6729) );
  NOR4_X1 U7659 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6017) );
  NOR4_X1 U7660 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n6016) );
  NOR4_X1 U7661 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n6015) );
  NOR4_X1 U7662 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n6014) );
  NAND4_X1 U7663 ( .A1(n6017), .A2(n6016), .A3(n6015), .A4(n6014), .ZN(n6022)
         );
  NOR2_X1 U7664 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .ZN(
        n9133) );
  NOR4_X1 U7665 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6020) );
  NOR4_X1 U7666 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6019) );
  NOR4_X1 U7667 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n6018) );
  NAND4_X1 U7668 ( .A1(n9133), .A2(n6020), .A3(n6019), .A4(n6018), .ZN(n6021)
         );
  OAI21_X1 U7669 ( .B1(n6022), .B2(n6021), .A(n10500), .ZN(n6727) );
  AND2_X1 U7670 ( .A1(n6729), .A2(n6727), .ZN(n6485) );
  INV_X1 U7671 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10512) );
  AND2_X1 U7672 ( .A1(n7653), .A2(n9122), .ZN(n10513) );
  AOI21_X1 U7673 ( .B1(n10512), .B2(n10500), .A(n10513), .ZN(n6484) );
  NAND2_X1 U7674 ( .A1(n6485), .A2(n6484), .ZN(n7732) );
  XNOR2_X1 U7675 ( .A(n6024), .B(n6023), .ZN(n6172) );
  NAND2_X1 U7676 ( .A1(n6025), .A2(n8915), .ZN(n6032) );
  OR3_X1 U7677 ( .A1(n10501), .A2(n6814), .A3(n9074), .ZN(n7731) );
  AND2_X1 U7678 ( .A1(n8340), .A2(n8339), .ZN(n6027) );
  NAND2_X1 U7679 ( .A1(n6025), .A2(n6027), .ZN(n9047) );
  NAND2_X1 U7680 ( .A1(n7732), .A2(n6482), .ZN(n6604) );
  NOR2_X1 U7681 ( .A1(n10501), .A2(n10528), .ZN(n6028) );
  AND2_X1 U7682 ( .A1(n6032), .A2(n6814), .ZN(n6086) );
  INV_X1 U7683 ( .A(n6086), .ZN(n6029) );
  AND3_X1 U7684 ( .A1(n6029), .A2(n6815), .A3(n6172), .ZN(n6030) );
  NAND2_X1 U7685 ( .A1(n6604), .A2(n6030), .ZN(n6031) );
  INV_X1 U7686 ( .A(n7732), .ZN(n6033) );
  NOR2_X1 U7687 ( .A1(n10501), .A2(n6032), .ZN(n8502) );
  INV_X1 U7688 ( .A(n6034), .ZN(n6035) );
  NOR2_X1 U7689 ( .A1(n8193), .A2(n8263), .ZN(n6044) );
  INV_X1 U7690 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6042) );
  INV_X1 U7691 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6036) );
  OAI21_X1 U7692 ( .B1(n6037), .B2(n6042), .A(n6036), .ZN(n6038) );
  INV_X1 U7693 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9226) );
  NAND2_X1 U7694 ( .A1(n8288), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6040) );
  NAND2_X1 U7695 ( .A1(n7743), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6039) );
  OAI211_X1 U7696 ( .C1(n9226), .C2(n5826), .A(n6040), .B(n6039), .ZN(n6041)
         );
  NAND2_X1 U7697 ( .A1(n6814), .A2(n6034), .ZN(n8926) );
  OAI22_X1 U7698 ( .A1(n8710), .A2(n8277), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6042), .ZN(n6043) );
  AOI211_X1 U7699 ( .C1(n8273), .C2(n8722), .A(n6044), .B(n6043), .ZN(n6045)
         );
  INV_X1 U7700 ( .A(n6046), .ZN(n6047) );
  NAND4_X1 U7701 ( .A1(n6065), .A2(n6053), .A3(n6052), .A4(n6051), .ZN(n6054)
         );
  NAND2_X1 U7702 ( .A1(n6058), .A2(n6059), .ZN(n6055) );
  INV_X1 U7703 ( .A(n6132), .ZN(n6061) );
  XNOR2_X1 U7704 ( .A(n6057), .B(n6056), .ZN(n7654) );
  XNOR2_X1 U7705 ( .A(n6058), .B(n6059), .ZN(n7525) );
  NAND2_X2 U7706 ( .A1(n6061), .A2(n6060), .ZN(n6520) );
  NAND2_X1 U7707 ( .A1(n4501), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6063) );
  XNOR2_X1 U7708 ( .A(n6063), .B(n6062), .ZN(n6519) );
  INV_X1 U7709 ( .A(n6519), .ZN(n7342) );
  NOR2_X1 U7710 ( .A1(n6520), .A2(n7342), .ZN(n6199) );
  AND2_X1 U7711 ( .A1(n6305), .A2(n6065), .ZN(n6066) );
  NAND2_X1 U7712 ( .A1(n6071), .A2(n6070), .ZN(n6067) );
  NAND2_X1 U7713 ( .A1(n6067), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6069) );
  INV_X1 U7714 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6068) );
  OR2_X1 U7715 ( .A1(n6667), .A2(n6393), .ZN(n6072) );
  NAND2_X1 U7716 ( .A1(n6072), .A2(n6519), .ZN(n6211) );
  NAND2_X1 U7717 ( .A1(n6079), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X2 U7718 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U7719 ( .A(n6815), .ZN(n6080) );
  NAND2_X2 U7720 ( .A1(n6080), .A2(n10514), .ZN(n8514) );
  NAND2_X1 U7721 ( .A1(n6605), .A2(n8362), .ZN(n8353) );
  NAND2_X2 U7722 ( .A1(n8528), .A2(n5254), .ZN(n8361) );
  NAND2_X1 U7723 ( .A1(n8353), .A2(n8361), .ZN(n7100) );
  INV_X1 U7724 ( .A(n7100), .ZN(n6082) );
  INV_X1 U7725 ( .A(n6081), .ZN(n6611) );
  NAND2_X1 U7726 ( .A1(n6081), .A2(n7104), .ZN(n8363) );
  INV_X1 U7727 ( .A(n7030), .ZN(n6092) );
  NAND2_X1 U7728 ( .A1(n6082), .A2(n6092), .ZN(n7098) );
  INV_X1 U7729 ( .A(n7108), .ZN(n6622) );
  NAND2_X1 U7730 ( .A1(n8527), .A2(n10523), .ZN(n7297) );
  AND2_X1 U7731 ( .A1(n7298), .A2(n7297), .ZN(n7262) );
  NOR2_X1 U7732 ( .A1(n8526), .A2(n7258), .ZN(n7299) );
  INV_X1 U7733 ( .A(n7299), .ZN(n8347) );
  NAND2_X1 U7734 ( .A1(n8347), .A2(n8370), .ZN(n7261) );
  INV_X1 U7735 ( .A(n7261), .ZN(n6095) );
  XNOR2_X1 U7736 ( .A(n7262), .B(n6095), .ZN(n6083) );
  INV_X1 U7737 ( .A(n6025), .ZN(n8497) );
  NAND2_X1 U7738 ( .A1(n8497), .A2(n8350), .ZN(n8314) );
  NAND2_X1 U7739 ( .A1(n6083), .A2(n8935), .ZN(n6085) );
  AOI22_X1 U7740 ( .A1(n8886), .A2(n8527), .B1(n8525), .B2(n8888), .ZN(n6084)
         );
  NAND2_X1 U7741 ( .A1(n6085), .A2(n6084), .ZN(n7075) );
  INV_X1 U7742 ( .A(n6729), .ZN(n6088) );
  NOR2_X1 U7743 ( .A1(n10501), .A2(n6086), .ZN(n6603) );
  AND2_X1 U7744 ( .A1(n6727), .A2(n6603), .ZN(n6087) );
  NAND3_X1 U7745 ( .A1(n6088), .A2(n6484), .A3(n6087), .ZN(n7048) );
  MUX2_X1 U7746 ( .A(n7075), .B(P2_REG2_REG_5__SCAN_IN), .S(n8958), .Z(n6112)
         );
  INV_X1 U7747 ( .A(n7050), .ZN(n6487) );
  NOR2_X1 U7748 ( .A1(n6617), .A2(n6487), .ZN(n6734) );
  INV_X1 U7749 ( .A(n6734), .ZN(n6089) );
  NAND2_X1 U7750 ( .A1(n6081), .A2(n10518), .ZN(n7027) );
  NAND2_X1 U7751 ( .A1(n6090), .A2(n5254), .ZN(n7029) );
  AND2_X1 U7752 ( .A1(n7027), .A2(n7029), .ZN(n6091) );
  NAND2_X1 U7753 ( .A1(n6092), .A2(n7027), .ZN(n6093) );
  NAND2_X1 U7754 ( .A1(n7108), .A2(n6094), .ZN(n6096) );
  NAND2_X1 U7755 ( .A1(n6098), .A2(n6096), .ZN(n7111) );
  NAND2_X1 U7756 ( .A1(n7111), .A2(n7110), .ZN(n7109) );
  NAND3_X1 U7757 ( .A1(n7109), .A2(n6095), .A3(n6097), .ZN(n6101) );
  NAND2_X1 U7758 ( .A1(n6101), .A2(n7290), .ZN(n7077) );
  XNOR2_X1 U7759 ( .A(n6102), .B(n8504), .ZN(n8910) );
  NAND2_X1 U7760 ( .A1(n8910), .A2(n8915), .ZN(n8931) );
  OR2_X1 U7761 ( .A1(n6102), .A2(n8915), .ZN(n7161) );
  NAND2_X1 U7762 ( .A1(n8931), .A2(n7161), .ZN(n6103) );
  AND2_X1 U7763 ( .A1(n7077), .A2(n8953), .ZN(n6111) );
  OR2_X1 U7764 ( .A1(n8949), .A2(n8340), .ZN(n8759) );
  OAI21_X1 U7765 ( .B1(n7113), .B2(n7258), .A(n9075), .ZN(n6106) );
  OR2_X1 U7766 ( .A1(n6106), .A2(n7269), .ZN(n7074) );
  NOR2_X1 U7767 ( .A1(n8759), .A2(n7074), .ZN(n6110) );
  NOR2_X1 U7768 ( .A1(n6107), .A2(n6025), .ZN(n6108) );
  OAI22_X1 U7769 ( .A1(n8894), .A2(n7258), .B1(n6116), .B2(n8954), .ZN(n6109)
         );
  OR4_X1 U7770 ( .A1(n6112), .A2(n6111), .A3(n6110), .A4(n6109), .ZN(P2_U3291)
         );
  INV_X2 U7771 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U7772 ( .A(n6900), .ZN(n6113) );
  AOI211_X1 U7773 ( .C1(n6115), .C2(n6114), .A(n8282), .B(n6113), .ZN(n6120)
         );
  NOR2_X1 U7774 ( .A1(n8254), .A2(n6116), .ZN(n6119) );
  OAI22_X1 U7775 ( .A1(n7451), .A2(n8277), .B1(n8263), .B2(n8316), .ZN(n6118)
         );
  OAI22_X1 U7776 ( .A1(n8268), .A2(n7258), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5588), .ZN(n6117) );
  OR4_X1 U7777 ( .A1(n6120), .A2(n6119), .A3(n6118), .A4(n6117), .ZN(P2_U3229)
         );
  AND2_X1 U7778 ( .A1(n4393), .A2(P2_U3152), .ZN(n9388) );
  INV_X2 U7779 ( .A(n9388), .ZN(n9120) );
  NOR2_X2 U7780 ( .A1(n5167), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9386) );
  OAI222_X1 U7781 ( .A1(P2_U3152), .A2(n6838), .B1(n9120), .B2(n6379), .C1(
        n6121), .C2(n9118), .ZN(P2_U3357) );
  OAI222_X1 U7782 ( .A1(n8559), .A2(P2_U3152), .B1(n9120), .B2(n6495), .C1(
        n5249), .C2(n9118), .ZN(P2_U3355) );
  OAI222_X1 U7783 ( .A1(P2_U3152), .A2(n8546), .B1(n9120), .B2(n6449), .C1(
        n6122), .C2(n9118), .ZN(P2_U3356) );
  OAI222_X1 U7784 ( .A1(n8568), .A2(P2_U3152), .B1(n9120), .B2(n6580), .C1(
        n6123), .C2(n9118), .ZN(P2_U3354) );
  NAND2_X1 U7785 ( .A1(n5167), .A2(P1_U3084), .ZN(n8008) );
  AND2_X1 U7786 ( .A1(n4395), .A2(P1_U3084), .ZN(n7341) );
  INV_X2 U7787 ( .A(n7341), .ZN(n8004) );
  INV_X1 U7788 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6148) );
  NAND2_X1 U7789 ( .A1(n6149), .A2(n6148), .ZN(n6147) );
  NAND2_X1 U7790 ( .A1(n6147), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6125) );
  INV_X1 U7791 ( .A(n10355), .ZN(n6126) );
  OAI222_X1 U7792 ( .A1(n8008), .A2(n6496), .B1(n8004), .B2(n6495), .C1(
        P1_U3084), .C2(n6126), .ZN(P1_U3350) );
  NAND2_X1 U7793 ( .A1(n6127), .A2(n4550), .ZN(n6150) );
  INV_X1 U7794 ( .A(n6150), .ZN(n6128) );
  NOR2_X1 U7795 ( .A1(n6129), .A2(n6128), .ZN(n6582) );
  INV_X1 U7796 ( .A(n6582), .ZN(n6560) );
  OAI222_X1 U7797 ( .A1(n8008), .A2(n6581), .B1(n8004), .B2(n6580), .C1(
        P1_U3084), .C2(n6560), .ZN(P1_U3349) );
  NAND2_X1 U7798 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6130) );
  XNOR2_X1 U7799 ( .A(n6130), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6382) );
  INV_X1 U7800 ( .A(n6382), .ZN(n6367) );
  INV_X1 U7801 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6381) );
  OAI222_X1 U7802 ( .A1(n6367), .A2(P1_U3084), .B1(n8004), .B2(n6379), .C1(
        n6381), .C2(n8008), .ZN(P1_U3352) );
  AND2_X1 U7803 ( .A1(n6519), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6131) );
  INV_X1 U7804 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6140) );
  AND3_X1 U7805 ( .A1(n7654), .A2(P1_B_REG_SCAN_IN), .A3(n7525), .ZN(n6136) );
  INV_X1 U7806 ( .A(n7525), .ZN(n6134) );
  INV_X1 U7807 ( .A(P1_B_REG_SCAN_IN), .ZN(n6133) );
  AND2_X1 U7808 ( .A1(n6134), .A2(n6133), .ZN(n6135) );
  OR2_X1 U7809 ( .A1(n10429), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6138) );
  NAND2_X1 U7810 ( .A1(n6132), .A2(n7654), .ZN(n6137) );
  NAND2_X1 U7811 ( .A1(n6138), .A2(n6137), .ZN(n6322) );
  INV_X1 U7812 ( .A(n6322), .ZN(n6400) );
  NAND2_X1 U7813 ( .A1(n6400), .A2(n10443), .ZN(n6139) );
  OAI21_X1 U7814 ( .B1(n10443), .B2(n6140), .A(n6139), .ZN(P1_U3441) );
  INV_X1 U7815 ( .A(n8587), .ZN(n6142) );
  INV_X1 U7816 ( .A(n6754), .ZN(n6145) );
  OAI222_X1 U7817 ( .A1(n6142), .A2(P2_U3152), .B1(n9120), .B2(n6145), .C1(
        n6141), .C2(n9118), .ZN(P2_U3353) );
  INV_X1 U7818 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6756) );
  NAND2_X1 U7819 ( .A1(n6150), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6143) );
  XNOR2_X1 U7820 ( .A(n6143), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6755) );
  INV_X1 U7821 ( .A(n6755), .ZN(n6144) );
  OAI222_X1 U7822 ( .A1(n8008), .A2(n6756), .B1(n8004), .B2(n6145), .C1(
        P1_U3084), .C2(n6144), .ZN(P1_U3348) );
  INV_X1 U7823 ( .A(n6773), .ZN(n6152) );
  AOI22_X1 U7824 ( .A1(n8600), .A2(P2_STATE_REG_SCAN_IN), .B1(n9386), .B2(
        P1_DATAO_REG_6__SCAN_IN), .ZN(n6146) );
  OAI21_X1 U7825 ( .B1(n6152), .B2(n9120), .A(n6146), .ZN(P2_U3352) );
  OAI222_X1 U7826 ( .A1(P1_U3084), .A2(n6546), .B1(n8004), .B2(n6449), .C1(
        n6448), .C2(n8008), .ZN(P1_U3351) );
  INV_X1 U7827 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6153) );
  NAND2_X1 U7828 ( .A1(n6155), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6151) );
  XNOR2_X1 U7829 ( .A(n6151), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6774) );
  INV_X1 U7830 ( .A(n6774), .ZN(n6230) );
  OAI222_X1 U7831 ( .A1(n8008), .A2(n6153), .B1(n8004), .B2(n6152), .C1(
        P1_U3084), .C2(n6230), .ZN(P1_U3347) );
  INV_X1 U7832 ( .A(n4780), .ZN(n6157) );
  AOI22_X1 U7833 ( .A1(n8614), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n9386), .ZN(n6154) );
  OAI21_X1 U7834 ( .B1(n6157), .B2(n9120), .A(n6154), .ZN(P2_U3351) );
  INV_X1 U7835 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6158) );
  OR2_X1 U7836 ( .A1(n6161), .A2(n10343), .ZN(n6156) );
  XNOR2_X1 U7837 ( .A(n6156), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6745) );
  INV_X1 U7838 ( .A(n6745), .ZN(n6300) );
  OAI222_X1 U7839 ( .A1(n8008), .A2(n6158), .B1(n8004), .B2(n6157), .C1(
        P1_U3084), .C2(n6300), .ZN(P1_U3346) );
  INV_X1 U7840 ( .A(n7171), .ZN(n6165) );
  AOI22_X1 U7841 ( .A1(n8627), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n9386), .ZN(n6159) );
  OAI21_X1 U7842 ( .B1(n6165), .B2(n9120), .A(n6159), .ZN(P2_U3350) );
  NAND2_X1 U7843 ( .A1(n6161), .A2(n6160), .ZN(n6163) );
  NAND2_X1 U7844 ( .A1(n6163), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6162) );
  MUX2_X1 U7845 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6162), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n6164) );
  AND2_X1 U7846 ( .A1(n6164), .A2(n6178), .ZN(n7172) );
  INV_X1 U7847 ( .A(n7172), .ZN(n6427) );
  OAI222_X1 U7848 ( .A1(n8008), .A2(n6166), .B1(n8004), .B2(n6165), .C1(
        P1_U3084), .C2(n6427), .ZN(P1_U3345) );
  INV_X1 U7849 ( .A(n7385), .ZN(n6171) );
  INV_X1 U7850 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n6167) );
  NAND2_X1 U7851 ( .A1(n6187), .A2(n6167), .ZN(n6191) );
  NAND2_X1 U7852 ( .A1(n6191), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6168) );
  INV_X1 U7853 ( .A(n8008), .ZN(n10349) );
  AOI22_X1 U7854 ( .A1(n7386), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n10349), .ZN(n6169) );
  OAI21_X1 U7855 ( .B1(n6171), .B2(n8004), .A(n6169), .ZN(P1_U3341) );
  AOI22_X1 U7856 ( .A1(n6918), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n9386), .ZN(n6170) );
  OAI21_X1 U7857 ( .B1(n6171), .B2(n9120), .A(n6170), .ZN(P2_U3346) );
  OR2_X1 U7858 ( .A1(n6172), .A2(P2_U3152), .ZN(n8506) );
  NAND2_X1 U7859 ( .A1(n10501), .A2(n8506), .ZN(n6174) );
  NAND2_X1 U7860 ( .A1(n6174), .A2(n6173), .ZN(n6177) );
  INV_X1 U7861 ( .A(n6814), .ZN(n6175) );
  OR2_X1 U7862 ( .A1(n10501), .A2(n6175), .ZN(n6176) );
  NOR2_X1 U7863 ( .A1(n8685), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U7864 ( .A(n9389), .ZN(n6181) );
  NAND2_X1 U7865 ( .A1(n6178), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6179) );
  XNOR2_X1 U7866 ( .A(n6179), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9862) );
  AOI22_X1 U7867 ( .A1(n9862), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n10349), .ZN(n6180) );
  OAI21_X1 U7868 ( .B1(n6181), .B2(n8004), .A(n6180), .ZN(P1_U3344) );
  INV_X1 U7869 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9354) );
  INV_X1 U7870 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8690) );
  NAND2_X1 U7871 ( .A1(n7743), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6184) );
  NAND2_X1 U7872 ( .A1(n6182), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6183) );
  OAI211_X1 U7873 ( .C1(n5545), .C2(n8690), .A(n6184), .B(n6183), .ZN(n8311)
         );
  NAND2_X1 U7874 ( .A1(n8311), .A2(P2_U3966), .ZN(n6185) );
  OAI21_X1 U7875 ( .B1(n9354), .B2(P2_U3966), .A(n6185), .ZN(P2_U3583) );
  INV_X1 U7876 ( .A(n7354), .ZN(n6189) );
  AOI22_X1 U7877 ( .A1(n8660), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n9386), .ZN(n6186) );
  OAI21_X1 U7878 ( .B1(n6189), .B2(n9120), .A(n6186), .ZN(P2_U3347) );
  OR2_X1 U7879 ( .A1(n6187), .A2(n10343), .ZN(n6188) );
  XNOR2_X1 U7880 ( .A(n6188), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7355) );
  INV_X1 U7881 ( .A(n7355), .ZN(n6446) );
  OAI222_X1 U7882 ( .A1(n8008), .A2(n6190), .B1(n8004), .B2(n6189), .C1(n6446), 
        .C2(P1_U3084), .ZN(P1_U3342) );
  INV_X1 U7883 ( .A(n7799), .ZN(n6267) );
  AOI22_X1 U7884 ( .A1(n7800), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n10349), .ZN(n6192) );
  OAI21_X1 U7885 ( .B1(n6267), .B2(n8004), .A(n6192), .ZN(P1_U3340) );
  INV_X1 U7886 ( .A(n7349), .ZN(n6196) );
  NAND2_X1 U7887 ( .A1(n6193), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6194) );
  XNOR2_X1 U7888 ( .A(n6194), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9873) );
  INV_X1 U7889 ( .A(n9873), .ZN(n6432) );
  OAI222_X1 U7890 ( .A1(n8008), .A2(n9207), .B1(n8004), .B2(n6196), .C1(n6432), 
        .C2(P1_U3084), .ZN(P1_U3343) );
  INV_X1 U7891 ( .A(n6858), .ZN(n6924) );
  OAI222_X1 U7892 ( .A1(P2_U3152), .A2(n6924), .B1(n9120), .B2(n6196), .C1(
        n6195), .C2(n9118), .ZN(P2_U3348) );
  NOR2_X1 U7893 ( .A1(n6533), .A2(P1_U3084), .ZN(n10348) );
  NAND2_X1 U7894 ( .A1(n6211), .A2(n10348), .ZN(n9930) );
  INV_X1 U7895 ( .A(n9930), .ZN(n6198) );
  AND2_X1 U7896 ( .A1(n6198), .A2(n6197), .ZN(n10418) );
  INV_X1 U7897 ( .A(n10418), .ZN(n9928) );
  OR2_X1 U7898 ( .A1(P1_U3083), .A2(n6199), .ZN(n10411) );
  INV_X1 U7899 ( .A(n10411), .ZN(n10426) );
  NAND2_X1 U7900 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7068) );
  INV_X1 U7901 ( .A(n7068), .ZN(n6214) );
  INV_X1 U7902 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6200) );
  MUX2_X1 U7903 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6200), .S(n10355), .Z(n10362) );
  INV_X1 U7904 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6412) );
  MUX2_X1 U7905 ( .A(n6412), .B(P1_REG1_REG_2__SCAN_IN), .S(n6546), .Z(n6202)
         );
  INV_X1 U7906 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6333) );
  MUX2_X1 U7907 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n6333), .S(n6382), .Z(n6360)
         );
  AND2_X1 U7908 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6361) );
  NAND2_X1 U7909 ( .A1(n6360), .A2(n6361), .ZN(n6538) );
  NAND2_X1 U7910 ( .A1(n6382), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6537) );
  NAND2_X1 U7911 ( .A1(n6538), .A2(n6537), .ZN(n6201) );
  NAND2_X1 U7912 ( .A1(n6202), .A2(n6201), .ZN(n6541) );
  OR2_X1 U7913 ( .A1(n6546), .A2(n6412), .ZN(n6203) );
  NAND2_X1 U7914 ( .A1(n6541), .A2(n6203), .ZN(n10363) );
  NAND2_X1 U7915 ( .A1(n10362), .A2(n10363), .ZN(n10361) );
  NAND2_X1 U7916 ( .A1(n10355), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6204) );
  INV_X1 U7917 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10491) );
  MUX2_X1 U7918 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10491), .S(n6582), .Z(n6551)
         );
  NAND2_X1 U7919 ( .A1(n6552), .A2(n6551), .ZN(n6550) );
  OR2_X1 U7920 ( .A1(n6582), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6205) );
  NAND2_X1 U7921 ( .A1(n6550), .A2(n6205), .ZN(n6256) );
  INV_X1 U7922 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7146) );
  MUX2_X1 U7923 ( .A(n7146), .B(P1_REG1_REG_5__SCAN_IN), .S(n6755), .Z(n6255)
         );
  OR2_X1 U7924 ( .A1(n6256), .A2(n6255), .ZN(n6253) );
  NAND2_X1 U7925 ( .A1(n6755), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6206) );
  INV_X1 U7926 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10493) );
  MUX2_X1 U7927 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n10493), .S(n6774), .Z(n6208)
         );
  NAND2_X1 U7928 ( .A1(n6207), .A2(n6208), .ZN(n6296) );
  INV_X1 U7929 ( .A(n6207), .ZN(n6210) );
  INV_X1 U7930 ( .A(n6208), .ZN(n6209) );
  NAND2_X1 U7931 ( .A1(n6210), .A2(n6209), .ZN(n6212) );
  NAND2_X1 U7932 ( .A1(n6211), .A2(n4506), .ZN(n10408) );
  INV_X1 U7933 ( .A(n6533), .ZN(n10403) );
  AOI21_X1 U7934 ( .B1(n6296), .B2(n6212), .A(n9923), .ZN(n6213) );
  AOI211_X1 U7935 ( .C1(n10426), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n6214), .B(
        n6213), .ZN(n6229) );
  OR2_X1 U7936 ( .A1(n9930), .A2(n6197), .ZN(n9924) );
  INV_X1 U7937 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6467) );
  MUX2_X1 U7938 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6467), .S(n10355), .Z(n10365) );
  INV_X1 U7939 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6215) );
  MUX2_X1 U7940 ( .A(n6215), .B(P1_REG2_REG_2__SCAN_IN), .S(n6546), .Z(n6544)
         );
  INV_X1 U7941 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6216) );
  XNOR2_X1 U7942 ( .A(n6382), .B(n6216), .ZN(n6365) );
  AND2_X1 U7943 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6217) );
  NAND2_X1 U7944 ( .A1(n6365), .A2(n6217), .ZN(n6363) );
  NAND2_X1 U7945 ( .A1(n6382), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6218) );
  NAND2_X1 U7946 ( .A1(n6363), .A2(n6218), .ZN(n6543) );
  NAND2_X1 U7947 ( .A1(n6544), .A2(n6543), .ZN(n6542) );
  OR2_X1 U7948 ( .A1(n6546), .A2(n6215), .ZN(n6219) );
  NAND2_X1 U7949 ( .A1(n6542), .A2(n6219), .ZN(n10366) );
  NAND2_X1 U7950 ( .A1(n10365), .A2(n10366), .ZN(n10364) );
  NAND2_X1 U7951 ( .A1(n10355), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6220) );
  AND2_X1 U7952 ( .A1(n10364), .A2(n6220), .ZN(n6553) );
  MUX2_X1 U7953 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n6512), .S(n6582), .Z(n6554)
         );
  NAND2_X1 U7954 ( .A1(n6553), .A2(n6554), .ZN(n6555) );
  OR2_X1 U7955 ( .A1(n6582), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6259) );
  NAND2_X1 U7956 ( .A1(n6555), .A2(n6259), .ZN(n6222) );
  INV_X1 U7957 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6221) );
  MUX2_X1 U7958 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n6221), .S(n6755), .Z(n6258)
         );
  OR2_X1 U7959 ( .A1(n6755), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6223) );
  INV_X1 U7960 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6224) );
  MUX2_X1 U7961 ( .A(n6224), .B(P1_REG2_REG_6__SCAN_IN), .S(n6774), .Z(n6225)
         );
  NAND2_X1 U7962 ( .A1(n6226), .A2(n6225), .ZN(n6227) );
  NAND3_X1 U7963 ( .A1(n10416), .A2(n6241), .A3(n6227), .ZN(n6228) );
  OAI211_X1 U7964 ( .C1(n9928), .C2(n6230), .A(n6229), .B(n6228), .ZN(P1_U3247) );
  INV_X1 U7965 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10497) );
  MUX2_X1 U7966 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10497), .S(n7172), .Z(n6236)
         );
  OR2_X1 U7967 ( .A1(n6745), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6235) );
  INV_X1 U7968 ( .A(n6235), .ZN(n6231) );
  NOR2_X1 U7969 ( .A1(n6236), .A2(n6231), .ZN(n6238) );
  OR2_X1 U7970 ( .A1(n6774), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6295) );
  NAND2_X1 U7971 ( .A1(n6296), .A2(n6295), .ZN(n6234) );
  NAND2_X1 U7972 ( .A1(n6745), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6232) );
  NAND2_X1 U7973 ( .A1(n6235), .A2(n6232), .ZN(n6294) );
  INV_X1 U7974 ( .A(n6294), .ZN(n6233) );
  NAND2_X1 U7975 ( .A1(n6234), .A2(n6233), .ZN(n6298) );
  NAND2_X1 U7976 ( .A1(n6298), .A2(n6235), .ZN(n6237) );
  NAND2_X1 U7977 ( .A1(n6237), .A2(n6236), .ZN(n6428) );
  INV_X1 U7978 ( .A(n6428), .ZN(n9857) );
  AOI21_X1 U7979 ( .B1(n6238), .B2(n6298), .A(n9857), .ZN(n6252) );
  AND2_X1 U7980 ( .A1(P1_U3084), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7255) );
  NOR2_X1 U7981 ( .A1(n10411), .A2(n4631), .ZN(n6239) );
  AOI211_X1 U7982 ( .C1(n10418), .C2(n7172), .A(n7255), .B(n6239), .ZN(n6251)
         );
  NAND2_X1 U7983 ( .A1(n6774), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6240) );
  INV_X1 U7984 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6993) );
  MUX2_X1 U7985 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n6993), .S(n6745), .Z(n6290)
         );
  NAND2_X1 U7986 ( .A1(n6289), .A2(n6290), .ZN(n6245) );
  INV_X1 U7987 ( .A(n6245), .ZN(n6291) );
  INV_X1 U7988 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6242) );
  MUX2_X1 U7989 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n6242), .S(n7172), .Z(n6246)
         );
  OR2_X1 U7990 ( .A1(n6745), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6244) );
  INV_X1 U7991 ( .A(n6244), .ZN(n6243) );
  NOR3_X1 U7992 ( .A1(n6291), .A2(n6246), .A3(n6243), .ZN(n6249) );
  NAND2_X1 U7993 ( .A1(n6245), .A2(n6244), .ZN(n6247) );
  INV_X1 U7994 ( .A(n6422), .ZN(n6248) );
  OAI21_X1 U7995 ( .B1(n6249), .B2(n6248), .A(n10416), .ZN(n6250) );
  OAI211_X1 U7996 ( .C1(n6252), .C2(n9923), .A(n6251), .B(n6250), .ZN(P1_U3249) );
  INV_X1 U7997 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6266) );
  INV_X1 U7998 ( .A(n6253), .ZN(n6254) );
  AOI211_X1 U7999 ( .C1(n6256), .C2(n6255), .A(n6254), .B(n9923), .ZN(n6257)
         );
  INV_X1 U8000 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9367) );
  NOR2_X1 U8001 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9367), .ZN(n6876) );
  NOR2_X1 U8002 ( .A1(n6257), .A2(n6876), .ZN(n6265) );
  INV_X1 U8003 ( .A(n6258), .ZN(n6260) );
  NAND3_X1 U8004 ( .A1(n6555), .A2(n6260), .A3(n6259), .ZN(n6261) );
  AOI21_X1 U8005 ( .B1(n6262), .B2(n6261), .A(n9924), .ZN(n6263) );
  AOI21_X1 U8006 ( .B1(n10418), .B2(n6755), .A(n6263), .ZN(n6264) );
  OAI211_X1 U8007 ( .C1(n10411), .C2(n6266), .A(n6265), .B(n6264), .ZN(
        P1_U3246) );
  INV_X1 U8008 ( .A(n6883), .ZN(n6867) );
  OAI222_X1 U8009 ( .A1(P2_U3152), .A2(n6867), .B1(n9120), .B2(n6267), .C1(
        n9294), .C2(n9118), .ZN(P2_U3345) );
  INV_X1 U8010 ( .A(n7015), .ZN(n7009) );
  INV_X1 U8011 ( .A(n7804), .ZN(n6274) );
  OAI222_X1 U8012 ( .A1(P2_U3152), .A2(n7009), .B1(n9120), .B2(n6274), .C1(
        n6268), .C2(n9118), .ZN(P2_U3344) );
  INV_X1 U8013 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n6269) );
  NAND2_X1 U8014 ( .A1(n6270), .A2(n6269), .ZN(n6271) );
  NAND2_X1 U8015 ( .A1(n6271), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6273) );
  INV_X1 U8016 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6272) );
  OAI222_X1 U8017 ( .A1(n8008), .A2(n7805), .B1(n8004), .B2(n6274), .C1(n7806), 
        .C2(P1_U3084), .ZN(P1_U3339) );
  INV_X1 U8018 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9176) );
  INV_X1 U8019 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10406) );
  NAND2_X2 U8020 ( .A1(n4749), .A2(n7720), .ZN(n6472) );
  INV_X1 U8021 ( .A(n6472), .ZN(n6341) );
  NAND2_X1 U8022 ( .A1(n6341), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6285) );
  INV_X1 U8023 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6283) );
  OR2_X1 U8024 ( .A1(n6468), .A2(n6283), .ZN(n6284) );
  NAND2_X1 U8025 ( .A1(n6654), .A2(P1_U4006), .ZN(n6288) );
  OAI21_X1 U8026 ( .B1(P1_U4006), .B2(n9176), .A(n6288), .ZN(P1_U3555) );
  INV_X1 U8027 ( .A(n6289), .ZN(n6293) );
  INV_X1 U8028 ( .A(n6290), .ZN(n6292) );
  AOI21_X1 U8029 ( .B1(n6293), .B2(n6292), .A(n6291), .ZN(n6304) );
  NAND3_X1 U8030 ( .A1(n6296), .A2(n6295), .A3(n6294), .ZN(n6297) );
  AOI21_X1 U8031 ( .B1(n6298), .B2(n6297), .A(n9923), .ZN(n6302) );
  AND2_X1 U8032 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6811) );
  INV_X1 U8033 ( .A(n6811), .ZN(n6299) );
  OAI21_X1 U8034 ( .B1(n9928), .B2(n6300), .A(n6299), .ZN(n6301) );
  AOI211_X1 U8035 ( .C1(n10426), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n6302), .B(
        n6301), .ZN(n6303) );
  OAI21_X1 U8036 ( .B1(n6304), .B2(n9924), .A(n6303), .ZN(P1_U3248) );
  INV_X1 U8037 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6306) );
  NAND2_X1 U8038 ( .A1(n6307), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6309) );
  INV_X1 U8039 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6308) );
  OR2_X1 U8040 ( .A1(n10429), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6311) );
  NAND2_X1 U8041 ( .A1(n6132), .A2(n7525), .ZN(n6310) );
  OR4_X1 U8042 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n6317) );
  NOR4_X1 U8043 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n6315) );
  NOR4_X1 U8044 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6314) );
  NOR4_X1 U8045 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_29__SCAN_IN), .ZN(n6313) );
  NOR4_X1 U8046 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_27__SCAN_IN), .ZN(n6312) );
  NAND4_X1 U8047 ( .A1(n6315), .A2(n6314), .A3(n6313), .A4(n6312), .ZN(n6316)
         );
  OR4_X1 U8048 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .A3(
        n6317), .A4(n6316), .ZN(n6320) );
  NOR4_X1 U8049 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n6319) );
  NOR4_X1 U8050 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n6318) );
  NAND2_X1 U8051 ( .A1(n6319), .A2(n6318), .ZN(n9141) );
  NOR2_X1 U8052 ( .A1(n6320), .A2(n9141), .ZN(n6321) );
  OR2_X1 U8053 ( .A1(n10429), .A2(n6321), .ZN(n6399) );
  AND2_X1 U8054 ( .A1(n6322), .A2(n6399), .ZN(n6323) );
  INV_X1 U8055 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6340) );
  INV_X1 U8056 ( .A(SI_0_), .ZN(n6326) );
  INV_X1 U8057 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6325) );
  OAI21_X1 U8058 ( .B1(n4393), .B2(n6326), .A(n6325), .ZN(n6328) );
  AND2_X1 U8059 ( .A1(n6328), .A2(n6327), .ZN(n10354) );
  MUX2_X1 U8060 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10354), .S(n6380), .Z(n7796)
         );
  INV_X1 U8061 ( .A(n6387), .ZN(n9787) );
  INV_X1 U8062 ( .A(n6329), .ZN(n6331) );
  NOR2_X1 U8063 ( .A1(n9787), .A2(n6331), .ZN(n6338) );
  NAND2_X1 U8064 ( .A1(n6654), .A2(n6705), .ZN(n9798) );
  NAND2_X1 U8065 ( .A1(n6697), .A2(n9798), .ZN(n9696) );
  NAND2_X1 U8066 ( .A1(n6788), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6337) );
  INV_X1 U8067 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6332) );
  INV_X1 U8068 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6706) );
  OR2_X1 U8069 ( .A1(n6593), .A2(n6706), .ZN(n6334) );
  INV_X1 U8070 ( .A(n6197), .ZN(n9786) );
  AOI22_X1 U8071 ( .A1(n6338), .A2(n9696), .B1(n6663), .B2(n10189), .ZN(n6635)
         );
  OAI21_X1 U8072 ( .B1(n6705), .B2(n6329), .A(n6635), .ZN(n10320) );
  NAND2_X1 U8073 ( .A1(n10320), .A2(n10488), .ZN(n6339) );
  OAI21_X1 U8074 ( .B1(n10488), .B2(n6340), .A(n6339), .ZN(P1_U3454) );
  INV_X1 U8075 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6348) );
  NAND2_X1 U8076 ( .A1(n7974), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6346) );
  INV_X1 U8077 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6342) );
  OR2_X1 U8078 ( .A1(n7944), .A2(n6342), .ZN(n6345) );
  INV_X1 U8079 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n6343) );
  OR2_X1 U8080 ( .A1(n9570), .A2(n6343), .ZN(n6344) );
  AND3_X1 U8081 ( .A1(n6346), .A2(n6345), .A3(n6344), .ZN(n9562) );
  INV_X1 U8082 ( .A(n9562), .ZN(n9936) );
  NAND2_X1 U8083 ( .A1(n9936), .A2(P1_U4006), .ZN(n6347) );
  OAI21_X1 U8084 ( .B1(P1_U4006), .B2(n6348), .A(n6347), .ZN(P1_U3586) );
  INV_X1 U8085 ( .A(n6766), .ZN(n6349) );
  INV_X1 U8086 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n7822) );
  INV_X1 U8087 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9481) );
  NAND2_X1 U8088 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n6352) );
  XNOR2_X1 U8089 ( .A(n7903), .B(P1_REG3_REG_22__SCAN_IN), .ZN(n10033) );
  NAND2_X1 U8090 ( .A1(n10033), .A2(n7955), .ZN(n6358) );
  INV_X1 U8091 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n6355) );
  NAND2_X1 U8092 ( .A1(n7974), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6354) );
  NAND2_X1 U8093 ( .A1(n6466), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6353) );
  OAI211_X1 U8094 ( .C1(n9570), .C2(n6355), .A(n6354), .B(n6353), .ZN(n6356)
         );
  INV_X1 U8095 ( .A(n6356), .ZN(n6357) );
  INV_X1 U8096 ( .A(P1_U4006), .ZN(n9843) );
  NAND2_X1 U8097 ( .A1(n9843), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6359) );
  OAI21_X1 U8098 ( .B1(n10055), .B2(n9843), .A(n6359), .ZN(P1_U3577) );
  OAI211_X1 U8099 ( .C1(n6361), .C2(n6360), .A(n10425), .B(n6538), .ZN(n6362)
         );
  OAI21_X1 U8100 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6706), .A(n6362), .ZN(n6369) );
  NAND2_X1 U8101 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n6532) );
  INV_X1 U8102 ( .A(n6532), .ZN(n6364) );
  OAI211_X1 U8103 ( .C1(n6365), .C2(n6364), .A(n10416), .B(n6363), .ZN(n6366)
         );
  OAI21_X1 U8104 ( .B1(n9928), .B2(n6367), .A(n6366), .ZN(n6368) );
  AOI211_X1 U8105 ( .C1(n10426), .C2(P1_ADDR_REG_1__SCAN_IN), .A(n6369), .B(
        n6368), .ZN(n6370) );
  INV_X1 U8106 ( .A(n6370), .ZN(P1_U3242) );
  INV_X1 U8107 ( .A(n7819), .ZN(n6418) );
  NAND2_X1 U8108 ( .A1(n6371), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6372) );
  MUX2_X1 U8109 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6372), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n6373) );
  AND2_X1 U8110 ( .A1(n6375), .A2(n6373), .ZN(n9891) );
  AOI22_X1 U8111 ( .A1(n9891), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n10349), .ZN(n6374) );
  OAI21_X1 U8112 ( .B1(n6418), .B2(n8004), .A(n6374), .ZN(P1_U3338) );
  INV_X1 U8113 ( .A(n7832), .ZN(n6420) );
  NAND2_X1 U8114 ( .A1(n6375), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6376) );
  XNOR2_X1 U8115 ( .A(n6376), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9906) );
  AOI22_X1 U8116 ( .A1(n9906), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n10349), .ZN(n6377) );
  OAI21_X1 U8117 ( .B1(n6420), .B2(n8004), .A(n6377), .ZN(P1_U3337) );
  OR2_X1 U8118 ( .A1(n6744), .A2(n6379), .ZN(n6385) );
  OR2_X1 U8119 ( .A1(n9680), .A2(n6381), .ZN(n6384) );
  NAND2_X2 U8120 ( .A1(n6696), .A2(n6520), .ZN(n8121) );
  NAND2_X2 U8121 ( .A1(n6696), .A2(n6661), .ZN(n6504) );
  XNOR2_X1 U8122 ( .A(n6388), .B(n6504), .ZN(n6459) );
  INV_X1 U8123 ( .A(n6459), .ZN(n6463) );
  OR2_X2 U8124 ( .A1(n6632), .A2(n8121), .ZN(n8123) );
  OAI21_X1 U8125 ( .B1(n6705), .B2(n8127), .A(n6389), .ZN(n6390) );
  AND2_X1 U8126 ( .A1(n6392), .A2(n6391), .ZN(n6531) );
  NAND2_X1 U8127 ( .A1(n6654), .A2(n8133), .ZN(n6395) );
  INV_X2 U8128 ( .A(n8121), .ZN(n8126) );
  AOI22_X1 U8129 ( .A1(n7796), .A2(n8126), .B1(P1_REG1_REG_0__SCAN_IN), .B2(
        n6393), .ZN(n6394) );
  NAND2_X1 U8130 ( .A1(n6395), .A2(n6394), .ZN(n6530) );
  NAND2_X1 U8131 ( .A1(n6531), .A2(n6530), .ZN(n6529) );
  INV_X1 U8132 ( .A(n10447), .ZN(n6708) );
  NAND2_X1 U8133 ( .A1(n6708), .A2(n8133), .ZN(n6396) );
  NAND2_X1 U8134 ( .A1(n6397), .A2(n6396), .ZN(n6458) );
  INV_X1 U8135 ( .A(n6458), .ZN(n6462) );
  XNOR2_X1 U8136 ( .A(n6461), .B(n6462), .ZN(n6398) );
  XNOR2_X1 U8137 ( .A(n6463), .B(n6398), .ZN(n6416) );
  INV_X1 U8138 ( .A(n6676), .ZN(n6401) );
  NAND2_X1 U8139 ( .A1(n6400), .A2(n6399), .ZN(n6628) );
  INV_X1 U8140 ( .A(n6408), .ZN(n6403) );
  INV_X1 U8141 ( .A(n6402), .ZN(n9832) );
  NOR2_X1 U8142 ( .A1(n6329), .A2(n7007), .ZN(n6631) );
  NAND2_X1 U8143 ( .A1(n6408), .A2(n6631), .ZN(n6405) );
  NAND2_X1 U8144 ( .A1(n10443), .A2(n10007), .ZN(n6404) );
  AND2_X1 U8145 ( .A1(n6631), .A2(n10443), .ZN(n6406) );
  NAND2_X1 U8146 ( .A1(n6407), .A2(n6406), .ZN(n6523) );
  NAND2_X1 U8147 ( .A1(n6407), .A2(n10480), .ZN(n6521) );
  INV_X1 U8148 ( .A(n6677), .ZN(n6518) );
  NAND4_X1 U8149 ( .A1(n6523), .A2(n6521), .A3(n10443), .A4(n6518), .ZN(n7795)
         );
  AOI22_X1 U8150 ( .A1(n9556), .A2(n6708), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n7795), .ZN(n6415) );
  AND2_X1 U8151 ( .A1(n6408), .A2(n9787), .ZN(n6413) );
  INV_X1 U8152 ( .A(n6413), .ZN(n6409) );
  INV_X1 U8153 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6410) );
  INV_X1 U8154 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6411) );
  AOI22_X1 U8155 ( .A1(n9551), .A2(n9853), .B1(n9511), .B2(n6654), .ZN(n6414)
         );
  OAI211_X1 U8156 ( .C1(n6416), .C2(n9558), .A(n6415), .B(n6414), .ZN(P1_U3220) );
  INV_X1 U8157 ( .A(n7503), .ZN(n7011) );
  OAI222_X1 U8158 ( .A1(n7011), .A2(P2_U3152), .B1(n9120), .B2(n6418), .C1(
        n6417), .C2(n9118), .ZN(P2_U3343) );
  OAI222_X1 U8159 ( .A1(P2_U3152), .A2(n7607), .B1(n9120), .B2(n6420), .C1(
        n6419), .C2(n9118), .ZN(P2_U3342) );
  INV_X1 U8160 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6440) );
  NOR2_X1 U8161 ( .A1(n9930), .A2(n6440), .ZN(n6435) );
  NAND2_X1 U8162 ( .A1(n6427), .A2(n6242), .ZN(n6421) );
  INV_X1 U8163 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9236) );
  MUX2_X1 U8164 ( .A(n9236), .B(P1_REG2_REG_9__SCAN_IN), .S(n9862), .Z(n6423)
         );
  NAND2_X1 U8165 ( .A1(n9862), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9875) );
  INV_X1 U8166 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7207) );
  MUX2_X1 U8167 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n7207), .S(n9873), .Z(n6424)
         );
  NAND2_X1 U8168 ( .A1(n9873), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6426) );
  NAND2_X1 U8169 ( .A1(n6427), .A2(n10497), .ZN(n9854) );
  NAND2_X1 U8170 ( .A1(n6428), .A2(n9854), .ZN(n6430) );
  OR2_X1 U8171 ( .A1(n9862), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6431) );
  NAND2_X1 U8172 ( .A1(n9862), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6429) );
  AND2_X1 U8173 ( .A1(n6431), .A2(n6429), .ZN(n9855) );
  NAND2_X1 U8174 ( .A1(n6430), .A2(n9855), .ZN(n9858) );
  NAND2_X1 U8175 ( .A1(n9858), .A2(n6431), .ZN(n9869) );
  INV_X1 U8176 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7208) );
  XNOR2_X1 U8177 ( .A(n9873), .B(n7208), .ZN(n9870) );
  NAND2_X1 U8178 ( .A1(n9869), .A2(n9870), .ZN(n9868) );
  NAND2_X1 U8179 ( .A1(n6432), .A2(n7208), .ZN(n6433) );
  NAND2_X1 U8180 ( .A1(n9868), .A2(n6433), .ZN(n6437) );
  INV_X1 U8181 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7358) );
  NOR3_X1 U8182 ( .A1(n6437), .A2(n7358), .A3(n9923), .ZN(n6434) );
  AOI211_X1 U8183 ( .C1(n6435), .C2(n6443), .A(n10418), .B(n6434), .ZN(n6447)
         );
  AND2_X1 U8184 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7539) );
  NOR2_X1 U8185 ( .A1(n7355), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6438) );
  NAND2_X1 U8186 ( .A1(n7355), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6436) );
  AOI21_X1 U8187 ( .B1(n6437), .B2(n6436), .A(n6438), .ZN(n6683) );
  AOI211_X1 U8188 ( .C1(n6438), .C2(n6437), .A(n9923), .B(n6683), .ZN(n6439)
         );
  AOI211_X1 U8189 ( .C1(n10426), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n7539), .B(
        n6439), .ZN(n6445) );
  NAND2_X1 U8190 ( .A1(n6446), .A2(n6440), .ZN(n6442) );
  AND2_X1 U8191 ( .A1(n7355), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6441) );
  OAI211_X1 U8192 ( .C1(n6443), .C2(n6442), .A(n6568), .B(n10416), .ZN(n6444)
         );
  OAI211_X1 U8193 ( .C1(n6447), .C2(n6446), .A(n6445), .B(n6444), .ZN(P1_U3252) );
  INV_X1 U8194 ( .A(n9853), .ZN(n6669) );
  OR2_X1 U8195 ( .A1(n8123), .A2(n6669), .ZN(n6454) );
  OR2_X1 U8196 ( .A1(n6744), .A2(n6449), .ZN(n6451) );
  NAND2_X1 U8197 ( .A1(n6945), .A2(n8133), .ZN(n6453) );
  AND2_X1 U8198 ( .A1(n6454), .A2(n6453), .ZN(n6509) );
  NAND2_X1 U8199 ( .A1(n9853), .A2(n8133), .ZN(n6456) );
  NAND2_X1 U8200 ( .A1(n6945), .A2(n8126), .ZN(n6455) );
  NAND2_X1 U8201 ( .A1(n6456), .A2(n6455), .ZN(n6457) );
  XNOR2_X1 U8202 ( .A(n6457), .B(n6504), .ZN(n6508) );
  XNOR2_X1 U8203 ( .A(n6509), .B(n6508), .ZN(n6506) );
  NAND2_X1 U8204 ( .A1(n6459), .A2(n6458), .ZN(n6460) );
  NAND2_X1 U8205 ( .A1(n6463), .A2(n6462), .ZN(n6464) );
  NAND2_X1 U8206 ( .A1(n6465), .A2(n6464), .ZN(n6507) );
  XOR2_X1 U8207 ( .A(n6506), .B(n6507), .Z(n6477) );
  AOI22_X1 U8208 ( .A1(n9556), .A2(n6945), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n7795), .ZN(n6476) );
  OR2_X1 U8209 ( .A1(n6468), .A2(n6467), .ZN(n6470) );
  INV_X1 U8210 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6473) );
  AOI22_X1 U8211 ( .A1(n9551), .A2(n6659), .B1(n9511), .B2(n6663), .ZN(n6475)
         );
  OAI211_X1 U8212 ( .C1(n6477), .C2(n9558), .A(n6476), .B(n6475), .ZN(P1_U3235) );
  INV_X1 U8213 ( .A(n7841), .ZN(n6481) );
  NAND2_X1 U8214 ( .A1(n4476), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6478) );
  XNOR2_X1 U8215 ( .A(n6478), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9920) );
  AOI22_X1 U8216 ( .A1(n9920), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n10349), .ZN(n6479) );
  OAI21_X1 U8217 ( .B1(n6481), .B2(n8004), .A(n6479), .ZN(P1_U3336) );
  INV_X1 U8218 ( .A(n7672), .ZN(n7616) );
  INV_X1 U8219 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6480) );
  OAI222_X1 U8220 ( .A1(P2_U3152), .A2(n7616), .B1(n9120), .B2(n6481), .C1(
        n6480), .C2(n9118), .ZN(P2_U3341) );
  NAND2_X1 U8221 ( .A1(n6603), .A2(n6482), .ZN(n6483) );
  INV_X1 U8222 ( .A(n6617), .ZN(n8529) );
  NAND2_X1 U8223 ( .A1(n8529), .A2(n6487), .ZN(n8351) );
  AND2_X1 U8224 ( .A1(n6605), .A2(n8351), .ZN(n8318) );
  OR2_X1 U8225 ( .A1(n8318), .A2(n7790), .ZN(n6489) );
  OR2_X1 U8226 ( .A1(n6090), .A2(n8926), .ZN(n6488) );
  AND2_X1 U8227 ( .A1(n6489), .A2(n6488), .ZN(n7046) );
  OR2_X1 U8228 ( .A1(n8318), .A2(n9079), .ZN(n6492) );
  NAND2_X1 U8229 ( .A1(n7050), .A2(n6490), .ZN(n6491) );
  AND3_X1 U8230 ( .A1(n7046), .A2(n6492), .A3(n6491), .ZN(n10516) );
  NAND2_X1 U8231 ( .A1(n10542), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6493) );
  OAI21_X1 U8232 ( .B1(n10542), .B2(n10516), .A(n6493), .ZN(P2_U3520) );
  INV_X1 U8233 ( .A(n6659), .ZN(n6494) );
  OR2_X1 U8234 ( .A1(n8123), .A2(n6494), .ZN(n6501) );
  OR2_X1 U8235 ( .A1(n6744), .A2(n6495), .ZN(n6499) );
  OR2_X1 U8236 ( .A1(n9680), .A2(n6496), .ZN(n6498) );
  NAND2_X1 U8237 ( .A1(n7858), .A2(n10355), .ZN(n6497) );
  INV_X1 U8238 ( .A(n6660), .ZN(n6961) );
  NAND2_X1 U8239 ( .A1(n6961), .A2(n8133), .ZN(n6500) );
  NAND2_X1 U8240 ( .A1(n6659), .A2(n8133), .ZN(n6503) );
  NAND2_X1 U8241 ( .A1(n6961), .A2(n8126), .ZN(n6502) );
  NAND2_X1 U8242 ( .A1(n6503), .A2(n6502), .ZN(n6505) );
  XNOR2_X1 U8243 ( .A(n6505), .B(n6504), .ZN(n6576) );
  XNOR2_X1 U8244 ( .A(n6577), .B(n6576), .ZN(n6574) );
  INV_X1 U8245 ( .A(n6508), .ZN(n6510) );
  NAND2_X1 U8246 ( .A1(n6510), .A2(n6509), .ZN(n6511) );
  XOR2_X1 U8247 ( .A(n6574), .B(n6575), .Z(n6528) );
  NAND2_X1 U8248 ( .A1(n6466), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6517) );
  INV_X1 U8249 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6512) );
  XNOR2_X1 U8250 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6719) );
  OR2_X1 U8251 ( .A1(n6593), .A2(n6719), .ZN(n6515) );
  INV_X1 U8252 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6513) );
  OR2_X1 U8253 ( .A1(n6472), .A2(n6513), .ZN(n6514) );
  AOI22_X1 U8254 ( .A1(n9551), .A2(n9852), .B1(n9511), .B2(n9853), .ZN(n6527)
         );
  INV_X1 U8255 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6960) );
  NOR2_X1 U8256 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6960), .ZN(n10356) );
  NAND4_X1 U8257 ( .A1(n6521), .A2(n6520), .A3(n6519), .A4(n6518), .ZN(n6522)
         );
  NAND2_X1 U8258 ( .A1(n6522), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6524) );
  NAND2_X1 U8259 ( .A1(n6524), .A2(n6523), .ZN(n9550) );
  NOR2_X1 U8260 ( .A1(n9531), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6525) );
  AOI211_X1 U8261 ( .C1(n6961), .C2(n9556), .A(n10356), .B(n6525), .ZN(n6526)
         );
  OAI211_X1 U8262 ( .C1(n6528), .C2(n9558), .A(n6527), .B(n6526), .ZN(P1_U3216) );
  OAI21_X1 U8263 ( .B1(n6531), .B2(n6530), .A(n6529), .ZN(n7794) );
  MUX2_X1 U8264 ( .A(n6532), .B(n7794), .S(n6533), .Z(n6536) );
  NOR2_X1 U8265 ( .A1(n6533), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6534) );
  OR2_X1 U8266 ( .A1(n6197), .A2(n6534), .ZN(n10401) );
  INV_X1 U8267 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10404) );
  NAND2_X1 U8268 ( .A1(n10401), .A2(n10404), .ZN(n6535) );
  OAI211_X1 U8269 ( .C1(n6536), .C2(n6197), .A(P1_U4006), .B(n6535), .ZN(n6564) );
  MUX2_X1 U8270 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n6412), .S(n6546), .Z(n6539)
         );
  NAND3_X1 U8271 ( .A1(n6539), .A2(n6538), .A3(n6537), .ZN(n6540) );
  AND3_X1 U8272 ( .A1(n10425), .A2(n6541), .A3(n6540), .ZN(n6548) );
  OAI211_X1 U8273 ( .C1(n6544), .C2(n6543), .A(n10416), .B(n6542), .ZN(n6545)
         );
  OAI21_X1 U8274 ( .B1(n9928), .B2(n6546), .A(n6545), .ZN(n6547) );
  AOI211_X1 U8275 ( .C1(P1_REG3_REG_2__SCAN_IN), .C2(P1_U3084), .A(n6548), .B(
        n6547), .ZN(n6549) );
  OAI211_X1 U8276 ( .C1(n10411), .C2(n10376), .A(n6564), .B(n6549), .ZN(
        P1_U3243) );
  INV_X1 U8277 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n6565) );
  OAI21_X1 U8278 ( .B1(n6552), .B2(n6551), .A(n6550), .ZN(n6562) );
  AND2_X1 U8279 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n6599) );
  INV_X1 U8280 ( .A(n6553), .ZN(n6558) );
  INV_X1 U8281 ( .A(n6554), .ZN(n6557) );
  INV_X1 U8282 ( .A(n6555), .ZN(n6556) );
  AOI21_X1 U8283 ( .B1(n6558), .B2(n6557), .A(n6556), .ZN(n6559) );
  OAI22_X1 U8284 ( .A1(n9928), .A2(n6560), .B1(n6559), .B2(n9924), .ZN(n6561)
         );
  AOI211_X1 U8285 ( .C1(n10425), .C2(n6562), .A(n6599), .B(n6561), .ZN(n6563)
         );
  OAI211_X1 U8286 ( .C1(n10411), .C2(n6565), .A(n6564), .B(n6563), .ZN(
        P1_U3245) );
  XNOR2_X1 U8287 ( .A(n7386), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n6682) );
  XOR2_X1 U8288 ( .A(n6682), .B(n6683), .Z(n6573) );
  NAND2_X1 U8289 ( .A1(n10418), .A2(n7386), .ZN(n6567) );
  AND2_X1 U8290 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9451) );
  INV_X1 U8291 ( .A(n9451), .ZN(n6566) );
  NAND2_X1 U8292 ( .A1(n6567), .A2(n6566), .ZN(n6571) );
  XNOR2_X1 U8293 ( .A(n7386), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n6569) );
  AOI211_X1 U8294 ( .C1(n6569), .C2(n6568), .A(n9924), .B(n6686), .ZN(n6570)
         );
  AOI211_X1 U8295 ( .C1(n10426), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n6571), .B(
        n6570), .ZN(n6572) );
  OAI21_X1 U8296 ( .B1(n9923), .B2(n6573), .A(n6572), .ZN(P1_U3253) );
  INV_X1 U8297 ( .A(n6576), .ZN(n6578) );
  NAND2_X1 U8298 ( .A1(n6578), .A2(n6577), .ZN(n6579) );
  NAND2_X1 U8299 ( .A1(n9852), .A2(n8133), .ZN(n6587) );
  OR2_X1 U8300 ( .A1(n6580), .A2(n6744), .ZN(n6585) );
  OR2_X1 U8301 ( .A1(n9680), .A2(n6581), .ZN(n6584) );
  NAND2_X1 U8302 ( .A1(n7858), .A2(n6582), .ZN(n6583) );
  NAND2_X1 U8303 ( .A1(n7000), .A2(n8126), .ZN(n6586) );
  NAND2_X1 U8304 ( .A1(n6587), .A2(n6586), .ZN(n6588) );
  XNOR2_X1 U8305 ( .A(n6588), .B(n8130), .ZN(n6750) );
  INV_X1 U8306 ( .A(n9852), .ZN(n6668) );
  OR2_X1 U8307 ( .A1(n8123), .A2(n6668), .ZN(n6590) );
  NAND2_X1 U8308 ( .A1(n7000), .A2(n8133), .ZN(n6589) );
  AND2_X1 U8309 ( .A1(n6590), .A2(n6589), .ZN(n6751) );
  XNOR2_X1 U8310 ( .A(n6750), .B(n6751), .ZN(n6748) );
  XOR2_X1 U8311 ( .A(n6749), .B(n6748), .Z(n6602) );
  NAND2_X1 U8312 ( .A1(n7974), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6597) );
  OR2_X1 U8313 ( .A1(n7944), .A2(n7146), .ZN(n6596) );
  OR2_X1 U8314 ( .A1(n6468), .A2(n6221), .ZN(n6595) );
  NAND2_X1 U8315 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6591) );
  NAND2_X1 U8316 ( .A1(n9367), .A2(n6591), .ZN(n6592) );
  NAND2_X1 U8317 ( .A1(n6766), .A2(n6592), .ZN(n7132) );
  OR2_X1 U8318 ( .A1(n6593), .A2(n7132), .ZN(n6594) );
  AOI22_X1 U8319 ( .A1(n9551), .A2(n9851), .B1(n9511), .B2(n6659), .ZN(n6601)
         );
  NOR2_X1 U8320 ( .A1(n9531), .A2(n6719), .ZN(n6598) );
  AOI211_X1 U8321 ( .C1(n7000), .C2(n9556), .A(n6599), .B(n6598), .ZN(n6600)
         );
  OAI211_X1 U8322 ( .C1(n6602), .C2(n9558), .A(n6601), .B(n6600), .ZN(P1_U3228) );
  NAND2_X1 U8323 ( .A1(n6604), .A2(n6603), .ZN(n6623) );
  INV_X1 U8324 ( .A(n6623), .ZN(n6610) );
  INV_X1 U8325 ( .A(n8277), .ZN(n8209) );
  AOI22_X1 U8326 ( .A1(n8209), .A2(n8528), .B1(n7050), .B2(n8280), .ZN(n6609)
         );
  INV_X1 U8327 ( .A(n6605), .ZN(n6736) );
  INV_X1 U8328 ( .A(n8351), .ZN(n6606) );
  MUX2_X1 U8329 ( .A(n6606), .B(n7050), .S(n4796), .Z(n6607) );
  OAI21_X1 U8330 ( .B1(n6736), .B2(n6607), .A(n7733), .ZN(n6608) );
  OAI211_X1 U8331 ( .C1(n6610), .C2(n7045), .A(n6609), .B(n6608), .ZN(P2_U3234) );
  AOI22_X1 U8332 ( .A1(n8209), .A2(n6611), .B1(n8280), .B2(n8950), .ZN(n6616)
         );
  AOI22_X1 U8333 ( .A1(n7733), .A2(n6614), .B1(n6623), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n6615) );
  OAI211_X1 U8334 ( .C1(n6617), .C2(n8263), .A(n6616), .B(n6615), .ZN(P2_U3224) );
  INV_X1 U8335 ( .A(n7848), .ZN(n6637) );
  XNOR2_X1 U8336 ( .A(n6618), .B(P1_IR_REG_18__SCAN_IN), .ZN(n10417) );
  AOI22_X1 U8337 ( .A1(n10417), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n10349), .ZN(n6619) );
  OAI21_X1 U8338 ( .B1(n6637), .B2(n8004), .A(n6619), .ZN(P1_U3335) );
  XNOR2_X1 U8339 ( .A(n6621), .B(n6620), .ZN(n6626) );
  INV_X1 U8340 ( .A(n8263), .ZN(n8274) );
  AOI22_X1 U8341 ( .A1(n8274), .A2(n8528), .B1(n8209), .B2(n6622), .ZN(n6625)
         );
  AOI22_X1 U8342 ( .A1(n8280), .A2(n7104), .B1(n6623), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n6624) );
  OAI211_X1 U8343 ( .C1(n6626), .C2(n8282), .A(n6625), .B(n6624), .ZN(P2_U3239) );
  NOR2_X1 U8344 ( .A1(n6628), .A2(n6627), .ZN(n6629) );
  NAND2_X1 U8345 ( .A1(n6630), .A2(n6629), .ZN(n6994) );
  INV_X2 U8346 ( .A(n10180), .ZN(n10170) );
  OAI21_X1 U8347 ( .B1(n10048), .B2(n10195), .A(n7796), .ZN(n6634) );
  INV_X1 U8348 ( .A(n10157), .ZN(n10178) );
  AOI22_X1 U8349 ( .A1(n10180), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n10178), .ZN(n6633) );
  OAI211_X1 U8350 ( .C1(n10118), .C2(n6635), .A(n6634), .B(n6633), .ZN(
        P1_U3291) );
  INV_X1 U8351 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6636) );
  OAI222_X1 U8352 ( .A1(n4764), .A2(P2_U3152), .B1(n9120), .B2(n6637), .C1(
        n6636), .C2(n9118), .ZN(P2_U3340) );
  XNOR2_X1 U8353 ( .A(n6639), .B(n6638), .ZN(n6643) );
  MUX2_X1 U8354 ( .A(n8273), .B(P2_U3152), .S(P2_REG3_REG_3__SCAN_IN), .Z(
        n6641) );
  OAI22_X1 U8355 ( .A1(n8268), .A2(n6094), .B1(n8277), .B2(n8316), .ZN(n6640)
         );
  AOI211_X1 U8356 ( .C1(n8274), .C2(n6611), .A(n6641), .B(n6640), .ZN(n6642)
         );
  OAI21_X1 U8357 ( .B1(n8282), .B2(n6643), .A(n6642), .ZN(P2_U3220) );
  NAND2_X1 U8358 ( .A1(n6646), .A2(n6645), .ZN(n6647) );
  XNOR2_X1 U8359 ( .A(n6648), .B(n6647), .ZN(n6653) );
  INV_X1 U8360 ( .A(n6649), .ZN(n7115) );
  NAND2_X1 U8361 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n8574) );
  OAI21_X1 U8362 ( .B1(n8268), .B2(n10523), .A(n8574), .ZN(n6651) );
  INV_X1 U8363 ( .A(n8526), .ZN(n7259) );
  OAI22_X1 U8364 ( .A1(n7259), .A2(n8277), .B1(n8263), .B2(n7108), .ZN(n6650)
         );
  AOI211_X1 U8365 ( .C1(n7115), .C2(n8273), .A(n6651), .B(n6650), .ZN(n6652)
         );
  OAI21_X1 U8366 ( .B1(n6653), .B2(n8282), .A(n6652), .ZN(P2_U3232) );
  NAND2_X1 U8367 ( .A1(n7721), .A2(n10007), .ZN(n9683) );
  OR2_X1 U8368 ( .A1(n9683), .A2(n9829), .ZN(n10468) );
  INV_X1 U8369 ( .A(n10468), .ZN(n10485) );
  NAND2_X1 U8370 ( .A1(n6654), .A2(n7796), .ZN(n6695) );
  NAND2_X1 U8371 ( .A1(n6695), .A2(n6655), .ZN(n6656) );
  NAND2_X1 U8372 ( .A1(n6657), .A2(n6656), .ZN(n6944) );
  NAND2_X1 U8373 ( .A1(n9853), .A2(n10452), .ZN(n9800) );
  OR2_X1 U8374 ( .A1(n9853), .A2(n6945), .ZN(n6658) );
  NAND2_X1 U8375 ( .A1(n6659), .A2(n6660), .ZN(n9741) );
  NAND2_X1 U8376 ( .A1(n9803), .A2(n9741), .ZN(n9695) );
  INV_X1 U8377 ( .A(n9695), .ZN(n6664) );
  XNOR2_X1 U8378 ( .A(n6712), .B(n6664), .ZN(n6673) );
  INV_X1 U8379 ( .A(n6673), .ZN(n6967) );
  OAI21_X1 U8380 ( .B1(n6948), .B2(n6660), .A(n6721), .ZN(n6963) );
  OAI22_X1 U8381 ( .A1(n6963), .A2(n10458), .B1(n6660), .B2(n10480), .ZN(n6674) );
  NAND2_X1 U8382 ( .A1(n9743), .A2(n6664), .ZN(n9605) );
  OAI21_X1 U8383 ( .B1(n6664), .B2(n9743), .A(n9605), .ZN(n6671) );
  NAND2_X1 U8384 ( .A1(n9789), .A2(n10007), .ZN(n6666) );
  NAND2_X1 U8385 ( .A1(n6378), .A2(n9829), .ZN(n6665) );
  OAI22_X1 U8386 ( .A1(n6669), .A2(n10167), .B1(n6668), .B2(n10169), .ZN(n6670) );
  AOI21_X1 U8387 ( .B1(n6671), .B2(n10192), .A(n6670), .ZN(n6672) );
  OAI21_X1 U8388 ( .B1(n6673), .B2(n6661), .A(n6672), .ZN(n6964) );
  AOI211_X1 U8389 ( .C1(n10485), .C2(n6967), .A(n6674), .B(n6964), .ZN(n6681)
         );
  NAND2_X1 U8390 ( .A1(n10486), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6675) );
  OAI21_X1 U8391 ( .B1(n6681), .B2(n10486), .A(n6675), .ZN(P1_U3463) );
  NAND2_X1 U8392 ( .A1(n6676), .A2(n10443), .ZN(n10441) );
  NOR2_X1 U8393 ( .A1(n6677), .A2(n10441), .ZN(n6678) );
  NAND2_X1 U8394 ( .A1(n10496), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6680) );
  OAI21_X1 U8395 ( .B1(n6681), .B2(n10496), .A(n6680), .ZN(P1_U3526) );
  OAI22_X1 U8396 ( .A1(n6683), .A2(n6682), .B1(n7386), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n7147) );
  XNOR2_X1 U8397 ( .A(n7800), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n7148) );
  XNOR2_X1 U8398 ( .A(n7147), .B(n7148), .ZN(n6693) );
  NAND2_X1 U8399 ( .A1(n10418), .A2(n7800), .ZN(n6685) );
  AND2_X1 U8400 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9510) );
  INV_X1 U8401 ( .A(n9510), .ZN(n6684) );
  NAND2_X1 U8402 ( .A1(n6685), .A2(n6684), .ZN(n6691) );
  AOI21_X1 U8403 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7386), .A(n6686), .ZN(
        n6689) );
  NAND2_X1 U8404 ( .A1(n7800), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6687) );
  OAI21_X1 U8405 ( .B1(n7800), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6687), .ZN(
        n6688) );
  NOR2_X1 U8406 ( .A1(n6689), .A2(n6688), .ZN(n7153) );
  AOI211_X1 U8407 ( .C1(n6689), .C2(n6688), .A(n9924), .B(n7153), .ZN(n6690)
         );
  AOI211_X1 U8408 ( .C1(n10426), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n6691), .B(
        n6690), .ZN(n6692) );
  OAI21_X1 U8409 ( .B1(n9923), .B2(n6693), .A(n6692), .ZN(P1_U3254) );
  NAND2_X1 U8410 ( .A1(n6694), .A2(n9799), .ZN(n9694) );
  XNOR2_X1 U8411 ( .A(n6695), .B(n9694), .ZN(n10444) );
  INV_X1 U8412 ( .A(n10444), .ZN(n6711) );
  INV_X1 U8413 ( .A(n6661), .ZN(n7431) );
  NAND2_X1 U8414 ( .A1(n10444), .A2(n7431), .ZN(n6704) );
  INV_X1 U8415 ( .A(n9799), .ZN(n6700) );
  INV_X1 U8416 ( .A(n6697), .ZN(n6698) );
  NAND2_X1 U8417 ( .A1(n9694), .A2(n6698), .ZN(n6699) );
  OAI211_X1 U8418 ( .C1(n9801), .C2(n6700), .A(n6699), .B(n10192), .ZN(n6702)
         );
  AOI22_X1 U8419 ( .A1(n10187), .A2(n6654), .B1(n9853), .B2(n10189), .ZN(n6701) );
  AND2_X1 U8420 ( .A1(n6702), .A2(n6701), .ZN(n6703) );
  NAND2_X1 U8421 ( .A1(n6704), .A2(n6703), .ZN(n10449) );
  OAI211_X1 U8422 ( .C1(n6705), .C2(n10447), .A(n10464), .B(n6946), .ZN(n10445) );
  OAI22_X1 U8423 ( .A1(n10445), .A2(n10007), .B1(n10157), .B2(n6706), .ZN(
        n6707) );
  OAI21_X1 U8424 ( .B1(n10449), .B2(n6707), .A(n10170), .ZN(n6710) );
  AOI22_X1 U8425 ( .A1(n10048), .A2(n6708), .B1(n10118), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n6709) );
  OAI211_X1 U8426 ( .C1(n6711), .C2(n10150), .A(n6710), .B(n6709), .ZN(
        P1_U3290) );
  OR2_X1 U8427 ( .A1(n6659), .A2(n6961), .ZN(n6713) );
  NAND2_X1 U8428 ( .A1(n9852), .A2(n10457), .ZN(n9742) );
  NAND2_X1 U8429 ( .A1(n9807), .A2(n9742), .ZN(n6998) );
  INV_X1 U8430 ( .A(n6998), .ZN(n9698) );
  XNOR2_X1 U8431 ( .A(n6999), .B(n9698), .ZN(n10456) );
  AOI22_X1 U8432 ( .A1(n10187), .A2(n6659), .B1(n9851), .B2(n10189), .ZN(n6717) );
  AND2_X1 U8433 ( .A1(n9803), .A2(n9605), .ZN(n6715) );
  NAND2_X1 U8434 ( .A1(n6715), .A2(n9698), .ZN(n7122) );
  OAI211_X1 U8435 ( .C1(n6715), .C2(n9698), .A(n7122), .B(n10192), .ZN(n6716)
         );
  OAI211_X1 U8436 ( .C1(n10456), .C2(n6661), .A(n6717), .B(n6716), .ZN(n10460)
         );
  NAND2_X1 U8437 ( .A1(n10460), .A2(n10170), .ZN(n6726) );
  NAND2_X1 U8438 ( .A1(n10180), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6718) );
  OAI21_X1 U8439 ( .B1(n10157), .B2(n6719), .A(n6718), .ZN(n6724) );
  INV_X1 U8440 ( .A(n10195), .ZN(n8000) );
  NAND2_X1 U8441 ( .A1(n6721), .A2(n7000), .ZN(n6722) );
  NAND2_X1 U8442 ( .A1(n7126), .A2(n6722), .ZN(n10459) );
  NOR2_X1 U8443 ( .A1(n8000), .A2(n10459), .ZN(n6723) );
  AOI211_X1 U8444 ( .C1(n10048), .C2(n7000), .A(n6724), .B(n6723), .ZN(n6725)
         );
  OAI211_X1 U8445 ( .C1(n10456), .C2(n10150), .A(n6726), .B(n6725), .ZN(
        P1_U3287) );
  INV_X1 U8446 ( .A(n6727), .ZN(n6728) );
  OR2_X1 U8447 ( .A1(n6729), .A2(n6728), .ZN(n6730) );
  INV_X1 U8448 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6742) );
  NAND2_X1 U8449 ( .A1(n4675), .A2(n6734), .ZN(n6735) );
  NAND2_X1 U8450 ( .A1(n6732), .A2(n6735), .ZN(n8952) );
  INV_X1 U8451 ( .A(n8952), .ZN(n6740) );
  XNOR2_X1 U8452 ( .A(n4675), .B(n6736), .ZN(n6737) );
  AOI222_X1 U8453 ( .A1(n8935), .A2(n6737), .B1(n6611), .B2(n8888), .C1(n8529), 
        .C2(n8886), .ZN(n8959) );
  AND2_X1 U8454 ( .A1(n8950), .A2(n7050), .ZN(n6738) );
  NOR2_X1 U8455 ( .A1(n7093), .A2(n6738), .ZN(n8956) );
  AOI22_X1 U8456 ( .A1(n8956), .A2(n9075), .B1(n9074), .B2(n8950), .ZN(n6739)
         );
  OAI211_X1 U8457 ( .C1(n9079), .C2(n6740), .A(n8959), .B(n6739), .ZN(n9081)
         );
  NAND2_X1 U8458 ( .A1(n9081), .A2(n10538), .ZN(n6741) );
  OAI21_X1 U8459 ( .B1(n10538), .B2(n6742), .A(n6741), .ZN(P2_U3454) );
  INV_X1 U8460 ( .A(n7857), .ZN(n8003) );
  OAI222_X1 U8461 ( .A1(n8915), .A2(P2_U3152), .B1(n9120), .B2(n8003), .C1(
        n6743), .C2(n9118), .ZN(P2_U3339) );
  NAND2_X1 U8462 ( .A1(n4780), .A2(n9677), .ZN(n6747) );
  AOI22_X1 U8463 ( .A1(n7859), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n7858), .B2(
        n6745), .ZN(n6746) );
  INV_X1 U8464 ( .A(n6750), .ZN(n6752) );
  NAND2_X1 U8465 ( .A1(n6752), .A2(n6751), .ZN(n6753) );
  NAND2_X1 U8466 ( .A1(n9851), .A2(n8133), .ZN(n6761) );
  NAND2_X1 U8467 ( .A1(n9677), .A2(n6754), .ZN(n6759) );
  NAND2_X1 U8468 ( .A1(n7858), .A2(n6755), .ZN(n6758) );
  OR2_X1 U8469 ( .A1(n9680), .A2(n6756), .ZN(n6757) );
  NAND2_X1 U8470 ( .A1(n7134), .A2(n8126), .ZN(n6760) );
  NAND2_X1 U8471 ( .A1(n6761), .A2(n6760), .ZN(n6762) );
  XNOR2_X1 U8472 ( .A(n6762), .B(n6504), .ZN(n6783) );
  INV_X1 U8473 ( .A(n9851), .ZN(n7221) );
  OR2_X1 U8474 ( .A1(n8123), .A2(n7221), .ZN(n6764) );
  NAND2_X1 U8475 ( .A1(n7134), .A2(n8133), .ZN(n6763) );
  NAND2_X1 U8476 ( .A1(n6764), .A2(n6763), .ZN(n6873) );
  NAND2_X1 U8477 ( .A1(n6466), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6772) );
  OR2_X1 U8478 ( .A1(n9570), .A2(n6224), .ZN(n6771) );
  INV_X1 U8479 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6765) );
  NAND2_X1 U8480 ( .A1(n6766), .A2(n6765), .ZN(n6767) );
  NAND2_X1 U8481 ( .A1(n4499), .A2(n6767), .ZN(n7227) );
  OR2_X1 U8482 ( .A1(n6593), .A2(n7227), .ZN(n6770) );
  INV_X1 U8483 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n6768) );
  OR2_X1 U8484 ( .A1(n6472), .A2(n6768), .ZN(n6769) );
  NAND2_X1 U8485 ( .A1(n9850), .A2(n8133), .ZN(n6778) );
  NAND2_X1 U8486 ( .A1(n6773), .A2(n9677), .ZN(n6776) );
  AOI22_X1 U8487 ( .A1(n7859), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n7858), .B2(
        n6774), .ZN(n6775) );
  AND2_X2 U8488 ( .A1(n6776), .A2(n6775), .ZN(n7228) );
  OR2_X1 U8489 ( .A1(n7228), .A2(n8121), .ZN(n6777) );
  NAND2_X1 U8490 ( .A1(n6778), .A2(n6777), .ZN(n6779) );
  XNOR2_X1 U8491 ( .A(n6779), .B(n6504), .ZN(n7063) );
  OR2_X1 U8492 ( .A1(n8123), .A2(n4709), .ZN(n6781) );
  OR2_X1 U8493 ( .A1(n7228), .A2(n8127), .ZN(n6780) );
  NAND2_X1 U8494 ( .A1(n6781), .A2(n6780), .ZN(n7062) );
  AOI22_X1 U8495 ( .A1(n6783), .A2(n6873), .B1(n7063), .B2(n7062), .ZN(n6782)
         );
  OAI21_X1 U8496 ( .B1(n6783), .B2(n6873), .A(n7062), .ZN(n6786) );
  INV_X1 U8497 ( .A(n7063), .ZN(n6785) );
  NOR2_X1 U8498 ( .A1(n7062), .A2(n6873), .ZN(n6784) );
  INV_X1 U8499 ( .A(n6783), .ZN(n7061) );
  AOI22_X1 U8500 ( .A1(n6786), .A2(n6785), .B1(n6784), .B2(n7061), .ZN(n6787)
         );
  NAND2_X1 U8501 ( .A1(n6788), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6796) );
  INV_X1 U8502 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6789) );
  OR2_X1 U8503 ( .A1(n7944), .A2(n6789), .ZN(n6795) );
  INV_X1 U8504 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6790) );
  NAND2_X1 U8505 ( .A1(n4499), .A2(n6790), .ZN(n6791) );
  NAND2_X1 U8506 ( .A1(n6804), .A2(n6791), .ZN(n6992) );
  OR2_X1 U8507 ( .A1(n6593), .A2(n6992), .ZN(n6794) );
  INV_X1 U8508 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n6792) );
  OR2_X1 U8509 ( .A1(n6472), .A2(n6792), .ZN(n6793) );
  NAND2_X1 U8510 ( .A1(n7232), .A2(n8126), .ZN(n6797) );
  OAI21_X1 U8511 ( .B1(n7253), .B2(n8127), .A(n6797), .ZN(n6798) );
  INV_X2 U8512 ( .A(n8096), .ZN(n8130) );
  XNOR2_X1 U8513 ( .A(n6798), .B(n8096), .ZN(n7177) );
  OR2_X1 U8514 ( .A1(n8123), .A2(n7253), .ZN(n6800) );
  NAND2_X1 U8515 ( .A1(n7232), .A2(n8133), .ZN(n6799) );
  AND2_X1 U8516 ( .A1(n6800), .A2(n6799), .ZN(n7202) );
  INV_X1 U8517 ( .A(n7202), .ZN(n7179) );
  XNOR2_X1 U8518 ( .A(n7177), .B(n7179), .ZN(n6801) );
  XNOR2_X1 U8519 ( .A(n7178), .B(n6801), .ZN(n6802) );
  NAND2_X1 U8520 ( .A1(n6802), .A2(n9507), .ZN(n6813) );
  NAND2_X1 U8521 ( .A1(n7974), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6809) );
  OR2_X1 U8522 ( .A1(n7944), .A2(n10497), .ZN(n6808) );
  OR2_X1 U8523 ( .A1(n9570), .A2(n6242), .ZN(n6807) );
  INV_X1 U8524 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6803) );
  NAND2_X1 U8525 ( .A1(n6804), .A2(n6803), .ZN(n6805) );
  NAND2_X1 U8526 ( .A1(n7186), .A2(n6805), .ZN(n7285) );
  OR2_X1 U8527 ( .A1(n6593), .A2(n7285), .ZN(n6806) );
  NAND4_X1 U8528 ( .A1(n6809), .A2(n6808), .A3(n6807), .A4(n6806), .ZN(n9848)
         );
  OAI22_X1 U8529 ( .A1(n9531), .A2(n6992), .B1(n9529), .B2(n7242), .ZN(n6810)
         );
  AOI211_X1 U8530 ( .C1(n9511), .C2(n9850), .A(n6811), .B(n6810), .ZN(n6812)
         );
  OAI211_X1 U8531 ( .C1(n10473), .C2(n9544), .A(n6813), .B(n6812), .ZN(
        P1_U3211) );
  NOR2_X1 U8532 ( .A1(n10501), .A2(n6814), .ZN(n6817) );
  OR2_X1 U8533 ( .A1(n6034), .A2(P2_U3152), .ZN(n9112) );
  OAI21_X1 U8534 ( .B1(n6815), .B2(n9112), .A(n8506), .ZN(n6816) );
  AND2_X1 U8535 ( .A1(n6861), .A2(n8687), .ZN(n6818) );
  INV_X1 U8536 ( .A(n8675), .ZN(n8679) );
  XNOR2_X1 U8537 ( .A(n6883), .B(n6819), .ZN(n6881) );
  MUX2_X1 U8538 ( .A(n5525), .B(P2_REG1_REG_2__SCAN_IN), .S(n8546), .Z(n8550)
         );
  XNOR2_X1 U8539 ( .A(n6838), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n8537) );
  AND2_X1 U8540 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n8536) );
  NAND2_X1 U8541 ( .A1(n8537), .A2(n8536), .ZN(n8535) );
  INV_X1 U8542 ( .A(n6838), .ZN(n8534) );
  NAND2_X1 U8543 ( .A1(n8534), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6820) );
  NAND2_X1 U8544 ( .A1(n8535), .A2(n6820), .ZN(n8549) );
  NAND2_X1 U8545 ( .A1(n8550), .A2(n8549), .ZN(n8548) );
  OR2_X1 U8546 ( .A1(n8546), .A2(n5525), .ZN(n6821) );
  NAND2_X1 U8547 ( .A1(n8548), .A2(n6821), .ZN(n8562) );
  XNOR2_X1 U8548 ( .A(n8559), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n8563) );
  NAND2_X1 U8549 ( .A1(n8562), .A2(n8563), .ZN(n8561) );
  OR2_X1 U8550 ( .A1(n8559), .A2(n5544), .ZN(n6822) );
  NAND2_X1 U8551 ( .A1(n8561), .A2(n6822), .ZN(n8577) );
  XNOR2_X1 U8552 ( .A(n8568), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n8578) );
  NAND2_X1 U8553 ( .A1(n8577), .A2(n8578), .ZN(n8576) );
  NAND2_X1 U8554 ( .A1(n8573), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6823) );
  NAND2_X1 U8555 ( .A1(n8576), .A2(n6823), .ZN(n8590) );
  INV_X1 U8556 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6824) );
  XNOR2_X1 U8557 ( .A(n8587), .B(n6824), .ZN(n8591) );
  NAND2_X1 U8558 ( .A1(n8590), .A2(n8591), .ZN(n8589) );
  NAND2_X1 U8559 ( .A1(n8587), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6825) );
  NAND2_X1 U8560 ( .A1(n8589), .A2(n6825), .ZN(n8604) );
  INV_X1 U8561 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6826) );
  XNOR2_X1 U8562 ( .A(n8600), .B(n6826), .ZN(n8605) );
  NAND2_X1 U8563 ( .A1(n8604), .A2(n8605), .ZN(n8603) );
  NAND2_X1 U8564 ( .A1(n8600), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6827) );
  NAND2_X1 U8565 ( .A1(n8603), .A2(n6827), .ZN(n8617) );
  INV_X1 U8566 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6828) );
  XNOR2_X1 U8567 ( .A(n8614), .B(n6828), .ZN(n8618) );
  NAND2_X1 U8568 ( .A1(n8617), .A2(n8618), .ZN(n8616) );
  NAND2_X1 U8569 ( .A1(n8614), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6829) );
  NAND2_X1 U8570 ( .A1(n8616), .A2(n6829), .ZN(n8631) );
  XNOR2_X1 U8571 ( .A(n8627), .B(n9238), .ZN(n8632) );
  NAND2_X1 U8572 ( .A1(n8631), .A2(n8632), .ZN(n8630) );
  NAND2_X1 U8573 ( .A1(n8627), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6830) );
  NAND2_X1 U8574 ( .A1(n8630), .A2(n6830), .ZN(n8646) );
  INV_X1 U8575 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6831) );
  XNOR2_X1 U8576 ( .A(n9387), .B(n6831), .ZN(n8645) );
  NAND2_X1 U8577 ( .A1(n8646), .A2(n8645), .ZN(n8644) );
  NAND2_X1 U8578 ( .A1(n9387), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6832) );
  NAND2_X1 U8579 ( .A1(n8644), .A2(n6832), .ZN(n6929) );
  XNOR2_X1 U8580 ( .A(n6858), .B(n9224), .ZN(n6928) );
  NAND2_X1 U8581 ( .A1(n6929), .A2(n6928), .ZN(n6927) );
  NAND2_X1 U8582 ( .A1(n6858), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6833) );
  NAND2_X1 U8583 ( .A1(n6927), .A2(n6833), .ZN(n8659) );
  INV_X1 U8584 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6834) );
  XNOR2_X1 U8585 ( .A(n8660), .B(n6834), .ZN(n8658) );
  NAND2_X1 U8586 ( .A1(n8659), .A2(n8658), .ZN(n8657) );
  NAND2_X1 U8587 ( .A1(n8660), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6835) );
  NAND2_X1 U8588 ( .A1(n8657), .A2(n6835), .ZN(n6910) );
  XNOR2_X1 U8589 ( .A(n6918), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n6911) );
  OR2_X1 U8590 ( .A1(n6918), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6836) );
  NAND2_X1 U8591 ( .A1(n6908), .A2(n6836), .ZN(n6882) );
  XOR2_X1 U8592 ( .A(n6881), .B(n6882), .Z(n6871) );
  NOR2_X1 U8593 ( .A1(n6883), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6886) );
  AOI21_X1 U8594 ( .B1(n6883), .B2(P2_REG2_REG_13__SCAN_IN), .A(n6886), .ZN(
        n6860) );
  MUX2_X1 U8595 ( .A(n6839), .B(P2_REG2_REG_1__SCAN_IN), .S(n6838), .Z(n8531)
         );
  AND2_X1 U8596 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n8532) );
  NAND2_X1 U8597 ( .A1(n8531), .A2(n8532), .ZN(n8530) );
  NAND2_X1 U8598 ( .A1(n8534), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6840) );
  NAND2_X1 U8599 ( .A1(n8530), .A2(n6840), .ZN(n8542) );
  NAND2_X1 U8600 ( .A1(n8543), .A2(n8542), .ZN(n8557) );
  OR2_X1 U8601 ( .A1(n8546), .A2(n6837), .ZN(n8556) );
  NAND2_X1 U8602 ( .A1(n8557), .A2(n8556), .ZN(n6841) );
  OR2_X1 U8603 ( .A1(n8559), .A2(n6842), .ZN(n8569) );
  MUX2_X1 U8604 ( .A(n6843), .B(P2_REG2_REG_4__SCAN_IN), .S(n8568), .Z(n6844)
         );
  NAND2_X1 U8605 ( .A1(n6845), .A2(n6844), .ZN(n8585) );
  NAND2_X1 U8606 ( .A1(n8573), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n8584) );
  NAND2_X1 U8607 ( .A1(n8585), .A2(n8584), .ZN(n6848) );
  MUX2_X1 U8608 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n6846), .S(n8587), .Z(n6847)
         );
  NAND2_X1 U8609 ( .A1(n8587), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8597) );
  NAND2_X1 U8610 ( .A1(n8598), .A2(n8597), .ZN(n6850) );
  MUX2_X1 U8611 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n7268), .S(n8600), .Z(n6849)
         );
  NAND2_X1 U8612 ( .A1(n6850), .A2(n6849), .ZN(n8612) );
  NAND2_X1 U8613 ( .A1(n8600), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n8611) );
  NAND2_X1 U8614 ( .A1(n8612), .A2(n8611), .ZN(n6853) );
  MUX2_X1 U8615 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n6851), .S(n8614), .Z(n6852)
         );
  NAND2_X1 U8616 ( .A1(n8614), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8624) );
  NAND2_X1 U8617 ( .A1(n8625), .A2(n8624), .ZN(n6855) );
  MUX2_X1 U8618 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n7310), .S(n8627), .Z(n6854)
         );
  NAND2_X1 U8619 ( .A1(n8627), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n8638) );
  MUX2_X1 U8620 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n6856), .S(n9387), .Z(n6857)
         );
  NAND2_X1 U8621 ( .A1(n9387), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6922) );
  MUX2_X1 U8622 ( .A(n5683), .B(P2_REG2_REG_10__SCAN_IN), .S(n6858), .Z(n6921)
         );
  MUX2_X1 U8623 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n7558), .S(n8660), .Z(n8653)
         );
  MUX2_X1 U8624 ( .A(n5727), .B(P2_REG2_REG_12__SCAN_IN), .S(n6918), .Z(n6914)
         );
  OAI21_X1 U8625 ( .B1(n6860), .B2(n6859), .A(n6890), .ZN(n6869) );
  NAND2_X1 U8626 ( .A1(n6862), .A2(n6861), .ZN(n6863) );
  NAND2_X1 U8627 ( .A1(n6863), .A2(n8514), .ZN(n6865) );
  NOR2_X1 U8628 ( .A1(n6034), .A2(n8687), .ZN(n6864) );
  NAND2_X1 U8629 ( .A1(n6865), .A2(n6864), .ZN(n8681) );
  NAND2_X1 U8630 ( .A1(n6865), .A2(n6034), .ZN(n8677) );
  NAND2_X1 U8631 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7519) );
  NAND2_X1 U8632 ( .A1(n8685), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n6866) );
  OAI211_X1 U8633 ( .C1(n8677), .C2(n6867), .A(n7519), .B(n6866), .ZN(n6868)
         );
  AOI21_X1 U8634 ( .B1(n6869), .B2(n8654), .A(n6868), .ZN(n6870) );
  OAI21_X1 U8635 ( .B1(n8679), .B2(n6871), .A(n6870), .ZN(P2_U3258) );
  XNOR2_X1 U8636 ( .A(n6872), .B(n7061), .ZN(n6874) );
  NOR2_X1 U8637 ( .A1(n6874), .A2(n6873), .ZN(n7060) );
  AOI21_X1 U8638 ( .B1(n6874), .B2(n6873), .A(n7060), .ZN(n6879) );
  AOI22_X1 U8639 ( .A1(n9551), .A2(n9850), .B1(n9511), .B2(n9852), .ZN(n6878)
         );
  NOR2_X1 U8640 ( .A1(n9531), .A2(n7132), .ZN(n6875) );
  AOI211_X1 U8641 ( .C1(n7134), .C2(n9556), .A(n6876), .B(n6875), .ZN(n6877)
         );
  OAI211_X1 U8642 ( .C1(n6879), .C2(n9558), .A(n6878), .B(n6877), .ZN(P1_U3225) );
  XNOR2_X1 U8643 ( .A(n7015), .B(n6880), .ZN(n7017) );
  NAND2_X1 U8644 ( .A1(n6882), .A2(n6881), .ZN(n6885) );
  OR2_X1 U8645 ( .A1(n6883), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6884) );
  NAND2_X1 U8646 ( .A1(n6885), .A2(n6884), .ZN(n7018) );
  XOR2_X1 U8647 ( .A(n7017), .B(n7018), .Z(n6896) );
  INV_X1 U8648 ( .A(n6886), .ZN(n6888) );
  MUX2_X1 U8649 ( .A(n6887), .B(P2_REG2_REG_14__SCAN_IN), .S(n7015), .Z(n6889)
         );
  AOI21_X1 U8650 ( .B1(n6890), .B2(n6888), .A(n6889), .ZN(n7008) );
  AND3_X1 U8651 ( .A1(n6890), .A2(n6889), .A3(n6888), .ZN(n6891) );
  OAI21_X1 U8652 ( .B1(n7008), .B2(n6891), .A(n8654), .ZN(n6895) );
  INV_X1 U8653 ( .A(n8685), .ZN(n7673) );
  INV_X1 U8654 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n6892) );
  NAND2_X1 U8655 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8155) );
  OAI21_X1 U8656 ( .B1(n7673), .B2(n6892), .A(n8155), .ZN(n6893) );
  AOI21_X1 U8657 ( .B1(n8661), .B2(n7015), .A(n6893), .ZN(n6894) );
  OAI211_X1 U8658 ( .C1(n6896), .C2(n8679), .A(n6895), .B(n6894), .ZN(P2_U3259) );
  XNOR2_X1 U8659 ( .A(n6898), .B(n6897), .ZN(n6902) );
  NAND2_X1 U8660 ( .A1(n6900), .A2(n6899), .ZN(n6901) );
  NOR2_X1 U8661 ( .A1(n6901), .A2(n6902), .ZN(n6936) );
  AOI21_X1 U8662 ( .B1(n6902), .B2(n6901), .A(n6936), .ZN(n6907) );
  INV_X1 U8663 ( .A(n7270), .ZN(n6905) );
  NAND2_X1 U8664 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n8601) );
  OAI21_X1 U8665 ( .B1(n8268), .B2(n10529), .A(n8601), .ZN(n6904) );
  OAI22_X1 U8666 ( .A1(n7259), .A2(n8263), .B1(n8277), .B2(n7305), .ZN(n6903)
         );
  AOI211_X1 U8667 ( .C1(n6905), .C2(n8273), .A(n6904), .B(n6903), .ZN(n6906)
         );
  OAI21_X1 U8668 ( .B1(n6907), .B2(n8282), .A(n6906), .ZN(P2_U3241) );
  INV_X1 U8669 ( .A(n6908), .ZN(n6909) );
  AOI21_X1 U8670 ( .B1(n6911), .B2(n6910), .A(n6909), .ZN(n6920) );
  INV_X1 U8671 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n6912) );
  NAND2_X1 U8672 ( .A1(P2_U3152), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7335) );
  OAI21_X1 U8673 ( .B1(n7673), .B2(n6912), .A(n7335), .ZN(n6917) );
  AOI211_X1 U8674 ( .C1(n6915), .C2(n6914), .A(n8681), .B(n6913), .ZN(n6916)
         );
  AOI211_X1 U8675 ( .C1(n8661), .C2(n6918), .A(n6917), .B(n6916), .ZN(n6919)
         );
  OAI21_X1 U8676 ( .B1(n6920), .B2(n8679), .A(n6919), .ZN(P2_U3257) );
  NAND3_X1 U8677 ( .A1(n8641), .A2(n6922), .A3(n6921), .ZN(n6923) );
  NAND2_X1 U8678 ( .A1(n8654), .A2(n6923), .ZN(n6932) );
  NOR2_X1 U8679 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9163), .ZN(n6926) );
  NOR2_X1 U8680 ( .A1(n8677), .A2(n6924), .ZN(n6925) );
  AOI211_X1 U8681 ( .C1(P2_ADDR_REG_10__SCAN_IN), .C2(n8685), .A(n6926), .B(
        n6925), .ZN(n6931) );
  OAI211_X1 U8682 ( .C1(n6929), .C2(n6928), .A(n6927), .B(n8675), .ZN(n6930)
         );
  OAI211_X1 U8683 ( .C1(n6933), .C2(n6932), .A(n6931), .B(n6930), .ZN(P2_U3255) );
  OAI21_X1 U8684 ( .B1(n6936), .B2(n6935), .A(n6934), .ZN(n6938) );
  NAND3_X1 U8685 ( .A1(n6938), .A2(n7733), .A3(n6937), .ZN(n6943) );
  INV_X1 U8686 ( .A(n6939), .ZN(n7542) );
  OAI22_X1 U8687 ( .A1(n8268), .A2(n7291), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5620), .ZN(n6941) );
  OAI22_X1 U8688 ( .A1(n7451), .A2(n8263), .B1(n8277), .B2(n7493), .ZN(n6940)
         );
  AOI211_X1 U8689 ( .C1(n7542), .C2(n8273), .A(n6941), .B(n6940), .ZN(n6942)
         );
  NAND2_X1 U8690 ( .A1(n6943), .A2(n6942), .ZN(P2_U3215) );
  INV_X1 U8691 ( .A(n10150), .ZN(n6968) );
  XNOR2_X1 U8692 ( .A(n9697), .B(n6944), .ZN(n10455) );
  AND2_X1 U8693 ( .A1(n6946), .A2(n6945), .ZN(n6947) );
  NOR2_X1 U8694 ( .A1(n6948), .A2(n6947), .ZN(n10450) );
  AOI22_X1 U8695 ( .A1(n10195), .A2(n10450), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n10178), .ZN(n6949) );
  OAI21_X1 U8696 ( .B1(n10452), .B2(n10182), .A(n6949), .ZN(n6958) );
  NAND2_X1 U8697 ( .A1(n10455), .A2(n7431), .ZN(n6956) );
  AOI22_X1 U8698 ( .A1(n6663), .A2(n10187), .B1(n10189), .B2(n6659), .ZN(n6955) );
  OAI21_X1 U8699 ( .B1(n6952), .B2(n6951), .A(n6950), .ZN(n6953) );
  NAND2_X1 U8700 ( .A1(n6953), .A2(n10192), .ZN(n6954) );
  NAND3_X1 U8701 ( .A1(n6956), .A2(n6955), .A3(n6954), .ZN(n10453) );
  MUX2_X1 U8702 ( .A(n10453), .B(P1_REG2_REG_2__SCAN_IN), .S(n10180), .Z(n6957) );
  AOI211_X1 U8703 ( .C1(n6968), .C2(n10455), .A(n6958), .B(n6957), .ZN(n6959)
         );
  INV_X1 U8704 ( .A(n6959), .ZN(P1_U3289) );
  AOI22_X1 U8705 ( .A1(n10048), .A2(n6961), .B1(n6960), .B2(n10178), .ZN(n6962) );
  OAI21_X1 U8706 ( .B1(n8000), .B2(n6963), .A(n6962), .ZN(n6966) );
  MUX2_X1 U8707 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6964), .S(n10170), .Z(n6965)
         );
  AOI211_X1 U8708 ( .C1(n6968), .C2(n6967), .A(n6966), .B(n6965), .ZN(n6969)
         );
  INV_X1 U8709 ( .A(n6969), .ZN(P1_U3288) );
  NAND2_X1 U8710 ( .A1(n8675), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6970) );
  OAI21_X1 U8711 ( .B1(n8681), .B2(n6971), .A(n6970), .ZN(n6975) );
  NAND2_X1 U8712 ( .A1(n8675), .A2(n6972), .ZN(n6973) );
  OAI211_X1 U8713 ( .C1(n8681), .C2(P2_REG2_REG_0__SCAN_IN), .A(n6973), .B(
        n8677), .ZN(n6974) );
  MUX2_X1 U8714 ( .A(n6975), .B(n6974), .S(P2_IR_REG_0__SCAN_IN), .Z(n6978) );
  INV_X1 U8715 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6976) );
  OAI22_X1 U8716 ( .A1(n7673), .A2(n6976), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7045), .ZN(n6977) );
  OR2_X1 U8717 ( .A1(n6978), .A2(n6977), .ZN(P2_U3245) );
  NAND2_X1 U8718 ( .A1(n6937), .A2(n6979), .ZN(n6983) );
  XNOR2_X1 U8719 ( .A(n6981), .B(n6980), .ZN(n6982) );
  NAND2_X1 U8720 ( .A1(n6983), .A2(n6982), .ZN(n7085) );
  OAI211_X1 U8721 ( .C1(n6983), .C2(n6982), .A(n7085), .B(n7733), .ZN(n6987)
         );
  NAND2_X1 U8722 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n8628) );
  OAI21_X1 U8723 ( .B1(n8277), .B2(n7582), .A(n8628), .ZN(n6985) );
  OAI22_X1 U8724 ( .A1(n8254), .A2(n7314), .B1(n7305), .B2(n8263), .ZN(n6984)
         );
  AOI211_X1 U8725 ( .C1(n8280), .C2(n7483), .A(n6985), .B(n6984), .ZN(n6986)
         );
  NAND2_X1 U8726 ( .A1(n6987), .A2(n6986), .ZN(P2_U3223) );
  OR2_X1 U8727 ( .A1(n7253), .A2(n7232), .ZN(n9607) );
  NAND2_X1 U8728 ( .A1(n7253), .A2(n7232), .ZN(n7279) );
  NAND2_X1 U8729 ( .A1(n9607), .A2(n7279), .ZN(n9703) );
  NAND2_X1 U8730 ( .A1(n9807), .A2(n9803), .ZN(n9601) );
  NAND2_X1 U8731 ( .A1(n9851), .A2(n6990), .ZN(n9810) );
  INV_X1 U8732 ( .A(n9741), .ZN(n6988) );
  NAND2_X1 U8733 ( .A1(n6988), .A2(n9807), .ZN(n6989) );
  NAND2_X1 U8734 ( .A1(n9850), .A2(n7228), .ZN(n9606) );
  XOR2_X1 U8735 ( .A(n7239), .B(n9703), .Z(n6991) );
  AOI222_X1 U8736 ( .A1(n10192), .A2(n6991), .B1(n9848), .B2(n10189), .C1(
        n9850), .C2(n10187), .ZN(n10472) );
  OAI22_X1 U8737 ( .A1(n10170), .A2(n6993), .B1(n6992), .B2(n10157), .ZN(n6997) );
  OAI211_X1 U8738 ( .C1(n7225), .C2(n10473), .A(n7278), .B(n10464), .ZN(n10471) );
  NOR2_X1 U8739 ( .A1(n6994), .A2(n10007), .ZN(n10161) );
  INV_X1 U8740 ( .A(n10161), .ZN(n6995) );
  NOR2_X1 U8741 ( .A1(n10471), .A2(n6995), .ZN(n6996) );
  AOI211_X1 U8742 ( .C1(n10048), .C2(n7232), .A(n6997), .B(n6996), .ZN(n7006)
         );
  NAND2_X1 U8743 ( .A1(n9851), .A2(n7134), .ZN(n7001) );
  NOR2_X1 U8744 ( .A1(n7236), .A2(n9603), .ZN(n7219) );
  NOR2_X1 U8745 ( .A1(n9850), .A2(n4710), .ZN(n7234) );
  NOR2_X1 U8746 ( .A1(n7219), .A2(n7234), .ZN(n7002) );
  XOR2_X1 U8747 ( .A(n9703), .B(n7002), .Z(n10475) );
  NAND2_X1 U8748 ( .A1(n6661), .A2(n10059), .ZN(n7003) );
  AND2_X1 U8749 ( .A1(n6504), .A2(n7003), .ZN(n7004) );
  INV_X1 U8750 ( .A(n10197), .ZN(n7411) );
  NAND2_X1 U8751 ( .A1(n10475), .A2(n7411), .ZN(n7005) );
  OAI211_X1 U8752 ( .C1(n10472), .C2(n10118), .A(n7006), .B(n7005), .ZN(
        P1_U3284) );
  INV_X1 U8753 ( .A(n7867), .ZN(n7081) );
  OAI222_X1 U8754 ( .A1(P1_U3084), .A2(n7007), .B1(n8004), .B2(n7081), .C1(
        n7868), .C2(n8008), .ZN(P1_U3333) );
  AOI21_X1 U8755 ( .B1(n6887), .B2(n7009), .A(n7008), .ZN(n7010) );
  AOI21_X1 U8756 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(n7012), .A(n7507), .ZN(
        n7025) );
  INV_X1 U8757 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7013) );
  NAND2_X1 U8758 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8275) );
  OAI21_X1 U8759 ( .B1(n7673), .B2(n7013), .A(n8275), .ZN(n7014) );
  AOI21_X1 U8760 ( .B1(n8661), .B2(n7503), .A(n7014), .ZN(n7024) );
  NOR2_X1 U8761 ( .A1(n7015), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7016) );
  AOI21_X1 U8762 ( .B1(n7018), .B2(n7017), .A(n7016), .ZN(n7504) );
  XNOR2_X1 U8763 ( .A(n7504), .B(n7503), .ZN(n7020) );
  INV_X1 U8764 ( .A(n7020), .ZN(n7022) );
  NOR2_X1 U8765 ( .A1(n7020), .A2(n7019), .ZN(n7502) );
  INV_X1 U8766 ( .A(n7502), .ZN(n7021) );
  OAI211_X1 U8767 ( .C1(P2_REG1_REG_15__SCAN_IN), .C2(n7022), .A(n7021), .B(
        n8675), .ZN(n7023) );
  OAI211_X1 U8768 ( .C1(n7025), .C2(n8681), .A(n7024), .B(n7023), .ZN(P2_U3260) );
  INV_X1 U8769 ( .A(n7027), .ZN(n7028) );
  NOR2_X1 U8770 ( .A1(n7026), .A2(n7028), .ZN(n7032) );
  NAND2_X1 U8771 ( .A1(n6732), .A2(n7029), .ZN(n7095) );
  NAND2_X1 U8772 ( .A1(n7095), .A2(n7030), .ZN(n7094) );
  INV_X1 U8773 ( .A(n6098), .ZN(n7031) );
  AOI21_X1 U8774 ( .B1(n7032), .B2(n7094), .A(n7031), .ZN(n7162) );
  OAI22_X1 U8775 ( .A1(n8316), .A2(n8926), .B1(n6081), .B2(n8924), .ZN(n7035)
         );
  NOR2_X1 U8776 ( .A1(n7162), .A2(n8931), .ZN(n7034) );
  AOI211_X1 U8777 ( .C1(n8935), .C2(n7036), .A(n7035), .B(n7034), .ZN(n7167)
         );
  INV_X1 U8778 ( .A(n7112), .ZN(n7037) );
  AOI21_X1 U8779 ( .B1(n7038), .B2(n7092), .A(n7037), .ZN(n7165) );
  AOI22_X1 U8780 ( .A1(n7165), .A2(n9075), .B1(n9074), .B2(n7038), .ZN(n7039)
         );
  OAI211_X1 U8781 ( .C1(n7162), .C2(n9047), .A(n7167), .B(n7039), .ZN(n7041)
         );
  NAND2_X1 U8782 ( .A1(n7041), .A2(n10544), .ZN(n7040) );
  OAI21_X1 U8783 ( .B1(n10544), .B2(n5544), .A(n7040), .ZN(P2_U3523) );
  INV_X1 U8784 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7043) );
  NAND2_X1 U8785 ( .A1(n7041), .A2(n10538), .ZN(n7042) );
  OAI21_X1 U8786 ( .B1(n10538), .B2(n7043), .A(n7042), .ZN(P2_U3460) );
  INV_X1 U8787 ( .A(n7880), .ZN(n7059) );
  INV_X1 U8788 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7044) );
  OAI222_X1 U8789 ( .A1(P2_U3152), .A2(n8337), .B1(n9120), .B2(n7059), .C1(
        n7044), .C2(n9118), .ZN(P2_U3337) );
  OAI22_X1 U8790 ( .A1(n8958), .A2(n7046), .B1(n7045), .B2(n8954), .ZN(n7047)
         );
  AOI21_X1 U8791 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n8958), .A(n7047), .ZN(
        n7052) );
  INV_X1 U8792 ( .A(n7048), .ZN(n7049) );
  OAI21_X1 U8793 ( .B1(n8951), .B2(n8957), .A(n7050), .ZN(n7051) );
  OAI211_X1 U8794 ( .C1(n8318), .C2(n8899), .A(n7052), .B(n7051), .ZN(P2_U3296) );
  XNOR2_X1 U8795 ( .A(n7054), .B(n7053), .ZN(n7058) );
  INV_X1 U8796 ( .A(n8520), .ZN(n7551) );
  OAI22_X1 U8797 ( .A1(n8277), .A2(n7551), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9163), .ZN(n7056) );
  OAI22_X1 U8798 ( .A1(n8254), .A2(n7643), .B1(n7582), .B2(n8263), .ZN(n7055)
         );
  AOI211_X1 U8799 ( .C1(n8280), .C2(n7645), .A(n7056), .B(n7055), .ZN(n7057)
         );
  OAI21_X1 U8800 ( .B1(n7058), .B2(n8282), .A(n7057), .ZN(P2_U3219) );
  INV_X1 U8801 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7881) );
  OAI222_X1 U8802 ( .A1(n8008), .A2(n7881), .B1(P1_U3084), .B2(n9690), .C1(
        n8004), .C2(n7059), .ZN(P1_U3332) );
  AOI21_X1 U8803 ( .B1(n7061), .B2(n6872), .A(n7060), .ZN(n7065) );
  XNOR2_X1 U8804 ( .A(n7063), .B(n7062), .ZN(n7064) );
  XNOR2_X1 U8805 ( .A(n7065), .B(n7064), .ZN(n7072) );
  INV_X1 U8806 ( .A(n7227), .ZN(n7066) );
  AOI22_X1 U8807 ( .A1(n9511), .A2(n9851), .B1(n7066), .B2(n9550), .ZN(n7070)
         );
  NAND2_X1 U8808 ( .A1(n9556), .A2(n4710), .ZN(n7069) );
  INV_X1 U8809 ( .A(n7253), .ZN(n9849) );
  NAND2_X1 U8810 ( .A1(n9551), .A2(n9849), .ZN(n7067) );
  NAND4_X1 U8811 ( .A1(n7070), .A2(n7069), .A3(n7068), .A4(n7067), .ZN(n7071)
         );
  AOI21_X1 U8812 ( .B1(n7072), .B2(n9507), .A(n7071), .ZN(n7073) );
  INV_X1 U8813 ( .A(n7073), .ZN(P1_U3237) );
  OAI21_X1 U8814 ( .B1(n7258), .B2(n10528), .A(n7074), .ZN(n7076) );
  AOI211_X1 U8815 ( .C1(n10536), .C2(n7077), .A(n7076), .B(n7075), .ZN(n7079)
         );
  OR2_X1 U8816 ( .A1(n7079), .A2(n10537), .ZN(n7078) );
  OAI21_X1 U8817 ( .B1(n10538), .B2(n5591), .A(n7078), .ZN(P2_U3466) );
  OR2_X1 U8818 ( .A1(n7079), .A2(n10542), .ZN(n7080) );
  OAI21_X1 U8819 ( .B1(n10544), .B2(n6824), .A(n7080), .ZN(P2_U3525) );
  OAI222_X1 U8820 ( .A1(P2_U3152), .A2(n6025), .B1(n9120), .B2(n7081), .C1(
        n9374), .C2(n9118), .ZN(P2_U3338) );
  NAND2_X1 U8821 ( .A1(n7083), .A2(n7082), .ZN(n7087) );
  NAND2_X1 U8822 ( .A1(n7085), .A2(n7084), .ZN(n7086) );
  XOR2_X1 U8823 ( .A(n7087), .B(n7086), .Z(n7091) );
  NAND2_X1 U8824 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n8642) );
  OAI21_X1 U8825 ( .B1(n8277), .B2(n7554), .A(n8642), .ZN(n7089) );
  OAI22_X1 U8826 ( .A1(n8254), .A2(n7565), .B1(n7493), .B2(n8263), .ZN(n7088)
         );
  AOI211_X1 U8827 ( .C1(n8280), .C2(n7567), .A(n7089), .B(n7088), .ZN(n7090)
         );
  OAI21_X1 U8828 ( .B1(n7091), .B2(n8282), .A(n7090), .ZN(P2_U3233) );
  OAI211_X1 U8829 ( .C1(n7093), .C2(n10518), .A(n9075), .B(n7092), .ZN(n10517)
         );
  OAI21_X1 U8830 ( .B1(n7095), .B2(n7030), .A(n7094), .ZN(n10521) );
  NAND2_X1 U8831 ( .A1(n8953), .A2(n10521), .ZN(n7097) );
  NAND2_X1 U8832 ( .A1(n8871), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n7096) );
  OAI211_X1 U8833 ( .C1(n8944), .C2(n10517), .A(n7097), .B(n7096), .ZN(n7103)
         );
  INV_X1 U8834 ( .A(n7098), .ZN(n7099) );
  AOI21_X1 U8835 ( .B1(n7030), .B2(n7100), .A(n7099), .ZN(n7101) );
  OAI222_X1 U8836 ( .A1(n8926), .A2(n7108), .B1(n8924), .B2(n6090), .C1(n7790), 
        .C2(n7101), .ZN(n10519) );
  MUX2_X1 U8837 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n10519), .S(n8940), .Z(n7102)
         );
  AOI211_X1 U8838 ( .C1(n8951), .C2(n7104), .A(n7103), .B(n7102), .ZN(n7105)
         );
  INV_X1 U8839 ( .A(n7105), .ZN(P2_U3294) );
  XNOR2_X1 U8840 ( .A(n7106), .B(n7110), .ZN(n7107) );
  OAI222_X1 U8841 ( .A1(n8926), .A2(n7259), .B1(n8924), .B2(n7108), .C1(n7790), 
        .C2(n7107), .ZN(n10525) );
  OAI21_X1 U8842 ( .B1(n7111), .B2(n7110), .A(n7109), .ZN(n10527) );
  AOI22_X1 U8843 ( .A1(n8953), .A2(n10527), .B1(n8951), .B2(n6099), .ZN(n7118)
         );
  AND2_X1 U8844 ( .A1(n7112), .A2(n6099), .ZN(n7114) );
  OR2_X1 U8845 ( .A1(n7114), .A2(n7113), .ZN(n10524) );
  INV_X1 U8846 ( .A(n10524), .ZN(n7116) );
  AOI22_X1 U8847 ( .A1(n8957), .A2(n7116), .B1(n7115), .B2(n8871), .ZN(n7117)
         );
  OAI211_X1 U8848 ( .C1(n6843), .C2(n8940), .A(n7118), .B(n7117), .ZN(n7119)
         );
  AOI21_X1 U8849 ( .B1(n10525), .B2(n8940), .A(n7119), .ZN(n7120) );
  INV_X1 U8850 ( .A(n7120), .ZN(P2_U3292) );
  INV_X1 U8851 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9296) );
  NAND2_X1 U8852 ( .A1(n6661), .A2(n10468), .ZN(n10476) );
  XNOR2_X1 U8853 ( .A(n9699), .B(n7121), .ZN(n7137) );
  NAND2_X1 U8854 ( .A1(n7122), .A2(n9742), .ZN(n7123) );
  XOR2_X1 U8855 ( .A(n9699), .B(n7123), .Z(n7124) );
  AOI222_X1 U8856 ( .A1(n10192), .A2(n7124), .B1(n9850), .B2(n10189), .C1(
        n9852), .C2(n10187), .ZN(n7131) );
  INV_X1 U8857 ( .A(n7226), .ZN(n7125) );
  AOI211_X1 U8858 ( .C1(n7134), .C2(n7126), .A(n10458), .B(n7125), .ZN(n7129)
         );
  AOI21_X1 U8859 ( .B1(n10463), .B2(n7134), .A(n7129), .ZN(n7127) );
  OAI211_X1 U8860 ( .C1(n10299), .C2(n7137), .A(n7131), .B(n7127), .ZN(n7144)
         );
  NAND2_X1 U8861 ( .A1(n7144), .A2(n10488), .ZN(n7128) );
  OAI21_X1 U8862 ( .B1(n10488), .B2(n9296), .A(n7128), .ZN(P1_U3469) );
  NAND2_X1 U8863 ( .A1(n7129), .A2(n10059), .ZN(n7130) );
  OAI211_X1 U8864 ( .C1(n10157), .C2(n7132), .A(n7131), .B(n7130), .ZN(n7133)
         );
  NAND2_X1 U8865 ( .A1(n7133), .A2(n10170), .ZN(n7136) );
  AOI22_X1 U8866 ( .A1(n10048), .A2(n7134), .B1(n10180), .B2(
        P1_REG2_REG_5__SCAN_IN), .ZN(n7135) );
  OAI211_X1 U8867 ( .C1(n7137), .C2(n10197), .A(n7136), .B(n7135), .ZN(
        P1_U3286) );
  XNOR2_X1 U8868 ( .A(n7138), .B(n7139), .ZN(n7143) );
  OAI22_X1 U8869 ( .A1(n8277), .A2(n7626), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5724), .ZN(n7141) );
  OAI22_X1 U8870 ( .A1(n8254), .A2(n7560), .B1(n7554), .B2(n8263), .ZN(n7140)
         );
  AOI211_X1 U8871 ( .C1(n8280), .C2(n9073), .A(n7141), .B(n7140), .ZN(n7142)
         );
  OAI21_X1 U8872 ( .B1(n7143), .B2(n8282), .A(n7142), .ZN(P2_U3238) );
  NAND2_X1 U8873 ( .A1(n7144), .A2(n10499), .ZN(n7145) );
  OAI21_X1 U8874 ( .B1(n10499), .B2(n7146), .A(n7145), .ZN(P1_U3528) );
  INV_X1 U8875 ( .A(n7147), .ZN(n7149) );
  OAI22_X1 U8876 ( .A1(n7149), .A2(n7148), .B1(n7800), .B2(
        P1_REG1_REG_13__SCAN_IN), .ZN(n7151) );
  XNOR2_X1 U8877 ( .A(n7806), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n7150) );
  NAND2_X1 U8878 ( .A1(n7150), .A2(n7151), .ZN(n7595) );
  OAI21_X1 U8879 ( .B1(n7151), .B2(n7150), .A(n7595), .ZN(n7152) );
  INV_X1 U8880 ( .A(n7152), .ZN(n7159) );
  NAND2_X1 U8881 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9408) );
  OAI21_X1 U8882 ( .B1(n9928), .B2(n7806), .A(n9408), .ZN(n7157) );
  INV_X1 U8883 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7154) );
  AOI211_X1 U8884 ( .C1(n7155), .C2(n7154), .A(n4552), .B(n9924), .ZN(n7156)
         );
  AOI211_X1 U8885 ( .C1(n10426), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n7157), .B(
        n7156), .ZN(n7158) );
  OAI21_X1 U8886 ( .B1(n7159), .B2(n9923), .A(n7158), .ZN(P1_U3255) );
  NAND2_X1 U8887 ( .A1(n8958), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7160) );
  OAI21_X1 U8888 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(n8954), .A(n7160), .ZN(
        n7164) );
  OR2_X1 U8889 ( .A1(n8949), .A2(n7161), .ZN(n8920) );
  OAI22_X1 U8890 ( .A1(n7162), .A2(n8920), .B1(n6094), .B2(n8894), .ZN(n7163)
         );
  AOI211_X1 U8891 ( .C1(n8957), .C2(n7165), .A(n7164), .B(n7163), .ZN(n7166)
         );
  OAI21_X1 U8892 ( .B1(n7167), .B2(n8949), .A(n7166), .ZN(P2_U3293) );
  NAND2_X1 U8893 ( .A1(n9389), .A2(n9677), .ZN(n7169) );
  AOI22_X1 U8894 ( .A1(n7859), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n7858), .B2(
        n9862), .ZN(n7168) );
  INV_X1 U8895 ( .A(n7184), .ZN(n9595) );
  NAND2_X1 U8896 ( .A1(n7171), .A2(n9677), .ZN(n7174) );
  AOI22_X1 U8897 ( .A1(n7859), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7858), .B2(
        n7172), .ZN(n7173) );
  NAND2_X1 U8898 ( .A1(n9590), .A2(n8133), .ZN(n7176) );
  OR2_X1 U8899 ( .A1(n8123), .A2(n7242), .ZN(n7175) );
  NAND2_X1 U8900 ( .A1(n7176), .A2(n7175), .ZN(n7463) );
  INV_X1 U8901 ( .A(n7463), .ZN(n7180) );
  NAND3_X1 U8902 ( .A1(n7465), .A2(n7180), .A3(n7475), .ZN(n7248) );
  NAND2_X1 U8903 ( .A1(n9590), .A2(n8126), .ZN(n7182) );
  NAND2_X1 U8904 ( .A1(n9848), .A2(n8133), .ZN(n7181) );
  NAND2_X1 U8905 ( .A1(n7182), .A2(n7181), .ZN(n7183) );
  XNOR2_X1 U8906 ( .A(n7183), .B(n8096), .ZN(n7473) );
  NAND2_X1 U8907 ( .A1(n7248), .A2(n4906), .ZN(n7251) );
  NAND2_X1 U8908 ( .A1(n7184), .A2(n8126), .ZN(n7194) );
  NAND2_X1 U8909 ( .A1(n6466), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7192) );
  OR2_X1 U8910 ( .A1(n9570), .A2(n9236), .ZN(n7191) );
  NAND2_X1 U8911 ( .A1(n7186), .A2(n7185), .ZN(n7187) );
  NAND2_X1 U8912 ( .A1(n7210), .A2(n7187), .ZN(n7323) );
  OR2_X1 U8913 ( .A1(n6593), .A2(n7323), .ZN(n7190) );
  INV_X1 U8914 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n7188) );
  OR2_X1 U8915 ( .A1(n6472), .A2(n7188), .ZN(n7189) );
  OR2_X1 U8916 ( .A1(n9591), .A2(n8127), .ZN(n7193) );
  NAND2_X1 U8917 ( .A1(n7194), .A2(n7193), .ZN(n7195) );
  XNOR2_X1 U8918 ( .A(n7195), .B(n8130), .ZN(n7201) );
  INV_X1 U8919 ( .A(n7201), .ZN(n7199) );
  NAND2_X1 U8920 ( .A1(n7184), .A2(n8133), .ZN(n7197) );
  OR2_X1 U8921 ( .A1(n8123), .A2(n9591), .ZN(n7196) );
  NAND2_X1 U8922 ( .A1(n7197), .A2(n7196), .ZN(n7200) );
  INV_X1 U8923 ( .A(n7200), .ZN(n7198) );
  AND2_X1 U8924 ( .A1(n7201), .A2(n7200), .ZN(n7466) );
  NOR2_X1 U8925 ( .A1(n7474), .A2(n7466), .ZN(n7204) );
  AND2_X1 U8926 ( .A1(n7457), .A2(n7463), .ZN(n7203) );
  NAND2_X1 U8927 ( .A1(n7203), .A2(n7458), .ZN(n7247) );
  NAND3_X1 U8928 ( .A1(n7251), .A2(n7204), .A3(n7247), .ZN(n7477) );
  INV_X1 U8929 ( .A(n7477), .ZN(n7206) );
  AOI21_X1 U8930 ( .B1(n7251), .B2(n7247), .A(n7204), .ZN(n7205) );
  OAI21_X1 U8931 ( .B1(n7206), .B2(n7205), .A(n9507), .ZN(n7218) );
  AND2_X1 U8932 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9861) );
  NAND2_X1 U8933 ( .A1(n7974), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n7215) );
  OR2_X1 U8934 ( .A1(n9570), .A2(n7207), .ZN(n7214) );
  OR2_X1 U8935 ( .A1(n7944), .A2(n7208), .ZN(n7213) );
  NAND2_X1 U8936 ( .A1(n7210), .A2(n7209), .ZN(n7211) );
  NAND2_X1 U8937 ( .A1(n7359), .A2(n7211), .ZN(n7479) );
  OR2_X1 U8938 ( .A1(n6593), .A2(n7479), .ZN(n7212) );
  OAI22_X1 U8939 ( .A1(n9531), .A2(n7323), .B1(n9529), .B2(n9596), .ZN(n7216)
         );
  AOI211_X1 U8940 ( .C1(n9511), .C2(n9848), .A(n9861), .B(n7216), .ZN(n7217)
         );
  OAI211_X1 U8941 ( .C1(n9595), .C2(n9544), .A(n7218), .B(n7217), .ZN(P1_U3229) );
  AOI21_X1 U8942 ( .B1(n9603), .B2(n7236), .A(n7219), .ZN(n10469) );
  OAI21_X1 U8943 ( .B1(n9603), .B2(n4507), .A(n7220), .ZN(n7224) );
  OAI22_X1 U8944 ( .A1(n7221), .A2(n10167), .B1(n7253), .B2(n10169), .ZN(n7223) );
  NOR2_X1 U8945 ( .A1(n10469), .A2(n6661), .ZN(n7222) );
  AOI211_X1 U8946 ( .C1(n10192), .C2(n7224), .A(n7223), .B(n7222), .ZN(n10467)
         );
  MUX2_X1 U8947 ( .A(n6224), .B(n10467), .S(n10170), .Z(n7231) );
  AOI21_X1 U8948 ( .B1(n4710), .B2(n7226), .A(n7225), .ZN(n10465) );
  OAI22_X1 U8949 ( .A1(n10182), .A2(n7228), .B1(n10157), .B2(n7227), .ZN(n7229) );
  AOI21_X1 U8950 ( .B1(n10465), .B2(n10195), .A(n7229), .ZN(n7230) );
  OAI211_X1 U8951 ( .C1(n10469), .C2(n10150), .A(n7231), .B(n7230), .ZN(
        P1_U3285) );
  NOR2_X1 U8952 ( .A1(n7232), .A2(n9849), .ZN(n7233) );
  AOI21_X1 U8953 ( .B1(n9703), .B2(n7234), .A(n7233), .ZN(n7235) );
  OR2_X2 U8954 ( .A1(n9590), .A2(n7242), .ZN(n9610) );
  NAND2_X1 U8955 ( .A1(n9590), .A2(n7242), .ZN(n9586) );
  NAND2_X1 U8956 ( .A1(n9610), .A2(n9586), .ZN(n9693) );
  NAND2_X1 U8957 ( .A1(n4498), .A2(n9693), .ZN(n7276) );
  NAND2_X1 U8958 ( .A1(n9590), .A2(n9848), .ZN(n7344) );
  NAND2_X1 U8959 ( .A1(n7276), .A2(n7344), .ZN(n7237) );
  OR2_X1 U8960 ( .A1(n7184), .A2(n9591), .ZN(n9612) );
  NAND2_X1 U8961 ( .A1(n7184), .A2(n9591), .ZN(n7427) );
  XNOR2_X1 U8962 ( .A(n7237), .B(n9708), .ZN(n7319) );
  AND2_X1 U8963 ( .A1(n5316), .A2(n7184), .ZN(n7238) );
  OR2_X1 U8964 ( .A1(n7238), .A2(n7438), .ZN(n7322) );
  OAI22_X1 U8965 ( .A1(n7322), .A2(n10458), .B1(n9595), .B2(n10480), .ZN(n7243) );
  AND2_X1 U8966 ( .A1(n9586), .A2(n7279), .ZN(n9733) );
  NAND2_X1 U8967 ( .A1(n7429), .A2(n9610), .ZN(n7240) );
  XNOR2_X1 U8968 ( .A(n7240), .B(n9708), .ZN(n7241) );
  OAI222_X1 U8969 ( .A1(n10167), .A2(n7242), .B1(n10169), .B2(n9596), .C1(
        n10165), .C2(n7241), .ZN(n7320) );
  AOI211_X1 U8970 ( .C1(n7319), .C2(n10476), .A(n7243), .B(n7320), .ZN(n7246)
         );
  NAND2_X1 U8971 ( .A1(n10486), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n7244) );
  OAI21_X1 U8972 ( .B1(n7246), .B2(n10486), .A(n7244), .ZN(P1_U3481) );
  NAND2_X1 U8973 ( .A1(n10496), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7245) );
  OAI21_X1 U8974 ( .B1(n7246), .B2(n10496), .A(n7245), .ZN(P1_U3532) );
  INV_X1 U8975 ( .A(n9590), .ZN(n10481) );
  INV_X1 U8976 ( .A(n7247), .ZN(n7252) );
  INV_X1 U8977 ( .A(n7248), .ZN(n7249) );
  OAI21_X1 U8978 ( .B1(n7249), .B2(n7252), .A(n7473), .ZN(n7250) );
  OAI211_X1 U8979 ( .C1(n7252), .C2(n7251), .A(n7250), .B(n9507), .ZN(n7257)
         );
  INV_X1 U8980 ( .A(n9591), .ZN(n9847) );
  OAI22_X1 U8981 ( .A1(n9554), .A2(n7253), .B1(n9531), .B2(n7285), .ZN(n7254)
         );
  AOI211_X1 U8982 ( .C1(n9551), .C2(n9847), .A(n7255), .B(n7254), .ZN(n7256)
         );
  OAI211_X1 U8983 ( .C1(n10481), .C2(n9544), .A(n7257), .B(n7256), .ZN(
        P1_U3219) );
  NAND2_X1 U8984 ( .A1(n7259), .A2(n7258), .ZN(n7289) );
  NAND2_X1 U8985 ( .A1(n7290), .A2(n7289), .ZN(n7260) );
  NAND2_X1 U8986 ( .A1(n7260), .A2(n8320), .ZN(n7445) );
  OAI21_X1 U8987 ( .B1(n7260), .B2(n8320), .A(n7445), .ZN(n10535) );
  INV_X1 U8988 ( .A(n10535), .ZN(n7275) );
  NOR2_X1 U8989 ( .A1(n7262), .A2(n7261), .ZN(n7264) );
  INV_X1 U8990 ( .A(n8370), .ZN(n7263) );
  NOR3_X1 U8991 ( .A1(n7264), .A2(n7263), .A3(n8320), .ZN(n7449) );
  INV_X1 U8992 ( .A(n7449), .ZN(n7266) );
  OAI21_X1 U8993 ( .B1(n7264), .B2(n7263), .A(n8320), .ZN(n7265) );
  NAND2_X1 U8994 ( .A1(n7266), .A2(n7265), .ZN(n7267) );
  INV_X1 U8995 ( .A(n7305), .ZN(n8524) );
  AOI222_X1 U8996 ( .A1(n8935), .A2(n7267), .B1(n8524), .B2(n8888), .C1(n8526), 
        .C2(n8886), .ZN(n10532) );
  MUX2_X1 U8997 ( .A(n7268), .B(n10532), .S(n8940), .Z(n7274) );
  NAND2_X1 U8998 ( .A1(n7269), .A2(n10529), .ZN(n7312) );
  OAI21_X1 U8999 ( .B1(n7269), .B2(n10529), .A(n7312), .ZN(n10531) );
  OAI22_X1 U9000 ( .A1(n8944), .A2(n10531), .B1(n7270), .B2(n8954), .ZN(n7271)
         );
  AOI21_X1 U9001 ( .B1(n8951), .B2(n7272), .A(n7271), .ZN(n7273) );
  OAI211_X1 U9002 ( .C1(n7275), .C2(n8899), .A(n7274), .B(n7273), .ZN(P2_U3290) );
  OAI21_X1 U9003 ( .B1(n4498), .B2(n9693), .A(n7276), .ZN(n10477) );
  INV_X1 U9004 ( .A(n5316), .ZN(n7277) );
  AOI211_X1 U9005 ( .C1(n9590), .C2(n7278), .A(n10458), .B(n7277), .ZN(n10478)
         );
  AOI22_X1 U9006 ( .A1(n10187), .A2(n9849), .B1(n9847), .B2(n10189), .ZN(n7283) );
  AOI21_X1 U9007 ( .B1(n9589), .B2(n9693), .A(n10165), .ZN(n7281) );
  OAI21_X1 U9008 ( .B1(n4399), .B2(n7429), .A(n7281), .ZN(n7282) );
  OAI211_X1 U9009 ( .C1(n10477), .C2(n6661), .A(n7283), .B(n7282), .ZN(n10482)
         );
  AOI21_X1 U9010 ( .B1(n10478), .B2(n10059), .A(n10482), .ZN(n7284) );
  MUX2_X1 U9011 ( .A(n6242), .B(n7284), .S(n10170), .Z(n7288) );
  INV_X1 U9012 ( .A(n7285), .ZN(n7286) );
  AOI22_X1 U9013 ( .A1(n10048), .A2(n9590), .B1(n10178), .B2(n7286), .ZN(n7287) );
  OAI211_X1 U9014 ( .C1(n10477), .C2(n10150), .A(n7288), .B(n7287), .ZN(
        P1_U3283) );
  NAND2_X1 U9015 ( .A1(n7451), .A2(n10529), .ZN(n7444) );
  NAND2_X1 U9016 ( .A1(n7290), .A2(n4462), .ZN(n7294) );
  INV_X1 U9017 ( .A(n7444), .ZN(n7292) );
  NAND2_X1 U9018 ( .A1(n7543), .A2(n7305), .ZN(n8379) );
  OAI21_X1 U9019 ( .B1(n8320), .B2(n7292), .A(n8321), .ZN(n7293) );
  NAND2_X1 U9020 ( .A1(n7291), .A2(n7305), .ZN(n7295) );
  OR2_X1 U9021 ( .A1(n7483), .A2(n7493), .ZN(n8385) );
  NAND2_X1 U9022 ( .A1(n7483), .A2(n7493), .ZN(n8386) );
  OAI21_X1 U9023 ( .B1(n7296), .B2(n8383), .A(n7485), .ZN(n7415) );
  AND2_X1 U9024 ( .A1(n8370), .A2(n7297), .ZN(n8369) );
  NAND3_X1 U9025 ( .A1(n7298), .A2(n8369), .A3(n8372), .ZN(n7301) );
  INV_X1 U9026 ( .A(n8321), .ZN(n8375) );
  NAND2_X1 U9027 ( .A1(n7299), .A2(n8372), .ZN(n7300) );
  NAND2_X1 U9028 ( .A1(n7301), .A2(n5318), .ZN(n7303) );
  AND2_X1 U9029 ( .A1(n7303), .A2(n8380), .ZN(n7304) );
  NAND2_X1 U9030 ( .A1(n7303), .A2(n7302), .ZN(n7491) );
  OAI21_X1 U9031 ( .B1(n7304), .B2(n8325), .A(n7491), .ZN(n7307) );
  OAI22_X1 U9032 ( .A1(n7582), .A2(n8926), .B1(n7305), .B2(n8924), .ZN(n7306)
         );
  AOI21_X1 U9033 ( .B1(n7307), .B2(n8935), .A(n7306), .ZN(n7309) );
  OR2_X1 U9034 ( .A1(n7415), .A2(n8931), .ZN(n7308) );
  NAND2_X1 U9035 ( .A1(n7309), .A2(n7308), .ZN(n7418) );
  INV_X1 U9036 ( .A(n7418), .ZN(n7311) );
  MUX2_X1 U9037 ( .A(n7311), .B(n7310), .S(n8949), .Z(n7318) );
  NAND2_X1 U9038 ( .A1(n7448), .A2(n7483), .ZN(n7313) );
  NAND2_X1 U9039 ( .A1(n7487), .A2(n7313), .ZN(n7417) );
  INV_X1 U9040 ( .A(n7417), .ZN(n7316) );
  INV_X1 U9041 ( .A(n7483), .ZN(n7416) );
  OAI22_X1 U9042 ( .A1(n8894), .A2(n7416), .B1(n8954), .B2(n7314), .ZN(n7315)
         );
  AOI21_X1 U9043 ( .B1(n7316), .B2(n8957), .A(n7315), .ZN(n7317) );
  OAI211_X1 U9044 ( .C1(n7415), .C2(n8920), .A(n7318), .B(n7317), .ZN(P2_U3288) );
  INV_X1 U9045 ( .A(n7319), .ZN(n7328) );
  INV_X1 U9046 ( .A(n7320), .ZN(n7321) );
  MUX2_X1 U9047 ( .A(n9236), .B(n7321), .S(n10170), .Z(n7327) );
  INV_X1 U9048 ( .A(n7322), .ZN(n7325) );
  OAI22_X1 U9049 ( .A1(n9595), .A2(n10182), .B1(n10157), .B2(n7323), .ZN(n7324) );
  AOI21_X1 U9050 ( .B1(n7325), .B2(n10195), .A(n7324), .ZN(n7326) );
  OAI211_X1 U9051 ( .C1(n10197), .C2(n7328), .A(n7327), .B(n7326), .ZN(
        P1_U3282) );
  INV_X1 U9052 ( .A(n7899), .ZN(n7330) );
  NAND2_X1 U9053 ( .A1(n9386), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7329) );
  OAI211_X1 U9054 ( .C1(n7330), .C2(n9120), .A(n8506), .B(n7329), .ZN(P2_U3335) );
  XNOR2_X1 U9055 ( .A(n7331), .B(n7332), .ZN(n7340) );
  INV_X1 U9056 ( .A(n7333), .ZN(n7659) );
  NAND2_X1 U9057 ( .A1(n8273), .A2(n7659), .ZN(n7334) );
  OAI21_X1 U9058 ( .B1(n8263), .B2(n7551), .A(n7334), .ZN(n7337) );
  OAI21_X1 U9059 ( .B1(n8277), .B2(n8156), .A(n7335), .ZN(n7336) );
  NOR2_X1 U9060 ( .A1(n7337), .A2(n7336), .ZN(n7339) );
  NAND2_X1 U9061 ( .A1(n8280), .A2(n9067), .ZN(n7338) );
  OAI211_X1 U9062 ( .C1(n7340), .C2(n8282), .A(n7339), .B(n7338), .ZN(P2_U3226) );
  NAND2_X1 U9063 ( .A1(n7899), .A2(n7341), .ZN(n7343) );
  NAND2_X1 U9064 ( .A1(n7342), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9830) );
  OAI211_X1 U9065 ( .C1(n7900), .C2(n8008), .A(n7343), .B(n9830), .ZN(P1_U3330) );
  OAI21_X1 U9066 ( .B1(n7184), .B2(n9847), .A(n9693), .ZN(n7348) );
  NAND2_X1 U9067 ( .A1(n7344), .A2(n9591), .ZN(n7346) );
  INV_X1 U9068 ( .A(n7344), .ZN(n7345) );
  AOI22_X1 U9069 ( .A1(n7184), .A2(n7346), .B1(n7345), .B2(n9847), .ZN(n7347)
         );
  NAND2_X1 U9070 ( .A1(n7349), .A2(n9677), .ZN(n7351) );
  AOI22_X1 U9071 ( .A1(n7859), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n7858), .B2(
        n9873), .ZN(n7350) );
  NAND2_X1 U9072 ( .A1(n7352), .A2(n9596), .ZN(n9618) );
  OR2_X1 U9073 ( .A1(n7352), .A2(n4701), .ZN(n7353) );
  NAND2_X1 U9074 ( .A1(n7354), .A2(n9677), .ZN(n7357) );
  AOI22_X1 U9075 ( .A1(n7858), .A2(n7355), .B1(n7859), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n7356) );
  NAND2_X1 U9076 ( .A1(n6788), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7365) );
  OR2_X1 U9077 ( .A1(n7944), .A2(n7358), .ZN(n7364) );
  INV_X1 U9078 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n9235) );
  NAND2_X1 U9079 ( .A1(n7359), .A2(n9235), .ZN(n7360) );
  NAND2_X1 U9080 ( .A1(n7370), .A2(n7360), .ZN(n7537) );
  OR2_X1 U9081 ( .A1(n6593), .A2(n7537), .ZN(n7363) );
  INV_X1 U9082 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7361) );
  OR2_X1 U9083 ( .A1(n6472), .A2(n7361), .ZN(n7362) );
  INV_X1 U9084 ( .A(n7981), .ZN(n7366) );
  AND2_X1 U9085 ( .A1(n5056), .A2(n7532), .ZN(n9624) );
  XNOR2_X1 U9086 ( .A(n7408), .B(n9711), .ZN(n10308) );
  NAND2_X1 U9087 ( .A1(n9618), .A2(n7427), .ZN(n7367) );
  NAND2_X1 U9088 ( .A1(n7367), .A2(n9611), .ZN(n9734) );
  XNOR2_X1 U9089 ( .A(n7389), .B(n9711), .ZN(n7378) );
  NAND2_X1 U9090 ( .A1(n7974), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n7376) );
  INV_X1 U9091 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7368) );
  OR2_X1 U9092 ( .A1(n7944), .A2(n7368), .ZN(n7375) );
  INV_X1 U9093 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7369) );
  NAND2_X1 U9094 ( .A1(n7370), .A2(n7369), .ZN(n7371) );
  NAND2_X1 U9095 ( .A1(n7394), .A2(n7371), .ZN(n9449) );
  OR2_X1 U9096 ( .A1(n6593), .A2(n9449), .ZN(n7374) );
  INV_X1 U9097 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7372) );
  OR2_X1 U9098 ( .A1(n9570), .A2(n7372), .ZN(n7373) );
  OAI22_X1 U9099 ( .A1(n9596), .A2(n10167), .B1(n8030), .B2(n10169), .ZN(n7377) );
  AOI21_X1 U9100 ( .B1(n7378), .B2(n10192), .A(n7377), .ZN(n7379) );
  OAI21_X1 U9101 ( .B1(n10308), .B2(n6661), .A(n7379), .ZN(n10311) );
  NAND2_X1 U9102 ( .A1(n10311), .A2(n10170), .ZN(n7384) );
  OAI22_X1 U9103 ( .A1(n10170), .A2(n6440), .B1(n7537), .B2(n10157), .ZN(n7382) );
  OR2_X1 U9104 ( .A1(n7439), .A2(n10309), .ZN(n7380) );
  NAND2_X1 U9105 ( .A1(n7402), .A2(n7380), .ZN(n10310) );
  NOR2_X1 U9106 ( .A1(n10310), .A2(n8000), .ZN(n7381) );
  AOI211_X1 U9107 ( .C1(n10048), .C2(n5056), .A(n7382), .B(n7381), .ZN(n7383)
         );
  OAI211_X1 U9108 ( .C1(n10308), .C2(n10150), .A(n7384), .B(n7383), .ZN(
        P1_U3280) );
  NAND2_X1 U9109 ( .A1(n7385), .A2(n9677), .ZN(n7388) );
  AOI22_X1 U9110 ( .A1(n7386), .A2(n7858), .B1(n7859), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n7387) );
  OR2_X1 U9111 ( .A1(n10303), .A2(n8030), .ZN(n9625) );
  NAND2_X1 U9112 ( .A1(n10303), .A2(n8030), .ZN(n9623) );
  INV_X1 U9113 ( .A(n7389), .ZN(n7391) );
  NAND2_X1 U9114 ( .A1(n7984), .A2(n7981), .ZN(n7392) );
  XOR2_X1 U9115 ( .A(n9707), .B(n7392), .Z(n7401) );
  NAND2_X1 U9116 ( .A1(n7974), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n7400) );
  INV_X1 U9117 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9348) );
  OR2_X1 U9118 ( .A1(n7944), .A2(n9348), .ZN(n7399) );
  NAND2_X1 U9119 ( .A1(n7394), .A2(n7393), .ZN(n7395) );
  NAND2_X1 U9120 ( .A1(n7812), .A2(n7395), .ZN(n10177) );
  OR2_X1 U9121 ( .A1(n6593), .A2(n10177), .ZN(n7398) );
  INV_X1 U9122 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7396) );
  OR2_X1 U9123 ( .A1(n9570), .A2(n7396), .ZN(n7397) );
  NAND4_X1 U9124 ( .A1(n7400), .A2(n7399), .A3(n7398), .A4(n7397), .ZN(n9845)
         );
  AOI222_X1 U9125 ( .A1(n10192), .A2(n7401), .B1(n9845), .B2(n10189), .C1(
        n9846), .C2(n10187), .ZN(n10305) );
  AOI21_X1 U9126 ( .B1(n7402), .B2(n10303), .A(n10458), .ZN(n7403) );
  AND2_X1 U9127 ( .A1(n7403), .A2(n10176), .ZN(n10302) );
  INV_X1 U9128 ( .A(n10303), .ZN(n7406) );
  NOR2_X1 U9129 ( .A1(n10157), .A2(n9449), .ZN(n7404) );
  AOI21_X1 U9130 ( .B1(n10180), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7404), .ZN(
        n7405) );
  OAI21_X1 U9131 ( .B1(n7406), .B2(n10182), .A(n7405), .ZN(n7407) );
  AOI21_X1 U9132 ( .B1(n10302), .B2(n10161), .A(n7407), .ZN(n7414) );
  INV_X1 U9133 ( .A(n10307), .ZN(n7412) );
  NAND2_X1 U9134 ( .A1(n7410), .A2(n9707), .ZN(n10301) );
  NAND3_X1 U9135 ( .A1(n7412), .A2(n7411), .A3(n10301), .ZN(n7413) );
  OAI211_X1 U9136 ( .C1(n10305), .C2(n10118), .A(n7414), .B(n7413), .ZN(
        P1_U3279) );
  INV_X1 U9137 ( .A(n9047), .ZN(n9062) );
  INV_X1 U9138 ( .A(n7415), .ZN(n7420) );
  OAI22_X1 U9139 ( .A1(n7417), .A2(n10530), .B1(n7416), .B2(n10528), .ZN(n7419) );
  AOI211_X1 U9140 ( .C1(n9062), .C2(n7420), .A(n7419), .B(n7418), .ZN(n7423)
         );
  NAND2_X1 U9141 ( .A1(n10542), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7421) );
  OAI21_X1 U9142 ( .B1(n7423), .B2(n10542), .A(n7421), .ZN(P2_U3528) );
  NAND2_X1 U9143 ( .A1(n10537), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n7422) );
  OAI21_X1 U9144 ( .B1(n7423), .B2(n10537), .A(n7422), .ZN(P2_U3475) );
  NAND2_X1 U9145 ( .A1(n7424), .A2(n9710), .ZN(n7425) );
  NAND2_X1 U9146 ( .A1(n7426), .A2(n7425), .ZN(n7432) );
  INV_X1 U9147 ( .A(n7432), .ZN(n10319) );
  INV_X1 U9148 ( .A(n7427), .ZN(n9588) );
  AOI21_X1 U9149 ( .B1(n7429), .B2(n7428), .A(n9588), .ZN(n7430) );
  XNOR2_X1 U9150 ( .A(n7430), .B(n9710), .ZN(n7436) );
  NAND2_X1 U9151 ( .A1(n7432), .A2(n7431), .ZN(n7435) );
  OAI22_X1 U9152 ( .A1(n7532), .A2(n10169), .B1(n9591), .B2(n10167), .ZN(n7433) );
  INV_X1 U9153 ( .A(n7433), .ZN(n7434) );
  OAI211_X1 U9154 ( .C1(n7436), .C2(n10165), .A(n7435), .B(n7434), .ZN(n10316)
         );
  MUX2_X1 U9155 ( .A(n10316), .B(P1_REG2_REG_10__SCAN_IN), .S(n10118), .Z(
        n7437) );
  INV_X1 U9156 ( .A(n7437), .ZN(n7443) );
  INV_X1 U9157 ( .A(n7438), .ZN(n7440) );
  AOI211_X1 U9158 ( .C1(n7352), .C2(n7440), .A(n10458), .B(n7439), .ZN(n10315)
         );
  OAI22_X1 U9159 ( .A1(n4702), .A2(n10182), .B1(n7479), .B2(n10157), .ZN(n7441) );
  AOI21_X1 U9160 ( .B1(n10315), .B2(n10161), .A(n7441), .ZN(n7442) );
  OAI211_X1 U9161 ( .C1(n10319), .C2(n10150), .A(n7443), .B(n7442), .ZN(
        P1_U3281) );
  NAND3_X1 U9162 ( .A1(n7445), .A2(n8375), .A3(n7444), .ZN(n7447) );
  NAND2_X1 U9163 ( .A1(n7447), .A2(n7446), .ZN(n7549) );
  OAI21_X1 U9164 ( .B1(n5265), .B2(n7291), .A(n7448), .ZN(n7545) );
  OAI22_X1 U9165 ( .A1(n7545), .A2(n10530), .B1(n7291), .B2(n10528), .ZN(n7453) );
  INV_X1 U9166 ( .A(n8376), .ZN(n8348) );
  NOR2_X1 U9167 ( .A1(n7449), .A2(n8348), .ZN(n7450) );
  XNOR2_X1 U9168 ( .A(n8375), .B(n7450), .ZN(n7452) );
  OAI222_X1 U9169 ( .A1(n8926), .A2(n7493), .B1(n7452), .B2(n7790), .C1(n8924), 
        .C2(n7451), .ZN(n7546) );
  AOI211_X1 U9170 ( .C1(n10536), .C2(n7549), .A(n7453), .B(n7546), .ZN(n7456)
         );
  NAND2_X1 U9171 ( .A1(n10537), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n7454) );
  OAI21_X1 U9172 ( .B1(n7456), .B2(n10537), .A(n7454), .ZN(P2_U3472) );
  NAND2_X1 U9173 ( .A1(n10542), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7455) );
  OAI21_X1 U9174 ( .B1(n7456), .B2(n10542), .A(n7455), .ZN(P2_U3527) );
  NAND4_X1 U9175 ( .A1(n7458), .A2(n7457), .A3(n4907), .A4(n7463), .ZN(n7472)
         );
  NAND2_X1 U9176 ( .A1(n7352), .A2(n8126), .ZN(n7460) );
  OR2_X1 U9177 ( .A1(n9596), .A2(n8127), .ZN(n7459) );
  NAND2_X1 U9178 ( .A1(n7460), .A2(n7459), .ZN(n7461) );
  XNOR2_X1 U9179 ( .A(n7461), .B(n8096), .ZN(n7530) );
  NOR2_X1 U9180 ( .A1(n8123), .A2(n9596), .ZN(n7462) );
  AOI21_X1 U9181 ( .B1(n7352), .B2(n8133), .A(n7462), .ZN(n7529) );
  XNOR2_X1 U9182 ( .A(n7530), .B(n7529), .ZN(n7476) );
  NOR2_X1 U9183 ( .A1(n7466), .A2(n7463), .ZN(n7464) );
  NAND2_X1 U9184 ( .A1(n7465), .A2(n7464), .ZN(n7469) );
  INV_X1 U9185 ( .A(n7466), .ZN(n7467) );
  AND3_X1 U9186 ( .A1(n7477), .A2(n7476), .A3(n4907), .ZN(n7478) );
  OAI21_X1 U9187 ( .B1(n7535), .B2(n7478), .A(n9507), .ZN(n7482) );
  AND2_X1 U9188 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9872) );
  OAI22_X1 U9189 ( .A1(n9554), .A2(n9591), .B1(n9531), .B2(n7479), .ZN(n7480)
         );
  AOI211_X1 U9190 ( .C1(n9551), .C2(n9846), .A(n9872), .B(n7480), .ZN(n7481)
         );
  OAI211_X1 U9191 ( .C1(n4702), .C2(n9544), .A(n7482), .B(n7481), .ZN(P1_U3215) );
  INV_X1 U9192 ( .A(n7493), .ZN(n8523) );
  NAND2_X1 U9193 ( .A1(n7483), .A2(n8523), .ZN(n7484) );
  OR2_X1 U9194 ( .A1(n7567), .A2(n7582), .ZN(n8391) );
  NAND2_X1 U9195 ( .A1(n7567), .A2(n7582), .ZN(n8389) );
  OAI21_X1 U9196 ( .B1(n7486), .B2(n7492), .A(n7553), .ZN(n7573) );
  INV_X1 U9197 ( .A(n7578), .ZN(n7489) );
  NAND2_X1 U9198 ( .A1(n7487), .A2(n7567), .ZN(n7488) );
  NAND2_X1 U9199 ( .A1(n7489), .A2(n7488), .ZN(n7569) );
  INV_X1 U9200 ( .A(n7567), .ZN(n7490) );
  OAI22_X1 U9201 ( .A1(n7569), .A2(n10530), .B1(n7490), .B2(n10528), .ZN(n7498) );
  XNOR2_X1 U9202 ( .A(n7556), .B(n7492), .ZN(n7497) );
  INV_X1 U9203 ( .A(n8931), .ZN(n7628) );
  NAND2_X1 U9204 ( .A1(n7573), .A2(n7628), .ZN(n7496) );
  OAI22_X1 U9205 ( .A1(n7554), .A2(n8926), .B1(n7493), .B2(n8924), .ZN(n7494)
         );
  INV_X1 U9206 ( .A(n7494), .ZN(n7495) );
  OAI211_X1 U9207 ( .C1(n7790), .C2(n7497), .A(n7496), .B(n7495), .ZN(n7570)
         );
  AOI211_X1 U9208 ( .C1(n9062), .C2(n7573), .A(n7498), .B(n7570), .ZN(n7501)
         );
  NAND2_X1 U9209 ( .A1(n10542), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7499) );
  OAI21_X1 U9210 ( .B1(n7501), .B2(n10542), .A(n7499), .ZN(P2_U3529) );
  NAND2_X1 U9211 ( .A1(n10537), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7500) );
  OAI21_X1 U9212 ( .B1(n7501), .B2(n10537), .A(n7500), .ZN(P2_U3478) );
  XNOR2_X1 U9213 ( .A(n7607), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n7506) );
  AOI21_X1 U9214 ( .B1(n7504), .B2(n7503), .A(n7502), .ZN(n7505) );
  NAND2_X1 U9215 ( .A1(n7505), .A2(n7506), .ZN(n7602) );
  OAI21_X1 U9216 ( .B1(n7506), .B2(n7505), .A(n7602), .ZN(n7513) );
  MUX2_X1 U9217 ( .A(n8939), .B(P2_REG2_REG_16__SCAN_IN), .S(n7607), .Z(n7509)
         );
  NAND2_X1 U9218 ( .A1(n4422), .A2(n7509), .ZN(n7606) );
  OAI211_X1 U9219 ( .C1(n4422), .C2(n7509), .A(n7606), .B(n8654), .ZN(n7511)
         );
  AND2_X1 U9220 ( .A1(P2_U3152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8208) );
  AOI21_X1 U9221 ( .B1(n8685), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8208), .ZN(
        n7510) );
  OAI211_X1 U9222 ( .C1(n8677), .C2(n7607), .A(n7511), .B(n7510), .ZN(n7512)
         );
  AOI21_X1 U9223 ( .B1(n8675), .B2(n7513), .A(n7512), .ZN(n7514) );
  INV_X1 U9224 ( .A(n7514), .ZN(P2_U3261) );
  XNOR2_X1 U9225 ( .A(n7515), .B(n7516), .ZN(n7524) );
  INV_X1 U9226 ( .A(n7637), .ZN(n7517) );
  NAND2_X1 U9227 ( .A1(n8273), .A2(n7517), .ZN(n7518) );
  OAI21_X1 U9228 ( .B1(n8263), .B2(n7626), .A(n7518), .ZN(n7521) );
  OAI21_X1 U9229 ( .B1(n8277), .B2(n7700), .A(n7519), .ZN(n7520) );
  NOR2_X1 U9230 ( .A1(n7521), .A2(n7520), .ZN(n7523) );
  NAND2_X1 U9231 ( .A1(n8280), .A2(n8407), .ZN(n7522) );
  OAI211_X1 U9232 ( .C1(n7524), .C2(n8282), .A(n7523), .B(n7522), .ZN(P2_U3236) );
  INV_X1 U9233 ( .A(n7911), .ZN(n7527) );
  OAI222_X1 U9234 ( .A1(P1_U3084), .A2(n7525), .B1(n8004), .B2(n7527), .C1(
        n7912), .C2(n8008), .ZN(P1_U3329) );
  OAI222_X1 U9235 ( .A1(n7528), .A2(P2_U3152), .B1(n9120), .B2(n7527), .C1(
        n7526), .C2(n9118), .ZN(P2_U3334) );
  AND2_X1 U9236 ( .A1(n7530), .A2(n7529), .ZN(n7534) );
  OAI22_X1 U9237 ( .A1(n10309), .A2(n8121), .B1(n7532), .B2(n8127), .ZN(n7531)
         );
  XNOR2_X1 U9238 ( .A(n7531), .B(n6504), .ZN(n8025) );
  OAI22_X1 U9239 ( .A1(n10309), .A2(n8127), .B1(n7532), .B2(n8123), .ZN(n8026)
         );
  XNOR2_X1 U9240 ( .A(n8025), .B(n8026), .ZN(n7533) );
  OAI21_X1 U9241 ( .B1(n7535), .B2(n7534), .A(n7533), .ZN(n7536) );
  NAND3_X1 U9242 ( .A1(n4617), .A2(n9507), .A3(n7536), .ZN(n7541) );
  OAI22_X1 U9243 ( .A1(n9554), .A2(n9596), .B1(n9531), .B2(n7537), .ZN(n7538)
         );
  AOI211_X1 U9244 ( .C1(n9551), .C2(n10188), .A(n7539), .B(n7538), .ZN(n7540)
         );
  OAI211_X1 U9245 ( .C1(n10309), .C2(n9544), .A(n7541), .B(n7540), .ZN(
        P1_U3234) );
  AOI22_X1 U9246 ( .A1(n8951), .A2(n7543), .B1(n7542), .B2(n8871), .ZN(n7544)
         );
  OAI21_X1 U9247 ( .B1(n8944), .B2(n7545), .A(n7544), .ZN(n7548) );
  MUX2_X1 U9248 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n7546), .S(n8940), .Z(n7547)
         );
  AOI211_X1 U9249 ( .C1(n8953), .C2(n7549), .A(n7548), .B(n7547), .ZN(n7550)
         );
  INV_X1 U9250 ( .A(n7550), .ZN(P2_U3289) );
  AND2_X1 U9251 ( .A1(n7561), .A2(n8520), .ZN(n7629) );
  INV_X1 U9252 ( .A(n7582), .ZN(n8522) );
  OR2_X1 U9253 ( .A1(n7567), .A2(n8522), .ZN(n7552) );
  NAND2_X1 U9254 ( .A1(n7645), .A2(n7554), .ZN(n8390) );
  NOR2_X1 U9255 ( .A1(n7622), .A2(n7575), .ZN(n7577) );
  INV_X1 U9256 ( .A(n7554), .ZN(n8521) );
  AND2_X1 U9257 ( .A1(n7645), .A2(n8521), .ZN(n7619) );
  NOR2_X1 U9258 ( .A1(n7577), .A2(n7619), .ZN(n7555) );
  XOR2_X1 U9259 ( .A(n8327), .B(n7555), .Z(n9080) );
  XNOR2_X1 U9260 ( .A(n7630), .B(n8327), .ZN(n7557) );
  INV_X1 U9261 ( .A(n7626), .ZN(n8519) );
  AOI222_X1 U9262 ( .A1(n8935), .A2(n7557), .B1(n8519), .B2(n8888), .C1(n8521), 
        .C2(n8886), .ZN(n9078) );
  MUX2_X1 U9263 ( .A(n7558), .B(n9078), .S(n8940), .Z(n7564) );
  INV_X1 U9264 ( .A(n7645), .ZN(n7579) );
  AOI21_X1 U9265 ( .B1(n9073), .B2(n7559), .A(n4572), .ZN(n9076) );
  OAI22_X1 U9266 ( .A1(n8894), .A2(n7561), .B1(n8954), .B2(n7560), .ZN(n7562)
         );
  AOI21_X1 U9267 ( .B1(n9076), .B2(n8957), .A(n7562), .ZN(n7563) );
  OAI211_X1 U9268 ( .C1(n9080), .C2(n8899), .A(n7564), .B(n7563), .ZN(P2_U3285) );
  INV_X1 U9269 ( .A(n8920), .ZN(n8946) );
  INV_X1 U9270 ( .A(n7565), .ZN(n7566) );
  AOI22_X1 U9271 ( .A1(n8951), .A2(n7567), .B1(n8871), .B2(n7566), .ZN(n7568)
         );
  OAI21_X1 U9272 ( .B1(n7569), .B2(n8944), .A(n7568), .ZN(n7572) );
  MUX2_X1 U9273 ( .A(n7570), .B(P2_REG2_REG_9__SCAN_IN), .S(n8958), .Z(n7571)
         );
  AOI211_X1 U9274 ( .C1(n8946), .C2(n7573), .A(n7572), .B(n7571), .ZN(n7574)
         );
  INV_X1 U9275 ( .A(n7574), .ZN(P2_U3287) );
  AND2_X1 U9276 ( .A1(n7622), .A2(n7575), .ZN(n7576) );
  OR2_X1 U9277 ( .A1(n7577), .A2(n7576), .ZN(n7587) );
  INV_X1 U9278 ( .A(n7587), .ZN(n7651) );
  OAI21_X1 U9279 ( .B1(n7578), .B2(n7579), .A(n7559), .ZN(n7647) );
  OAI22_X1 U9280 ( .A1(n7647), .A2(n10530), .B1(n7579), .B2(n10528), .ZN(n7588) );
  AOI21_X1 U9281 ( .B1(n7580), .B2(n8328), .A(n7790), .ZN(n7585) );
  NAND2_X1 U9282 ( .A1(n8520), .A2(n8888), .ZN(n7581) );
  OAI21_X1 U9283 ( .B1(n7582), .B2(n8924), .A(n7581), .ZN(n7583) );
  AOI21_X1 U9284 ( .B1(n7585), .B2(n7584), .A(n7583), .ZN(n7586) );
  OAI21_X1 U9285 ( .B1(n7587), .B2(n8931), .A(n7586), .ZN(n7648) );
  AOI211_X1 U9286 ( .C1(n9062), .C2(n7651), .A(n7588), .B(n7648), .ZN(n7591)
         );
  NAND2_X1 U9287 ( .A1(n10542), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7589) );
  OAI21_X1 U9288 ( .B1(n7591), .B2(n10542), .A(n7589), .ZN(P2_U3530) );
  NAND2_X1 U9289 ( .A1(n10537), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n7590) );
  OAI21_X1 U9290 ( .B1(n7591), .B2(n10537), .A(n7590), .ZN(P2_U3481) );
  XOR2_X1 U9291 ( .A(n9891), .B(n9883), .Z(n7594) );
  INV_X1 U9292 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7593) );
  AOI211_X1 U9293 ( .C1(n7594), .C2(n7593), .A(n9924), .B(n9884), .ZN(n7601)
         );
  INV_X1 U9294 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7825) );
  INV_X1 U9295 ( .A(n7806), .ZN(n7596) );
  OAI21_X1 U9296 ( .B1(n7596), .B2(P1_REG1_REG_14__SCAN_IN), .A(n7595), .ZN(
        n9889) );
  XOR2_X1 U9297 ( .A(n9891), .B(n9889), .Z(n7597) );
  NOR2_X1 U9298 ( .A1(n7597), .A2(n7825), .ZN(n9890) );
  AOI211_X1 U9299 ( .C1(n7825), .C2(n7597), .A(n9923), .B(n9890), .ZN(n7600)
         );
  NAND2_X1 U9300 ( .A1(n10418), .A2(n9891), .ZN(n7598) );
  NAND2_X1 U9301 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9552) );
  OAI211_X1 U9302 ( .C1(n10411), .C2(n4628), .A(n7598), .B(n9552), .ZN(n7599)
         );
  OR3_X1 U9303 ( .A1(n7601), .A2(n7600), .A3(n7599), .ZN(P1_U3256) );
  XNOR2_X1 U9304 ( .A(n7672), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n7605) );
  OAI21_X1 U9305 ( .B1(n7603), .B2(P2_REG1_REG_16__SCAN_IN), .A(n7602), .ZN(
        n7604) );
  NOR2_X1 U9306 ( .A1(n7604), .A2(n7605), .ZN(n7671) );
  AOI211_X1 U9307 ( .C1(n7605), .C2(n7604), .A(n8679), .B(n7671), .ZN(n7618)
         );
  INV_X1 U9308 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n7608) );
  MUX2_X1 U9309 ( .A(n7608), .B(P2_REG2_REG_17__SCAN_IN), .S(n7672), .Z(n7609)
         );
  INV_X1 U9310 ( .A(n7609), .ZN(n7610) );
  OAI211_X1 U9311 ( .C1(n7611), .C2(n7610), .A(n8654), .B(n7668), .ZN(n7615)
         );
  NOR2_X1 U9312 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7612), .ZN(n7613) );
  AOI21_X1 U9313 ( .B1(n8685), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n7613), .ZN(
        n7614) );
  OAI211_X1 U9314 ( .C1(n8677), .C2(n7616), .A(n7615), .B(n7614), .ZN(n7617)
         );
  OR2_X1 U9315 ( .A1(n7618), .A2(n7617), .ZN(P2_U3262) );
  NAND2_X1 U9316 ( .A1(n8328), .A2(n8327), .ZN(n7621) );
  AND2_X1 U9317 ( .A1(n9067), .A2(n7626), .ZN(n7631) );
  INV_X1 U9318 ( .A(n7631), .ZN(n8403) );
  NAND2_X1 U9319 ( .A1(n7624), .A2(n8406), .ZN(n7625) );
  OAI22_X1 U9320 ( .A1(n7700), .A2(n8926), .B1(n7626), .B2(n8924), .ZN(n7627)
         );
  AOI21_X1 U9321 ( .B1(n9063), .B2(n7628), .A(n7627), .ZN(n7634) );
  XNOR2_X1 U9322 ( .A(n7681), .B(n7680), .ZN(n7632) );
  NAND2_X1 U9323 ( .A1(n7632), .A2(n8935), .ZN(n7633) );
  NOR2_X1 U9324 ( .A1(n7635), .A2(n9059), .ZN(n7636) );
  OR2_X1 U9325 ( .A1(n7686), .A2(n7636), .ZN(n9060) );
  INV_X1 U9326 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7638) );
  OAI22_X1 U9327 ( .A1(n8940), .A2(n7638), .B1(n7637), .B2(n8954), .ZN(n7639)
         );
  AOI21_X1 U9328 ( .B1(n8951), .B2(n8407), .A(n7639), .ZN(n7640) );
  OAI21_X1 U9329 ( .B1(n9060), .B2(n8944), .A(n7640), .ZN(n7641) );
  AOI21_X1 U9330 ( .B1(n9063), .B2(n8946), .A(n7641), .ZN(n7642) );
  OAI21_X1 U9331 ( .B1(n9065), .B2(n8949), .A(n7642), .ZN(P2_U3283) );
  INV_X1 U9332 ( .A(n7643), .ZN(n7644) );
  AOI22_X1 U9333 ( .A1(n8951), .A2(n7645), .B1(n7644), .B2(n8871), .ZN(n7646)
         );
  OAI21_X1 U9334 ( .B1(n7647), .B2(n8944), .A(n7646), .ZN(n7650) );
  MUX2_X1 U9335 ( .A(n7648), .B(P2_REG2_REG_10__SCAN_IN), .S(n8949), .Z(n7649)
         );
  AOI211_X1 U9336 ( .C1(n7651), .C2(n8946), .A(n7650), .B(n7649), .ZN(n7652)
         );
  INV_X1 U9337 ( .A(n7652), .ZN(P2_U3286) );
  INV_X1 U9338 ( .A(n7924), .ZN(n7655) );
  OAI222_X1 U9339 ( .A1(P2_U3152), .A2(n7653), .B1(n9120), .B2(n7655), .C1(
        n9253), .C2(n9118), .ZN(P2_U3333) );
  OAI222_X1 U9340 ( .A1(n8008), .A2(n7925), .B1(n8004), .B2(n7655), .C1(
        P1_U3084), .C2(n7654), .ZN(P1_U3328) );
  XNOR2_X1 U9341 ( .A(n7656), .B(n8323), .ZN(n9066) );
  INV_X1 U9342 ( .A(n7635), .ZN(n7658) );
  NAND2_X1 U9343 ( .A1(n5327), .A2(n9067), .ZN(n7657) );
  NAND2_X1 U9344 ( .A1(n7658), .A2(n7657), .ZN(n9070) );
  AOI22_X1 U9345 ( .A1(n8951), .A2(n9067), .B1(n7659), .B2(n8871), .ZN(n7660)
         );
  OAI21_X1 U9346 ( .B1(n9070), .B2(n8944), .A(n7660), .ZN(n7666) );
  XNOR2_X1 U9347 ( .A(n7661), .B(n8323), .ZN(n7662) );
  NAND2_X1 U9348 ( .A1(n7662), .A2(n8935), .ZN(n7664) );
  AOI22_X1 U9349 ( .A1(n8518), .A2(n8888), .B1(n8886), .B2(n8520), .ZN(n7663)
         );
  NAND2_X1 U9350 ( .A1(n7664), .A2(n7663), .ZN(n9071) );
  MUX2_X1 U9351 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n9071), .S(n8940), .Z(n7665)
         );
  AOI211_X1 U9352 ( .C1(n9066), .C2(n8953), .A(n7666), .B(n7665), .ZN(n7667)
         );
  INV_X1 U9353 ( .A(n7667), .ZN(P2_U3284) );
  NAND2_X1 U9354 ( .A1(n7672), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7669) );
  NAND2_X1 U9355 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n7670), .ZN(n8668) );
  OAI211_X1 U9356 ( .C1(n7670), .C2(P2_REG2_REG_18__SCAN_IN), .A(n8654), .B(
        n8668), .ZN(n7677) );
  INV_X1 U9357 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9251) );
  XNOR2_X1 U9358 ( .A(n8670), .B(n9251), .ZN(n8673) );
  AOI21_X1 U9359 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n7672), .A(n7671), .ZN(
        n8672) );
  XNOR2_X1 U9360 ( .A(n8673), .B(n8672), .ZN(n7675) );
  INV_X1 U9361 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10584) );
  NAND2_X1 U9362 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8252) );
  OAI21_X1 U9363 ( .B1(n7673), .B2(n10584), .A(n8252), .ZN(n7674) );
  AOI21_X1 U9364 ( .B1(n8675), .B2(n7675), .A(n7674), .ZN(n7676) );
  OAI211_X1 U9365 ( .C1(n8677), .C2(n4764), .A(n7677), .B(n7676), .ZN(P2_U3263) );
  NAND2_X1 U9366 ( .A1(n8407), .A2(n8518), .ZN(n7678) );
  NAND2_X1 U9367 ( .A1(n9054), .A2(n7700), .ZN(n8419) );
  NAND2_X1 U9368 ( .A1(n8413), .A2(n8419), .ZN(n8411) );
  XNOR2_X1 U9369 ( .A(n7701), .B(n8411), .ZN(n9058) );
  AOI21_X1 U9370 ( .B1(n7682), .B2(n8411), .A(n7790), .ZN(n7685) );
  OAI22_X1 U9371 ( .A1(n8925), .A2(n8926), .B1(n8156), .B2(n8924), .ZN(n7684)
         );
  AOI21_X1 U9372 ( .B1(n7685), .B2(n7694), .A(n7684), .ZN(n9057) );
  OR2_X1 U9373 ( .A1(n9057), .A2(n8949), .ZN(n7693) );
  INV_X1 U9374 ( .A(n9054), .ZN(n7690) );
  OR2_X1 U9375 ( .A1(n7686), .A2(n7690), .ZN(n7687) );
  AND2_X1 U9376 ( .A1(n7704), .A2(n7687), .ZN(n9055) );
  NOR2_X1 U9377 ( .A1(n8954), .A2(n8157), .ZN(n7688) );
  AOI21_X1 U9378 ( .B1(n8958), .B2(P2_REG2_REG_14__SCAN_IN), .A(n7688), .ZN(
        n7689) );
  OAI21_X1 U9379 ( .B1(n7690), .B2(n8894), .A(n7689), .ZN(n7691) );
  AOI21_X1 U9380 ( .B1(n9055), .B2(n8957), .A(n7691), .ZN(n7692) );
  OAI211_X1 U9381 ( .C1(n9058), .C2(n8899), .A(n7693), .B(n7692), .ZN(P2_U3282) );
  INV_X1 U9382 ( .A(n7697), .ZN(n7696) );
  NAND2_X1 U9383 ( .A1(n9049), .A2(n8925), .ZN(n7695) );
  AOI21_X1 U9384 ( .B1(n7696), .B2(n7702), .A(n7790), .ZN(n7699) );
  OAI22_X1 U9385 ( .A1(n8278), .A2(n8926), .B1(n7700), .B2(n8924), .ZN(n7698)
         );
  AOI21_X1 U9386 ( .B1(n7699), .B2(n7781), .A(n7698), .ZN(n9052) );
  INV_X1 U9387 ( .A(n7700), .ZN(n8517) );
  OAI21_X1 U9388 ( .B1(n7703), .B2(n7702), .A(n7760), .ZN(n9048) );
  INV_X1 U9389 ( .A(n5322), .ZN(n7705) );
  AOI21_X1 U9390 ( .B1(n9049), .B2(n7704), .A(n7705), .ZN(n9050) );
  NAND2_X1 U9391 ( .A1(n9050), .A2(n8957), .ZN(n7707) );
  AOI22_X1 U9392 ( .A1(n8958), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8272), .B2(
        n8871), .ZN(n7706) );
  OAI211_X1 U9393 ( .C1(n4778), .C2(n8894), .A(n7707), .B(n7706), .ZN(n7708)
         );
  AOI21_X1 U9394 ( .B1(n9048), .B2(n8953), .A(n7708), .ZN(n7709) );
  OAI21_X1 U9395 ( .B1(n9052), .B2(n8949), .A(n7709), .ZN(P2_U3281) );
  INV_X1 U9396 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9679) );
  INV_X1 U9397 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7714) );
  INV_X1 U9398 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8007) );
  MUX2_X1 U9399 ( .A(n7714), .B(n8007), .S(n4395), .Z(n7716) );
  XNOR2_X1 U9400 ( .A(n7716), .B(SI_28_), .ZN(n7724) );
  INV_X1 U9401 ( .A(SI_28_), .ZN(n7715) );
  NAND2_X1 U9402 ( .A1(n7716), .A2(n7715), .ZN(n7717) );
  MUX2_X1 U9403 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n4396), .Z(n8009) );
  INV_X1 U9404 ( .A(SI_29_), .ZN(n9317) );
  XNOR2_X1 U9405 ( .A(n8009), .B(n9317), .ZN(n7719) );
  INV_X1 U9406 ( .A(n9678), .ZN(n9110) );
  OAI222_X1 U9407 ( .A1(n8008), .A2(n9679), .B1(P1_U3084), .B2(n7720), .C1(
        n8004), .C2(n9110), .ZN(P1_U3324) );
  INV_X1 U9408 ( .A(n7893), .ZN(n7723) );
  OAI222_X1 U9409 ( .A1(n8008), .A2(n7894), .B1(n8004), .B2(n7723), .C1(
        P1_U3084), .C2(n7721), .ZN(P1_U3331) );
  OAI222_X1 U9410 ( .A1(n8339), .A2(P2_U3152), .B1(n9120), .B2(n7723), .C1(
        n7722), .C2(n9118), .ZN(P2_U3336) );
  NAND2_X1 U9411 ( .A1(n8006), .A2(n8307), .ZN(n7727) );
  NAND2_X1 U9412 ( .A1(n8308), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n7726) );
  OR2_X1 U9413 ( .A1(n8710), .A2(n4796), .ZN(n7730) );
  XNOR2_X1 U9414 ( .A(n4746), .B(n7730), .ZN(n7738) );
  INV_X1 U9415 ( .A(n7738), .ZN(n7736) );
  NOR2_X1 U9416 ( .A1(n7732), .A2(n7731), .ZN(n7733) );
  AOI21_X1 U9417 ( .B1(n8978), .B2(n8280), .A(n7733), .ZN(n7740) );
  INV_X1 U9418 ( .A(n7740), .ZN(n7735) );
  NAND3_X1 U9419 ( .A1(n8978), .A2(n10528), .A3(n7736), .ZN(n7734) );
  OAI211_X1 U9420 ( .C1(n8978), .C2(n7736), .A(n7735), .B(n7734), .ZN(n7757)
         );
  NAND3_X1 U9421 ( .A1(n8978), .A2(n7738), .A3(n10528), .ZN(n7737) );
  OAI21_X1 U9422 ( .B1(n7738), .B2(n8978), .A(n7737), .ZN(n7739) );
  NOR3_X1 U9423 ( .A1(n7740), .A2(n7741), .A3(n7739), .ZN(n7755) );
  INV_X1 U9424 ( .A(n7741), .ZN(n7753) );
  NOR2_X1 U9425 ( .A1(n8742), .A2(n8263), .ZN(n7751) );
  INV_X1 U9426 ( .A(n7742), .ZN(n8703) );
  INV_X1 U9427 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n9320) );
  NAND2_X1 U9428 ( .A1(n7743), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n7745) );
  NAND2_X1 U9429 ( .A1(n8288), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n7744) );
  OAI211_X1 U9430 ( .C1(n5826), .C2(n9320), .A(n7745), .B(n7744), .ZN(n7746)
         );
  AOI21_X1 U9431 ( .B1(n8703), .B2(n7747), .A(n7746), .ZN(n8508) );
  NAND2_X1 U9432 ( .A1(P2_U3152), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n7749) );
  NAND2_X1 U9433 ( .A1(n7777), .A2(n8273), .ZN(n7748) );
  OAI211_X1 U9434 ( .C1(n8508), .C2(n8277), .A(n7749), .B(n7748), .ZN(n7750)
         );
  NOR2_X1 U9435 ( .A1(n7751), .A2(n7750), .ZN(n7752) );
  OAI21_X1 U9436 ( .B1(n7757), .B2(n7753), .A(n7752), .ZN(n7754) );
  AOI21_X1 U9437 ( .B1(n7758), .B2(n7755), .A(n7754), .ZN(n7756) );
  INV_X1 U9438 ( .A(n8925), .ZN(n8516) );
  OR2_X1 U9439 ( .A1(n9049), .A2(n8516), .ZN(n7759) );
  NAND2_X1 U9440 ( .A1(n8942), .A2(n8278), .ZN(n8421) );
  OR2_X1 U9441 ( .A1(n9037), .A2(n8927), .ZN(n7784) );
  NAND2_X1 U9442 ( .A1(n9037), .A2(n8927), .ZN(n8422) );
  INV_X1 U9443 ( .A(n8903), .ZN(n8907) );
  NAND2_X1 U9444 ( .A1(n8942), .A2(n8515), .ZN(n8902) );
  AND2_X1 U9445 ( .A1(n8907), .A2(n8902), .ZN(n7761) );
  INV_X1 U9446 ( .A(n8927), .ZN(n8887) );
  OR2_X1 U9447 ( .A1(n9037), .A2(n8887), .ZN(n7762) );
  INV_X1 U9448 ( .A(n8214), .ZN(n8865) );
  NOR2_X1 U9449 ( .A1(n9032), .A2(n8865), .ZN(n7763) );
  INV_X1 U9450 ( .A(n9032), .ZN(n8895) );
  AND2_X1 U9451 ( .A1(n9028), .A2(n8889), .ZN(n7765) );
  OR2_X1 U9452 ( .A1(n9028), .A2(n8889), .ZN(n7764) );
  NAND2_X1 U9453 ( .A1(n9022), .A2(n8182), .ZN(n8442) );
  NAND2_X1 U9454 ( .A1(n8441), .A2(n8442), .ZN(n8857) );
  INV_X1 U9455 ( .A(n8182), .ZN(n8866) );
  OR2_X1 U9456 ( .A1(n9015), .A2(n8513), .ZN(n7766) );
  NAND2_X1 U9457 ( .A1(n9015), .A2(n8513), .ZN(n7767) );
  AND2_X1 U9458 ( .A1(n9010), .A2(n8453), .ZN(n7786) );
  INV_X1 U9459 ( .A(n7786), .ZN(n8444) );
  NAND2_X1 U9460 ( .A1(n9005), .A2(n8824), .ZN(n8447) );
  NAND2_X1 U9461 ( .A1(n8459), .A2(n8447), .ZN(n8803) );
  INV_X1 U9462 ( .A(n8803), .ZN(n8795) );
  INV_X1 U9463 ( .A(n8824), .ZN(n8512) );
  NAND2_X1 U9464 ( .A1(n9005), .A2(n8512), .ZN(n7769) );
  NAND2_X1 U9465 ( .A1(n9000), .A2(n8192), .ZN(n8462) );
  INV_X1 U9466 ( .A(n8192), .ZN(n8799) );
  OR2_X1 U9467 ( .A1(n9000), .A2(n8799), .ZN(n7770) );
  NAND2_X1 U9468 ( .A1(n8772), .A2(n7770), .ZN(n8757) );
  NAND2_X1 U9469 ( .A1(n8996), .A2(n8741), .ZN(n8468) );
  INV_X1 U9470 ( .A(n8741), .ZN(n8511) );
  OR2_X1 U9471 ( .A1(n8996), .A2(n8511), .ZN(n7771) );
  NAND2_X1 U9472 ( .A1(n8756), .A2(n7771), .ZN(n8733) );
  NAND2_X1 U9473 ( .A1(n8746), .A2(n8193), .ZN(n8472) );
  NAND2_X1 U9474 ( .A1(n8724), .A2(n8742), .ZN(n7773) );
  NAND2_X1 U9475 ( .A1(n8978), .A2(n8710), .ZN(n8478) );
  AND2_X2 U9476 ( .A1(n8479), .A2(n8478), .ZN(n8476) );
  INV_X1 U9477 ( .A(n9010), .ZN(n8820) );
  INV_X1 U9478 ( .A(n9005), .ZN(n8811) );
  INV_X1 U9479 ( .A(n9000), .ZN(n8782) );
  INV_X1 U9480 ( .A(n8720), .ZN(n7776) );
  INV_X1 U9481 ( .A(n8700), .ZN(n7775) );
  AOI21_X1 U9482 ( .B1(n8978), .B2(n7776), .A(n7775), .ZN(n8979) );
  AOI22_X1 U9483 ( .A1(n7777), .A2(n8871), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n8949), .ZN(n7778) );
  OAI21_X1 U9484 ( .B1(n7779), .B2(n8894), .A(n7778), .ZN(n7792) );
  INV_X1 U9485 ( .A(n8935), .ZN(n7790) );
  OR2_X1 U9486 ( .A1(n9032), .A2(n8214), .ZN(n8438) );
  NAND2_X1 U9487 ( .A1(n9032), .A2(n8214), .ZN(n8431) );
  NAND2_X1 U9488 ( .A1(n8438), .A2(n8431), .ZN(n8882) );
  INV_X1 U9489 ( .A(n7784), .ZN(n8883) );
  NOR2_X1 U9490 ( .A1(n8882), .A2(n8883), .ZN(n7785) );
  OR2_X1 U9491 ( .A1(n9028), .A2(n8848), .ZN(n8440) );
  NAND2_X1 U9492 ( .A1(n9028), .A2(n8848), .ZN(n8846) );
  INV_X1 U9493 ( .A(n8846), .ZN(n8437) );
  OR2_X1 U9494 ( .A1(n9015), .A2(n8850), .ZN(n8434) );
  OAI211_X1 U9495 ( .C1(n8823), .C2(n7786), .A(n8459), .B(n8794), .ZN(n7787)
         );
  AND2_X1 U9496 ( .A1(n7787), .A2(n8447), .ZN(n7788) );
  NOR2_X1 U9497 ( .A1(n8981), .A2(n8949), .ZN(n7791) );
  AOI211_X1 U9498 ( .C1(n8957), .C2(n8979), .A(n7792), .B(n7791), .ZN(n7793)
         );
  OAI21_X1 U9499 ( .B1(n8983), .B2(n8899), .A(n7793), .ZN(P2_U3268) );
  NAND2_X1 U9500 ( .A1(n7794), .A2(n9507), .ZN(n7798) );
  AOI22_X1 U9501 ( .A1(n9556), .A2(n7796), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n7795), .ZN(n7797) );
  OAI211_X1 U9502 ( .C1(n6655), .C2(n9529), .A(n7798), .B(n7797), .ZN(P1_U3230) );
  NAND2_X1 U9503 ( .A1(n7799), .A2(n9677), .ZN(n7802) );
  AOI22_X1 U9504 ( .A1(n7800), .A2(n7858), .B1(n7859), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n7801) );
  NOR2_X1 U9505 ( .A1(n10295), .A2(n9845), .ZN(n7803) );
  NAND2_X1 U9506 ( .A1(n7804), .A2(n9677), .ZN(n7809) );
  INV_X1 U9507 ( .A(n7807), .ZN(n7808) );
  NAND2_X1 U9508 ( .A1(n7974), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n7817) );
  OR2_X1 U9509 ( .A1(n9570), .A2(n7154), .ZN(n7816) );
  INV_X1 U9510 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7810) );
  OR2_X1 U9511 ( .A1(n7944), .A2(n7810), .ZN(n7815) );
  INV_X1 U9512 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7811) );
  NAND2_X1 U9513 ( .A1(n7812), .A2(n7811), .ZN(n7813) );
  NAND2_X1 U9514 ( .A1(n7823), .A2(n7813), .ZN(n10158) );
  OR2_X1 U9515 ( .A1(n6593), .A2(n10158), .ZN(n7814) );
  NOR2_X1 U9516 ( .A1(n10156), .A2(n10138), .ZN(n7818) );
  NAND2_X1 U9517 ( .A1(n7819), .A2(n9677), .ZN(n7821) );
  AOI22_X1 U9518 ( .A1(n7859), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n7858), .B2(
        n9891), .ZN(n7820) );
  NAND2_X1 U9519 ( .A1(n7823), .A2(n7822), .ZN(n7824) );
  AND2_X1 U9520 ( .A1(n7836), .A2(n7824), .ZN(n10147) );
  NAND2_X1 U9521 ( .A1(n7955), .A2(n10147), .ZN(n7830) );
  OR2_X1 U9522 ( .A1(n7944), .A2(n7825), .ZN(n7829) );
  INV_X1 U9523 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n7826) );
  OR2_X1 U9524 ( .A1(n6472), .A2(n7826), .ZN(n7828) );
  OR2_X1 U9525 ( .A1(n9570), .A2(n7593), .ZN(n7827) );
  NAND4_X1 U9526 ( .A1(n7830), .A2(n7829), .A3(n7828), .A4(n7827), .ZN(n9844)
         );
  NOR2_X1 U9527 ( .A1(n10285), .A2(n9844), .ZN(n7831) );
  AOI22_X1 U9528 ( .A1(n7859), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n7858), .B2(
        n9906), .ZN(n7833) );
  INV_X1 U9529 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9352) );
  OR2_X1 U9530 ( .A1(n7944), .A2(n9352), .ZN(n7835) );
  INV_X1 U9531 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n10128) );
  OR2_X1 U9532 ( .A1(n9570), .A2(n10128), .ZN(n7834) );
  AND2_X1 U9533 ( .A1(n7835), .A2(n7834), .ZN(n7840) );
  INV_X1 U9534 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9473) );
  NAND2_X1 U9535 ( .A1(n7836), .A2(n9473), .ZN(n7837) );
  NAND2_X1 U9536 ( .A1(n7844), .A2(n7837), .ZN(n10127) );
  OR2_X1 U9537 ( .A1(n10127), .A2(n6593), .ZN(n7839) );
  INV_X1 U9538 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9316) );
  OR2_X1 U9539 ( .A1(n6472), .A2(n9316), .ZN(n7838) );
  NAND2_X1 U9540 ( .A1(n10282), .A2(n10139), .ZN(n9636) );
  NAND2_X1 U9541 ( .A1(n7841), .A2(n9677), .ZN(n7843) );
  AOI22_X1 U9542 ( .A1(n7859), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n7858), .B2(
        n9920), .ZN(n7842) );
  NAND2_X1 U9543 ( .A1(n7844), .A2(n9481), .ZN(n7845) );
  NAND2_X1 U9544 ( .A1(n7852), .A2(n7845), .ZN(n10109) );
  AOI22_X1 U9545 ( .A1(n6788), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n6466), .B2(
        P1_REG1_REG_17__SCAN_IN), .ZN(n7847) );
  NAND2_X1 U9546 ( .A1(n7974), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n7846) );
  OAI211_X1 U9547 ( .C1(n10109), .C2(n6593), .A(n7847), .B(n7846), .ZN(n10102)
         );
  INV_X1 U9548 ( .A(n10275), .ZN(n10112) );
  INV_X1 U9549 ( .A(n10102), .ZN(n10134) );
  NAND2_X1 U9550 ( .A1(n7848), .A2(n9677), .ZN(n7850) );
  AOI22_X1 U9551 ( .A1(n7859), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n7858), .B2(
        n10417), .ZN(n7849) );
  INV_X1 U9552 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n7851) );
  NAND2_X1 U9553 ( .A1(n7852), .A2(n7851), .ZN(n7853) );
  NAND2_X1 U9554 ( .A1(n7871), .A2(n7853), .ZN(n10094) );
  OR2_X1 U9555 ( .A1(n10094), .A2(n6593), .ZN(n7856) );
  AOI22_X1 U9556 ( .A1(n6788), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n6466), .B2(
        P1_REG1_REG_18__SCAN_IN), .ZN(n7855) );
  NAND2_X1 U9557 ( .A1(n7974), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n7854) );
  NAND2_X1 U9558 ( .A1(n10270), .A2(n9482), .ZN(n9760) );
  NAND2_X1 U9559 ( .A1(n9643), .A2(n9760), .ZN(n10100) );
  INV_X1 U9560 ( .A(n9482), .ZN(n10116) );
  NAND2_X1 U9561 ( .A1(n7857), .A2(n9677), .ZN(n7861) );
  AOI22_X1 U9562 ( .A1(n7859), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n10007), 
        .B2(n7858), .ZN(n7860) );
  XNOR2_X1 U9563 ( .A(n7871), .B(P1_REG3_REG_19__SCAN_IN), .ZN(n10082) );
  NAND2_X1 U9564 ( .A1(n10082), .A2(n7955), .ZN(n7866) );
  INV_X1 U9565 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9369) );
  NAND2_X1 U9566 ( .A1(n6788), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n7863) );
  NAND2_X1 U9567 ( .A1(n7974), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n7862) );
  OAI211_X1 U9568 ( .C1(n7944), .C2(n9369), .A(n7863), .B(n7862), .ZN(n7864)
         );
  INV_X1 U9569 ( .A(n7864), .ZN(n7865) );
  NAND2_X1 U9570 ( .A1(n7866), .A2(n7865), .ZN(n10103) );
  NAND2_X1 U9571 ( .A1(n7867), .A2(n9677), .ZN(n7870) );
  OR2_X1 U9572 ( .A1(n9680), .A2(n7868), .ZN(n7869) );
  INV_X1 U9573 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9433) );
  INV_X1 U9574 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9498) );
  OAI21_X1 U9575 ( .B1(n7871), .B2(n9433), .A(n9498), .ZN(n7872) );
  AND2_X1 U9576 ( .A1(n7872), .A2(n7884), .ZN(n10069) );
  NAND2_X1 U9577 ( .A1(n10069), .A2(n7955), .ZN(n7878) );
  INV_X1 U9578 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n7875) );
  NAND2_X1 U9579 ( .A1(n6788), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n7874) );
  NAND2_X1 U9580 ( .A1(n6466), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n7873) );
  OAI211_X1 U9581 ( .C1(n7875), .C2(n6472), .A(n7874), .B(n7873), .ZN(n7876)
         );
  INV_X1 U9582 ( .A(n7876), .ZN(n7877) );
  NAND2_X1 U9583 ( .A1(n7880), .A2(n9677), .ZN(n7883) );
  OR2_X1 U9584 ( .A1(n9680), .A2(n7881), .ZN(n7882) );
  INV_X1 U9585 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9372) );
  NAND2_X1 U9586 ( .A1(n7884), .A2(n9372), .ZN(n7885) );
  NAND2_X1 U9587 ( .A1(n7903), .A2(n7885), .ZN(n10061) );
  OR2_X1 U9588 ( .A1(n10061), .A2(n6593), .ZN(n7890) );
  INV_X1 U9589 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9196) );
  NAND2_X1 U9590 ( .A1(n6466), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n7887) );
  NAND2_X1 U9591 ( .A1(n7974), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n7886) );
  OAI211_X1 U9592 ( .C1(n9196), .C2(n9570), .A(n7887), .B(n7886), .ZN(n7888)
         );
  INV_X1 U9593 ( .A(n7888), .ZN(n7889) );
  NAND2_X1 U9594 ( .A1(n10256), .A2(n9521), .ZN(n9655) );
  NAND2_X1 U9595 ( .A1(n10046), .A2(n10047), .ZN(n7892) );
  NAND2_X1 U9596 ( .A1(n10256), .A2(n10074), .ZN(n7891) );
  NAND2_X1 U9597 ( .A1(n7892), .A2(n7891), .ZN(n10030) );
  NAND2_X1 U9598 ( .A1(n7893), .A2(n9677), .ZN(n7896) );
  OR2_X1 U9599 ( .A1(n9680), .A2(n7894), .ZN(n7895) );
  NOR2_X1 U9600 ( .A1(n10035), .A2(n10055), .ZN(n7898) );
  NAND2_X1 U9601 ( .A1(n10035), .A2(n10055), .ZN(n7897) );
  NAND2_X1 U9602 ( .A1(n7899), .A2(n9677), .ZN(n7902) );
  OR2_X1 U9603 ( .A1(n9680), .A2(n7900), .ZN(n7901) );
  INV_X1 U9604 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9519) );
  INV_X1 U9605 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9420) );
  OAI21_X1 U9606 ( .B1(n7903), .B2(n9519), .A(n9420), .ZN(n7904) );
  AND2_X1 U9607 ( .A1(n7904), .A2(n7915), .ZN(n10018) );
  NAND2_X1 U9608 ( .A1(n10018), .A2(n7955), .ZN(n7909) );
  INV_X1 U9609 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9222) );
  NAND2_X1 U9610 ( .A1(n6466), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n7906) );
  NAND2_X1 U9611 ( .A1(n6788), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n7905) );
  OAI211_X1 U9612 ( .C1(n9222), .C2(n6472), .A(n7906), .B(n7905), .ZN(n7907)
         );
  INV_X1 U9613 ( .A(n7907), .ZN(n7908) );
  NOR2_X1 U9614 ( .A1(n10248), .A2(n10041), .ZN(n7910) );
  NAND2_X1 U9615 ( .A1(n10248), .A2(n10041), .ZN(n9578) );
  NAND2_X1 U9616 ( .A1(n7911), .A2(n9677), .ZN(n7914) );
  OR2_X1 U9617 ( .A1(n9680), .A2(n7912), .ZN(n7913) );
  INV_X1 U9618 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9188) );
  NAND2_X1 U9619 ( .A1(n7915), .A2(n9188), .ZN(n7916) );
  NAND2_X1 U9620 ( .A1(n7930), .A2(n7916), .ZN(n10006) );
  INV_X1 U9621 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n7919) );
  NAND2_X1 U9622 ( .A1(n6466), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n7918) );
  NAND2_X1 U9623 ( .A1(n7974), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n7917) );
  OAI211_X1 U9624 ( .C1(n7919), .C2(n9570), .A(n7918), .B(n7917), .ZN(n7920)
         );
  INV_X1 U9625 ( .A(n7920), .ZN(n7921) );
  NOR2_X1 U9626 ( .A1(n9577), .A2(n10025), .ZN(n7923) );
  NAND2_X1 U9627 ( .A1(n7924), .A2(n9677), .ZN(n7927) );
  OR2_X1 U9628 ( .A1(n9680), .A2(n7925), .ZN(n7926) );
  INV_X1 U9629 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n7929) );
  NAND2_X1 U9630 ( .A1(n7930), .A2(n7929), .ZN(n7931) );
  NAND2_X1 U9631 ( .A1(n7942), .A2(n7931), .ZN(n9998) );
  INV_X1 U9632 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9319) );
  NAND2_X1 U9633 ( .A1(n6466), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n7933) );
  NAND2_X1 U9634 ( .A1(n6788), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n7932) );
  OAI211_X1 U9635 ( .C1(n6472), .C2(n9319), .A(n7933), .B(n7932), .ZN(n7934)
         );
  INV_X1 U9636 ( .A(n7934), .ZN(n7935) );
  NAND2_X1 U9637 ( .A1(n10238), .A2(n10013), .ZN(n9665) );
  NAND2_X1 U9638 ( .A1(n8111), .A2(n10013), .ZN(n7937) );
  OR2_X1 U9639 ( .A1(n9680), .A2(n10352), .ZN(n7939) );
  INV_X1 U9640 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n7941) );
  NAND2_X1 U9641 ( .A1(n7942), .A2(n7941), .ZN(n7943) );
  NAND2_X1 U9642 ( .A1(n9982), .A2(n7955), .ZN(n7950) );
  INV_X1 U9643 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n7947) );
  NAND2_X1 U9644 ( .A1(n7974), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n7946) );
  INV_X1 U9645 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9283) );
  OR2_X1 U9646 ( .A1(n7944), .A2(n9283), .ZN(n7945) );
  OAI211_X1 U9647 ( .C1(n9570), .C2(n7947), .A(n7946), .B(n7945), .ZN(n7948)
         );
  INV_X1 U9648 ( .A(n7948), .ZN(n7949) );
  NOR2_X1 U9649 ( .A1(n10231), .A2(n9841), .ZN(n7952) );
  NAND2_X1 U9650 ( .A1(n10231), .A2(n9841), .ZN(n7951) );
  NAND2_X1 U9651 ( .A1(n9114), .A2(n9677), .ZN(n7954) );
  OR2_X1 U9652 ( .A1(n9680), .A2(n9351), .ZN(n7953) );
  XNOR2_X1 U9653 ( .A(n7967), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9970) );
  NAND2_X1 U9654 ( .A1(n9970), .A2(n7955), .ZN(n7960) );
  INV_X1 U9655 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n9159) );
  NAND2_X1 U9656 ( .A1(n6466), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n7957) );
  NAND2_X1 U9657 ( .A1(n7974), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n7956) );
  OAI211_X1 U9658 ( .C1(n9159), .C2(n9570), .A(n7957), .B(n7956), .ZN(n7958)
         );
  INV_X1 U9659 ( .A(n7958), .ZN(n7959) );
  NAND2_X1 U9660 ( .A1(n10226), .A2(n8138), .ZN(n9726) );
  INV_X1 U9661 ( .A(n10226), .ZN(n9973) );
  NAND2_X1 U9662 ( .A1(n9973), .A2(n8138), .ZN(n7961) );
  NAND2_X1 U9663 ( .A1(n8006), .A2(n9677), .ZN(n7963) );
  OR2_X1 U9664 ( .A1(n9680), .A2(n8007), .ZN(n7962) );
  INV_X1 U9665 ( .A(n7967), .ZN(n7965) );
  AND2_X1 U9666 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n7964) );
  NAND2_X1 U9667 ( .A1(n7965), .A2(n7964), .ZN(n9948) );
  INV_X1 U9668 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9398) );
  INV_X1 U9669 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n7966) );
  INV_X1 U9670 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n7997) );
  NAND2_X1 U9671 ( .A1(n7974), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n7969) );
  NAND2_X1 U9672 ( .A1(n6466), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n7968) );
  OAI211_X1 U9673 ( .C1(n9570), .C2(n7997), .A(n7969), .B(n7968), .ZN(n7970)
         );
  NAND2_X1 U9674 ( .A1(n9943), .A2(n9966), .ZN(n9951) );
  INV_X1 U9675 ( .A(n9576), .ZN(n7971) );
  OR2_X1 U9676 ( .A1(n9948), .A2(n6593), .ZN(n7980) );
  INV_X1 U9677 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n7977) );
  NAND2_X1 U9678 ( .A1(n7974), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n7976) );
  NAND2_X1 U9679 ( .A1(n6466), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n7975) );
  OAI211_X1 U9680 ( .C1(n9570), .C2(n7977), .A(n7976), .B(n7975), .ZN(n7978)
         );
  INV_X1 U9681 ( .A(n7978), .ZN(n7979) );
  INV_X1 U9682 ( .A(n10208), .ZN(n10211) );
  INV_X1 U9683 ( .A(n9623), .ZN(n7983) );
  NAND2_X1 U9684 ( .A1(n7981), .A2(n9625), .ZN(n7982) );
  NAND2_X1 U9685 ( .A1(n7982), .A2(n9623), .ZN(n9749) );
  OR2_X1 U9686 ( .A1(n10295), .A2(n10166), .ZN(n9627) );
  NAND2_X1 U9687 ( .A1(n10295), .A2(n10166), .ZN(n9753) );
  NAND2_X1 U9688 ( .A1(n9627), .A2(n9753), .ZN(n10184) );
  XNOR2_X1 U9689 ( .A(n10292), .B(n10138), .ZN(n10162) );
  NOR2_X1 U9690 ( .A1(n10285), .A2(n10168), .ZN(n9581) );
  NAND2_X1 U9691 ( .A1(n10285), .A2(n10168), .ZN(n9737) );
  INV_X1 U9692 ( .A(n10131), .ZN(n9715) );
  AND2_X1 U9693 ( .A1(n10275), .A2(n10134), .ZN(n9638) );
  OR2_X1 U9694 ( .A1(n10275), .A2(n10134), .ZN(n10098) );
  AND2_X1 U9695 ( .A1(n9643), .A2(n10098), .ZN(n9761) );
  INV_X1 U9696 ( .A(n10103), .ZN(n9530) );
  OR2_X1 U9697 ( .A1(n10265), .A2(n9530), .ZN(n9657) );
  NAND2_X1 U9698 ( .A1(n10265), .A2(n9530), .ZN(n9766) );
  OR2_X1 U9699 ( .A1(n10260), .A2(n10054), .ZN(n9692) );
  AND2_X1 U9700 ( .A1(n10260), .A2(n10054), .ZN(n9653) );
  NOR2_X1 U9701 ( .A1(n10047), .A2(n9653), .ZN(n7988) );
  NAND2_X1 U9702 ( .A1(n10051), .A2(n7988), .ZN(n10036) );
  NAND2_X1 U9703 ( .A1(n5048), .A2(n10055), .ZN(n10021) );
  NAND2_X1 U9704 ( .A1(n9746), .A2(n10021), .ZN(n10037) );
  INV_X1 U9705 ( .A(n9768), .ZN(n10038) );
  NOR2_X1 U9706 ( .A1(n10037), .A2(n10038), .ZN(n7989) );
  INV_X1 U9707 ( .A(n10041), .ZN(n10012) );
  NAND2_X1 U9708 ( .A1(n10248), .A2(n10012), .ZN(n9773) );
  NAND2_X1 U9709 ( .A1(n9747), .A2(n9773), .ZN(n10022) );
  INV_X1 U9710 ( .A(n10021), .ZN(n7990) );
  NOR2_X1 U9711 ( .A1(n10022), .A2(n7990), .ZN(n7991) );
  NAND2_X1 U9712 ( .A1(n10039), .A2(n7991), .ZN(n7992) );
  XNOR2_X1 U9713 ( .A(n10243), .B(n9842), .ZN(n10009) );
  OR2_X1 U9714 ( .A1(n10231), .A2(n9997), .ZN(n9651) );
  NAND2_X1 U9715 ( .A1(n10231), .A2(n9997), .ZN(n9727) );
  NAND2_X1 U9716 ( .A1(n9968), .A2(n9781), .ZN(n7996) );
  INV_X1 U9717 ( .A(n9781), .ZN(n9728) );
  NOR2_X1 U9718 ( .A1(n9576), .A2(n9728), .ZN(n7995) );
  NAND2_X1 U9719 ( .A1(n10155), .A2(n10149), .ZN(n10123) );
  INV_X1 U9720 ( .A(n10270), .ZN(n10097) );
  NAND2_X1 U9721 ( .A1(n10108), .A2(n10097), .ZN(n10080) );
  OAI21_X1 U9722 ( .B1(n4458), .B2(n10221), .A(n9945), .ZN(n10222) );
  OAI22_X1 U9723 ( .A1(n8139), .A2(n10157), .B1(n7997), .B2(n10170), .ZN(n7998) );
  AOI21_X1 U9724 ( .B1(n9943), .B2(n10048), .A(n7998), .ZN(n7999) );
  OAI21_X1 U9725 ( .B1(n10222), .B2(n8000), .A(n7999), .ZN(n8001) );
  AOI21_X1 U9726 ( .B1(n10224), .B2(n10170), .A(n8001), .ZN(n8002) );
  OAI21_X1 U9727 ( .B1(n10225), .B2(n10197), .A(n8002), .ZN(P1_U3263) );
  OAI222_X1 U9728 ( .A1(n8008), .A2(n8005), .B1(n8004), .B2(n8003), .C1(n10059), .C2(P1_U3084), .ZN(P1_U3334) );
  INV_X1 U9729 ( .A(n8006), .ZN(n9113) );
  OAI222_X1 U9730 ( .A1(n8008), .A2(n8007), .B1(P1_U3084), .B2(n6197), .C1(
        n8004), .C2(n9113), .ZN(P1_U3325) );
  INV_X1 U9731 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9564) );
  NAND2_X1 U9732 ( .A1(n8011), .A2(n9317), .ZN(n8010) );
  MUX2_X1 U9733 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n4397), .Z(n8301) );
  XNOR2_X1 U9734 ( .A(n8301), .B(SI_30_), .ZN(n8012) );
  INV_X1 U9735 ( .A(n9563), .ZN(n9108) );
  OAI222_X1 U9736 ( .A1(n8008), .A2(n9564), .B1(n8004), .B2(n9108), .C1(n4749), 
        .C2(P1_U3084), .ZN(P1_U3323) );
  NAND2_X1 U9737 ( .A1(n9943), .A2(n8126), .ZN(n8015) );
  NAND2_X1 U9738 ( .A1(n9956), .A2(n8133), .ZN(n8014) );
  NAND2_X1 U9739 ( .A1(n8015), .A2(n8014), .ZN(n8016) );
  XNOR2_X1 U9740 ( .A(n8016), .B(n8130), .ZN(n8018) );
  AOI22_X1 U9741 ( .A1(n9943), .A2(n8133), .B1(n8084), .B2(n9956), .ZN(n8017)
         );
  XNOR2_X1 U9742 ( .A(n8018), .B(n8017), .ZN(n8144) );
  INV_X1 U9743 ( .A(n8144), .ZN(n8019) );
  NAND2_X1 U9744 ( .A1(n8019), .A2(n9507), .ZN(n8150) );
  NAND2_X1 U9745 ( .A1(n10282), .A2(n8133), .ZN(n8021) );
  NAND2_X1 U9746 ( .A1(n8084), .A2(n10115), .ZN(n8020) );
  NAND2_X1 U9747 ( .A1(n8021), .A2(n8020), .ZN(n8048) );
  INV_X1 U9748 ( .A(n8048), .ZN(n8046) );
  NAND2_X1 U9749 ( .A1(n10285), .A2(n8133), .ZN(n8023) );
  OR2_X1 U9750 ( .A1(n10168), .A2(n8123), .ZN(n8022) );
  NAND2_X1 U9751 ( .A1(n8023), .A2(n8022), .ZN(n9467) );
  INV_X1 U9752 ( .A(n9467), .ZN(n9548) );
  OAI22_X1 U9753 ( .A1(n10156), .A2(n8121), .B1(n10138), .B2(n8127), .ZN(n8024) );
  XNOR2_X1 U9754 ( .A(n8024), .B(n8130), .ZN(n9404) );
  INV_X1 U9755 ( .A(n9404), .ZN(n8038) );
  NAND2_X1 U9756 ( .A1(n10303), .A2(n8126), .ZN(n8028) );
  OR2_X1 U9757 ( .A1(n8030), .A2(n8127), .ZN(n8027) );
  NAND2_X1 U9758 ( .A1(n8028), .A2(n8027), .ZN(n8029) );
  XNOR2_X1 U9759 ( .A(n8029), .B(n8096), .ZN(n8033) );
  NOR2_X1 U9760 ( .A1(n8123), .A2(n8030), .ZN(n8031) );
  AOI21_X1 U9761 ( .B1(n10303), .B2(n8133), .A(n8031), .ZN(n8032) );
  OR2_X1 U9762 ( .A1(n8033), .A2(n8032), .ZN(n9447) );
  OAI22_X1 U9763 ( .A1(n10183), .A2(n8121), .B1(n10166), .B2(n8127), .ZN(n8034) );
  OAI22_X1 U9764 ( .A1(n10183), .A2(n8127), .B1(n10166), .B2(n8123), .ZN(n9504) );
  AOI22_X1 U9765 ( .A1(n10292), .A2(n8133), .B1(n8084), .B2(n10190), .ZN(n8036) );
  INV_X1 U9766 ( .A(n8036), .ZN(n9405) );
  NAND2_X1 U9767 ( .A1(n8035), .A2(n9405), .ZN(n9462) );
  INV_X1 U9768 ( .A(n8047), .ZN(n8037) );
  NAND2_X1 U9769 ( .A1(n10282), .A2(n8126), .ZN(n8040) );
  NAND2_X1 U9770 ( .A1(n10115), .A2(n8133), .ZN(n8039) );
  NAND2_X1 U9771 ( .A1(n8040), .A2(n8039), .ZN(n8041) );
  XNOR2_X1 U9772 ( .A(n8041), .B(n8130), .ZN(n8049) );
  INV_X1 U9773 ( .A(n8049), .ZN(n8042) );
  NAND2_X1 U9774 ( .A1(n8042), .A2(n8046), .ZN(n9478) );
  OAI22_X1 U9775 ( .A1(n10149), .A2(n8121), .B1(n10168), .B2(n8127), .ZN(n8043) );
  XOR2_X1 U9776 ( .A(n6504), .B(n8043), .Z(n9463) );
  INV_X1 U9777 ( .A(n9463), .ZN(n9465) );
  NAND3_X1 U9778 ( .A1(n9466), .A2(n9478), .A3(n9465), .ZN(n8045) );
  OAI21_X1 U9779 ( .B1(n8048), .B2(n9467), .A(n8049), .ZN(n8044) );
  NAND2_X1 U9780 ( .A1(n8047), .A2(n9404), .ZN(n9464) );
  NAND2_X1 U9781 ( .A1(n8049), .A2(n8048), .ZN(n9470) );
  NAND4_X1 U9782 ( .A1(n9464), .A2(n9463), .A3(n9462), .A4(n9470), .ZN(n8053)
         );
  NAND2_X1 U9783 ( .A1(n10275), .A2(n8126), .ZN(n8051) );
  NAND2_X1 U9784 ( .A1(n10102), .A2(n8133), .ZN(n8050) );
  NAND2_X1 U9785 ( .A1(n8051), .A2(n8050), .ZN(n8052) );
  XNOR2_X1 U9786 ( .A(n8052), .B(n6504), .ZN(n8055) );
  OAI22_X1 U9787 ( .A1(n10112), .A2(n8127), .B1(n10134), .B2(n8123), .ZN(n8054) );
  XNOR2_X1 U9788 ( .A(n8055), .B(n8054), .ZN(n9477) );
  NAND2_X1 U9789 ( .A1(n10265), .A2(n8126), .ZN(n8058) );
  NAND2_X1 U9790 ( .A1(n10103), .A2(n8133), .ZN(n8057) );
  NAND2_X1 U9791 ( .A1(n8058), .A2(n8057), .ZN(n8059) );
  XNOR2_X1 U9792 ( .A(n8059), .B(n8130), .ZN(n9430) );
  AOI22_X1 U9793 ( .A1(n10265), .A2(n8133), .B1(n8084), .B2(n10103), .ZN(n8065) );
  INV_X1 U9794 ( .A(n8065), .ZN(n9429) );
  NOR2_X1 U9795 ( .A1(n9482), .A2(n8123), .ZN(n8060) );
  AOI21_X1 U9796 ( .B1(n10270), .B2(n8133), .A(n8060), .ZN(n9526) );
  INV_X1 U9797 ( .A(n9526), .ZN(n8064) );
  NAND2_X1 U9798 ( .A1(n10270), .A2(n8126), .ZN(n8062) );
  OR2_X1 U9799 ( .A1(n9482), .A2(n8127), .ZN(n8061) );
  NAND2_X1 U9800 ( .A1(n8062), .A2(n8061), .ZN(n8063) );
  XNOR2_X1 U9801 ( .A(n8063), .B(n8096), .ZN(n9527) );
  INV_X1 U9802 ( .A(n9527), .ZN(n9428) );
  AOI22_X1 U9803 ( .A1(n9430), .A2(n9429), .B1(n8064), .B2(n9428), .ZN(n8069)
         );
  AOI21_X1 U9804 ( .B1(n9527), .B2(n9526), .A(n8065), .ZN(n8067) );
  NAND2_X1 U9805 ( .A1(n8065), .A2(n9526), .ZN(n8066) );
  OAI22_X1 U9806 ( .A1(n8067), .A2(n9430), .B1(n9428), .B2(n8066), .ZN(n8068)
         );
  NAND2_X1 U9807 ( .A1(n10260), .A2(n8126), .ZN(n8071) );
  NAND2_X1 U9808 ( .A1(n10086), .A2(n8133), .ZN(n8070) );
  NAND2_X1 U9809 ( .A1(n8071), .A2(n8070), .ZN(n8072) );
  XNOR2_X1 U9810 ( .A(n8072), .B(n8130), .ZN(n8074) );
  OAI22_X1 U9811 ( .A1(n10071), .A2(n8127), .B1(n10054), .B2(n8123), .ZN(n8073) );
  XNOR2_X1 U9812 ( .A(n8074), .B(n8073), .ZN(n9497) );
  NAND2_X1 U9813 ( .A1(n10256), .A2(n8126), .ZN(n8076) );
  NAND2_X1 U9814 ( .A1(n10074), .A2(n8133), .ZN(n8075) );
  NAND2_X1 U9815 ( .A1(n8076), .A2(n8075), .ZN(n8077) );
  XNOR2_X1 U9816 ( .A(n8077), .B(n8130), .ZN(n8078) );
  AOI22_X1 U9817 ( .A1(n10256), .A2(n8133), .B1(n8084), .B2(n10074), .ZN(n8079) );
  XNOR2_X1 U9818 ( .A(n8078), .B(n8079), .ZN(n9440) );
  INV_X1 U9819 ( .A(n8078), .ZN(n8080) );
  NAND2_X1 U9820 ( .A1(n8080), .A2(n8079), .ZN(n8081) );
  AND2_X1 U9821 ( .A1(n10041), .A2(n8133), .ZN(n8083) );
  AOI21_X1 U9822 ( .B1(n10248), .B2(n8126), .A(n8083), .ZN(n8098) );
  XNOR2_X1 U9823 ( .A(n8098), .B(n6504), .ZN(n9417) );
  AND2_X1 U9824 ( .A1(n10041), .A2(n8084), .ZN(n8085) );
  AOI21_X1 U9825 ( .B1(n10248), .B2(n8133), .A(n8085), .ZN(n9416) );
  NOR2_X1 U9826 ( .A1(n9417), .A2(n9416), .ZN(n8090) );
  OR2_X1 U9827 ( .A1(n10035), .A2(n8121), .ZN(n8087) );
  OR2_X1 U9828 ( .A1(n10055), .A2(n8127), .ZN(n8086) );
  XNOR2_X1 U9829 ( .A(n8095), .B(n8096), .ZN(n9517) );
  OR2_X1 U9830 ( .A1(n10035), .A2(n8127), .ZN(n8089) );
  OR2_X1 U9831 ( .A1(n10055), .A2(n8123), .ZN(n8088) );
  INV_X1 U9832 ( .A(n9417), .ZN(n8092) );
  OAI21_X1 U9833 ( .B1(n9517), .B2(n9414), .A(n8092), .ZN(n8102) );
  OR2_X1 U9834 ( .A1(n8095), .A2(n6504), .ZN(n8094) );
  INV_X1 U9835 ( .A(n8098), .ZN(n8093) );
  OAI21_X1 U9836 ( .B1(n8094), .B2(n9414), .A(n8093), .ZN(n8101) );
  INV_X1 U9837 ( .A(n8095), .ZN(n8097) );
  OR2_X1 U9838 ( .A1(n8097), .A2(n8096), .ZN(n8099) );
  OAI21_X1 U9839 ( .B1(n8099), .B2(n9414), .A(n8098), .ZN(n8100) );
  AOI22_X1 U9840 ( .A1(n8102), .A2(n9416), .B1(n8101), .B2(n8100), .ZN(n9487)
         );
  OAI22_X1 U9841 ( .A1(n9577), .A2(n8121), .B1(n10025), .B2(n8127), .ZN(n8103)
         );
  XNOR2_X1 U9842 ( .A(n8103), .B(n8130), .ZN(n8107) );
  INV_X1 U9843 ( .A(n8107), .ZN(n8105) );
  OAI22_X1 U9844 ( .A1(n9577), .A2(n8127), .B1(n10025), .B2(n8123), .ZN(n8108)
         );
  INV_X1 U9845 ( .A(n8108), .ZN(n8104) );
  NAND2_X1 U9846 ( .A1(n8105), .A2(n8104), .ZN(n8106) );
  AND2_X1 U9847 ( .A1(n9487), .A2(n8106), .ZN(n8110) );
  INV_X1 U9848 ( .A(n8106), .ZN(n8109) );
  XOR2_X1 U9849 ( .A(n8108), .B(n8107), .Z(n9490) );
  OAI22_X1 U9850 ( .A1(n8111), .A2(n8127), .B1(n10013), .B2(n8123), .ZN(n8116)
         );
  NAND2_X1 U9851 ( .A1(n10238), .A2(n8126), .ZN(n8113) );
  NAND2_X1 U9852 ( .A1(n9989), .A2(n8133), .ZN(n8112) );
  NAND2_X1 U9853 ( .A1(n8113), .A2(n8112), .ZN(n8114) );
  XNOR2_X1 U9854 ( .A(n8114), .B(n8130), .ZN(n8115) );
  XOR2_X1 U9855 ( .A(n8116), .B(n8115), .Z(n9456) );
  INV_X1 U9856 ( .A(n8115), .ZN(n8118) );
  INV_X1 U9857 ( .A(n8116), .ZN(n8117) );
  NAND2_X1 U9858 ( .A1(n8118), .A2(n8117), .ZN(n8119) );
  OAI22_X1 U9859 ( .A1(n9984), .A2(n8121), .B1(n9997), .B2(n8127), .ZN(n8122)
         );
  XNOR2_X1 U9860 ( .A(n8122), .B(n8130), .ZN(n8125) );
  OAI22_X1 U9861 ( .A1(n9984), .A2(n8127), .B1(n9997), .B2(n8123), .ZN(n8124)
         );
  XNOR2_X1 U9862 ( .A(n8125), .B(n8124), .ZN(n9536) );
  NAND2_X1 U9863 ( .A1(n10226), .A2(n8126), .ZN(n8129) );
  OR2_X1 U9864 ( .A1(n8138), .A2(n8127), .ZN(n8128) );
  NAND2_X1 U9865 ( .A1(n8129), .A2(n8128), .ZN(n8131) );
  XNOR2_X1 U9866 ( .A(n8131), .B(n8130), .ZN(n9394) );
  INV_X1 U9867 ( .A(n9394), .ZN(n8134) );
  NOR2_X1 U9868 ( .A1(n8138), .A2(n8123), .ZN(n8132) );
  AOI21_X1 U9869 ( .B1(n10226), .B2(n8133), .A(n8132), .ZN(n9393) );
  NAND2_X1 U9870 ( .A1(n8134), .A2(n9393), .ZN(n8135) );
  INV_X1 U9871 ( .A(n9393), .ZN(n8136) );
  NAND2_X1 U9872 ( .A1(n9394), .A2(n8136), .ZN(n8143) );
  AND2_X1 U9873 ( .A1(n8144), .A2(n5333), .ZN(n8137) );
  NAND2_X1 U9874 ( .A1(n8149), .A2(n8137), .ZN(n8148) );
  NAND2_X1 U9875 ( .A1(n9990), .A2(n9511), .ZN(n8142) );
  INV_X1 U9876 ( .A(n8139), .ZN(n8140) );
  AOI22_X1 U9877 ( .A1(n8140), .A2(n9550), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n8141) );
  OAI211_X1 U9878 ( .C1(n10211), .C2(n9529), .A(n8142), .B(n8141), .ZN(n8146)
         );
  NOR3_X1 U9879 ( .A1(n8144), .A2(n9558), .A3(n8143), .ZN(n8145) );
  AOI211_X1 U9880 ( .C1(n9943), .C2(n9556), .A(n8146), .B(n8145), .ZN(n8147)
         );
  OAI211_X1 U9881 ( .C1(n8150), .C2(n8149), .A(n8148), .B(n8147), .ZN(P1_U3218) );
  INV_X1 U9882 ( .A(n8151), .ZN(n8152) );
  AOI21_X1 U9883 ( .B1(n8154), .B2(n8153), .A(n8152), .ZN(n8161) );
  OAI21_X1 U9884 ( .B1(n8277), .B2(n8925), .A(n8155), .ZN(n8159) );
  OAI22_X1 U9885 ( .A1(n8254), .A2(n8157), .B1(n8156), .B2(n8263), .ZN(n8158)
         );
  AOI211_X1 U9886 ( .C1(n8280), .C2(n9054), .A(n8159), .B(n8158), .ZN(n8160)
         );
  OAI21_X1 U9887 ( .B1(n8161), .B2(n8282), .A(n8160), .ZN(P2_U3217) );
  NOR2_X1 U9888 ( .A1(n8163), .A2(n8219), .ZN(n8165) );
  XNOR2_X1 U9889 ( .A(n8165), .B(n8164), .ZN(n8170) );
  OAI22_X1 U9890 ( .A1(n8192), .A2(n8277), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8166), .ZN(n8168) );
  OAI22_X1 U9891 ( .A1(n8254), .A2(n8807), .B1(n8453), .B2(n8263), .ZN(n8167)
         );
  AOI211_X1 U9892 ( .C1(n9005), .C2(n8280), .A(n8168), .B(n8167), .ZN(n8169)
         );
  OAI21_X1 U9893 ( .B1(n8170), .B2(n8282), .A(n8169), .ZN(P2_U3218) );
  INV_X1 U9894 ( .A(n8172), .ZN(n8173) );
  AOI21_X1 U9895 ( .B1(n8171), .B2(n8174), .A(n8173), .ZN(n8178) );
  AND2_X1 U9896 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8684) );
  OAI22_X1 U9897 ( .A1(n8254), .A2(n8870), .B1(n8214), .B2(n8263), .ZN(n8175)
         );
  AOI211_X1 U9898 ( .C1(n8209), .C2(n8866), .A(n8684), .B(n8175), .ZN(n8177)
         );
  NAND2_X1 U9899 ( .A1(n9028), .A2(n8280), .ZN(n8176) );
  OAI211_X1 U9900 ( .C1(n8178), .C2(n8282), .A(n8177), .B(n8176), .ZN(P2_U3221) );
  XNOR2_X1 U9901 ( .A(n8180), .B(n8179), .ZN(n8187) );
  OAI22_X1 U9902 ( .A1(n8277), .A2(n8453), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8181), .ZN(n8185) );
  INV_X1 U9903 ( .A(n8834), .ZN(n8183) );
  OAI22_X1 U9904 ( .A1(n8254), .A2(n8183), .B1(n8182), .B2(n8263), .ZN(n8184)
         );
  AOI211_X1 U9905 ( .C1(n9015), .C2(n8280), .A(n8185), .B(n8184), .ZN(n8186)
         );
  OAI21_X1 U9906 ( .B1(n8187), .B2(n8282), .A(n8186), .ZN(P2_U3225) );
  XNOR2_X1 U9907 ( .A(n8189), .B(n8188), .ZN(n8190) );
  XNOR2_X1 U9908 ( .A(n8191), .B(n8190), .ZN(n8198) );
  INV_X1 U9909 ( .A(n8762), .ZN(n8195) );
  OAI22_X1 U9910 ( .A1(n8193), .A2(n8926), .B1(n8192), .B2(n8924), .ZN(n8767)
         );
  AOI22_X1 U9911 ( .A1(n8767), .A2(n8227), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8194) );
  OAI21_X1 U9912 ( .B1(n8195), .B2(n8254), .A(n8194), .ZN(n8196) );
  AOI21_X1 U9913 ( .B1(n8996), .B2(n8280), .A(n8196), .ZN(n8197) );
  OAI21_X1 U9914 ( .B1(n8198), .B2(n8282), .A(n8197), .ZN(P2_U3227) );
  INV_X1 U9915 ( .A(n8942), .ZN(n9041) );
  NAND2_X1 U9916 ( .A1(n8200), .A2(n8199), .ZN(n8201) );
  OAI21_X1 U9917 ( .B1(n8200), .B2(n8199), .A(n8201), .ZN(n8270) );
  NOR2_X1 U9918 ( .A1(n8270), .A2(n8271), .ZN(n8269) );
  INV_X1 U9919 ( .A(n8201), .ZN(n8203) );
  NOR3_X1 U9920 ( .A1(n8269), .A2(n8203), .A3(n8202), .ZN(n8206) );
  INV_X1 U9921 ( .A(n8204), .ZN(n8205) );
  OAI21_X1 U9922 ( .B1(n8206), .B2(n8205), .A(n7733), .ZN(n8211) );
  OAI22_X1 U9923 ( .A1(n8254), .A2(n8938), .B1(n8925), .B2(n8263), .ZN(n8207)
         );
  AOI211_X1 U9924 ( .C1(n8209), .C2(n8887), .A(n8208), .B(n8207), .ZN(n8210)
         );
  OAI211_X1 U9925 ( .C1(n9041), .C2(n8268), .A(n8211), .B(n8210), .ZN(P2_U3228) );
  XNOR2_X1 U9926 ( .A(n8213), .B(n8212), .ZN(n8218) );
  OAI22_X1 U9927 ( .A1(n8214), .A2(n8926), .B1(n8278), .B2(n8924), .ZN(n8908)
         );
  AOI22_X1 U9928 ( .A1(n8227), .A2(n8908), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3152), .ZN(n8215) );
  OAI21_X1 U9929 ( .B1(n8254), .B2(n8916), .A(n8215), .ZN(n8216) );
  AOI21_X1 U9930 ( .B1(n9037), .B2(n8280), .A(n8216), .ZN(n8217) );
  OAI21_X1 U9931 ( .B1(n8218), .B2(n8282), .A(n8217), .ZN(P2_U3230) );
  NOR2_X1 U9932 ( .A1(n8220), .A2(n8219), .ZN(n8224) );
  XNOR2_X1 U9933 ( .A(n8222), .B(n8221), .ZN(n8223) );
  XNOR2_X1 U9934 ( .A(n8224), .B(n8223), .ZN(n8231) );
  OR2_X1 U9935 ( .A1(n8741), .A2(n8926), .ZN(n8226) );
  NAND2_X1 U9936 ( .A1(n8512), .A2(n8886), .ZN(n8225) );
  NAND2_X1 U9937 ( .A1(n8226), .A2(n8225), .ZN(n8785) );
  AOI22_X1 U9938 ( .A1(n8785), .A2(n8227), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3152), .ZN(n8228) );
  OAI21_X1 U9939 ( .B1(n8779), .B2(n8254), .A(n8228), .ZN(n8229) );
  AOI21_X1 U9940 ( .B1(n9000), .B2(n8280), .A(n8229), .ZN(n8230) );
  OAI21_X1 U9941 ( .B1(n8231), .B2(n8282), .A(n8230), .ZN(P2_U3231) );
  XNOR2_X1 U9942 ( .A(n8233), .B(n8232), .ZN(n8239) );
  OAI22_X1 U9943 ( .A1(n8277), .A2(n8850), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8234), .ZN(n8237) );
  INV_X1 U9944 ( .A(n8853), .ZN(n8235) );
  OAI22_X1 U9945 ( .A1(n8254), .A2(n8235), .B1(n8848), .B2(n8263), .ZN(n8236)
         );
  AOI211_X1 U9946 ( .C1(n9022), .C2(n8280), .A(n8237), .B(n8236), .ZN(n8238)
         );
  OAI21_X1 U9947 ( .B1(n8239), .B2(n8282), .A(n8238), .ZN(P2_U3235) );
  INV_X1 U9948 ( .A(n8240), .ZN(n8241) );
  NOR2_X1 U9949 ( .A1(n4486), .A2(n8241), .ZN(n8245) );
  XNOR2_X1 U9950 ( .A(n8243), .B(n8242), .ZN(n8244) );
  XNOR2_X1 U9951 ( .A(n8245), .B(n8244), .ZN(n8249) );
  OAI22_X1 U9952 ( .A1(n8277), .A2(n8824), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9325), .ZN(n8247) );
  OAI22_X1 U9953 ( .A1(n8254), .A2(n8817), .B1(n8850), .B2(n8263), .ZN(n8246)
         );
  AOI211_X1 U9954 ( .C1(n9010), .C2(n8280), .A(n8247), .B(n8246), .ZN(n8248)
         );
  OAI21_X1 U9955 ( .B1(n8249), .B2(n8282), .A(n8248), .ZN(P2_U3237) );
  XNOR2_X1 U9956 ( .A(n8251), .B(n8250), .ZN(n8258) );
  OAI21_X1 U9957 ( .B1(n8277), .B2(n8848), .A(n8252), .ZN(n8256) );
  INV_X1 U9958 ( .A(n8253), .ZN(n8891) );
  OAI22_X1 U9959 ( .A1(n8254), .A2(n8891), .B1(n8927), .B2(n8263), .ZN(n8255)
         );
  AOI211_X1 U9960 ( .C1(n9032), .C2(n8280), .A(n8256), .B(n8255), .ZN(n8257)
         );
  OAI21_X1 U9961 ( .B1(n8258), .B2(n8282), .A(n8257), .ZN(P2_U3240) );
  OAI211_X1 U9962 ( .C1(n8261), .C2(n8260), .A(n8259), .B(n7733), .ZN(n8267)
         );
  INV_X1 U9963 ( .A(n8262), .ZN(n8750) );
  OAI22_X1 U9964 ( .A1(n8741), .A2(n8263), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9254), .ZN(n8265) );
  NOR2_X1 U9965 ( .A1(n8742), .A2(n8277), .ZN(n8264) );
  AOI211_X1 U9966 ( .C1(n8273), .C2(n8750), .A(n8265), .B(n8264), .ZN(n8266)
         );
  OAI211_X1 U9967 ( .C1(n5269), .C2(n8268), .A(n8267), .B(n8266), .ZN(P2_U3242) );
  AOI21_X1 U9968 ( .B1(n8271), .B2(n8270), .A(n8269), .ZN(n8283) );
  AOI22_X1 U9969 ( .A1(n8274), .A2(n8517), .B1(n8273), .B2(n8272), .ZN(n8276)
         );
  OAI211_X1 U9970 ( .C1(n8278), .C2(n8277), .A(n8276), .B(n8275), .ZN(n8279)
         );
  AOI21_X1 U9971 ( .B1(n8280), .B2(n9049), .A(n8279), .ZN(n8281) );
  OAI21_X1 U9972 ( .B1(n8283), .B2(n8282), .A(n8281), .ZN(P2_U3243) );
  NAND2_X1 U9973 ( .A1(n9678), .A2(n8307), .ZN(n8286) );
  NAND2_X1 U9974 ( .A1(n8308), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8285) );
  NAND2_X1 U9975 ( .A1(n8971), .A2(n8508), .ZN(n8482) );
  INV_X1 U9976 ( .A(n8482), .ZN(n8287) );
  OR2_X1 U9977 ( .A1(n8311), .A2(n8337), .ZN(n8294) );
  INV_X1 U9978 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9281) );
  NAND2_X1 U9979 ( .A1(n8288), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8290) );
  NAND2_X1 U9980 ( .A1(n6182), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8289) );
  OAI211_X1 U9981 ( .C1(n5641), .C2(n9281), .A(n8290), .B(n8289), .ZN(n8507)
         );
  NAND2_X1 U9982 ( .A1(n9563), .A2(n8307), .ZN(n8292) );
  NAND2_X1 U9983 ( .A1(n8308), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8291) );
  NAND2_X1 U9984 ( .A1(n8295), .A2(n8294), .ZN(n8296) );
  NAND2_X1 U9985 ( .A1(n8297), .A2(n8296), .ZN(n8313) );
  NAND2_X1 U9986 ( .A1(n8301), .A2(SI_30_), .ZN(n8298) );
  INV_X1 U9987 ( .A(n8301), .ZN(n8303) );
  INV_X1 U9988 ( .A(SI_30_), .ZN(n8302) );
  NAND2_X1 U9989 ( .A1(n8303), .A2(n8302), .ZN(n8304) );
  MUX2_X1 U9990 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n4394), .Z(n8305) );
  XNOR2_X1 U9991 ( .A(n8305), .B(n9309), .ZN(n8306) );
  NAND2_X1 U9992 ( .A1(n9560), .A2(n8307), .ZN(n8310) );
  NAND2_X1 U9993 ( .A1(n8308), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8309) );
  INV_X1 U9994 ( .A(n8311), .ZN(n8689) );
  INV_X1 U9995 ( .A(n8507), .ZN(n8709) );
  NAND2_X1 U9996 ( .A1(n8694), .A2(n8709), .ZN(n8312) );
  NAND2_X1 U9997 ( .A1(n5575), .A2(n8314), .ZN(n8501) );
  OR2_X1 U9998 ( .A1(n8694), .A2(n8709), .ZN(n8487) );
  INV_X1 U9999 ( .A(n8823), .ZN(n8443) );
  INV_X1 U10000 ( .A(n8864), .ZN(n8875) );
  NOR3_X1 U10001 ( .A1(n7026), .A2(n7030), .A3(n6025), .ZN(n8319) );
  NAND2_X1 U10002 ( .A1(n8316), .A2(n6099), .ZN(n8317) );
  AND2_X1 U10003 ( .A1(n8347), .A2(n8317), .ZN(n8342) );
  NAND4_X1 U10004 ( .A1(n8319), .A2(n8342), .A3(n8318), .A4(n4675), .ZN(n8322)
         );
  INV_X1 U10005 ( .A(n8369), .ZN(n8343) );
  NOR4_X1 U10006 ( .A1(n8322), .A2(n8321), .A3(n8343), .A4(n8320), .ZN(n8326)
         );
  NAND4_X1 U10007 ( .A1(n8326), .A2(n8325), .A3(n8324), .A4(n8323), .ZN(n8329)
         );
  NAND4_X1 U10008 ( .A1(n8928), .A2(n8420), .A3(n8330), .A4(n8406), .ZN(n8331)
         );
  NAND4_X1 U10009 ( .A1(n8792), .A2(n5223), .A3(n8839), .A4(n8332), .ZN(n8333)
         );
  NOR4_X1 U10010 ( .A1(n8765), .A2(n4587), .A3(n8803), .A4(n8333), .ZN(n8334)
         );
  INV_X1 U10011 ( .A(n8717), .ZN(n8725) );
  NAND4_X1 U10012 ( .A1(n8476), .A2(n7789), .A3(n8334), .A4(n8725), .ZN(n8335)
         );
  XNOR2_X1 U10013 ( .A(n8336), .B(n8915), .ZN(n8338) );
  NAND2_X1 U10014 ( .A1(n8338), .A2(n8337), .ZN(n8500) );
  OR2_X1 U10015 ( .A1(n8459), .A2(n8481), .ZN(n8436) );
  MUX2_X1 U10016 ( .A(n8421), .B(n5331), .S(n8494), .Z(n8341) );
  AND2_X1 U10017 ( .A1(n8903), .A2(n8341), .ZN(n8417) );
  INV_X1 U10018 ( .A(n8342), .ZN(n8345) );
  MUX2_X1 U10019 ( .A(n8343), .B(n8345), .S(n8494), .Z(n8371) );
  NOR2_X1 U10020 ( .A1(n8345), .A2(n5143), .ZN(n8346) );
  AOI21_X1 U10021 ( .B1(n8371), .B2(n8347), .A(n8346), .ZN(n8349) );
  OAI21_X1 U10022 ( .B1(n8349), .B2(n8348), .A(n8481), .ZN(n8359) );
  INV_X1 U10023 ( .A(n8371), .ZN(n8357) );
  AND2_X1 U10024 ( .A1(n8351), .A2(n8350), .ZN(n8360) );
  OAI211_X1 U10025 ( .C1(n8353), .C2(n8360), .A(n8352), .B(n8361), .ZN(n8354)
         );
  NAND3_X1 U10026 ( .A1(n8354), .A2(n8363), .A3(n8481), .ZN(n8355) );
  NAND3_X1 U10027 ( .A1(n8357), .A2(n8356), .A3(n8355), .ZN(n8358) );
  INV_X1 U10028 ( .A(n8360), .ZN(n8365) );
  INV_X1 U10029 ( .A(n8361), .ZN(n8364) );
  OAI211_X1 U10030 ( .C1(n8365), .C2(n8364), .A(n8363), .B(n8362), .ZN(n8366)
         );
  NAND3_X1 U10031 ( .A1(n8366), .A2(n8494), .A3(n8352), .ZN(n8367) );
  AOI22_X1 U10032 ( .A1(n8371), .A2(n8370), .B1(n8369), .B2(n8368), .ZN(n8374)
         );
  INV_X1 U10033 ( .A(n8372), .ZN(n8373) );
  OAI21_X1 U10034 ( .B1(n8374), .B2(n8373), .A(n8494), .ZN(n8378) );
  OAI21_X1 U10035 ( .B1(n8376), .B2(n8481), .A(n8375), .ZN(n8377) );
  INV_X1 U10036 ( .A(n8379), .ZN(n8382) );
  INV_X1 U10037 ( .A(n8380), .ZN(n8381) );
  MUX2_X1 U10038 ( .A(n8382), .B(n8381), .S(n8494), .Z(n8384) );
  MUX2_X1 U10039 ( .A(n8386), .B(n8385), .S(n8481), .Z(n8387) );
  NAND3_X1 U10040 ( .A1(n8388), .A2(n8389), .A3(n8387), .ZN(n8397) );
  INV_X1 U10041 ( .A(n8391), .ZN(n8392) );
  NAND2_X1 U10042 ( .A1(n8393), .A2(n8392), .ZN(n8395) );
  NAND3_X1 U10043 ( .A1(n8395), .A2(n8398), .A3(n8394), .ZN(n8396) );
  NAND2_X1 U10044 ( .A1(n8398), .A2(n8402), .ZN(n8401) );
  NAND2_X1 U10045 ( .A1(n8399), .A2(n8403), .ZN(n8400) );
  MUX2_X1 U10046 ( .A(n8401), .B(n8400), .S(n8481), .Z(n8405) );
  MUX2_X1 U10047 ( .A(n8403), .B(n8402), .S(n8481), .Z(n8404) );
  MUX2_X1 U10048 ( .A(n8518), .B(n8407), .S(n8481), .Z(n8409) );
  NOR2_X1 U10049 ( .A1(n8407), .A2(n8518), .ZN(n8408) );
  NOR2_X1 U10050 ( .A1(n8409), .A2(n8408), .ZN(n8410) );
  NOR2_X1 U10051 ( .A1(n8411), .A2(n8410), .ZN(n8412) );
  AND2_X1 U10052 ( .A1(n8413), .A2(n8494), .ZN(n8414) );
  AND2_X1 U10053 ( .A1(n8516), .A2(n8481), .ZN(n8416) );
  NOR2_X1 U10054 ( .A1(n8516), .A2(n8481), .ZN(n8415) );
  MUX2_X1 U10055 ( .A(n8416), .B(n8415), .S(n9049), .Z(n8418) );
  INV_X1 U10056 ( .A(n8928), .ZN(n8922) );
  OAI21_X1 U10057 ( .B1(n8418), .B2(n8922), .A(n8417), .ZN(n8430) );
  AND4_X1 U10058 ( .A1(n8421), .A2(n8420), .A3(n8419), .A4(n8481), .ZN(n8423)
         );
  NAND3_X1 U10059 ( .A1(n8424), .A2(n8423), .A3(n8422), .ZN(n8429) );
  AND2_X1 U10060 ( .A1(n8887), .A2(n8481), .ZN(n8426) );
  OAI21_X1 U10061 ( .B1(n8887), .B2(n8481), .A(n9037), .ZN(n8425) );
  OAI21_X1 U10062 ( .B1(n8426), .B2(n9037), .A(n8425), .ZN(n8427) );
  AND3_X1 U10063 ( .A1(n8438), .A2(n8431), .A3(n8427), .ZN(n8428) );
  NAND3_X1 U10064 ( .A1(n8439), .A2(n8431), .A3(n8846), .ZN(n8433) );
  INV_X1 U10065 ( .A(n8442), .ZN(n8432) );
  AOI21_X1 U10066 ( .B1(n8433), .B2(n8440), .A(n8432), .ZN(n8435) );
  AOI21_X1 U10067 ( .B1(n8439), .B2(n8438), .A(n8437), .ZN(n8446) );
  NAND2_X1 U10068 ( .A1(n8441), .A2(n8440), .ZN(n8445) );
  INV_X1 U10069 ( .A(n8447), .ZN(n8458) );
  NAND2_X1 U10070 ( .A1(n8513), .A2(n8494), .ZN(n8448) );
  OAI22_X1 U10071 ( .A1(n9015), .A2(n8448), .B1(n8453), .B2(n8481), .ZN(n8450)
         );
  INV_X1 U10072 ( .A(n9015), .ZN(n8836) );
  NOR2_X1 U10073 ( .A1(n8453), .A2(n8448), .ZN(n8449) );
  AOI22_X1 U10074 ( .A1(n8820), .A2(n8450), .B1(n8836), .B2(n8449), .ZN(n8457)
         );
  NOR2_X1 U10075 ( .A1(n8513), .A2(n8494), .ZN(n8451) );
  NAND2_X1 U10076 ( .A1(n9015), .A2(n8451), .ZN(n8452) );
  OAI21_X1 U10077 ( .B1(n8494), .B2(n8841), .A(n8452), .ZN(n8455) );
  INV_X1 U10078 ( .A(n8452), .ZN(n8454) );
  AOI22_X1 U10079 ( .A1(n8455), .A2(n9010), .B1(n8454), .B2(n8453), .ZN(n8456)
         );
  OAI21_X1 U10080 ( .B1(n8458), .B2(n8457), .A(n8456), .ZN(n8460) );
  NAND2_X1 U10081 ( .A1(n8460), .A2(n8459), .ZN(n8461) );
  NAND3_X1 U10082 ( .A1(n8467), .A2(n8462), .A3(n8465), .ZN(n8464) );
  NAND2_X1 U10083 ( .A1(n8469), .A2(n8468), .ZN(n8471) );
  OAI21_X1 U10084 ( .B1(n8472), .B2(n8481), .A(n8725), .ZN(n8477) );
  NAND2_X1 U10085 ( .A1(n8510), .A2(n8494), .ZN(n8474) );
  OR2_X1 U10086 ( .A1(n8510), .A2(n8494), .ZN(n8473) );
  MUX2_X1 U10087 ( .A(n8474), .B(n8473), .S(n8984), .Z(n8475) );
  MUX2_X1 U10088 ( .A(n8479), .B(n8478), .S(n8494), .Z(n8480) );
  MUX2_X1 U10089 ( .A(n8483), .B(n8482), .S(n8481), .Z(n8484) );
  AOI22_X1 U10090 ( .A1(n8489), .A2(n8488), .B1(n8486), .B2(n8485), .ZN(n8496)
         );
  INV_X1 U10091 ( .A(n8487), .ZN(n8491) );
  OAI21_X1 U10092 ( .B1(n8491), .B2(n8490), .A(n8489), .ZN(n8493) );
  NAND2_X1 U10093 ( .A1(n8493), .A2(n8492), .ZN(n8495) );
  OAI21_X1 U10094 ( .B1(n8497), .B2(n4741), .A(n10530), .ZN(n8498) );
  INV_X1 U10095 ( .A(n8687), .ZN(n9115) );
  NAND3_X1 U10096 ( .A1(n8502), .A2(n9115), .A3(n8886), .ZN(n8503) );
  OAI211_X1 U10097 ( .C1(n8504), .C2(n8506), .A(n8503), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8505) );
  MUX2_X1 U10098 ( .A(n8507), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8514), .Z(
        P2_U3582) );
  INV_X1 U10099 ( .A(n8508), .ZN(n8509) );
  MUX2_X1 U10100 ( .A(n8509), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8514), .Z(
        P2_U3581) );
  INV_X1 U10101 ( .A(n8710), .ZN(n8728) );
  MUX2_X1 U10102 ( .A(n8728), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8514), .Z(
        P2_U3580) );
  MUX2_X1 U10103 ( .A(n8510), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8514), .Z(
        P2_U3579) );
  MUX2_X1 U10104 ( .A(n8727), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8514), .Z(
        P2_U3578) );
  MUX2_X1 U10105 ( .A(n8511), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8514), .Z(
        P2_U3577) );
  MUX2_X1 U10106 ( .A(n8799), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8514), .Z(
        P2_U3576) );
  MUX2_X1 U10107 ( .A(n8512), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8514), .Z(
        P2_U3575) );
  MUX2_X1 U10108 ( .A(n8841), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8514), .Z(
        P2_U3574) );
  MUX2_X1 U10109 ( .A(n8513), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8514), .Z(
        P2_U3573) );
  MUX2_X1 U10110 ( .A(n8866), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8514), .Z(
        P2_U3572) );
  MUX2_X1 U10111 ( .A(n8889), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8514), .Z(
        P2_U3571) );
  MUX2_X1 U10112 ( .A(n8865), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8514), .Z(
        P2_U3570) );
  MUX2_X1 U10113 ( .A(n8887), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8514), .Z(
        P2_U3569) );
  MUX2_X1 U10114 ( .A(n8515), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8514), .Z(
        P2_U3568) );
  MUX2_X1 U10115 ( .A(n8516), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8514), .Z(
        P2_U3567) );
  MUX2_X1 U10116 ( .A(n8517), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8514), .Z(
        P2_U3566) );
  MUX2_X1 U10117 ( .A(n8518), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8514), .Z(
        P2_U3565) );
  MUX2_X1 U10118 ( .A(n8519), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8514), .Z(
        P2_U3564) );
  MUX2_X1 U10119 ( .A(n8520), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8514), .Z(
        P2_U3563) );
  MUX2_X1 U10120 ( .A(n8521), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8514), .Z(
        P2_U3562) );
  MUX2_X1 U10121 ( .A(n8522), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8514), .Z(
        P2_U3561) );
  MUX2_X1 U10122 ( .A(n8523), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8514), .Z(
        P2_U3560) );
  MUX2_X1 U10123 ( .A(n8524), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8514), .Z(
        P2_U3559) );
  MUX2_X1 U10124 ( .A(n8525), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8514), .Z(
        P2_U3558) );
  MUX2_X1 U10125 ( .A(n8526), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8514), .Z(
        P2_U3557) );
  MUX2_X1 U10126 ( .A(n8527), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8514), .Z(
        P2_U3556) );
  MUX2_X1 U10127 ( .A(n6622), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8514), .Z(
        P2_U3555) );
  MUX2_X1 U10128 ( .A(n6611), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8514), .Z(
        P2_U3554) );
  MUX2_X1 U10129 ( .A(n8528), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8514), .Z(
        P2_U3553) );
  MUX2_X1 U10130 ( .A(n8529), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8514), .Z(
        P2_U3552) );
  OAI211_X1 U10131 ( .C1(n8532), .C2(n8531), .A(n8654), .B(n8530), .ZN(n8541)
         );
  NOR2_X1 U10132 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5500), .ZN(n8533) );
  AOI21_X1 U10133 ( .B1(n8685), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n8533), .ZN(
        n8540) );
  NAND2_X1 U10134 ( .A1(n8661), .A2(n8534), .ZN(n8539) );
  OAI211_X1 U10135 ( .C1(n8537), .C2(n8536), .A(n8675), .B(n8535), .ZN(n8538)
         );
  NAND4_X1 U10136 ( .A1(n8541), .A2(n8540), .A3(n8539), .A4(n8538), .ZN(
        P2_U3246) );
  OAI211_X1 U10137 ( .C1(n8543), .C2(n8542), .A(n8654), .B(n8557), .ZN(n8554)
         );
  NOR2_X1 U10138 ( .A1(n8544), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8545) );
  AOI21_X1 U10139 ( .B1(n8685), .B2(P2_ADDR_REG_2__SCAN_IN), .A(n8545), .ZN(
        n8553) );
  INV_X1 U10140 ( .A(n8546), .ZN(n8547) );
  NAND2_X1 U10141 ( .A1(n8661), .A2(n8547), .ZN(n8552) );
  OAI211_X1 U10142 ( .C1(n8550), .C2(n8549), .A(n8675), .B(n8548), .ZN(n8551)
         );
  NAND4_X1 U10143 ( .A1(n8554), .A2(n8553), .A3(n8552), .A4(n8551), .ZN(
        P2_U3247) );
  MUX2_X1 U10144 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6842), .S(n8559), .Z(n8555)
         );
  NAND3_X1 U10145 ( .A1(n8557), .A2(n8556), .A3(n8555), .ZN(n8558) );
  NAND3_X1 U10146 ( .A1(n8654), .A2(n8570), .A3(n8558), .ZN(n8567) );
  INV_X1 U10147 ( .A(n8559), .ZN(n8560) );
  NAND2_X1 U10148 ( .A1(n8661), .A2(n8560), .ZN(n8566) );
  AOI22_X1 U10149 ( .A1(n8685), .A2(P2_ADDR_REG_3__SCAN_IN), .B1(
        P2_REG3_REG_3__SCAN_IN), .B2(P2_U3152), .ZN(n8565) );
  OAI211_X1 U10150 ( .C1(n8563), .C2(n8562), .A(n8675), .B(n8561), .ZN(n8564)
         );
  NAND4_X1 U10151 ( .A1(n8567), .A2(n8566), .A3(n8565), .A4(n8564), .ZN(
        P2_U3248) );
  MUX2_X1 U10152 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6843), .S(n8568), .Z(n8571)
         );
  NAND3_X1 U10153 ( .A1(n8571), .A2(n8570), .A3(n8569), .ZN(n8572) );
  NAND3_X1 U10154 ( .A1(n8654), .A2(n8585), .A3(n8572), .ZN(n8582) );
  NAND2_X1 U10155 ( .A1(n8661), .A2(n8573), .ZN(n8581) );
  INV_X1 U10156 ( .A(n8574), .ZN(n8575) );
  AOI21_X1 U10157 ( .B1(n8685), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n8575), .ZN(
        n8580) );
  OAI211_X1 U10158 ( .C1(n8578), .C2(n8577), .A(n8675), .B(n8576), .ZN(n8579)
         );
  NAND4_X1 U10159 ( .A1(n8582), .A2(n8581), .A3(n8580), .A4(n8579), .ZN(
        P2_U3249) );
  MUX2_X1 U10160 ( .A(n6846), .B(P2_REG2_REG_5__SCAN_IN), .S(n8587), .Z(n8583)
         );
  NAND3_X1 U10161 ( .A1(n8585), .A2(n8584), .A3(n8583), .ZN(n8586) );
  NAND3_X1 U10162 ( .A1(n8654), .A2(n8598), .A3(n8586), .ZN(n8595) );
  NAND2_X1 U10163 ( .A1(n8661), .A2(n8587), .ZN(n8594) );
  NOR2_X1 U10164 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5588), .ZN(n8588) );
  AOI21_X1 U10165 ( .B1(n8685), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n8588), .ZN(
        n8593) );
  OAI211_X1 U10166 ( .C1(n8591), .C2(n8590), .A(n8675), .B(n8589), .ZN(n8592)
         );
  NAND4_X1 U10167 ( .A1(n8595), .A2(n8594), .A3(n8593), .A4(n8592), .ZN(
        P2_U3250) );
  MUX2_X1 U10168 ( .A(n7268), .B(P2_REG2_REG_6__SCAN_IN), .S(n8600), .Z(n8596)
         );
  NAND3_X1 U10169 ( .A1(n8598), .A2(n8597), .A3(n8596), .ZN(n8599) );
  NAND3_X1 U10170 ( .A1(n8654), .A2(n8612), .A3(n8599), .ZN(n8609) );
  NAND2_X1 U10171 ( .A1(n8661), .A2(n8600), .ZN(n8608) );
  INV_X1 U10172 ( .A(n8601), .ZN(n8602) );
  AOI21_X1 U10173 ( .B1(n8685), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n8602), .ZN(
        n8607) );
  OAI211_X1 U10174 ( .C1(n8605), .C2(n8604), .A(n8675), .B(n8603), .ZN(n8606)
         );
  NAND4_X1 U10175 ( .A1(n8609), .A2(n8608), .A3(n8607), .A4(n8606), .ZN(
        P2_U3251) );
  MUX2_X1 U10176 ( .A(n6851), .B(P2_REG2_REG_7__SCAN_IN), .S(n8614), .Z(n8610)
         );
  NAND3_X1 U10177 ( .A1(n8612), .A2(n8611), .A3(n8610), .ZN(n8613) );
  NAND3_X1 U10178 ( .A1(n8654), .A2(n8625), .A3(n8613), .ZN(n8622) );
  NAND2_X1 U10179 ( .A1(n8661), .A2(n8614), .ZN(n8621) );
  NOR2_X1 U10180 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5620), .ZN(n8615) );
  AOI21_X1 U10181 ( .B1(n8685), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n8615), .ZN(
        n8620) );
  OAI211_X1 U10182 ( .C1(n8618), .C2(n8617), .A(n8675), .B(n8616), .ZN(n8619)
         );
  NAND4_X1 U10183 ( .A1(n8622), .A2(n8621), .A3(n8620), .A4(n8619), .ZN(
        P2_U3252) );
  MUX2_X1 U10184 ( .A(n7310), .B(P2_REG2_REG_8__SCAN_IN), .S(n8627), .Z(n8623)
         );
  NAND3_X1 U10185 ( .A1(n8625), .A2(n8624), .A3(n8623), .ZN(n8626) );
  NAND3_X1 U10186 ( .A1(n8654), .A2(n8639), .A3(n8626), .ZN(n8636) );
  NAND2_X1 U10187 ( .A1(n8661), .A2(n8627), .ZN(n8635) );
  INV_X1 U10188 ( .A(n8628), .ZN(n8629) );
  AOI21_X1 U10189 ( .B1(n8685), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n8629), .ZN(
        n8634) );
  OAI211_X1 U10190 ( .C1(n8632), .C2(n8631), .A(n8675), .B(n8630), .ZN(n8633)
         );
  NAND4_X1 U10191 ( .A1(n8636), .A2(n8635), .A3(n8634), .A4(n8633), .ZN(
        P2_U3253) );
  MUX2_X1 U10192 ( .A(n6856), .B(P2_REG2_REG_9__SCAN_IN), .S(n9387), .Z(n8637)
         );
  NAND3_X1 U10193 ( .A1(n8639), .A2(n8638), .A3(n8637), .ZN(n8640) );
  NAND3_X1 U10194 ( .A1(n8654), .A2(n8641), .A3(n8640), .ZN(n8650) );
  NAND2_X1 U10195 ( .A1(n8661), .A2(n9387), .ZN(n8649) );
  INV_X1 U10196 ( .A(n8642), .ZN(n8643) );
  AOI21_X1 U10197 ( .B1(n8685), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n8643), .ZN(
        n8648) );
  OAI211_X1 U10198 ( .C1(n8646), .C2(n8645), .A(n8644), .B(n8675), .ZN(n8647)
         );
  NAND4_X1 U10199 ( .A1(n8650), .A2(n8649), .A3(n8648), .A4(n8647), .ZN(
        P2_U3254) );
  OAI21_X1 U10200 ( .B1(n8653), .B2(n8652), .A(n8651), .ZN(n8655) );
  NAND2_X1 U10201 ( .A1(n8655), .A2(n8654), .ZN(n8665) );
  NOR2_X1 U10202 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5724), .ZN(n8656) );
  AOI21_X1 U10203 ( .B1(n8685), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n8656), .ZN(
        n8664) );
  OAI211_X1 U10204 ( .C1(n8659), .C2(n8658), .A(n8657), .B(n8675), .ZN(n8663)
         );
  NAND2_X1 U10205 ( .A1(n8661), .A2(n8660), .ZN(n8662) );
  NAND4_X1 U10206 ( .A1(n8665), .A2(n8664), .A3(n8663), .A4(n8662), .ZN(
        P2_U3256) );
  NAND2_X1 U10207 ( .A1(n8666), .A2(n8670), .ZN(n8667) );
  NAND2_X1 U10208 ( .A1(n8668), .A2(n8667), .ZN(n8669) );
  XNOR2_X1 U10209 ( .A(n8669), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8682) );
  INV_X1 U10210 ( .A(n8682), .ZN(n8678) );
  NOR2_X1 U10211 ( .A1(n8670), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8671) );
  AOI21_X1 U10212 ( .B1(n8673), .B2(n8672), .A(n8671), .ZN(n8674) );
  XNOR2_X1 U10213 ( .A(n8674), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8680) );
  NAND2_X1 U10214 ( .A1(n8675), .A2(n8680), .ZN(n8676) );
  OAI211_X1 U10215 ( .C1(n8678), .C2(n8681), .A(n8677), .B(n8676), .ZN(n8683)
         );
  INV_X1 U10216 ( .A(P2_B_REG_SCAN_IN), .ZN(n8686) );
  NOR2_X1 U10217 ( .A1(n8687), .A2(n8686), .ZN(n8688) );
  OR2_X1 U10218 ( .A1(n8926), .A2(n8688), .ZN(n8708) );
  NOR2_X1 U10219 ( .A1(n8689), .A2(n8708), .ZN(n8968) );
  NAND2_X1 U10220 ( .A1(n8940), .A2(n8968), .ZN(n8695) );
  OAI21_X1 U10221 ( .B1(n8940), .B2(n8690), .A(n8695), .ZN(n8691) );
  AOI21_X1 U10222 ( .B1(n8963), .B2(n8951), .A(n8691), .ZN(n8692) );
  OAI21_X1 U10223 ( .B1(n8965), .B2(n8944), .A(n8692), .ZN(P2_U3265) );
  INV_X1 U10224 ( .A(n8693), .ZN(n8967) );
  NAND2_X1 U10225 ( .A1(n8702), .A2(n8694), .ZN(n8966) );
  NAND3_X1 U10226 ( .A1(n8967), .A2(n8957), .A3(n8966), .ZN(n8698) );
  INV_X1 U10227 ( .A(n8695), .ZN(n8696) );
  AOI21_X1 U10228 ( .B1(n8958), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8696), .ZN(
        n8697) );
  OAI211_X1 U10229 ( .C1(n8293), .C2(n8894), .A(n8698), .B(n8697), .ZN(
        P2_U3266) );
  NOR2_X1 U10230 ( .A1(n8976), .A2(n8973), .ZN(n8699) );
  XNOR2_X1 U10231 ( .A(n8699), .B(n5018), .ZN(n8715) );
  NAND2_X1 U10232 ( .A1(n8700), .A2(n8971), .ZN(n8701) );
  INV_X1 U10233 ( .A(n8971), .ZN(n8705) );
  AOI22_X1 U10234 ( .A1(n8703), .A2(n8871), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n8949), .ZN(n8704) );
  OAI21_X1 U10235 ( .B1(n8705), .B2(n8894), .A(n8704), .ZN(n8714) );
  NOR2_X1 U10236 ( .A1(n8706), .A2(n8975), .ZN(n8707) );
  OAI22_X1 U10237 ( .A1(n8710), .A2(n8924), .B1(n8709), .B2(n8708), .ZN(n8711)
         );
  INV_X1 U10238 ( .A(n8711), .ZN(n8712) );
  OAI21_X1 U10239 ( .B1(n8718), .B2(n8717), .A(n8716), .ZN(n8719) );
  INV_X1 U10240 ( .A(n8719), .ZN(n8988) );
  INV_X1 U10241 ( .A(n8748), .ZN(n8721) );
  AOI21_X1 U10242 ( .B1(n8984), .B2(n8721), .A(n8720), .ZN(n8985) );
  AOI22_X1 U10243 ( .A1(n8722), .A2(n8871), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n8949), .ZN(n8723) );
  OAI21_X1 U10244 ( .B1(n8724), .B2(n8894), .A(n8723), .ZN(n8731) );
  XNOR2_X1 U10245 ( .A(n8726), .B(n8725), .ZN(n8729) );
  AOI222_X1 U10246 ( .A1(n8935), .A2(n8729), .B1(n8728), .B2(n8888), .C1(n8727), .C2(n8886), .ZN(n8987) );
  NOR2_X1 U10247 ( .A1(n8987), .A2(n8949), .ZN(n8730) );
  AOI211_X1 U10248 ( .C1(n8985), .C2(n8957), .A(n8731), .B(n8730), .ZN(n8732)
         );
  OAI21_X1 U10249 ( .B1(n8988), .B2(n8899), .A(n8732), .ZN(P2_U3269) );
  OR2_X1 U10250 ( .A1(n8733), .A2(n8738), .ZN(n8734) );
  NAND2_X1 U10251 ( .A1(n8735), .A2(n8734), .ZN(n8989) );
  INV_X1 U10252 ( .A(n8989), .ZN(n8755) );
  NAND2_X1 U10253 ( .A1(n8737), .A2(n8738), .ZN(n8739) );
  NAND2_X1 U10254 ( .A1(n8736), .A2(n8739), .ZN(n8740) );
  NAND2_X1 U10255 ( .A1(n8740), .A2(n8935), .ZN(n8745) );
  OAI22_X1 U10256 ( .A1(n8742), .A2(n8926), .B1(n8741), .B2(n8924), .ZN(n8743)
         );
  INV_X1 U10257 ( .A(n8743), .ZN(n8744) );
  NAND2_X1 U10258 ( .A1(n8745), .A2(n8744), .ZN(n8992) );
  NAND2_X1 U10259 ( .A1(n8760), .A2(n8746), .ZN(n8747) );
  NAND2_X1 U10260 ( .A1(n8747), .A2(n9075), .ZN(n8749) );
  OR2_X1 U10261 ( .A1(n8749), .A2(n8748), .ZN(n8990) );
  NOR2_X1 U10262 ( .A1(n8990), .A2(n8759), .ZN(n8753) );
  AOI22_X1 U10263 ( .A1(n8750), .A2(n8871), .B1(P2_REG2_REG_26__SCAN_IN), .B2(
        n8949), .ZN(n8751) );
  OAI21_X1 U10264 ( .B1(n5269), .B2(n8894), .A(n8751), .ZN(n8752) );
  AOI211_X1 U10265 ( .C1(n8992), .C2(n8940), .A(n8753), .B(n8752), .ZN(n8754)
         );
  OAI21_X1 U10266 ( .B1(n8755), .B2(n8899), .A(n8754), .ZN(P2_U3270) );
  OAI21_X1 U10267 ( .B1(n8757), .B2(n8765), .A(n8756), .ZN(n8758) );
  INV_X1 U10268 ( .A(n8758), .ZN(n8999) );
  INV_X1 U10269 ( .A(n8759), .ZN(n8878) );
  INV_X1 U10270 ( .A(n8760), .ZN(n8761) );
  AOI211_X1 U10271 ( .C1(n8996), .C2(n8776), .A(n10530), .B(n8761), .ZN(n8995)
         );
  INV_X1 U10272 ( .A(n8996), .ZN(n8764) );
  AOI22_X1 U10273 ( .A1(n8762), .A2(n8871), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n8949), .ZN(n8763) );
  OAI21_X1 U10274 ( .B1(n8764), .B2(n8894), .A(n8763), .ZN(n8770) );
  XNOR2_X1 U10275 ( .A(n8766), .B(n8765), .ZN(n8768) );
  AOI21_X1 U10276 ( .B1(n8768), .B2(n8935), .A(n8767), .ZN(n8998) );
  NOR2_X1 U10277 ( .A1(n8998), .A2(n8958), .ZN(n8769) );
  AOI211_X1 U10278 ( .C1(n8878), .C2(n8995), .A(n8770), .B(n8769), .ZN(n8771)
         );
  OAI21_X1 U10279 ( .B1(n8999), .B2(n8899), .A(n8771), .ZN(P2_U3271) );
  INV_X1 U10280 ( .A(n8772), .ZN(n8773) );
  AOI21_X1 U10281 ( .B1(n8775), .B2(n8774), .A(n8773), .ZN(n9004) );
  INV_X1 U10282 ( .A(n8806), .ZN(n8778) );
  INV_X1 U10283 ( .A(n8776), .ZN(n8777) );
  AOI21_X1 U10284 ( .B1(n9000), .B2(n8778), .A(n8777), .ZN(n9001) );
  INV_X1 U10285 ( .A(n8779), .ZN(n8780) );
  AOI22_X1 U10286 ( .A1(n8780), .A2(n8871), .B1(n8949), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n8781) );
  OAI21_X1 U10287 ( .B1(n8782), .B2(n8894), .A(n8781), .ZN(n8789) );
  INV_X1 U10288 ( .A(n8783), .ZN(n8784) );
  AOI21_X1 U10289 ( .B1(n8784), .B2(n4587), .A(n7790), .ZN(n8787) );
  AOI21_X1 U10290 ( .B1(n8787), .B2(n8786), .A(n8785), .ZN(n9003) );
  NOR2_X1 U10291 ( .A1(n9003), .A2(n8958), .ZN(n8788) );
  AOI211_X1 U10292 ( .C1(n9001), .C2(n8957), .A(n8789), .B(n8788), .ZN(n8790)
         );
  OAI21_X1 U10293 ( .B1(n9004), .B2(n8899), .A(n8790), .ZN(P2_U3272) );
  NOR2_X1 U10294 ( .A1(n8791), .A2(n8831), .ZN(n8837) );
  NOR3_X1 U10295 ( .A1(n8837), .A2(n8823), .A3(n8822), .ZN(n8821) );
  INV_X1 U10296 ( .A(n8794), .ZN(n8793) );
  OAI21_X1 U10297 ( .B1(n8821), .B2(n8793), .A(n8803), .ZN(n8798) );
  INV_X1 U10298 ( .A(n8821), .ZN(n8796) );
  NAND3_X1 U10299 ( .A1(n8796), .A2(n8795), .A3(n8794), .ZN(n8797) );
  NAND2_X1 U10300 ( .A1(n8798), .A2(n8797), .ZN(n8800) );
  AOI222_X1 U10301 ( .A1(n8935), .A2(n8800), .B1(n8799), .B2(n8888), .C1(n8841), .C2(n8886), .ZN(n9008) );
  OAI21_X1 U10302 ( .B1(n8801), .B2(n8803), .A(n8802), .ZN(n9009) );
  INV_X1 U10303 ( .A(n9009), .ZN(n8813) );
  NOR2_X1 U10304 ( .A1(n8804), .A2(n8811), .ZN(n8805) );
  NOR2_X1 U10305 ( .A1(n8806), .A2(n8805), .ZN(n9006) );
  NAND2_X1 U10306 ( .A1(n9006), .A2(n8957), .ZN(n8810) );
  INV_X1 U10307 ( .A(n8807), .ZN(n8808) );
  AOI22_X1 U10308 ( .A1(n8958), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8808), .B2(
        n8871), .ZN(n8809) );
  OAI211_X1 U10309 ( .C1(n8811), .C2(n8894), .A(n8810), .B(n8809), .ZN(n8812)
         );
  AOI21_X1 U10310 ( .B1(n8813), .B2(n8953), .A(n8812), .ZN(n8814) );
  OAI21_X1 U10311 ( .B1(n4398), .B2(n8949), .A(n8814), .ZN(P2_U3273) );
  XNOR2_X1 U10312 ( .A(n8815), .B(n8822), .ZN(n9014) );
  INV_X1 U10313 ( .A(n8833), .ZN(n8816) );
  AOI21_X1 U10314 ( .B1(n9010), .B2(n8816), .A(n8804), .ZN(n9011) );
  INV_X1 U10315 ( .A(n8817), .ZN(n8818) );
  AOI22_X1 U10316 ( .A1(n8949), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8818), .B2(
        n8871), .ZN(n8819) );
  OAI21_X1 U10317 ( .B1(n8820), .B2(n8894), .A(n8819), .ZN(n8829) );
  NOR2_X1 U10318 ( .A1(n8821), .A2(n7790), .ZN(n8827) );
  OAI21_X1 U10319 ( .B1(n8837), .B2(n8823), .A(n8822), .ZN(n8826) );
  OAI22_X1 U10320 ( .A1(n8824), .A2(n8926), .B1(n8850), .B2(n8924), .ZN(n8825)
         );
  AOI21_X1 U10321 ( .B1(n8827), .B2(n8826), .A(n8825), .ZN(n9013) );
  NOR2_X1 U10322 ( .A1(n9013), .A2(n8949), .ZN(n8828) );
  AOI211_X1 U10323 ( .C1(n9011), .C2(n8957), .A(n8829), .B(n8828), .ZN(n8830)
         );
  OAI21_X1 U10324 ( .B1(n8899), .B2(n9014), .A(n8830), .ZN(P2_U3274) );
  XNOR2_X1 U10325 ( .A(n8832), .B(n8831), .ZN(n9019) );
  AOI21_X1 U10326 ( .B1(n9015), .B2(n8852), .A(n8833), .ZN(n9016) );
  AOI22_X1 U10327 ( .A1(n8949), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8834), .B2(
        n8871), .ZN(n8835) );
  OAI21_X1 U10328 ( .B1(n8836), .B2(n8894), .A(n8835), .ZN(n8844) );
  INV_X1 U10329 ( .A(n8837), .ZN(n8838) );
  OAI21_X1 U10330 ( .B1(n8840), .B2(n8839), .A(n8838), .ZN(n8842) );
  AOI222_X1 U10331 ( .A1(n8935), .A2(n8842), .B1(n8841), .B2(n8888), .C1(n8866), .C2(n8886), .ZN(n9018) );
  NOR2_X1 U10332 ( .A1(n9018), .A2(n8958), .ZN(n8843) );
  AOI211_X1 U10333 ( .C1(n9016), .C2(n8957), .A(n8844), .B(n8843), .ZN(n8845)
         );
  OAI21_X1 U10334 ( .B1(n8899), .B2(n9019), .A(n8845), .ZN(P2_U3275) );
  NAND2_X1 U10335 ( .A1(n8862), .A2(n8846), .ZN(n8847) );
  XNOR2_X1 U10336 ( .A(n8847), .B(n8857), .ZN(n8849) );
  OAI222_X1 U10337 ( .A1(n8926), .A2(n8850), .B1(n8849), .B2(n7790), .C1(n8924), .C2(n8848), .ZN(n9025) );
  NAND2_X1 U10338 ( .A1(n8869), .A2(n9022), .ZN(n8851) );
  NAND2_X1 U10339 ( .A1(n8852), .A2(n8851), .ZN(n9023) );
  AOI22_X1 U10340 ( .A1(n8958), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8853), .B2(
        n8871), .ZN(n8855) );
  NAND2_X1 U10341 ( .A1(n9022), .A2(n8951), .ZN(n8854) );
  OAI211_X1 U10342 ( .C1(n9023), .C2(n8944), .A(n8855), .B(n8854), .ZN(n8860)
         );
  NOR2_X1 U10343 ( .A1(n8856), .A2(n8857), .ZN(n9021) );
  INV_X1 U10344 ( .A(n8858), .ZN(n9020) );
  NOR3_X1 U10345 ( .A1(n9021), .A2(n9020), .A3(n8899), .ZN(n8859) );
  AOI211_X1 U10346 ( .C1(n8940), .C2(n9025), .A(n8860), .B(n8859), .ZN(n8861)
         );
  INV_X1 U10347 ( .A(n8861), .ZN(P2_U3276) );
  OAI21_X1 U10348 ( .B1(n8864), .B2(n8863), .A(n8862), .ZN(n8867) );
  AOI222_X1 U10349 ( .A1(n8935), .A2(n8867), .B1(n8866), .B2(n8888), .C1(n8865), .C2(n8886), .ZN(n9030) );
  AOI211_X1 U10350 ( .C1(n9028), .C2(n8868), .A(n10530), .B(n4582), .ZN(n9027)
         );
  INV_X1 U10351 ( .A(n8870), .ZN(n8872) );
  AOI22_X1 U10352 ( .A1(n8949), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8872), .B2(
        n8871), .ZN(n8873) );
  OAI21_X1 U10353 ( .B1(n4776), .B2(n8894), .A(n8873), .ZN(n8877) );
  XNOR2_X1 U10354 ( .A(n8874), .B(n8875), .ZN(n9031) );
  NOR2_X1 U10355 ( .A1(n9031), .A2(n8899), .ZN(n8876) );
  AOI211_X1 U10356 ( .C1(n9027), .C2(n8878), .A(n8877), .B(n8876), .ZN(n8879)
         );
  OAI21_X1 U10357 ( .B1(n8958), .B2(n9030), .A(n8879), .ZN(P2_U3277) );
  XOR2_X1 U10358 ( .A(n8882), .B(n8880), .Z(n9036) );
  INV_X1 U10359 ( .A(n8881), .ZN(n8906) );
  OAI21_X1 U10360 ( .B1(n8906), .B2(n8883), .A(n8882), .ZN(n8885) );
  NAND2_X1 U10361 ( .A1(n8885), .A2(n8884), .ZN(n8890) );
  AOI222_X1 U10362 ( .A1(n8935), .A2(n8890), .B1(n8889), .B2(n8888), .C1(n8887), .C2(n8886), .ZN(n9035) );
  OAI21_X1 U10363 ( .B1(n8891), .B2(n8954), .A(n9035), .ZN(n8892) );
  NAND2_X1 U10364 ( .A1(n8892), .A2(n8940), .ZN(n8898) );
  AOI21_X1 U10365 ( .B1(n9032), .B2(n4430), .A(n5259), .ZN(n9033) );
  INV_X1 U10366 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8893) );
  OAI22_X1 U10367 ( .A1(n8895), .A2(n8894), .B1(n8940), .B2(n8893), .ZN(n8896)
         );
  AOI21_X1 U10368 ( .B1(n9033), .B2(n8957), .A(n8896), .ZN(n8897) );
  OAI211_X1 U10369 ( .C1(n9036), .C2(n8899), .A(n8898), .B(n8897), .ZN(
        P2_U3278) );
  NAND2_X1 U10370 ( .A1(n8901), .A2(n8902), .ZN(n8904) );
  NAND2_X1 U10371 ( .A1(n8904), .A2(n8903), .ZN(n8905) );
  NAND2_X1 U10372 ( .A1(n8900), .A2(n8905), .ZN(n9038) );
  INV_X1 U10373 ( .A(n9038), .ZN(n8921) );
  AOI211_X1 U10374 ( .C1(n4423), .C2(n8907), .A(n7790), .B(n8906), .ZN(n8909)
         );
  OR2_X1 U10375 ( .A1(n8909), .A2(n8908), .ZN(n8914) );
  INV_X1 U10376 ( .A(n8910), .ZN(n8912) );
  XNOR2_X1 U10377 ( .A(n8936), .B(n9037), .ZN(n8911) );
  AOI21_X1 U10378 ( .B1(n9075), .B2(n8911), .A(n8914), .ZN(n9040) );
  OAI21_X1 U10379 ( .B1(n8921), .B2(n8912), .A(n9040), .ZN(n8913) );
  OAI211_X1 U10380 ( .C1(n8915), .C2(n8914), .A(n8913), .B(n8940), .ZN(n8919)
         );
  OAI22_X1 U10381 ( .A1(n8940), .A2(n7608), .B1(n8916), .B2(n8954), .ZN(n8917)
         );
  AOI21_X1 U10382 ( .B1(n9037), .B2(n8951), .A(n8917), .ZN(n8918) );
  OAI211_X1 U10383 ( .C1(n8921), .C2(n8920), .A(n8919), .B(n8918), .ZN(
        P2_U3279) );
  XNOR2_X1 U10384 ( .A(n8923), .B(n8922), .ZN(n8934) );
  OAI22_X1 U10385 ( .A1(n8927), .A2(n8926), .B1(n8925), .B2(n8924), .ZN(n8933)
         );
  NAND2_X1 U10386 ( .A1(n8929), .A2(n8928), .ZN(n8930) );
  NAND2_X1 U10387 ( .A1(n8901), .A2(n8930), .ZN(n9046) );
  NOR2_X1 U10388 ( .A1(n9046), .A2(n8931), .ZN(n8932) );
  AOI211_X1 U10389 ( .C1(n8935), .C2(n8934), .A(n8933), .B(n8932), .ZN(n9045)
         );
  INV_X1 U10390 ( .A(n9046), .ZN(n8947) );
  AND2_X1 U10391 ( .A1(n5322), .A2(n8942), .ZN(n8937) );
  OR2_X1 U10392 ( .A1(n8937), .A2(n8936), .ZN(n9042) );
  OAI22_X1 U10393 ( .A1(n8940), .A2(n8939), .B1(n8938), .B2(n8954), .ZN(n8941)
         );
  AOI21_X1 U10394 ( .B1(n8942), .B2(n8951), .A(n8941), .ZN(n8943) );
  OAI21_X1 U10395 ( .B1(n9042), .B2(n8944), .A(n8943), .ZN(n8945) );
  AOI21_X1 U10396 ( .B1(n8947), .B2(n8946), .A(n8945), .ZN(n8948) );
  OAI21_X1 U10397 ( .B1(n9045), .B2(n8949), .A(n8948), .ZN(P2_U3280) );
  AOI22_X1 U10398 ( .A1(n8953), .A2(n8952), .B1(n8951), .B2(n8950), .ZN(n8962)
         );
  NOR2_X1 U10399 ( .A1(n8954), .A2(n5500), .ZN(n8955) );
  AOI21_X1 U10400 ( .B1(n8957), .B2(n8956), .A(n8955), .ZN(n8961) );
  MUX2_X1 U10401 ( .A(n8959), .B(n6839), .S(n8958), .Z(n8960) );
  NAND3_X1 U10402 ( .A1(n8962), .A2(n8961), .A3(n8960), .ZN(P2_U3295) );
  AOI21_X1 U10403 ( .B1(n8963), .B2(n9074), .A(n8968), .ZN(n8964) );
  OAI21_X1 U10404 ( .B1(n8965), .B2(n10530), .A(n8964), .ZN(n9082) );
  MUX2_X1 U10405 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9082), .S(n10544), .Z(
        P2_U3551) );
  NAND3_X1 U10406 ( .A1(n8967), .A2(n9075), .A3(n8966), .ZN(n8970) );
  INV_X1 U10407 ( .A(n8968), .ZN(n8969) );
  OAI211_X1 U10408 ( .C1(n8293), .C2(n10528), .A(n8970), .B(n8969), .ZN(n9083)
         );
  MUX2_X1 U10409 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9083), .S(n10544), .Z(
        P2_U3550) );
  AOI22_X1 U10410 ( .A1(n8972), .A2(n9075), .B1(n9074), .B2(n8971), .ZN(n8974)
         );
  NAND3_X1 U10411 ( .A1(n8976), .A2(n5018), .A3(n10536), .ZN(n8977) );
  AOI22_X1 U10412 ( .A1(n8979), .A2(n9075), .B1(n9074), .B2(n8978), .ZN(n8980)
         );
  MUX2_X1 U10413 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9085), .S(n10544), .Z(
        P2_U3548) );
  AOI22_X1 U10414 ( .A1(n8985), .A2(n9075), .B1(n9074), .B2(n8984), .ZN(n8986)
         );
  OAI211_X1 U10415 ( .C1(n8988), .C2(n9079), .A(n8987), .B(n8986), .ZN(n9086)
         );
  MUX2_X1 U10416 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9086), .S(n10544), .Z(
        P2_U3547) );
  NAND2_X1 U10417 ( .A1(n8989), .A2(n10536), .ZN(n8994) );
  OAI21_X1 U10418 ( .B1(n5269), .B2(n10528), .A(n8990), .ZN(n8991) );
  NOR2_X1 U10419 ( .A1(n8992), .A2(n8991), .ZN(n8993) );
  NAND2_X1 U10420 ( .A1(n8994), .A2(n8993), .ZN(n9087) );
  MUX2_X1 U10421 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9087), .S(n10544), .Z(
        P2_U3546) );
  AOI21_X1 U10422 ( .B1(n9074), .B2(n8996), .A(n8995), .ZN(n8997) );
  OAI211_X1 U10423 ( .C1(n8999), .C2(n9079), .A(n8998), .B(n8997), .ZN(n9088)
         );
  MUX2_X1 U10424 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9088), .S(n10544), .Z(
        P2_U3545) );
  AOI22_X1 U10425 ( .A1(n9001), .A2(n9075), .B1(n9074), .B2(n9000), .ZN(n9002)
         );
  OAI211_X1 U10426 ( .C1(n9004), .C2(n9079), .A(n9003), .B(n9002), .ZN(n9089)
         );
  MUX2_X1 U10427 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9089), .S(n10544), .Z(
        P2_U3544) );
  AOI22_X1 U10428 ( .A1(n9006), .A2(n9075), .B1(n9074), .B2(n9005), .ZN(n9007)
         );
  OAI211_X1 U10429 ( .C1(n9079), .C2(n9009), .A(n4398), .B(n9007), .ZN(n9090)
         );
  MUX2_X1 U10430 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9090), .S(n10544), .Z(
        P2_U3543) );
  AOI22_X1 U10431 ( .A1(n9011), .A2(n9075), .B1(n9074), .B2(n9010), .ZN(n9012)
         );
  OAI211_X1 U10432 ( .C1(n9079), .C2(n9014), .A(n9013), .B(n9012), .ZN(n9091)
         );
  MUX2_X1 U10433 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9091), .S(n10544), .Z(
        P2_U3542) );
  AOI22_X1 U10434 ( .A1(n9016), .A2(n9075), .B1(n9074), .B2(n9015), .ZN(n9017)
         );
  OAI211_X1 U10435 ( .C1(n9079), .C2(n9019), .A(n9018), .B(n9017), .ZN(n9092)
         );
  MUX2_X1 U10436 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9092), .S(n10544), .Z(
        P2_U3541) );
  NOR3_X1 U10437 ( .A1(n9021), .A2(n9020), .A3(n9079), .ZN(n9026) );
  OAI22_X1 U10438 ( .A1(n9023), .A2(n10530), .B1(n4581), .B2(n10528), .ZN(
        n9024) );
  MUX2_X1 U10439 ( .A(n9093), .B(P2_REG1_REG_20__SCAN_IN), .S(n10542), .Z(
        P2_U3540) );
  AOI21_X1 U10440 ( .B1(n9074), .B2(n9028), .A(n9027), .ZN(n9029) );
  OAI211_X1 U10441 ( .C1(n9079), .C2(n9031), .A(n9030), .B(n9029), .ZN(n9094)
         );
  MUX2_X1 U10442 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9094), .S(n10544), .Z(
        P2_U3539) );
  AOI22_X1 U10443 ( .A1(n9033), .A2(n9075), .B1(n9074), .B2(n9032), .ZN(n9034)
         );
  OAI211_X1 U10444 ( .C1(n9079), .C2(n9036), .A(n9035), .B(n9034), .ZN(n9095)
         );
  MUX2_X1 U10445 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9095), .S(n10544), .Z(
        P2_U3538) );
  AOI22_X1 U10446 ( .A1(n9038), .A2(n10536), .B1(n9074), .B2(n9037), .ZN(n9039) );
  NAND2_X1 U10447 ( .A1(n9040), .A2(n9039), .ZN(n9096) );
  MUX2_X1 U10448 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9096), .S(n10544), .Z(
        P2_U3537) );
  OAI22_X1 U10449 ( .A1(n9042), .A2(n10530), .B1(n9041), .B2(n10528), .ZN(
        n9043) );
  INV_X1 U10450 ( .A(n9043), .ZN(n9044) );
  OAI211_X1 U10451 ( .C1(n9047), .C2(n9046), .A(n9045), .B(n9044), .ZN(n9097)
         );
  MUX2_X1 U10452 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9097), .S(n10544), .Z(
        P2_U3536) );
  INV_X1 U10453 ( .A(n9048), .ZN(n9053) );
  AOI22_X1 U10454 ( .A1(n9050), .A2(n9075), .B1(n9074), .B2(n9049), .ZN(n9051)
         );
  OAI211_X1 U10455 ( .C1(n9079), .C2(n9053), .A(n9052), .B(n9051), .ZN(n9098)
         );
  MUX2_X1 U10456 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9098), .S(n10544), .Z(
        P2_U3535) );
  AOI22_X1 U10457 ( .A1(n9055), .A2(n9075), .B1(n9074), .B2(n9054), .ZN(n9056)
         );
  OAI211_X1 U10458 ( .C1(n9079), .C2(n9058), .A(n9057), .B(n9056), .ZN(n9099)
         );
  MUX2_X1 U10459 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n9099), .S(n10544), .Z(
        P2_U3534) );
  OAI22_X1 U10460 ( .A1(n9060), .A2(n10530), .B1(n9059), .B2(n10528), .ZN(
        n9061) );
  AOI21_X1 U10461 ( .B1(n9063), .B2(n9062), .A(n9061), .ZN(n9064) );
  NAND2_X1 U10462 ( .A1(n9065), .A2(n9064), .ZN(n9100) );
  MUX2_X1 U10463 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n9100), .S(n10544), .Z(
        P2_U3533) );
  NAND2_X1 U10464 ( .A1(n9066), .A2(n10536), .ZN(n9069) );
  NAND2_X1 U10465 ( .A1(n9067), .A2(n9074), .ZN(n9068) );
  OAI211_X1 U10466 ( .C1(n10530), .C2(n9070), .A(n9069), .B(n9068), .ZN(n9072)
         );
  OR2_X1 U10467 ( .A1(n9072), .A2(n9071), .ZN(n9101) );
  MUX2_X1 U10468 ( .A(n9101), .B(P2_REG1_REG_12__SCAN_IN), .S(n10542), .Z(
        P2_U3532) );
  AOI22_X1 U10469 ( .A1(n9076), .A2(n9075), .B1(n9074), .B2(n9073), .ZN(n9077)
         );
  OAI211_X1 U10470 ( .C1(n9080), .C2(n9079), .A(n9078), .B(n9077), .ZN(n9102)
         );
  MUX2_X1 U10471 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n9102), .S(n10544), .Z(
        P2_U3531) );
  MUX2_X1 U10472 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n9081), .S(n10544), .Z(
        P2_U3521) );
  MUX2_X1 U10473 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9082), .S(n10538), .Z(
        P2_U3519) );
  MUX2_X1 U10474 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n9083), .S(n10538), .Z(
        P2_U3518) );
  MUX2_X1 U10475 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9086), .S(n10538), .Z(
        P2_U3515) );
  MUX2_X1 U10476 ( .A(n9087), .B(P2_REG0_REG_26__SCAN_IN), .S(n10537), .Z(
        P2_U3514) );
  MUX2_X1 U10477 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9088), .S(n10538), .Z(
        P2_U3513) );
  MUX2_X1 U10478 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9089), .S(n10538), .Z(
        P2_U3512) );
  MUX2_X1 U10479 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9090), .S(n10538), .Z(
        P2_U3511) );
  MUX2_X1 U10480 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9091), .S(n10538), .Z(
        P2_U3510) );
  MUX2_X1 U10481 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9092), .S(n10538), .Z(
        P2_U3509) );
  MUX2_X1 U10482 ( .A(n9093), .B(P2_REG0_REG_20__SCAN_IN), .S(n10537), .Z(
        P2_U3508) );
  MUX2_X1 U10483 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9094), .S(n10538), .Z(
        P2_U3507) );
  MUX2_X1 U10484 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9095), .S(n10538), .Z(
        P2_U3505) );
  MUX2_X1 U10485 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9096), .S(n10538), .Z(
        P2_U3502) );
  MUX2_X1 U10486 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9097), .S(n10538), .Z(
        P2_U3499) );
  MUX2_X1 U10487 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9098), .S(n10538), .Z(
        P2_U3496) );
  MUX2_X1 U10488 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n9099), .S(n10538), .Z(
        P2_U3493) );
  MUX2_X1 U10489 ( .A(n9100), .B(P2_REG0_REG_13__SCAN_IN), .S(n10537), .Z(
        P2_U3490) );
  MUX2_X1 U10490 ( .A(n9101), .B(P2_REG0_REG_12__SCAN_IN), .S(n10537), .Z(
        P2_U3487) );
  MUX2_X1 U10491 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n9102), .S(n10538), .Z(
        P2_U3484) );
  INV_X1 U10492 ( .A(n9560), .ZN(n10347) );
  NOR4_X1 U10493 ( .A1(n5040), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3152), .A4(
        n9103), .ZN(n9104) );
  AOI21_X1 U10494 ( .B1(n9386), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9104), .ZN(
        n9105) );
  OAI21_X1 U10495 ( .B1(n10347), .B2(n9120), .A(n9105), .ZN(P2_U3327) );
  AOI22_X1 U10496 ( .A1(n9106), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n9386), .ZN(n9107) );
  OAI21_X1 U10497 ( .B1(n9108), .B2(n9120), .A(n9107), .ZN(P2_U3328) );
  AOI22_X1 U10498 ( .A1(n5359), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n9386), .ZN(n9109) );
  OAI21_X1 U10499 ( .B1(n9110), .B2(n9120), .A(n9109), .ZN(P2_U3329) );
  NAND2_X1 U10500 ( .A1(n9386), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9111) );
  OAI211_X1 U10501 ( .C1(n9113), .C2(n9120), .A(n9112), .B(n9111), .ZN(
        P2_U3330) );
  INV_X1 U10502 ( .A(n9114), .ZN(n10351) );
  AOI22_X1 U10503 ( .A1(n9115), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n9386), .ZN(n9116) );
  OAI21_X1 U10504 ( .B1(n10351), .B2(n9120), .A(n9116), .ZN(P2_U3331) );
  INV_X1 U10505 ( .A(n9117), .ZN(n10353) );
  OAI222_X1 U10506 ( .A1(n9122), .A2(P2_U3152), .B1(n9120), .B2(n10353), .C1(
        n9119), .C2(n9118), .ZN(P2_U3332) );
  NAND4_X1 U10507 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), 
        .A3(P2_D_REG_24__SCAN_IN), .A4(P2_REG2_REG_9__SCAN_IN), .ZN(n9123) );
  NOR3_X1 U10508 ( .A1(SI_21_), .A2(P2_REG3_REG_22__SCAN_IN), .A3(n9123), .ZN(
        n9132) );
  NOR4_X1 U10509 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_REG2_REG_28__SCAN_IN), 
        .A3(SI_31_), .A4(n9327), .ZN(n9124) );
  NAND3_X1 U10510 ( .A1(SI_27_), .A2(n9124), .A3(n9296), .ZN(n9130) );
  INV_X1 U10511 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n10435) );
  NOR4_X1 U10512 ( .A1(P2_REG0_REG_13__SCAN_IN), .A2(P2_REG0_REG_2__SCAN_IN), 
        .A3(n9294), .A4(n10435), .ZN(n9128) );
  NOR4_X1 U10513 ( .A1(P1_REG2_REG_26__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), 
        .A3(n5874), .A4(n9185), .ZN(n9127) );
  NAND4_X1 U10514 ( .A1(n9188), .A2(P1_IR_REG_17__SCAN_IN), .A3(
        P1_REG3_REG_28__SCAN_IN), .A4(P2_REG3_REG_2__SCAN_IN), .ZN(n9125) );
  NOR4_X1 U10515 ( .A1(n9125), .A2(n9175), .A3(P1_REG2_REG_21__SCAN_IN), .A4(
        P2_REG2_REG_31__SCAN_IN), .ZN(n9126) );
  NAND4_X1 U10516 ( .A1(n9128), .A2(n9127), .A3(n9126), .A4(
        P2_D_REG_1__SCAN_IN), .ZN(n9129) );
  NOR4_X1 U10517 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(n6467), .A3(n9130), .A4(
        n9129), .ZN(n9131) );
  NAND4_X1 U10518 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n9132), .A3(n9131), 
        .A4(n9372), .ZN(n9171) );
  INV_X1 U10519 ( .A(n9133), .ZN(n9140) );
  NOR4_X1 U10520 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P2_ADDR_REG_17__SCAN_IN), 
        .A3(P1_ADDR_REG_7__SCAN_IN), .A4(n10584), .ZN(n9135) );
  NAND2_X1 U10521 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10375) );
  INV_X1 U10522 ( .A(n10375), .ZN(n9134) );
  NAND3_X1 U10523 ( .A1(n9227), .A2(n9135), .A3(n9134), .ZN(n9136) );
  NOR3_X1 U10524 ( .A1(n9136), .A2(P2_DATAO_REG_2__SCAN_IN), .A3(
        P2_DATAO_REG_6__SCAN_IN), .ZN(n9138) );
  NAND4_X1 U10525 ( .A1(n9138), .A2(n9137), .A3(P2_REG3_REG_6__SCAN_IN), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n9139) );
  NOR3_X1 U10526 ( .A1(n9141), .A2(n9140), .A3(n9139), .ZN(n9144) );
  NOR4_X1 U10527 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_5__SCAN_IN), .A4(n10377), .ZN(n9143) );
  INV_X1 U10528 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n9173) );
  INV_X1 U10529 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9262) );
  NOR4_X1 U10530 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(P2_ADDR_REG_13__SCAN_IN), 
        .A3(n9173), .A4(n9262), .ZN(n9142) );
  AND3_X1 U10531 ( .A1(n9144), .A2(n9143), .A3(n9142), .ZN(n9169) );
  NOR4_X1 U10532 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), 
        .A3(P2_WR_REG_SCAN_IN), .A4(n6789), .ZN(n9145) );
  NAND3_X1 U10533 ( .A1(n9145), .A2(n9283), .A3(n9281), .ZN(n9154) );
  NAND4_X1 U10534 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .A3(n6473), .A4(n9316), .ZN(n9146) );
  NOR3_X1 U10535 ( .A1(P1_REG1_REG_13__SCAN_IN), .A2(SI_29_), .A3(n9146), .ZN(
        n9152) );
  NAND4_X1 U10536 ( .A1(SI_23_), .A2(P1_REG0_REG_25__SCAN_IN), .A3(
        P1_REG0_REG_1__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n9150) );
  INV_X1 U10537 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9286) );
  INV_X1 U10538 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9569) );
  NAND4_X1 U10539 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(P2_REG0_REG_29__SCAN_IN), 
        .A3(n9286), .A4(n9569), .ZN(n9149) );
  INV_X1 U10540 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9358) );
  NAND4_X1 U10541 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(n9356), .A3(n9369), .A4(
        n9358), .ZN(n9148) );
  NAND4_X1 U10542 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(P2_REG1_REG_6__SCAN_IN), 
        .A3(P2_DATAO_REG_31__SCAN_IN), .A4(n9352), .ZN(n9147) );
  NOR4_X1 U10543 ( .A1(n9150), .A2(n9149), .A3(n9148), .A4(n9147), .ZN(n9151)
         );
  NAND4_X1 U10544 ( .A1(SI_17_), .A2(n9152), .A3(n9151), .A4(n7558), .ZN(n9153) );
  NOR4_X1 U10545 ( .A1(SI_2_), .A2(n9176), .A3(n9154), .A4(n9153), .ZN(n9168)
         );
  NAND4_X1 U10546 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(P2_REG1_REG_4__SCAN_IN), 
        .A3(n9253), .A4(n9235), .ZN(n9158) );
  NAND4_X1 U10547 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9236), .A3(n9240), .A4(
        n9238), .ZN(n9157) );
  NAND4_X1 U10548 ( .A1(n9249), .A2(n5886), .A3(n9248), .A4(
        P2_REG0_REG_24__SCAN_IN), .ZN(n9156) );
  NAND4_X1 U10549 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P2_REG2_REG_23__SCAN_IN), 
        .A3(P1_WR_REG_SCAN_IN), .A4(n9251), .ZN(n9155) );
  NOR4_X1 U10550 ( .A1(n9158), .A2(n9157), .A3(n9156), .A4(n9155), .ZN(n9167)
         );
  NOR4_X1 U10551 ( .A1(n9159), .A2(P1_IR_REG_0__SCAN_IN), .A3(
        P1_IR_REG_28__SCAN_IN), .A4(P1_REG0_REG_20__SCAN_IN), .ZN(n9165) );
  NAND4_X1 U10552 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .A3(P2_DATAO_REG_10__SCAN_IN), .A4(n9226), .ZN(n9161) );
  NAND4_X1 U10553 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_REG1_REG_10__SCAN_IN), 
        .A3(n9222), .A4(n10497), .ZN(n9160) );
  NOR4_X1 U10554 ( .A1(n9162), .A2(n9161), .A3(n9160), .A4(
        P1_IR_REG_19__SCAN_IN), .ZN(n9164) );
  AND4_X1 U10555 ( .A1(n9165), .A2(P2_REG2_REG_19__SCAN_IN), .A3(n9164), .A4(
        n9163), .ZN(n9166) );
  NAND4_X1 U10556 ( .A1(n9169), .A2(n9168), .A3(n9167), .A4(n9166), .ZN(n9170)
         );
  OAI21_X1 U10557 ( .B1(n9171), .B2(n9170), .A(P2_IR_REG_23__SCAN_IN), .ZN(
        n9279) );
  AOI22_X1 U10558 ( .A1(n9173), .A2(keyinput91), .B1(n10512), .B2(keyinput115), 
        .ZN(n9172) );
  OAI221_X1 U10559 ( .B1(n9173), .B2(keyinput91), .C1(n10512), .C2(keyinput115), .A(n9172), .ZN(n9183) );
  AOI22_X1 U10560 ( .A1(n9176), .A2(keyinput83), .B1(keyinput122), .B2(n9175), 
        .ZN(n9174) );
  OAI221_X1 U10561 ( .B1(n9176), .B2(keyinput83), .C1(n9175), .C2(keyinput122), 
        .A(n9174), .ZN(n9182) );
  XOR2_X1 U10562 ( .A(n8690), .B(keyinput123), .Z(n9180) );
  XOR2_X1 U10563 ( .A(n6008), .B(keyinput29), .Z(n9179) );
  XNOR2_X1 U10564 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput26), .ZN(n9178) );
  XNOR2_X1 U10565 ( .A(P2_IR_REG_9__SCAN_IN), .B(keyinput107), .ZN(n9177) );
  NAND4_X1 U10566 ( .A1(n9180), .A2(n9179), .A3(n9178), .A4(n9177), .ZN(n9181)
         );
  NOR3_X1 U10567 ( .A1(n9183), .A2(n9182), .A3(n9181), .ZN(n9219) );
  AOI22_X1 U10568 ( .A1(n5874), .A2(keyinput63), .B1(keyinput87), .B2(n9185), 
        .ZN(n9184) );
  OAI221_X1 U10569 ( .B1(n5874), .B2(keyinput63), .C1(n9185), .C2(keyinput87), 
        .A(n9184), .ZN(n9194) );
  INV_X1 U10570 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n10505) );
  INV_X1 U10571 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10432) );
  AOI22_X1 U10572 ( .A1(n10505), .A2(keyinput16), .B1(n10432), .B2(keyinput106), .ZN(n9186) );
  OAI221_X1 U10573 ( .B1(n10505), .B2(keyinput16), .C1(n10432), .C2(
        keyinput106), .A(n9186), .ZN(n9193) );
  AOI22_X1 U10574 ( .A1(n7947), .A2(keyinput31), .B1(n9188), .B2(keyinput127), 
        .ZN(n9187) );
  OAI221_X1 U10575 ( .B1(n7947), .B2(keyinput31), .C1(n9188), .C2(keyinput127), 
        .A(n9187), .ZN(n9192) );
  XNOR2_X1 U10576 ( .A(P1_REG3_REG_28__SCAN_IN), .B(keyinput114), .ZN(n9190)
         );
  XNOR2_X1 U10577 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput77), .ZN(n9189) );
  NAND2_X1 U10578 ( .A1(n9190), .A2(n9189), .ZN(n9191) );
  NOR4_X1 U10579 ( .A1(n9194), .A2(n9193), .A3(n9192), .A4(n9191), .ZN(n9218)
         );
  INV_X1 U10580 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10436) );
  AOI22_X1 U10581 ( .A1(n9196), .A2(keyinput76), .B1(n10436), .B2(keyinput103), 
        .ZN(n9195) );
  OAI221_X1 U10582 ( .B1(n9196), .B2(keyinput76), .C1(n10436), .C2(keyinput103), .A(n9195), .ZN(n9205) );
  INV_X1 U10583 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n9198) );
  AOI22_X1 U10584 ( .A1(n10584), .A2(keyinput58), .B1(n9198), .B2(keyinput90), 
        .ZN(n9197) );
  OAI221_X1 U10585 ( .B1(n10584), .B2(keyinput58), .C1(n9198), .C2(keyinput90), 
        .A(n9197), .ZN(n9204) );
  XOR2_X1 U10586 ( .A(n9159), .B(keyinput118), .Z(n9201) );
  XNOR2_X1 U10587 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput15), .ZN(n9200) );
  XNOR2_X1 U10588 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(keyinput53), .ZN(n9199) );
  NAND3_X1 U10589 ( .A1(n9201), .A2(n9200), .A3(n9199), .ZN(n9203) );
  XNOR2_X1 U10590 ( .A(n10377), .B(keyinput60), .ZN(n9202) );
  NOR4_X1 U10591 ( .A1(n9205), .A2(n9204), .A3(n9203), .A4(n9202), .ZN(n9217)
         );
  AOI22_X1 U10592 ( .A1(n6308), .A2(keyinput105), .B1(keyinput30), .B2(n9162), 
        .ZN(n9206) );
  OAI221_X1 U10593 ( .B1(n6308), .B2(keyinput105), .C1(n9162), .C2(keyinput30), 
        .A(n9206), .ZN(n9215) );
  XOR2_X1 U10594 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput8), .Z(n9214) );
  XNOR2_X1 U10595 ( .A(n9207), .B(keyinput36), .ZN(n9213) );
  XNOR2_X1 U10596 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput0), .ZN(n9211) );
  XNOR2_X1 U10597 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput92), .ZN(n9210) );
  XNOR2_X1 U10598 ( .A(P1_REG0_REG_20__SCAN_IN), .B(keyinput3), .ZN(n9209) );
  XNOR2_X1 U10599 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput55), .ZN(n9208) );
  NAND4_X1 U10600 ( .A1(n9211), .A2(n9210), .A3(n9209), .A4(n9208), .ZN(n9212)
         );
  NOR4_X1 U10601 ( .A1(n9215), .A2(n9214), .A3(n9213), .A4(n9212), .ZN(n9216)
         );
  NAND4_X1 U10602 ( .A1(n9219), .A2(n9218), .A3(n9217), .A4(n9216), .ZN(n9278)
         );
  INV_X1 U10603 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9221) );
  AOI22_X1 U10604 ( .A1(n9222), .A2(keyinput38), .B1(keyinput67), .B2(n9221), 
        .ZN(n9220) );
  OAI221_X1 U10605 ( .B1(n9222), .B2(keyinput38), .C1(n9221), .C2(keyinput67), 
        .A(n9220), .ZN(n9233) );
  INV_X1 U10606 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10438) );
  AOI22_X1 U10607 ( .A1(n9224), .A2(keyinput32), .B1(n10438), .B2(keyinput112), 
        .ZN(n9223) );
  OAI221_X1 U10608 ( .B1(n9224), .B2(keyinput32), .C1(n10438), .C2(keyinput112), .A(n9223), .ZN(n9232) );
  AOI22_X1 U10609 ( .A1(n9226), .A2(keyinput74), .B1(n6056), .B2(keyinput52), 
        .ZN(n9225) );
  OAI221_X1 U10610 ( .B1(n9226), .B2(keyinput74), .C1(n6056), .C2(keyinput52), 
        .A(n9225), .ZN(n9231) );
  XOR2_X1 U10611 ( .A(n9227), .B(keyinput73), .Z(n9229) );
  XNOR2_X1 U10612 ( .A(P2_IR_REG_25__SCAN_IN), .B(keyinput75), .ZN(n9228) );
  NAND2_X1 U10613 ( .A1(n9229), .A2(n9228), .ZN(n9230) );
  NOR4_X1 U10614 ( .A1(n9233), .A2(n9232), .A3(n9231), .A4(n9230), .ZN(n9276)
         );
  AOI22_X1 U10615 ( .A1(n9236), .A2(keyinput22), .B1(n9235), .B2(keyinput2), 
        .ZN(n9234) );
  OAI221_X1 U10616 ( .B1(n9236), .B2(keyinput22), .C1(n9235), .C2(keyinput2), 
        .A(n9234), .ZN(n9246) );
  AOI22_X1 U10617 ( .A1(n10497), .A2(keyinput125), .B1(keyinput116), .B2(n9238), .ZN(n9237) );
  OAI221_X1 U10618 ( .B1(n10497), .B2(keyinput125), .C1(n9238), .C2(
        keyinput116), .A(n9237), .ZN(n9245) );
  INV_X1 U10619 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n10507) );
  AOI22_X1 U10620 ( .A1(n10507), .A2(keyinput85), .B1(keyinput121), .B2(n9240), 
        .ZN(n9239) );
  OAI221_X1 U10621 ( .B1(n10507), .B2(keyinput85), .C1(n9240), .C2(keyinput121), .A(n9239), .ZN(n9244) );
  XNOR2_X1 U10622 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(keyinput13), .ZN(n9242) );
  XNOR2_X1 U10623 ( .A(SI_2_), .B(keyinput82), .ZN(n9241) );
  NAND2_X1 U10624 ( .A1(n9242), .A2(n9241), .ZN(n9243) );
  NOR4_X1 U10625 ( .A1(n9246), .A2(n9245), .A3(n9244), .A4(n9243), .ZN(n9275)
         );
  AOI22_X1 U10626 ( .A1(n9249), .A2(keyinput66), .B1(keyinput64), .B2(n9248), 
        .ZN(n9247) );
  OAI221_X1 U10627 ( .B1(n9249), .B2(keyinput66), .C1(n9248), .C2(keyinput64), 
        .A(n9247), .ZN(n9260) );
  AOI22_X1 U10628 ( .A1(n5924), .A2(keyinput117), .B1(n9251), .B2(keyinput104), 
        .ZN(n9250) );
  OAI221_X1 U10629 ( .B1(n5924), .B2(keyinput117), .C1(n9251), .C2(keyinput104), .A(n9250), .ZN(n9259) );
  AOI22_X1 U10630 ( .A1(n9254), .A2(keyinput1), .B1(n9253), .B2(keyinput11), 
        .ZN(n9252) );
  OAI221_X1 U10631 ( .B1(n9254), .B2(keyinput1), .C1(n9253), .C2(keyinput11), 
        .A(n9252), .ZN(n9258) );
  INV_X1 U10632 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10540) );
  XOR2_X1 U10633 ( .A(n10540), .B(keyinput119), .Z(n9256) );
  XNOR2_X1 U10634 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput126), .ZN(n9255) );
  NAND2_X1 U10635 ( .A1(n9256), .A2(n9255), .ZN(n9257) );
  NOR4_X1 U10636 ( .A1(n9260), .A2(n9259), .A3(n9258), .A4(n9257), .ZN(n9274)
         );
  INV_X1 U10637 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n9263) );
  AOI22_X1 U10638 ( .A1(n9263), .A2(keyinput78), .B1(keyinput42), .B2(n9262), 
        .ZN(n9261) );
  OAI221_X1 U10639 ( .B1(n9263), .B2(keyinput78), .C1(n9262), .C2(keyinput42), 
        .A(n9261), .ZN(n9272) );
  INV_X1 U10640 ( .A(P1_WR_REG_SCAN_IN), .ZN(n10400) );
  AOI22_X1 U10641 ( .A1(n10400), .A2(keyinput41), .B1(n5886), .B2(keyinput28), 
        .ZN(n9264) );
  OAI221_X1 U10642 ( .B1(n10400), .B2(keyinput41), .C1(n5886), .C2(keyinput28), 
        .A(n9264), .ZN(n9271) );
  INV_X1 U10643 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n9265) );
  XOR2_X1 U10644 ( .A(n9265), .B(keyinput35), .Z(n9269) );
  XNOR2_X1 U10645 ( .A(P1_REG3_REG_6__SCAN_IN), .B(keyinput21), .ZN(n9268) );
  XNOR2_X1 U10646 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput71), .ZN(n9267) );
  XNOR2_X1 U10647 ( .A(P2_REG0_REG_24__SCAN_IN), .B(keyinput54), .ZN(n9266) );
  NAND4_X1 U10648 ( .A1(n9269), .A2(n9268), .A3(n9267), .A4(n9266), .ZN(n9270)
         );
  NOR3_X1 U10649 ( .A1(n9272), .A2(n9271), .A3(n9270), .ZN(n9273) );
  NAND4_X1 U10650 ( .A1(n9276), .A2(n9275), .A3(n9274), .A4(n9273), .ZN(n9277)
         );
  AOI211_X1 U10651 ( .C1(keyinput102), .C2(n9279), .A(n9278), .B(n9277), .ZN(
        n9385) );
  NAND2_X1 U10652 ( .A1(n9281), .A2(keyinput70), .ZN(n9280) );
  OAI221_X1 U10653 ( .B1(n6023), .B2(keyinput102), .C1(n9281), .C2(keyinput70), 
        .A(n9280), .ZN(n9291) );
  INV_X1 U10654 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9284) );
  AOI22_X1 U10655 ( .A1(n9284), .A2(keyinput19), .B1(n9283), .B2(keyinput124), 
        .ZN(n9282) );
  OAI221_X1 U10656 ( .B1(n9284), .B2(keyinput19), .C1(n9283), .C2(keyinput124), 
        .A(n9282), .ZN(n9290) );
  AOI22_X1 U10657 ( .A1(n6565), .A2(keyinput56), .B1(n9286), .B2(keyinput18), 
        .ZN(n9285) );
  OAI221_X1 U10658 ( .B1(n6565), .B2(keyinput56), .C1(n9286), .C2(keyinput18), 
        .A(n9285), .ZN(n9289) );
  INV_X1 U10659 ( .A(P2_WR_REG_SCAN_IN), .ZN(n10399) );
  AOI22_X1 U10660 ( .A1(n10399), .A2(keyinput89), .B1(n6789), .B2(keyinput23), 
        .ZN(n9287) );
  OAI221_X1 U10661 ( .B1(n10399), .B2(keyinput89), .C1(n6789), .C2(keyinput23), 
        .A(n9287), .ZN(n9288) );
  NOR4_X1 U10662 ( .A1(n9291), .A2(n9290), .A3(n9289), .A4(n9288), .ZN(n9384)
         );
  AOI22_X1 U10663 ( .A1(n9294), .A2(keyinput12), .B1(keyinput84), .B2(n9293), 
        .ZN(n9292) );
  OAI221_X1 U10664 ( .B1(n9294), .B2(keyinput12), .C1(n9293), .C2(keyinput84), 
        .A(n9292), .ZN(n9304) );
  AOI22_X1 U10665 ( .A1(n9297), .A2(keyinput39), .B1(keyinput5), .B2(n9296), 
        .ZN(n9295) );
  OAI221_X1 U10666 ( .B1(n9297), .B2(keyinput39), .C1(n9296), .C2(keyinput5), 
        .A(n9295), .ZN(n9303) );
  INV_X1 U10667 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n10576) );
  AOI22_X1 U10668 ( .A1(n10435), .A2(keyinput40), .B1(keyinput6), .B2(n10576), 
        .ZN(n9298) );
  OAI221_X1 U10669 ( .B1(n10435), .B2(keyinput40), .C1(n10576), .C2(keyinput6), 
        .A(n9298), .ZN(n9302) );
  INV_X1 U10670 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n9300) );
  INV_X1 U10671 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10522) );
  AOI22_X1 U10672 ( .A1(n9300), .A2(keyinput10), .B1(n10522), .B2(keyinput100), 
        .ZN(n9299) );
  OAI221_X1 U10673 ( .B1(n9300), .B2(keyinput10), .C1(n10522), .C2(keyinput100), .A(n9299), .ZN(n9301) );
  NOR4_X1 U10674 ( .A1(n9304), .A2(n9303), .A3(n9302), .A4(n9301), .ZN(n9383)
         );
  INV_X1 U10675 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n10437) );
  AOI22_X1 U10676 ( .A1(n10437), .A2(keyinput24), .B1(n6068), .B2(keyinput88), 
        .ZN(n9305) );
  OAI221_X1 U10677 ( .B1(n10437), .B2(keyinput24), .C1(n6068), .C2(keyinput88), 
        .A(n9305), .ZN(n9313) );
  INV_X1 U10678 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n10502) );
  INV_X1 U10679 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n10504) );
  AOI22_X1 U10680 ( .A1(n10502), .A2(keyinput51), .B1(n10504), .B2(keyinput61), 
        .ZN(n9306) );
  OAI221_X1 U10681 ( .B1(n10502), .B2(keyinput51), .C1(n10504), .C2(keyinput61), .A(n9306), .ZN(n9312) );
  INV_X1 U10682 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n10506) );
  AOI22_X1 U10683 ( .A1(n10506), .A2(keyinput7), .B1(n6332), .B2(keyinput37), 
        .ZN(n9307) );
  OAI221_X1 U10684 ( .B1(n10506), .B2(keyinput7), .C1(n6332), .C2(keyinput37), 
        .A(n9307), .ZN(n9311) );
  INV_X1 U10685 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10549) );
  INV_X1 U10686 ( .A(SI_31_), .ZN(n9309) );
  AOI22_X1 U10687 ( .A1(n10549), .A2(keyinput79), .B1(n9309), .B2(keyinput80), 
        .ZN(n9308) );
  OAI221_X1 U10688 ( .B1(n10549), .B2(keyinput79), .C1(n9309), .C2(keyinput80), 
        .A(n9308), .ZN(n9310) );
  NOR4_X1 U10689 ( .A1(n9313), .A2(n9312), .A3(n9311), .A4(n9310), .ZN(n9346)
         );
  INV_X1 U10690 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n10430) );
  AOI22_X1 U10691 ( .A1(n10430), .A2(keyinput27), .B1(keyinput94), .B2(n10376), 
        .ZN(n9314) );
  OAI221_X1 U10692 ( .B1(n10430), .B2(keyinput27), .C1(n10376), .C2(keyinput94), .A(n9314), .ZN(n9323) );
  AOI22_X1 U10693 ( .A1(n9317), .A2(keyinput4), .B1(n9316), .B2(keyinput86), 
        .ZN(n9315) );
  OAI221_X1 U10694 ( .B1(n9317), .B2(keyinput4), .C1(n9316), .C2(keyinput86), 
        .A(n9315), .ZN(n9322) );
  AOI22_X1 U10695 ( .A1(n9320), .A2(keyinput14), .B1(n9319), .B2(keyinput46), 
        .ZN(n9318) );
  OAI221_X1 U10696 ( .B1(n9320), .B2(keyinput14), .C1(n9319), .C2(keyinput46), 
        .A(n9318), .ZN(n9321) );
  NOR3_X1 U10697 ( .A1(n9323), .A2(n9322), .A3(n9321), .ZN(n9345) );
  AOI22_X1 U10698 ( .A1(n9325), .A2(keyinput96), .B1(keyinput33), .B2(n6856), 
        .ZN(n9324) );
  OAI221_X1 U10699 ( .B1(n9325), .B2(keyinput96), .C1(n6856), .C2(keyinput33), 
        .A(n9324), .ZN(n9333) );
  AOI22_X1 U10700 ( .A1(n7997), .A2(keyinput109), .B1(keyinput34), .B2(n9327), 
        .ZN(n9326) );
  OAI221_X1 U10701 ( .B1(n7997), .B2(keyinput109), .C1(n9327), .C2(keyinput34), 
        .A(n9326), .ZN(n9332) );
  XNOR2_X1 U10702 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput20), .ZN(n9330) );
  XNOR2_X1 U10703 ( .A(P1_REG2_REG_0__SCAN_IN), .B(keyinput81), .ZN(n9329) );
  XNOR2_X1 U10704 ( .A(keyinput47), .B(P1_REG0_REG_3__SCAN_IN), .ZN(n9328) );
  NAND3_X1 U10705 ( .A1(n9330), .A2(n9329), .A3(n9328), .ZN(n9331) );
  NOR3_X1 U10706 ( .A1(n9333), .A2(n9332), .A3(n9331), .ZN(n9344) );
  AOI22_X1 U10707 ( .A1(n6266), .A2(keyinput99), .B1(n9335), .B2(keyinput62), 
        .ZN(n9334) );
  OAI221_X1 U10708 ( .B1(n6266), .B2(keyinput99), .C1(n9335), .C2(keyinput62), 
        .A(n9334), .ZN(n9342) );
  INV_X1 U10709 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10431) );
  XNOR2_X1 U10710 ( .A(n10431), .B(keyinput113), .ZN(n9341) );
  XNOR2_X1 U10711 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput108), .ZN(n9339) );
  XNOR2_X1 U10712 ( .A(P1_REG2_REG_30__SCAN_IN), .B(keyinput98), .ZN(n9338) );
  XNOR2_X1 U10713 ( .A(P2_REG1_REG_0__SCAN_IN), .B(keyinput25), .ZN(n9337) );
  XNOR2_X1 U10714 ( .A(keyinput50), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9336) );
  NAND4_X1 U10715 ( .A1(n9339), .A2(n9338), .A3(n9337), .A4(n9336), .ZN(n9340)
         );
  NOR3_X1 U10716 ( .A1(n9342), .A2(n9341), .A3(n9340), .ZN(n9343) );
  NAND4_X1 U10717 ( .A1(n9346), .A2(n9345), .A3(n9344), .A4(n9343), .ZN(n9381)
         );
  INV_X1 U10718 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10434) );
  OAI22_X1 U10719 ( .A1(n10434), .A2(keyinput120), .B1(n9348), .B2(keyinput69), 
        .ZN(n9347) );
  AOI221_X1 U10720 ( .B1(n10434), .B2(keyinput120), .C1(keyinput69), .C2(n9348), .A(n9347), .ZN(n9365) );
  OAI22_X1 U10721 ( .A1(n5464), .A2(keyinput44), .B1(n7558), .B2(keyinput72), 
        .ZN(n9349) );
  AOI221_X1 U10722 ( .B1(n5464), .B2(keyinput44), .C1(keyinput72), .C2(n7558), 
        .A(n9349), .ZN(n9364) );
  AOI22_X1 U10723 ( .A1(n9352), .A2(keyinput17), .B1(n9351), .B2(keyinput110), 
        .ZN(n9350) );
  OAI221_X1 U10724 ( .B1(n9352), .B2(keyinput17), .C1(n9351), .C2(keyinput110), 
        .A(n9350), .ZN(n9362) );
  AOI22_X1 U10725 ( .A1(n6277), .A2(keyinput101), .B1(keyinput65), .B2(n9354), 
        .ZN(n9353) );
  OAI221_X1 U10726 ( .B1(n6277), .B2(keyinput101), .C1(n9354), .C2(keyinput65), 
        .A(n9353), .ZN(n9361) );
  INV_X1 U10727 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10574) );
  AOI22_X1 U10728 ( .A1(n10574), .A2(keyinput59), .B1(n9356), .B2(keyinput97), 
        .ZN(n9355) );
  OAI221_X1 U10729 ( .B1(n10574), .B2(keyinput59), .C1(n9356), .C2(keyinput97), 
        .A(n9355), .ZN(n9360) );
  AOI22_X1 U10730 ( .A1(n6826), .A2(keyinput57), .B1(n9358), .B2(keyinput49), 
        .ZN(n9357) );
  OAI221_X1 U10731 ( .B1(n6826), .B2(keyinput57), .C1(n9358), .C2(keyinput49), 
        .A(n9357), .ZN(n9359) );
  NOR4_X1 U10732 ( .A1(n9362), .A2(n9361), .A3(n9360), .A4(n9359), .ZN(n9363)
         );
  NAND3_X1 U10733 ( .A1(n9365), .A2(n9364), .A3(n9363), .ZN(n9380) );
  INV_X1 U10734 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n10503) );
  AOI22_X1 U10735 ( .A1(n9367), .A2(keyinput111), .B1(keyinput68), .B2(n10503), 
        .ZN(n9366) );
  OAI221_X1 U10736 ( .B1(n9367), .B2(keyinput111), .C1(n10503), .C2(keyinput68), .A(n9366), .ZN(n9378) );
  INV_X1 U10737 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10433) );
  AOI22_X1 U10738 ( .A1(n10433), .A2(keyinput95), .B1(keyinput48), .B2(n9369), 
        .ZN(n9368) );
  OAI221_X1 U10739 ( .B1(n10433), .B2(keyinput95), .C1(n9369), .C2(keyinput48), 
        .A(n9368), .ZN(n9377) );
  INV_X1 U10740 ( .A(SI_21_), .ZN(n9371) );
  AOI22_X1 U10741 ( .A1(n9372), .A2(keyinput93), .B1(n9371), .B2(keyinput45), 
        .ZN(n9370) );
  OAI221_X1 U10742 ( .B1(n9372), .B2(keyinput93), .C1(n9371), .C2(keyinput45), 
        .A(n9370), .ZN(n9376) );
  AOI22_X1 U10743 ( .A1(n9473), .A2(keyinput43), .B1(n9374), .B2(keyinput9), 
        .ZN(n9373) );
  OAI221_X1 U10744 ( .B1(n9473), .B2(keyinput43), .C1(n9374), .C2(keyinput9), 
        .A(n9373), .ZN(n9375) );
  OR4_X1 U10745 ( .A1(n9378), .A2(n9377), .A3(n9376), .A4(n9375), .ZN(n9379)
         );
  NOR3_X1 U10746 ( .A1(n9381), .A2(n9380), .A3(n9379), .ZN(n9382) );
  NAND4_X1 U10747 ( .A1(n9385), .A2(n9384), .A3(n9383), .A4(n9382), .ZN(n9391)
         );
  AOI222_X1 U10748 ( .A1(n9389), .A2(n9388), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9387), .C1(P1_DATAO_REG_9__SCAN_IN), .C2(n9386), .ZN(n9390) );
  XOR2_X1 U10749 ( .A(n9391), .B(n9390), .Z(P2_U3349) );
  MUX2_X1 U10750 ( .A(n9392), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  XNOR2_X1 U10751 ( .A(n9394), .B(n9393), .ZN(n9395) );
  XNOR2_X1 U10752 ( .A(n9396), .B(n9395), .ZN(n9403) );
  NAND2_X1 U10753 ( .A1(n9841), .A2(n9511), .ZN(n9397) );
  OAI21_X1 U10754 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n9398), .A(n9397), .ZN(
        n9399) );
  AOI21_X1 U10755 ( .B1(n9970), .B2(n9550), .A(n9399), .ZN(n9400) );
  OAI21_X1 U10756 ( .B1(n9966), .B2(n9529), .A(n9400), .ZN(n9401) );
  AOI21_X1 U10757 ( .B1(n10226), .B2(n9556), .A(n9401), .ZN(n9402) );
  OAI21_X1 U10758 ( .B1(n9403), .B2(n9558), .A(n9402), .ZN(P1_U3212) );
  XNOR2_X1 U10759 ( .A(n9405), .B(n9404), .ZN(n9406) );
  XNOR2_X1 U10760 ( .A(n9407), .B(n9406), .ZN(n9412) );
  OAI22_X1 U10761 ( .A1(n9531), .A2(n10158), .B1(n9529), .B2(n10168), .ZN(
        n9410) );
  OAI21_X1 U10762 ( .B1(n9554), .B2(n10166), .A(n9408), .ZN(n9409) );
  AOI211_X1 U10763 ( .C1(n10292), .C2(n9556), .A(n9410), .B(n9409), .ZN(n9411)
         );
  OAI21_X1 U10764 ( .B1(n9412), .B2(n9558), .A(n9411), .ZN(P1_U3213) );
  INV_X1 U10765 ( .A(n9414), .ZN(n9415) );
  NOR2_X1 U10766 ( .A1(n9413), .A2(n9415), .ZN(n9516) );
  NAND2_X1 U10767 ( .A1(n9413), .A2(n9415), .ZN(n9514) );
  OAI21_X1 U10768 ( .B1(n9516), .B2(n9517), .A(n9514), .ZN(n9419) );
  XNOR2_X1 U10769 ( .A(n9417), .B(n9416), .ZN(n9418) );
  XNOR2_X1 U10770 ( .A(n9419), .B(n9418), .ZN(n9425) );
  OAI22_X1 U10771 ( .A1(n10025), .A2(n9529), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9420), .ZN(n9421) );
  AOI21_X1 U10772 ( .B1(n10018), .B2(n9550), .A(n9421), .ZN(n9422) );
  OAI21_X1 U10773 ( .B1(n10055), .B2(n9554), .A(n9422), .ZN(n9423) );
  AOI21_X1 U10774 ( .B1(n10248), .B2(n9556), .A(n9423), .ZN(n9424) );
  OAI21_X1 U10775 ( .B1(n9425), .B2(n9558), .A(n9424), .ZN(P1_U3214) );
  OAI21_X1 U10776 ( .B1(n9426), .B2(n9527), .A(n9526), .ZN(n9427) );
  OAI21_X1 U10777 ( .B1(n5194), .B2(n9428), .A(n9427), .ZN(n9432) );
  XNOR2_X1 U10778 ( .A(n9430), .B(n9429), .ZN(n9431) );
  XNOR2_X1 U10779 ( .A(n9432), .B(n9431), .ZN(n9438) );
  OAI22_X1 U10780 ( .A1(n10054), .A2(n9529), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9433), .ZN(n9436) );
  INV_X1 U10781 ( .A(n10082), .ZN(n9434) );
  OAI22_X1 U10782 ( .A1(n9554), .A2(n9482), .B1(n9531), .B2(n9434), .ZN(n9435)
         );
  AOI211_X1 U10783 ( .C1(n10265), .C2(n9556), .A(n9436), .B(n9435), .ZN(n9437)
         );
  OAI21_X1 U10784 ( .B1(n9438), .B2(n9558), .A(n9437), .ZN(P1_U3217) );
  XOR2_X1 U10785 ( .A(n9440), .B(n9439), .Z(n9445) );
  NOR2_X1 U10786 ( .A1(n10055), .A2(n9529), .ZN(n9443) );
  AOI22_X1 U10787 ( .A1(n9511), .A2(n10086), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9441) );
  OAI21_X1 U10788 ( .B1(n9531), .B2(n10061), .A(n9441), .ZN(n9442) );
  AOI211_X1 U10789 ( .C1(n10256), .C2(n9556), .A(n9443), .B(n9442), .ZN(n9444)
         );
  OAI21_X1 U10790 ( .B1(n9445), .B2(n9558), .A(n9444), .ZN(P1_U3221) );
  NAND2_X1 U10791 ( .A1(n5183), .A2(n9447), .ZN(n9448) );
  XNOR2_X1 U10792 ( .A(n4442), .B(n9448), .ZN(n9454) );
  OAI22_X1 U10793 ( .A1(n9531), .A2(n9449), .B1(n9529), .B2(n10166), .ZN(n9450) );
  AOI211_X1 U10794 ( .C1(n9511), .C2(n9846), .A(n9451), .B(n9450), .ZN(n9453)
         );
  NAND2_X1 U10795 ( .A1(n10303), .A2(n9556), .ZN(n9452) );
  OAI211_X1 U10796 ( .C1(n9454), .C2(n9558), .A(n9453), .B(n9452), .ZN(
        P1_U3222) );
  XOR2_X1 U10797 ( .A(n9456), .B(n9455), .Z(n9461) );
  NAND2_X1 U10798 ( .A1(n9841), .A2(n9551), .ZN(n9458) );
  AOI22_X1 U10799 ( .A1(n9842), .A2(n9511), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n9457) );
  OAI211_X1 U10800 ( .C1(n9531), .C2(n9998), .A(n9458), .B(n9457), .ZN(n9459)
         );
  AOI21_X1 U10801 ( .B1(n10238), .B2(n9556), .A(n9459), .ZN(n9460) );
  OAI21_X1 U10802 ( .B1(n9461), .B2(n9558), .A(n9460), .ZN(P1_U3223) );
  INV_X1 U10803 ( .A(n10282), .ZN(n10126) );
  NAND3_X1 U10804 ( .A1(n9464), .A2(n9463), .A3(n9462), .ZN(n9547) );
  AND2_X1 U10805 ( .A1(n9466), .A2(n9465), .ZN(n9545) );
  AOI21_X1 U10806 ( .B1(n9547), .B2(n9467), .A(n9545), .ZN(n9469) );
  NAND2_X1 U10807 ( .A1(n9469), .A2(n9470), .ZN(n9479) );
  INV_X1 U10808 ( .A(n9478), .ZN(n9468) );
  NOR2_X1 U10809 ( .A1(n9479), .A2(n9468), .ZN(n9472) );
  AOI21_X1 U10810 ( .B1(n9478), .B2(n9470), .A(n9469), .ZN(n9471) );
  OAI21_X1 U10811 ( .B1(n9472), .B2(n9471), .A(n9507), .ZN(n9476) );
  NOR2_X1 U10812 ( .A1(n9473), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9895) );
  OAI22_X1 U10813 ( .A1(n9554), .A2(n10168), .B1(n9531), .B2(n10127), .ZN(
        n9474) );
  AOI211_X1 U10814 ( .C1(n9551), .C2(n10102), .A(n9895), .B(n9474), .ZN(n9475)
         );
  OAI211_X1 U10815 ( .C1(n10126), .C2(n9544), .A(n9476), .B(n9475), .ZN(
        P1_U3224) );
  AND3_X1 U10816 ( .A1(n9479), .A2(n9478), .A3(n9477), .ZN(n9480) );
  OAI21_X1 U10817 ( .B1(n9480), .B2(n4444), .A(n9507), .ZN(n9486) );
  OAI22_X1 U10818 ( .A1(n9529), .A2(n9482), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9481), .ZN(n9484) );
  OAI22_X1 U10819 ( .A1(n9554), .A2(n10139), .B1(n9531), .B2(n10109), .ZN(
        n9483) );
  AOI211_X1 U10820 ( .C1(n10275), .C2(n9556), .A(n9484), .B(n9483), .ZN(n9485)
         );
  NAND2_X1 U10821 ( .A1(n9486), .A2(n9485), .ZN(P1_U3226) );
  NAND2_X1 U10822 ( .A1(n9488), .A2(n9487), .ZN(n9489) );
  XOR2_X1 U10823 ( .A(n9490), .B(n9489), .Z(n9495) );
  NAND2_X1 U10824 ( .A1(n9989), .A2(n9551), .ZN(n9492) );
  AOI22_X1 U10825 ( .A1(n10041), .A2(n9511), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9491) );
  OAI211_X1 U10826 ( .C1(n9531), .C2(n10006), .A(n9492), .B(n9491), .ZN(n9493)
         );
  AOI21_X1 U10827 ( .B1(n10243), .B2(n9556), .A(n9493), .ZN(n9494) );
  OAI21_X1 U10828 ( .B1(n9495), .B2(n9558), .A(n9494), .ZN(P1_U3227) );
  XOR2_X1 U10829 ( .A(n9497), .B(n9496), .Z(n9503) );
  OAI22_X1 U10830 ( .A1(n9521), .A2(n9529), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9498), .ZN(n9501) );
  INV_X1 U10831 ( .A(n10069), .ZN(n9499) );
  OAI22_X1 U10832 ( .A1(n9554), .A2(n9530), .B1(n9531), .B2(n9499), .ZN(n9500)
         );
  AOI211_X1 U10833 ( .C1(n10260), .C2(n9556), .A(n9501), .B(n9500), .ZN(n9502)
         );
  OAI21_X1 U10834 ( .B1(n9503), .B2(n9558), .A(n9502), .ZN(P1_U3231) );
  XNOR2_X1 U10835 ( .A(n5328), .B(n9504), .ZN(n9505) );
  XNOR2_X1 U10836 ( .A(n9506), .B(n9505), .ZN(n9508) );
  NAND2_X1 U10837 ( .A1(n9508), .A2(n9507), .ZN(n9513) );
  OAI22_X1 U10838 ( .A1(n9531), .A2(n10177), .B1(n9529), .B2(n10138), .ZN(
        n9509) );
  AOI211_X1 U10839 ( .C1(n9511), .C2(n10188), .A(n9510), .B(n9509), .ZN(n9512)
         );
  OAI211_X1 U10840 ( .C1(n10183), .C2(n9544), .A(n9513), .B(n9512), .ZN(
        P1_U3232) );
  INV_X1 U10841 ( .A(n9514), .ZN(n9515) );
  NOR2_X1 U10842 ( .A1(n9516), .A2(n9515), .ZN(n9518) );
  XNOR2_X1 U10843 ( .A(n9518), .B(n9517), .ZN(n9525) );
  OAI22_X1 U10844 ( .A1(n10012), .A2(n9529), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9519), .ZN(n9523) );
  INV_X1 U10845 ( .A(n10033), .ZN(n9520) );
  OAI22_X1 U10846 ( .A1(n9521), .A2(n9554), .B1(n9520), .B2(n9531), .ZN(n9522)
         );
  AOI211_X1 U10847 ( .C1(n5048), .C2(n9556), .A(n9523), .B(n9522), .ZN(n9524)
         );
  OAI21_X1 U10848 ( .B1(n9525), .B2(n9558), .A(n9524), .ZN(P1_U3233) );
  XNOR2_X1 U10849 ( .A(n9527), .B(n9526), .ZN(n9528) );
  XNOR2_X1 U10850 ( .A(n9426), .B(n9528), .ZN(n9535) );
  NAND2_X1 U10851 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10419)
         );
  OAI21_X1 U10852 ( .B1(n9530), .B2(n9529), .A(n10419), .ZN(n9533) );
  OAI22_X1 U10853 ( .A1(n9554), .A2(n10134), .B1(n9531), .B2(n10094), .ZN(
        n9532) );
  AOI211_X1 U10854 ( .C1(n10270), .C2(n9556), .A(n9533), .B(n9532), .ZN(n9534)
         );
  OAI21_X1 U10855 ( .B1(n9535), .B2(n9558), .A(n9534), .ZN(P1_U3236) );
  AOI21_X1 U10856 ( .B1(n9537), .B2(n9536), .A(n9558), .ZN(n9539) );
  NAND2_X1 U10857 ( .A1(n9539), .A2(n9538), .ZN(n9543) );
  AOI22_X1 U10858 ( .A1(n9982), .A2(n9550), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9540) );
  OAI21_X1 U10859 ( .B1(n10013), .B2(n9554), .A(n9540), .ZN(n9541) );
  AOI21_X1 U10860 ( .B1(n9990), .B2(n9551), .A(n9541), .ZN(n9542) );
  OAI211_X1 U10861 ( .C1(n9984), .C2(n9544), .A(n9543), .B(n9542), .ZN(
        P1_U3238) );
  INV_X1 U10862 ( .A(n9545), .ZN(n9546) );
  NAND2_X1 U10863 ( .A1(n9547), .A2(n9546), .ZN(n9549) );
  XNOR2_X1 U10864 ( .A(n9549), .B(n9548), .ZN(n9559) );
  AOI22_X1 U10865 ( .A1(n9551), .A2(n10115), .B1(n10147), .B2(n9550), .ZN(
        n9553) );
  OAI211_X1 U10866 ( .C1(n10138), .C2(n9554), .A(n9553), .B(n9552), .ZN(n9555)
         );
  AOI21_X1 U10867 ( .B1(n10285), .B2(n9556), .A(n9555), .ZN(n9557) );
  OAI21_X1 U10868 ( .B1(n9559), .B2(n9558), .A(n9557), .ZN(P1_U3239) );
  INV_X1 U10869 ( .A(n9683), .ZN(n9688) );
  MUX2_X1 U10870 ( .A(n9560), .B(P2_DATAO_REG_31__SCAN_IN), .S(n5167), .Z(
        n9561) );
  NAND2_X1 U10871 ( .A1(n9689), .A2(n9562), .ZN(n9685) );
  NAND2_X1 U10872 ( .A1(n9563), .A2(n9677), .ZN(n9566) );
  OR2_X1 U10873 ( .A1(n9680), .A2(n9564), .ZN(n9565) );
  NAND2_X1 U10874 ( .A1(n6466), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n9568) );
  NAND2_X1 U10875 ( .A1(n7974), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n9567) );
  OAI211_X1 U10876 ( .C1(n9570), .C2(n9569), .A(n9568), .B(n9567), .ZN(n9954)
         );
  INV_X1 U10877 ( .A(n9954), .ZN(n9691) );
  OR2_X1 U10878 ( .A1(n9939), .A2(n9691), .ZN(n9571) );
  NAND2_X1 U10879 ( .A1(n9685), .A2(n9571), .ZN(n9722) );
  NAND2_X1 U10880 ( .A1(n9722), .A2(n9689), .ZN(n9784) );
  NAND2_X1 U10881 ( .A1(n9954), .A2(n9936), .ZN(n9572) );
  NAND2_X1 U10882 ( .A1(n9939), .A2(n9572), .ZN(n9783) );
  NAND2_X1 U10883 ( .A1(n9784), .A2(n9783), .ZN(n9687) );
  INV_X1 U10884 ( .A(n9726), .ZN(n9573) );
  MUX2_X1 U10885 ( .A(n9573), .B(n9728), .S(n9683), .Z(n9575) );
  MUX2_X1 U10886 ( .A(n9724), .B(n9951), .S(n9683), .Z(n9574) );
  OAI21_X1 U10887 ( .B1(n9575), .B2(n9576), .A(n9574), .ZN(n9674) );
  OR2_X1 U10888 ( .A1(n9577), .A2(n9842), .ZN(n9580) );
  NAND2_X1 U10889 ( .A1(n9580), .A2(n9774), .ZN(n9661) );
  INV_X1 U10890 ( .A(n9578), .ZN(n9579) );
  OR2_X1 U10891 ( .A1(n9661), .A2(n9579), .ZN(n9664) );
  AND2_X1 U10892 ( .A1(n9665), .A2(n9580), .ZN(n9777) );
  INV_X1 U10893 ( .A(n9581), .ZN(n9755) );
  NAND4_X1 U10894 ( .A1(n9761), .A2(n9756), .A3(n9683), .A4(n9755), .ZN(n9585)
         );
  NAND3_X1 U10895 ( .A1(n9636), .A2(n9688), .A3(n9737), .ZN(n9582) );
  NOR2_X1 U10896 ( .A1(n9638), .A2(n9582), .ZN(n9583) );
  NAND2_X1 U10897 ( .A1(n9583), .A2(n9760), .ZN(n9584) );
  NAND2_X1 U10898 ( .A1(n9585), .A2(n9584), .ZN(n9642) );
  INV_X1 U10899 ( .A(n9586), .ZN(n9587) );
  NAND4_X1 U10900 ( .A1(n9611), .A2(n9591), .A3(n9688), .A4(n7184), .ZN(n9599)
         );
  NAND2_X1 U10901 ( .A1(n9848), .A2(n9683), .ZN(n9592) );
  OAI22_X1 U10902 ( .A1(n9590), .A2(n9592), .B1(n9591), .B2(n9688), .ZN(n9594)
         );
  NOR2_X1 U10903 ( .A1(n9592), .A2(n9591), .ZN(n9593) );
  AOI22_X1 U10904 ( .A1(n9595), .A2(n9594), .B1(n10481), .B2(n9593), .ZN(n9598) );
  OR3_X1 U10905 ( .A1(n7352), .A2(n9596), .A3(n9688), .ZN(n9597) );
  AND3_X1 U10906 ( .A1(n9599), .A2(n9598), .A3(n9597), .ZN(n9616) );
  INV_X1 U10907 ( .A(n9602), .ZN(n9604) );
  INV_X1 U10908 ( .A(n9808), .ZN(n9600) );
  AOI21_X1 U10909 ( .B1(n9602), .B2(n9601), .A(n9600), .ZN(n9745) );
  OAI211_X1 U10910 ( .C1(n9605), .C2(n9604), .A(n9603), .B(n9745), .ZN(n9608)
         );
  AND2_X1 U10911 ( .A1(n9607), .A2(n9606), .ZN(n9764) );
  NAND2_X1 U10912 ( .A1(n9608), .A2(n9764), .ZN(n9609) );
  NAND2_X1 U10913 ( .A1(n9609), .A2(n9733), .ZN(n9614) );
  AND2_X1 U10914 ( .A1(n9610), .A2(n9688), .ZN(n9613) );
  NAND4_X1 U10915 ( .A1(n9614), .A2(n9613), .A3(n9612), .A4(n9611), .ZN(n9615)
         );
  NAND4_X1 U10916 ( .A1(n9617), .A2(n9616), .A3(n9618), .A4(n9615), .ZN(n9622)
         );
  NOR2_X1 U10917 ( .A1(n9618), .A2(n9688), .ZN(n9619) );
  NOR2_X1 U10918 ( .A1(n9620), .A2(n9619), .ZN(n9621) );
  NOR2_X1 U10919 ( .A1(n9624), .A2(n7983), .ZN(n9735) );
  NAND2_X1 U10920 ( .A1(n9634), .A2(n9735), .ZN(n9626) );
  OR2_X1 U10921 ( .A1(n10156), .A2(n10190), .ZN(n9736) );
  NAND2_X1 U10922 ( .A1(n9633), .A2(n9627), .ZN(n9752) );
  NAND3_X1 U10923 ( .A1(n9752), .A2(n9688), .A3(n9736), .ZN(n9630) );
  AND2_X1 U10924 ( .A1(n9627), .A2(n9683), .ZN(n9632) );
  INV_X1 U10925 ( .A(n9753), .ZN(n9628) );
  NAND3_X1 U10926 ( .A1(n9633), .A2(n9632), .A3(n9628), .ZN(n9629) );
  OAI211_X1 U10927 ( .C1(n9688), .C2(n9736), .A(n9630), .B(n9629), .ZN(n9631)
         );
  INV_X1 U10928 ( .A(n9631), .ZN(n9635) );
  XNOR2_X1 U10929 ( .A(n10285), .B(n9844), .ZN(n10140) );
  INV_X1 U10930 ( .A(n9636), .ZN(n9637) );
  OR2_X1 U10931 ( .A1(n9638), .A2(n9637), .ZN(n9731) );
  NAND4_X1 U10932 ( .A1(n9643), .A2(n10098), .A3(n9731), .A4(n9683), .ZN(n9641) );
  NAND2_X1 U10933 ( .A1(n10098), .A2(n9756), .ZN(n9639) );
  NAND4_X1 U10934 ( .A1(n9760), .A2(n9688), .A3(n7986), .A4(n9639), .ZN(n9640)
         );
  NAND3_X1 U10935 ( .A1(n9656), .A2(n9657), .A3(n9643), .ZN(n9644) );
  INV_X1 U10936 ( .A(n9653), .ZN(n10050) );
  NAND3_X1 U10937 ( .A1(n9644), .A2(n10050), .A3(n9766), .ZN(n9646) );
  INV_X1 U10938 ( .A(n9655), .ZN(n9645) );
  AOI21_X1 U10939 ( .B1(n9646), .B2(n9692), .A(n9645), .ZN(n9648) );
  NAND2_X1 U10940 ( .A1(n9746), .A2(n9768), .ZN(n9647) );
  OAI21_X1 U10941 ( .B1(n9648), .B2(n9647), .A(n10021), .ZN(n9649) );
  OAI211_X1 U10942 ( .C1(n9664), .C2(n5044), .A(n9777), .B(n9650), .ZN(n9652)
         );
  NAND4_X1 U10943 ( .A1(n9652), .A2(n9651), .A3(n9688), .A4(n9985), .ZN(n9671)
         );
  AND2_X1 U10944 ( .A1(n9985), .A2(n9774), .ZN(n9663) );
  NAND2_X1 U10945 ( .A1(n9768), .A2(n9653), .ZN(n9654) );
  NAND3_X1 U10946 ( .A1(n10021), .A2(n9655), .A3(n9654), .ZN(n9775) );
  INV_X1 U10947 ( .A(n9656), .ZN(n9659) );
  NAND2_X1 U10948 ( .A1(n9766), .A2(n9760), .ZN(n9658) );
  AND2_X1 U10949 ( .A1(n9692), .A2(n9657), .ZN(n9769) );
  OAI211_X1 U10950 ( .C1(n9659), .C2(n9658), .A(n9769), .B(n9768), .ZN(n9660)
         );
  OAI211_X1 U10951 ( .C1(n9664), .C2(n10012), .A(n9663), .B(n9662), .ZN(n9666)
         );
  NAND4_X1 U10952 ( .A1(n9666), .A2(n9665), .A3(n9683), .A4(n9727), .ZN(n9670)
         );
  AND2_X1 U10953 ( .A1(n9841), .A2(n9683), .ZN(n9668) );
  OAI21_X1 U10954 ( .B1(n9841), .B2(n9683), .A(n10231), .ZN(n9667) );
  OAI21_X1 U10955 ( .B1(n9668), .B2(n10231), .A(n9667), .ZN(n9669) );
  NAND3_X1 U10956 ( .A1(n9671), .A2(n9670), .A3(n9669), .ZN(n9672) );
  NAND3_X1 U10957 ( .A1(n7971), .A2(n9820), .A3(n9672), .ZN(n9673) );
  INV_X1 U10958 ( .A(n9676), .ZN(n9675) );
  NAND2_X1 U10959 ( .A1(n9678), .A2(n9677), .ZN(n9682) );
  OR2_X1 U10960 ( .A1(n9680), .A2(n9679), .ZN(n9681) );
  INV_X1 U10961 ( .A(n9783), .ZN(n9684) );
  NAND3_X1 U10962 ( .A1(n9685), .A2(n9684), .A3(n9683), .ZN(n9686) );
  AND2_X1 U10963 ( .A1(n10200), .A2(n9936), .ZN(n9826) );
  AND2_X1 U10964 ( .A1(n9939), .A2(n9691), .ZN(n9821) );
  INV_X1 U10965 ( .A(n10047), .ZN(n10049) );
  INV_X1 U10966 ( .A(n9693), .ZN(n9706) );
  NOR2_X1 U10967 ( .A1(n9695), .A2(n9694), .ZN(n9701) );
  NOR2_X1 U10968 ( .A1(n9697), .A2(n9696), .ZN(n9700) );
  NAND4_X1 U10969 ( .A1(n9701), .A2(n9700), .A3(n9699), .A4(n9698), .ZN(n9704)
         );
  NOR3_X1 U10970 ( .A1(n9704), .A2(n9703), .A3(n9702), .ZN(n9705) );
  NAND4_X1 U10971 ( .A1(n9708), .A2(n9707), .A3(n9706), .A4(n9705), .ZN(n9709)
         );
  NOR2_X1 U10972 ( .A1(n9709), .A2(n10184), .ZN(n9712) );
  NAND3_X1 U10973 ( .A1(n9712), .A2(n9711), .A3(n9710), .ZN(n9713) );
  NOR2_X1 U10974 ( .A1(n9713), .A2(n10162), .ZN(n9714) );
  NAND4_X1 U10975 ( .A1(n10113), .A2(n9715), .A3(n9714), .A4(n10140), .ZN(
        n9716) );
  NOR2_X1 U10976 ( .A1(n9716), .A2(n10100), .ZN(n9717) );
  NAND4_X1 U10977 ( .A1(n10049), .A2(n10072), .A3(n10084), .A4(n9717), .ZN(
        n9718) );
  OR3_X1 U10978 ( .A1(n10022), .A2(n10037), .A3(n9718), .ZN(n9719) );
  NOR3_X1 U10979 ( .A1(n9996), .A2(n4720), .A3(n9719), .ZN(n9720) );
  XNOR2_X1 U10980 ( .A(n10231), .B(n9841), .ZN(n9988) );
  NAND4_X1 U10981 ( .A1(n7971), .A2(n9820), .A3(n9720), .A4(n9988), .ZN(n9721)
         );
  NOR4_X1 U10982 ( .A1(n9826), .A2(n9821), .A3(n10219), .A4(n9721), .ZN(n9723)
         );
  INV_X1 U10983 ( .A(n9722), .ZN(n9828) );
  AOI21_X1 U10984 ( .B1(n9723), .B2(n9828), .A(n6378), .ZN(n9794) );
  OR2_X1 U10985 ( .A1(n10209), .A2(n10211), .ZN(n9725) );
  AND2_X1 U10986 ( .A1(n9725), .A2(n9724), .ZN(n9796) );
  OAI211_X1 U10987 ( .C1(n9728), .C2(n9727), .A(n9951), .B(n9726), .ZN(n9730)
         );
  AND2_X1 U10988 ( .A1(n10209), .A2(n10211), .ZN(n9729) );
  AOI21_X1 U10989 ( .B1(n9796), .B2(n9730), .A(n9729), .ZN(n9823) );
  INV_X1 U10990 ( .A(n9731), .ZN(n9732) );
  NAND2_X1 U10991 ( .A1(n9732), .A2(n9760), .ZN(n9763) );
  NAND2_X1 U10992 ( .A1(n9753), .A2(n9733), .ZN(n9738) );
  NAND2_X1 U10993 ( .A1(n9735), .A2(n9734), .ZN(n9751) );
  NAND2_X1 U10994 ( .A1(n9737), .A2(n9736), .ZN(n9757) );
  OR4_X1 U10995 ( .A1(n9763), .A2(n9738), .A3(n9751), .A4(n9757), .ZN(n9765)
         );
  NAND2_X1 U10996 ( .A1(n9766), .A2(n9739), .ZN(n9740) );
  NOR2_X1 U10997 ( .A1(n9765), .A2(n9740), .ZN(n9813) );
  AND2_X1 U10998 ( .A1(n9742), .A2(n9741), .ZN(n9805) );
  NAND3_X1 U10999 ( .A1(n9743), .A2(n9805), .A3(n9810), .ZN(n9744) );
  AND3_X1 U11000 ( .A1(n9813), .A2(n9745), .A3(n9744), .ZN(n9779) );
  AND2_X1 U11001 ( .A1(n9747), .A2(n9746), .ZN(n9748) );
  AND2_X1 U11002 ( .A1(n9774), .A2(n9748), .ZN(n9776) );
  INV_X1 U11003 ( .A(n9776), .ZN(n9772) );
  OAI21_X1 U11004 ( .B1(n9751), .B2(n9750), .A(n9749), .ZN(n9754) );
  AOI21_X1 U11005 ( .B1(n9754), .B2(n9753), .A(n9752), .ZN(n9758) );
  OAI211_X1 U11006 ( .C1(n9758), .C2(n9757), .A(n9756), .B(n9755), .ZN(n9759)
         );
  INV_X1 U11007 ( .A(n9759), .ZN(n9762) );
  OAI222_X1 U11008 ( .A1(n9765), .A2(n9764), .B1(n9763), .B2(n9762), .C1(n9761), .C2(n5068), .ZN(n9767) );
  NAND2_X1 U11009 ( .A1(n9767), .A2(n9766), .ZN(n9770) );
  NAND3_X1 U11010 ( .A1(n9770), .A2(n9769), .A3(n9768), .ZN(n9771) );
  OR2_X1 U11011 ( .A1(n9772), .A2(n9771), .ZN(n9797) );
  AOI22_X1 U11012 ( .A1(n9776), .A2(n9775), .B1(n4891), .B2(n9774), .ZN(n9778)
         );
  AND2_X1 U11013 ( .A1(n9778), .A2(n9777), .ZN(n9817) );
  OAI21_X1 U11014 ( .B1(n9779), .B2(n9797), .A(n9817), .ZN(n9780) );
  NAND4_X1 U11015 ( .A1(n9796), .A2(n9819), .A3(n9781), .A4(n9780), .ZN(n9782)
         );
  NAND4_X1 U11016 ( .A1(n9823), .A2(n6378), .A3(n9783), .A4(n9782), .ZN(n9785)
         );
  OAI211_X1 U11017 ( .C1(n9826), .C2(n9785), .A(n9784), .B(n10059), .ZN(n9790)
         );
  NAND4_X1 U11018 ( .A1(n9787), .A2(n10403), .A3(n9786), .A4(n10443), .ZN(
        n9788) );
  OAI211_X1 U11019 ( .C1(n9789), .C2(n9830), .A(n9788), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9831) );
  OAI211_X1 U11020 ( .C1(n9794), .C2(n9790), .A(n9829), .B(n9831), .ZN(n9791)
         );
  NOR2_X1 U11021 ( .A1(n9792), .A2(n9791), .ZN(n9840) );
  NOR3_X1 U11022 ( .A1(n9793), .A2(n9826), .A3(n6330), .ZN(n9795) );
  OAI21_X1 U11023 ( .B1(n9795), .B2(n9794), .A(n10007), .ZN(n9839) );
  INV_X1 U11024 ( .A(n9796), .ZN(n9825) );
  INV_X1 U11025 ( .A(n9797), .ZN(n9815) );
  AND2_X1 U11026 ( .A1(n9798), .A2(n6378), .ZN(n9802) );
  OAI211_X1 U11027 ( .C1(n9802), .C2(n9801), .A(n9800), .B(n9799), .ZN(n9804)
         );
  NAND3_X1 U11028 ( .A1(n9804), .A2(n6662), .A3(n9803), .ZN(n9806) );
  NAND2_X1 U11029 ( .A1(n9806), .A2(n9805), .ZN(n9809) );
  NAND3_X1 U11030 ( .A1(n9809), .A2(n9808), .A3(n9807), .ZN(n9811) );
  NAND2_X1 U11031 ( .A1(n9811), .A2(n9810), .ZN(n9812) );
  NAND2_X1 U11032 ( .A1(n9813), .A2(n9812), .ZN(n9814) );
  NAND2_X1 U11033 ( .A1(n9815), .A2(n9814), .ZN(n9816) );
  NAND2_X1 U11034 ( .A1(n9817), .A2(n9816), .ZN(n9818) );
  NAND3_X1 U11035 ( .A1(n9820), .A2(n9819), .A3(n9818), .ZN(n9824) );
  INV_X1 U11036 ( .A(n9821), .ZN(n9822) );
  OAI211_X1 U11037 ( .C1(n9825), .C2(n9824), .A(n9823), .B(n9822), .ZN(n9827)
         );
  AOI21_X1 U11038 ( .B1(n9828), .B2(n9827), .A(n9826), .ZN(n9833) );
  INV_X1 U11039 ( .A(n9831), .ZN(n9835) );
  NOR4_X1 U11040 ( .A1(n9833), .A2(n9835), .A3(n9829), .A4(n10059), .ZN(n9838)
         );
  INV_X1 U11041 ( .A(n9830), .ZN(n9836) );
  NAND3_X1 U11042 ( .A1(n9833), .A2(n9832), .A3(n9831), .ZN(n9834) );
  OAI21_X1 U11043 ( .B1(n9836), .B2(n9835), .A(n9834), .ZN(n9837) );
  AOI211_X1 U11044 ( .C1(n9840), .C2(n9839), .A(n9838), .B(n9837), .ZN(
        P1_U3240) );
  MUX2_X1 U11045 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9954), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U11046 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n10208), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U11047 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9956), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U11048 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9990), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U11049 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9841), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U11050 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9989), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U11051 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9842), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U11052 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n10041), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U11053 ( .A(n10074), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9843), .Z(
        P1_U3576) );
  MUX2_X1 U11054 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n10086), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U11055 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n10103), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U11056 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n10116), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U11057 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n10102), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U11058 ( .A(n10115), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9843), .Z(
        P1_U3571) );
  MUX2_X1 U11059 ( .A(n9844), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9843), .Z(
        P1_U3570) );
  MUX2_X1 U11060 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n10190), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U11061 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9845), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U11062 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n10188), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U11063 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9846), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U11064 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n4701), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U11065 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9847), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U11066 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9848), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U11067 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9849), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U11068 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9850), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U11069 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9851), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U11070 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9852), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U11071 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n6659), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U11072 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9853), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U11073 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6663), .S(P1_U4006), .Z(
        P1_U3556) );
  INV_X1 U11074 ( .A(n9854), .ZN(n9856) );
  NOR3_X1 U11075 ( .A1(n9857), .A2(n9856), .A3(n9855), .ZN(n9860) );
  INV_X1 U11076 ( .A(n9858), .ZN(n9859) );
  OAI21_X1 U11077 ( .B1(n9860), .B2(n9859), .A(n10425), .ZN(n9867) );
  AOI21_X1 U11078 ( .B1(n10418), .B2(n9862), .A(n9861), .ZN(n9866) );
  MUX2_X1 U11079 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n9236), .S(n9862), .Z(n9863)
         );
  OAI211_X1 U11080 ( .C1(n4505), .C2(n9863), .A(n10416), .B(n9876), .ZN(n9865)
         );
  NAND2_X1 U11081 ( .A1(n10426), .A2(P1_ADDR_REG_9__SCAN_IN), .ZN(n9864) );
  NAND4_X1 U11082 ( .A1(n9867), .A2(n9866), .A3(n9865), .A4(n9864), .ZN(
        P1_U3250) );
  OAI21_X1 U11083 ( .B1(n9870), .B2(n9869), .A(n9868), .ZN(n9871) );
  NAND2_X1 U11084 ( .A1(n9871), .A2(n10425), .ZN(n9882) );
  AOI21_X1 U11085 ( .B1(n10418), .B2(n9873), .A(n9872), .ZN(n9881) );
  MUX2_X1 U11086 ( .A(n7207), .B(P1_REG2_REG_10__SCAN_IN), .S(n9873), .Z(n9874) );
  NAND3_X1 U11087 ( .A1(n9876), .A2(n9875), .A3(n9874), .ZN(n9877) );
  NAND3_X1 U11088 ( .A1(n9878), .A2(n10416), .A3(n9877), .ZN(n9880) );
  NAND2_X1 U11089 ( .A1(n10426), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n9879) );
  NAND4_X1 U11090 ( .A1(n9882), .A2(n9881), .A3(n9880), .A4(n9879), .ZN(
        P1_U3251) );
  INV_X1 U11091 ( .A(n9883), .ZN(n9885) );
  NAND2_X1 U11092 ( .A1(n9906), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9886) );
  OAI21_X1 U11093 ( .B1(n9906), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9886), .ZN(
        n9887) );
  AOI211_X1 U11094 ( .C1(n9888), .C2(n9887), .A(n9900), .B(n9924), .ZN(n9899)
         );
  INV_X1 U11095 ( .A(n9889), .ZN(n9892) );
  XNOR2_X1 U11096 ( .A(n9906), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n9893) );
  NOR2_X1 U11097 ( .A1(n9894), .A2(n9893), .ZN(n9905) );
  AOI211_X1 U11098 ( .C1(n9894), .C2(n9893), .A(n9905), .B(n9923), .ZN(n9898)
         );
  AOI21_X1 U11099 ( .B1(n10418), .B2(n9906), .A(n9895), .ZN(n9896) );
  OAI21_X1 U11100 ( .B1(n10411), .B2(n9221), .A(n9896), .ZN(n9897) );
  OR3_X1 U11101 ( .A1(n9899), .A2(n9898), .A3(n9897), .ZN(P1_U3257) );
  NAND2_X1 U11102 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9920), .ZN(n9901) );
  OAI21_X1 U11103 ( .B1(n9920), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9901), .ZN(
        n9902) );
  NOR2_X1 U11104 ( .A1(n9903), .A2(n9902), .ZN(n9915) );
  AOI211_X1 U11105 ( .C1(n9903), .C2(n9902), .A(n9915), .B(n9924), .ZN(n9904)
         );
  AOI21_X1 U11106 ( .B1(n10418), .B2(n9920), .A(n9904), .ZN(n9913) );
  NAND2_X1 U11107 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3084), .ZN(n9912) );
  NAND2_X1 U11108 ( .A1(n10426), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n9911) );
  AOI21_X1 U11109 ( .B1(n9906), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9905), .ZN(
        n9908) );
  XNOR2_X1 U11110 ( .A(n9920), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9907) );
  NOR2_X1 U11111 ( .A1(n9908), .A2(n9907), .ZN(n9919) );
  AOI211_X1 U11112 ( .C1(n9908), .C2(n9907), .A(n9919), .B(n9923), .ZN(n9909)
         );
  INV_X1 U11113 ( .A(n9909), .ZN(n9910) );
  NAND4_X1 U11114 ( .A1(n9913), .A2(n9912), .A3(n9911), .A4(n9910), .ZN(
        P1_U3258) );
  NAND2_X1 U11115 ( .A1(n10417), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9916) );
  OR2_X1 U11116 ( .A1(n10417), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9914) );
  NAND2_X1 U11117 ( .A1(n9916), .A2(n9914), .ZN(n10413) );
  INV_X1 U11118 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9917) );
  INV_X1 U11119 ( .A(n9929), .ZN(n9925) );
  INV_X1 U11120 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9918) );
  XNOR2_X1 U11121 ( .A(n10417), .B(n9918), .ZN(n10423) );
  NOR2_X1 U11122 ( .A1(n10417), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9921) );
  AOI21_X1 U11123 ( .B1(n10423), .B2(n10422), .A(n9921), .ZN(n9922) );
  XNOR2_X1 U11124 ( .A(n9922), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9926) );
  OAI22_X1 U11125 ( .A1(n9925), .A2(n9924), .B1(n9923), .B2(n9926), .ZN(n9932)
         );
  NAND2_X1 U11126 ( .A1(n10425), .A2(n9926), .ZN(n9927) );
  OAI211_X1 U11127 ( .C1(n9930), .C2(n9929), .A(n9928), .B(n9927), .ZN(n9931)
         );
  NAND2_X1 U11128 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3084), .ZN(n9933) );
  NAND2_X1 U11129 ( .A1(n9947), .A2(n10204), .ZN(n9934) );
  XNOR2_X1 U11130 ( .A(n9934), .B(n10200), .ZN(n10198) );
  NAND2_X1 U11131 ( .A1(n10198), .A2(n10195), .ZN(n9938) );
  AND2_X1 U11132 ( .A1(n10403), .A2(P1_B_REG_SCAN_IN), .ZN(n9935) );
  NOR2_X1 U11133 ( .A1(n10169), .A2(n9935), .ZN(n9955) );
  NAND2_X1 U11134 ( .A1(n9936), .A2(n9955), .ZN(n10202) );
  NOR2_X1 U11135 ( .A1(n10180), .A2(n10202), .ZN(n9940) );
  AOI21_X1 U11136 ( .B1(n10180), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9940), .ZN(
        n9937) );
  OAI211_X1 U11137 ( .C1(n10182), .C2(n10200), .A(n9938), .B(n9937), .ZN(
        P1_U3261) );
  XNOR2_X1 U11138 ( .A(n9947), .B(n9939), .ZN(n10201) );
  NAND2_X1 U11139 ( .A1(n10201), .A2(n10195), .ZN(n9942) );
  AOI21_X1 U11140 ( .B1(n10118), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9940), .ZN(
        n9941) );
  OAI211_X1 U11141 ( .C1(n10204), .C2(n10182), .A(n9942), .B(n9941), .ZN(
        P1_U3262) );
  INV_X1 U11142 ( .A(n10207), .ZN(n10220) );
  NAND2_X1 U11143 ( .A1(n9943), .A2(n9956), .ZN(n10218) );
  NAND2_X1 U11144 ( .A1(n10220), .A2(n10218), .ZN(n9944) );
  XNOR2_X1 U11145 ( .A(n9944), .B(n10219), .ZN(n9962) );
  NOR2_X1 U11146 ( .A1(n9947), .A2(n9946), .ZN(n10215) );
  INV_X1 U11147 ( .A(n9948), .ZN(n9949) );
  AOI22_X1 U11148 ( .A1(n9949), .A2(n10178), .B1(P1_REG2_REG_29__SCAN_IN), 
        .B2(n10118), .ZN(n9950) );
  OAI21_X1 U11149 ( .B1(n5156), .B2(n10182), .A(n9950), .ZN(n9960) );
  NAND2_X1 U11150 ( .A1(n9952), .A2(n9951), .ZN(n9953) );
  XNOR2_X1 U11151 ( .A(n9953), .B(n10205), .ZN(n9959) );
  AOI22_X1 U11152 ( .A1(n9956), .A2(n10187), .B1(n9955), .B2(n9954), .ZN(n9957) );
  OAI21_X1 U11153 ( .B1(n9962), .B2(n10197), .A(n9961), .ZN(P1_U3355) );
  XNOR2_X1 U11154 ( .A(n9963), .B(n9964), .ZN(n10230) );
  AOI21_X1 U11155 ( .B1(n9965), .B2(n9964), .A(n10165), .ZN(n9969) );
  OAI22_X1 U11156 ( .A1(n9966), .A2(n10169), .B1(n9997), .B2(n10167), .ZN(
        n9967) );
  AOI21_X1 U11157 ( .B1(n9969), .B2(n9968), .A(n9967), .ZN(n10229) );
  INV_X1 U11158 ( .A(n10229), .ZN(n9975) );
  AOI21_X1 U11159 ( .B1(n10226), .B2(n9979), .A(n4458), .ZN(n10227) );
  NAND2_X1 U11160 ( .A1(n10227), .A2(n10195), .ZN(n9972) );
  AOI22_X1 U11161 ( .A1(n9970), .A2(n10178), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n10118), .ZN(n9971) );
  OAI211_X1 U11162 ( .C1(n9973), .C2(n10182), .A(n9972), .B(n9971), .ZN(n9974)
         );
  AOI21_X1 U11163 ( .B1(n9975), .B2(n10170), .A(n9974), .ZN(n9976) );
  OAI21_X1 U11164 ( .B1(n10230), .B2(n10197), .A(n9976), .ZN(P1_U3264) );
  XNOR2_X1 U11165 ( .A(n9977), .B(n9988), .ZN(n10235) );
  INV_X1 U11166 ( .A(n9978), .ZN(n9981) );
  INV_X1 U11167 ( .A(n9979), .ZN(n9980) );
  AOI21_X1 U11168 ( .B1(n10231), .B2(n9981), .A(n9980), .ZN(n10232) );
  AOI22_X1 U11169 ( .A1(n9982), .A2(n10178), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n10118), .ZN(n9983) );
  OAI21_X1 U11170 ( .B1(n9984), .B2(n10182), .A(n9983), .ZN(n9992) );
  NAND2_X1 U11171 ( .A1(n9986), .A2(n9985), .ZN(n9987) );
  NOR2_X1 U11172 ( .A1(n10234), .A2(n10118), .ZN(n9991) );
  AOI211_X1 U11173 ( .C1(n10232), .C2(n10195), .A(n9992), .B(n9991), .ZN(n9993) );
  OAI21_X1 U11174 ( .B1(n10235), .B2(n10197), .A(n9993), .ZN(P1_U3265) );
  XOR2_X1 U11175 ( .A(n9996), .B(n9994), .Z(n10240) );
  AOI22_X1 U11176 ( .A1(n10238), .A2(n10048), .B1(n10180), .B2(
        P1_REG2_REG_25__SCAN_IN), .ZN(n10002) );
  AOI211_X1 U11177 ( .C1(n10238), .C2(n10004), .A(n10458), .B(n9978), .ZN(
        n10237) );
  INV_X1 U11178 ( .A(n10237), .ZN(n9999) );
  OAI22_X1 U11179 ( .A1(n9999), .A2(n10007), .B1(n10157), .B2(n9998), .ZN(
        n10000) );
  OAI21_X1 U11180 ( .B1(n10236), .B2(n10000), .A(n10170), .ZN(n10001) );
  OAI211_X1 U11181 ( .C1(n10240), .C2(n10197), .A(n10002), .B(n10001), .ZN(
        P1_U3266) );
  XNOR2_X1 U11182 ( .A(n10003), .B(n4720), .ZN(n10245) );
  AOI22_X1 U11183 ( .A1(n10243), .A2(n10048), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n10118), .ZN(n10016) );
  INV_X1 U11184 ( .A(n10004), .ZN(n10005) );
  AOI211_X1 U11185 ( .C1(n10243), .C2(n4526), .A(n10458), .B(n10005), .ZN(
        n10242) );
  INV_X1 U11186 ( .A(n10242), .ZN(n10008) );
  OAI22_X1 U11187 ( .A1(n10008), .A2(n10007), .B1(n10157), .B2(n10006), .ZN(
        n10014) );
  XNOR2_X1 U11188 ( .A(n10010), .B(n10009), .ZN(n10011) );
  OAI222_X1 U11189 ( .A1(n10169), .A2(n10013), .B1(n10167), .B2(n10012), .C1(
        n10011), .C2(n10165), .ZN(n10241) );
  OAI21_X1 U11190 ( .B1(n10014), .B2(n10241), .A(n10170), .ZN(n10015) );
  OAI211_X1 U11191 ( .C1(n10245), .C2(n10197), .A(n10016), .B(n10015), .ZN(
        P1_U3267) );
  XOR2_X1 U11192 ( .A(n10017), .B(n10022), .Z(n10250) );
  INV_X1 U11193 ( .A(n10018), .ZN(n10020) );
  INV_X1 U11194 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n10019) );
  OAI22_X1 U11195 ( .A1(n10020), .A2(n10157), .B1(n10019), .B2(n10170), .ZN(
        n10028) );
  AOI211_X1 U11196 ( .C1(n10248), .C2(n10031), .A(n10458), .B(n4523), .ZN(
        n10247) );
  NAND2_X1 U11197 ( .A1(n10039), .A2(n10021), .ZN(n10023) );
  XNOR2_X1 U11198 ( .A(n10023), .B(n10022), .ZN(n10024) );
  OAI222_X1 U11199 ( .A1(n10169), .A2(n10025), .B1(n10167), .B2(n10055), .C1(
        n10024), .C2(n10165), .ZN(n10246) );
  AOI21_X1 U11200 ( .B1(n10247), .B2(n10059), .A(n10246), .ZN(n10026) );
  NOR2_X1 U11201 ( .A1(n10026), .A2(n10118), .ZN(n10027) );
  AOI211_X1 U11202 ( .C1(n10048), .C2(n10248), .A(n10028), .B(n10027), .ZN(
        n10029) );
  OAI21_X1 U11203 ( .B1(n10250), .B2(n10197), .A(n10029), .ZN(P1_U3268) );
  XNOR2_X1 U11204 ( .A(n10030), .B(n10037), .ZN(n10254) );
  INV_X1 U11205 ( .A(n10031), .ZN(n10032) );
  AOI21_X1 U11206 ( .B1(n5048), .B2(n5049), .A(n10032), .ZN(n10251) );
  AOI22_X1 U11207 ( .A1(n10033), .A2(n10178), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n10118), .ZN(n10034) );
  OAI21_X1 U11208 ( .B1(n10035), .B2(n10182), .A(n10034), .ZN(n10044) );
  INV_X1 U11209 ( .A(n10036), .ZN(n10053) );
  OAI21_X1 U11210 ( .B1(n10053), .B2(n10038), .A(n10037), .ZN(n10040) );
  NAND2_X1 U11211 ( .A1(n10040), .A2(n10039), .ZN(n10042) );
  AOI222_X1 U11212 ( .A1(n10192), .A2(n10042), .B1(n10041), .B2(n10189), .C1(
        n10074), .C2(n10187), .ZN(n10253) );
  NOR2_X1 U11213 ( .A1(n10253), .A2(n10118), .ZN(n10043) );
  AOI211_X1 U11214 ( .C1(n10251), .C2(n10195), .A(n10044), .B(n10043), .ZN(
        n10045) );
  OAI21_X1 U11215 ( .B1(n10254), .B2(n10197), .A(n10045), .ZN(P1_U3269) );
  XNOR2_X1 U11216 ( .A(n10046), .B(n10047), .ZN(n10259) );
  AOI22_X1 U11217 ( .A1(n10256), .A2(n10048), .B1(n10180), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n10064) );
  AOI21_X1 U11218 ( .B1(n10051), .B2(n10050), .A(n10049), .ZN(n10052) );
  NOR3_X1 U11219 ( .A1(n10053), .A2(n10052), .A3(n10165), .ZN(n10057) );
  OAI22_X1 U11220 ( .A1(n10055), .A2(n10169), .B1(n10054), .B2(n10167), .ZN(
        n10056) );
  NOR2_X1 U11221 ( .A1(n10057), .A2(n10056), .ZN(n10258) );
  AOI211_X1 U11222 ( .C1(n10256), .C2(n10066), .A(n10458), .B(n10058), .ZN(
        n10255) );
  NAND2_X1 U11223 ( .A1(n10255), .A2(n10059), .ZN(n10060) );
  OAI211_X1 U11224 ( .C1(n10157), .C2(n10061), .A(n10258), .B(n10060), .ZN(
        n10062) );
  NAND2_X1 U11225 ( .A1(n10062), .A2(n10170), .ZN(n10063) );
  OAI211_X1 U11226 ( .C1(n10259), .C2(n10197), .A(n10064), .B(n10063), .ZN(
        P1_U3270) );
  XOR2_X1 U11227 ( .A(n10065), .B(n10072), .Z(n10264) );
  INV_X1 U11228 ( .A(n10081), .ZN(n10068) );
  INV_X1 U11229 ( .A(n10066), .ZN(n10067) );
  AOI21_X1 U11230 ( .B1(n10260), .B2(n10068), .A(n10067), .ZN(n10261) );
  AOI22_X1 U11231 ( .A1(n10180), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n10069), 
        .B2(n10178), .ZN(n10070) );
  OAI21_X1 U11232 ( .B1(n10071), .B2(n10182), .A(n10070), .ZN(n10077) );
  XNOR2_X1 U11233 ( .A(n10073), .B(n10072), .ZN(n10075) );
  AOI222_X1 U11234 ( .A1(n10192), .A2(n10075), .B1(n10074), .B2(n10189), .C1(
        n10103), .C2(n10187), .ZN(n10263) );
  NOR2_X1 U11235 ( .A1(n10263), .A2(n10118), .ZN(n10076) );
  AOI211_X1 U11236 ( .C1(n10261), .C2(n10195), .A(n10077), .B(n10076), .ZN(
        n10078) );
  OAI21_X1 U11237 ( .B1(n10264), .B2(n10197), .A(n10078), .ZN(P1_U3271) );
  XNOR2_X1 U11238 ( .A(n10079), .B(n10084), .ZN(n10269) );
  AOI21_X1 U11239 ( .B1(n10265), .B2(n10080), .A(n10081), .ZN(n10266) );
  AOI22_X1 U11240 ( .A1(n10180), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n10082), 
        .B2(n10178), .ZN(n10083) );
  OAI21_X1 U11241 ( .B1(n4525), .B2(n10182), .A(n10083), .ZN(n10089) );
  XNOR2_X1 U11242 ( .A(n10085), .B(n10084), .ZN(n10087) );
  AOI222_X1 U11243 ( .A1(n10192), .A2(n10087), .B1(n10086), .B2(n10189), .C1(
        n10116), .C2(n10187), .ZN(n10268) );
  NOR2_X1 U11244 ( .A1(n10268), .A2(n10118), .ZN(n10088) );
  AOI211_X1 U11245 ( .C1(n10266), .C2(n10195), .A(n10089), .B(n10088), .ZN(
        n10090) );
  OAI21_X1 U11246 ( .B1(n10269), .B2(n10197), .A(n10090), .ZN(P1_U3272) );
  XNOR2_X1 U11247 ( .A(n10091), .B(n10100), .ZN(n10274) );
  INV_X1 U11248 ( .A(n10108), .ZN(n10093) );
  INV_X1 U11249 ( .A(n10080), .ZN(n10092) );
  AOI21_X1 U11250 ( .B1(n10270), .B2(n10093), .A(n10092), .ZN(n10271) );
  INV_X1 U11251 ( .A(n10094), .ZN(n10095) );
  AOI22_X1 U11252 ( .A1(n10180), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n10095), 
        .B2(n10178), .ZN(n10096) );
  OAI21_X1 U11253 ( .B1(n10097), .B2(n10182), .A(n10096), .ZN(n10106) );
  NAND2_X1 U11254 ( .A1(n10099), .A2(n10098), .ZN(n10101) );
  XNOR2_X1 U11255 ( .A(n10101), .B(n10100), .ZN(n10104) );
  AOI222_X1 U11256 ( .A1(n10192), .A2(n10104), .B1(n10103), .B2(n10189), .C1(
        n10102), .C2(n10187), .ZN(n10273) );
  NOR2_X1 U11257 ( .A1(n10273), .A2(n10118), .ZN(n10105) );
  AOI211_X1 U11258 ( .C1(n10271), .C2(n10195), .A(n10106), .B(n10105), .ZN(
        n10107) );
  OAI21_X1 U11259 ( .B1(n10274), .B2(n10197), .A(n10107), .ZN(P1_U3273) );
  XNOR2_X1 U11260 ( .A(n4488), .B(n10113), .ZN(n10279) );
  AOI21_X1 U11261 ( .B1(n10275), .B2(n10124), .A(n10108), .ZN(n10276) );
  INV_X1 U11262 ( .A(n10109), .ZN(n10110) );
  AOI22_X1 U11263 ( .A1(n10180), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n10110), 
        .B2(n10178), .ZN(n10111) );
  OAI21_X1 U11264 ( .B1(n10112), .B2(n10182), .A(n10111), .ZN(n10120) );
  XNOR2_X1 U11265 ( .A(n10114), .B(n10113), .ZN(n10117) );
  AOI222_X1 U11266 ( .A1(n10192), .A2(n10117), .B1(n10116), .B2(n10189), .C1(
        n10115), .C2(n10187), .ZN(n10278) );
  NOR2_X1 U11267 ( .A1(n10278), .A2(n10118), .ZN(n10119) );
  AOI211_X1 U11268 ( .C1(n10276), .C2(n10195), .A(n10120), .B(n10119), .ZN(
        n10121) );
  OAI21_X1 U11269 ( .B1(n10197), .B2(n10279), .A(n10121), .ZN(P1_U3274) );
  XNOR2_X1 U11270 ( .A(n10122), .B(n10131), .ZN(n10284) );
  INV_X1 U11271 ( .A(n10124), .ZN(n10125) );
  AOI211_X1 U11272 ( .C1(n10282), .C2(n10123), .A(n10458), .B(n10125), .ZN(
        n10281) );
  NOR2_X1 U11273 ( .A1(n10126), .A2(n10182), .ZN(n10130) );
  OAI22_X1 U11274 ( .A1(n10170), .A2(n10128), .B1(n10127), .B2(n10157), .ZN(
        n10129) );
  AOI211_X1 U11275 ( .C1(n10281), .C2(n10161), .A(n10130), .B(n10129), .ZN(
        n10136) );
  XNOR2_X1 U11276 ( .A(n10132), .B(n10131), .ZN(n10133) );
  OAI222_X1 U11277 ( .A1(n10169), .A2(n10134), .B1(n10167), .B2(n10168), .C1(
        n10133), .C2(n10165), .ZN(n10280) );
  NAND2_X1 U11278 ( .A1(n10280), .A2(n10170), .ZN(n10135) );
  OAI211_X1 U11279 ( .C1(n10284), .C2(n10197), .A(n10136), .B(n10135), .ZN(
        P1_U3275) );
  XOR2_X1 U11280 ( .A(n10137), .B(n10140), .Z(n10144) );
  OAI22_X1 U11281 ( .A1(n10139), .A2(n10169), .B1(n10138), .B2(n10167), .ZN(
        n10143) );
  XNOR2_X1 U11282 ( .A(n10141), .B(n10140), .ZN(n10289) );
  NOR2_X1 U11283 ( .A1(n10289), .A2(n6661), .ZN(n10142) );
  AOI211_X1 U11284 ( .C1(n10144), .C2(n10192), .A(n10143), .B(n10142), .ZN(
        n10288) );
  INV_X1 U11285 ( .A(n10155), .ZN(n10146) );
  INV_X1 U11286 ( .A(n10123), .ZN(n10145) );
  AOI21_X1 U11287 ( .B1(n10285), .B2(n10146), .A(n10145), .ZN(n10286) );
  AOI22_X1 U11288 ( .A1(n10180), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n10147), 
        .B2(n10178), .ZN(n10148) );
  OAI21_X1 U11289 ( .B1(n10149), .B2(n10182), .A(n10148), .ZN(n10152) );
  NOR2_X1 U11290 ( .A1(n10289), .A2(n10150), .ZN(n10151) );
  AOI211_X1 U11291 ( .C1(n10286), .C2(n10195), .A(n10152), .B(n10151), .ZN(
        n10153) );
  OAI21_X1 U11292 ( .B1(n10288), .B2(n10118), .A(n10153), .ZN(P1_U3276) );
  XNOR2_X1 U11293 ( .A(n10154), .B(n10162), .ZN(n10294) );
  AOI211_X1 U11294 ( .C1(n10292), .C2(n10174), .A(n10458), .B(n10155), .ZN(
        n10291) );
  NOR2_X1 U11295 ( .A1(n10156), .A2(n10182), .ZN(n10160) );
  OAI22_X1 U11296 ( .A1(n10170), .A2(n7154), .B1(n10158), .B2(n10157), .ZN(
        n10159) );
  AOI211_X1 U11297 ( .C1(n10291), .C2(n10161), .A(n10160), .B(n10159), .ZN(
        n10172) );
  XNOR2_X1 U11298 ( .A(n10163), .B(n10162), .ZN(n10164) );
  OAI222_X1 U11299 ( .A1(n10169), .A2(n10168), .B1(n10167), .B2(n10166), .C1(
        n10165), .C2(n10164), .ZN(n10290) );
  NAND2_X1 U11300 ( .A1(n10290), .A2(n10170), .ZN(n10171) );
  OAI211_X1 U11301 ( .C1(n10294), .C2(n10197), .A(n10172), .B(n10171), .ZN(
        P1_U3277) );
  XOR2_X1 U11302 ( .A(n10184), .B(n10173), .Z(n10300) );
  INV_X1 U11303 ( .A(n10174), .ZN(n10175) );
  AOI21_X1 U11304 ( .B1(n10295), .B2(n10176), .A(n10175), .ZN(n10296) );
  INV_X1 U11305 ( .A(n10177), .ZN(n10179) );
  AOI22_X1 U11306 ( .A1(n10180), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n10179), 
        .B2(n10178), .ZN(n10181) );
  OAI21_X1 U11307 ( .B1(n10183), .B2(n10182), .A(n10181), .ZN(n10194) );
  OAI21_X1 U11308 ( .B1(n10186), .B2(n7985), .A(n10185), .ZN(n10191) );
  AOI222_X1 U11309 ( .A1(n10192), .A2(n10191), .B1(n10190), .B2(n10189), .C1(
        n10188), .C2(n10187), .ZN(n10298) );
  NOR2_X1 U11310 ( .A1(n10298), .A2(n10118), .ZN(n10193) );
  AOI211_X1 U11311 ( .C1(n10296), .C2(n10195), .A(n10194), .B(n10193), .ZN(
        n10196) );
  OAI21_X1 U11312 ( .B1(n10197), .B2(n10300), .A(n10196), .ZN(P1_U3278) );
  NAND2_X1 U11313 ( .A1(n10198), .A2(n10464), .ZN(n10199) );
  OAI211_X1 U11314 ( .C1(n10200), .C2(n10480), .A(n10199), .B(n10202), .ZN(
        n10321) );
  MUX2_X1 U11315 ( .A(n10321), .B(P1_REG1_REG_31__SCAN_IN), .S(n10496), .Z(
        P1_U3554) );
  NAND2_X1 U11316 ( .A1(n10201), .A2(n10464), .ZN(n10203) );
  OAI211_X1 U11317 ( .C1(n10204), .C2(n10480), .A(n10203), .B(n10202), .ZN(
        n10322) );
  MUX2_X1 U11318 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n10322), .S(n10499), .Z(
        P1_U3553) );
  NAND2_X1 U11319 ( .A1(n10208), .A2(n10476), .ZN(n10210) );
  OAI211_X1 U11320 ( .C1(n10218), .C2(n10210), .A(n10209), .B(n10480), .ZN(
        n10214) );
  NAND2_X1 U11321 ( .A1(n10211), .A2(n10476), .ZN(n10212) );
  OAI21_X1 U11322 ( .B1(n10218), .B2(n10212), .A(n5156), .ZN(n10213) );
  OAI22_X1 U11323 ( .A1(n10222), .A2(n10458), .B1(n10221), .B2(n10480), .ZN(
        n10223) );
  MUX2_X1 U11324 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n10324), .S(n10499), .Z(
        P1_U3551) );
  AOI22_X1 U11325 ( .A1(n10227), .A2(n10464), .B1(n10463), .B2(n10226), .ZN(
        n10228) );
  OAI211_X1 U11326 ( .C1(n10230), .C2(n10299), .A(n10229), .B(n10228), .ZN(
        n10325) );
  MUX2_X1 U11327 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10325), .S(n10499), .Z(
        P1_U3550) );
  AOI22_X1 U11328 ( .A1(n10232), .A2(n10464), .B1(n10463), .B2(n10231), .ZN(
        n10233) );
  OAI211_X1 U11329 ( .C1(n10235), .C2(n10299), .A(n10234), .B(n10233), .ZN(
        n10326) );
  MUX2_X1 U11330 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10326), .S(n10499), .Z(
        P1_U3549) );
  AOI211_X1 U11331 ( .C1(n10463), .C2(n10238), .A(n10237), .B(n10236), .ZN(
        n10239) );
  AOI211_X1 U11332 ( .C1(n10463), .C2(n10243), .A(n10242), .B(n10241), .ZN(
        n10244) );
  OAI21_X1 U11333 ( .B1(n10245), .B2(n10299), .A(n10244), .ZN(n10328) );
  MUX2_X1 U11334 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10328), .S(n10499), .Z(
        P1_U3547) );
  AOI211_X1 U11335 ( .C1(n10463), .C2(n10248), .A(n10247), .B(n10246), .ZN(
        n10249) );
  OAI21_X1 U11336 ( .B1(n10250), .B2(n10299), .A(n10249), .ZN(n10329) );
  MUX2_X1 U11337 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10329), .S(n10499), .Z(
        P1_U3546) );
  AOI22_X1 U11338 ( .A1(n10251), .A2(n10464), .B1(n10463), .B2(n5048), .ZN(
        n10252) );
  OAI211_X1 U11339 ( .C1(n10254), .C2(n10299), .A(n10253), .B(n10252), .ZN(
        n10330) );
  MUX2_X1 U11340 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10330), .S(n10499), .Z(
        P1_U3545) );
  AOI21_X1 U11341 ( .B1(n10463), .B2(n10256), .A(n10255), .ZN(n10257) );
  OAI211_X1 U11342 ( .C1(n10259), .C2(n10299), .A(n10258), .B(n10257), .ZN(
        n10331) );
  MUX2_X1 U11343 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10331), .S(n10499), .Z(
        P1_U3544) );
  AOI22_X1 U11344 ( .A1(n10261), .A2(n10464), .B1(n10463), .B2(n10260), .ZN(
        n10262) );
  OAI211_X1 U11345 ( .C1(n10264), .C2(n10299), .A(n10263), .B(n10262), .ZN(
        n10332) );
  MUX2_X1 U11346 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10332), .S(n10499), .Z(
        P1_U3543) );
  AOI22_X1 U11347 ( .A1(n10266), .A2(n10464), .B1(n10463), .B2(n10265), .ZN(
        n10267) );
  OAI211_X1 U11348 ( .C1(n10269), .C2(n10299), .A(n10268), .B(n10267), .ZN(
        n10333) );
  MUX2_X1 U11349 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10333), .S(n10499), .Z(
        P1_U3542) );
  AOI22_X1 U11350 ( .A1(n10271), .A2(n10464), .B1(n10463), .B2(n10270), .ZN(
        n10272) );
  OAI211_X1 U11351 ( .C1(n10274), .C2(n10299), .A(n10273), .B(n10272), .ZN(
        n10334) );
  MUX2_X1 U11352 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10334), .S(n10499), .Z(
        P1_U3541) );
  AOI22_X1 U11353 ( .A1(n10276), .A2(n10464), .B1(n10463), .B2(n10275), .ZN(
        n10277) );
  OAI211_X1 U11354 ( .C1(n10279), .C2(n10299), .A(n10278), .B(n10277), .ZN(
        n10335) );
  MUX2_X1 U11355 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10335), .S(n10499), .Z(
        P1_U3540) );
  AOI211_X1 U11356 ( .C1(n10463), .C2(n10282), .A(n10281), .B(n10280), .ZN(
        n10283) );
  OAI21_X1 U11357 ( .B1(n10284), .B2(n10299), .A(n10283), .ZN(n10336) );
  MUX2_X1 U11358 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10336), .S(n10499), .Z(
        P1_U3539) );
  AOI22_X1 U11359 ( .A1(n10286), .A2(n10464), .B1(n10463), .B2(n10285), .ZN(
        n10287) );
  OAI211_X1 U11360 ( .C1(n10468), .C2(n10289), .A(n10288), .B(n10287), .ZN(
        n10337) );
  MUX2_X1 U11361 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n10337), .S(n10499), .Z(
        P1_U3538) );
  AOI211_X1 U11362 ( .C1(n10463), .C2(n10292), .A(n10291), .B(n10290), .ZN(
        n10293) );
  OAI21_X1 U11363 ( .B1(n10294), .B2(n10299), .A(n10293), .ZN(n10338) );
  MUX2_X1 U11364 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10338), .S(n10499), .Z(
        P1_U3537) );
  AOI22_X1 U11365 ( .A1(n10296), .A2(n10464), .B1(n10463), .B2(n10295), .ZN(
        n10297) );
  OAI211_X1 U11366 ( .C1(n10300), .C2(n10299), .A(n10298), .B(n10297), .ZN(
        n10339) );
  MUX2_X1 U11367 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n10339), .S(n10499), .Z(
        P1_U3536) );
  NAND2_X1 U11368 ( .A1(n10301), .A2(n10476), .ZN(n10306) );
  AOI21_X1 U11369 ( .B1(n10463), .B2(n10303), .A(n10302), .ZN(n10304) );
  OAI211_X1 U11370 ( .C1(n10307), .C2(n10306), .A(n10305), .B(n10304), .ZN(
        n10340) );
  MUX2_X1 U11371 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10340), .S(n10499), .Z(
        P1_U3535) );
  INV_X1 U11372 ( .A(n10308), .ZN(n10313) );
  OAI22_X1 U11373 ( .A1(n10310), .A2(n10458), .B1(n10309), .B2(n10480), .ZN(
        n10312) );
  AOI211_X1 U11374 ( .C1(n10485), .C2(n10313), .A(n10312), .B(n10311), .ZN(
        n10314) );
  INV_X1 U11375 ( .A(n10314), .ZN(n10341) );
  MUX2_X1 U11376 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10341), .S(n10499), .Z(
        P1_U3534) );
  AOI21_X1 U11377 ( .B1(n10463), .B2(n7352), .A(n10315), .ZN(n10318) );
  INV_X1 U11378 ( .A(n10316), .ZN(n10317) );
  OAI211_X1 U11379 ( .C1(n10319), .C2(n10468), .A(n10318), .B(n10317), .ZN(
        n10342) );
  MUX2_X1 U11380 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n10342), .S(n10499), .Z(
        P1_U3533) );
  MUX2_X1 U11381 ( .A(n10320), .B(P1_REG1_REG_0__SCAN_IN), .S(n10496), .Z(
        P1_U3523) );
  MUX2_X1 U11382 ( .A(n10321), .B(P1_REG0_REG_31__SCAN_IN), .S(n10486), .Z(
        P1_U3522) );
  MUX2_X1 U11383 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n10322), .S(n10488), .Z(
        P1_U3521) );
  MUX2_X1 U11384 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n10324), .S(n10488), .Z(
        P1_U3519) );
  MUX2_X1 U11385 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10325), .S(n10488), .Z(
        P1_U3518) );
  MUX2_X1 U11386 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10326), .S(n10488), .Z(
        P1_U3517) );
  MUX2_X1 U11387 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10327), .S(n10488), .Z(
        P1_U3516) );
  MUX2_X1 U11388 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10328), .S(n10488), .Z(
        P1_U3515) );
  MUX2_X1 U11389 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10329), .S(n10488), .Z(
        P1_U3514) );
  MUX2_X1 U11390 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10330), .S(n10488), .Z(
        P1_U3513) );
  MUX2_X1 U11391 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10331), .S(n10488), .Z(
        P1_U3512) );
  MUX2_X1 U11392 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10332), .S(n10488), .Z(
        P1_U3511) );
  MUX2_X1 U11393 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10333), .S(n10488), .Z(
        P1_U3510) );
  MUX2_X1 U11394 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10334), .S(n10488), .Z(
        P1_U3508) );
  MUX2_X1 U11395 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10335), .S(n10488), .Z(
        P1_U3505) );
  MUX2_X1 U11396 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10336), .S(n10488), .Z(
        P1_U3502) );
  MUX2_X1 U11397 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n10337), .S(n10488), .Z(
        P1_U3499) );
  MUX2_X1 U11398 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10338), .S(n10488), .Z(
        P1_U3496) );
  MUX2_X1 U11399 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n10339), .S(n10488), .Z(
        P1_U3493) );
  MUX2_X1 U11400 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n10340), .S(n10488), .Z(
        P1_U3490) );
  MUX2_X1 U11401 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n10341), .S(n10488), .Z(
        P1_U3487) );
  MUX2_X1 U11402 ( .A(P1_REG0_REG_10__SCAN_IN), .B(n10342), .S(n10488), .Z(
        P1_U3484) );
  NOR4_X1 U11403 ( .A1(n10344), .A2(P1_IR_REG_30__SCAN_IN), .A3(n10343), .A4(
        P1_U3084), .ZN(n10345) );
  AOI21_X1 U11404 ( .B1(n10349), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n10345), 
        .ZN(n10346) );
  OAI21_X1 U11405 ( .B1(n10347), .B2(n8004), .A(n10346), .ZN(P1_U3322) );
  AOI21_X1 U11406 ( .B1(n10349), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n10348), 
        .ZN(n10350) );
  OAI21_X1 U11407 ( .B1(n10351), .B2(n8004), .A(n10350), .ZN(P1_U3326) );
  OAI222_X1 U11408 ( .A1(P1_U3084), .A2(n6132), .B1(n8004), .B2(n10353), .C1(
        n10352), .C2(n8008), .ZN(P1_U3327) );
  MUX2_X1 U11409 ( .A(n10354), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  INV_X1 U11410 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n10359) );
  NAND2_X1 U11411 ( .A1(n10418), .A2(n10355), .ZN(n10358) );
  INV_X1 U11412 ( .A(n10356), .ZN(n10357) );
  OAI211_X1 U11413 ( .C1(n10411), .C2(n10359), .A(n10358), .B(n10357), .ZN(
        n10360) );
  INV_X1 U11414 ( .A(n10360), .ZN(n10369) );
  OAI211_X1 U11415 ( .C1(n10363), .C2(n10362), .A(n10425), .B(n10361), .ZN(
        n10368) );
  OAI211_X1 U11416 ( .C1(n10366), .C2(n10365), .A(n10416), .B(n10364), .ZN(
        n10367) );
  NAND3_X1 U11417 ( .A1(n10369), .A2(n10368), .A3(n10367), .ZN(P1_U3244) );
  NOR2_X1 U11418 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(P2_ADDR_REG_17__SCAN_IN), 
        .ZN(n10370) );
  AOI21_X1 U11419 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10370), .ZN(n10552) );
  NOR2_X1 U11420 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(P2_ADDR_REG_16__SCAN_IN), 
        .ZN(n10371) );
  AOI21_X1 U11421 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10371), .ZN(n10555) );
  NOR2_X1 U11422 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10372) );
  AOI21_X1 U11423 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n10372), .ZN(n10558) );
  NOR2_X1 U11424 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10373) );
  AOI21_X1 U11425 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n10373), .ZN(n10561) );
  NOR2_X1 U11426 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10374) );
  AOI21_X1 U11427 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n10374), .ZN(n10564) );
  OAI21_X1 U11428 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10375), .ZN(n10593) );
  NAND2_X1 U11429 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n10381) );
  XOR2_X1 U11430 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10591) );
  NAND2_X1 U11431 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n10380) );
  AOI21_X1 U11432 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10545) );
  INV_X1 U11433 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10378) );
  NAND3_X1 U11434 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10547) );
  OAI21_X1 U11435 ( .B1(n10545), .B2(n10378), .A(n10547), .ZN(n10589) );
  NAND2_X1 U11436 ( .A1(n4451), .A2(n10589), .ZN(n10379) );
  NAND2_X1 U11437 ( .A1(n10380), .A2(n10379), .ZN(n10590) );
  NOR2_X1 U11438 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10382), .ZN(n10578) );
  NAND2_X1 U11439 ( .A1(n10383), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n10385) );
  NAND2_X1 U11440 ( .A1(n10385), .A2(n10384), .ZN(n10386) );
  NAND2_X1 U11441 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10386), .ZN(n10387) );
  NAND2_X1 U11442 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n10388), .ZN(n10390) );
  NAND2_X1 U11443 ( .A1(n10581), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n10389) );
  NAND2_X1 U11444 ( .A1(n10390), .A2(n10389), .ZN(n10391) );
  AND2_X1 U11445 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10391), .ZN(n10392) );
  INV_X1 U11446 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10588) );
  XNOR2_X1 U11447 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n10391), .ZN(n10587) );
  NAND2_X1 U11448 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n10393) );
  OAI21_X1 U11449 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n10393), .ZN(n10572) );
  NAND2_X1 U11450 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n10394) );
  OAI21_X1 U11451 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n10394), .ZN(n10569) );
  NOR2_X1 U11452 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10395) );
  AOI21_X1 U11453 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n10395), .ZN(n10566) );
  NAND2_X1 U11454 ( .A1(n10564), .A2(n10563), .ZN(n10562) );
  NAND2_X1 U11455 ( .A1(n10561), .A2(n10560), .ZN(n10559) );
  NAND2_X1 U11456 ( .A1(n10552), .A2(n10551), .ZN(n10550) );
  NOR2_X1 U11457 ( .A1(n10584), .A2(n10583), .ZN(n10396) );
  NAND2_X1 U11458 ( .A1(n10584), .A2(n10583), .ZN(n10582) );
  OAI21_X1 U11459 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n10396), .A(n10582), 
        .ZN(n10398) );
  XOR2_X1 U11460 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .Z(n10397) );
  XNOR2_X1 U11461 ( .A(n10398), .B(n10397), .ZN(ADD_1071_U4) );
  AOI22_X1 U11462 ( .A1(P2_WR_REG_SCAN_IN), .A2(n10400), .B1(P1_WR_REG_SCAN_IN), .B2(n10399), .ZN(U123) );
  XNOR2_X1 U11463 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U11464 ( .A(n10401), .ZN(n10402) );
  OAI21_X1 U11465 ( .B1(n10403), .B2(P1_REG1_REG_0__SCAN_IN), .A(n10402), .ZN(
        n10405) );
  XNOR2_X1 U11466 ( .A(n10405), .B(n10404), .ZN(n10407) );
  OAI22_X1 U11467 ( .A1(n10408), .A2(n10407), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10406), .ZN(n10409) );
  INV_X1 U11468 ( .A(n10409), .ZN(n10410) );
  OAI21_X1 U11469 ( .B1(n10411), .B2(n10549), .A(n10410), .ZN(P1_U3241) );
  NAND2_X1 U11470 ( .A1(n10413), .A2(n10412), .ZN(n10414) );
  NAND3_X1 U11471 ( .A1(n10416), .A2(n10415), .A3(n10414), .ZN(n10421) );
  NAND2_X1 U11472 ( .A1(n10418), .A2(n10417), .ZN(n10420) );
  AND3_X1 U11473 ( .A1(n10421), .A2(n10420), .A3(n10419), .ZN(n10428) );
  XNOR2_X1 U11474 ( .A(n10423), .B(n10422), .ZN(n10424) );
  AOI22_X1 U11475 ( .A1(n10426), .A2(P1_ADDR_REG_18__SCAN_IN), .B1(n10425), 
        .B2(n10424), .ZN(n10427) );
  NAND2_X1 U11476 ( .A1(n10428), .A2(n10427), .ZN(P1_U3259) );
  AND2_X1 U11477 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10440), .ZN(P1_U3292) );
  AND2_X1 U11478 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10440), .ZN(P1_U3293) );
  AND2_X1 U11479 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10440), .ZN(P1_U3294) );
  AND2_X1 U11480 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10440), .ZN(P1_U3295) );
  AND2_X1 U11481 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10440), .ZN(P1_U3296) );
  AND2_X1 U11482 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10440), .ZN(P1_U3297) );
  AND2_X1 U11483 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10440), .ZN(P1_U3298) );
  AND2_X1 U11484 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10440), .ZN(P1_U3299) );
  AND2_X1 U11485 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10440), .ZN(P1_U3300) );
  NOR2_X1 U11486 ( .A1(n10439), .A2(n10430), .ZN(P1_U3301) );
  AND2_X1 U11487 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10440), .ZN(P1_U3302) );
  NOR2_X1 U11488 ( .A1(n10439), .A2(n10431), .ZN(P1_U3303) );
  NOR2_X1 U11489 ( .A1(n10439), .A2(n10432), .ZN(P1_U3304) );
  NOR2_X1 U11490 ( .A1(n10439), .A2(n10433), .ZN(P1_U3305) );
  NOR2_X1 U11491 ( .A1(n10439), .A2(n10434), .ZN(P1_U3306) );
  AND2_X1 U11492 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10440), .ZN(P1_U3307) );
  AND2_X1 U11493 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10440), .ZN(P1_U3308) );
  NOR2_X1 U11494 ( .A1(n10439), .A2(n10435), .ZN(P1_U3309) );
  AND2_X1 U11495 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10440), .ZN(P1_U3310) );
  AND2_X1 U11496 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10440), .ZN(P1_U3311) );
  NOR2_X1 U11497 ( .A1(n10439), .A2(n10436), .ZN(P1_U3312) );
  AND2_X1 U11498 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10440), .ZN(P1_U3313) );
  AND2_X1 U11499 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10440), .ZN(P1_U3314) );
  AND2_X1 U11500 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10440), .ZN(P1_U3315) );
  AND2_X1 U11501 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10440), .ZN(P1_U3316) );
  NOR2_X1 U11502 ( .A1(n10439), .A2(n10437), .ZN(P1_U3317) );
  AND2_X1 U11503 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10440), .ZN(P1_U3318) );
  NOR2_X1 U11504 ( .A1(n10439), .A2(n10438), .ZN(P1_U3319) );
  AND2_X1 U11505 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10440), .ZN(P1_U3320) );
  AND2_X1 U11506 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10440), .ZN(P1_U3321) );
  INV_X1 U11507 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10442) );
  OAI21_X1 U11508 ( .B1(n10443), .B2(n10442), .A(n10441), .ZN(P1_U3440) );
  NAND2_X1 U11509 ( .A1(n10444), .A2(n10485), .ZN(n10446) );
  OAI211_X1 U11510 ( .C1(n10447), .C2(n10480), .A(n10446), .B(n10445), .ZN(
        n10448) );
  NOR2_X1 U11511 ( .A1(n10449), .A2(n10448), .ZN(n10489) );
  AOI22_X1 U11512 ( .A1(n10488), .A2(n10489), .B1(n6332), .B2(n10486), .ZN(
        P1_U3457) );
  NAND2_X1 U11513 ( .A1(n10450), .A2(n10464), .ZN(n10451) );
  OAI21_X1 U11514 ( .B1(n10452), .B2(n10480), .A(n10451), .ZN(n10454) );
  AOI211_X1 U11515 ( .C1(n10485), .C2(n10455), .A(n10454), .B(n10453), .ZN(
        n10490) );
  AOI22_X1 U11516 ( .A1(n10488), .A2(n10490), .B1(n6410), .B2(n10486), .ZN(
        P1_U3460) );
  INV_X1 U11517 ( .A(n10456), .ZN(n10462) );
  OAI22_X1 U11518 ( .A1(n10459), .A2(n10458), .B1(n10457), .B2(n10480), .ZN(
        n10461) );
  AOI211_X1 U11519 ( .C1(n10485), .C2(n10462), .A(n10461), .B(n10460), .ZN(
        n10492) );
  AOI22_X1 U11520 ( .A1(n10488), .A2(n10492), .B1(n6513), .B2(n10486), .ZN(
        P1_U3466) );
  AOI22_X1 U11521 ( .A1(n10465), .A2(n10464), .B1(n10463), .B2(n4710), .ZN(
        n10466) );
  OAI211_X1 U11522 ( .C1(n10469), .C2(n10468), .A(n10467), .B(n10466), .ZN(
        n10470) );
  INV_X1 U11523 ( .A(n10470), .ZN(n10494) );
  AOI22_X1 U11524 ( .A1(n10488), .A2(n10494), .B1(n6768), .B2(n10486), .ZN(
        P1_U3472) );
  OAI211_X1 U11525 ( .C1(n10473), .C2(n10480), .A(n10472), .B(n10471), .ZN(
        n10474) );
  AOI21_X1 U11526 ( .B1(n10476), .B2(n10475), .A(n10474), .ZN(n10495) );
  AOI22_X1 U11527 ( .A1(n10488), .A2(n10495), .B1(n6792), .B2(n10486), .ZN(
        P1_U3475) );
  INV_X1 U11528 ( .A(n10477), .ZN(n10484) );
  INV_X1 U11529 ( .A(n10478), .ZN(n10479) );
  OAI21_X1 U11530 ( .B1(n10481), .B2(n10480), .A(n10479), .ZN(n10483) );
  AOI211_X1 U11531 ( .C1(n10485), .C2(n10484), .A(n10483), .B(n10482), .ZN(
        n10498) );
  INV_X1 U11532 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10487) );
  AOI22_X1 U11533 ( .A1(n10488), .A2(n10498), .B1(n10487), .B2(n10486), .ZN(
        P1_U3478) );
  AOI22_X1 U11534 ( .A1(n10499), .A2(n10489), .B1(n6333), .B2(n10496), .ZN(
        P1_U3524) );
  AOI22_X1 U11535 ( .A1(n10499), .A2(n10490), .B1(n6412), .B2(n10496), .ZN(
        P1_U3525) );
  AOI22_X1 U11536 ( .A1(n10499), .A2(n10492), .B1(n10491), .B2(n10496), .ZN(
        P1_U3527) );
  AOI22_X1 U11537 ( .A1(n10499), .A2(n10494), .B1(n10493), .B2(n10496), .ZN(
        P1_U3529) );
  AOI22_X1 U11538 ( .A1(n10499), .A2(n10495), .B1(n6789), .B2(n10496), .ZN(
        P1_U3530) );
  AOI22_X1 U11539 ( .A1(n10499), .A2(n10498), .B1(n10497), .B2(n10496), .ZN(
        P1_U3531) );
  AND2_X1 U11540 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10511), .ZN(P2_U3297) );
  AND2_X1 U11541 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10511), .ZN(P2_U3298) );
  AND2_X1 U11542 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10511), .ZN(P2_U3299) );
  AND2_X1 U11543 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10511), .ZN(P2_U3300) );
  AND2_X1 U11544 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10511), .ZN(P2_U3301) );
  AND2_X1 U11545 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10511), .ZN(P2_U3302) );
  AND2_X1 U11546 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10511), .ZN(P2_U3303) );
  NOR2_X1 U11547 ( .A1(n10508), .A2(n10502), .ZN(P2_U3304) );
  AND2_X1 U11548 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10511), .ZN(P2_U3305) );
  AND2_X1 U11549 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10511), .ZN(P2_U3306) );
  AND2_X1 U11550 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10511), .ZN(P2_U3307) );
  AND2_X1 U11551 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10511), .ZN(P2_U3308) );
  AND2_X1 U11552 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10511), .ZN(P2_U3309) );
  AND2_X1 U11553 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10511), .ZN(P2_U3310) );
  AND2_X1 U11554 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10511), .ZN(P2_U3311) );
  NOR2_X1 U11555 ( .A1(n10508), .A2(n10503), .ZN(P2_U3312) );
  AND2_X1 U11556 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10511), .ZN(P2_U3313) );
  AND2_X1 U11557 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10511), .ZN(P2_U3314) );
  NOR2_X1 U11558 ( .A1(n10508), .A2(n10504), .ZN(P2_U3315) );
  NOR2_X1 U11559 ( .A1(n10508), .A2(n10505), .ZN(P2_U3316) );
  AND2_X1 U11560 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10511), .ZN(P2_U3317) );
  NOR2_X1 U11561 ( .A1(n10508), .A2(n10506), .ZN(P2_U3318) );
  AND2_X1 U11562 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10511), .ZN(P2_U3319) );
  AND2_X1 U11563 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10511), .ZN(P2_U3320) );
  AND2_X1 U11564 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10511), .ZN(P2_U3321) );
  AND2_X1 U11565 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10511), .ZN(P2_U3322) );
  AND2_X1 U11566 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10511), .ZN(P2_U3323) );
  NOR2_X1 U11567 ( .A1(n10508), .A2(n10507), .ZN(P2_U3324) );
  AND2_X1 U11568 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10511), .ZN(P2_U3325) );
  AND2_X1 U11569 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10511), .ZN(P2_U3326) );
  AOI22_X1 U11570 ( .A1(n10514), .A2(n10510), .B1(n10509), .B2(n10511), .ZN(
        P2_U3437) );
  AOI22_X1 U11571 ( .A1(n10514), .A2(n10513), .B1(n10512), .B2(n10511), .ZN(
        P2_U3438) );
  INV_X1 U11572 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10515) );
  AOI22_X1 U11573 ( .A1(n10538), .A2(n10516), .B1(n10515), .B2(n10537), .ZN(
        P2_U3451) );
  OAI21_X1 U11574 ( .B1(n10518), .B2(n10528), .A(n10517), .ZN(n10520) );
  AOI211_X1 U11575 ( .C1(n10536), .C2(n10521), .A(n10520), .B(n10519), .ZN(
        n10539) );
  AOI22_X1 U11576 ( .A1(n10538), .A2(n10539), .B1(n10522), .B2(n10537), .ZN(
        P2_U3457) );
  OAI22_X1 U11577 ( .A1(n10524), .A2(n10530), .B1(n10523), .B2(n10528), .ZN(
        n10526) );
  AOI211_X1 U11578 ( .C1(n10536), .C2(n10527), .A(n10526), .B(n10525), .ZN(
        n10541) );
  AOI22_X1 U11579 ( .A1(n10538), .A2(n10541), .B1(n5570), .B2(n10537), .ZN(
        P2_U3463) );
  OAI22_X1 U11580 ( .A1(n10531), .A2(n10530), .B1(n10529), .B2(n10528), .ZN(
        n10534) );
  INV_X1 U11581 ( .A(n10532), .ZN(n10533) );
  AOI211_X1 U11582 ( .C1(n10536), .C2(n10535), .A(n10534), .B(n10533), .ZN(
        n10543) );
  AOI22_X1 U11583 ( .A1(n10538), .A2(n10543), .B1(n5608), .B2(n10537), .ZN(
        P2_U3469) );
  AOI22_X1 U11584 ( .A1(n10544), .A2(n10539), .B1(n5525), .B2(n10542), .ZN(
        P2_U3522) );
  AOI22_X1 U11585 ( .A1(n10544), .A2(n10541), .B1(n10540), .B2(n10542), .ZN(
        P2_U3524) );
  AOI22_X1 U11586 ( .A1(n10544), .A2(n10543), .B1(n6826), .B2(n10542), .ZN(
        P2_U3526) );
  INV_X1 U11587 ( .A(n10545), .ZN(n10546) );
  NAND2_X1 U11588 ( .A1(n10547), .A2(n10546), .ZN(n10548) );
  XNOR2_X1 U11589 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10548), .ZN(ADD_1071_U5)
         );
  AOI22_X1 U11590 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .B1(n10549), .B2(n6976), .ZN(ADD_1071_U46) );
  OAI21_X1 U11591 ( .B1(n10552), .B2(n10551), .A(n10550), .ZN(ADD_1071_U56) );
  OAI21_X1 U11592 ( .B1(n10555), .B2(n10554), .A(n10553), .ZN(ADD_1071_U57) );
  OAI21_X1 U11593 ( .B1(n10558), .B2(n10557), .A(n10556), .ZN(ADD_1071_U58) );
  OAI21_X1 U11594 ( .B1(n10561), .B2(n10560), .A(n10559), .ZN(ADD_1071_U59) );
  OAI21_X1 U11595 ( .B1(n10564), .B2(n10563), .A(n10562), .ZN(ADD_1071_U60) );
  OAI21_X1 U11596 ( .B1(n10567), .B2(n10566), .A(n10565), .ZN(ADD_1071_U61) );
  AOI21_X1 U11597 ( .B1(n10570), .B2(n10569), .A(n10568), .ZN(ADD_1071_U62) );
  AOI21_X1 U11598 ( .B1(n10573), .B2(n10572), .A(n10571), .ZN(ADD_1071_U63) );
  XNOR2_X1 U11599 ( .A(n10575), .B(n10574), .ZN(ADD_1071_U49) );
  XNOR2_X1 U11600 ( .A(n10577), .B(n10576), .ZN(ADD_1071_U50) );
  NOR2_X1 U11601 ( .A1(n10579), .A2(n10578), .ZN(n10580) );
  XNOR2_X1 U11602 ( .A(n10580), .B(n6266), .ZN(ADD_1071_U51) );
  XOR2_X1 U11603 ( .A(n10581), .B(P2_ADDR_REG_8__SCAN_IN), .Z(ADD_1071_U48) );
  OAI21_X1 U11604 ( .B1(n10584), .B2(n10583), .A(n10582), .ZN(n10585) );
  XNOR2_X1 U11605 ( .A(n10585), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11606 ( .B1(n10588), .B2(n10587), .A(n10586), .ZN(ADD_1071_U47) );
  XOR2_X1 U11607 ( .A(n4451), .B(n10589), .Z(ADD_1071_U54) );
  XOR2_X1 U11608 ( .A(n10591), .B(n10590), .Z(ADD_1071_U53) );
  XNOR2_X1 U11609 ( .A(n10593), .B(n10592), .ZN(ADD_1071_U52) );
endmodule

