

module b22_C_AntiSAT_k_256_1 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, SUB_1596_U4, SUB_1596_U62, 
        SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, 
        SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, 
        SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, 
        SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, 
        P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, 
        P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, 
        P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, 
        P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, 
        P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, 
        P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, 
        P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, 
        P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, 
        P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, 
        P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, 
        P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, 
        P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, 
        P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, 
        P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, 
        P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, 
        P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, 
        P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, 
        P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, 
        P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, 
        P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, 
        P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, 
        P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, 
        P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, 
        P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, 
        P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, 
        P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, 
        P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, 
        P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, 
        P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, 
        P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, 
        P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, 
        P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, 
        P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, 
        P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, 
        P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, 
        P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, 
        P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, 
        P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, 
        P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, 
        P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, 
        P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, 
        P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, 
        P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, 
        P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, 
        P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, 
        P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, 
        P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, 
        P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, 
        P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, 
        P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, 
        P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, 
        P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, 
        P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, 
        P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, 
        P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, 
        P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, 
        P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, 
        P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, 
        P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, 
        P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, 
        P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, 
        P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, 
        P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, 
        P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, 
        P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, 
        P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, 
        P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, 
        P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, 
        P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, 
        P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, 
        P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, 
        P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, 
        P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, 
        P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, 
        P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, 
        P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, 
        P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, 
        P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, 
        P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, 
        P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, 
        P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, 
        P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, 
        P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, 
        P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, 
        P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, 
        P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, 
        P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, 
        P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, 
        P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, 
        P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, 
        P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127,
         keyinput128, keyinput129, keyinput130, keyinput131, keyinput132,
         keyinput133, keyinput134, keyinput135, keyinput136, keyinput137,
         keyinput138, keyinput139, keyinput140, keyinput141, keyinput142,
         keyinput143, keyinput144, keyinput145, keyinput146, keyinput147,
         keyinput148, keyinput149, keyinput150, keyinput151, keyinput152,
         keyinput153, keyinput154, keyinput155, keyinput156, keyinput157,
         keyinput158, keyinput159, keyinput160, keyinput161, keyinput162,
         keyinput163, keyinput164, keyinput165, keyinput166, keyinput167,
         keyinput168, keyinput169, keyinput170, keyinput171, keyinput172,
         keyinput173, keyinput174, keyinput175, keyinput176, keyinput177,
         keyinput178, keyinput179, keyinput180, keyinput181, keyinput182,
         keyinput183, keyinput184, keyinput185, keyinput186, keyinput187,
         keyinput188, keyinput189, keyinput190, keyinput191, keyinput192,
         keyinput193, keyinput194, keyinput195, keyinput196, keyinput197,
         keyinput198, keyinput199, keyinput200, keyinput201, keyinput202,
         keyinput203, keyinput204, keyinput205, keyinput206, keyinput207,
         keyinput208, keyinput209, keyinput210, keyinput211, keyinput212,
         keyinput213, keyinput214, keyinput215, keyinput216, keyinput217,
         keyinput218, keyinput219, keyinput220, keyinput221, keyinput222,
         keyinput223, keyinput224, keyinput225, keyinput226, keyinput227,
         keyinput228, keyinput229, keyinput230, keyinput231, keyinput232,
         keyinput233, keyinput234, keyinput235, keyinput236, keyinput237,
         keyinput238, keyinput239, keyinput240, keyinput241, keyinput242,
         keyinput243, keyinput244, keyinput245, keyinput246, keyinput247,
         keyinput248, keyinput249, keyinput250, keyinput251, keyinput252,
         keyinput253, keyinput254, keyinput255;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616;

  NAND2_X1 U7388 ( .A1(n7600), .A2(n7599), .ZN(n12536) );
  INV_X1 U7389 ( .A(n12013), .ZN(n8079) );
  CLKBUF_X2 U7390 ( .A(n12027), .Z(n6986) );
  AND4_X1 U7391 ( .A1(n8583), .A2(n8582), .A3(n8581), .A4(n8580), .ZN(n10587)
         );
  INV_X1 U7393 ( .A(n7773), .ZN(n8281) );
  NAND2_X1 U7394 ( .A1(n8065), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n7755) );
  AND2_X1 U7395 ( .A1(n8537), .A2(n8538), .ZN(n8578) );
  AND2_X1 U7396 ( .A1(n11822), .A2(n8537), .ZN(n8927) );
  CLKBUF_X1 U7397 ( .A(n9136), .Z(n9507) );
  CLKBUF_X2 U7398 ( .A(n9085), .Z(n9466) );
  NOR2_X1 U7399 ( .A1(n8724), .A2(n7379), .ZN(n7382) );
  NAND2_X1 U7401 ( .A1(n9825), .A2(n8205), .ZN(n8611) );
  CLKBUF_X3 U7402 ( .A(n8611), .Z(n11550) );
  NAND2_X1 U7403 ( .A1(n8409), .A2(n8408), .ZN(n8411) );
  INV_X1 U7404 ( .A(n9642), .ZN(n8078) );
  INV_X1 U7405 ( .A(n13407), .ZN(n10014) );
  NAND2_X1 U7406 ( .A1(n10008), .A2(n11825), .ZN(n10299) );
  INV_X1 U7407 ( .A(n10299), .ZN(n10013) );
  INV_X4 U7408 ( .A(n12220), .ZN(n12273) );
  CLKBUF_X3 U7409 ( .A(n8927), .Z(n8828) );
  AND2_X1 U7410 ( .A1(n11822), .A2(n12783), .ZN(n8565) );
  BUF_X1 U7411 ( .A(n7742), .Z(n9642) );
  INV_X1 U7412 ( .A(n7792), .ZN(n8282) );
  NOR2_X1 U7413 ( .A1(n13979), .A2(n13810), .ZN(n13792) );
  NAND2_X1 U7414 ( .A1(n8413), .A2(n8412), .ZN(n8752) );
  NAND2_X1 U7415 ( .A1(n7937), .A2(n7936), .ZN(n14329) );
  NAND2_X1 U7416 ( .A1(n7922), .A2(n7921), .ZN(n11919) );
  AND4_X1 U7417 ( .A1(n9089), .A2(n9088), .A3(n9087), .A4(n9086), .ZN(n11092)
         );
  NAND2_X1 U7418 ( .A1(n13726), .A2(n7132), .ZN(n13945) );
  NOR2_X1 U7419 ( .A1(n10298), .A2(n10008), .ZN(n10012) );
  OR2_X2 U7420 ( .A1(n8645), .A2(n8397), .ZN(n8399) );
  NAND2_X2 U7421 ( .A1(n7919), .A2(n7918), .ZN(n7932) );
  NAND2_X2 U7422 ( .A1(n7610), .A2(n7611), .ZN(n7919) );
  AOI22_X2 U7424 ( .A1(n11119), .A2(n6655), .B1(n7125), .B2(n6645), .ZN(n14531) );
  NAND2_X1 U7425 ( .A1(n10785), .A2(n15156), .ZN(n11589) );
  OAI22_X2 U7426 ( .A1(n12067), .A2(n9915), .B1(n12944), .B2(n9920), .ZN(
        n10044) );
  XNOR2_X2 U7427 ( .A(n8072), .B(n8096), .ZN(n10920) );
  AND3_X2 U7428 ( .A1(n8987), .A2(n9197), .A3(n8986), .ZN(n7688) );
  AND4_X4 U7429 ( .A1(n9037), .A2(n9036), .A3(n9035), .A4(n9034), .ZN(n10152)
         );
  NAND2_X2 U7430 ( .A1(n13540), .A2(n6919), .ZN(n13457) );
  OAI21_X2 U7431 ( .B1(n10570), .B2(n7512), .A(n7509), .ZN(n10840) );
  NAND2_X4 U7432 ( .A1(n8923), .A2(n8922), .ZN(n12670) );
  OAI211_X2 U7433 ( .C1(n11550), .C2(SI_2_), .A(n8575), .B(n8574), .ZN(n10593)
         );
  INV_X1 U7434 ( .A(n8829), .ZN(n6640) );
  NAND2_X2 U7435 ( .A1(n9908), .A2(n8564), .ZN(n11567) );
  NOR4_X2 U7436 ( .A1(n11745), .A2(n11744), .A3(n11743), .A4(n11742), .ZN(
        n11746) );
  NAND4_X4 U7437 ( .A1(n7758), .A2(n7757), .A3(n7756), .A4(n7755), .ZN(n12942)
         );
  CLKBUF_X1 U7438 ( .A(n13611), .Z(n6641) );
  XNOR2_X1 U7439 ( .A(n9030), .B(n9029), .ZN(n13611) );
  INV_X1 U7440 ( .A(n12500), .ZN(n12507) );
  NAND2_X1 U7441 ( .A1(n10547), .A2(n10546), .ZN(n10550) );
  NAND2_X1 U7442 ( .A1(n10466), .A2(n10465), .ZN(n10467) );
  AOI21_X1 U7443 ( .B1(n10439), .B2(n10438), .A(n10437), .ZN(n12257) );
  NAND2_X1 U7444 ( .A1(n7848), .A2(n7847), .ZN(n11890) );
  NAND3_X1 U7445 ( .A1(n8597), .A2(n8596), .A3(n7390), .ZN(n12406) );
  INV_X1 U7446 ( .A(n10899), .ZN(n10898) );
  AND4_X2 U7447 ( .A1(n8549), .A2(n8548), .A3(n8547), .A4(n8546), .ZN(n10586)
         );
  CLKBUF_X2 U7448 ( .A(P2_U3947), .Z(n6642) );
  INV_X1 U7449 ( .A(n10593), .ZN(n10083) );
  BUF_X2 U7450 ( .A(n8578), .Z(n8934) );
  CLKBUF_X2 U7451 ( .A(n10532), .Z(n12154) );
  CLKBUF_X2 U7452 ( .A(n9310), .Z(n6935) );
  AND2_X1 U7453 ( .A1(n8538), .A2(n12783), .ZN(n8579) );
  INV_X1 U7454 ( .A(n7792), .ZN(n8065) );
  NAND2_X1 U7455 ( .A1(n10299), .A2(n10451), .ZN(n13393) );
  NAND3_X2 U7456 ( .A1(n14038), .A2(n11331), .A3(n9992), .ZN(n10451) );
  CLKBUF_X2 U7457 ( .A(n7763), .Z(n8209) );
  OR2_X1 U7458 ( .A1(n8501), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n8503) );
  XNOR2_X1 U7459 ( .A(n9561), .B(P1_IR_REG_26__SCAN_IN), .ZN(n14038) );
  AND2_X1 U7460 ( .A1(n7606), .A2(n8478), .ZN(n7605) );
  NOR2_X2 U7461 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n8572) );
  INV_X2 U7462 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  AND2_X1 U7463 ( .A1(n11751), .A2(n11750), .ZN(n7113) );
  NAND2_X1 U7464 ( .A1(n12501), .A2(n12500), .ZN(n12499) );
  AND2_X1 U7465 ( .A1(n12516), .A2(n8933), .ZN(n12501) );
  NOR2_X1 U7466 ( .A1(n13474), .A2(n7579), .ZN(n7578) );
  OR2_X1 U7467 ( .A1(n13766), .A2(n13765), .ZN(n13764) );
  CLKBUF_X1 U7468 ( .A(n12603), .Z(n12616) );
  NAND2_X1 U7469 ( .A1(n12815), .A2(n12130), .ZN(n12132) );
  NAND2_X1 U7470 ( .A1(n12209), .A2(n6775), .ZN(n12346) );
  NOR2_X1 U7471 ( .A1(n14178), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n6918) );
  XNOR2_X1 U7472 ( .A(n13390), .B(n13389), .ZN(n13566) );
  XNOR2_X1 U7473 ( .A(n8253), .B(n8252), .ZN(n13351) );
  NAND2_X1 U7474 ( .A1(n8909), .A2(n8908), .ZN(n12675) );
  OAI21_X1 U7475 ( .B1(n8921), .B2(n8444), .A(n8445), .ZN(n8543) );
  OAI21_X1 U7476 ( .B1(n8328), .B2(n7518), .A(n7516), .ZN(n8331) );
  AOI21_X1 U7477 ( .B1(n6968), .B2(n7014), .A(n14128), .ZN(n14426) );
  NAND2_X1 U7478 ( .A1(n6863), .A2(n12321), .ZN(n12366) );
  NAND2_X1 U7479 ( .A1(n8886), .A2(n8885), .ZN(n12683) );
  AOI21_X1 U7480 ( .B1(n7150), .B2(n7155), .A(n7149), .ZN(n7148) );
  NAND2_X1 U7481 ( .A1(n12197), .A2(n12196), .ZN(n12323) );
  NAND2_X1 U7482 ( .A1(n11401), .A2(n7526), .ZN(n12113) );
  NAND2_X1 U7483 ( .A1(n6872), .A2(n12194), .ZN(n12310) );
  OAI21_X1 U7484 ( .B1(n11490), .B2(n7253), .A(n7251), .ZN(n6872) );
  OR2_X1 U7485 ( .A1(n8173), .A2(n8172), .ZN(n8187) );
  NAND2_X1 U7486 ( .A1(n13922), .A2(n11761), .ZN(n13908) );
  NAND2_X1 U7487 ( .A1(n14267), .A2(n8735), .ZN(n14255) );
  NAND2_X1 U7488 ( .A1(n8081), .A2(n8080), .ZN(n13278) );
  NAND2_X1 U7489 ( .A1(n8317), .A2(n8316), .ZN(n14310) );
  NAND2_X1 U7490 ( .A1(n10761), .A2(n10760), .ZN(n11008) );
  NOR2_X1 U7491 ( .A1(n15039), .A2(n15329), .ZN(n15038) );
  NAND2_X1 U7492 ( .A1(n7993), .A2(n7992), .ZN(n13336) );
  NAND2_X1 U7493 ( .A1(n12183), .A2(n12182), .ZN(n12181) );
  NOR2_X1 U7494 ( .A1(n12085), .A2(n7439), .ZN(n7438) );
  AND2_X1 U7495 ( .A1(n14563), .A2(n14642), .ZN(n14560) );
  OAI21_X1 U7496 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n15282), .A(n14064), .ZN(
        n14065) );
  OAI21_X1 U7497 ( .B1(n11084), .B2(n7117), .A(n7115), .ZN(n10894) );
  NAND2_X1 U7498 ( .A1(n7869), .A2(n7868), .ZN(n11895) );
  XNOR2_X1 U7499 ( .A(n10801), .B(n14993), .ZN(n14999) );
  XNOR2_X1 U7500 ( .A(n8411), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n8736) );
  INV_X1 U7501 ( .A(n10587), .ZN(n12407) );
  NAND2_X2 U7502 ( .A1(n7520), .A2(n7519), .ZN(n14891) );
  OR2_X1 U7503 ( .A1(n7790), .A2(n7789), .ZN(n11870) );
  INV_X1 U7504 ( .A(n10313), .ZN(n14574) );
  CLKBUF_X1 U7505 ( .A(n10021), .Z(n13903) );
  INV_X1 U7506 ( .A(n6672), .ZN(n10976) );
  NAND2_X2 U7507 ( .A1(n7139), .A2(n7138), .ZN(n10313) );
  OAI21_X1 U7508 ( .B1(n7787), .B2(n7788), .A(n7802), .ZN(n9603) );
  INV_X2 U7509 ( .A(n11711), .ZN(n11697) );
  NAND4_X1 U7510 ( .A1(n9062), .A2(n9061), .A3(n9060), .A4(n9059), .ZN(n13597)
         );
  NAND4_X1 U7511 ( .A1(n7741), .A2(n7740), .A3(n7739), .A4(n7738), .ZN(n12943)
         );
  INV_X2 U7512 ( .A(n11318), .ZN(n13476) );
  NAND2_X1 U7513 ( .A1(n7784), .A2(n7287), .ZN(n9608) );
  BUF_X2 U7514 ( .A(n11181), .Z(n12126) );
  INV_X1 U7515 ( .A(n13393), .ZN(n6643) );
  INV_X1 U7516 ( .A(n12783), .ZN(n8537) );
  INV_X1 U7517 ( .A(n14313), .ZN(n11181) );
  NAND2_X1 U7518 ( .A1(n7736), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7723) );
  AND2_X1 U7519 ( .A1(n9016), .A2(n11829), .ZN(n9057) );
  BUF_X2 U7520 ( .A(n7832), .Z(n12008) );
  INV_X1 U7521 ( .A(n10008), .ZN(n7399) );
  NAND2_X1 U7522 ( .A1(n8535), .A2(n12777), .ZN(n12783) );
  AND2_X1 U7523 ( .A1(n7770), .A2(n6742), .ZN(n7519) );
  XNOR2_X1 U7524 ( .A(n8500), .B(P3_IR_REG_22__SCAN_IN), .ZN(n11756) );
  INV_X1 U7525 ( .A(n7737), .ZN(n7792) );
  NAND2_X1 U7526 ( .A1(n9017), .A2(n14037), .ZN(n9491) );
  NAND2_X4 U7527 ( .A1(n9570), .A2(n13611), .ZN(n9043) );
  AND2_X2 U7528 ( .A1(n9555), .A2(n8993), .ZN(n10008) );
  AND2_X1 U7529 ( .A1(n12058), .A2(n8343), .ZN(n14883) );
  INV_X1 U7530 ( .A(n12058), .ZN(n12105) );
  NAND2_X1 U7531 ( .A1(n9013), .A2(n9014), .ZN(n14037) );
  OAI21_X1 U7532 ( .B1(n7750), .B2(n6894), .A(n7749), .ZN(n7035) );
  NAND2_X1 U7533 ( .A1(n7443), .A2(n7445), .ZN(n13348) );
  NAND2_X1 U7534 ( .A1(n8271), .A2(n8077), .ZN(n12983) );
  MUX2_X1 U7535 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9012), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n9013) );
  NAND2_X1 U7536 ( .A1(n7444), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n7443) );
  XNOR2_X1 U7537 ( .A(n8508), .B(n8507), .ZN(n10326) );
  XNOR2_X1 U7538 ( .A(n8479), .B(n8478), .ZN(n10959) );
  NOR2_X1 U7539 ( .A1(n8277), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n8360) );
  NAND2_X1 U7540 ( .A1(n7361), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9030) );
  INV_X2 U7541 ( .A(n9042), .ZN(n9371) );
  NAND2_X1 U7542 ( .A1(n7654), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7720) );
  AOI21_X1 U7543 ( .B1(n8584), .B2(n7312), .A(n7311), .ZN(n7309) );
  NAND2_X1 U7544 ( .A1(n7013), .A2(n7544), .ZN(n14076) );
  AND2_X1 U7545 ( .A1(n8386), .A2(n8385), .ZN(n8570) );
  AND3_X1 U7546 ( .A1(n7478), .A2(n7477), .A3(n7761), .ZN(n7701) );
  AND4_X1 U7547 ( .A1(n8455), .A2(n8781), .A3(n15342), .A4(n8454), .ZN(n8456)
         );
  AND3_X1 U7548 ( .A1(n8450), .A2(n8449), .A3(n8448), .ZN(n8719) );
  AND3_X1 U7549 ( .A1(n8722), .A2(n8452), .A3(n8616), .ZN(n8453) );
  NOR2_X1 U7550 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6812) );
  INV_X4 U7551 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NOR2_X1 U7552 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n7269) );
  INV_X1 U7553 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9556) );
  INV_X1 U7554 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7718) );
  INV_X1 U7555 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n12988) );
  INV_X4 U7556 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7557 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n7886) );
  NOR2_X1 U7558 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n7478) );
  NOR2_X1 U7559 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n7477) );
  INV_X1 U7560 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9006) );
  INV_X1 U7561 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8268) );
  INV_X1 U7562 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9596) );
  NOR2_X1 U7563 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n7695) );
  NOR2_X1 U7564 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n7694) );
  NOR2_X1 U7565 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n8986) );
  INV_X1 U7566 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n7933) );
  INV_X1 U7567 ( .A(n8538), .ZN(n11822) );
  NAND2_X1 U7568 ( .A1(n8997), .A2(n8996), .ZN(n11825) );
  NOR2_X2 U7569 ( .A1(n12491), .A2(n6961), .ZN(n9584) );
  OAI21_X2 U7570 ( .B1(n8955), .B2(n14264), .A(n8954), .ZN(n12491) );
  NOR2_X2 U7571 ( .A1(n8036), .A2(n7699), .ZN(n7702) );
  XNOR2_X2 U7572 ( .A(n12132), .B(n12131), .ZN(n12873) );
  OAI22_X2 U7573 ( .A1(n12582), .A2(n8866), .B1(n12568), .B2(n12747), .ZN(
        n12566) );
  OAI21_X2 U7574 ( .B1(n8843), .B2(n7596), .A(n7595), .ZN(n12582) );
  XNOR2_X2 U7575 ( .A(n7385), .B(P3_IR_REG_30__SCAN_IN), .ZN(n8538) );
  OR2_X2 U7576 ( .A1(n8536), .A2(n8598), .ZN(n7385) );
  AND2_X1 U7577 ( .A1(n10796), .A2(n7474), .ZN(n10797) );
  NAND2_X1 U7578 ( .A1(n10814), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7474) );
  NAND2_X1 U7579 ( .A1(n12603), .A2(n12605), .ZN(n8843) );
  NAND2_X1 U7580 ( .A1(n7707), .A2(n7658), .ZN(n7657) );
  INV_X1 U7581 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n7658) );
  NAND2_X1 U7582 ( .A1(n12346), .A2(n7261), .ZN(n12295) );
  NOR2_X1 U7583 ( .A1(n12298), .A2(n7262), .ZN(n7261) );
  INV_X1 U7584 ( .A(n12213), .ZN(n7262) );
  INV_X1 U7585 ( .A(n8579), .ZN(n8594) );
  OR2_X1 U7586 ( .A1(n15057), .A2(n15056), .ZN(n15054) );
  NAND2_X1 U7587 ( .A1(n6686), .A2(n7166), .ZN(n7167) );
  NAND2_X1 U7588 ( .A1(n7742), .A2(n9042), .ZN(n7769) );
  NAND2_X1 U7589 ( .A1(n13759), .A2(n6699), .ZN(n13698) );
  INV_X1 U7590 ( .A(n13941), .ZN(n7288) );
  NAND2_X1 U7591 ( .A1(n13958), .A2(n6711), .ZN(n13726) );
  INV_X1 U7592 ( .A(n9485), .ZN(n9488) );
  NAND2_X1 U7593 ( .A1(n7003), .A2(n6748), .ZN(n6835) );
  AOI22_X1 U7594 ( .A1(n12941), .A2(n12031), .B1(n11870), .B2(n12051), .ZN(
        n11871) );
  OAI21_X1 U7595 ( .B1(n11886), .B2(n12051), .A(n11885), .ZN(n11887) );
  OAI21_X1 U7596 ( .B1(n6673), .B2(n11913), .A(n11917), .ZN(n7676) );
  INV_X1 U7597 ( .A(n11935), .ZN(n7671) );
  NOR2_X1 U7598 ( .A1(n8098), .A2(n7650), .ZN(n7649) );
  INV_X1 U7599 ( .A(n8055), .ZN(n7650) );
  INV_X1 U7600 ( .A(n11559), .ZN(n11566) );
  NOR2_X1 U7601 ( .A1(n13283), .A2(n13278), .ZN(n7230) );
  NAND2_X1 U7602 ( .A1(n8004), .A2(n8003), .ZN(n13183) );
  INV_X1 U7603 ( .A(n7970), .ZN(n7634) );
  OR2_X1 U7604 ( .A1(n7260), .A2(n11747), .ZN(n6869) );
  AND2_X1 U7605 ( .A1(n7336), .A2(n7335), .ZN(n12463) );
  NAND2_X1 U7606 ( .A1(n15033), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7335) );
  OR2_X1 U7607 ( .A1(n12547), .A2(n12227), .ZN(n11689) );
  OR2_X1 U7608 ( .A1(n12343), .A2(n12210), .ZN(n11665) );
  AND3_X1 U7609 ( .A1(n8684), .A2(n8683), .A3(n8682), .ZN(n11139) );
  NAND2_X1 U7610 ( .A1(n8651), .A2(n8650), .ZN(n10945) );
  NAND2_X1 U7611 ( .A1(n8702), .A2(n8701), .ZN(n14291) );
  NAND2_X1 U7612 ( .A1(n11559), .A2(n9578), .ZN(n11747) );
  INV_X1 U7613 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8455) );
  INV_X1 U7614 ( .A(n7333), .ZN(n7332) );
  OAI21_X1 U7615 ( .B1(n8692), .B2(n7334), .A(n8406), .ZN(n7333) );
  OR2_X1 U7616 ( .A1(n8629), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n8721) );
  INV_X1 U7617 ( .A(n12806), .ZN(n7156) );
  INV_X1 U7618 ( .A(n12112), .ZN(n7165) );
  INV_X1 U7619 ( .A(n13348), .ZN(n7713) );
  AND2_X1 U7620 ( .A1(n8251), .A2(n8250), .ZN(n12095) );
  OR2_X1 U7621 ( .A1(n11910), .A2(n11909), .ZN(n11902) );
  NOR2_X1 U7622 ( .A1(n7857), .A2(n7434), .ZN(n7433) );
  INV_X1 U7623 ( .A(n7837), .ZN(n7434) );
  NOR2_X1 U7624 ( .A1(n6669), .A2(n8209), .ZN(n7620) );
  INV_X1 U7625 ( .A(n7626), .ZN(n7623) );
  NAND2_X1 U7626 ( .A1(n7625), .A2(n7627), .ZN(n7624) );
  NOR3_X1 U7627 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .A3(
        P2_IR_REG_24__SCAN_IN), .ZN(n7705) );
  INV_X1 U7628 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n7697) );
  AND2_X1 U7629 ( .A1(n13490), .A2(n7571), .ZN(n7566) );
  INV_X1 U7630 ( .A(n7130), .ZN(n7129) );
  OAI21_X1 U7631 ( .B1(n13808), .B2(n7131), .A(n11773), .ZN(n7130) );
  NAND2_X1 U7632 ( .A1(n7280), .A2(n11770), .ZN(n7279) );
  INV_X1 U7633 ( .A(n13823), .ZN(n7280) );
  AND2_X1 U7634 ( .A1(n13832), .A2(n11768), .ZN(n7281) );
  NAND2_X1 U7635 ( .A1(n6814), .A2(n11764), .ZN(n13865) );
  OR2_X1 U7636 ( .A1(n14383), .A2(n13912), .ZN(n11780) );
  NOR2_X1 U7637 ( .A1(n7682), .A2(n7189), .ZN(n7188) );
  INV_X1 U7638 ( .A(n9043), .ZN(n9310) );
  NAND2_X1 U7639 ( .A1(n8223), .A2(n8222), .ZN(n8238) );
  NAND2_X1 U7640 ( .A1(n8187), .A2(n7641), .ZN(n7643) );
  NOR2_X1 U7641 ( .A1(n8201), .A2(n7642), .ZN(n7641) );
  INV_X1 U7642 ( .A(n8186), .ZN(n7642) );
  INV_X1 U7643 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9005) );
  AND2_X1 U7644 ( .A1(n7421), .A2(n9006), .ZN(n7420) );
  INV_X1 U7645 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9004) );
  NAND2_X1 U7646 ( .A1(n9371), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6892) );
  INV_X1 U7647 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7616) );
  XNOR2_X1 U7648 ( .A(n14052), .B(P3_ADDR_REG_4__SCAN_IN), .ZN(n6862) );
  OAI21_X1 U7649 ( .B1(n7257), .B2(n10740), .A(n6865), .ZN(n12183) );
  AOI21_X1 U7650 ( .B1(n7256), .B2(n7255), .A(n6687), .ZN(n6865) );
  INV_X1 U7651 ( .A(n10739), .ZN(n7255) );
  OR2_X1 U7652 ( .A1(n10443), .A2(n10444), .ZN(n10564) );
  NAND2_X1 U7653 ( .A1(n12295), .A2(n12215), .ZN(n12218) );
  NOR2_X1 U7654 ( .A1(n11715), .A2(n11714), .ZN(n11751) );
  NAND2_X1 U7655 ( .A1(n7098), .A2(n6723), .ZN(n7097) );
  OAI21_X1 U7656 ( .B1(n11529), .B2(n7099), .A(n11557), .ZN(n7098) );
  AND2_X1 U7657 ( .A1(n10797), .A2(n14962), .ZN(n10798) );
  OR2_X1 U7658 ( .A1(n14996), .A2(n15195), .ZN(n6831) );
  NOR2_X1 U7659 ( .A1(n15009), .A2(n7061), .ZN(n12412) );
  NOR2_X1 U7660 ( .A1(n15015), .A2(n10803), .ZN(n7061) );
  NAND2_X1 U7661 ( .A1(n12649), .A2(n6776), .ZN(n12630) );
  INV_X1 U7662 ( .A(n7088), .ZN(n7087) );
  OAI21_X1 U7663 ( .B1(n7089), .B2(n11630), .A(n11642), .ZN(n7088) );
  AND2_X1 U7664 ( .A1(n9579), .A2(n11558), .ZN(n14264) );
  INV_X1 U7665 ( .A(n11756), .ZN(n8975) );
  INV_X1 U7666 ( .A(n11550), .ZN(n8823) );
  INV_X2 U7667 ( .A(n8679), .ZN(n11549) );
  INV_X1 U7668 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8452) );
  AND2_X1 U7669 ( .A1(n8403), .A2(n8402), .ZN(n8675) );
  AOI21_X1 U7670 ( .B1(n8662), .B2(n7307), .A(n7306), .ZN(n7305) );
  INV_X1 U7671 ( .A(n8401), .ZN(n7306) );
  INV_X1 U7672 ( .A(n8398), .ZN(n7307) );
  INV_X1 U7673 ( .A(n8662), .ZN(n7308) );
  INV_X1 U7674 ( .A(n7322), .ZN(n7321) );
  OAI21_X1 U7675 ( .B1(n7323), .B2(n8393), .A(n8395), .ZN(n7322) );
  AND2_X1 U7676 ( .A1(n11402), .A2(n11400), .ZN(n7526) );
  NAND2_X1 U7677 ( .A1(n12120), .A2(n7158), .ZN(n7157) );
  INV_X1 U7678 ( .A(n12121), .ZN(n7158) );
  INV_X1 U7679 ( .A(n12921), .ZN(n12827) );
  NAND2_X1 U7680 ( .A1(n7505), .A2(n7504), .ZN(n7503) );
  INV_X1 U7681 ( .A(n12842), .ZN(n7504) );
  NAND2_X1 U7682 ( .A1(n7742), .A2(n8205), .ZN(n7763) );
  NAND2_X1 U7683 ( .A1(n12834), .A2(n6656), .ZN(n7502) );
  AND2_X1 U7684 ( .A1(n7713), .A2(n13346), .ZN(n7736) );
  AND2_X1 U7685 ( .A1(n13348), .A2(n7712), .ZN(n7832) );
  AND2_X1 U7686 ( .A1(n13346), .A2(n13348), .ZN(n7737) );
  NAND2_X1 U7687 ( .A1(n7426), .A2(n7424), .ZN(n13090) );
  NOR2_X1 U7688 ( .A1(n13094), .A2(n7425), .ZN(n7424) );
  INV_X1 U7689 ( .A(n7427), .ZN(n7425) );
  NAND2_X1 U7690 ( .A1(n13158), .A2(n8324), .ZN(n13137) );
  NAND2_X1 U7691 ( .A1(n13165), .A2(n8322), .ZN(n7508) );
  NAND2_X1 U7692 ( .A1(n13169), .A2(n8050), .ZN(n13148) );
  OR2_X1 U7693 ( .A1(n7036), .A2(n11103), .ZN(n7037) );
  INV_X1 U7694 ( .A(n7438), .ZN(n7036) );
  AOI21_X1 U7695 ( .B1(n7438), .B2(n12082), .A(n6685), .ZN(n7038) );
  NOR2_X1 U7696 ( .A1(n8314), .A2(n7495), .ZN(n7494) );
  NOR2_X1 U7697 ( .A1(n11910), .A2(n12935), .ZN(n7495) );
  CLKBUF_X1 U7698 ( .A(n11181), .Z(n13049) );
  INV_X1 U7699 ( .A(n14304), .ZN(n13171) );
  NAND2_X1 U7700 ( .A1(n6905), .A2(n12014), .ZN(n13224) );
  CLKBUF_X2 U7701 ( .A(n7769), .Z(n12013) );
  XNOR2_X1 U7702 ( .A(n7711), .B(P2_IR_REG_30__SCAN_IN), .ZN(n7712) );
  OR2_X1 U7703 ( .A1(n7710), .A2(n8268), .ZN(n7711) );
  NOR2_X1 U7704 ( .A1(n7577), .A2(n7574), .ZN(n7573) );
  INV_X1 U7705 ( .A(n13499), .ZN(n7574) );
  INV_X1 U7706 ( .A(n7578), .ZN(n7577) );
  AND2_X1 U7707 ( .A1(n11829), .A2(n14037), .ZN(n9085) );
  NAND2_X1 U7708 ( .A1(n11235), .A2(n11234), .ZN(n11315) );
  CLKBUF_X3 U7709 ( .A(n9057), .Z(n9492) );
  NAND2_X1 U7710 ( .A1(n6815), .A2(n11774), .ZN(n13766) );
  NAND2_X1 U7711 ( .A1(n13769), .A2(n13772), .ZN(n6815) );
  OR2_X1 U7712 ( .A1(n13973), .A2(n13789), .ZN(n11793) );
  AOI21_X1 U7713 ( .B1(n13923), .B2(n7357), .A(n6653), .ZN(n7178) );
  OR2_X1 U7714 ( .A1(n14375), .A2(n13899), .ZN(n11782) );
  NAND2_X1 U7715 ( .A1(n7267), .A2(n11200), .ZN(n11258) );
  NAND2_X1 U7716 ( .A1(n14531), .A2(n14534), .ZN(n7267) );
  NAND2_X1 U7717 ( .A1(n9472), .A2(n9471), .ZN(n13941) );
  NAND2_X1 U7718 ( .A1(n10309), .A2(n10308), .ZN(n14554) );
  NOR2_X1 U7719 ( .A1(n9506), .A2(n6786), .ZN(n7626) );
  OAI21_X1 U7720 ( .B1(n8253), .B2(n6790), .A(n6887), .ZN(n9504) );
  AOI21_X1 U7721 ( .B1(n9482), .B2(n6888), .A(n6802), .ZN(n6887) );
  XNOR2_X1 U7722 ( .A(n9015), .B(P1_IR_REG_30__SCAN_IN), .ZN(n9017) );
  NAND2_X1 U7723 ( .A1(n9014), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9015) );
  AND2_X1 U7724 ( .A1(n7589), .A2(n7283), .ZN(n7282) );
  INV_X1 U7725 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n7283) );
  NAND3_X1 U7726 ( .A1(n8204), .A2(n8222), .A3(n6897), .ZN(n8223) );
  INV_X1 U7727 ( .A(n8206), .ZN(n6897) );
  AOI21_X1 U7728 ( .B1(n7612), .B2(n7882), .A(n7903), .ZN(n7611) );
  AND2_X1 U7729 ( .A1(n7546), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n14078) );
  OAI21_X1 U7730 ( .B1(n14106), .B2(n15462), .A(n14147), .ZN(n14107) );
  NAND2_X1 U7731 ( .A1(n14409), .A2(n6867), .ZN(n14116) );
  NAND2_X1 U7732 ( .A1(n6868), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n6867) );
  OR2_X1 U7733 ( .A1(n14425), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n7016) );
  NAND2_X1 U7734 ( .A1(n15054), .A2(n6787), .ZN(n7457) );
  AND2_X1 U7735 ( .A1(n12506), .A2(n12505), .ZN(n12667) );
  AOI21_X1 U7736 ( .B1(n8294), .B2(n14304), .A(n8293), .ZN(n11841) );
  INV_X1 U7737 ( .A(n13995), .ZN(n13536) );
  NOR2_X1 U7738 ( .A1(n13714), .A2(n7133), .ZN(n7132) );
  INV_X1 U7739 ( .A(n11778), .ZN(n7133) );
  OAI21_X1 U7740 ( .B1(n9499), .B2(n10302), .A(n9033), .ZN(n9069) );
  NAND2_X1 U7741 ( .A1(n9499), .A2(n9032), .ZN(n9033) );
  OAI22_X1 U7742 ( .A1(n11862), .A2(n11863), .B1(n11860), .B2(n11861), .ZN(
        n11867) );
  OR2_X1 U7743 ( .A1(n7003), .A2(n6748), .ZN(n6837) );
  OAI21_X1 U7744 ( .B1(n11873), .B2(n7663), .A(n7001), .ZN(n11880) );
  NAND2_X1 U7745 ( .A1(n11887), .A2(n6701), .ZN(n7673) );
  INV_X1 U7746 ( .A(n11575), .ZN(n6983) );
  AND2_X1 U7747 ( .A1(n11572), .A2(n11573), .ZN(n6984) );
  NAND2_X1 U7748 ( .A1(n6681), .A2(n7671), .ZN(n7670) );
  NOR3_X1 U7749 ( .A1(n11614), .A2(n11613), .A3(n11612), .ZN(n11624) );
  NAND2_X1 U7750 ( .A1(n7006), .A2(n7005), .ZN(n7004) );
  INV_X1 U7751 ( .A(n11951), .ZN(n7005) );
  INV_X1 U7752 ( .A(n11952), .ZN(n7006) );
  OR2_X1 U7753 ( .A1(n9363), .A2(n7412), .ZN(n7411) );
  INV_X1 U7754 ( .A(n9362), .ZN(n7412) );
  OAI21_X1 U7755 ( .B1(n11640), .B2(n11639), .A(n11641), .ZN(n11647) );
  INV_X1 U7756 ( .A(n6840), .ZN(n6839) );
  OAI21_X1 U7757 ( .B1(n7674), .B2(n6696), .A(n11978), .ZN(n6840) );
  NAND2_X1 U7758 ( .A1(n6969), .A2(n6838), .ZN(n6841) );
  AND2_X1 U7759 ( .A1(n7674), .A2(n6696), .ZN(n6838) );
  AOI21_X1 U7760 ( .B1(n11679), .B2(n12687), .A(n11678), .ZN(n11687) );
  OR2_X1 U7761 ( .A1(n10298), .A2(n10878), .ZN(n9003) );
  INV_X1 U7762 ( .A(n8051), .ZN(n7647) );
  NAND2_X1 U7763 ( .A1(n12408), .A2(n10593), .ZN(n11573) );
  NAND2_X1 U7764 ( .A1(n8462), .A2(n7380), .ZN(n7379) );
  INV_X1 U7765 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8462) );
  INV_X1 U7766 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n7380) );
  NAND2_X1 U7767 ( .A1(n6736), .A2(n7660), .ZN(n7659) );
  NAND2_X1 U7768 ( .A1(n13045), .A2(n8334), .ZN(n7531) );
  INV_X1 U7769 ( .A(n8334), .ZN(n7528) );
  AND2_X1 U7770 ( .A1(n11766), .A2(n11765), .ZN(n11784) );
  AOI21_X1 U7771 ( .B1(n7931), .B2(n7930), .A(n7640), .ZN(n7639) );
  INV_X1 U7772 ( .A(n7949), .ZN(n7640) );
  OR2_X1 U7773 ( .A1(n12372), .A2(n7249), .ZN(n7248) );
  OAI211_X1 U7774 ( .C1(n9825), .C2(n9836), .A(n8555), .B(n8554), .ZN(n10028)
         );
  OR2_X1 U7775 ( .A1(n8679), .A2(n9591), .ZN(n8554) );
  OR2_X1 U7776 ( .A1(n12722), .A2(n12486), .ZN(n11713) );
  AND2_X1 U7777 ( .A1(n8496), .A2(n8480), .ZN(n9589) );
  NAND2_X1 U7778 ( .A1(n9854), .A2(n6722), .ZN(n7337) );
  NAND2_X1 U7779 ( .A1(n6817), .A2(n6816), .ZN(n12469) );
  AOI21_X1 U7780 ( .B1(n12465), .B2(n6818), .A(n6796), .ZN(n6816) );
  NAND2_X1 U7781 ( .A1(n15042), .A2(n6818), .ZN(n6817) );
  OR2_X1 U7782 ( .A1(n12513), .A2(n12231), .ZN(n11700) );
  INV_X1 U7783 ( .A(n7111), .ZN(n7106) );
  OR2_X1 U7784 ( .A1(n12596), .A2(n12354), .ZN(n11669) );
  OR2_X1 U7785 ( .A1(n12759), .A2(n12392), .ZN(n11660) );
  OR2_X1 U7786 ( .A1(n8760), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8772) );
  NAND2_X1 U7787 ( .A1(n10507), .A2(n11729), .ZN(n7594) );
  NAND2_X1 U7788 ( .A1(n11585), .A2(n11586), .ZN(n8622) );
  AND3_X1 U7789 ( .A1(n8621), .A2(n8620), .A3(n8619), .ZN(n10559) );
  NAND2_X1 U7790 ( .A1(n10586), .A2(n10028), .ZN(n11570) );
  NAND2_X1 U7791 ( .A1(n11567), .A2(n11570), .ZN(n15115) );
  XNOR2_X1 U7792 ( .A(n12406), .B(n15147), .ZN(n11729) );
  NAND2_X1 U7793 ( .A1(n8482), .A2(n8496), .ZN(n8494) );
  INV_X1 U7794 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8467) );
  INV_X1 U7795 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7381) );
  INV_X1 U7796 ( .A(n7379), .ZN(n7378) );
  INV_X1 U7797 ( .A(n8405), .ZN(n7334) );
  INV_X1 U7798 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8616) );
  INV_X1 U7799 ( .A(n8386), .ZN(n7312) );
  NAND2_X1 U7800 ( .A1(n10195), .A2(n7172), .ZN(n10532) );
  NAND2_X1 U7801 ( .A1(n12105), .A2(n12983), .ZN(n7172) );
  AOI21_X1 U7802 ( .B1(n7436), .B2(n8336), .A(n7025), .ZN(n7031) );
  INV_X1 U7803 ( .A(n8251), .ZN(n7025) );
  INV_X1 U7804 ( .A(n8329), .ZN(n7518) );
  OAI21_X1 U7805 ( .B1(n6679), .B2(n7518), .A(n13074), .ZN(n7517) );
  NOR2_X1 U7806 ( .A1(n13183), .A2(n13198), .ZN(n7053) );
  NAND2_X1 U7807 ( .A1(n7909), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7941) );
  INV_X1 U7808 ( .A(n8310), .ZN(n7513) );
  OAI22_X1 U7809 ( .A1(n14301), .A2(n7985), .B1(n7984), .B2(n14308), .ZN(
        n13203) );
  XNOR2_X1 U7810 ( .A(n7213), .B(P2_IR_REG_28__SCAN_IN), .ZN(n8286) );
  AOI21_X1 U7811 ( .B1(n7720), .B2(n7721), .A(n8268), .ZN(n7213) );
  NAND4_X1 U7812 ( .A1(n8075), .A2(n7704), .A3(n8269), .A4(n7703), .ZN(n8272)
         );
  INV_X1 U7813 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n7704) );
  NAND2_X1 U7814 ( .A1(n13413), .A2(n13414), .ZN(n7557) );
  INV_X1 U7815 ( .A(n9491), .ZN(n9058) );
  OAI22_X1 U7816 ( .A1(n10144), .A2(n13407), .B1(n14574), .B2(n13393), .ZN(
        n10146) );
  NAND2_X1 U7817 ( .A1(n14342), .A2(n13387), .ZN(n13390) );
  NOR2_X1 U7818 ( .A1(n13943), .A2(n7290), .ZN(n7289) );
  INV_X1 U7819 ( .A(n11772), .ZN(n7131) );
  INV_X1 U7820 ( .A(n7355), .ZN(n7197) );
  AND2_X1 U7821 ( .A1(n13850), .A2(n11785), .ZN(n7198) );
  NOR2_X1 U7822 ( .A1(n14383), .A2(n14169), .ZN(n7295) );
  INV_X1 U7823 ( .A(n7122), .ZN(n7121) );
  OAI21_X1 U7824 ( .B1(n7189), .B2(n7123), .A(n11353), .ZN(n7122) );
  INV_X1 U7825 ( .A(n11259), .ZN(n7123) );
  NAND2_X1 U7826 ( .A1(n10867), .A2(n10889), .ZN(n10868) );
  NOR2_X1 U7827 ( .A1(n10888), .A2(n11072), .ZN(n7116) );
  XNOR2_X1 U7828 ( .A(n13597), .B(n11088), .ZN(n11090) );
  NAND2_X1 U7829 ( .A1(n10865), .A2(n10864), .ZN(n11091) );
  NAND2_X1 U7830 ( .A1(n7174), .A2(n7175), .ZN(n13868) );
  AOI21_X1 U7831 ( .B1(n6644), .B2(n7179), .A(n6658), .ZN(n7175) );
  INV_X1 U7832 ( .A(n11784), .ZN(n13867) );
  INV_X1 U7833 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9010) );
  NAND2_X1 U7834 ( .A1(n6883), .A2(n8155), .ZN(n8157) );
  NOR2_X1 U7835 ( .A1(n8153), .A2(n6885), .ZN(n6884) );
  NAND2_X1 U7836 ( .A1(n8122), .A2(SI_21_), .ZN(n8138) );
  AOI21_X1 U7837 ( .B1(n7645), .B2(n7648), .A(n6783), .ZN(n7644) );
  NAND2_X1 U7838 ( .A1(n8103), .A2(n8104), .ZN(n6896) );
  INV_X1 U7839 ( .A(n8105), .ZN(n8104) );
  OR2_X1 U7840 ( .A1(n8099), .A2(n15288), .ZN(n8070) );
  NAND2_X1 U7841 ( .A1(n6880), .A2(n6878), .ZN(n8031) );
  AND2_X1 U7842 ( .A1(n6879), .A2(n8012), .ZN(n6878) );
  NAND2_X1 U7843 ( .A1(n6674), .A2(n6882), .ZN(n6879) );
  AOI21_X1 U7844 ( .B1(n7883), .B2(n7614), .A(n7613), .ZN(n7612) );
  INV_X1 U7845 ( .A(n7879), .ZN(n7614) );
  INV_X1 U7846 ( .A(n7900), .ZN(n7613) );
  NAND2_X1 U7847 ( .A1(n7787), .A2(n6936), .ZN(n7608) );
  OAI21_X1 U7848 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n15040), .A(n14069), .ZN(
        n14113) );
  OAI21_X1 U7849 ( .B1(n7239), .B2(n7238), .A(n6738), .ZN(n7236) );
  NAND2_X1 U7850 ( .A1(n8524), .A2(n15313), .ZN(n8861) );
  OR2_X1 U7851 ( .A1(n11489), .A2(n7253), .ZN(n7252) );
  INV_X1 U7852 ( .A(n11493), .ZN(n7253) );
  OR2_X1 U7853 ( .A1(n11150), .A2(n11151), .ZN(n11339) );
  NOR2_X1 U7854 ( .A1(n12411), .A2(n10056), .ZN(n15113) );
  NAND2_X1 U7855 ( .A1(n6908), .A2(n6907), .ZN(n10081) );
  NAND2_X1 U7856 ( .A1(n10588), .A2(n12220), .ZN(n6907) );
  NAND2_X1 U7857 ( .A1(n12273), .A2(n11570), .ZN(n6908) );
  AOI21_X2 U7858 ( .B1(n12353), .B2(n12568), .A(n12219), .ZN(n12333) );
  OR2_X1 U7859 ( .A1(n12773), .A2(n9589), .ZN(n11755) );
  AND3_X1 U7860 ( .A1(n8842), .A2(n8841), .A3(n8840), .ZN(n12210) );
  AND4_X1 U7861 ( .A1(n8818), .A2(n8817), .A3(n8816), .A4(n8815), .ZN(n12324)
         );
  AND4_X1 U7862 ( .A1(n8804), .A2(n8803), .A3(n8802), .A4(n8801), .ZN(n12199)
         );
  AND4_X1 U7863 ( .A1(n8777), .A2(n8776), .A3(n8775), .A4(n8774), .ZN(n12192)
         );
  AND4_X1 U7864 ( .A1(n8658), .A2(n8657), .A3(n8656), .A4(n8655), .ZN(n11146)
         );
  OAI21_X1 U7865 ( .B1(n8594), .B2(n7392), .A(n8595), .ZN(n7391) );
  NAND2_X1 U7866 ( .A1(n9973), .A2(n6930), .ZN(n14948) );
  OR2_X1 U7867 ( .A1(n7337), .A2(n9983), .ZN(n6930) );
  NOR2_X1 U7868 ( .A1(n14948), .A2(n15566), .ZN(n14947) );
  OR2_X1 U7869 ( .A1(n10806), .A2(n14962), .ZN(n6823) );
  NOR2_X1 U7870 ( .A1(n10800), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7471) );
  AND2_X1 U7871 ( .A1(n7473), .A2(n7063), .ZN(n10801) );
  NAND2_X1 U7872 ( .A1(n10812), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7063) );
  NAND2_X1 U7873 ( .A1(n7062), .A2(n7461), .ZN(n15009) );
  NAND2_X1 U7874 ( .A1(n10802), .A2(n7465), .ZN(n7461) );
  OR2_X1 U7875 ( .A1(n14999), .A2(n7462), .ZN(n7062) );
  NAND2_X1 U7876 ( .A1(n7465), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7462) );
  OR2_X1 U7877 ( .A1(n14999), .A2(n15000), .ZN(n7464) );
  NAND2_X1 U7878 ( .A1(n6831), .A2(n6675), .ZN(n7341) );
  NAND2_X1 U7879 ( .A1(n7341), .A2(n7340), .ZN(n7339) );
  INV_X1 U7880 ( .A(n15007), .ZN(n7340) );
  NAND2_X1 U7881 ( .A1(n7453), .A2(n7451), .ZN(n7070) );
  INV_X1 U7882 ( .A(n7452), .ZN(n7451) );
  OAI21_X1 U7883 ( .B1(n12414), .B2(P3_REG2_REG_9__SCAN_IN), .A(n7456), .ZN(
        n7452) );
  XNOR2_X1 U7884 ( .A(n12463), .B(n12464), .ZN(n15043) );
  NOR2_X1 U7885 ( .A1(n15043), .A2(n15044), .ZN(n15042) );
  NAND2_X1 U7886 ( .A1(n7070), .A2(n7069), .ZN(n7068) );
  NAND2_X1 U7887 ( .A1(n15033), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7069) );
  INV_X1 U7888 ( .A(n15041), .ZN(n12464) );
  OR2_X1 U7889 ( .A1(n15077), .A2(n15078), .ZN(n6997) );
  XNOR2_X1 U7890 ( .A(n12469), .B(n12468), .ZN(n15077) );
  NOR2_X1 U7891 ( .A1(n14203), .A2(n14202), .ZN(n14201) );
  NOR2_X1 U7892 ( .A1(n14201), .A2(n6980), .ZN(n14217) );
  AND2_X1 U7893 ( .A1(n12444), .A2(n14198), .ZN(n6980) );
  NOR2_X1 U7894 ( .A1(n14226), .A2(n12479), .ZN(n14246) );
  OAI21_X1 U7895 ( .B1(n14224), .B2(n7469), .A(n7468), .ZN(n14240) );
  NAND2_X1 U7896 ( .A1(n7470), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n7469) );
  NAND2_X1 U7897 ( .A1(n12424), .A2(n7470), .ZN(n7468) );
  INV_X1 U7898 ( .A(n14241), .ZN(n7470) );
  NOR2_X1 U7899 ( .A1(n14246), .A2(n14245), .ZN(n14244) );
  AOI21_X1 U7900 ( .B1(n6649), .B2(n8895), .A(n6731), .ZN(n7599) );
  NOR2_X1 U7901 ( .A1(n7371), .A2(n6660), .ZN(n7093) );
  INV_X1 U7902 ( .A(n11673), .ZN(n7094) );
  OR2_X1 U7903 ( .A1(n8966), .A2(n7095), .ZN(n7092) );
  INV_X1 U7904 ( .A(n7096), .ZN(n7095) );
  OR2_X1 U7905 ( .A1(n12553), .A2(n8895), .ZN(n7602) );
  NAND2_X1 U7906 ( .A1(n12557), .A2(n11685), .ZN(n12541) );
  OR2_X1 U7907 ( .A1(n8873), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8887) );
  OR2_X1 U7908 ( .A1(n12687), .A2(n12355), .ZN(n11681) );
  AOI21_X1 U7909 ( .B1(n7597), .B2(n7109), .A(n6726), .ZN(n7595) );
  INV_X1 U7910 ( .A(n7597), .ZN(n7596) );
  NOR2_X1 U7911 ( .A1(n12593), .A2(n7598), .ZN(n7597) );
  INV_X1 U7912 ( .A(n8844), .ZN(n7598) );
  NOR2_X1 U7913 ( .A1(n6646), .A2(n11651), .ZN(n7111) );
  INV_X1 U7914 ( .A(n7384), .ZN(n7383) );
  OAI21_X1 U7915 ( .B1(n6651), .B2(n6646), .A(n11660), .ZN(n7384) );
  NAND2_X1 U7916 ( .A1(n8843), .A2(n12604), .ZN(n12607) );
  NAND2_X1 U7917 ( .A1(n12644), .A2(n6651), .ZN(n12629) );
  NAND2_X1 U7918 ( .A1(n12645), .A2(n12647), .ZN(n12644) );
  NAND2_X1 U7919 ( .A1(n8805), .A2(n11651), .ZN(n12649) );
  AOI21_X1 U7920 ( .B1(n11378), .B2(n7087), .A(n7084), .ZN(n7083) );
  NAND2_X1 U7921 ( .A1(n7085), .A2(n11737), .ZN(n7084) );
  NAND2_X1 U7922 ( .A1(n7087), .A2(n7089), .ZN(n7085) );
  NAND2_X1 U7923 ( .A1(n11441), .A2(n7090), .ZN(n7089) );
  NAND2_X1 U7924 ( .A1(n11735), .A2(n11630), .ZN(n7090) );
  OR2_X1 U7925 ( .A1(n11474), .A2(n11631), .ZN(n11440) );
  OAI21_X1 U7926 ( .B1(n14259), .B2(n11625), .A(n11627), .ZN(n11378) );
  OR2_X1 U7927 ( .A1(n14291), .A2(n14290), .ZN(n7604) );
  NAND2_X1 U7928 ( .A1(n7604), .A2(n7603), .ZN(n14267) );
  AND2_X1 U7929 ( .A1(n8734), .A2(n8716), .ZN(n7603) );
  INV_X1 U7930 ( .A(n14272), .ZN(n8734) );
  AND2_X1 U7931 ( .A1(n11620), .A2(n11621), .ZN(n14272) );
  AND2_X1 U7932 ( .A1(n14290), .A2(n8961), .ZN(n7389) );
  AOI21_X1 U7933 ( .B1(n7077), .B2(n7079), .A(n7075), .ZN(n7074) );
  INV_X1 U7934 ( .A(n7077), .ZN(n7076) );
  OR2_X1 U7935 ( .A1(n11024), .A2(n11605), .ZN(n11025) );
  OR2_X1 U7936 ( .A1(n10945), .A2(n11720), .ZN(n10947) );
  AND4_X1 U7937 ( .A1(n8674), .A2(n8673), .A3(n8672), .A4(n8671), .ZN(n11336)
         );
  NOR2_X1 U7938 ( .A1(n8638), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8652) );
  NAND2_X1 U7939 ( .A1(n7594), .A2(n7593), .ZN(n10706) );
  AND2_X1 U7940 ( .A1(n8622), .A2(n8604), .ZN(n7593) );
  NAND2_X1 U7941 ( .A1(n10585), .A2(n11719), .ZN(n10584) );
  AND4_X1 U7942 ( .A1(n8569), .A2(n8568), .A3(n8567), .A4(n8566), .ZN(n15118)
         );
  NAND2_X1 U7943 ( .A1(n8837), .A2(n8836), .ZN(n12343) );
  AND2_X1 U7944 ( .A1(n8944), .A2(n11711), .ZN(n12375) );
  NAND2_X1 U7945 ( .A1(n11534), .A2(n11533), .ZN(n11548) );
  OR2_X1 U7946 ( .A1(n11532), .A2(n11531), .ZN(n11534) );
  NAND2_X1 U7947 ( .A1(n8443), .A2(n8442), .ZN(n8921) );
  INV_X1 U7948 ( .A(n8943), .ZN(n11753) );
  OR2_X1 U7949 ( .A1(n8437), .A2(n11333), .ZN(n8438) );
  AND2_X1 U7950 ( .A1(n8461), .A2(n8456), .ZN(n7606) );
  AND4_X1 U7951 ( .A1(n8460), .A2(n8459), .A3(n8458), .A4(n8457), .ZN(n8461)
         );
  INV_X1 U7952 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8458) );
  INV_X1 U7953 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8457) );
  INV_X1 U7954 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8478) );
  XNOR2_X1 U7955 ( .A(n8473), .B(n15330), .ZN(n9939) );
  OAI21_X1 U7956 ( .B1(n8503), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8473) );
  NAND2_X1 U7957 ( .A1(n8471), .A2(n8472), .ZN(n8509) );
  NAND2_X1 U7958 ( .A1(n8423), .A2(n8422), .ZN(n8808) );
  NAND2_X1 U7959 ( .A1(n7325), .A2(n7324), .ZN(n8780) );
  AOI21_X1 U7960 ( .B1(n7327), .B2(n7329), .A(n6782), .ZN(n7324) );
  AND2_X1 U7961 ( .A1(n8725), .A2(n8724), .ZN(n12466) );
  AND2_X1 U7962 ( .A1(n8405), .A2(n8404), .ZN(n8692) );
  NAND2_X1 U7963 ( .A1(n8693), .A2(n8692), .ZN(n8695) );
  OR2_X1 U7964 ( .A1(n8696), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n8711) );
  INV_X1 U7965 ( .A(n8675), .ZN(n7303) );
  OR2_X1 U7966 ( .A1(n8680), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n8696) );
  NOR2_X1 U7967 ( .A1(n8721), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n8660) );
  NAND2_X1 U7968 ( .A1(n8613), .A2(n8612), .ZN(n8615) );
  AND2_X1 U7969 ( .A1(n8572), .A2(n8451), .ZN(n8617) );
  NOR2_X1 U7970 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n8451) );
  NAND2_X1 U7971 ( .A1(n8571), .A2(n8570), .ZN(n7313) );
  INV_X1 U7972 ( .A(n12917), .ZN(n12793) );
  NAND2_X1 U7973 ( .A1(n7499), .A2(n6712), .ZN(n11288) );
  INV_X1 U7974 ( .A(n8084), .ZN(n8082) );
  AND2_X1 U7975 ( .A1(n7503), .A2(n6759), .ZN(n7501) );
  AND2_X1 U7976 ( .A1(n12885), .A2(n12145), .ZN(n7535) );
  NAND2_X1 U7977 ( .A1(n12113), .A2(n6707), .ZN(n7159) );
  NOR2_X1 U7978 ( .A1(n12097), .A2(n12096), .ZN(n6954) );
  AND2_X1 U7979 ( .A1(n8219), .A2(n8218), .ZN(n12828) );
  AND2_X1 U7980 ( .A1(n8197), .A2(n8196), .ZN(n12890) );
  INV_X1 U7981 ( .A(n8259), .ZN(n11832) );
  OR2_X1 U7982 ( .A1(n13046), .A2(n13045), .ZN(n13048) );
  NAND2_X1 U7983 ( .A1(n8328), .A2(n6679), .ZN(n13093) );
  NAND2_X1 U7984 ( .A1(n7059), .A2(n7054), .ZN(n7426) );
  NOR2_X1 U7985 ( .A1(n7060), .A2(n7057), .ZN(n7054) );
  INV_X1 U7986 ( .A(n8137), .ZN(n7060) );
  AOI21_X1 U7987 ( .B1(n8137), .B2(n7428), .A(n6719), .ZN(n7427) );
  INV_X1 U7988 ( .A(n8119), .ZN(n7428) );
  INV_X1 U7989 ( .A(n12091), .ZN(n13094) );
  OR2_X1 U7990 ( .A1(n8110), .A2(n12864), .ZN(n8130) );
  INV_X1 U7991 ( .A(n7059), .ZN(n7055) );
  NAND2_X1 U7992 ( .A1(n7059), .A2(n7056), .ZN(n13118) );
  NAND2_X1 U7993 ( .A1(n13137), .A2(n12064), .ZN(n7539) );
  NOR2_X1 U7994 ( .A1(n13161), .A2(n7507), .ZN(n7506) );
  INV_X1 U7995 ( .A(n8323), .ZN(n7507) );
  NAND2_X1 U7996 ( .A1(n7961), .A2(n7960), .ZN(n11934) );
  AOI21_X1 U7997 ( .B1(n7489), .B2(n7488), .A(n6734), .ZN(n7487) );
  INV_X1 U7998 ( .A(n7494), .ZN(n7488) );
  INV_X1 U7999 ( .A(n7927), .ZN(n7439) );
  NAND2_X1 U8000 ( .A1(n11101), .A2(n7927), .ZN(n11161) );
  INV_X1 U8001 ( .A(n10962), .ZN(n7498) );
  NOR2_X1 U8002 ( .A1(n7442), .A2(n7441), .ZN(n7440) );
  NAND2_X1 U8003 ( .A1(n11103), .A2(n11102), .ZN(n11101) );
  OR2_X1 U8004 ( .A1(n10601), .A2(n7432), .ZN(n7049) );
  NAND2_X1 U8005 ( .A1(n10569), .A2(n7514), .ZN(n10986) );
  NAND2_X1 U8006 ( .A1(n10569), .A2(n8308), .ZN(n10984) );
  NAND2_X1 U8007 ( .A1(n10369), .A2(n10372), .ZN(n7537) );
  NAND2_X1 U8008 ( .A1(n7024), .A2(n7791), .ZN(n10399) );
  INV_X1 U8009 ( .A(n12073), .ZN(n10398) );
  NAND2_X1 U8010 ( .A1(n8280), .A2(n8279), .ZN(n14304) );
  NOR2_X1 U8011 ( .A1(n13049), .A2(n12983), .ZN(n9813) );
  NAND2_X1 U8012 ( .A1(n7437), .A2(n7436), .ZN(n13006) );
  NAND2_X1 U8013 ( .A1(n8176), .A2(n8175), .ZN(n13066) );
  OR2_X1 U8014 ( .A1(n8209), .A2(n11334), .ZN(n8176) );
  NAND2_X1 U8015 ( .A1(n8160), .A2(n8159), .ZN(n13257) );
  OR2_X1 U8016 ( .A1(n10723), .A2(n8209), .ZN(n8062) );
  NAND2_X1 U8017 ( .A1(n8040), .A2(n8039), .ZN(n13289) );
  XNOR2_X1 U8018 ( .A(n10195), .B(n12105), .ZN(n7173) );
  AND2_X1 U8019 ( .A1(n7709), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7444) );
  NAND2_X1 U8020 ( .A1(n7708), .A2(n7525), .ZN(n7524) );
  INV_X1 U8021 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7525) );
  XNOR2_X1 U8022 ( .A(n8356), .B(P2_IR_REG_26__SCAN_IN), .ZN(n8373) );
  NAND2_X1 U8023 ( .A1(n7705), .A2(n7422), .ZN(n7706) );
  INV_X1 U8024 ( .A(n8272), .ZN(n7422) );
  NOR2_X1 U8025 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n8273) );
  AND3_X1 U8026 ( .A1(n7702), .A2(n7866), .A3(n7703), .ZN(n8076) );
  INV_X1 U8027 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8075) );
  OR2_X1 U8028 ( .A1(n7583), .A2(n13557), .ZN(n7582) );
  INV_X1 U8029 ( .A(n7584), .ZN(n7583) );
  INV_X1 U8030 ( .A(n13588), .ZN(n11415) );
  OR2_X1 U8031 ( .A1(n7554), .A2(n7552), .ZN(n7551) );
  INV_X1 U8032 ( .A(n7557), .ZN(n7552) );
  AND2_X1 U8033 ( .A1(n13551), .A2(n7555), .ZN(n7554) );
  OR2_X1 U8034 ( .A1(n7556), .A2(n13518), .ZN(n7555) );
  NAND2_X1 U8035 ( .A1(n7557), .A2(n13404), .ZN(n7553) );
  NAND2_X1 U8036 ( .A1(n9043), .A2(n6718), .ZN(n9045) );
  NAND2_X1 U8037 ( .A1(n10150), .A2(n13476), .ZN(n10151) );
  NAND2_X1 U8038 ( .A1(n13508), .A2(n13509), .ZN(n13507) );
  NAND2_X1 U8039 ( .A1(n7567), .A2(n7566), .ZN(n13488) );
  INV_X1 U8040 ( .A(n13538), .ZN(n7567) );
  AND2_X1 U8041 ( .A1(n13542), .A2(n7565), .ZN(n7564) );
  OR2_X1 U8042 ( .A1(n7566), .A2(n7570), .ZN(n7565) );
  NAND2_X1 U8043 ( .A1(n13498), .A2(n13499), .ZN(n7585) );
  NAND3_X1 U8044 ( .A1(n6913), .A2(n6912), .A3(n6689), .ZN(n6911) );
  AND4_X1 U8045 ( .A1(n9164), .A2(n9163), .A3(n9162), .A4(n9161), .ZN(n11207)
         );
  NOR2_X1 U8046 ( .A1(n14459), .A2(n14460), .ZN(n14458) );
  NAND2_X1 U8047 ( .A1(n13339), .A2(n9488), .ZN(n9509) );
  NAND2_X1 U8048 ( .A1(n13759), .A2(n7289), .ZN(n13708) );
  NAND2_X1 U8049 ( .A1(n13759), .A2(n13743), .ZN(n13735) );
  NAND2_X1 U8050 ( .A1(n13764), .A2(n11775), .ZN(n13747) );
  OR2_X1 U8051 ( .A1(n11795), .A2(n13736), .ZN(n7684) );
  OR2_X1 U8052 ( .A1(n13751), .A2(n11794), .ZN(n13752) );
  NAND2_X1 U8053 ( .A1(n7194), .A2(n7193), .ZN(n7350) );
  AOI21_X1 U8054 ( .B1(n13808), .B2(n11790), .A(n13786), .ZN(n7193) );
  NAND2_X1 U8055 ( .A1(n7296), .A2(n13983), .ZN(n13810) );
  OR2_X1 U8056 ( .A1(n13803), .A2(n13808), .ZN(n13801) );
  OAI21_X1 U8057 ( .B1(n11769), .B2(n7279), .A(n7277), .ZN(n13809) );
  INV_X1 U8058 ( .A(n7278), .ZN(n7277) );
  OAI21_X1 U8059 ( .B1(n7281), .B2(n7279), .A(n11771), .ZN(n7278) );
  NAND2_X1 U8060 ( .A1(n13809), .A2(n13808), .ZN(n13807) );
  NAND2_X1 U8061 ( .A1(n11769), .A2(n7281), .ZN(n13837) );
  NOR2_X1 U8062 ( .A1(n13832), .A2(n7356), .ZN(n7355) );
  INV_X1 U8063 ( .A(n11787), .ZN(n7356) );
  NAND2_X1 U8064 ( .A1(n13868), .A2(n13867), .ZN(n13866) );
  NAND2_X1 U8065 ( .A1(n13866), .A2(n7198), .ZN(n13849) );
  OAI21_X1 U8066 ( .B1(n13865), .B2(n11767), .A(n11766), .ZN(n13848) );
  OR2_X1 U8067 ( .A1(n13904), .A2(n14015), .ZN(n13888) );
  INV_X1 U8068 ( .A(n13919), .ZN(n7177) );
  INV_X1 U8069 ( .A(n11782), .ZN(n7358) );
  NAND2_X1 U8070 ( .A1(n13919), .A2(n13918), .ZN(n13917) );
  AND2_X1 U8071 ( .A1(n7679), .A2(n11760), .ZN(n7685) );
  NAND2_X1 U8072 ( .A1(n7685), .A2(n13923), .ZN(n13922) );
  NAND2_X1 U8073 ( .A1(n14170), .A2(n14171), .ZN(n6810) );
  AND2_X1 U8074 ( .A1(n11780), .A2(n9266), .ZN(n11426) );
  NAND2_X1 U8075 ( .A1(n7184), .A2(n7183), .ZN(n11358) );
  AND2_X1 U8076 ( .A1(n7185), .A2(n11263), .ZN(n7184) );
  OR2_X1 U8077 ( .A1(n7188), .A2(n7186), .ZN(n7185) );
  INV_X1 U8078 ( .A(n14539), .ZN(n13913) );
  NAND2_X1 U8079 ( .A1(n7187), .A2(n7188), .ZN(n11262) );
  AND4_X1 U8080 ( .A1(n9149), .A2(n9148), .A3(n9147), .A4(n9146), .ZN(n14536)
         );
  NOR2_X1 U8081 ( .A1(n14533), .A2(n14534), .ZN(n14532) );
  INV_X1 U8082 ( .A(n11199), .ZN(n14534) );
  NAND2_X1 U8083 ( .A1(n14548), .A2(n14549), .ZN(n7348) );
  NAND2_X1 U8084 ( .A1(n11119), .A2(n11118), .ZN(n14550) );
  NOR2_X1 U8085 ( .A1(n10906), .A2(n14631), .ZN(n14563) );
  NAND2_X1 U8086 ( .A1(n10894), .A2(n10893), .ZN(n10896) );
  AOI21_X1 U8087 ( .B1(n10902), .B2(n10901), .A(n7681), .ZN(n11129) );
  NAND2_X1 U8088 ( .A1(n13596), .A2(n10898), .ZN(n10901) );
  NAND2_X1 U8089 ( .A1(n10023), .A2(n13614), .ZN(n14537) );
  NAND2_X1 U8090 ( .A1(n10023), .A2(n9571), .ZN(n14539) );
  NAND2_X1 U8091 ( .A1(n9312), .A2(n9311), .ZN(n14009) );
  OR2_X1 U8092 ( .A1(n10723), .A2(n9485), .ZN(n9312) );
  NAND2_X1 U8093 ( .A1(n9222), .A2(n9221), .ZN(n14156) );
  AND2_X1 U8094 ( .A1(n9168), .A2(n9167), .ZN(n14658) );
  AOI21_X1 U8095 ( .B1(n7626), .B2(n9503), .A(n6789), .ZN(n7625) );
  NAND2_X1 U8096 ( .A1(n7628), .A2(n9506), .ZN(n7627) );
  XNOR2_X1 U8097 ( .A(n9504), .B(n7628), .ZN(n12012) );
  NAND2_X1 U8098 ( .A1(n9028), .A2(n9027), .ZN(n9570) );
  MUX2_X1 U8099 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9025), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n9028) );
  NAND2_X1 U8100 ( .A1(n6813), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9025) );
  NAND2_X1 U8101 ( .A1(n8241), .A2(n8240), .ZN(n8253) );
  NAND2_X1 U8102 ( .A1(n8238), .A2(n8237), .ZN(n8241) );
  NAND2_X1 U8103 ( .A1(n9564), .A2(n9010), .ZN(n9567) );
  NAND2_X1 U8104 ( .A1(n7643), .A2(n6670), .ZN(n8222) );
  NAND2_X1 U8105 ( .A1(n8187), .A2(n8186), .ZN(n8202) );
  INV_X1 U8106 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n9007) );
  OR2_X1 U8107 ( .A1(n8157), .A2(n8156), .ZN(n8169) );
  AND2_X1 U8108 ( .A1(n8991), .A2(n6757), .ZN(n8999) );
  INV_X1 U8109 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n7419) );
  AND2_X1 U8110 ( .A1(n9307), .A2(n9005), .ZN(n7421) );
  OR2_X1 U8111 ( .A1(n8102), .A2(n10325), .ZN(n8120) );
  INV_X1 U8112 ( .A(n6896), .ZN(n6895) );
  OR2_X1 U8113 ( .A1(n8057), .A2(n8094), .ZN(n8071) );
  AND2_X2 U8114 ( .A1(n9294), .A2(n9004), .ZN(n8991) );
  INV_X1 U8115 ( .A(n7612), .ZN(n6991) );
  NAND2_X1 U8116 ( .A1(n7860), .A2(n7859), .ZN(n7864) );
  AND2_X1 U8117 ( .A1(n7192), .A2(n7783), .ZN(n6910) );
  AND2_X1 U8118 ( .A1(n7801), .A2(n7764), .ZN(n7192) );
  INV_X1 U8119 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9064) );
  INV_X1 U8120 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7587) );
  NAND2_X1 U8121 ( .A1(n7035), .A2(n7033), .ZN(n7765) );
  AND3_X1 U8122 ( .A1(n6988), .A2(n6892), .A3(n6891), .ZN(n6894) );
  NAND2_X1 U8123 ( .A1(n6988), .A2(n6892), .ZN(n7730) );
  NAND2_X1 U8124 ( .A1(n7545), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n7544) );
  XNOR2_X1 U8125 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), 
        .ZN(n14075) );
  XNOR2_X1 U8126 ( .A(n6862), .B(P1_ADDR_REG_4__SCAN_IN), .ZN(n14087) );
  NAND2_X1 U8127 ( .A1(n14090), .A2(n14055), .ZN(n14056) );
  OAI21_X1 U8128 ( .B1(n15608), .B2(n15609), .A(n6682), .ZN(n7020) );
  AND3_X1 U8129 ( .A1(n8649), .A2(n8648), .A3(n8647), .ZN(n12184) );
  NAND2_X1 U8130 ( .A1(n6874), .A2(n6873), .ZN(n11490) );
  AND3_X1 U8131 ( .A1(n8591), .A2(n8590), .A3(n8589), .ZN(n12258) );
  NAND2_X1 U8132 ( .A1(n12181), .A2(n11144), .ZN(n12285) );
  NAND2_X1 U8133 ( .A1(n12346), .A2(n12213), .ZN(n12297) );
  NAND2_X1 U8134 ( .A1(n10564), .A2(n10563), .ZN(n10740) );
  NAND2_X1 U8135 ( .A1(n8800), .A2(n8799), .ZN(n12653) );
  XNOR2_X1 U8136 ( .A(n12218), .B(n12216), .ZN(n12353) );
  AND4_X1 U8137 ( .A1(n8708), .A2(n8707), .A3(n8706), .A4(n8705), .ZN(n12249)
         );
  AND2_X1 U8138 ( .A1(n8715), .A2(n8714), .ZN(n14288) );
  NAND2_X1 U8139 ( .A1(n6652), .A2(n11752), .ZN(n7114) );
  NAND2_X1 U8140 ( .A1(n8917), .A2(n8916), .ZN(n12387) );
  INV_X1 U8141 ( .A(n12210), .ZN(n12391) );
  NAND4_X1 U8142 ( .A1(n8691), .A2(n8690), .A3(n8689), .A4(n8688), .ZN(n12400)
         );
  INV_X1 U8143 ( .A(n11146), .ZN(n12402) );
  AND2_X1 U8144 ( .A1(n10799), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n14965) );
  OR2_X1 U8145 ( .A1(n10804), .A2(n10826), .ZN(n7454) );
  INV_X1 U8146 ( .A(n6978), .ZN(n12461) );
  XNOR2_X1 U8147 ( .A(n7068), .B(n15041), .ZN(n15039) );
  AND2_X1 U8148 ( .A1(n7460), .A2(n6683), .ZN(n15091) );
  AND2_X1 U8149 ( .A1(n15054), .A2(n12418), .ZN(n12419) );
  AND2_X1 U8150 ( .A1(n15025), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n6996) );
  AND2_X1 U8151 ( .A1(n15016), .A2(n12483), .ZN(n7345) );
  XNOR2_X1 U8152 ( .A(n6825), .B(n6824), .ZN(n7067) );
  INV_X1 U8153 ( .A(n12481), .ZN(n6824) );
  NOR2_X1 U8154 ( .A1(n14244), .A2(n6959), .ZN(n6825) );
  NOR2_X1 U8155 ( .A1(n12480), .A2(n12712), .ZN(n6959) );
  OAI21_X1 U8156 ( .B1(n10701), .B2(n7079), .A(n7077), .ZN(n10924) );
  AND2_X1 U8157 ( .A1(n12496), .A2(n14289), .ZN(n6961) );
  INV_X1 U8158 ( .A(n12513), .ZN(n12732) );
  AND2_X1 U8159 ( .A1(n12668), .A2(n12667), .ZN(n12730) );
  MUX2_X1 U8160 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8464), .S(
        P3_IR_REG_28__SCAN_IN), .Z(n8465) );
  NAND2_X1 U8161 ( .A1(n8503), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8500) );
  OR2_X1 U8162 ( .A1(n10531), .A2(n10530), .ZN(n7484) );
  AND2_X1 U8163 ( .A1(n11401), .A2(n11400), .ZN(n11403) );
  NAND2_X1 U8164 ( .A1(n12877), .A2(n7157), .ZN(n12808) );
  NAND2_X1 U8165 ( .A1(n7147), .A2(n7145), .ZN(n12815) );
  AOI21_X1 U8166 ( .B1(n7148), .B2(n7151), .A(n7146), .ZN(n7145) );
  INV_X1 U8167 ( .A(n12816), .ZN(n7146) );
  NAND2_X1 U8168 ( .A1(n7144), .A2(n7148), .ZN(n12817) );
  OR2_X1 U8169 ( .A1(n12877), .A2(n7151), .ZN(n7144) );
  INV_X1 U8170 ( .A(n7141), .ZN(n7140) );
  NAND2_X1 U8171 ( .A1(n7152), .A2(n7153), .ZN(n12862) );
  NAND2_X1 U8172 ( .A1(n12877), .A2(n7154), .ZN(n7152) );
  NAND2_X1 U8173 ( .A1(n8141), .A2(n8140), .ZN(n13262) );
  NAND2_X1 U8174 ( .A1(n9819), .A2(n9818), .ZN(n12908) );
  AND2_X1 U8175 ( .A1(n12053), .A2(n12054), .ZN(n7629) );
  NOR3_X1 U8176 ( .A1(n12035), .A2(n12038), .A3(n12034), .ZN(n12055) );
  INV_X1 U8177 ( .A(n12828), .ZN(n12919) );
  NAND2_X1 U8178 ( .A1(n7737), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n7714) );
  NAND2_X1 U8179 ( .A1(n7736), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7715) );
  NAND2_X1 U8180 ( .A1(n7228), .A2(n7227), .ZN(n13223) );
  NOR2_X1 U8181 ( .A1(n12996), .A2(n13049), .ZN(n7227) );
  OR2_X1 U8182 ( .A1(n14041), .A2(n8209), .ZN(n8211) );
  NAND2_X1 U8183 ( .A1(n7491), .A2(n7492), .ZN(n11159) );
  NAND2_X1 U8184 ( .A1(n10962), .A2(n7494), .ZN(n7491) );
  NAND2_X1 U8185 ( .A1(n7908), .A2(n7907), .ZN(n11910) );
  OR2_X1 U8186 ( .A1(n9791), .A2(n8209), .ZN(n7908) );
  NAND2_X1 U8187 ( .A1(n7891), .A2(n7890), .ZN(n11905) );
  AND2_X2 U8188 ( .A1(n8978), .A2(n10190), .ZN(n14934) );
  NAND2_X1 U8189 ( .A1(n13223), .A2(n13222), .ZN(n13309) );
  AND2_X1 U8190 ( .A1(n8346), .A2(n11837), .ZN(n7045) );
  INV_X1 U8191 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n15387) );
  NAND2_X1 U8192 ( .A1(n9445), .A2(n9444), .ZN(n13951) );
  NAND2_X1 U8193 ( .A1(n11830), .A2(n9488), .ZN(n9445) );
  AND2_X1 U8194 ( .A1(n13379), .A2(n13378), .ZN(n14343) );
  NAND2_X1 U8195 ( .A1(n13424), .A2(n13425), .ZN(n6919) );
  NAND2_X1 U8196 ( .A1(n9388), .A2(n9387), .ZN(n13979) );
  NAND2_X1 U8197 ( .A1(n9187), .A2(n9186), .ZN(n14357) );
  NAND2_X1 U8198 ( .A1(n7572), .A2(n7575), .ZN(n13482) );
  AOI21_X1 U8199 ( .B1(n7578), .B2(n7576), .A(n6733), .ZN(n7575) );
  NAND2_X1 U8200 ( .A1(n11315), .A2(n6661), .ZN(n11388) );
  NAND2_X1 U8201 ( .A1(n9404), .A2(n9403), .ZN(n13973) );
  NAND2_X1 U8202 ( .A1(n9203), .A2(n9202), .ZN(n11356) );
  INV_X1 U8203 ( .A(n13737), .ZN(n13704) );
  NAND3_X1 U8204 ( .A1(n10011), .A2(n10010), .A3(n14665), .ZN(n13564) );
  NAND2_X1 U8205 ( .A1(n7585), .A2(n13444), .ZN(n6976) );
  INV_X1 U8206 ( .A(n13557), .ZN(n6975) );
  OR2_X1 U8207 ( .A1(n14041), .A2(n9485), .ZN(n9433) );
  AND2_X1 U8208 ( .A1(n11017), .A2(n14632), .ZN(n14358) );
  INV_X1 U8209 ( .A(n11092), .ZN(n10867) );
  AND2_X1 U8210 ( .A1(n13649), .A2(n7212), .ZN(n10240) );
  NAND2_X1 U8211 ( .A1(n13645), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n7212) );
  AND2_X1 U8212 ( .A1(n13646), .A2(n6949), .ZN(n10233) );
  NAND2_X1 U8213 ( .A1(n13645), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6949) );
  AND2_X1 U8214 ( .A1(n7211), .A2(n7210), .ZN(n10179) );
  NAND2_X1 U8215 ( .A1(n10235), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n7210) );
  INV_X1 U8216 ( .A(n7201), .ZN(n14503) );
  NAND2_X1 U8217 ( .A1(n6807), .A2(n13726), .ZN(n6806) );
  NAND2_X1 U8218 ( .A1(n13727), .A2(n13728), .ZN(n6807) );
  NAND2_X1 U8219 ( .A1(n13958), .A2(n11776), .ZN(n13727) );
  AND2_X1 U8220 ( .A1(n9348), .A2(n9347), .ZN(n13995) );
  AOI21_X1 U8221 ( .B1(n13936), .B2(n14554), .A(n7180), .ZN(n7276) );
  NAND2_X1 U8222 ( .A1(n7182), .A2(n7181), .ZN(n7180) );
  AOI21_X1 U8223 ( .B1(n13941), .B2(n14632), .A(n13940), .ZN(n7181) );
  OAI211_X1 U8224 ( .C1(n13945), .C2(n11801), .A(n7134), .B(n6728), .ZN(n13942) );
  NOR2_X1 U8225 ( .A1(n11800), .A2(n7274), .ZN(n7273) );
  NOR2_X1 U8226 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n7284) );
  INV_X1 U8227 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10725) );
  NAND2_X1 U8228 ( .A1(n15615), .A2(n15616), .ZN(n14081) );
  XNOR2_X1 U8229 ( .A(n14098), .B(P2_ADDR_REG_7__SCAN_IN), .ZN(n15608) );
  XNOR2_X1 U8230 ( .A(n7020), .B(n14102), .ZN(n14146) );
  NAND2_X1 U8231 ( .A1(n14110), .A2(n14109), .ZN(n6926) );
  XNOR2_X1 U8232 ( .A(n14116), .B(n14115), .ZN(n14413) );
  NOR2_X1 U8233 ( .A1(n6678), .A2(n14124), .ZN(n14425) );
  INV_X1 U8234 ( .A(n14124), .ZN(n6968) );
  NAND2_X1 U8235 ( .A1(n9499), .A2(n12178), .ZN(n7396) );
  NAND2_X1 U8236 ( .A1(n9109), .A2(n7417), .ZN(n7416) );
  NAND2_X1 U8237 ( .A1(n9140), .A2(n9142), .ZN(n7407) );
  NAND2_X1 U8238 ( .A1(n9878), .A2(n7214), .ZN(n6985) );
  NAND2_X1 U8239 ( .A1(n7664), .A2(n7665), .ZN(n7662) );
  INV_X1 U8240 ( .A(n11872), .ZN(n7664) );
  INV_X1 U8241 ( .A(n11867), .ZN(n6836) );
  AND2_X1 U8242 ( .A1(n11872), .A2(n11871), .ZN(n7663) );
  AND2_X1 U8243 ( .A1(n7662), .A2(n6750), .ZN(n7001) );
  NAND2_X1 U8244 ( .A1(n9188), .A2(n7415), .ZN(n7414) );
  NAND2_X1 U8245 ( .A1(n6673), .A2(n11916), .ZN(n7677) );
  OAI22_X1 U8246 ( .A1(n6857), .A2(n6856), .B1(n11892), .B2(n11891), .ZN(
        n11899) );
  NOR2_X1 U8247 ( .A1(n7002), .A2(n7000), .ZN(n6856) );
  INV_X1 U8248 ( .A(n11892), .ZN(n7000) );
  NAND2_X1 U8249 ( .A1(n9240), .A2(n7410), .ZN(n7409) );
  INV_X1 U8250 ( .A(n11931), .ZN(n6946) );
  INV_X1 U8251 ( .A(n11930), .ZN(n6945) );
  NAND2_X1 U8252 ( .A1(n11584), .A2(n11721), .ZN(n6932) );
  AND2_X1 U8253 ( .A1(n11580), .A2(n11579), .ZN(n6933) );
  NAND2_X1 U8254 ( .A1(n13850), .A2(n6943), .ZN(n6942) );
  AND2_X1 U8255 ( .A1(n9320), .A2(n13884), .ZN(n6943) );
  OAI21_X1 U8256 ( .B1(n11939), .B2(n6844), .A(n6843), .ZN(n11948) );
  NAND2_X1 U8257 ( .A1(n6845), .A2(n6703), .ZN(n6843) );
  NOR2_X1 U8258 ( .A1(n6845), .A2(n6703), .ZN(n6844) );
  NAND2_X1 U8259 ( .A1(n11948), .A2(n11947), .ZN(n11945) );
  INV_X1 U8260 ( .A(n11948), .ZN(n6928) );
  INV_X1 U8261 ( .A(n11947), .ZN(n6927) );
  OAI21_X1 U8262 ( .B1(n11957), .B2(n6855), .A(n6854), .ZN(n11964) );
  NAND2_X1 U8263 ( .A1(n11956), .A2(n6774), .ZN(n6854) );
  NOR2_X1 U8264 ( .A1(n11956), .A2(n6774), .ZN(n6855) );
  NAND2_X1 U8265 ( .A1(n11964), .A2(n11965), .ZN(n11963) );
  NAND2_X1 U8266 ( .A1(n9405), .A2(n9407), .ZN(n7393) );
  NAND2_X1 U8267 ( .A1(n11983), .A2(n6773), .ZN(n7667) );
  OR2_X1 U8268 ( .A1(n9435), .A2(n7405), .ZN(n7403) );
  INV_X1 U8269 ( .A(n11992), .ZN(n6851) );
  INV_X1 U8270 ( .A(n11993), .ZN(n6848) );
  INV_X1 U8271 ( .A(n6853), .ZN(n6849) );
  INV_X1 U8272 ( .A(n9499), .ZN(n9108) );
  INV_X1 U8273 ( .A(n15058), .ZN(n6818) );
  INV_X1 U8274 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8781) );
  NAND2_X1 U8275 ( .A1(n9461), .A2(n9463), .ZN(n7400) );
  INV_X1 U8276 ( .A(n8152), .ZN(n8154) );
  INV_X1 U8277 ( .A(n8138), .ZN(n6885) );
  AND2_X1 U8278 ( .A1(n7646), .A2(n8097), .ZN(n7645) );
  NAND2_X1 U8279 ( .A1(n7649), .A2(n7647), .ZN(n7646) );
  INV_X1 U8280 ( .A(n7649), .ZN(n7648) );
  INV_X1 U8281 ( .A(n7974), .ZN(n6882) );
  AND2_X1 U8282 ( .A1(n7633), .A2(n6674), .ZN(n6877) );
  NAND2_X1 U8283 ( .A1(n14050), .A2(n14051), .ZN(n14052) );
  NAND2_X1 U8284 ( .A1(n14085), .A2(n14049), .ZN(n14050) );
  NAND2_X1 U8285 ( .A1(n6861), .A2(n7011), .ZN(n14048) );
  NOR2_X1 U8286 ( .A1(n8494), .A2(n8493), .ZN(n9936) );
  INV_X1 U8287 ( .A(n10746), .ZN(n7258) );
  NAND2_X1 U8288 ( .A1(n11707), .A2(n11697), .ZN(n7317) );
  INV_X1 U8289 ( .A(n11712), .ZN(n7315) );
  OAI21_X1 U8290 ( .B1(n11710), .B2(n11709), .A(n11711), .ZN(n7318) );
  INV_X1 U8291 ( .A(n11707), .ZN(n7099) );
  INV_X1 U8292 ( .A(n15010), .ZN(n7465) );
  NOR2_X1 U8293 ( .A1(n14972), .A2(n6929), .ZN(n10807) );
  NOR2_X1 U8294 ( .A1(n14982), .A2(n15193), .ZN(n6929) );
  AND2_X1 U8295 ( .A1(n7339), .A2(n7338), .ZN(n12459) );
  NAND2_X1 U8296 ( .A1(n10808), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n7338) );
  NAND2_X1 U8297 ( .A1(n6820), .A2(n6819), .ZN(n7336) );
  NAND2_X1 U8298 ( .A1(n10809), .A2(n6647), .ZN(n6819) );
  AOI21_X1 U8299 ( .B1(n6647), .B2(n15199), .A(n15030), .ZN(n6820) );
  NAND2_X1 U8300 ( .A1(n15097), .A2(n12472), .ZN(n6830) );
  NOR2_X1 U8301 ( .A1(n14210), .A2(n12476), .ZN(n12477) );
  AND2_X1 U8302 ( .A1(n14214), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n12476) );
  OR2_X1 U8303 ( .A1(n8926), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n12487) );
  OR2_X1 U8304 ( .A1(n8967), .A2(n7373), .ZN(n7372) );
  INV_X1 U8305 ( .A(n11685), .ZN(n7373) );
  NOR2_X1 U8306 ( .A1(n7372), .A2(n11675), .ZN(n7096) );
  OR2_X1 U8307 ( .A1(n8788), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8813) );
  NAND2_X1 U8308 ( .A1(n8520), .A2(n8519), .ZN(n8788) );
  INV_X1 U8309 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n8519) );
  INV_X1 U8310 ( .A(n8772), .ZN(n8520) );
  INV_X1 U8311 ( .A(n11604), .ZN(n7075) );
  NOR2_X1 U8312 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), .ZN(
        n8459) );
  INV_X1 U8313 ( .A(n7328), .ZN(n7327) );
  OAI21_X1 U8314 ( .B1(n8751), .B2(n7329), .A(n8416), .ZN(n7328) );
  INV_X1 U8315 ( .A(n8415), .ZN(n7329) );
  INV_X1 U8316 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n8410) );
  INV_X1 U8317 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8722) );
  INV_X1 U8318 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8659) );
  AND2_X1 U8319 ( .A1(n8612), .A2(n8394), .ZN(n7320) );
  INV_X1 U8320 ( .A(n12843), .ZN(n7505) );
  AND2_X1 U8321 ( .A1(n7222), .A2(n7221), .ZN(n7220) );
  NOR2_X1 U8322 ( .A1(n13232), .A2(n13238), .ZN(n7222) );
  NAND2_X1 U8323 ( .A1(n7042), .A2(n13058), .ZN(n7041) );
  INV_X1 U8324 ( .A(n8091), .ZN(n7058) );
  NAND2_X1 U8325 ( .A1(n8041), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8063) );
  NAND2_X1 U8326 ( .A1(n8021), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8042) );
  INV_X1 U8327 ( .A(n8022), .ZN(n8021) );
  INV_X1 U8328 ( .A(n7899), .ZN(n7441) );
  NAND2_X1 U8329 ( .A1(n13015), .A2(n13020), .ZN(n7437) );
  AOI21_X1 U8330 ( .B1(n7530), .B2(n7528), .A(n6721), .ZN(n7527) );
  AND2_X1 U8331 ( .A1(n8335), .A2(n7531), .ZN(n7530) );
  NAND2_X1 U8332 ( .A1(n13175), .A2(n6714), .ZN(n13109) );
  AND2_X1 U8333 ( .A1(n13175), .A2(n6662), .ZN(n13126) );
  NAND2_X1 U8334 ( .A1(n13175), .A2(n7230), .ZN(n13138) );
  NAND2_X1 U8335 ( .A1(n7217), .A2(n7216), .ZN(n13190) );
  INV_X1 U8336 ( .A(n13336), .ZN(n7216) );
  INV_X1 U8337 ( .A(n14312), .ZN(n7217) );
  INV_X1 U8338 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n7761) );
  INV_X1 U8339 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7700) );
  NOR2_X1 U8340 ( .A1(n9550), .A2(n11800), .ZN(n6912) );
  XNOR2_X1 U8341 ( .A(n13695), .B(n9516), .ZN(n9551) );
  NAND2_X1 U8342 ( .A1(n6916), .A2(n6914), .ZN(n9526) );
  NAND2_X1 U8343 ( .A1(n6915), .A2(n9473), .ZN(n6914) );
  NAND2_X1 U8344 ( .A1(n9511), .A2(n9510), .ZN(n6916) );
  NAND2_X1 U8345 ( .A1(n13695), .A2(n9516), .ZN(n6915) );
  NOR2_X1 U8346 ( .A1(n9551), .A2(n9528), .ZN(n9521) );
  NOR2_X1 U8347 ( .A1(n13951), .A2(n13957), .ZN(n7291) );
  OR2_X1 U8348 ( .A1(n14009), .A2(n13853), .ZN(n11766) );
  NOR2_X1 U8349 ( .A1(n14375), .A2(n7294), .ZN(n7293) );
  INV_X1 U8350 ( .A(n7295), .ZN(n7294) );
  INV_X1 U8351 ( .A(n9482), .ZN(n6889) );
  INV_X1 U8352 ( .A(n8256), .ZN(n6888) );
  AND2_X1 U8353 ( .A1(n7589), .A2(n7363), .ZN(n7137) );
  AND2_X1 U8354 ( .A1(n9010), .A2(n9011), .ZN(n7590) );
  INV_X1 U8355 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9011) );
  NAND2_X1 U8356 ( .A1(n7651), .A2(n8055), .ZN(n8099) );
  INV_X1 U8357 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n8988) );
  NAND2_X1 U8358 ( .A1(n6881), .A2(n7974), .ZN(n8007) );
  NAND2_X1 U8359 ( .A1(n7635), .A2(n7633), .ZN(n6881) );
  INV_X1 U8360 ( .A(n7639), .ZN(n7638) );
  AOI21_X1 U8361 ( .B1(n7639), .B2(n7637), .A(n6732), .ZN(n7636) );
  INV_X1 U8362 ( .A(n7930), .ZN(n7637) );
  OR3_X1 U8363 ( .A1(n9200), .A2(n9199), .A3(n9198), .ZN(n9219) );
  OAI21_X1 U8364 ( .B1(n9371), .B2(n9614), .A(n6909), .ZN(n7803) );
  NAND2_X1 U8365 ( .A1(n9371), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n6909) );
  INV_X1 U8366 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n8985) );
  INV_X1 U8367 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6811) );
  OAI21_X1 U8368 ( .B1(n9371), .B2(n9602), .A(n6944), .ZN(n7785) );
  OR2_X1 U8369 ( .A1(n9042), .A2(n9599), .ZN(n6944) );
  OAI21_X1 U8370 ( .B1(n9042), .B2(n9596), .A(n6972), .ZN(n7766) );
  NAND2_X1 U8371 ( .A1(n9042), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n6972) );
  NAND2_X1 U8372 ( .A1(n6971), .A2(n7783), .ZN(n6937) );
  OR2_X1 U8373 ( .A1(n7766), .A2(SI_3_), .ZN(n6971) );
  OAI21_X1 U8374 ( .B1(n9042), .B2(n9600), .A(n6940), .ZN(n7752) );
  NAND2_X1 U8375 ( .A1(n9042), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n6940) );
  XNOR2_X1 U8376 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(P3_ADDR_REG_1__SCAN_IN), 
        .ZN(n14077) );
  NAND2_X1 U8377 ( .A1(n14076), .A2(n14075), .ZN(n6861) );
  NAND2_X1 U8378 ( .A1(n7012), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n7011) );
  XNOR2_X1 U8379 ( .A(n14054), .B(n6939), .ZN(n14090) );
  INV_X1 U8380 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n6939) );
  OAI21_X1 U8381 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(n14989), .A(n14058), .ZN(
        n14059) );
  INV_X1 U8382 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n15282) );
  AND2_X1 U8383 ( .A1(n7240), .A2(n6761), .ZN(n7239) );
  NAND2_X1 U8384 ( .A1(n7243), .A2(n7241), .ZN(n7240) );
  INV_X1 U8385 ( .A(n12372), .ZN(n7245) );
  INV_X1 U8386 ( .A(n12271), .ZN(n7238) );
  INV_X1 U8387 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n15313) );
  INV_X1 U8388 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n11152) );
  NAND2_X1 U8389 ( .A1(n8523), .A2(n12348), .ZN(n8849) );
  NAND2_X1 U8390 ( .A1(n7263), .A2(n7264), .ZN(n11477) );
  AOI21_X1 U8391 ( .B1(n6648), .B2(n11151), .A(n6702), .ZN(n7264) );
  NAND2_X1 U8392 ( .A1(n7254), .A2(n10081), .ZN(n10082) );
  AND2_X1 U8393 ( .A1(n10032), .A2(n10029), .ZN(n7254) );
  NAND2_X1 U8394 ( .A1(n10740), .A2(n10739), .ZN(n7259) );
  AND2_X1 U8395 ( .A1(n12304), .A2(n7247), .ZN(n7246) );
  NAND2_X1 U8396 ( .A1(n12225), .A2(n12224), .ZN(n7247) );
  INV_X1 U8397 ( .A(n7249), .ZN(n7242) );
  NOR2_X1 U8398 ( .A1(n11748), .A2(n11747), .ZN(n11749) );
  AND2_X1 U8399 ( .A1(n11546), .A2(n11545), .ZN(n12486) );
  AND3_X1 U8400 ( .A1(n8853), .A2(n8852), .A3(n8851), .ZN(n12354) );
  AND4_X1 U8401 ( .A1(n8765), .A2(n8764), .A3(n8763), .A4(n8762), .ZN(n11631)
         );
  AND4_X1 U8402 ( .A1(n8733), .A2(n8732), .A3(n8731), .A4(n8730), .ZN(n11430)
         );
  AND4_X1 U8403 ( .A1(n8610), .A2(n8609), .A3(n8608), .A4(n8607), .ZN(n10742)
         );
  NAND2_X1 U8404 ( .A1(n6827), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n9851) );
  NAND2_X1 U8405 ( .A1(n9967), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n9850) );
  NAND2_X1 U8406 ( .A1(n9855), .A2(n9856), .ZN(n9854) );
  AND2_X1 U8407 ( .A1(n9862), .A2(n9861), .ZN(n9979) );
  OR2_X1 U8408 ( .A1(n14946), .A2(n14945), .ZN(n7072) );
  INV_X1 U8409 ( .A(n7072), .ZN(n14944) );
  INV_X1 U8410 ( .A(n9975), .ZN(n6955) );
  NAND2_X1 U8411 ( .A1(n6822), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n6821) );
  NOR2_X1 U8412 ( .A1(n6690), .A2(n14973), .ZN(n14972) );
  OR2_X1 U8413 ( .A1(n10809), .A2(n15199), .ZN(n6978) );
  INV_X1 U8414 ( .A(n7336), .ZN(n15029) );
  OR2_X1 U8415 ( .A1(n15089), .A2(n12420), .ZN(n7066) );
  AND2_X1 U8416 ( .A1(n6830), .A2(n14198), .ZN(n12474) );
  OAI21_X1 U8417 ( .B1(n14195), .B2(n7342), .A(n6829), .ZN(n14210) );
  NAND2_X1 U8418 ( .A1(n7343), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n7342) );
  NAND2_X1 U8419 ( .A1(n12474), .A2(n7343), .ZN(n6829) );
  INV_X1 U8420 ( .A(n14211), .ZN(n7343) );
  NOR2_X1 U8421 ( .A1(n14195), .A2(n14194), .ZN(n14193) );
  NOR2_X1 U8422 ( .A1(n14208), .A2(n7064), .ZN(n12423) );
  AND2_X1 U8423 ( .A1(n14214), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n7064) );
  NOR2_X1 U8424 ( .A1(n14247), .A2(n12451), .ZN(n12455) );
  OAI21_X1 U8425 ( .B1(n12508), .B2(n8968), .A(n11700), .ZN(n11529) );
  AND2_X1 U8426 ( .A1(n8932), .A2(n8931), .ZN(n12502) );
  OR2_X1 U8427 ( .A1(n8910), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8924) );
  NAND2_X1 U8428 ( .A1(n7091), .A2(n11691), .ZN(n12524) );
  NAND2_X1 U8429 ( .A1(n8525), .A2(n15304), .ZN(n8901) );
  INV_X1 U8430 ( .A(n8887), .ZN(n8525) );
  NAND2_X1 U8431 ( .A1(n12565), .A2(n6680), .ZN(n12557) );
  NAND2_X1 U8432 ( .A1(n8966), .A2(n11673), .ZN(n12563) );
  NAND2_X1 U8433 ( .A1(n12563), .A2(n12567), .ZN(n12565) );
  AOI21_X1 U8434 ( .B1(n7107), .B2(n7106), .A(n7105), .ZN(n7104) );
  INV_X1 U8435 ( .A(n11665), .ZN(n7105) );
  CLKBUF_X1 U8436 ( .A(n11504), .Z(n11505) );
  NOR2_X1 U8437 ( .A1(n8728), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8740) );
  OR2_X1 U8438 ( .A1(n8703), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8728) );
  AOI21_X1 U8439 ( .B1(n7389), .B2(n11605), .A(n7388), .ZN(n7387) );
  INV_X1 U8440 ( .A(n11615), .ZN(n7388) );
  AOI21_X1 U8441 ( .B1(n11720), .B2(n8685), .A(n6663), .ZN(n7591) );
  NAND2_X1 U8442 ( .A1(n7078), .A2(n6650), .ZN(n7077) );
  INV_X1 U8443 ( .A(n7081), .ZN(n7078) );
  AOI21_X1 U8444 ( .B1(n11718), .B2(n7082), .A(n6740), .ZN(n7081) );
  NAND2_X1 U8445 ( .A1(n11718), .A2(n6650), .ZN(n7079) );
  INV_X1 U8446 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n12286) );
  INV_X1 U8447 ( .A(n7080), .ZN(n10943) );
  AOI21_X1 U8448 ( .B1(n10701), .B2(n11589), .A(n11142), .ZN(n7080) );
  OR2_X1 U8449 ( .A1(n8623), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8638) );
  INV_X1 U8450 ( .A(n8958), .ZN(n11725) );
  NAND2_X1 U8451 ( .A1(n7594), .A2(n8604), .ZN(n10618) );
  INV_X1 U8452 ( .A(n8622), .ZN(n11721) );
  NAND2_X1 U8453 ( .A1(n11723), .A2(n7102), .ZN(n7100) );
  INV_X1 U8454 ( .A(n11568), .ZN(n7102) );
  NAND2_X1 U8455 ( .A1(n8576), .A2(n8956), .ZN(n10590) );
  AND2_X1 U8456 ( .A1(n10326), .A2(n12483), .ZN(n11750) );
  NAND2_X1 U8457 ( .A1(n15115), .A2(n15116), .ZN(n15114) );
  CLKBUF_X1 U8458 ( .A(n15115), .Z(n6960) );
  CLKBUF_X1 U8459 ( .A(n8564), .Z(n15112) );
  OR2_X1 U8460 ( .A1(n11379), .A2(n15179), .ZN(n14289) );
  INV_X1 U8461 ( .A(n15146), .ZN(n15157) );
  INV_X1 U8462 ( .A(n8494), .ZN(n9709) );
  OAI21_X1 U8463 ( .B1(n8543), .B2(n8446), .A(n8447), .ZN(n11532) );
  NOR2_X1 U8464 ( .A1(n8724), .A2(n7376), .ZN(n7375) );
  NAND2_X1 U8465 ( .A1(n7378), .A2(n7377), .ZN(n7376) );
  AND2_X1 U8466 ( .A1(n8467), .A2(n7381), .ZN(n7377) );
  XNOR2_X1 U8467 ( .A(n8475), .B(P3_IR_REG_26__SCAN_IN), .ZN(n8496) );
  AND2_X1 U8468 ( .A1(n8435), .A2(n8434), .ZN(n8867) );
  AND2_X1 U8469 ( .A1(n8433), .A2(n8432), .ZN(n8854) );
  INV_X1 U8470 ( .A(n8506), .ZN(n8505) );
  NAND2_X1 U8471 ( .A1(n8471), .A2(n6866), .ZN(n8506) );
  NOR2_X1 U8472 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), .ZN(
        n6866) );
  INV_X1 U8473 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8507) );
  OR2_X1 U8474 ( .A1(n8784), .A2(P3_IR_REG_16__SCAN_IN), .ZN(n8797) );
  INV_X1 U8475 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n15342) );
  AOI21_X1 U8476 ( .B1(n7332), .B2(n7334), .A(n6739), .ZN(n7330) );
  AND2_X1 U8477 ( .A1(n8398), .A2(n8396), .ZN(n8644) );
  INV_X1 U8478 ( .A(n8388), .ZN(n7311) );
  OAI21_X1 U8479 ( .B1(n12824), .B2(n7534), .A(n7532), .ZN(n12790) );
  AOI21_X1 U8480 ( .B1(n7535), .B2(n7533), .A(n6737), .ZN(n7532) );
  INV_X1 U8481 ( .A(n7535), .ZN(n7534) );
  INV_X1 U8482 ( .A(n12826), .ZN(n7533) );
  OR2_X1 U8483 ( .A1(n8161), .A2(n12802), .ZN(n8178) );
  OR2_X1 U8484 ( .A1(n8063), .A2(n14818), .ZN(n8084) );
  NOR2_X1 U8485 ( .A1(n10683), .A2(n7480), .ZN(n7479) );
  INV_X1 U8486 ( .A(n10529), .ZN(n7480) );
  NAND2_X1 U8487 ( .A1(n10530), .A2(n10529), .ZN(n7485) );
  NAND2_X1 U8488 ( .A1(n9873), .A2(n7429), .ZN(n9874) );
  INV_X1 U8489 ( .A(n12860), .ZN(n7149) );
  NAND2_X1 U8490 ( .A1(n11183), .A2(n11182), .ZN(n7499) );
  INV_X1 U8491 ( .A(n12852), .ZN(n7142) );
  NAND2_X1 U8492 ( .A1(n12834), .A2(n12833), .ZN(n12844) );
  INV_X1 U8493 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7892) );
  NAND2_X1 U8494 ( .A1(n7156), .A2(n6772), .ZN(n7153) );
  OR2_X1 U8495 ( .A1(n7941), .A2(n7940), .ZN(n7963) );
  NOR2_X1 U8496 ( .A1(n7161), .A2(n12909), .ZN(n7160) );
  INV_X1 U8497 ( .A(n7164), .ZN(n7161) );
  NAND2_X1 U8498 ( .A1(n12114), .A2(n7165), .ZN(n7164) );
  NAND2_X1 U8499 ( .A1(n12002), .A2(n12001), .ZN(n12003) );
  OR2_X1 U8500 ( .A1(n12097), .A2(n12049), .ZN(n6924) );
  NAND2_X1 U8501 ( .A1(n12048), .A2(n12030), .ZN(n12038) );
  NAND2_X1 U8502 ( .A1(n12037), .A2(n12036), .ZN(n7631) );
  NAND2_X1 U8503 ( .A1(n12040), .A2(n12039), .ZN(n7632) );
  AND2_X1 U8504 ( .A1(n8234), .A2(n8233), .ZN(n12892) );
  OR2_X1 U8505 ( .A1(n13023), .A2(n8229), .ZN(n8234) );
  AND4_X1 U8506 ( .A1(n7916), .A2(n7915), .A3(n7914), .A4(n7913), .ZN(n11909)
         );
  OR2_X1 U8507 ( .A1(n7888), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n8037) );
  OAI21_X1 U8508 ( .B1(n12096), .B2(n7031), .A(n7028), .ZN(n7027) );
  OR2_X1 U8509 ( .A1(n7436), .A2(n12096), .ZN(n7026) );
  NAND2_X1 U8510 ( .A1(n7436), .A2(n12096), .ZN(n7030) );
  NAND2_X1 U8511 ( .A1(n13051), .A2(n7222), .ZN(n13018) );
  AND2_X1 U8512 ( .A1(n13051), .A2(n13036), .ZN(n13032) );
  INV_X1 U8513 ( .A(n7517), .ZN(n7516) );
  OR2_X1 U8514 ( .A1(n13262), .A2(n13109), .ZN(n13095) );
  NAND2_X1 U8515 ( .A1(n8129), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n8143) );
  AND2_X1 U8516 ( .A1(n12065), .A2(n12064), .ZN(n13136) );
  OAI21_X1 U8517 ( .B1(n13148), .B2(n8068), .A(n8069), .ZN(n13133) );
  NAND2_X1 U8518 ( .A1(n13175), .A2(n13157), .ZN(n13152) );
  OAI21_X1 U8519 ( .B1(n7053), .B2(n7052), .A(n8048), .ZN(n13169) );
  INV_X1 U8520 ( .A(n13166), .ZN(n7052) );
  INV_X1 U8521 ( .A(n7053), .ZN(n13184) );
  AND2_X1 U8522 ( .A1(n9816), .A2(n8287), .ZN(n12902) );
  AND2_X1 U8523 ( .A1(n9816), .A2(n8291), .ZN(n12901) );
  NAND2_X1 U8524 ( .A1(n7219), .A2(n7218), .ZN(n14312) );
  NAND2_X1 U8525 ( .A1(n7039), .A2(n7969), .ZN(n14301) );
  OR2_X1 U8526 ( .A1(n7978), .A2(n11405), .ZN(n7995) );
  AOI21_X1 U8527 ( .B1(n7494), .B2(n8313), .A(n6654), .ZN(n7492) );
  AND2_X1 U8528 ( .A1(n10845), .A2(n10939), .ZN(n10968) );
  NAND2_X1 U8529 ( .A1(n10841), .A2(n7899), .ZN(n10963) );
  NAND2_X1 U8530 ( .A1(n7046), .A2(n7049), .ZN(n7048) );
  AND2_X1 U8531 ( .A1(n7430), .A2(n6743), .ZN(n7046) );
  NAND2_X1 U8532 ( .A1(n7048), .A2(n7047), .ZN(n10841) );
  NOR2_X1 U8533 ( .A1(n12080), .A2(n7051), .ZN(n7047) );
  AOI21_X1 U8534 ( .B1(n7511), .B2(n7510), .A(n7513), .ZN(n7509) );
  INV_X1 U8535 ( .A(n7514), .ZN(n7512) );
  AND2_X1 U8536 ( .A1(n12076), .A2(n8308), .ZN(n7511) );
  NAND2_X1 U8537 ( .A1(n10570), .A2(n10571), .ZN(n10569) );
  AND2_X1 U8538 ( .A1(n10378), .A2(n10370), .ZN(n10403) );
  AND2_X1 U8539 ( .A1(n10403), .A2(n14901), .ZN(n10606) );
  NAND2_X1 U8540 ( .A1(n7772), .A2(n7771), .ZN(n10373) );
  INV_X1 U8541 ( .A(n8209), .ZN(n7521) );
  INV_X1 U8542 ( .A(n9608), .ZN(n7522) );
  NAND2_X1 U8543 ( .A1(n7215), .A2(n7214), .ZN(n10049) );
  OAI211_X1 U8544 ( .C1(n9504), .C2(n7621), .A(n7619), .B(n12006), .ZN(n12989)
         );
  NAND2_X1 U8545 ( .A1(n7624), .A2(n12011), .ZN(n7621) );
  INV_X1 U8546 ( .A(n14915), .ZN(n14892) );
  NOR2_X1 U8547 ( .A1(n10189), .A2(n8376), .ZN(n8978) );
  CLKBUF_X1 U8548 ( .A(n8286), .Z(n8287) );
  NOR2_X1 U8549 ( .A1(n7706), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n7655) );
  INV_X1 U8550 ( .A(n8059), .ZN(n7656) );
  INV_X1 U8551 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8359) );
  NAND2_X1 U8552 ( .A1(n8059), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8060) );
  OR2_X1 U8553 ( .A1(n7990), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n7991) );
  AND2_X1 U8554 ( .A1(n7959), .A2(n7990), .ZN(n10335) );
  INV_X1 U8555 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n7810) );
  OR2_X1 U8556 ( .A1(n7781), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n7809) );
  CLKBUF_X1 U8557 ( .A(n7745), .Z(n7746) );
  AND2_X1 U8558 ( .A1(n7584), .A2(n13444), .ZN(n7581) );
  INV_X1 U8559 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n15558) );
  INV_X1 U8560 ( .A(n7582), .ZN(n7579) );
  INV_X1 U8561 ( .A(n7581), .ZN(n7576) );
  AND2_X1 U8562 ( .A1(n13392), .A2(n13391), .ZN(n6920) );
  CLKBUF_X1 U8563 ( .A(n13393), .Z(n6962) );
  NAND2_X1 U8564 ( .A1(n7558), .A2(n10548), .ZN(n10658) );
  INV_X1 U8565 ( .A(n10550), .ZN(n7558) );
  NAND2_X1 U8566 ( .A1(n10550), .A2(n10549), .ZN(n10655) );
  NAND2_X1 U8567 ( .A1(n10016), .A2(n10015), .ZN(n10147) );
  INV_X1 U8568 ( .A(n13405), .ZN(n6977) );
  OR2_X1 U8569 ( .A1(n9315), .A2(n9288), .ZN(n9341) );
  NAND2_X1 U8570 ( .A1(n13517), .A2(n13518), .ZN(n13516) );
  NAND2_X1 U8571 ( .A1(n9313), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9315) );
  AND2_X1 U8572 ( .A1(n10657), .A2(n7560), .ZN(n7559) );
  NAND2_X1 U8573 ( .A1(n10654), .A2(n10548), .ZN(n7560) );
  NOR2_X1 U8574 ( .A1(n10654), .A2(n10548), .ZN(n7561) );
  OR2_X1 U8575 ( .A1(n10240), .A2(n10239), .ZN(n7211) );
  NOR2_X1 U8576 ( .A1(n10423), .A2(n7205), .ZN(n14434) );
  AND2_X1 U8577 ( .A1(n10424), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7205) );
  NOR2_X1 U8578 ( .A1(n14434), .A2(n14433), .ZN(n14432) );
  AOI21_X1 U8579 ( .B1(n10424), .B2(P1_REG1_REG_10__SCAN_IN), .A(n10414), .ZN(
        n14430) );
  NAND2_X1 U8580 ( .A1(n14428), .A2(n6947), .ZN(n10416) );
  OR2_X1 U8581 ( .A1(n10426), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6947) );
  NAND2_X1 U8582 ( .A1(n10416), .A2(n10417), .ZN(n13670) );
  NOR2_X1 U8583 ( .A1(n14444), .A2(n7208), .ZN(n14459) );
  AND2_X1 U8584 ( .A1(n14449), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7208) );
  AOI21_X1 U8585 ( .B1(n14449), .B2(P1_REG1_REG_13__SCAN_IN), .A(n14441), .ZN(
        n14455) );
  XNOR2_X1 U8586 ( .A(n14478), .B(n13674), .ZN(n14470) );
  INV_X1 U8587 ( .A(n13661), .ZN(n13662) );
  NOR2_X1 U8588 ( .A1(n14458), .A2(n7207), .ZN(n13661) );
  AND2_X1 U8589 ( .A1(n14453), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7207) );
  AOI21_X1 U8590 ( .B1(n14493), .B2(P1_REG1_REG_16__SCAN_IN), .A(n14484), .ZN(
        n14499) );
  OR2_X1 U8591 ( .A1(n14488), .A2(n7202), .ZN(n7201) );
  NOR2_X1 U8592 ( .A1(n7203), .A2(n15332), .ZN(n7202) );
  INV_X1 U8593 ( .A(n14493), .ZN(n7203) );
  AND2_X1 U8594 ( .A1(n7201), .A2(n7200), .ZN(n14502) );
  INV_X1 U8595 ( .A(n14504), .ZN(n7200) );
  AOI21_X1 U8596 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n13676), .A(n14498), .ZN(
        n13677) );
  NOR2_X1 U8597 ( .A1(n14502), .A2(n7199), .ZN(n13665) );
  AND2_X1 U8598 ( .A1(n13676), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7199) );
  INV_X1 U8599 ( .A(n7367), .ZN(n7366) );
  OAI22_X1 U8600 ( .A1(n11796), .A2(n7368), .B1(n13957), .B2(n13719), .ZN(
        n7367) );
  NAND2_X1 U8601 ( .A1(n11794), .A2(n7684), .ZN(n7368) );
  NOR2_X1 U8602 ( .A1(n11796), .A2(n7370), .ZN(n7369) );
  INV_X1 U8603 ( .A(n7684), .ZN(n7370) );
  AOI21_X1 U8604 ( .B1(n7129), .B2(n7131), .A(n6724), .ZN(n7128) );
  NAND2_X1 U8605 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(n9365), .ZN(n9382) );
  AND2_X1 U8606 ( .A1(n9354), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9365) );
  OAI21_X1 U8607 ( .B1(n13866), .B2(n7197), .A(n7195), .ZN(n13824) );
  AND2_X1 U8608 ( .A1(n7196), .A2(n11788), .ZN(n7195) );
  OR2_X1 U8609 ( .A1(n7198), .A2(n7197), .ZN(n7196) );
  INV_X1 U8610 ( .A(n14009), .ZN(n13878) );
  AND2_X1 U8611 ( .A1(n9300), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9313) );
  NAND2_X1 U8612 ( .A1(n14173), .A2(n7293), .ZN(n13924) );
  AND4_X1 U8613 ( .A1(n9253), .A2(n9252), .A3(n9251), .A4(n9250), .ZN(n13912)
         );
  OR2_X1 U8614 ( .A1(n14169), .A2(n11415), .ZN(n11411) );
  NAND2_X1 U8615 ( .A1(n14173), .A2(n14391), .ZN(n14172) );
  NOR2_X1 U8616 ( .A1(n9230), .A2(n9229), .ZN(n9248) );
  NAND2_X1 U8617 ( .A1(n11358), .A2(n11357), .ZN(n11360) );
  OR2_X1 U8618 ( .A1(n11356), .A2(n11355), .ZN(n11357) );
  AOI21_X1 U8619 ( .B1(n7121), .B2(n7123), .A(n6725), .ZN(n7119) );
  INV_X1 U8620 ( .A(n11421), .ZN(n11359) );
  OR2_X1 U8621 ( .A1(n9213), .A2(n9212), .ZN(n9230) );
  OR2_X1 U8622 ( .A1(n9159), .A2(n9156), .ZN(n9174) );
  OAI21_X1 U8623 ( .B1(n11120), .B2(n7126), .A(n11196), .ZN(n7125) );
  AND2_X1 U8624 ( .A1(n11130), .A2(n6688), .ZN(n7347) );
  AND2_X1 U8625 ( .A1(n14560), .A2(n11123), .ZN(n14543) );
  OAI22_X1 U8626 ( .A1(n11129), .A2(n11128), .B1(n13595), .B2(n11127), .ZN(
        n14548) );
  OR2_X1 U8627 ( .A1(n9130), .A2(n10764), .ZN(n9159) );
  OR2_X1 U8628 ( .A1(n13903), .A2(n13685), .ZN(n10873) );
  AND3_X1 U8629 ( .A1(n6744), .A2(n7352), .A3(n7351), .ZN(n10897) );
  OR2_X1 U8630 ( .A1(n11066), .A2(n10899), .ZN(n10906) );
  NOR2_X1 U8631 ( .A1(n10889), .A2(n11092), .ZN(n7117) );
  AOI21_X1 U8632 ( .B1(n6741), .B2(n11092), .A(n7116), .ZN(n7115) );
  NAND2_X1 U8633 ( .A1(n11091), .A2(n11090), .ZN(n7353) );
  NAND2_X1 U8634 ( .A1(n7292), .A2(n10889), .ZN(n11066) );
  INV_X1 U8635 ( .A(n11085), .ZN(n7292) );
  NAND2_X1 U8636 ( .A1(n6935), .A2(n7286), .ZN(n7285) );
  NAND2_X1 U8637 ( .A1(n10350), .A2(n10295), .ZN(n10296) );
  NAND2_X1 U8638 ( .A1(n10296), .A2(n10307), .ZN(n10886) );
  NAND2_X1 U8639 ( .A1(n13599), .A2(n12178), .ZN(n10303) );
  NAND2_X1 U8640 ( .A1(n10346), .A2(n10353), .ZN(n10350) );
  NAND2_X1 U8641 ( .A1(n11803), .A2(n13698), .ZN(n7182) );
  INV_X1 U8642 ( .A(n11779), .ZN(n7274) );
  NAND2_X1 U8643 ( .A1(n13807), .A2(n11772), .ZN(n13796) );
  NAND2_X1 U8644 ( .A1(n9361), .A2(n9360), .ZN(n13990) );
  NAND2_X1 U8645 ( .A1(n9299), .A2(n9298), .ZN(n14015) );
  OAI21_X1 U8646 ( .B1(n9632), .B2(n9485), .A(n9115), .ZN(n14631) );
  INV_X1 U8647 ( .A(n14632), .ZN(n14665) );
  AND2_X1 U8648 ( .A1(n9793), .A2(n9569), .ZN(n10871) );
  AND2_X1 U8649 ( .A1(n10451), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9569) );
  AND2_X1 U8650 ( .A1(n7590), .A2(n9029), .ZN(n7589) );
  XNOR2_X1 U8651 ( .A(n9483), .B(n9482), .ZN(n13347) );
  NAND2_X1 U8652 ( .A1(n6890), .A2(n8256), .ZN(n9483) );
  OR2_X1 U8653 ( .A1(n8253), .A2(n8252), .ZN(n6890) );
  NOR2_X1 U8654 ( .A1(n7364), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n7362) );
  INV_X1 U8655 ( .A(n7590), .ZN(n7364) );
  XNOR2_X1 U8656 ( .A(n8238), .B(n8224), .ZN(n11830) );
  NAND2_X1 U8657 ( .A1(n6876), .A2(n8170), .ZN(n8173) );
  NAND2_X1 U8658 ( .A1(n8169), .A2(n10647), .ZN(n6876) );
  NAND2_X1 U8659 ( .A1(n8139), .A2(n8138), .ZN(n6886) );
  NAND2_X1 U8660 ( .A1(n6896), .A2(n8120), .ZN(n8125) );
  INV_X1 U8661 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9242) );
  OAI21_X1 U8662 ( .B1(n7932), .B2(n7931), .A(n7930), .ZN(n7950) );
  NAND2_X1 U8663 ( .A1(n7823), .A2(n7822), .ZN(n7839) );
  CLKBUF_X1 U8664 ( .A(n9095), .Z(n9096) );
  INV_X1 U8665 ( .A(n7608), .ZN(n7607) );
  INV_X1 U8666 ( .A(n6937), .ZN(n7767) );
  NAND2_X1 U8667 ( .A1(n7765), .A2(n7764), .ZN(n7768) );
  NAND2_X1 U8668 ( .A1(n7768), .A2(n7767), .ZN(n7784) );
  AND2_X1 U8669 ( .A1(n7034), .A2(n7764), .ZN(n7033) );
  OR2_X1 U8670 ( .A1(n7752), .A2(SI_2_), .ZN(n7034) );
  OAI211_X1 U8671 ( .C1(n6861), .C2(P3_ADDR_REG_3__SCAN_IN), .A(n6859), .B(
        n6858), .ZN(n14085) );
  NAND2_X1 U8672 ( .A1(n6860), .A2(n15493), .ZN(n6859) );
  NAND2_X1 U8673 ( .A1(n6861), .A2(n6720), .ZN(n6858) );
  INV_X1 U8674 ( .A(n7011), .ZN(n6860) );
  XNOR2_X1 U8675 ( .A(n14090), .B(n14055), .ZN(n14091) );
  NOR2_X1 U8676 ( .A1(n14088), .A2(n14089), .ZN(n14092) );
  NAND2_X1 U8677 ( .A1(n6875), .A2(n14096), .ZN(n14098) );
  XOR2_X1 U8678 ( .A(n14059), .B(P3_ADDR_REG_7__SCAN_IN), .Z(n14097) );
  OAI21_X1 U8679 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n15366), .A(n14063), .ZN(
        n14104) );
  OAI21_X1 U8680 ( .B1(n14151), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n6926), .ZN(
        n6925) );
  OAI21_X1 U8681 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n15062), .A(n14070), .ZN(
        n14073) );
  AND2_X1 U8682 ( .A1(n7010), .A2(n7008), .ZN(n14122) );
  NOR2_X1 U8683 ( .A1(n14422), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n14124) );
  AND2_X1 U8684 ( .A1(n8880), .A2(n8879), .ZN(n12355) );
  NAND2_X1 U8685 ( .A1(n11339), .A2(n11338), .ZN(n12244) );
  NAND2_X1 U8686 ( .A1(n11339), .A2(n6648), .ZN(n12245) );
  INV_X1 U8687 ( .A(n7234), .ZN(n12275) );
  OAI21_X1 U8688 ( .B1(n12333), .B2(n7237), .A(n7235), .ZN(n7234) );
  OR2_X1 U8689 ( .A1(n7244), .A2(n7238), .ZN(n7237) );
  INV_X1 U8690 ( .A(n7236), .ZN(n7235) );
  NAND2_X1 U8691 ( .A1(n8848), .A2(n8847), .ZN(n12596) );
  NAND2_X1 U8692 ( .A1(n8900), .A2(n8899), .ZN(n12547) );
  AND2_X1 U8693 ( .A1(n12190), .A2(n7252), .ZN(n7251) );
  NAND2_X1 U8694 ( .A1(n8787), .A2(n8786), .ZN(n12317) );
  INV_X1 U8695 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n12348) );
  NAND2_X1 U8696 ( .A1(n9949), .A2(n9948), .ZN(n12376) );
  INV_X1 U8697 ( .A(n12208), .ZN(n6864) );
  NAND2_X1 U8698 ( .A1(n12209), .A2(n12208), .ZN(n12345) );
  NAND2_X1 U8699 ( .A1(n8860), .A2(n8859), .ZN(n12361) );
  NAND2_X1 U8700 ( .A1(n7259), .A2(n10744), .ZN(n10745) );
  AND4_X1 U8701 ( .A1(n8643), .A2(n8642), .A3(n8641), .A4(n8640), .ZN(n10948)
         );
  INV_X1 U8702 ( .A(n7231), .ZN(n12371) );
  AOI21_X1 U8703 ( .B1(n12333), .B2(n7233), .A(n7232), .ZN(n7231) );
  NOR2_X1 U8704 ( .A1(n7242), .A2(n7241), .ZN(n7233) );
  NOR2_X1 U8705 ( .A1(n7246), .A2(n7242), .ZN(n7232) );
  NAND2_X1 U8706 ( .A1(n7250), .A2(n11493), .ZN(n12191) );
  NAND2_X1 U8707 ( .A1(n11490), .A2(n11489), .ZN(n7250) );
  INV_X1 U8708 ( .A(n11759), .ZN(n7301) );
  AND2_X1 U8709 ( .A1(n11546), .A2(n8951), .ZN(n11554) );
  INV_X1 U8710 ( .A(n12355), .ZN(n12388) );
  INV_X1 U8711 ( .A(n11336), .ZN(n12401) );
  INV_X1 U8712 ( .A(n10948), .ZN(n12403) );
  INV_X1 U8713 ( .A(n10785), .ZN(n12404) );
  INV_X1 U8714 ( .A(n10742), .ZN(n12405) );
  INV_X1 U8715 ( .A(n7391), .ZN(n7390) );
  INV_X1 U8716 ( .A(n15118), .ZN(n12408) );
  OR2_X1 U8717 ( .A1(n9940), .A2(n12773), .ZN(n12410) );
  AOI22_X1 U8718 ( .A1(n14951), .A2(n14952), .B1(n14956), .B2(n9972), .ZN(
        n10817) );
  INV_X1 U8719 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n14989) );
  NOR2_X1 U8720 ( .A1(n14965), .A2(n10800), .ZN(n14976) );
  INV_X1 U8721 ( .A(n7464), .ZN(n15001) );
  INV_X1 U8722 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n15366) );
  INV_X1 U8723 ( .A(n10802), .ZN(n7463) );
  INV_X1 U8724 ( .A(n7341), .ZN(n15008) );
  INV_X1 U8725 ( .A(n7339), .ZN(n15006) );
  INV_X1 U8726 ( .A(n7070), .ZN(n15023) );
  OR2_X1 U8727 ( .A1(n15059), .A2(n15058), .ZN(n15061) );
  NOR2_X1 U8728 ( .A1(n15042), .A2(n12465), .ZN(n15059) );
  INV_X1 U8729 ( .A(n7068), .ZN(n12415) );
  INV_X1 U8730 ( .A(n6997), .ZN(n15076) );
  XNOR2_X1 U8731 ( .A(n7066), .B(n14198), .ZN(n14191) );
  NOR2_X1 U8732 ( .A1(n14191), .A2(n14192), .ZN(n14190) );
  OAI21_X1 U8733 ( .B1(n14191), .B2(n7466), .A(n7065), .ZN(n14208) );
  NAND2_X1 U8734 ( .A1(n7467), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7466) );
  NAND2_X1 U8735 ( .A1(n12421), .A2(n7467), .ZN(n7065) );
  INV_X1 U8736 ( .A(n14209), .ZN(n7467) );
  XNOR2_X1 U8737 ( .A(n12423), .B(n12478), .ZN(n14224) );
  NOR2_X1 U8738 ( .A1(n14224), .A2(n14225), .ZN(n14223) );
  OAI21_X1 U8739 ( .B1(n14217), .B2(n14218), .A(n6979), .ZN(n14236) );
  OR2_X1 U8740 ( .A1(n12446), .A2(n12447), .ZN(n6979) );
  XNOR2_X1 U8741 ( .A(n11529), .B(n11743), .ZN(n12496) );
  NAND2_X1 U8742 ( .A1(n7092), .A2(n7093), .ZN(n12530) );
  NAND2_X1 U8743 ( .A1(n7602), .A2(n6649), .ZN(n12543) );
  NAND2_X1 U8744 ( .A1(n8872), .A2(n8871), .ZN(n12687) );
  NAND2_X1 U8745 ( .A1(n12607), .A2(n8844), .ZN(n12592) );
  NAND2_X1 U8746 ( .A1(n7110), .A2(n7383), .ZN(n12602) );
  NAND2_X1 U8747 ( .A1(n12645), .A2(n7111), .ZN(n7110) );
  NAND2_X1 U8748 ( .A1(n12629), .A2(n11648), .ZN(n12615) );
  NAND2_X1 U8749 ( .A1(n12649), .A2(n8806), .ZN(n12632) );
  NAND2_X1 U8750 ( .A1(n12644), .A2(n11650), .ZN(n12627) );
  NAND2_X1 U8751 ( .A1(n8812), .A2(n8811), .ZN(n12709) );
  OAI21_X1 U8752 ( .B1(n11378), .B2(n7089), .A(n7087), .ZN(n11503) );
  OR2_X1 U8753 ( .A1(n10392), .A2(n15146), .ZN(n15593) );
  INV_X1 U8754 ( .A(n7086), .ZN(n11438) );
  OAI21_X1 U8755 ( .B1(n11378), .B2(n11735), .A(n11630), .ZN(n11439) );
  AOI21_X1 U8756 ( .B1(n11378), .B2(n11630), .A(n7089), .ZN(n7086) );
  NAND2_X1 U8757 ( .A1(n8750), .A2(n8749), .ZN(n11372) );
  NAND2_X1 U8758 ( .A1(n7604), .A2(n8716), .ZN(n14265) );
  NAND2_X1 U8759 ( .A1(n11025), .A2(n7389), .ZN(n14287) );
  NAND2_X1 U8760 ( .A1(n12576), .A2(n11380), .ZN(n15600) );
  NAND2_X1 U8761 ( .A1(n9959), .A2(n9958), .ZN(n14270) );
  NAND2_X1 U8762 ( .A1(n10947), .A2(n8685), .ZN(n10926) );
  NAND2_X1 U8763 ( .A1(n10584), .A2(n11568), .ZN(n10382) );
  INV_X1 U8764 ( .A(n14270), .ZN(n15591) );
  NAND2_X1 U8765 ( .A1(n11540), .A2(n11539), .ZN(n12722) );
  INV_X1 U8766 ( .A(n12343), .ZN(n12755) );
  NAND2_X1 U8767 ( .A1(n8825), .A2(n8824), .ZN(n12759) );
  NAND2_X1 U8768 ( .A1(n8759), .A2(n8758), .ZN(n11474) );
  NAND2_X1 U8769 ( .A1(n9939), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12773) );
  XNOR2_X1 U8770 ( .A(n8921), .B(n8920), .ZN(n11178) );
  NAND2_X1 U8771 ( .A1(n7266), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8479) );
  NAND2_X1 U8772 ( .A1(n7606), .A2(n8753), .ZN(n7266) );
  INV_X1 U8773 ( .A(SI_19_), .ZN(n9965) );
  INV_X1 U8774 ( .A(SI_18_), .ZN(n15288) );
  NAND2_X1 U8775 ( .A1(n7326), .A2(n8415), .ZN(n8768) );
  NAND2_X1 U8776 ( .A1(n8752), .A2(n8751), .ZN(n7326) );
  NAND2_X1 U8777 ( .A1(n8724), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8737) );
  INV_X1 U8778 ( .A(SI_11_), .ZN(n15428) );
  NAND2_X1 U8779 ( .A1(n8695), .A2(n8405), .ZN(n8710) );
  XNOR2_X1 U8780 ( .A(n8698), .B(n8697), .ZN(n15033) );
  OAI21_X1 U8781 ( .B1(n8399), .B2(n7308), .A(n7305), .ZN(n8676) );
  NAND2_X1 U8782 ( .A1(n8663), .A2(n8662), .ZN(n8665) );
  NAND2_X1 U8783 ( .A1(n8399), .A2(n8398), .ZN(n8663) );
  XNOR2_X1 U8784 ( .A(n8646), .B(P3_IR_REG_7__SCAN_IN), .ZN(n14993) );
  NAND2_X1 U8785 ( .A1(n8615), .A2(n8393), .ZN(n8632) );
  XNOR2_X1 U8786 ( .A(n8618), .B(P3_IR_REG_5__SCAN_IN), .ZN(n14962) );
  XNOR2_X1 U8787 ( .A(n8599), .B(P3_IR_REG_4__SCAN_IN), .ZN(n10795) );
  NAND2_X1 U8788 ( .A1(n8584), .A2(n8585), .ZN(n8587) );
  NAND2_X1 U8789 ( .A1(n7313), .A2(n8386), .ZN(n8585) );
  NAND2_X1 U8790 ( .A1(n8550), .A2(n8598), .ZN(n6828) );
  NAND2_X1 U8791 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n8551) );
  OR2_X1 U8792 ( .A1(n8368), .A2(n11335), .ZN(n9643) );
  INV_X1 U8793 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n11405) );
  NAND2_X1 U8794 ( .A1(n7482), .A2(n7481), .ZN(n10692) );
  NAND2_X1 U8795 ( .A1(n7483), .A2(n7486), .ZN(n7481) );
  NAND2_X1 U8796 ( .A1(n10531), .A2(n7479), .ZN(n7482) );
  INV_X1 U8797 ( .A(n10683), .ZN(n7486) );
  NAND2_X1 U8798 ( .A1(n7499), .A2(n11184), .ZN(n11187) );
  NAND2_X1 U8799 ( .A1(n7502), .A2(n7503), .ZN(n12846) );
  NAND2_X1 U8800 ( .A1(n12798), .A2(n12137), .ZN(n12853) );
  NAND2_X1 U8801 ( .A1(n12853), .A2(n12852), .ZN(n12851) );
  NAND2_X1 U8802 ( .A1(n7429), .A2(n9871), .ZN(n9821) );
  NAND2_X1 U8803 ( .A1(n11297), .A2(n11296), .ZN(n11401) );
  NAND2_X1 U8804 ( .A1(n9900), .A2(n9901), .ZN(n9926) );
  OR2_X1 U8805 ( .A1(n7769), .A2(n9600), .ZN(n7653) );
  OR2_X1 U8806 ( .A1(n9610), .A2(n7763), .ZN(n7652) );
  AND2_X1 U8807 ( .A1(n12878), .A2(n7501), .ZN(n7500) );
  AND2_X1 U8808 ( .A1(n7502), .A2(n7501), .ZN(n12879) );
  NAND2_X1 U8809 ( .A1(n12825), .A2(n7535), .ZN(n12884) );
  AND2_X1 U8810 ( .A1(n12825), .A2(n12145), .ZN(n12886) );
  NAND2_X1 U8811 ( .A1(n8271), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6938) );
  XNOR2_X1 U8812 ( .A(n6953), .B(n12983), .ZN(n12099) );
  NAND2_X1 U8813 ( .A1(n6659), .A2(n6713), .ZN(n6953) );
  INV_X1 U8814 ( .A(n12108), .ZN(n6967) );
  NAND2_X1 U8815 ( .A1(n8249), .A2(n8248), .ZN(n12917) );
  INV_X1 U8816 ( .A(n12890), .ZN(n12920) );
  INV_X1 U8817 ( .A(n12983), .ZN(n13195) );
  NAND2_X1 U8818 ( .A1(n13048), .A2(n8334), .ZN(n13038) );
  OAI21_X1 U8819 ( .B1(n13075), .B2(n13058), .A(n7042), .ZN(n13042) );
  NAND2_X1 U8820 ( .A1(n13075), .A2(n8168), .ZN(n13059) );
  NAND2_X1 U8821 ( .A1(n13093), .A2(n8329), .ZN(n13073) );
  NAND2_X1 U8822 ( .A1(n7426), .A2(n7427), .ZN(n13087) );
  NAND2_X1 U8823 ( .A1(n13118), .A2(n8119), .ZN(n13104) );
  NOR2_X1 U8824 ( .A1(n7055), .A2(n8091), .ZN(n13119) );
  NAND2_X1 U8825 ( .A1(n7539), .A2(n12065), .ZN(n13117) );
  NAND2_X1 U8826 ( .A1(n7508), .A2(n8323), .ZN(n13160) );
  NAND2_X1 U8827 ( .A1(n8020), .A2(n8019), .ZN(n13294) );
  NAND2_X1 U8828 ( .A1(n7037), .A2(n7038), .ZN(n11246) );
  NAND2_X1 U8829 ( .A1(n11101), .A2(n7438), .ZN(n11164) );
  NAND2_X1 U8830 ( .A1(n7496), .A2(n7493), .ZN(n11100) );
  INV_X1 U8831 ( .A(n7495), .ZN(n7493) );
  NAND2_X1 U8832 ( .A1(n7498), .A2(n7497), .ZN(n7496) );
  OR2_X1 U8833 ( .A1(n13211), .A2(n10200), .ZN(n14835) );
  NAND2_X1 U8834 ( .A1(n7049), .A2(n7430), .ZN(n10991) );
  NAND2_X1 U8835 ( .A1(n7435), .A2(n7837), .ZN(n10572) );
  NAND2_X1 U8836 ( .A1(n10601), .A2(n12075), .ZN(n7435) );
  NAND2_X1 U8837 ( .A1(n7537), .A2(n8304), .ZN(n10397) );
  INV_X1 U8838 ( .A(n13213), .ZN(n14315) );
  OR2_X1 U8839 ( .A1(n10201), .A2(n13195), .ZN(n13213) );
  INV_X1 U8840 ( .A(n13182), .ZN(n14316) );
  NAND2_X1 U8841 ( .A1(n14881), .A2(n9813), .ZN(n13194) );
  INV_X1 U8842 ( .A(n14835), .ZN(n14307) );
  NAND2_X1 U8843 ( .A1(n7429), .A2(n11846), .ZN(n14884) );
  INV_X1 U8844 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n7225) );
  INV_X1 U8845 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n7542) );
  INV_X1 U8846 ( .A(n13319), .ZN(n13248) );
  NAND2_X1 U8847 ( .A1(n8128), .A2(n8127), .ZN(n13270) );
  OR2_X1 U8848 ( .A1(n10999), .A2(n8209), .ZN(n8128) );
  AND2_X1 U8849 ( .A1(n14934), .A2(n14892), .ZN(n13304) );
  INV_X1 U8850 ( .A(n13224), .ZN(n13312) );
  OR2_X1 U8851 ( .A1(n14924), .A2(n8246), .ZN(n7447) );
  NAND2_X1 U8852 ( .A1(n7450), .A2(n14905), .ZN(n7449) );
  INV_X1 U8853 ( .A(n13066), .ZN(n13323) );
  INV_X1 U8854 ( .A(n11870), .ZN(n10378) );
  AND2_X2 U8855 ( .A1(n8978), .A2(n9808), .ZN(n14924) );
  NOR2_X1 U8856 ( .A1(n14849), .A2(n14879), .ZN(n14872) );
  CLKBUF_X1 U8857 ( .A(n14872), .Z(n14876) );
  NOR2_X1 U8858 ( .A1(n9930), .A2(P2_U3088), .ZN(n14881) );
  NOR2_X1 U8859 ( .A1(P2_IR_REG_29__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n7446) );
  OAI21_X1 U8860 ( .B1(n8271), .B2(P2_IR_REG_20__SCAN_IN), .A(n8270), .ZN(
        n8275) );
  NOR2_X1 U8861 ( .A1(n7143), .A2(n8273), .ZN(n8274) );
  NOR2_X1 U8862 ( .A1(n8269), .A2(n8268), .ZN(n8270) );
  INV_X1 U8863 ( .A(n8342), .ZN(n12066) );
  INV_X1 U8864 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n15311) );
  INV_X1 U8865 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10521) );
  INV_X1 U8866 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10091) );
  INV_X1 U8867 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9888) );
  INV_X1 U8868 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9743) );
  INV_X1 U8869 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9705) );
  INV_X1 U8870 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9635) );
  INV_X1 U8871 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9630) );
  INV_X1 U8872 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9613) );
  XNOR2_X1 U8873 ( .A(n9557), .B(n9556), .ZN(n9793) );
  OAI21_X1 U8874 ( .B1(n9555), .B2(P1_IR_REG_22__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9557) );
  INV_X1 U8875 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n10764) );
  INV_X1 U8876 ( .A(n13474), .ZN(n6981) );
  NAND2_X1 U8877 ( .A1(n14343), .A2(n14344), .ZN(n14342) );
  NAND2_X1 U8878 ( .A1(n9247), .A2(n9246), .ZN(n14383) );
  CLKBUF_X1 U8879 ( .A(n14349), .Z(n14351) );
  AOI21_X1 U8880 ( .B1(n7551), .B2(n7553), .A(n7549), .ZN(n7548) );
  INV_X1 U8881 ( .A(n13465), .ZN(n7549) );
  NAND2_X1 U8882 ( .A1(n7547), .A2(n7551), .ZN(n13466) );
  OR2_X1 U8883 ( .A1(n13517), .A2(n7553), .ZN(n7547) );
  NAND2_X1 U8884 ( .A1(n11008), .A2(n11007), .ZN(n11010) );
  NAND2_X1 U8885 ( .A1(n9057), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9049) );
  OR2_X1 U8886 ( .A1(n13437), .A2(n13436), .ZN(n6999) );
  NAND2_X1 U8887 ( .A1(n9415), .A2(n9414), .ZN(n13965) );
  NAND2_X1 U8888 ( .A1(n11388), .A2(n11387), .ZN(n11394) );
  NAND2_X1 U8889 ( .A1(n13488), .A2(n7569), .ZN(n13541) );
  NAND2_X1 U8890 ( .A1(n13516), .A2(n13404), .ZN(n13550) );
  INV_X1 U8891 ( .A(n14365), .ZN(n13573) );
  OR2_X1 U8892 ( .A1(n9491), .A2(n10117), .ZN(n9060) );
  NAND2_X1 U8893 ( .A1(n13634), .A2(n13635), .ZN(n13633) );
  NAND2_X1 U8894 ( .A1(n13647), .A2(n13648), .ZN(n13646) );
  INV_X1 U8895 ( .A(n7211), .ZN(n10238) );
  NOR2_X1 U8896 ( .A1(n10177), .A2(n6695), .ZN(n10167) );
  NOR2_X1 U8897 ( .A1(n10167), .A2(n10166), .ZN(n10165) );
  AOI21_X1 U8898 ( .B1(n10183), .B2(P1_REG1_REG_6__SCAN_IN), .A(n10180), .ZN(
        n10170) );
  NOR2_X1 U8899 ( .A1(n10165), .A2(n7204), .ZN(n10227) );
  AND2_X1 U8900 ( .A1(n10171), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7204) );
  NOR2_X1 U8901 ( .A1(n10227), .A2(n10226), .ZN(n10225) );
  NAND2_X1 U8902 ( .A1(n10219), .A2(n6948), .ZN(n10206) );
  OR2_X1 U8903 ( .A1(n10222), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6948) );
  NAND2_X1 U8904 ( .A1(n10206), .A2(n10207), .ZN(n10205) );
  NOR2_X1 U8905 ( .A1(n10212), .A2(n7206), .ZN(n10126) );
  AND2_X1 U8906 ( .A1(n10208), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7206) );
  NOR2_X1 U8907 ( .A1(n10126), .A2(n10125), .ZN(n10423) );
  NOR2_X1 U8908 ( .A1(n14490), .A2(n14489), .ZN(n14488) );
  AND2_X1 U8909 ( .A1(n10139), .A2(n10124), .ZN(n14521) );
  AOI21_X1 U8910 ( .B1(n12012), .B2(n9488), .A(n9487), .ZN(n13935) );
  INV_X1 U8911 ( .A(n7182), .ZN(n13939) );
  NAND2_X1 U8912 ( .A1(n13726), .A2(n11778), .ZN(n13715) );
  AOI21_X1 U8913 ( .B1(n13707), .B2(n14554), .A(n13706), .ZN(n13949) );
  NAND2_X1 U8914 ( .A1(n13752), .A2(n7684), .ZN(n13732) );
  INV_X1 U8915 ( .A(n13792), .ZN(n13774) );
  AND2_X1 U8916 ( .A1(n13770), .A2(n11792), .ZN(n7349) );
  NAND2_X1 U8917 ( .A1(n7350), .A2(n11792), .ZN(n13773) );
  NAND2_X1 U8918 ( .A1(n13801), .A2(n11790), .ZN(n13787) );
  NAND2_X1 U8919 ( .A1(n11769), .A2(n11768), .ZN(n13839) );
  NAND2_X1 U8920 ( .A1(n13849), .A2(n7355), .ZN(n13835) );
  NAND2_X1 U8921 ( .A1(n13849), .A2(n11787), .ZN(n13833) );
  NAND2_X1 U8922 ( .A1(n7176), .A2(n7178), .ZN(n13885) );
  NAND2_X1 U8923 ( .A1(n7177), .A2(n7357), .ZN(n7176) );
  NAND2_X1 U8924 ( .A1(n13917), .A2(n11782), .ZN(n13897) );
  NOR2_X1 U8925 ( .A1(n11426), .A2(n6809), .ZN(n6808) );
  INV_X1 U8926 ( .A(n11425), .ZN(n6809) );
  NAND2_X1 U8927 ( .A1(n6810), .A2(n11425), .ZN(n11427) );
  NAND2_X1 U8928 ( .A1(n11262), .A2(n11261), .ZN(n11264) );
  NAND2_X1 U8929 ( .A1(n11258), .A2(n7189), .ZN(n7120) );
  NOR2_X1 U8930 ( .A1(n14532), .A2(n7682), .ZN(n11209) );
  INV_X1 U8931 ( .A(n14658), .ZN(n14541) );
  NAND2_X1 U8932 ( .A1(n14550), .A2(n11120), .ZN(n7124) );
  INV_X1 U8933 ( .A(n14631), .ZN(n11127) );
  NAND2_X1 U8934 ( .A1(n11084), .A2(n10888), .ZN(n11065) );
  INV_X1 U8935 ( .A(n14557), .ZN(n14573) );
  INV_X1 U8936 ( .A(n13857), .ZN(n14569) );
  INV_X1 U8937 ( .A(n13896), .ZN(n14175) );
  INV_X1 U8938 ( .A(n14688), .ZN(n14686) );
  INV_X1 U8939 ( .A(n6806), .ZN(n13954) );
  AND2_X1 U8940 ( .A1(n9568), .A2(n9567), .ZN(n9992) );
  OAI211_X1 U8941 ( .C1(n9504), .C2(n7627), .A(n7622), .B(n7625), .ZN(n13339)
         );
  OR2_X1 U8942 ( .A1(n9026), .A2(n8998), .ZN(n9012) );
  CLKBUF_X1 U8943 ( .A(n9570), .Z(n9571) );
  NAND2_X1 U8944 ( .A1(n8223), .A2(n8208), .ZN(n14041) );
  NAND2_X1 U8945 ( .A1(n8204), .A2(n8222), .ZN(n8207) );
  INV_X1 U8946 ( .A(n9992), .ZN(n11463) );
  XNOR2_X1 U8947 ( .A(n9563), .B(P1_IR_REG_24__SCAN_IN), .ZN(n11331) );
  NAND2_X1 U8948 ( .A1(n7135), .A2(n9009), .ZN(n9562) );
  XNOR2_X1 U8949 ( .A(n8158), .B(SI_23_), .ZN(n11308) );
  OR2_X1 U8950 ( .A1(n8999), .A2(n8998), .ZN(n9000) );
  INV_X1 U8951 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11827) );
  MUX2_X1 U8952 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8995), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n8997) );
  NAND2_X1 U8953 ( .A1(n8991), .A2(n7421), .ZN(n8994) );
  NAND2_X1 U8954 ( .A1(n6895), .A2(n8120), .ZN(n8121) );
  NAND2_X1 U8955 ( .A1(n8120), .A2(n8103), .ZN(n8106) );
  NAND2_X1 U8956 ( .A1(n8071), .A2(n8058), .ZN(n10723) );
  INV_X1 U8957 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n15494) );
  INV_X1 U8958 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10519) );
  INV_X1 U8959 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9886) );
  INV_X1 U8960 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9788) );
  OAI21_X1 U8961 ( .B1(n7880), .B2(n7882), .A(n6990), .ZN(n7905) );
  NOR2_X1 U8962 ( .A1(n6991), .A2(n7904), .ZN(n6990) );
  NAND2_X1 U8963 ( .A1(n7884), .A2(n7883), .ZN(n7901) );
  NAND2_X1 U8964 ( .A1(n7880), .A2(n7879), .ZN(n7884) );
  INV_X1 U8965 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9740) );
  INV_X1 U8966 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9706) );
  INV_X1 U8967 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9636) );
  INV_X1 U8968 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9631) );
  AND2_X1 U8969 ( .A1(n7190), .A2(n7191), .ZN(n7806) );
  AND2_X1 U8970 ( .A1(n7586), .A2(n7588), .ZN(n9077) );
  AND2_X1 U8971 ( .A1(n9064), .A2(n7587), .ZN(n7586) );
  XNOR2_X1 U8972 ( .A(n7209), .B(n9064), .ZN(n13630) );
  OR2_X1 U8973 ( .A1(n9063), .A2(n8998), .ZN(n7209) );
  AND2_X1 U8974 ( .A1(n7588), .A2(n7587), .ZN(n9063) );
  NAND2_X1 U8975 ( .A1(n7765), .A2(n7032), .ZN(n9610) );
  OR2_X1 U8976 ( .A1(n7033), .A2(n7035), .ZN(n7032) );
  NAND2_X1 U8977 ( .A1(n6893), .A2(n7749), .ZN(n7751) );
  INV_X1 U8978 ( .A(n6894), .ZN(n6893) );
  INV_X1 U8979 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n14079) );
  XNOR2_X1 U8980 ( .A(n14080), .B(n6970), .ZN(n15615) );
  INV_X1 U8981 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6970) );
  AOI21_X1 U8982 ( .B1(n14084), .B2(n14083), .A(n14140), .ZN(n15611) );
  NAND2_X1 U8983 ( .A1(n6871), .A2(n14103), .ZN(n14149) );
  NAND2_X1 U8984 ( .A1(n14146), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n6871) );
  INV_X1 U8985 ( .A(n7020), .ZN(n14101) );
  OAI21_X1 U8986 ( .B1(n14413), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n6698), .ZN(
        n7022) );
  NOR2_X1 U8987 ( .A1(n14414), .A2(n6870), .ZN(n14420) );
  AOI21_X1 U8988 ( .B1(n14416), .B2(n14415), .A(P2_ADDR_REG_13__SCAN_IN), .ZN(
        n6870) );
  OR2_X1 U8989 ( .A1(n14420), .A2(n14419), .ZN(n7010) );
  AND2_X1 U8990 ( .A1(n14122), .A2(n14123), .ZN(n14422) );
  AND2_X1 U8991 ( .A1(n7017), .A2(n7016), .ZN(n14178) );
  INV_X1 U8992 ( .A(n14132), .ZN(n6923) );
  INV_X1 U8993 ( .A(n14426), .ZN(n7015) );
  OR2_X1 U8994 ( .A1(n11758), .A2(n11757), .ZN(n7299) );
  INV_X1 U8995 ( .A(n7454), .ZN(n12413) );
  OR2_X1 U8996 ( .A1(n14252), .A2(n6995), .ZN(P3_U3200) );
  OAI21_X1 U8997 ( .B1(n14254), .B2(n15110), .A(n6797), .ZN(n6995) );
  OR2_X1 U8998 ( .A1(n12484), .A2(n15110), .ZN(n6957) );
  NOR2_X1 U8999 ( .A1(n12482), .A2(n7345), .ZN(n7344) );
  INV_X1 U9000 ( .A(n6899), .ZN(n6898) );
  OAI21_X1 U9001 ( .B1(n12732), .B2(n12721), .A(n6900), .ZN(n6899) );
  OR2_X1 U9002 ( .A1(n15202), .A2(n12669), .ZN(n6900) );
  NOR2_X1 U9003 ( .A1(n6777), .A2(n6974), .ZN(n6973) );
  NOR2_X1 U9004 ( .A1(n15181), .A2(n9585), .ZN(n6974) );
  INV_X1 U9005 ( .A(n6902), .ZN(n6901) );
  OAI22_X1 U9006 ( .A1(n12732), .A2(n12771), .B1(n15181), .B2(n12731), .ZN(
        n6902) );
  NAND2_X1 U9007 ( .A1(n7484), .A2(n10529), .ZN(n10685) );
  AOI21_X1 U9008 ( .B1(n13309), .B2(n14934), .A(n7223), .ZN(n13225) );
  NAND2_X1 U9009 ( .A1(n7226), .A2(n7224), .ZN(n7223) );
  OR2_X1 U9010 ( .A1(n14934), .A2(n7225), .ZN(n7224) );
  NAND2_X1 U9011 ( .A1(n7543), .A2(n7540), .ZN(P2_U3527) );
  AOI21_X1 U9012 ( .B1(n13229), .B2(n13304), .A(n7541), .ZN(n7540) );
  NAND2_X1 U9013 ( .A1(n13313), .A2(n14934), .ZN(n7543) );
  NOR2_X1 U9014 ( .A1(n14934), .A2(n7542), .ZN(n7541) );
  AOI21_X1 U9015 ( .B1(n12022), .B2(n8982), .A(n8981), .ZN(n8983) );
  NAND2_X1 U9016 ( .A1(n7448), .A2(n6921), .ZN(P2_U3495) );
  INV_X1 U9017 ( .A(n6922), .ZN(n6921) );
  NAND2_X1 U9018 ( .A1(n13313), .A2(n14924), .ZN(n7448) );
  OAI21_X1 U9019 ( .B1(n7221), .B2(n13329), .A(n7447), .ZN(n6922) );
  XNOR2_X1 U9020 ( .A(n6976), .B(n6975), .ZN(n13562) );
  NAND2_X1 U9021 ( .A1(n14671), .A2(n14675), .ZN(n7272) );
  INV_X1 U9022 ( .A(n7271), .ZN(n7270) );
  OAI21_X1 U9023 ( .B1(n7276), .B2(n14673), .A(n7275), .ZN(n7271) );
  INV_X1 U9024 ( .A(n6926), .ZN(n14152) );
  AND2_X1 U9025 ( .A1(n7178), .A2(n13884), .ZN(n6644) );
  OR2_X1 U9026 ( .A1(n11198), .A2(n13593), .ZN(n6645) );
  OR2_X1 U9027 ( .A1(n11662), .A2(n11649), .ZN(n6646) );
  OR2_X1 U9028 ( .A1(n12460), .A2(n12459), .ZN(n6647) );
  AND2_X1 U9029 ( .A1(n7265), .A2(n11338), .ZN(n6648) );
  AND2_X1 U9030 ( .A1(n7601), .A2(n8896), .ZN(n6649) );
  OR2_X1 U9031 ( .A1(n8959), .A2(n11720), .ZN(n6650) );
  AND2_X1 U9032 ( .A1(n12633), .A2(n11650), .ZN(n6651) );
  XNOR2_X1 U9033 ( .A(n13232), .B(n12918), .ZN(n13020) );
  INV_X1 U9034 ( .A(n13020), .ZN(n8336) );
  XOR2_X1 U9035 ( .A(n7097), .B(n9966), .Z(n6652) );
  XNOR2_X1 U9036 ( .A(n6830), .B(n14198), .ZN(n14195) );
  MUX2_X1 U9037 ( .A(P2_IR_REG_0__SCAN_IN), .B(n13361), .S(n7742), .Z(n14882)
         );
  INV_X1 U9038 ( .A(n14882), .ZN(n7214) );
  AND2_X1 U9039 ( .A1(n14367), .A2(n13570), .ZN(n6653) );
  AND2_X1 U9040 ( .A1(n11919), .A2(n12934), .ZN(n6654) );
  AND3_X1 U9041 ( .A1(n6645), .A2(n11118), .A3(n11121), .ZN(n6655) );
  AND2_X1 U9042 ( .A1(n7505), .A2(n12833), .ZN(n6656) );
  AND2_X1 U9043 ( .A1(n7663), .A2(n7662), .ZN(n6657) );
  AND2_X1 U9044 ( .A1(n14043), .A2(n9043), .ZN(n13812) );
  INV_X1 U9045 ( .A(n13812), .ZN(n13983) );
  AND2_X1 U9046 ( .A1(n8226), .A2(n8225), .ZN(n13019) );
  INV_X1 U9047 ( .A(n13019), .ZN(n13232) );
  AND2_X1 U9048 ( .A1(n13893), .A2(n13585), .ZN(n6658) );
  XOR2_X1 U9049 ( .A(n13312), .B(n12915), .Z(n6659) );
  AND2_X1 U9050 ( .A1(n7096), .A2(n7094), .ZN(n6660) );
  AND2_X1 U9051 ( .A1(n11323), .A2(n11314), .ZN(n6661) );
  AND2_X1 U9052 ( .A1(n7230), .A2(n7229), .ZN(n6662) );
  AND2_X1 U9053 ( .A1(n12401), .A2(n11139), .ZN(n6663) );
  INV_X1 U9054 ( .A(n12076), .ZN(n10571) );
  NAND2_X1 U9055 ( .A1(n9509), .A2(n9508), .ZN(n13695) );
  INV_X1 U9056 ( .A(n13695), .ZN(n6998) );
  INV_X1 U9057 ( .A(n11717), .ZN(n7374) );
  NOR2_X1 U9058 ( .A1(n11890), .A2(n7858), .ZN(n6664) );
  AND2_X1 U9059 ( .A1(n7041), .A2(n13045), .ZN(n6665) );
  AND2_X1 U9060 ( .A1(n11009), .A2(n11007), .ZN(n6666) );
  AND2_X1 U9061 ( .A1(n6806), .A2(n6805), .ZN(n6667) );
  NOR2_X1 U9062 ( .A1(n7358), .A2(n7359), .ZN(n7357) );
  OAI21_X1 U9063 ( .B1(n13908), .B2(n6779), .A(n11762), .ZN(n13883) );
  INV_X1 U9064 ( .A(n10878), .ZN(n13685) );
  NAND2_X1 U9065 ( .A1(n7977), .A2(n7976), .ZN(n14308) );
  INV_X1 U9066 ( .A(n14308), .ZN(n7218) );
  OR2_X1 U9067 ( .A1(n8200), .A2(SI_25_), .ZN(n6668) );
  AND2_X1 U9068 ( .A1(n7625), .A2(n7623), .ZN(n6669) );
  NAND2_X1 U9069 ( .A1(n7348), .A2(n7347), .ZN(n11206) );
  AND2_X1 U9070 ( .A1(n6668), .A2(SI_26_), .ZN(n6670) );
  AND2_X1 U9071 ( .A1(n7459), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n6671) );
  INV_X1 U9072 ( .A(n9082), .ZN(n9343) );
  AND3_X1 U9073 ( .A1(n9047), .A2(n9046), .A3(n9045), .ZN(n6672) );
  NAND2_X1 U9074 ( .A1(n13133), .A2(n8092), .ZN(n7059) );
  NAND2_X1 U9075 ( .A1(n11915), .A2(n11908), .ZN(n6673) );
  OAI211_X1 U9076 ( .C1(n8551), .C2(n8550), .A(n8552), .B(n6828), .ZN(n9836)
         );
  NOR2_X1 U9077 ( .A1(n8724), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n8753) );
  INV_X1 U9078 ( .A(n12224), .ZN(n7241) );
  CLKBUF_X3 U9079 ( .A(n10014), .Z(n13445) );
  XNOR2_X1 U9080 ( .A(n13066), .B(n12827), .ZN(n13058) );
  AND2_X1 U9081 ( .A1(n8010), .A2(n8006), .ZN(n6674) );
  OR2_X1 U9082 ( .A1(n8343), .A2(n8342), .ZN(n10195) );
  INV_X1 U9083 ( .A(n13943), .ZN(n13709) );
  NAND2_X1 U9084 ( .A1(n9460), .A2(n9459), .ZN(n13943) );
  XNOR2_X1 U9085 ( .A(n8588), .B(P3_IR_REG_3__SCAN_IN), .ZN(n14956) );
  AND2_X1 U9086 ( .A1(n8189), .A2(n8188), .ZN(n13319) );
  XNOR2_X1 U9087 ( .A(n6938), .B(P2_IR_REG_20__SCAN_IN), .ZN(n8342) );
  INV_X1 U9088 ( .A(n11208), .ZN(n7189) );
  NOR2_X1 U9089 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n7588) );
  NAND2_X1 U9090 ( .A1(n8545), .A2(n8544), .ZN(n12513) );
  NAND2_X1 U9091 ( .A1(n7605), .A2(n7382), .ZN(n8474) );
  XNOR2_X1 U9092 ( .A(n12022), .B(n8267), .ZN(n12096) );
  OR2_X1 U9093 ( .A1(n14993), .A2(n10807), .ZN(n6675) );
  AND2_X1 U9094 ( .A1(n13759), .A2(n7291), .ZN(n6676) );
  AND2_X1 U9095 ( .A1(n13090), .A2(n8151), .ZN(n6677) );
  OR2_X1 U9096 ( .A1(n14423), .A2(n7018), .ZN(n6678) );
  AND2_X1 U9097 ( .A1(n13094), .A2(n8327), .ZN(n6679) );
  AND2_X1 U9098 ( .A1(n7374), .A2(n11681), .ZN(n6680) );
  NAND2_X1 U9099 ( .A1(n9433), .A2(n9432), .ZN(n13957) );
  AND2_X1 U9100 ( .A1(n11933), .A2(n11932), .ZN(n6681) );
  NAND4_X1 U9101 ( .A1(n7717), .A2(n7715), .A3(n7714), .A4(n7716), .ZN(n11843)
         );
  NOR2_X1 U9102 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n9039) );
  INV_X1 U9103 ( .A(n10302), .ZN(n10304) );
  OR2_X1 U9104 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n14098), .ZN(n6682) );
  NAND2_X1 U9105 ( .A1(n8076), .A2(n8075), .ZN(n8271) );
  INV_X1 U9106 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n15493) );
  OR2_X1 U9107 ( .A1(n15074), .A2(n12419), .ZN(n6683) );
  AND2_X1 U9108 ( .A1(n13051), .A2(n7220), .ZN(n6684) );
  NOR2_X1 U9109 ( .A1(n14329), .A2(n7948), .ZN(n6685) );
  AND2_X1 U9110 ( .A1(n11648), .A2(n11653), .ZN(n12633) );
  AND2_X1 U9111 ( .A1(n12113), .A2(n12112), .ZN(n6686) );
  AND2_X1 U9112 ( .A1(n12404), .A2(n11141), .ZN(n6687) );
  OR2_X1 U9113 ( .A1(n13594), .A2(n14642), .ZN(n6688) );
  INV_X1 U9114 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6989) );
  INV_X1 U9115 ( .A(n7151), .ZN(n7150) );
  NAND2_X1 U9116 ( .A1(n7153), .A2(n6788), .ZN(n7151) );
  XOR2_X1 U9117 ( .A(n13935), .B(n13577), .Z(n6689) );
  AND2_X1 U9118 ( .A1(n6823), .A2(n6821), .ZN(n6690) );
  AND4_X1 U9119 ( .A1(n12095), .A2(n12094), .A3(n13020), .A4(n13037), .ZN(
        n6691) );
  NOR2_X1 U9120 ( .A1(n13422), .A2(n13423), .ZN(n7570) );
  NAND2_X1 U9121 ( .A1(n13837), .A2(n11770), .ZN(n13817) );
  OR2_X1 U9122 ( .A1(n15074), .A2(n12470), .ZN(n6692) );
  NAND2_X1 U9123 ( .A1(n9284), .A2(n9283), .ZN(n14367) );
  INV_X1 U9124 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n12778) );
  NOR2_X1 U9125 ( .A1(n9981), .A2(n14956), .ZN(n9986) );
  NAND2_X1 U9126 ( .A1(n9239), .A2(n9238), .ZN(n14169) );
  AND2_X1 U9127 ( .A1(n8328), .A2(n8327), .ZN(n13092) );
  OR3_X1 U9128 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n6693) );
  OR2_X1 U9129 ( .A1(n11876), .A2(n12940), .ZN(n6694) );
  AND2_X1 U9130 ( .A1(n10183), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6695) );
  INV_X1 U9131 ( .A(n11371), .ZN(n11735) );
  INV_X1 U9132 ( .A(n9189), .ZN(n7415) );
  INV_X1 U9133 ( .A(n9241), .ZN(n7410) );
  AND2_X1 U9134 ( .A1(n11976), .A2(n11975), .ZN(n6696) );
  AND2_X1 U9135 ( .A1(n12101), .A2(n12062), .ZN(n6697) );
  NAND2_X1 U9136 ( .A1(n8062), .A2(n8061), .ZN(n13283) );
  OR2_X1 U9137 ( .A1(n14116), .A2(n14115), .ZN(n6698) );
  AND2_X1 U9138 ( .A1(n7289), .A2(n7288), .ZN(n6699) );
  INV_X1 U9139 ( .A(n7244), .ZN(n7243) );
  NAND2_X1 U9140 ( .A1(n7246), .A2(n7245), .ZN(n7244) );
  NAND2_X1 U9141 ( .A1(n10097), .A2(n10096), .ZN(n6700) );
  AND2_X1 U9142 ( .A1(n11883), .A2(n11882), .ZN(n6701) );
  AND2_X1 U9143 ( .A1(n11615), .A2(n11616), .ZN(n14290) );
  AND2_X1 U9144 ( .A1(n11340), .A2(n12400), .ZN(n6702) );
  AND2_X1 U9145 ( .A1(n11937), .A2(n11936), .ZN(n6703) );
  OR2_X1 U9146 ( .A1(n12709), .A2(n12324), .ZN(n11648) );
  NOR2_X1 U9147 ( .A1(n14190), .A2(n12421), .ZN(n6704) );
  NOR2_X1 U9148 ( .A1(n14193), .A2(n12474), .ZN(n6705) );
  NOR2_X1 U9149 ( .A1(n14223), .A2(n12424), .ZN(n6706) );
  NOR2_X1 U9150 ( .A1(n12114), .A2(n7165), .ZN(n6707) );
  INV_X1 U9151 ( .A(n7296), .ZN(n13818) );
  NOR2_X1 U9152 ( .A1(n13841), .A2(n13990), .ZN(n7296) );
  AND2_X1 U9153 ( .A1(n7365), .A2(n7366), .ZN(n6708) );
  AND2_X1 U9154 ( .A1(n12565), .A2(n11681), .ZN(n6709) );
  NAND2_X1 U9155 ( .A1(n14329), .A2(n12933), .ZN(n6710) );
  INV_X1 U9156 ( .A(n14375), .ZN(n13925) );
  NAND2_X1 U9157 ( .A1(n9258), .A2(n9257), .ZN(n14375) );
  AND2_X1 U9158 ( .A1(n8211), .A2(n8210), .ZN(n13036) );
  INV_X1 U9159 ( .A(n13036), .ZN(n13238) );
  AND2_X1 U9160 ( .A1(n11777), .A2(n11776), .ZN(n6711) );
  AND2_X1 U9161 ( .A1(n11185), .A2(n11184), .ZN(n6712) );
  INV_X1 U9162 ( .A(n8313), .ZN(n7497) );
  AND2_X1 U9163 ( .A1(n6954), .A2(n6691), .ZN(n6713) );
  AND2_X1 U9164 ( .A1(n6662), .A2(n13330), .ZN(n6714) );
  AND2_X1 U9165 ( .A1(n12607), .A2(n7597), .ZN(n6715) );
  OR2_X1 U9166 ( .A1(n12230), .A2(n12387), .ZN(n6716) );
  INV_X1 U9167 ( .A(n7155), .ZN(n7154) );
  NAND2_X1 U9168 ( .A1(n7156), .A2(n7157), .ZN(n7155) );
  OR2_X1 U9169 ( .A1(n11989), .A2(n11988), .ZN(n6717) );
  AND2_X1 U9170 ( .A1(n9044), .A2(n9042), .ZN(n6718) );
  AND2_X1 U9171 ( .A1(n13270), .A2(n11982), .ZN(n6719) );
  INV_X1 U9172 ( .A(n7357), .ZN(n7179) );
  INV_X1 U9173 ( .A(n7143), .ZN(n8277) );
  NOR2_X1 U9174 ( .A1(n8059), .A2(n8272), .ZN(n7143) );
  AND2_X1 U9175 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n7011), .ZN(n6720) );
  AND2_X1 U9176 ( .A1(n13036), .A2(n12828), .ZN(n6721) );
  INV_X1 U9177 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8598) );
  NAND2_X1 U9178 ( .A1(n9980), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n6722) );
  NAND2_X1 U9179 ( .A1(n11744), .A2(n12722), .ZN(n6723) );
  OAI21_X1 U9180 ( .B1(n6680), .B2(n7372), .A(n11689), .ZN(n7371) );
  INV_X1 U9181 ( .A(n7051), .ZN(n7050) );
  NOR2_X1 U9182 ( .A1(n14909), .A2(n12937), .ZN(n7051) );
  NOR2_X1 U9183 ( .A1(n13979), .A2(n13582), .ZN(n6724) );
  NOR2_X1 U9184 ( .A1(n11356), .A2(n13590), .ZN(n6725) );
  NOR2_X1 U9185 ( .A1(n12596), .A2(n12390), .ZN(n6726) );
  XOR2_X1 U9186 ( .A(P3_ADDR_REG_19__SCAN_IN), .B(n14186), .Z(n6727) );
  OR2_X1 U9187 ( .A1(n11801), .A2(n11779), .ZN(n6728) );
  OR2_X1 U9188 ( .A1(n11934), .A2(n11245), .ZN(n6729) );
  INV_X1 U9189 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8269) );
  AND2_X1 U9190 ( .A1(n7602), .A2(n8896), .ZN(n6730) );
  AND2_X1 U9191 ( .A1(n12547), .A2(n12373), .ZN(n6731) );
  INV_X1 U9192 ( .A(n13923), .ZN(n13918) );
  AND2_X1 U9193 ( .A1(n7952), .A2(n15490), .ZN(n6732) );
  NOR2_X1 U9194 ( .A1(n13473), .A2(n13472), .ZN(n6733) );
  NOR2_X1 U9195 ( .A1(n14329), .A2(n12933), .ZN(n6734) );
  NAND2_X1 U9196 ( .A1(n7605), .A2(n8753), .ZN(n6735) );
  INV_X1 U9197 ( .A(n7057), .ZN(n7056) );
  NAND2_X1 U9198 ( .A1(n7058), .A2(n13120), .ZN(n7057) );
  AND2_X1 U9199 ( .A1(n11995), .A2(n11994), .ZN(n6736) );
  AND2_X1 U9200 ( .A1(n12148), .A2(n12147), .ZN(n6737) );
  INV_X1 U9201 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n7363) );
  INV_X1 U9202 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9614) );
  NAND2_X1 U9203 ( .A1(n12270), .A2(n12502), .ZN(n6738) );
  AND2_X1 U9204 ( .A1(n9886), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n6739) );
  NAND2_X1 U9205 ( .A1(n11594), .A2(n11598), .ZN(n6740) );
  AND2_X1 U9206 ( .A1(n11689), .A2(n11692), .ZN(n12542) );
  INV_X1 U9207 ( .A(n12542), .ZN(n7601) );
  INV_X1 U9208 ( .A(n7257), .ZN(n7256) );
  NAND2_X1 U9209 ( .A1(n7258), .A2(n10744), .ZN(n7257) );
  NAND2_X1 U9210 ( .A1(n10888), .A2(n11072), .ZN(n6741) );
  INV_X1 U9211 ( .A(n12114), .ZN(n7166) );
  AND2_X1 U9212 ( .A1(n12095), .A2(n8235), .ZN(n7436) );
  OR2_X1 U9213 ( .A1(n13229), .A2(n12793), .ZN(n8251) );
  NAND2_X1 U9214 ( .A1(n8991), .A2(n7420), .ZN(n8996) );
  NAND2_X1 U9215 ( .A1(n8243), .A2(n8242), .ZN(n13229) );
  INV_X1 U9216 ( .A(n13229), .ZN(n7221) );
  OR2_X1 U9217 ( .A1(n9642), .A2(n9686), .ZN(n6742) );
  AND2_X1 U9218 ( .A1(n11598), .A2(n11599), .ZN(n11720) );
  INV_X1 U9219 ( .A(n10889), .ZN(n11072) );
  AND3_X1 U9220 ( .A1(n9081), .A2(n9080), .A3(n9079), .ZN(n10889) );
  OR2_X1 U9221 ( .A1(n11895), .A2(n7878), .ZN(n6743) );
  OR2_X1 U9222 ( .A1(n10867), .A2(n10889), .ZN(n6744) );
  OR2_X1 U9223 ( .A1(n14188), .A2(n14187), .ZN(n6745) );
  OR2_X1 U9224 ( .A1(n14092), .A2(n14091), .ZN(n6746) );
  OR2_X1 U9225 ( .A1(n6773), .A2(n11983), .ZN(n6747) );
  AND2_X1 U9226 ( .A1(n11865), .A2(n11864), .ZN(n6748) );
  AND4_X1 U9227 ( .A1(n9021), .A2(n9020), .A3(n9019), .A4(n9018), .ZN(n10351)
         );
  OR2_X1 U9228 ( .A1(n11974), .A2(n6752), .ZN(n6749) );
  AND2_X1 U9229 ( .A1(n11875), .A2(n11874), .ZN(n6750) );
  AND2_X1 U9230 ( .A1(n7093), .A2(n11688), .ZN(n6751) );
  AND2_X1 U9231 ( .A1(n11971), .A2(n11970), .ZN(n6752) );
  INV_X1 U9232 ( .A(n10152), .ZN(n13599) );
  AND2_X1 U9233 ( .A1(n7293), .A2(n13515), .ZN(n6753) );
  AND2_X1 U9234 ( .A1(n7038), .A2(n6729), .ZN(n6754) );
  OR2_X1 U9235 ( .A1(n11751), .A2(n11716), .ZN(n6755) );
  OR2_X1 U9236 ( .A1(n11887), .A2(n6701), .ZN(n6756) );
  INV_X1 U9237 ( .A(n8308), .ZN(n7515) );
  INV_X1 U9238 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7719) );
  INV_X1 U9239 ( .A(n7783), .ZN(n7609) );
  NAND2_X1 U9240 ( .A1(n7766), .A2(SI_3_), .ZN(n7783) );
  INV_X1 U9241 ( .A(n11261), .ZN(n7186) );
  INV_X1 U9242 ( .A(n11121), .ZN(n7126) );
  AND2_X1 U9243 ( .A1(n7420), .A2(n7419), .ZN(n6757) );
  INV_X1 U9244 ( .A(n7043), .ZN(n7042) );
  OAI21_X1 U9245 ( .B1(n13058), .B2(n8168), .A(n8185), .ZN(n7043) );
  OR2_X1 U9246 ( .A1(n9364), .A2(n9362), .ZN(n6758) );
  NAND2_X1 U9247 ( .A1(n12119), .A2(n12118), .ZN(n6759) );
  OR2_X1 U9248 ( .A1(n9142), .A2(n9140), .ZN(n6760) );
  INV_X1 U9249 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7703) );
  INV_X1 U9250 ( .A(n8394), .ZN(n7323) );
  AND2_X1 U9251 ( .A1(n7248), .A2(n6716), .ZN(n6761) );
  OR2_X1 U9252 ( .A1(n7415), .A2(n9188), .ZN(n6762) );
  AND2_X1 U9253 ( .A1(n7589), .A2(n7284), .ZN(n6763) );
  OR2_X1 U9254 ( .A1(n9240), .A2(n7410), .ZN(n6764) );
  OR2_X1 U9255 ( .A1(n7660), .A2(n6736), .ZN(n6765) );
  INV_X1 U9256 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9029) );
  NAND2_X1 U9257 ( .A1(n11951), .A2(n11952), .ZN(n6766) );
  NAND2_X1 U9258 ( .A1(n9462), .A2(n7402), .ZN(n6767) );
  INV_X1 U9259 ( .A(n13728), .ZN(n11777) );
  AND2_X1 U9260 ( .A1(n11797), .A2(n9534), .ZN(n13728) );
  INV_X1 U9261 ( .A(n7571), .ZN(n7568) );
  NAND2_X1 U9262 ( .A1(n13418), .A2(n13419), .ZN(n7571) );
  INV_X1 U9263 ( .A(n7570), .ZN(n7569) );
  NAND2_X1 U9264 ( .A1(n8258), .A2(n8257), .ZN(n12022) );
  INV_X1 U9265 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n8990) );
  OR2_X1 U9266 ( .A1(n6681), .A2(n7671), .ZN(n6768) );
  NAND2_X1 U9267 ( .A1(n9406), .A2(n7395), .ZN(n6769) );
  NAND2_X1 U9268 ( .A1(n9435), .A2(n7405), .ZN(n6770) );
  INV_X1 U9269 ( .A(n7490), .ZN(n7489) );
  NAND2_X1 U9270 ( .A1(n7492), .A2(n6710), .ZN(n7490) );
  INV_X1 U9271 ( .A(n7108), .ZN(n7107) );
  NAND2_X1 U9272 ( .A1(n7383), .A2(n7109), .ZN(n7108) );
  INV_X1 U9273 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9599) );
  INV_X2 U9274 ( .A(n8829), .ZN(n8654) );
  INV_X1 U9275 ( .A(n13884), .ZN(n7346) );
  INV_X1 U9276 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n6827) );
  NAND2_X1 U9277 ( .A1(n6810), .A2(n6808), .ZN(n7679) );
  AND2_X1 U9278 ( .A1(n14173), .A2(n7295), .ZN(n6771) );
  INV_X1 U9279 ( .A(n12604), .ZN(n7109) );
  INV_X1 U9280 ( .A(SI_1_), .ZN(n6891) );
  INV_X1 U9281 ( .A(n15015), .ZN(n10808) );
  XNOR2_X1 U9282 ( .A(n8661), .B(P3_IR_REG_8__SCAN_IN), .ZN(n15015) );
  AND2_X1 U9283 ( .A1(n12123), .A2(n12122), .ZN(n6772) );
  NAND3_X1 U9284 ( .A1(n8989), .A2(n7680), .A3(n7688), .ZN(n9254) );
  INV_X1 U9285 ( .A(n9254), .ZN(n7135) );
  AND2_X1 U9286 ( .A1(n11980), .A2(n11979), .ZN(n6773) );
  AND2_X1 U9287 ( .A1(n11954), .A2(n11953), .ZN(n6774) );
  NOR2_X1 U9288 ( .A1(n12344), .A2(n6864), .ZN(n6775) );
  INV_X1 U9289 ( .A(n11651), .ZN(n12647) );
  AND2_X1 U9290 ( .A1(n8819), .A2(n8806), .ZN(n6776) );
  AND2_X1 U9291 ( .A1(n8941), .A2(n9586), .ZN(n6777) );
  AND2_X1 U9292 ( .A1(n13917), .A2(n7357), .ZN(n6778) );
  NOR2_X1 U9293 ( .A1(n14367), .A2(n13914), .ZN(n6779) );
  INV_X1 U9294 ( .A(n13404), .ZN(n7556) );
  AND2_X1 U9295 ( .A1(n13431), .A2(n13430), .ZN(n6780) );
  AND2_X1 U9296 ( .A1(n7110), .A2(n7107), .ZN(n6781) );
  AND2_X1 U9297 ( .A1(n8753), .A2(n8456), .ZN(n8471) );
  AND2_X1 U9298 ( .A1(n10519), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n6782) );
  AND2_X1 U9299 ( .A1(n8101), .A2(n9965), .ZN(n6783) );
  AND2_X1 U9300 ( .A1(n13866), .A2(n11785), .ZN(n6784) );
  INV_X1 U9301 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n7392) );
  AND2_X1 U9302 ( .A1(n7693), .A2(n8380), .ZN(n6785) );
  NAND2_X1 U9303 ( .A1(n7702), .A2(n7866), .ZN(n8059) );
  INV_X1 U9304 ( .A(n13785), .ZN(n6805) );
  INV_X1 U9305 ( .A(n11783), .ZN(n7359) );
  NAND2_X1 U9306 ( .A1(n7656), .A2(n7655), .ZN(n8355) );
  AND2_X1 U9307 ( .A1(n9502), .A2(SI_30_), .ZN(n6786) );
  AND2_X1 U9308 ( .A1(n12418), .A2(n15074), .ZN(n6787) );
  NAND2_X1 U9309 ( .A1(n8962), .A2(n11621), .ZN(n14259) );
  NAND2_X1 U9310 ( .A1(n7124), .A2(n11121), .ZN(n11197) );
  NAND2_X1 U9311 ( .A1(n7120), .A2(n11259), .ZN(n11354) );
  OR2_X1 U9312 ( .A1(n12125), .A2(n12124), .ZN(n6788) );
  NAND2_X1 U9313 ( .A1(n8109), .A2(n8108), .ZN(n13273) );
  INV_X1 U9314 ( .A(n13273), .ZN(n7229) );
  AND2_X1 U9315 ( .A1(n9506), .A2(n6786), .ZN(n6789) );
  OR2_X1 U9316 ( .A1(n6889), .A2(n8252), .ZN(n6790) );
  OR2_X1 U9317 ( .A1(n8059), .A2(n7706), .ZN(n6791) );
  NAND2_X1 U9318 ( .A1(n11315), .A2(n11314), .ZN(n11321) );
  INV_X1 U9319 ( .A(n8209), .ZN(n12011) );
  INV_X1 U9320 ( .A(n7260), .ZN(n12774) );
  OAI21_X1 U9321 ( .B1(n8494), .B2(P3_D_REG_0__SCAN_IN), .A(n8499), .ZN(n7260)
         );
  AND2_X1 U9322 ( .A1(n11025), .A2(n8961), .ZN(n6792) );
  AND2_X1 U9323 ( .A1(n7259), .A2(n7256), .ZN(n6793) );
  AND2_X1 U9324 ( .A1(n7454), .A2(n7455), .ZN(n6794) );
  AND2_X1 U9325 ( .A1(n7464), .A2(n7463), .ZN(n6795) );
  AND2_X1 U9326 ( .A1(n15063), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n6796) );
  NAND2_X1 U9327 ( .A1(n11252), .A2(n14325), .ZN(n14311) );
  INV_X1 U9328 ( .A(n14311), .ZN(n7219) );
  NOR2_X1 U9329 ( .A1(n14253), .A2(n6996), .ZN(n6797) );
  AND2_X1 U9330 ( .A1(n7048), .A2(n7050), .ZN(n6798) );
  INV_X1 U9331 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n7707) );
  AND2_X1 U9332 ( .A1(n7348), .A2(n6688), .ZN(n6799) );
  AND2_X1 U9333 ( .A1(n6978), .A2(n6647), .ZN(n6800) );
  NAND2_X1 U9334 ( .A1(n7173), .A2(n12983), .ZN(n9870) );
  INV_X1 U9335 ( .A(n12075), .ZN(n7431) );
  INV_X1 U9336 ( .A(n9503), .ZN(n7628) );
  BUF_X1 U9337 ( .A(n11854), .Z(n9920) );
  INV_X1 U9338 ( .A(n9920), .ZN(n7215) );
  NAND2_X1 U9339 ( .A1(n9835), .A2(n12452), .ZN(n15095) );
  NAND2_X1 U9340 ( .A1(n9926), .A2(n9925), .ZN(n10092) );
  AND2_X1 U9341 ( .A1(n6823), .A2(n6822), .ZN(n6801) );
  AND2_X1 U9342 ( .A1(n14551), .A2(n14636), .ZN(n14018) );
  AND2_X1 U9343 ( .A1(n9484), .A2(n12786), .ZN(n6802) );
  AND2_X1 U9344 ( .A1(n7354), .A2(n7353), .ZN(n6803) );
  AND2_X1 U9345 ( .A1(n10081), .A2(n10029), .ZN(n6804) );
  XNOR2_X1 U9346 ( .A(n8510), .B(P3_IR_REG_19__SCAN_IN), .ZN(n12483) );
  INV_X1 U9347 ( .A(n12483), .ZN(n9966) );
  INV_X1 U9348 ( .A(n12480), .ZN(n14243) );
  NAND2_X1 U9349 ( .A1(n7337), .A2(n9983), .ZN(n9973) );
  INV_X1 U9350 ( .A(n9973), .ZN(n9974) );
  INV_X1 U9351 ( .A(n13630), .ZN(n7286) );
  INV_X1 U9352 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7545) );
  INV_X1 U9353 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7012) );
  INV_X1 U9354 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7546) );
  INV_X1 U9355 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7476) );
  OR2_X1 U9356 ( .A1(n15054), .A2(n15074), .ZN(n7458) );
  OR2_X1 U9357 ( .A1(n12418), .A2(n15074), .ZN(n7459) );
  NAND4_X1 U9358 ( .A1(n6812), .A2(n8985), .A3(n6811), .A4(n9064), .ZN(n9095)
         );
  NAND3_X1 U9359 ( .A1(n7135), .A2(n7137), .A3(n9009), .ZN(n6813) );
  NAND2_X1 U9360 ( .A1(n10886), .A2(n10885), .ZN(n11082) );
  NAND2_X1 U9361 ( .A1(n13883), .A2(n11763), .ZN(n6814) );
  NAND2_X1 U9362 ( .A1(n10806), .A2(n14962), .ZN(n6822) );
  INV_X1 U9363 ( .A(n9851), .ZN(n14936) );
  NAND2_X1 U9364 ( .A1(n9830), .A2(n6826), .ZN(n9831) );
  NAND2_X1 U9365 ( .A1(n9836), .A2(n9851), .ZN(n6826) );
  INV_X1 U9366 ( .A(n6831), .ZN(n14995) );
  XNOR2_X1 U9367 ( .A(n10807), .B(n14993), .ZN(n14996) );
  NAND2_X1 U9368 ( .A1(n6832), .A2(n6835), .ZN(n11873) );
  NAND2_X1 U9369 ( .A1(n6837), .A2(n6836), .ZN(n6832) );
  OAI211_X1 U9370 ( .C1(n6837), .C2(n6834), .A(n6833), .B(n7662), .ZN(n7661)
         );
  NAND2_X1 U9371 ( .A1(n11867), .A2(n6835), .ZN(n6833) );
  INV_X1 U9372 ( .A(n6835), .ZN(n6834) );
  OAI21_X1 U9373 ( .B1(n6969), .B2(n6696), .A(n6839), .ZN(n6842) );
  NAND3_X1 U9374 ( .A1(n6842), .A2(n6747), .A3(n6841), .ZN(n7666) );
  INV_X1 U9375 ( .A(n11938), .ZN(n6845) );
  NAND2_X1 U9376 ( .A1(n6846), .A2(n7659), .ZN(n11999) );
  NAND3_X1 U9377 ( .A1(n6850), .A2(n6847), .A3(n6765), .ZN(n6846) );
  NAND2_X1 U9378 ( .A1(n6849), .A2(n6848), .ZN(n6847) );
  NAND2_X1 U9379 ( .A1(n6852), .A2(n6851), .ZN(n6850) );
  NAND2_X1 U9380 ( .A1(n6853), .A2(n11993), .ZN(n6852) );
  NAND2_X1 U9381 ( .A1(n6992), .A2(n6717), .ZN(n6853) );
  AND2_X2 U9382 ( .A1(n7701), .A2(n7745), .ZN(n7866) );
  NAND2_X1 U9383 ( .A1(n7672), .A2(n7673), .ZN(n6857) );
  OAI21_X1 U9384 ( .B1(n6862), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n14053), .ZN(
        n14054) );
  NAND2_X1 U9385 ( .A1(n12366), .A2(n12201), .ZN(n12204) );
  NAND2_X1 U9386 ( .A1(n12323), .A2(n12320), .ZN(n6863) );
  NAND2_X1 U9387 ( .A1(n6925), .A2(n6917), .ZN(n6868) );
  NAND2_X1 U9388 ( .A1(n14410), .A2(n14411), .ZN(n14409) );
  AND2_X4 U9389 ( .A1(n10027), .A2(n6869), .ZN(n12220) );
  NAND2_X4 U9390 ( .A1(n8504), .A2(n8503), .ZN(n11559) );
  NAND2_X1 U9391 ( .A1(n11452), .A2(n11483), .ZN(n6873) );
  OAI21_X1 U9392 ( .B1(n11452), .B2(n11483), .A(n11451), .ZN(n6874) );
  INV_X1 U9393 ( .A(n7023), .ZN(n14093) );
  NAND2_X1 U9394 ( .A1(n14145), .A2(n14144), .ZN(n6875) );
  XNOR2_X1 U9395 ( .A(n7023), .B(P2_ADDR_REG_6__SCAN_IN), .ZN(n14145) );
  NAND2_X1 U9396 ( .A1(n7635), .A2(n6877), .ZN(n6880) );
  NAND2_X1 U9397 ( .A1(n8139), .A2(n6884), .ZN(n6883) );
  XNOR2_X1 U9398 ( .A(n6886), .B(SI_22_), .ZN(n9372) );
  NAND2_X1 U9399 ( .A1(n7819), .A2(n7818), .ZN(n7823) );
  NAND3_X1 U9400 ( .A1(n7190), .A2(n7191), .A3(n7805), .ZN(n7819) );
  INV_X1 U9401 ( .A(SI_26_), .ZN(n11136) );
  NAND2_X1 U9402 ( .A1(n8778), .A2(n11732), .ZN(n11507) );
  AOI21_X1 U9403 ( .B1(n12536), .B2(n8919), .A(n8918), .ZN(n12517) );
  NAND2_X1 U9404 ( .A1(n10386), .A2(n8593), .ZN(n10507) );
  OAI21_X1 U9405 ( .B1(n12730), .B2(n8976), .A(n6898), .ZN(P3_U3487) );
  OAI21_X1 U9406 ( .B1(n12730), .B2(n15183), .A(n6901), .ZN(P3_U3455) );
  NAND2_X1 U9407 ( .A1(n10692), .A2(n10691), .ZN(n10775) );
  INV_X1 U9408 ( .A(n10093), .ZN(n10098) );
  NAND2_X1 U9409 ( .A1(n7163), .A2(n12114), .ZN(n7162) );
  OAI21_X2 U9410 ( .B1(n12798), .B2(n7142), .A(n7140), .ZN(n12824) );
  NAND3_X1 U9411 ( .A1(n6904), .A2(n6903), .A3(n6764), .ZN(n7408) );
  NAND2_X1 U9412 ( .A1(n9228), .A2(n9227), .ZN(n6903) );
  NAND2_X1 U9413 ( .A1(n9224), .A2(n9223), .ZN(n6904) );
  OR2_X1 U9414 ( .A1(n9497), .A2(n7399), .ZN(n7398) );
  NAND2_X1 U9415 ( .A1(n7401), .A2(n7400), .ZN(n9476) );
  NAND2_X1 U9416 ( .A1(n7404), .A2(n7403), .ZN(n9448) );
  NAND2_X1 U9417 ( .A1(n7394), .A2(n7393), .ZN(n9418) );
  OR3_X2 U9418 ( .A1(n9519), .A2(n9522), .A3(n9520), .ZN(n7689) );
  NAND2_X1 U9419 ( .A1(n9127), .A2(n9126), .ZN(n9128) );
  AOI21_X1 U9420 ( .B1(n9322), .B2(n9321), .A(n6942), .ZN(n9323) );
  BUF_X4 U9421 ( .A(n9108), .Z(n9473) );
  NAND2_X1 U9422 ( .A1(n7765), .A2(n6910), .ZN(n7191) );
  NAND2_X1 U9423 ( .A1(n12012), .A2(n12011), .ZN(n6905) );
  NAND2_X1 U9424 ( .A1(n7785), .A2(SI_4_), .ZN(n7801) );
  NAND2_X1 U9425 ( .A1(n6906), .A2(n7644), .ZN(n8102) );
  NAND2_X1 U9426 ( .A1(n8052), .A2(n7645), .ZN(n6906) );
  NAND2_X1 U9427 ( .A1(n9042), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n6988) );
  INV_X1 U9428 ( .A(n7786), .ZN(n7787) );
  NAND2_X1 U9429 ( .A1(n7843), .A2(n7842), .ZN(n7860) );
  NAND2_X1 U9430 ( .A1(n7617), .A2(n7616), .ZN(n7615) );
  NAND2_X1 U9431 ( .A1(n6937), .A2(n7783), .ZN(n6936) );
  NAND2_X1 U9432 ( .A1(n7839), .A2(n7838), .ZN(n7843) );
  NAND2_X1 U9433 ( .A1(n8035), .A2(n8034), .ZN(n8052) );
  NAND3_X1 U9434 ( .A1(n13728), .A2(n7366), .A3(n7365), .ZN(n13718) );
  XNOR2_X1 U9435 ( .A(n6911), .B(n13685), .ZN(n9553) );
  INV_X1 U9436 ( .A(n9551), .ZN(n6913) );
  NAND2_X1 U9437 ( .A1(n8979), .A2(n14934), .ZN(n7044) );
  INV_X1 U9438 ( .A(n14411), .ZN(n6917) );
  INV_X1 U9439 ( .A(n6925), .ZN(n14410) );
  NOR2_X1 U9440 ( .A1(n14179), .A2(n6918), .ZN(n14188) );
  AOI21_X2 U9441 ( .B1(n13457), .B2(n13458), .A(n6780), .ZN(n13523) );
  NOR2_X2 U9442 ( .A1(n13563), .A2(n6920), .ZN(n13508) );
  NAND2_X1 U9443 ( .A1(n10469), .A2(n10468), .ZN(n10547) );
  NAND2_X1 U9444 ( .A1(n12171), .A2(n10157), .ZN(n10158) );
  NAND2_X1 U9445 ( .A1(n6934), .A2(n10151), .ZN(n12172) );
  OAI21_X1 U9446 ( .B1(n10550), .B2(n7561), .A(n7559), .ZN(n7562) );
  NAND2_X2 U9447 ( .A1(n6643), .A2(n10021), .ZN(n13405) );
  OAI21_X1 U9448 ( .B1(n11899), .B2(n11898), .A(n7677), .ZN(n6987) );
  NAND2_X1 U9449 ( .A1(n10590), .A2(n8592), .ZN(n10386) );
  NOR2_X1 U9450 ( .A1(n7113), .A2(n11749), .ZN(n7112) );
  OAI21_X1 U9451 ( .B1(n9584), .B2(n8976), .A(n8977), .ZN(P3_U3488) );
  OAI21_X1 U9452 ( .B1(n9584), .B2(n15183), .A(n6973), .ZN(P3_U3456) );
  NOR2_X1 U9453 ( .A1(n11710), .A2(n7317), .ZN(n7316) );
  NAND2_X1 U9454 ( .A1(n6998), .A2(n13694), .ZN(n9511) );
  INV_X1 U9455 ( .A(n12093), .ZN(n13045) );
  INV_X1 U9456 ( .A(n7530), .ZN(n7529) );
  INV_X1 U9457 ( .A(n13228), .ZN(n7450) );
  NAND3_X1 U9458 ( .A1(n7449), .A2(n13227), .A3(n13226), .ZN(n13313) );
  AOI21_X1 U9459 ( .B1(n7016), .B2(n7015), .A(n6923), .ZN(n14179) );
  NAND2_X1 U9460 ( .A1(n12048), .A2(n6924), .ZN(n12050) );
  NAND2_X1 U9461 ( .A1(n12025), .A2(n12041), .ZN(n12048) );
  XNOR2_X1 U9462 ( .A(n14188), .B(n14187), .ZN(n14189) );
  NAND2_X1 U9463 ( .A1(n12517), .A2(n12518), .ZN(n12516) );
  OAI21_X1 U9464 ( .B1(n12055), .B2(n7630), .A(n7629), .ZN(n12101) );
  OAI21_X1 U9465 ( .B1(n11897), .B2(n6987), .A(n7675), .ZN(n11924) );
  NAND2_X1 U9466 ( .A1(n6928), .A2(n6927), .ZN(n7007) );
  AOI21_X1 U9467 ( .B1(n6956), .B2(n9973), .A(n6955), .ZN(n10805) );
  NAND3_X1 U9468 ( .A1(n11946), .A2(n7007), .A3(n6766), .ZN(n6931) );
  NAND2_X1 U9469 ( .A1(n6931), .A2(n7004), .ZN(n11957) );
  NAND3_X1 U9470 ( .A1(n11693), .A2(n11741), .A3(n11692), .ZN(n11696) );
  AOI21_X1 U9471 ( .B1(n11581), .B2(n6933), .A(n6932), .ZN(n11593) );
  AOI21_X1 U9472 ( .B1(n11574), .B2(n6984), .A(n6983), .ZN(n11576) );
  AOI21_X1 U9473 ( .B1(n6994), .B2(n6993), .A(n11743), .ZN(n11710) );
  NOR2_X1 U9474 ( .A1(n7316), .A2(n7315), .ZN(n7314) );
  AOI21_X1 U9475 ( .B1(n12432), .B2(n12431), .A(n12430), .ZN(n15027) );
  AOI21_X1 U9476 ( .B1(n12440), .B2(n15074), .A(n15079), .ZN(n15107) );
  AOI21_X1 U9477 ( .B1(n12437), .B2(n12464), .A(n15045), .ZN(n15068) );
  NAND3_X1 U9478 ( .A1(n6958), .A2(n7344), .A3(n6957), .ZN(P3_U3201) );
  NAND2_X1 U9479 ( .A1(n10148), .A2(n10149), .ZN(n6934) );
  NAND2_X1 U9480 ( .A1(n6977), .A2(n10017), .ZN(n10016) );
  NAND2_X1 U9481 ( .A1(n11008), .A2(n6666), .ZN(n11220) );
  INV_X1 U9482 ( .A(n8991), .ZN(n9306) );
  NOR2_X2 U9483 ( .A1(n13566), .A2(n13565), .ZN(n13563) );
  AND2_X1 U9484 ( .A1(n9053), .A2(n9054), .ZN(n7138) );
  NOR2_X1 U9485 ( .A1(n14426), .A2(n14132), .ZN(n7017) );
  INV_X1 U9486 ( .A(n7022), .ZN(n14416) );
  XNOR2_X1 U9487 ( .A(n14092), .B(n14091), .ZN(n15607) );
  OAI21_X1 U9488 ( .B1(n14189), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n6745), .ZN(
        n7021) );
  NAND2_X1 U9489 ( .A1(n6946), .A2(n6945), .ZN(n7669) );
  INV_X1 U9490 ( .A(n11929), .ZN(n6951) );
  NAND2_X1 U9491 ( .A1(n11974), .A2(n6752), .ZN(n7674) );
  MUX2_X1 U9492 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(P2_DATAO_REG_0__SCAN_IN), 
        .S(n9042), .Z(n7731) );
  AND2_X4 U9493 ( .A1(n7618), .A2(n7615), .ZN(n9042) );
  NOR2_X1 U9494 ( .A1(n6657), .A2(n6750), .ZN(n6965) );
  NAND2_X1 U9495 ( .A1(n6941), .A2(n7411), .ZN(n9376) );
  NAND3_X1 U9496 ( .A1(n9353), .A2(n9352), .A3(n6758), .ZN(n6941) );
  NAND2_X1 U9497 ( .A1(n9379), .A2(n9378), .ZN(n9380) );
  OAI21_X1 U9498 ( .B1(n8898), .B2(n8440), .A(n8441), .ZN(n8907) );
  NAND2_X1 U9499 ( .A1(n8868), .A2(n8867), .ZN(n8870) );
  NAND2_X1 U9500 ( .A1(n7319), .A2(n7321), .ZN(n8645) );
  NAND2_X1 U9501 ( .A1(n7304), .A2(n7302), .ZN(n8678) );
  INV_X1 U9502 ( .A(n11705), .ZN(n6993) );
  NAND2_X1 U9503 ( .A1(n6963), .A2(n7301), .ZN(n7300) );
  NAND3_X1 U9504 ( .A1(n6950), .A2(n7669), .A3(n6768), .ZN(n7668) );
  NAND2_X1 U9505 ( .A1(n7072), .A2(n9982), .ZN(n7071) );
  NAND2_X1 U9506 ( .A1(n9853), .A2(n9852), .ZN(n9855) );
  NAND2_X1 U9507 ( .A1(n8552), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8573) );
  AOI21_X1 U9508 ( .B1(P3_REG1_REG_4__SCAN_IN), .B2(n10814), .A(n10805), .ZN(
        n10806) );
  NOR2_X2 U9509 ( .A1(n10797), .A2(n14962), .ZN(n10800) );
  CLKBUF_X2 U9510 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n14044) );
  NAND2_X1 U9511 ( .A1(n9041), .A2(n9040), .ZN(n10128) );
  NOR2_X1 U9512 ( .A1(n7710), .A2(n7446), .ZN(n7445) );
  NAND2_X1 U9513 ( .A1(n11848), .A2(n11847), .ZN(n11857) );
  NAND2_X1 U9514 ( .A1(n6952), .A2(n6951), .ZN(n6950) );
  NAND2_X1 U9515 ( .A1(n11842), .A2(n12058), .ZN(n12027) );
  INV_X1 U9516 ( .A(n11891), .ZN(n7002) );
  OAI22_X1 U9517 ( .A1(n11857), .A2(n11856), .B1(n11859), .B2(n11858), .ZN(
        n11863) );
  NAND2_X1 U9518 ( .A1(n11851), .A2(n12027), .ZN(n11852) );
  OAI211_X1 U9519 ( .C1(n7214), .C2(n12051), .A(n11844), .B(n6985), .ZN(n11848) );
  NAND2_X1 U9520 ( .A1(n11931), .A2(n11930), .ZN(n6952) );
  NAND2_X1 U9521 ( .A1(n8125), .A2(n8124), .ZN(n8139) );
  INV_X1 U9522 ( .A(n7291), .ZN(n7290) );
  OAI21_X1 U9523 ( .B1(n14018), .B2(n13942), .A(n7276), .ZN(n14022) );
  OAI21_X1 U9524 ( .B1(n12101), .B2(n8342), .A(n12100), .ZN(n12107) );
  INV_X1 U9525 ( .A(n14947), .ZN(n6956) );
  NAND2_X1 U9526 ( .A1(n7067), .A2(n14966), .ZN(n6958) );
  NAND2_X1 U9527 ( .A1(n12630), .A2(n8834), .ZN(n12603) );
  NAND2_X4 U9528 ( .A1(n10013), .A2(n10451), .ZN(n13407) );
  NOR2_X2 U9529 ( .A1(n7136), .A2(n9254), .ZN(n9564) );
  NAND2_X1 U9530 ( .A1(n8439), .A2(n8438), .ZN(n8898) );
  AOI21_X1 U9531 ( .B1(n7305), .B2(n7308), .A(n7303), .ZN(n7302) );
  NAND2_X1 U9532 ( .A1(n8870), .A2(n8435), .ZN(n8437) );
  NAND3_X1 U9533 ( .A1(n7112), .A2(n7114), .A3(n6755), .ZN(n6963) );
  NAND2_X1 U9534 ( .A1(n8907), .A2(n8906), .ZN(n8443) );
  NAND2_X1 U9535 ( .A1(n8420), .A2(n8419), .ZN(n8796) );
  NAND2_X1 U9536 ( .A1(n7298), .A2(n8425), .ZN(n8821) );
  NAND2_X1 U9537 ( .A1(n8857), .A2(n8433), .ZN(n8868) );
  NAND2_X1 U9538 ( .A1(n7331), .A2(n7330), .ZN(n8718) );
  NAND2_X1 U9539 ( .A1(n7585), .A2(n7581), .ZN(n7580) );
  XNOR2_X1 U9540 ( .A(n6982), .B(n6981), .ZN(n13456) );
  OAI21_X2 U9541 ( .B1(n8835), .B2(P2_DATAO_REG_20__SCAN_IN), .A(n8428), .ZN(
        n8846) );
  INV_X1 U9542 ( .A(n11866), .ZN(n7003) );
  NAND2_X1 U9543 ( .A1(n6964), .A2(n11879), .ZN(n11881) );
  NAND2_X1 U9544 ( .A1(n7661), .A2(n6965), .ZN(n6964) );
  INV_X4 U9545 ( .A(n12027), .ZN(n12031) );
  NAND4_X2 U9546 ( .A1(n7702), .A2(n7423), .A3(n7866), .A4(n7705), .ZN(n7654)
         );
  OAI211_X1 U9547 ( .C1(n6697), .C2(n6966), .A(n12107), .B(n12106), .ZN(
        P2_U3328) );
  OAI21_X1 U9548 ( .B1(n12101), .B2(n12063), .A(n6967), .ZN(n6966) );
  NAND3_X1 U9549 ( .A1(n11969), .A2(n11968), .A3(n6749), .ZN(n6969) );
  NAND2_X1 U9550 ( .A1(n14077), .A2(n14078), .ZN(n7013) );
  XNOR2_X1 U9551 ( .A(n7021), .B(n6727), .ZN(SUB_1596_U4) );
  NAND2_X1 U9552 ( .A1(n11841), .A2(n7045), .ZN(n8979) );
  NAND2_X1 U9553 ( .A1(n7608), .A2(n7801), .ZN(n7190) );
  NAND2_X1 U9554 ( .A1(n7044), .A2(n6785), .ZN(P2_U3528) );
  NAND2_X1 U9555 ( .A1(n7592), .A2(n7591), .ZN(n11027) );
  NAND2_X1 U9556 ( .A1(n7605), .A2(n7375), .ZN(n8463) );
  NAND2_X1 U9557 ( .A1(n7580), .A2(n7582), .ZN(n6982) );
  NAND2_X1 U9558 ( .A1(n7550), .A2(n7548), .ZN(n13464) );
  OAI211_X1 U9559 ( .C1(n12038), .C2(n7632), .A(n12050), .B(n7631), .ZN(n7630)
         );
  NAND2_X1 U9560 ( .A1(n15012), .A2(n15013), .ZN(n10825) );
  NAND2_X1 U9561 ( .A1(n14990), .A2(n10821), .ZN(n15012) );
  NAND2_X1 U9562 ( .A1(n6692), .A2(n6997), .ZN(n15092) );
  NAND2_X1 U9563 ( .A1(n8505), .A2(n8507), .ZN(n8501) );
  NAND2_X1 U9564 ( .A1(n11706), .A2(n12507), .ZN(n6994) );
  AND2_X4 U9565 ( .A1(n7713), .A2(n7712), .ZN(n7997) );
  NAND2_X1 U9566 ( .A1(n7523), .A2(n7708), .ZN(n7709) );
  NAND2_X1 U9567 ( .A1(n8275), .A2(n8274), .ZN(n8343) );
  AOI21_X1 U9568 ( .B1(n11989), .B2(n11988), .A(n11986), .ZN(n11987) );
  NOR2_X1 U9569 ( .A1(n10195), .A2(n12983), .ZN(n11842) );
  INV_X1 U9570 ( .A(n7676), .ZN(n7675) );
  INV_X1 U9571 ( .A(n11987), .ZN(n6992) );
  NAND2_X1 U9572 ( .A1(n8991), .A2(n9307), .ZN(n9001) );
  INV_X1 U9573 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9607) );
  XNOR2_X2 U9574 ( .A(n12670), .B(n12502), .ZN(n12518) );
  XNOR2_X1 U9575 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8553) );
  NAND2_X1 U9576 ( .A1(n8780), .A2(n8417), .ZN(n8420) );
  NAND2_X1 U9577 ( .A1(n8796), .A2(n8421), .ZN(n8423) );
  NAND2_X1 U9578 ( .A1(n8855), .A2(n8854), .ZN(n8857) );
  NAND2_X1 U9579 ( .A1(n7300), .A2(n7299), .ZN(P3_U3296) );
  AOI21_X1 U9580 ( .B1(n7318), .B2(n7314), .A(n11744), .ZN(n11715) );
  NAND2_X2 U9581 ( .A1(n7864), .A2(n7863), .ZN(n7880) );
  NAND4_X1 U9582 ( .A1(n7689), .A2(n9531), .A3(n9554), .A4(n9532), .ZN(n9560)
         );
  OAI21_X2 U9583 ( .B1(n13523), .B2(n13524), .A(n6999), .ZN(n13498) );
  NAND2_X2 U9584 ( .A1(n13507), .A2(n13397), .ZN(n13517) );
  NAND2_X1 U9585 ( .A1(n7563), .A2(n7564), .ZN(n13540) );
  NOR2_X1 U9586 ( .A1(n14228), .A2(n14227), .ZN(n14226) );
  NAND2_X1 U9587 ( .A1(n15092), .A2(n12471), .ZN(n15097) );
  NAND2_X1 U9588 ( .A1(n7784), .A2(n7783), .ZN(n7788) );
  AOI21_X1 U9589 ( .B1(n11999), .B2(n12000), .A(n11997), .ZN(n11998) );
  INV_X1 U9590 ( .A(n7010), .ZN(n14418) );
  NAND2_X1 U9591 ( .A1(n7009), .A2(n14117), .ZN(n7008) );
  NAND2_X1 U9592 ( .A1(n14420), .A2(n14419), .ZN(n7009) );
  INV_X1 U9593 ( .A(n14423), .ZN(n7014) );
  INV_X1 U9594 ( .A(n14128), .ZN(n7018) );
  INV_X1 U9595 ( .A(n14107), .ZN(n14110) );
  AND2_X1 U9596 ( .A1(n14107), .A2(n7019), .ZN(n14151) );
  INV_X1 U9597 ( .A(n14109), .ZN(n7019) );
  OAI21_X1 U9598 ( .B1(n15607), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6746), .ZN(
        n7023) );
  NAND2_X1 U9599 ( .A1(n10399), .A2(n10398), .ZN(n7817) );
  NAND2_X1 U9600 ( .A1(n10373), .A2(n12070), .ZN(n7024) );
  NAND2_X1 U9601 ( .A1(n7031), .A2(n7026), .ZN(n7028) );
  OAI211_X1 U9602 ( .C1(n13015), .C2(n7030), .A(n7029), .B(n7027), .ZN(n8294)
         );
  NAND3_X1 U9603 ( .A1(n13015), .A2(n7031), .A3(n8340), .ZN(n7029) );
  NAND2_X1 U9604 ( .A1(n7037), .A2(n6754), .ZN(n7039) );
  INV_X1 U9605 ( .A(n13075), .ZN(n7040) );
  OAI21_X1 U9606 ( .B1(n7040), .B2(n7043), .A(n6665), .ZN(n8199) );
  AND2_X1 U9607 ( .A1(n7066), .A2(n14198), .ZN(n12421) );
  NAND2_X1 U9608 ( .A1(n7071), .A2(n9985), .ZN(n10796) );
  INV_X1 U9609 ( .A(n10701), .ZN(n7073) );
  OAI21_X1 U9610 ( .B1(n7073), .B2(n7076), .A(n7074), .ZN(n8960) );
  INV_X1 U9611 ( .A(n11589), .ZN(n7082) );
  INV_X1 U9612 ( .A(n7083), .ZN(n11502) );
  NAND2_X1 U9613 ( .A1(n7092), .A2(n6751), .ZN(n7091) );
  NAND3_X1 U9614 ( .A1(n7101), .A2(n11575), .A3(n7100), .ZN(n10504) );
  NAND3_X1 U9615 ( .A1(n11723), .A2(n10585), .A3(n11719), .ZN(n7101) );
  OR2_X1 U9616 ( .A1(n12645), .A2(n7108), .ZN(n7103) );
  NAND2_X1 U9617 ( .A1(n7103), .A2(n7104), .ZN(n12591) );
  NAND3_X1 U9618 ( .A1(n7382), .A2(n7381), .A3(n7605), .ZN(n8466) );
  NAND2_X1 U9619 ( .A1(n11258), .A2(n7121), .ZN(n7118) );
  NAND2_X1 U9620 ( .A1(n7118), .A2(n7119), .ZN(n11422) );
  NAND2_X1 U9621 ( .A1(n13809), .A2(n7129), .ZN(n7127) );
  NAND2_X1 U9622 ( .A1(n7127), .A2(n7128), .ZN(n13769) );
  NAND2_X1 U9623 ( .A1(n13945), .A2(n7273), .ZN(n7134) );
  NAND2_X1 U9624 ( .A1(n9009), .A2(n7363), .ZN(n7136) );
  OR2_X1 U9625 ( .A1(n9610), .A2(n9485), .ZN(n7139) );
  NAND2_X2 U9626 ( .A1(n9043), .A2(n9042), .ZN(n9485) );
  OAI21_X1 U9627 ( .B1(n12137), .B2(n7142), .A(n12141), .ZN(n7141) );
  NAND2_X1 U9628 ( .A1(n12824), .A2(n12826), .ZN(n12825) );
  NAND2_X1 U9629 ( .A1(n12877), .A2(n7148), .ZN(n7147) );
  INV_X1 U9630 ( .A(n12113), .ZN(n7163) );
  NAND3_X1 U9631 ( .A1(n7162), .A2(n7164), .A3(n7159), .ZN(n12910) );
  NAND3_X1 U9632 ( .A1(n7162), .A2(n7160), .A3(n7159), .ZN(n7168) );
  INV_X1 U9633 ( .A(n7168), .ZN(n12907) );
  AND2_X2 U9634 ( .A1(n7168), .A2(n7167), .ZN(n12834) );
  NAND2_X1 U9635 ( .A1(n7170), .A2(n7169), .ZN(n10105) );
  NAND3_X1 U9636 ( .A1(n9900), .A2(n6700), .A3(n9901), .ZN(n7169) );
  NAND2_X1 U9637 ( .A1(n7171), .A2(n6700), .ZN(n7170) );
  NAND2_X1 U9638 ( .A1(n10098), .A2(n9925), .ZN(n7171) );
  INV_X2 U9639 ( .A(n10532), .ZN(n9889) );
  NAND2_X1 U9640 ( .A1(n13919), .A2(n6644), .ZN(n7174) );
  INV_X1 U9641 ( .A(n14532), .ZN(n7187) );
  NAND2_X1 U9642 ( .A1(n14532), .A2(n11261), .ZN(n7183) );
  NAND2_X1 U9643 ( .A1(n13803), .A2(n11790), .ZN(n7194) );
  NAND2_X1 U9644 ( .A1(n7824), .A2(n7839), .ZN(n9632) );
  MUX2_X1 U9645 ( .A(n10117), .B(P1_REG2_REG_3__SCAN_IN), .S(n13630), .Z(
        n13635) );
  NOR2_X2 U9646 ( .A1(n10273), .A2(n14891), .ZN(n10370) );
  OR2_X2 U9647 ( .A1(n10049), .A2(n11851), .ZN(n10273) );
  NOR2_X2 U9648 ( .A1(n11168), .A2(n14329), .ZN(n11252) );
  NAND3_X1 U9649 ( .A1(n13051), .A2(n11833), .A3(n7220), .ZN(n12995) );
  NAND2_X1 U9650 ( .A1(n13224), .A2(n13304), .ZN(n7226) );
  INV_X1 U9651 ( .A(n12997), .ZN(n7228) );
  OAI21_X1 U9652 ( .B1(n12333), .B2(n7244), .A(n7239), .ZN(n12272) );
  OAI21_X1 U9653 ( .B1(n12333), .B2(n12225), .A(n12224), .ZN(n12303) );
  NAND2_X1 U9654 ( .A1(n12226), .A2(n12227), .ZN(n7249) );
  OAI211_X1 U9655 ( .C1(n6804), .C2(n15116), .A(n10082), .B(n10033), .ZN(
        n10034) );
  NAND2_X1 U9656 ( .A1(n11150), .A2(n6648), .ZN(n7263) );
  INV_X1 U9657 ( .A(n12243), .ZN(n7265) );
  NOR2_X2 U9658 ( .A1(n7268), .A2(n9008), .ZN(n9009) );
  NAND4_X1 U9659 ( .A1(n7269), .A2(n9007), .A3(n9556), .A4(n8990), .ZN(n7268)
         );
  NAND2_X2 U9660 ( .A1(n13747), .A2(n13746), .ZN(n13958) );
  OAI21_X1 U9661 ( .B1(n13942), .B2(n7272), .A(n7270), .ZN(P1_U3525) );
  OR2_X1 U9662 ( .A1(n14675), .A2(n15292), .ZN(n7275) );
  AND2_X1 U9663 ( .A1(n9564), .A2(n7282), .ZN(n9026) );
  NAND2_X1 U9664 ( .A1(n9564), .A2(n6763), .ZN(n9014) );
  OAI211_X2 U9665 ( .C1(n9608), .C2(n9485), .A(n9065), .B(n7285), .ZN(n11088)
         );
  OR2_X1 U9666 ( .A1(n7768), .A2(n7767), .ZN(n7287) );
  NAND2_X1 U9667 ( .A1(n6753), .A2(n14173), .ZN(n13904) );
  XNOR2_X1 U9668 ( .A(n8437), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n8884) );
  NAND2_X2 U9669 ( .A1(n7297), .A2(n8426), .ZN(n8427) );
  NAND2_X1 U9670 ( .A1(n8821), .A2(n8820), .ZN(n7297) );
  NAND2_X1 U9671 ( .A1(n8808), .A2(n8424), .ZN(n7298) );
  NAND2_X1 U9672 ( .A1(n8399), .A2(n7305), .ZN(n7304) );
  NAND2_X1 U9673 ( .A1(n7310), .A2(n7309), .ZN(n8601) );
  NAND3_X1 U9674 ( .A1(n8571), .A2(n8584), .A3(n8570), .ZN(n7310) );
  NAND2_X1 U9675 ( .A1(n8613), .A2(n7320), .ZN(n7319) );
  NAND2_X1 U9676 ( .A1(n8752), .A2(n7327), .ZN(n7325) );
  NAND2_X1 U9677 ( .A1(n8693), .A2(n7332), .ZN(n7331) );
  OAI21_X2 U9678 ( .B1(n8846), .B2(n8845), .A(n8430), .ZN(n8855) );
  OR2_X2 U9679 ( .A1(n10607), .A2(n11890), .ZN(n10575) );
  NOR2_X4 U9680 ( .A1(n13191), .A2(n13289), .ZN(n13175) );
  NAND2_X1 U9681 ( .A1(n7350), .A2(n7349), .ZN(n13771) );
  NAND3_X1 U9682 ( .A1(n11091), .A2(n11090), .A3(n10868), .ZN(n7352) );
  INV_X1 U9683 ( .A(n10866), .ZN(n7354) );
  NAND2_X1 U9684 ( .A1(n10868), .A2(n10866), .ZN(n7351) );
  AND2_X1 U9685 ( .A1(n9009), .A2(n7362), .ZN(n7360) );
  NAND2_X1 U9686 ( .A1(n7135), .A2(n7360), .ZN(n7361) );
  NAND2_X1 U9687 ( .A1(n13751), .A2(n7369), .ZN(n7365) );
  AND2_X2 U9688 ( .A1(n8534), .A2(n8533), .ZN(n8536) );
  NAND2_X1 U9689 ( .A1(n11024), .A2(n7389), .ZN(n7386) );
  NAND2_X1 U9690 ( .A1(n7386), .A2(n7387), .ZN(n14273) );
  INV_X2 U9691 ( .A(n8594), .ZN(n11541) );
  NAND3_X1 U9692 ( .A1(n9396), .A2(n9395), .A3(n6769), .ZN(n7394) );
  INV_X1 U9693 ( .A(n9405), .ZN(n7395) );
  NAND2_X1 U9694 ( .A1(n9497), .A2(n11825), .ZN(n7397) );
  OAI21_X1 U9695 ( .B1(n13599), .B2(n9499), .A(n7396), .ZN(n9056) );
  NAND2_X4 U9696 ( .A1(n7398), .A2(n7397), .ZN(n9499) );
  NAND3_X1 U9697 ( .A1(n9453), .A2(n9452), .A3(n6767), .ZN(n7401) );
  INV_X1 U9698 ( .A(n9461), .ZN(n7402) );
  NAND3_X1 U9699 ( .A1(n9423), .A2(n9422), .A3(n6770), .ZN(n7404) );
  INV_X1 U9700 ( .A(n9434), .ZN(n7405) );
  NAND2_X1 U9701 ( .A1(n7406), .A2(n7407), .ZN(n9151) );
  NAND3_X1 U9702 ( .A1(n9129), .A2(n9128), .A3(n6760), .ZN(n7406) );
  NAND2_X1 U9703 ( .A1(n7408), .A2(n7409), .ZN(n9270) );
  NAND2_X1 U9704 ( .A1(n7413), .A2(n7414), .ZN(n9206) );
  NAND3_X1 U9705 ( .A1(n9173), .A2(n6762), .A3(n9172), .ZN(n7413) );
  NAND2_X1 U9706 ( .A1(n7418), .A2(n7416), .ZN(n9124) );
  INV_X1 U9707 ( .A(n9110), .ZN(n7417) );
  OAI211_X1 U9708 ( .C1(n9109), .C2(n7417), .A(n9093), .B(n9094), .ZN(n7418)
         );
  NAND4_X1 U9709 ( .A1(n8989), .A2(n7680), .A3(n7688), .A4(n8990), .ZN(n9281)
         );
  NOR2_X1 U9710 ( .A1(n8272), .A2(n7657), .ZN(n7423) );
  INV_X1 U9711 ( .A(n9917), .ZN(n7429) );
  AND2_X1 U9712 ( .A1(n9878), .A2(n14882), .ZN(n9917) );
  AOI21_X1 U9713 ( .B1(n7431), .B2(n7433), .A(n6664), .ZN(n7430) );
  INV_X1 U9714 ( .A(n7433), .ZN(n7432) );
  NAND2_X1 U9715 ( .A1(n7437), .A2(n8235), .ZN(n13004) );
  NAND2_X1 U9716 ( .A1(n10841), .A2(n7440), .ZN(n7917) );
  INV_X1 U9717 ( .A(n11902), .ZN(n7442) );
  NAND2_X1 U9718 ( .A1(n7455), .A2(n10804), .ZN(n7453) );
  XNOR2_X1 U9719 ( .A(n12412), .B(n12460), .ZN(n10804) );
  INV_X1 U9720 ( .A(n12414), .ZN(n7455) );
  INV_X1 U9721 ( .A(n15024), .ZN(n7456) );
  NAND3_X1 U9722 ( .A1(n7458), .A2(n7459), .A3(n7457), .ZN(n15073) );
  NAND3_X1 U9723 ( .A1(n7458), .A2(n6671), .A3(n7457), .ZN(n7460) );
  INV_X1 U9724 ( .A(n7460), .ZN(n15072) );
  NOR2_X1 U9725 ( .A1(n7471), .A2(n14975), .ZN(n7472) );
  OAI21_X1 U9726 ( .B1(n10799), .B2(n10800), .A(n7472), .ZN(n7473) );
  INV_X1 U9727 ( .A(n7473), .ZN(n14974) );
  INV_X1 U9728 ( .A(n10799), .ZN(n14964) );
  NAND2_X1 U9729 ( .A1(n7475), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n7618) );
  NAND3_X1 U9730 ( .A1(n12988), .A2(n7718), .A3(n7476), .ZN(n7475) );
  NAND2_X1 U9731 ( .A1(n7485), .A2(n10684), .ZN(n7483) );
  NAND2_X1 U9732 ( .A1(n10775), .A2(n10774), .ZN(n10776) );
  OAI21_X1 U9733 ( .B1(n10962), .B2(n7490), .A(n7487), .ZN(n11251) );
  NAND2_X2 U9734 ( .A1(n7502), .A2(n7500), .ZN(n12877) );
  NAND2_X1 U9735 ( .A1(n7508), .A2(n7506), .ZN(n13158) );
  INV_X1 U9736 ( .A(n12078), .ZN(n7510) );
  NOR2_X1 U9737 ( .A1(n12078), .A2(n7515), .ZN(n7514) );
  XNOR2_X1 U9738 ( .A(n10095), .B(n10094), .ZN(n10093) );
  XNOR2_X1 U9739 ( .A(n9889), .B(n14891), .ZN(n10094) );
  NAND2_X1 U9740 ( .A1(n7522), .A2(n7521), .ZN(n7520) );
  AOI21_X2 U9741 ( .B1(n13209), .B2(n13208), .A(n8320), .ZN(n13199) );
  OAI21_X2 U9742 ( .B1(n14310), .B2(n8318), .A(n8319), .ZN(n13209) );
  INV_X1 U9743 ( .A(n7654), .ZN(n7523) );
  NOR2_X2 U9744 ( .A1(n7654), .A2(n7524), .ZN(n7710) );
  OAI21_X1 U9745 ( .B1(n13046), .B2(n7529), .A(n7527), .ZN(n13021) );
  NAND2_X1 U9746 ( .A1(n7537), .A2(n7536), .ZN(n8306) );
  AND2_X1 U9747 ( .A1(n6694), .A2(n8304), .ZN(n7536) );
  NAND2_X1 U9748 ( .A1(n7539), .A2(n7538), .ZN(n8326) );
  AND2_X1 U9749 ( .A1(n12065), .A2(n7690), .ZN(n7538) );
  INV_X2 U9750 ( .A(n7736), .ZN(n7773) );
  NAND2_X1 U9751 ( .A1(n13517), .A2(n7551), .ZN(n7550) );
  AND2_X2 U9752 ( .A1(n7562), .A2(n10662), .ZN(n10754) );
  NAND2_X1 U9753 ( .A1(n13538), .A2(n7569), .ZN(n7563) );
  NOR2_X1 U9754 ( .A1(n13538), .A2(n7568), .ZN(n13489) );
  NAND2_X1 U9755 ( .A1(n13498), .A2(n7573), .ZN(n7572) );
  NAND2_X1 U9756 ( .A1(n13451), .A2(n13450), .ZN(n7584) );
  NAND2_X1 U9757 ( .A1(n10945), .A2(n8685), .ZN(n7592) );
  NAND2_X1 U9758 ( .A1(n11442), .A2(n11440), .ZN(n8778) );
  NAND2_X1 U9759 ( .A1(n12553), .A2(n6649), .ZN(n7600) );
  OAI21_X1 U9760 ( .B1(n7768), .B2(n7609), .A(n7607), .ZN(n7802) );
  NAND2_X1 U9761 ( .A1(n7880), .A2(n7612), .ZN(n7610) );
  NAND3_X1 U9762 ( .A1(n14139), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n7617) );
  NAND2_X1 U9763 ( .A1(n9504), .A2(n7626), .ZN(n7622) );
  NAND2_X1 U9764 ( .A1(n9504), .A2(n7620), .ZN(n7619) );
  NAND2_X1 U9765 ( .A1(n7932), .A2(n7636), .ZN(n7635) );
  OAI21_X1 U9766 ( .B1(n7932), .B2(n7638), .A(n7636), .ZN(n7971) );
  AOI21_X1 U9767 ( .B1(n7636), .B2(n7638), .A(n7634), .ZN(n7633) );
  NAND2_X1 U9768 ( .A1(n7643), .A2(n6668), .ZN(n8203) );
  NAND2_X1 U9769 ( .A1(n8052), .A2(n8051), .ZN(n7651) );
  OAI211_X2 U9770 ( .C1(n9642), .C2(n14714), .A(n7653), .B(n7652), .ZN(n11851)
         );
  NAND2_X2 U9771 ( .A1(n8286), .A2(n8288), .ZN(n7742) );
  INV_X1 U9772 ( .A(n11996), .ZN(n7660) );
  INV_X1 U9773 ( .A(n11871), .ZN(n7665) );
  NAND2_X1 U9774 ( .A1(n7666), .A2(n7667), .ZN(n11989) );
  NAND2_X1 U9775 ( .A1(n7668), .A2(n7670), .ZN(n11939) );
  NAND3_X1 U9776 ( .A1(n11881), .A2(n6756), .A3(n11880), .ZN(n7672) );
  NAND2_X1 U9777 ( .A1(n9394), .A2(n9393), .ZN(n9395) );
  NAND2_X1 U9778 ( .A1(n8157), .A2(n8156), .ZN(n8170) );
  NOR2_X2 U9779 ( .A1(n13080), .A2(n13066), .ZN(n13065) );
  NAND2_X1 U9780 ( .A1(n9421), .A2(n9420), .ZN(n9422) );
  INV_X1 U9781 ( .A(n12134), .ZN(n12136) );
  NAND2_X1 U9782 ( .A1(n13718), .A2(n11797), .ZN(n13703) );
  NAND2_X1 U9783 ( .A1(n13771), .A2(n11793), .ZN(n13751) );
  OAI21_X1 U9784 ( .B1(n9351), .B2(n9350), .A(n9349), .ZN(n9353) );
  AND4_X2 U9785 ( .A1(n9051), .A2(n9050), .A3(n9049), .A4(n9048), .ZN(n10144)
         );
  AND2_X1 U9786 ( .A1(n9530), .A2(n9529), .ZN(n9531) );
  NAND2_X1 U9787 ( .A1(n9273), .A2(n9272), .ZN(n9322) );
  NAND2_X1 U9788 ( .A1(n13703), .A2(n11798), .ZN(n11799) );
  INV_X1 U9789 ( .A(n14037), .ZN(n9016) );
  NAND2_X1 U9790 ( .A1(n8979), .A2(n14924), .ZN(n8984) );
  INV_X1 U9791 ( .A(n9095), .ZN(n8989) );
  NAND2_X1 U9792 ( .A1(n10304), .A2(n10303), .ZN(n10306) );
  CLKBUF_X1 U9793 ( .A(n10547), .Z(n10470) );
  NOR2_X1 U9794 ( .A1(n9486), .A2(n11828), .ZN(n9487) );
  CLKBUF_X1 U9795 ( .A(n9294), .Z(n9295) );
  INV_X1 U9796 ( .A(n10353), .ZN(n10347) );
  AND2_X1 U9797 ( .A1(n10012), .A2(n10009), .ZN(n14632) );
  XNOR2_X1 U9798 ( .A(n12944), .B(n11854), .ZN(n12067) );
  XNOR2_X1 U9799 ( .A(n11802), .B(n11801), .ZN(n13936) );
  NAND2_X1 U9800 ( .A1(n11799), .A2(n7683), .ZN(n11802) );
  NOR2_X2 U9801 ( .A1(n10357), .A2(n10313), .ZN(n11086) );
  CLKBUF_X1 U9802 ( .A(n9908), .Z(n12409) );
  INV_X1 U9803 ( .A(n10586), .ZN(n9908) );
  AND2_X2 U9804 ( .A1(n13531), .A2(n13530), .ZN(n13538) );
  OAI21_X1 U9805 ( .B1(n11982), .B2(n12031), .A(n11981), .ZN(n11983) );
  OAI21_X1 U9806 ( .B1(n11973), .B2(n12031), .A(n11972), .ZN(n11974) );
  XNOR2_X2 U9807 ( .A(n8341), .B(n8340), .ZN(n11839) );
  XNOR2_X1 U9808 ( .A(n7720), .B(n7721), .ZN(n8288) );
  INV_X1 U9809 ( .A(n10897), .ZN(n10902) );
  AND2_X2 U9810 ( .A1(n9016), .A2(n9017), .ZN(n9082) );
  INV_X1 U9811 ( .A(n8343), .ZN(n12098) );
  NAND2_X1 U9812 ( .A1(n8312), .A2(n8311), .ZN(n10962) );
  OR2_X1 U9813 ( .A1(n11251), .A2(n8315), .ZN(n8317) );
  NOR2_X2 U9814 ( .A1(n13874), .A2(n13852), .ZN(n13851) );
  AND2_X1 U9815 ( .A1(n8728), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7678) );
  INV_X1 U9816 ( .A(n12633), .ZN(n8819) );
  NAND2_X1 U9817 ( .A1(n10285), .A2(n14270), .ZN(n12657) );
  INV_X2 U9818 ( .A(n12657), .ZN(n15595) );
  INV_X1 U9819 ( .A(n15202), .ZN(n8976) );
  OR2_X1 U9820 ( .A1(n15183), .A2(n15146), .ZN(n12771) );
  INV_X1 U9821 ( .A(n12771), .ZN(n9586) );
  AND3_X1 U9822 ( .A1(n9196), .A2(n8988), .A3(n9242), .ZN(n7680) );
  AND2_X1 U9823 ( .A1(n10900), .A2(n10899), .ZN(n7681) );
  AND2_X1 U9824 ( .A1(n14541), .A2(n11207), .ZN(n7682) );
  OR2_X1 U9825 ( .A1(n13709), .A2(n13579), .ZN(n7683) );
  AND2_X1 U9826 ( .A1(n12033), .A2(n12032), .ZN(n7686) );
  OR3_X1 U9827 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .A3(
        n15429), .ZN(n7687) );
  INV_X1 U9828 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8361) );
  OR2_X1 U9829 ( .A1(n13273), .A2(n12925), .ZN(n7690) );
  AND2_X1 U9830 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n7691) );
  AND2_X1 U9831 ( .A1(n10862), .A2(n9068), .ZN(n7692) );
  INV_X4 U9832 ( .A(n9042), .ZN(n8205) );
  NAND2_X1 U9833 ( .A1(n12022), .A2(n13304), .ZN(n7693) );
  INV_X1 U9834 ( .A(n12022), .ZN(n11833) );
  INV_X1 U9835 ( .A(n8670), .ZN(n8829) );
  AND2_X1 U9836 ( .A1(n10976), .A2(n13599), .ZN(n9068) );
  NAND2_X1 U9837 ( .A1(n9069), .A2(n7692), .ZN(n9070) );
  AOI22_X1 U9838 ( .A1(n12943), .A2(n12051), .B1(n11851), .B2(n12031), .ZN(
        n11859) );
  INV_X1 U9839 ( .A(n9141), .ZN(n9142) );
  NAND2_X1 U9840 ( .A1(n9209), .A2(n9208), .ZN(n9210) );
  NAND2_X1 U9841 ( .A1(n11926), .A2(n11925), .ZN(n11931) );
  OAI21_X1 U9842 ( .B1(n11943), .B2(n12031), .A(n11942), .ZN(n11944) );
  INV_X1 U9843 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8454) );
  INV_X1 U9844 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n7698) );
  INV_X1 U9845 ( .A(n9473), .ZN(n9510) );
  NAND2_X1 U9846 ( .A1(n9967), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n9858) );
  INV_X1 U9847 ( .A(n12469), .ZN(n12470) );
  INV_X1 U9848 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n8472) );
  AND2_X1 U9849 ( .A1(n7719), .A2(n7721), .ZN(n7708) );
  INV_X1 U9850 ( .A(n10472), .ZN(n10468) );
  INV_X1 U9851 ( .A(n14357), .ZN(n11260) );
  INV_X1 U9852 ( .A(n8813), .ZN(n8522) );
  OAI21_X1 U9853 ( .B1(n9967), .B2(P3_REG1_REG_2__SCAN_IN), .A(n9850), .ZN(
        n9856) );
  INV_X1 U9854 ( .A(n15074), .ZN(n12468) );
  NAND2_X1 U9855 ( .A1(n8527), .A2(n8526), .ZN(n8910) );
  INV_X1 U9856 ( .A(n11675), .ZN(n12567) );
  NAND2_X1 U9857 ( .A1(n12407), .A2(n11578), .ZN(n11572) );
  NAND2_X1 U9858 ( .A1(n12127), .A2(n12129), .ZN(n12130) );
  INV_X1 U9859 ( .A(n7911), .ZN(n7909) );
  INV_X1 U9860 ( .A(n8130), .ZN(n8129) );
  INV_X1 U9861 ( .A(n13074), .ZN(n8167) );
  INV_X1 U9862 ( .A(n9606), .ZN(n9044) );
  INV_X1 U9863 ( .A(n9486), .ZN(n9136) );
  INV_X1 U9864 ( .A(SI_16_), .ZN(n8032) );
  NAND2_X1 U9865 ( .A1(n8522), .A2(n8521), .ZN(n8826) );
  INV_X1 U9866 ( .A(n8849), .ZN(n8524) );
  INV_X1 U9867 ( .A(n8838), .ZN(n8523) );
  INV_X1 U9868 ( .A(n8828), .ZN(n8949) );
  OR2_X1 U9869 ( .A1(n8861), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8873) );
  INV_X1 U9870 ( .A(n15093), .ZN(n12471) );
  AND2_X1 U9871 ( .A1(n10281), .A2(n10280), .ZN(n10282) );
  NOR2_X1 U9872 ( .A1(n8953), .A2(n8952), .ZN(n8954) );
  INV_X1 U9873 ( .A(n15119), .ZN(n12374) );
  INV_X1 U9874 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n8418) );
  AND2_X1 U9875 ( .A1(n8393), .A2(n8392), .ZN(n8612) );
  INV_X1 U9876 ( .A(n11188), .ZN(n11185) );
  INV_X1 U9877 ( .A(n7963), .ZN(n7962) );
  AND2_X1 U9878 ( .A1(n12098), .A2(n12105), .ZN(n9816) );
  OR2_X1 U9879 ( .A1(n8212), .A2(n12893), .ZN(n8227) );
  OR2_X1 U9880 ( .A1(n8143), .A2(n8142), .ZN(n8161) );
  NAND2_X1 U9881 ( .A1(n8082), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8110) );
  OR2_X1 U9882 ( .A1(n14762), .A2(n14761), .ZN(n14782) );
  AND2_X1 U9883 ( .A1(n8227), .A2(n8213), .ZN(n13034) );
  INV_X1 U9884 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n8379) );
  NOR2_X1 U9885 ( .A1(n9341), .A2(n9340), .ZN(n9354) );
  INV_X1 U9886 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9101) );
  NAND2_X1 U9887 ( .A1(n9519), .A2(n9518), .ZN(n9532) );
  INV_X1 U9888 ( .A(n13935), .ZN(n13690) );
  INV_X1 U9889 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n9229) );
  INV_X1 U9890 ( .A(n14537), .ZN(n13854) );
  INV_X1 U9891 ( .A(n10007), .ZN(n10023) );
  OR2_X1 U9892 ( .A1(n9219), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n9220) );
  INV_X1 U9893 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9112) );
  OR2_X1 U9894 ( .A1(n8686), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8703) );
  OR2_X1 U9895 ( .A1(n8826), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8838) );
  INV_X1 U9896 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n15315) );
  INV_X1 U9897 ( .A(n12305), .ZN(n12569) );
  NAND2_X1 U9898 ( .A1(n8668), .A2(n11152), .ZN(n8686) );
  INV_X1 U9899 ( .A(n12387), .ZN(n12228) );
  AND2_X1 U9900 ( .A1(n11546), .A2(n8940), .ZN(n12503) );
  INV_X1 U9901 ( .A(n15033), .ZN(n12462) );
  INV_X1 U9902 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n15040) );
  INV_X1 U9903 ( .A(n15016), .ZN(n15101) );
  AND2_X1 U9904 ( .A1(n9827), .A2(n9828), .ZN(n9835) );
  AND2_X1 U9905 ( .A1(n11669), .A2(n11670), .ZN(n12593) );
  INV_X1 U9906 ( .A(n8963), .ZN(n11737) );
  INV_X1 U9907 ( .A(n12375), .ZN(n15117) );
  INV_X1 U9908 ( .A(n14288), .ZN(n15594) );
  AND2_X1 U9909 ( .A1(n8652), .A2(n12286), .ZN(n8668) );
  INV_X1 U9910 ( .A(n9825), .ZN(n8822) );
  NOR2_X1 U9911 ( .A1(n9947), .A2(n11755), .ZN(n9954) );
  INV_X1 U9912 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n15330) );
  AND2_X1 U9913 ( .A1(n8401), .A2(n8400), .ZN(n8662) );
  AND2_X1 U9914 ( .A1(n8390), .A2(n8389), .ZN(n8600) );
  INV_X1 U9915 ( .A(n12789), .ZN(n12151) );
  NAND2_X1 U9916 ( .A1(n12136), .A2(n12135), .ZN(n12137) );
  OR2_X1 U9917 ( .A1(n7893), .A2(n7892), .ZN(n7911) );
  NAND2_X1 U9918 ( .A1(n7962), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7978) );
  NOR2_X1 U9919 ( .A1(n8227), .A2(n12794), .ZN(n8259) );
  OR2_X1 U9920 ( .A1(n13053), .A2(n8229), .ZN(n8197) );
  INV_X1 U9921 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n14818) );
  OR2_X1 U9922 ( .A1(n7995), .A2(n7994), .ZN(n8022) );
  INV_X1 U9923 ( .A(n12901), .ZN(n12889) );
  INV_X1 U9924 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8980) );
  INV_X1 U9925 ( .A(n12070), .ZN(n10372) );
  INV_X1 U9926 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7721) );
  NOR2_X1 U9927 ( .A1(n9174), .A2(n15558), .ZN(n9190) );
  NOR2_X1 U9928 ( .A1(n9275), .A2(n9274), .ZN(n9300) );
  INV_X1 U9929 ( .A(n9409), .ZN(n9408) );
  OR2_X1 U9930 ( .A1(n9553), .A2(n9552), .ZN(n9554) );
  AND2_X1 U9931 ( .A1(n9465), .A2(n9439), .ZN(n13723) );
  INV_X1 U9932 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14049) );
  INV_X1 U9933 ( .A(n13770), .ZN(n13772) );
  NOR2_X1 U9934 ( .A1(n15432), .A2(n9382), .ZN(n9397) );
  OR2_X1 U9935 ( .A1(n9260), .A2(n9259), .ZN(n9275) );
  NAND2_X1 U9936 ( .A1(n10298), .A2(n10878), .ZN(n10309) );
  OR2_X1 U9937 ( .A1(n10873), .A2(n10872), .ZN(n13857) );
  INV_X1 U9938 ( .A(n14554), .ZN(n14666) );
  INV_X1 U9939 ( .A(n12278), .ZN(n12289) );
  NAND2_X1 U9940 ( .A1(n9960), .A2(n14270), .ZN(n12380) );
  NAND2_X1 U9941 ( .A1(n8894), .A2(n8893), .ZN(n12305) );
  AND4_X1 U9942 ( .A1(n8793), .A2(n8792), .A3(n8791), .A4(n8790), .ZN(n12326)
         );
  INV_X1 U9943 ( .A(n15082), .ZN(n15104) );
  AND2_X1 U9944 ( .A1(n9835), .A2(n9834), .ZN(n14998) );
  OR2_X1 U9945 ( .A1(n10285), .A2(n11750), .ZN(n10392) );
  AND2_X1 U9946 ( .A1(n12629), .A2(n12628), .ZN(n12711) );
  INV_X1 U9947 ( .A(n14264), .ZN(n15122) );
  INV_X1 U9948 ( .A(n10392), .ZN(n14276) );
  INV_X1 U9949 ( .A(n11750), .ZN(n15126) );
  INV_X1 U9950 ( .A(n8514), .ZN(n8515) );
  NAND2_X1 U9951 ( .A1(n8975), .A2(n11559), .ZN(n15146) );
  AND2_X1 U9952 ( .A1(n8975), .A2(n11750), .ZN(n15179) );
  OR2_X1 U9953 ( .A1(n9957), .A2(n9580), .ZN(n9583) );
  AND2_X1 U9954 ( .A1(n8498), .A2(n8497), .ZN(n10279) );
  INV_X1 U9955 ( .A(n12908), .ZN(n12887) );
  AND3_X1 U9956 ( .A1(n8285), .A2(n8284), .A3(n8283), .ZN(n12018) );
  INV_X1 U9957 ( .A(n7997), .ZN(n8229) );
  INV_X1 U9958 ( .A(n12008), .ZN(n8262) );
  AND2_X1 U9959 ( .A1(n9658), .A2(n9657), .ZN(n14811) );
  INV_X1 U9960 ( .A(n12095), .ZN(n13003) );
  INV_X1 U9961 ( .A(n12089), .ZN(n13120) );
  INV_X1 U9962 ( .A(n12082), .ZN(n11102) );
  INV_X1 U9963 ( .A(n13211), .ZN(n14837) );
  INV_X1 U9964 ( .A(n13194), .ZN(n14841) );
  INV_X1 U9965 ( .A(n13329), .ZN(n8982) );
  INV_X1 U9966 ( .A(n14905), .ZN(n14895) );
  NAND2_X1 U9967 ( .A1(n9870), .A2(n9916), .ZN(n14905) );
  INV_X1 U9968 ( .A(n10190), .ZN(n9808) );
  AND2_X1 U9969 ( .A1(n8373), .A2(n8364), .ZN(n14849) );
  INV_X1 U9970 ( .A(n13546), .ZN(n14359) );
  INV_X1 U9971 ( .A(n13564), .ZN(n14350) );
  INV_X1 U9972 ( .A(n11305), .ZN(n9559) );
  AND3_X1 U9973 ( .A1(n9346), .A2(n9345), .A3(n9344), .ZN(n13827) );
  AND4_X1 U9974 ( .A1(n9265), .A2(n9264), .A3(n9263), .A4(n9262), .ZN(n13899)
         );
  INV_X1 U9975 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14047) );
  INV_X1 U9976 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n14066) );
  INV_X1 U9977 ( .A(n14483), .ZN(n14517) );
  INV_X1 U9978 ( .A(n14525), .ZN(n14494) );
  INV_X1 U9979 ( .A(n13903), .ZN(n14561) );
  NAND2_X1 U9980 ( .A1(n14163), .A2(n11411), .ZN(n11412) );
  NAND2_X1 U9981 ( .A1(n13857), .A2(n11808), .ZN(n13902) );
  AOI21_X1 U9982 ( .B1(n10006), .B2(n10005), .A(n10004), .ZN(n10318) );
  OR2_X1 U9983 ( .A1(n10298), .A2(n10297), .ZN(n14636) );
  INV_X1 U9984 ( .A(n14551), .ZN(n14639) );
  INV_X1 U9985 ( .A(n14018), .ZN(n14671) );
  NAND2_X1 U9986 ( .A1(n9745), .A2(n14038), .ZN(n10003) );
  AND2_X1 U9987 ( .A1(n9829), .A2(n9828), .ZN(n15025) );
  INV_X1 U9988 ( .A(n12380), .ZN(n12352) );
  INV_X1 U9989 ( .A(n12502), .ZN(n12386) );
  AND4_X1 U9990 ( .A1(n8746), .A2(n8745), .A3(n8744), .A4(n8743), .ZN(n11483)
         );
  INV_X1 U9991 ( .A(n14998), .ZN(n15110) );
  INV_X1 U9992 ( .A(n15600), .ZN(n12659) );
  NAND2_X1 U9993 ( .A1(n12657), .A2(n10383), .ZN(n12576) );
  AOI21_X1 U9994 ( .B1(n8941), .B2(n8517), .A(n8516), .ZN(n8977) );
  NAND2_X1 U9995 ( .A1(n15202), .A2(n15157), .ZN(n12721) );
  AND2_X2 U9996 ( .A1(n10283), .A2(n8515), .ZN(n15202) );
  INV_X1 U9997 ( .A(n12361), .ZN(n12747) );
  INV_X2 U9998 ( .A(n15183), .ZN(n15181) );
  AND2_X1 U9999 ( .A1(n9583), .A2(n9582), .ZN(n15183) );
  INV_X1 U10000 ( .A(SI_20_), .ZN(n10325) );
  INV_X1 U10001 ( .A(SI_12_), .ZN(n15490) );
  INV_X1 U10002 ( .A(n14982), .ZN(n10812) );
  INV_X1 U10003 ( .A(n11876), .ZN(n14901) );
  INV_X1 U10004 ( .A(n11934), .ZN(n14325) );
  AND2_X1 U10005 ( .A1(n9814), .A2(n13194), .ZN(n12900) );
  INV_X1 U10006 ( .A(n12892), .ZN(n12918) );
  OR2_X1 U10007 ( .A1(n8027), .A2(n8026), .ZN(n12929) );
  INV_X1 U10008 ( .A(n11909), .ZN(n12935) );
  OR2_X1 U10009 ( .A1(n14696), .A2(P2_U3088), .ZN(n14833) );
  OR2_X1 U10010 ( .A1(n9658), .A2(P2_U3088), .ZN(n14817) );
  OR2_X1 U10011 ( .A1(n13211), .A2(n10264), .ZN(n13182) );
  AND2_X1 U10012 ( .A1(n10201), .A2(n13194), .ZN(n13211) );
  INV_X1 U10013 ( .A(n14934), .ZN(n14932) );
  INV_X1 U10014 ( .A(n12989), .ZN(n13308) );
  INV_X1 U10015 ( .A(n13270), .ZN(n13330) );
  AND2_X1 U10016 ( .A1(n14335), .A2(n14334), .ZN(n14341) );
  INV_X1 U10017 ( .A(n14924), .ZN(n14922) );
  INV_X1 U10018 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n13354) );
  XNOR2_X1 U10019 ( .A(n8362), .B(n8361), .ZN(n11335) );
  INV_X1 U10020 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10524) );
  INV_X1 U10021 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9792) );
  AND2_X1 U10022 ( .A1(n10454), .A2(n11305), .ZN(n14365) );
  INV_X1 U10023 ( .A(n14169), .ZN(n14391) );
  NAND4_X1 U10024 ( .A1(n9431), .A2(n9430), .A3(n9429), .A4(n9428), .ZN(n13580) );
  INV_X1 U10025 ( .A(n13827), .ZN(n13855) );
  NAND2_X1 U10026 ( .A1(n9799), .A2(n9797), .ZN(n14529) );
  INV_X1 U10027 ( .A(n14567), .ZN(n13927) );
  AND2_X1 U10028 ( .A1(n14167), .A2(n14166), .ZN(n14390) );
  INV_X1 U10029 ( .A(n13902), .ZN(n13930) );
  AND2_X2 U10030 ( .A1(n10319), .A2(n10318), .ZN(n14688) );
  INV_X1 U10031 ( .A(n14675), .ZN(n14673) );
  AND2_X2 U10032 ( .A1(n10319), .A2(n10874), .ZN(n14675) );
  AND2_X2 U10033 ( .A1(n10871), .A2(n10003), .ZN(n14606) );
  NAND2_X1 U10034 ( .A1(n9558), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11305) );
  INV_X1 U10035 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10043) );
  INV_X2 U10036 ( .A(n12410), .ZN(P3_U3897) );
  NOR2_X1 U10037 ( .A1(n9643), .A2(n9587), .ZN(P2_U3947) );
  NAND2_X1 U10038 ( .A1(n8984), .A2(n8983), .ZN(P2_U3496) );
  AND2_X2 U10039 ( .A1(n9793), .A2(n9588), .ZN(P1_U4016) );
  NOR2_X1 U10040 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), 
        .ZN(n7696) );
  NAND4_X1 U10041 ( .A1(n7696), .A2(n7695), .A3(n7694), .A4(n7933), .ZN(n8036)
         );
  NAND3_X1 U10042 ( .A1(n7886), .A2(n7698), .A3(n7697), .ZN(n7699) );
  NOR2_X2 U10043 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n7727) );
  AND2_X2 U10044 ( .A1(n7727), .A2(n7700), .ZN(n7745) );
  NAND2_X1 U10045 ( .A1(n7997), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7717) );
  NAND2_X1 U10046 ( .A1(n7832), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7716) );
  INV_X1 U10047 ( .A(n7712), .ZN(n13346) );
  INV_X1 U10048 ( .A(n11843), .ZN(n9878) );
  NAND2_X1 U10049 ( .A1(n8205), .A2(SI_0_), .ZN(n8562) );
  XNOR2_X1 U10050 ( .A(n8562), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n13361) );
  NAND2_X1 U10051 ( .A1(n7997), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n7725) );
  NAND2_X1 U10052 ( .A1(n7737), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n7724) );
  NAND2_X1 U10053 ( .A1(n7832), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7722) );
  NAND4_X4 U10054 ( .A1(n7725), .A2(n7724), .A3(n7723), .A4(n7722), .ZN(n12944) );
  NAND2_X1 U10055 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n7726) );
  MUX2_X1 U10056 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7726), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n7729) );
  INV_X1 U10057 ( .A(n7727), .ZN(n7728) );
  NAND2_X1 U10058 ( .A1(n7729), .A2(n7728), .ZN(n9659) );
  NAND2_X1 U10059 ( .A1(n7730), .A2(SI_1_), .ZN(n7749) );
  NAND2_X1 U10060 ( .A1(n7731), .A2(SI_0_), .ZN(n7750) );
  XNOR2_X1 U10061 ( .A(n7751), .B(n7750), .ZN(n9606) );
  OR2_X1 U10062 ( .A1(n7763), .A2(n9606), .ZN(n7733) );
  OR2_X1 U10063 ( .A1(n7769), .A2(n6989), .ZN(n7732) );
  OAI211_X1 U10064 ( .C1(n7742), .C2(n9659), .A(n7733), .B(n7732), .ZN(n11854)
         );
  NAND2_X1 U10065 ( .A1(n9917), .A2(n12067), .ZN(n7735) );
  INV_X1 U10066 ( .A(n12944), .ZN(n9815) );
  NAND2_X1 U10067 ( .A1(n9815), .A2(n9920), .ZN(n7734) );
  NAND2_X1 U10068 ( .A1(n7735), .A2(n7734), .ZN(n10045) );
  NAND2_X1 U10069 ( .A1(n7997), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n7741) );
  NAND2_X1 U10070 ( .A1(n7832), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7740) );
  NAND2_X1 U10071 ( .A1(n7736), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7739) );
  NAND2_X1 U10072 ( .A1(n7737), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n7738) );
  NOR2_X1 U10073 ( .A1(n7727), .A2(n8268), .ZN(n7743) );
  MUX2_X1 U10074 ( .A(n8268), .B(n7743), .S(P2_IR_REG_2__SCAN_IN), .Z(n7744)
         );
  INV_X1 U10075 ( .A(n7744), .ZN(n7748) );
  INV_X1 U10076 ( .A(n7746), .ZN(n7747) );
  NAND2_X1 U10077 ( .A1(n7748), .A2(n7747), .ZN(n14714) );
  NAND2_X1 U10078 ( .A1(n7752), .A2(SI_2_), .ZN(n7764) );
  INV_X1 U10079 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9600) );
  XNOR2_X1 U10080 ( .A(n12943), .B(n11851), .ZN(n12069) );
  NAND2_X1 U10081 ( .A1(n10045), .A2(n12069), .ZN(n7754) );
  INV_X1 U10082 ( .A(n12943), .ZN(n9877) );
  NAND2_X1 U10083 ( .A1(n9877), .A2(n11851), .ZN(n7753) );
  NAND2_X1 U10084 ( .A1(n7754), .A2(n7753), .ZN(n10266) );
  INV_X1 U10085 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10270) );
  NAND2_X1 U10086 ( .A1(n7997), .A2(n10270), .ZN(n7758) );
  NAND2_X1 U10087 ( .A1(n7832), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7757) );
  INV_X2 U10088 ( .A(n7773), .ZN(n12007) );
  NAND2_X1 U10089 ( .A1(n12007), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7756) );
  NOR2_X1 U10090 ( .A1(n7746), .A2(n8268), .ZN(n7759) );
  MUX2_X1 U10091 ( .A(n8268), .B(n7759), .S(P2_IR_REG_3__SCAN_IN), .Z(n7760)
         );
  INV_X1 U10092 ( .A(n7760), .ZN(n7762) );
  NAND2_X1 U10093 ( .A1(n7746), .A2(n7761), .ZN(n7781) );
  NAND2_X1 U10094 ( .A1(n7762), .A2(n7781), .ZN(n9686) );
  OR2_X1 U10095 ( .A1(n7769), .A2(n9596), .ZN(n7770) );
  XNOR2_X1 U10096 ( .A(n12942), .B(n14891), .ZN(n12068) );
  NAND2_X1 U10097 ( .A1(n10266), .A2(n12068), .ZN(n7772) );
  INV_X1 U10098 ( .A(n12942), .ZN(n8300) );
  NAND2_X1 U10099 ( .A1(n8300), .A2(n14891), .ZN(n7771) );
  NAND2_X1 U10100 ( .A1(n8065), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n7779) );
  NAND2_X1 U10101 ( .A1(n8281), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7778) );
  INV_X1 U10102 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n7774) );
  NAND2_X1 U10103 ( .A1(n10270), .A2(n7774), .ZN(n7775) );
  NAND2_X1 U10104 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7795) );
  AND2_X1 U10105 ( .A1(n7775), .A2(n7795), .ZN(n10488) );
  NAND2_X1 U10106 ( .A1(n7997), .A2(n10488), .ZN(n7777) );
  NAND2_X1 U10107 ( .A1(n12008), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7776) );
  NAND4_X1 U10108 ( .A1(n7779), .A2(n7778), .A3(n7777), .A4(n7776), .ZN(n12941) );
  NAND2_X1 U10109 ( .A1(n7781), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7780) );
  MUX2_X1 U10110 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7780), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n7782) );
  NAND2_X1 U10111 ( .A1(n7782), .A2(n7809), .ZN(n9687) );
  OAI22_X1 U10112 ( .A1(n12013), .A2(n9599), .B1(n9642), .B2(n9687), .ZN(n7790) );
  OAI21_X1 U10113 ( .B1(n7785), .B2(SI_4_), .A(n7801), .ZN(n7786) );
  NOR2_X1 U10114 ( .A1(n9603), .A2(n8209), .ZN(n7789) );
  XNOR2_X1 U10115 ( .A(n12941), .B(n11870), .ZN(n12070) );
  INV_X1 U10116 ( .A(n12941), .ZN(n8303) );
  NAND2_X1 U10117 ( .A1(n8303), .A2(n11870), .ZN(n7791) );
  NAND2_X1 U10118 ( .A1(n8282), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n7800) );
  NAND2_X1 U10119 ( .A1(n12007), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7799) );
  INV_X1 U10120 ( .A(n7795), .ZN(n7793) );
  NAND2_X1 U10121 ( .A1(n7793), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7830) );
  INV_X1 U10122 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7794) );
  NAND2_X1 U10123 ( .A1(n7795), .A2(n7794), .ZN(n7796) );
  AND2_X1 U10124 ( .A1(n7830), .A2(n7796), .ZN(n10405) );
  NAND2_X1 U10125 ( .A1(n7997), .A2(n10405), .ZN(n7798) );
  NAND2_X1 U10126 ( .A1(n12008), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7797) );
  NAND4_X1 U10127 ( .A1(n7800), .A2(n7799), .A3(n7798), .A4(n7797), .ZN(n12940) );
  INV_X1 U10128 ( .A(n12940), .ZN(n7815) );
  NAND2_X1 U10129 ( .A1(n7803), .A2(SI_5_), .ZN(n7818) );
  OAI21_X1 U10130 ( .B1(n7803), .B2(SI_5_), .A(n7818), .ZN(n7804) );
  INV_X1 U10131 ( .A(n7804), .ZN(n7805) );
  OR2_X1 U10132 ( .A1(n7806), .A2(n7805), .ZN(n7807) );
  NAND2_X1 U10133 ( .A1(n7819), .A2(n7807), .ZN(n9615) );
  OR2_X1 U10134 ( .A1(n9615), .A2(n8209), .ZN(n7814) );
  NAND2_X1 U10135 ( .A1(n7809), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7808) );
  MUX2_X1 U10136 ( .A(n7808), .B(P2_IR_REG_31__SCAN_IN), .S(n7810), .Z(n7812)
         );
  INV_X1 U10137 ( .A(n7809), .ZN(n7811) );
  NAND2_X1 U10138 ( .A1(n7811), .A2(n7810), .ZN(n7845) );
  NAND2_X1 U10139 ( .A1(n7812), .A2(n7845), .ZN(n9695) );
  INV_X1 U10140 ( .A(n9695), .ZN(n9766) );
  AOI22_X1 U10141 ( .A1(n8079), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n8078), .B2(
        n9766), .ZN(n7813) );
  NAND2_X1 U10142 ( .A1(n7814), .A2(n7813), .ZN(n11876) );
  XNOR2_X1 U10143 ( .A(n7815), .B(n11876), .ZN(n12073) );
  NAND2_X1 U10144 ( .A1(n7815), .A2(n11876), .ZN(n7816) );
  NAND2_X1 U10145 ( .A1(n7817), .A2(n7816), .ZN(n10601) );
  MUX2_X1 U10146 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n9371), .Z(n7820) );
  NAND2_X1 U10147 ( .A1(n7820), .A2(SI_6_), .ZN(n7838) );
  OAI21_X1 U10148 ( .B1(n7820), .B2(SI_6_), .A(n7838), .ZN(n7821) );
  INV_X1 U10149 ( .A(n7821), .ZN(n7822) );
  OR2_X1 U10150 ( .A1(n7823), .A2(n7822), .ZN(n7824) );
  OR2_X1 U10151 ( .A1(n9632), .A2(n8209), .ZN(n7827) );
  NAND2_X1 U10152 ( .A1(n7845), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7825) );
  XNOR2_X1 U10153 ( .A(n7825), .B(P2_IR_REG_6__SCAN_IN), .ZN(n9769) );
  AOI22_X1 U10154 ( .A1(n8079), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8078), .B2(
        n9769), .ZN(n7826) );
  NAND2_X1 U10155 ( .A1(n7827), .A2(n7826), .ZN(n11884) );
  NAND2_X1 U10156 ( .A1(n8065), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n7836) );
  NAND2_X1 U10157 ( .A1(n8281), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7835) );
  INV_X1 U10158 ( .A(n7830), .ZN(n7828) );
  NAND2_X1 U10159 ( .A1(n7828), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7851) );
  INV_X1 U10160 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7829) );
  NAND2_X1 U10161 ( .A1(n7830), .A2(n7829), .ZN(n7831) );
  AND2_X1 U10162 ( .A1(n7851), .A2(n7831), .ZN(n10478) );
  NAND2_X1 U10163 ( .A1(n7997), .A2(n10478), .ZN(n7834) );
  NAND2_X1 U10164 ( .A1(n12008), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7833) );
  NAND4_X1 U10165 ( .A1(n7836), .A2(n7835), .A3(n7834), .A4(n7833), .ZN(n12939) );
  XNOR2_X1 U10166 ( .A(n11884), .B(n12939), .ZN(n12075) );
  INV_X1 U10167 ( .A(n12939), .ZN(n11886) );
  NAND2_X1 U10168 ( .A1(n11884), .A2(n11886), .ZN(n7837) );
  MUX2_X1 U10169 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n9371), .Z(n7840) );
  NAND2_X1 U10170 ( .A1(n7840), .A2(SI_7_), .ZN(n7859) );
  OAI21_X1 U10171 ( .B1(n7840), .B2(SI_7_), .A(n7859), .ZN(n7841) );
  INV_X1 U10172 ( .A(n7841), .ZN(n7842) );
  OR2_X1 U10173 ( .A1(n7843), .A2(n7842), .ZN(n7844) );
  NAND2_X1 U10174 ( .A1(n7860), .A2(n7844), .ZN(n9637) );
  OR2_X1 U10175 ( .A1(n9637), .A2(n8209), .ZN(n7848) );
  OAI21_X1 U10176 ( .B1(n7845), .B2(P2_IR_REG_6__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7846) );
  XNOR2_X1 U10177 ( .A(n7846), .B(P2_IR_REG_7__SCAN_IN), .ZN(n12951) );
  AOI22_X1 U10178 ( .A1(n8079), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8078), .B2(
        n12951), .ZN(n7847) );
  NAND2_X1 U10179 ( .A1(n8065), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n7856) );
  NAND2_X1 U10180 ( .A1(n12007), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7855) );
  INV_X1 U10181 ( .A(n7851), .ZN(n7849) );
  NAND2_X1 U10182 ( .A1(n7849), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7872) );
  INV_X1 U10183 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7850) );
  NAND2_X1 U10184 ( .A1(n7851), .A2(n7850), .ZN(n7852) );
  AND2_X1 U10185 ( .A1(n7872), .A2(n7852), .ZN(n10577) );
  NAND2_X1 U10186 ( .A1(n7997), .A2(n10577), .ZN(n7854) );
  NAND2_X1 U10187 ( .A1(n12008), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7853) );
  NAND4_X1 U10188 ( .A1(n7856), .A2(n7855), .A3(n7854), .A4(n7853), .ZN(n12938) );
  INV_X1 U10189 ( .A(n12938), .ZN(n7858) );
  AND2_X1 U10190 ( .A1(n11890), .A2(n7858), .ZN(n7857) );
  MUX2_X1 U10191 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n9371), .Z(n7861) );
  NAND2_X1 U10192 ( .A1(n7861), .A2(SI_8_), .ZN(n7879) );
  OAI21_X1 U10193 ( .B1(n7861), .B2(SI_8_), .A(n7879), .ZN(n7862) );
  INV_X1 U10194 ( .A(n7862), .ZN(n7863) );
  OR2_X1 U10195 ( .A1(n7864), .A2(n7863), .ZN(n7865) );
  NAND2_X1 U10196 ( .A1(n7880), .A2(n7865), .ZN(n9707) );
  OR2_X1 U10197 ( .A1(n9707), .A2(n8209), .ZN(n7869) );
  OR2_X1 U10198 ( .A1(n7866), .A2(n8268), .ZN(n7867) );
  XNOR2_X1 U10199 ( .A(n7867), .B(P2_IR_REG_8__SCAN_IN), .ZN(n14740) );
  AOI22_X1 U10200 ( .A1(n8079), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8078), .B2(
        n14740), .ZN(n7868) );
  NAND2_X1 U10201 ( .A1(n8281), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7877) );
  NAND2_X1 U10202 ( .A1(n8065), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n7876) );
  INV_X1 U10203 ( .A(n7872), .ZN(n7870) );
  NAND2_X1 U10204 ( .A1(n7870), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7893) );
  INV_X1 U10205 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7871) );
  NAND2_X1 U10206 ( .A1(n7872), .A2(n7871), .ZN(n7873) );
  AND2_X1 U10207 ( .A1(n7893), .A2(n7873), .ZN(n10989) );
  NAND2_X1 U10208 ( .A1(n7997), .A2(n10989), .ZN(n7875) );
  NAND2_X1 U10209 ( .A1(n12008), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7874) );
  NAND4_X1 U10210 ( .A1(n7877), .A2(n7876), .A3(n7875), .A4(n7874), .ZN(n12937) );
  INV_X1 U10211 ( .A(n12937), .ZN(n7878) );
  INV_X1 U10212 ( .A(n11895), .ZN(n14909) );
  MUX2_X1 U10213 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n8205), .Z(n7881) );
  NAND2_X1 U10214 ( .A1(n7881), .A2(SI_9_), .ZN(n7900) );
  OAI21_X1 U10215 ( .B1(n7881), .B2(SI_9_), .A(n7900), .ZN(n7882) );
  INV_X1 U10216 ( .A(n7882), .ZN(n7883) );
  OR2_X1 U10217 ( .A1(n7884), .A2(n7883), .ZN(n7885) );
  NAND2_X1 U10218 ( .A1(n7901), .A2(n7885), .ZN(n9742) );
  OR2_X1 U10219 ( .A1(n9742), .A2(n8209), .ZN(n7891) );
  NAND2_X1 U10220 ( .A1(n7866), .A2(n7886), .ZN(n7888) );
  NAND2_X1 U10221 ( .A1(n7888), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7887) );
  MUX2_X1 U10222 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7887), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n7889) );
  AND2_X1 U10223 ( .A1(n7889), .A2(n8037), .ZN(n9776) );
  AOI22_X1 U10224 ( .A1(n8079), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n8078), .B2(
        n9776), .ZN(n7890) );
  NAND2_X1 U10225 ( .A1(n12007), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7898) );
  NAND2_X1 U10226 ( .A1(n8065), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7897) );
  NAND2_X1 U10227 ( .A1(n7893), .A2(n7892), .ZN(n7894) );
  AND2_X1 U10228 ( .A1(n7911), .A2(n7894), .ZN(n10846) );
  NAND2_X1 U10229 ( .A1(n7997), .A2(n10846), .ZN(n7896) );
  NAND2_X1 U10230 ( .A1(n12008), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7895) );
  NAND4_X1 U10231 ( .A1(n7898), .A2(n7897), .A3(n7896), .A4(n7895), .ZN(n12936) );
  INV_X1 U10232 ( .A(n12936), .ZN(n11907) );
  XNOR2_X1 U10233 ( .A(n11905), .B(n11907), .ZN(n12080) );
  OR2_X1 U10234 ( .A1(n11905), .A2(n11907), .ZN(n7899) );
  MUX2_X1 U10235 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n8205), .Z(n7902) );
  NAND2_X1 U10236 ( .A1(n7902), .A2(SI_10_), .ZN(n7918) );
  OAI21_X1 U10237 ( .B1(n7902), .B2(SI_10_), .A(n7918), .ZN(n7903) );
  INV_X1 U10238 ( .A(n7903), .ZN(n7904) );
  NAND2_X1 U10239 ( .A1(n7919), .A2(n7905), .ZN(n9791) );
  NAND2_X1 U10240 ( .A1(n8037), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7906) );
  XNOR2_X1 U10241 ( .A(n7906), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10069) );
  AOI22_X1 U10242 ( .A1(n8079), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n8078), 
        .B2(n10069), .ZN(n7907) );
  NAND2_X1 U10243 ( .A1(n8281), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7916) );
  INV_X1 U10244 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7910) );
  NAND2_X1 U10245 ( .A1(n7911), .A2(n7910), .ZN(n7912) );
  AND2_X1 U10246 ( .A1(n7941), .A2(n7912), .ZN(n10969) );
  NAND2_X1 U10247 ( .A1(n7997), .A2(n10969), .ZN(n7915) );
  NAND2_X1 U10248 ( .A1(n8282), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n7914) );
  NAND2_X1 U10249 ( .A1(n12008), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7913) );
  NAND2_X1 U10250 ( .A1(n11910), .A2(n11909), .ZN(n10960) );
  NAND2_X1 U10251 ( .A1(n7917), .A2(n10960), .ZN(n11103) );
  MUX2_X1 U10252 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n8205), .Z(n7928) );
  XNOR2_X1 U10253 ( .A(n7928), .B(SI_11_), .ZN(n7931) );
  XNOR2_X1 U10254 ( .A(n7932), .B(n7931), .ZN(n9885) );
  NAND2_X1 U10255 ( .A1(n9885), .A2(n12011), .ZN(n7922) );
  NOR2_X1 U10256 ( .A1(n8037), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n7934) );
  OR2_X1 U10257 ( .A1(n7934), .A2(n8268), .ZN(n7920) );
  XNOR2_X1 U10258 ( .A(n7920), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10073) );
  AOI22_X1 U10259 ( .A1(n8079), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n8078), 
        .B2(n10073), .ZN(n7921) );
  NAND2_X1 U10260 ( .A1(n12007), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7926) );
  NAND2_X1 U10261 ( .A1(n8065), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n7925) );
  XNOR2_X1 U10262 ( .A(n7941), .B(P2_REG3_REG_11__SCAN_IN), .ZN(n11109) );
  NAND2_X1 U10263 ( .A1(n7997), .A2(n11109), .ZN(n7924) );
  NAND2_X1 U10264 ( .A1(n12008), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7923) );
  NAND4_X1 U10265 ( .A1(n7926), .A2(n7925), .A3(n7924), .A4(n7923), .ZN(n12934) );
  INV_X1 U10266 ( .A(n12934), .ZN(n11921) );
  XNOR2_X1 U10267 ( .A(n11919), .B(n11921), .ZN(n12082) );
  NAND2_X1 U10268 ( .A1(n11919), .A2(n11921), .ZN(n7927) );
  INV_X1 U10269 ( .A(n7928), .ZN(n7929) );
  NAND2_X1 U10270 ( .A1(n7929), .A2(n15428), .ZN(n7930) );
  MUX2_X1 U10271 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(P1_DATAO_REG_12__SCAN_IN), 
        .S(n8205), .Z(n7951) );
  XNOR2_X1 U10272 ( .A(n7951), .B(n15490), .ZN(n7949) );
  XNOR2_X1 U10273 ( .A(n7950), .B(n7949), .ZN(n10040) );
  NAND2_X1 U10274 ( .A1(n10040), .A2(n12011), .ZN(n7937) );
  AND2_X1 U10275 ( .A1(n7934), .A2(n7933), .ZN(n7954) );
  OR2_X1 U10276 ( .A1(n7954), .A2(n8268), .ZN(n7935) );
  XNOR2_X1 U10277 ( .A(n7935), .B(P2_IR_REG_12__SCAN_IN), .ZN(n14786) );
  AOI22_X1 U10278 ( .A1(n8079), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8078), 
        .B2(n14786), .ZN(n7936) );
  NAND2_X1 U10279 ( .A1(n8281), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7946) );
  NAND2_X1 U10280 ( .A1(n8282), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n7945) );
  INV_X1 U10281 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7939) );
  INV_X1 U10282 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7938) );
  OAI21_X1 U10283 ( .B1(n7941), .B2(n7939), .A(n7938), .ZN(n7942) );
  NAND2_X1 U10284 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_REG3_REG_12__SCAN_IN), 
        .ZN(n7940) );
  AND2_X1 U10285 ( .A1(n7942), .A2(n7963), .ZN(n11189) );
  NAND2_X1 U10286 ( .A1(n7997), .A2(n11189), .ZN(n7944) );
  NAND2_X1 U10287 ( .A1(n12008), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7943) );
  NAND4_X1 U10288 ( .A1(n7946), .A2(n7945), .A3(n7944), .A4(n7943), .ZN(n12933) );
  INV_X1 U10289 ( .A(n12933), .ZN(n7948) );
  XNOR2_X1 U10290 ( .A(n14329), .B(n7948), .ZN(n12085) );
  INV_X1 U10291 ( .A(n12085), .ZN(n7947) );
  INV_X1 U10292 ( .A(n7951), .ZN(n7952) );
  MUX2_X1 U10293 ( .A(n8410), .B(n10091), .S(n8205), .Z(n7973) );
  XNOR2_X1 U10294 ( .A(n7973), .B(SI_13_), .ZN(n7970) );
  XNOR2_X1 U10295 ( .A(n7971), .B(n7970), .ZN(n10059) );
  NAND2_X1 U10296 ( .A1(n10059), .A2(n12011), .ZN(n7961) );
  INV_X1 U10297 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n7953) );
  AND2_X1 U10298 ( .A1(n7954), .A2(n7953), .ZN(n7958) );
  NOR2_X1 U10299 ( .A1(n7958), .A2(n8268), .ZN(n7955) );
  MUX2_X1 U10300 ( .A(n8268), .B(n7955), .S(P2_IR_REG_13__SCAN_IN), .Z(n7956)
         );
  INV_X1 U10301 ( .A(n7956), .ZN(n7959) );
  INV_X1 U10302 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n7957) );
  NAND2_X1 U10303 ( .A1(n7958), .A2(n7957), .ZN(n7990) );
  AOI22_X1 U10304 ( .A1(n8079), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n10335), 
        .B2(n8078), .ZN(n7960) );
  NAND2_X1 U10305 ( .A1(n12007), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7968) );
  NAND2_X1 U10306 ( .A1(n8282), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n7967) );
  INV_X1 U10307 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n11299) );
  NAND2_X1 U10308 ( .A1(n7963), .A2(n11299), .ZN(n7964) );
  AND2_X1 U10309 ( .A1(n7978), .A2(n7964), .ZN(n11302) );
  NAND2_X1 U10310 ( .A1(n7997), .A2(n11302), .ZN(n7966) );
  NAND2_X1 U10311 ( .A1(n12008), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7965) );
  NAND4_X1 U10312 ( .A1(n7968), .A2(n7967), .A3(n7966), .A4(n7965), .ZN(n12932) );
  INV_X1 U10313 ( .A(n12932), .ZN(n11245) );
  NAND2_X1 U10314 ( .A1(n11934), .A2(n11245), .ZN(n7969) );
  INV_X1 U10315 ( .A(SI_13_), .ZN(n7972) );
  NAND2_X1 U10316 ( .A1(n7973), .A2(n7972), .ZN(n7974) );
  INV_X1 U10317 ( .A(SI_14_), .ZN(n9738) );
  XNOR2_X1 U10318 ( .A(n8007), .B(n9738), .ZN(n7987) );
  MUX2_X1 U10319 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n8205), .Z(n8008) );
  XNOR2_X1 U10320 ( .A(n7987), .B(n8008), .ZN(n10367) );
  NAND2_X1 U10321 ( .A1(n10367), .A2(n12011), .ZN(n7977) );
  NAND2_X1 U10322 ( .A1(n7990), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7975) );
  XNOR2_X1 U10323 ( .A(n7975), .B(P2_IR_REG_14__SCAN_IN), .ZN(n10732) );
  AOI22_X1 U10324 ( .A1(n8079), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8078), 
        .B2(n10732), .ZN(n7976) );
  NAND2_X1 U10325 ( .A1(n8282), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n7983) );
  NAND2_X1 U10326 ( .A1(n7978), .A2(n11405), .ZN(n7979) );
  AND2_X1 U10327 ( .A1(n7995), .A2(n7979), .ZN(n14306) );
  NAND2_X1 U10328 ( .A1(n7997), .A2(n14306), .ZN(n7982) );
  NAND2_X1 U10329 ( .A1(n8281), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7981) );
  NAND2_X1 U10330 ( .A1(n12008), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7980) );
  NAND4_X1 U10331 ( .A1(n7983), .A2(n7982), .A3(n7981), .A4(n7980), .ZN(n12931) );
  INV_X1 U10332 ( .A(n12931), .ZN(n7984) );
  AND2_X1 U10333 ( .A1(n14308), .A2(n7984), .ZN(n7985) );
  INV_X1 U10334 ( .A(n8007), .ZN(n7986) );
  OAI22_X1 U10335 ( .A1(n7987), .A2(n8008), .B1(n7986), .B2(SI_14_), .ZN(n7989) );
  MUX2_X1 U10336 ( .A(n10519), .B(n10521), .S(n8205), .Z(n8009) );
  XNOR2_X1 U10337 ( .A(n8009), .B(SI_15_), .ZN(n7988) );
  XNOR2_X1 U10338 ( .A(n7989), .B(n7988), .ZN(n10518) );
  NAND2_X1 U10339 ( .A1(n10518), .A2(n12011), .ZN(n7993) );
  NAND2_X1 U10340 ( .A1(n7991), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8014) );
  XNOR2_X1 U10341 ( .A(n8014), .B(P2_IR_REG_15__SCAN_IN), .ZN(n12970) );
  AOI22_X1 U10342 ( .A1(n8079), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n12970), 
        .B2(n8078), .ZN(n7992) );
  NAND2_X1 U10343 ( .A1(n12007), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8001) );
  NAND2_X1 U10344 ( .A1(n8282), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n8000) );
  INV_X1 U10345 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n7994) );
  NAND2_X1 U10346 ( .A1(n7995), .A2(n7994), .ZN(n7996) );
  AND2_X1 U10347 ( .A1(n8022), .A2(n7996), .ZN(n13207) );
  NAND2_X1 U10348 ( .A1(n7997), .A2(n13207), .ZN(n7999) );
  NAND2_X1 U10349 ( .A1(n12008), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n7998) );
  NAND4_X1 U10350 ( .A1(n8001), .A2(n8000), .A3(n7999), .A4(n7998), .ZN(n12930) );
  INV_X1 U10351 ( .A(n12930), .ZN(n11943) );
  XNOR2_X1 U10352 ( .A(n13336), .B(n11943), .ZN(n13208) );
  INV_X1 U10353 ( .A(n13208), .ZN(n8002) );
  NAND2_X1 U10354 ( .A1(n13203), .A2(n8002), .ZN(n8004) );
  OR2_X1 U10355 ( .A1(n13336), .A2(n11943), .ZN(n8003) );
  INV_X1 U10356 ( .A(n8009), .ZN(n8005) );
  NAND2_X1 U10357 ( .A1(n8005), .A2(SI_15_), .ZN(n8010) );
  NAND2_X1 U10358 ( .A1(n8008), .A2(SI_14_), .ZN(n8006) );
  NOR2_X1 U10359 ( .A1(n8008), .A2(SI_14_), .ZN(n8011) );
  INV_X1 U10360 ( .A(SI_15_), .ZN(n9751) );
  AOI22_X1 U10361 ( .A1(n8011), .A2(n8010), .B1(n8009), .B2(n9751), .ZN(n8012)
         );
  MUX2_X1 U10362 ( .A(n8418), .B(n15311), .S(n8205), .Z(n8033) );
  XNOR2_X1 U10363 ( .A(n8033), .B(SI_16_), .ZN(n8030) );
  XNOR2_X1 U10364 ( .A(n8031), .B(n8030), .ZN(n10344) );
  NAND2_X1 U10365 ( .A1(n10344), .A2(n12011), .ZN(n8020) );
  INV_X1 U10366 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n8013) );
  NAND2_X1 U10367 ( .A1(n8014), .A2(n8013), .ZN(n8015) );
  NAND2_X1 U10368 ( .A1(n8015), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8017) );
  INV_X1 U10369 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8016) );
  XNOR2_X1 U10370 ( .A(n8017), .B(n8016), .ZN(n14801) );
  OAI22_X1 U10371 ( .A1(n14801), .A2(n9642), .B1(n12013), .B2(n15311), .ZN(
        n8018) );
  INV_X1 U10372 ( .A(n8018), .ZN(n8019) );
  INV_X1 U10373 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n12836) );
  NAND2_X1 U10374 ( .A1(n8022), .A2(n12836), .ZN(n8023) );
  NAND2_X1 U10375 ( .A1(n8042), .A2(n8023), .ZN(n13193) );
  INV_X1 U10376 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n15405) );
  OAI22_X1 U10377 ( .A1(n13193), .A2(n8229), .B1(n8262), .B2(n15405), .ZN(
        n8027) );
  INV_X1 U10378 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8025) );
  INV_X1 U10379 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8024) );
  OAI22_X1 U10380 ( .A1(n7773), .A2(n8025), .B1(n7792), .B2(n8024), .ZN(n8026)
         );
  INV_X1 U10381 ( .A(n12929), .ZN(n8028) );
  NAND2_X1 U10382 ( .A1(n13294), .A2(n8028), .ZN(n13166) );
  OR2_X1 U10383 ( .A1(n13294), .A2(n8028), .ZN(n8029) );
  NAND2_X1 U10384 ( .A1(n13166), .A2(n8029), .ZN(n13198) );
  NAND2_X1 U10385 ( .A1(n8031), .A2(n8030), .ZN(n8035) );
  NAND2_X1 U10386 ( .A1(n8033), .A2(n8032), .ZN(n8034) );
  MUX2_X1 U10387 ( .A(n15494), .B(n10524), .S(n8205), .Z(n8054) );
  XNOR2_X1 U10388 ( .A(n8054), .B(SI_17_), .ZN(n8051) );
  XNOR2_X1 U10389 ( .A(n8052), .B(n8051), .ZN(n10522) );
  NAND2_X1 U10390 ( .A1(n10522), .A2(n12011), .ZN(n8040) );
  OAI21_X1 U10391 ( .B1(n8037), .B2(n8036), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n8038) );
  XNOR2_X1 U10392 ( .A(n8038), .B(P2_IR_REG_17__SCAN_IN), .ZN(n14808) );
  AOI22_X1 U10393 ( .A1(n8079), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8078), 
        .B2(n14808), .ZN(n8039) );
  INV_X1 U10394 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n12967) );
  INV_X1 U10395 ( .A(n8042), .ZN(n8041) );
  INV_X1 U10396 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n14802) );
  NAND2_X1 U10397 ( .A1(n8042), .A2(n14802), .ZN(n8043) );
  NAND2_X1 U10398 ( .A1(n8063), .A2(n8043), .ZN(n12847) );
  OR2_X1 U10399 ( .A1(n12847), .A2(n8229), .ZN(n8047) );
  NAND2_X1 U10400 ( .A1(n12007), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8045) );
  NAND2_X1 U10401 ( .A1(n8282), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n8044) );
  AND2_X1 U10402 ( .A1(n8045), .A2(n8044), .ZN(n8046) );
  OAI211_X1 U10403 ( .C1(n8262), .C2(n12967), .A(n8047), .B(n8046), .ZN(n12928) );
  INV_X1 U10404 ( .A(n12928), .ZN(n8049) );
  XNOR2_X1 U10405 ( .A(n13289), .B(n8049), .ZN(n13167) );
  INV_X1 U10406 ( .A(n13167), .ZN(n8048) );
  NAND2_X1 U10407 ( .A1(n13289), .A2(n8049), .ZN(n8050) );
  INV_X1 U10408 ( .A(SI_17_), .ZN(n8053) );
  NAND2_X1 U10409 ( .A1(n8054), .A2(n8053), .ZN(n8055) );
  NAND2_X1 U10410 ( .A1(n8099), .A2(n15288), .ZN(n8056) );
  NAND2_X1 U10411 ( .A1(n8070), .A2(n8056), .ZN(n8057) );
  MUX2_X1 U10412 ( .A(n10725), .B(n15387), .S(n8205), .Z(n8094) );
  NAND2_X1 U10413 ( .A1(n8057), .A2(n8094), .ZN(n8058) );
  XNOR2_X1 U10414 ( .A(n8060), .B(P2_IR_REG_18__SCAN_IN), .ZN(n12975) );
  AOI22_X1 U10415 ( .A1(n8079), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8078), 
        .B2(n12975), .ZN(n8061) );
  NAND2_X1 U10416 ( .A1(n8063), .A2(n14818), .ZN(n8064) );
  NAND2_X1 U10417 ( .A1(n8084), .A2(n8064), .ZN(n12880) );
  AOI22_X1 U10418 ( .A1(n12007), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n8065), 
        .B2(P2_REG0_REG_18__SCAN_IN), .ZN(n8067) );
  NAND2_X1 U10419 ( .A1(n12008), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8066) );
  OAI211_X1 U10420 ( .C1(n12880), .C2(n8229), .A(n8067), .B(n8066), .ZN(n12927) );
  INV_X1 U10421 ( .A(n12927), .ZN(n12809) );
  AND2_X1 U10422 ( .A1(n13283), .A2(n12809), .ZN(n8068) );
  OR2_X1 U10423 ( .A1(n13283), .A2(n12809), .ZN(n8069) );
  NAND2_X1 U10424 ( .A1(n8071), .A2(n8070), .ZN(n8072) );
  MUX2_X1 U10425 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n8205), .Z(n8100) );
  XNOR2_X1 U10426 ( .A(n8100), .B(SI_19_), .ZN(n8096) );
  NAND2_X1 U10427 ( .A1(n10920), .A2(n12011), .ZN(n8081) );
  INV_X1 U10428 ( .A(n8076), .ZN(n8073) );
  NAND2_X1 U10429 ( .A1(n8073), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8074) );
  MUX2_X1 U10430 ( .A(n8074), .B(P2_IR_REG_31__SCAN_IN), .S(n8075), .Z(n8077)
         );
  AOI22_X1 U10431 ( .A1(n8079), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8078), 
        .B2(n13195), .ZN(n8080) );
  INV_X1 U10432 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8083) );
  NAND2_X1 U10433 ( .A1(n8084), .A2(n8083), .ZN(n8085) );
  NAND2_X1 U10434 ( .A1(n8110), .A2(n8085), .ZN(n13140) );
  OR2_X1 U10435 ( .A1(n13140), .A2(n8229), .ZN(n8090) );
  INV_X1 U10436 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n15340) );
  NAND2_X1 U10437 ( .A1(n8282), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8087) );
  NAND2_X1 U10438 ( .A1(n12008), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8086) );
  OAI211_X1 U10439 ( .C1(n7773), .C2(n15340), .A(n8087), .B(n8086), .ZN(n8088)
         );
  INV_X1 U10440 ( .A(n8088), .ZN(n8089) );
  NAND2_X1 U10441 ( .A1(n8090), .A2(n8089), .ZN(n12926) );
  INV_X1 U10442 ( .A(n12926), .ZN(n11973) );
  NAND2_X1 U10443 ( .A1(n13278), .A2(n11973), .ZN(n8092) );
  NOR2_X1 U10444 ( .A1(n13278), .A2(n11973), .ZN(n8091) );
  INV_X1 U10445 ( .A(n8094), .ZN(n8093) );
  NOR2_X1 U10446 ( .A1(n8093), .A2(SI_18_), .ZN(n8098) );
  NOR2_X1 U10447 ( .A1(n8094), .A2(n15288), .ZN(n8095) );
  NOR2_X1 U10448 ( .A1(n8096), .A2(n8095), .ZN(n8097) );
  INV_X1 U10449 ( .A(n8100), .ZN(n8101) );
  NAND2_X1 U10450 ( .A1(n8102), .A2(n10325), .ZN(n8103) );
  INV_X1 U10451 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n10782) );
  MUX2_X1 U10452 ( .A(n11827), .B(n10782), .S(n8205), .Z(n8105) );
  NAND2_X1 U10453 ( .A1(n8106), .A2(n8105), .ZN(n8107) );
  NAND2_X1 U10454 ( .A1(n8121), .A2(n8107), .ZN(n11826) );
  OR2_X1 U10455 ( .A1(n11826), .A2(n8209), .ZN(n8109) );
  OR2_X1 U10456 ( .A1(n12013), .A2(n10782), .ZN(n8108) );
  INV_X1 U10457 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n12864) );
  NAND2_X1 U10458 ( .A1(n8110), .A2(n12864), .ZN(n8111) );
  AND2_X1 U10459 ( .A1(n8130), .A2(n8111), .ZN(n13127) );
  NAND2_X1 U10460 ( .A1(n13127), .A2(n7997), .ZN(n8117) );
  INV_X1 U10461 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8114) );
  NAND2_X1 U10462 ( .A1(n8281), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8113) );
  NAND2_X1 U10463 ( .A1(n8282), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n8112) );
  OAI211_X1 U10464 ( .C1(n8114), .C2(n8262), .A(n8113), .B(n8112), .ZN(n8115)
         );
  INV_X1 U10465 ( .A(n8115), .ZN(n8116) );
  NAND2_X1 U10466 ( .A1(n8117), .A2(n8116), .ZN(n12925) );
  INV_X1 U10467 ( .A(n12925), .ZN(n12810) );
  NAND2_X1 U10468 ( .A1(n13273), .A2(n12810), .ZN(n8119) );
  OR2_X1 U10469 ( .A1(n13273), .A2(n12810), .ZN(n8118) );
  NAND2_X1 U10470 ( .A1(n8119), .A2(n8118), .ZN(n12089) );
  MUX2_X1 U10471 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n8205), .Z(n8122) );
  OAI21_X1 U10472 ( .B1(n8122), .B2(SI_21_), .A(n8138), .ZN(n8123) );
  INV_X1 U10473 ( .A(n8123), .ZN(n8124) );
  OR2_X1 U10474 ( .A1(n8125), .A2(n8124), .ZN(n8126) );
  NAND2_X1 U10475 ( .A1(n8139), .A2(n8126), .ZN(n10999) );
  INV_X1 U10476 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11000) );
  OR2_X1 U10477 ( .A1(n12013), .A2(n11000), .ZN(n8127) );
  INV_X1 U10478 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n12820) );
  NAND2_X1 U10479 ( .A1(n8130), .A2(n12820), .ZN(n8131) );
  NAND2_X1 U10480 ( .A1(n8143), .A2(n8131), .ZN(n13107) );
  OR2_X1 U10481 ( .A1(n13107), .A2(n8229), .ZN(n8136) );
  INV_X1 U10482 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n15473) );
  NAND2_X1 U10483 ( .A1(n8281), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8133) );
  NAND2_X1 U10484 ( .A1(n12008), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8132) );
  OAI211_X1 U10485 ( .C1(n7792), .C2(n15473), .A(n8133), .B(n8132), .ZN(n8134)
         );
  INV_X1 U10486 ( .A(n8134), .ZN(n8135) );
  NAND2_X1 U10487 ( .A1(n8136), .A2(n8135), .ZN(n12924) );
  INV_X1 U10488 ( .A(n12924), .ZN(n11982) );
  OR2_X1 U10489 ( .A1(n13270), .A2(n11982), .ZN(n8137) );
  MUX2_X1 U10490 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n8205), .Z(n8152) );
  XNOR2_X1 U10491 ( .A(n9372), .B(n8152), .ZN(n11175) );
  NAND2_X1 U10492 ( .A1(n11175), .A2(n12011), .ZN(n8141) );
  INV_X1 U10493 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11177) );
  OR2_X1 U10494 ( .A1(n12013), .A2(n11177), .ZN(n8140) );
  INV_X1 U10495 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8142) );
  NAND2_X1 U10496 ( .A1(n8143), .A2(n8142), .ZN(n8144) );
  AND2_X1 U10497 ( .A1(n8161), .A2(n8144), .ZN(n13097) );
  NAND2_X1 U10498 ( .A1(n13097), .A2(n7997), .ZN(n8149) );
  INV_X1 U10499 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n15487) );
  NAND2_X1 U10500 ( .A1(n12008), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8146) );
  NAND2_X1 U10501 ( .A1(n8282), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8145) );
  OAI211_X1 U10502 ( .C1(n7773), .C2(n15487), .A(n8146), .B(n8145), .ZN(n8147)
         );
  INV_X1 U10503 ( .A(n8147), .ZN(n8148) );
  NAND2_X1 U10504 ( .A1(n8149), .A2(n8148), .ZN(n12923) );
  NAND2_X1 U10505 ( .A1(n13262), .A2(n12923), .ZN(n8329) );
  OR2_X1 U10506 ( .A1(n13262), .A2(n12923), .ZN(n8150) );
  NAND2_X1 U10507 ( .A1(n8329), .A2(n8150), .ZN(n12091) );
  INV_X1 U10508 ( .A(n12923), .ZN(n12801) );
  OR2_X1 U10509 ( .A1(n13262), .A2(n12801), .ZN(n8151) );
  INV_X1 U10510 ( .A(SI_22_), .ZN(n8858) );
  NOR2_X1 U10511 ( .A1(n8154), .A2(n8858), .ZN(n8153) );
  NAND2_X1 U10512 ( .A1(n8154), .A2(n8858), .ZN(n8155) );
  INV_X1 U10513 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11307) );
  INV_X1 U10514 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11311) );
  MUX2_X1 U10515 ( .A(n11307), .B(n11311), .S(n8205), .Z(n8156) );
  NAND2_X1 U10516 ( .A1(n8169), .A2(n8170), .ZN(n8158) );
  NAND2_X1 U10517 ( .A1(n11308), .A2(n12011), .ZN(n8160) );
  OR2_X1 U10518 ( .A1(n12013), .A2(n11311), .ZN(n8159) );
  INV_X1 U10519 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n12802) );
  NAND2_X1 U10520 ( .A1(n8161), .A2(n12802), .ZN(n8162) );
  NAND2_X1 U10521 ( .A1(n8178), .A2(n8162), .ZN(n13078) );
  INV_X1 U10522 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n13082) );
  NAND2_X1 U10523 ( .A1(n12007), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8164) );
  NAND2_X1 U10524 ( .A1(n8282), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8163) );
  OAI211_X1 U10525 ( .C1(n13082), .C2(n8262), .A(n8164), .B(n8163), .ZN(n8165)
         );
  INV_X1 U10526 ( .A(n8165), .ZN(n8166) );
  OAI21_X1 U10527 ( .B1(n13078), .B2(n8229), .A(n8166), .ZN(n12922) );
  INV_X1 U10528 ( .A(n12922), .ZN(n12854) );
  XNOR2_X1 U10529 ( .A(n13257), .B(n12854), .ZN(n13074) );
  NAND2_X1 U10530 ( .A1(n6677), .A2(n8167), .ZN(n13075) );
  NAND2_X1 U10531 ( .A1(n13257), .A2(n12854), .ZN(n8168) );
  INV_X1 U10532 ( .A(SI_23_), .ZN(n10647) );
  MUX2_X1 U10533 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n8205), .Z(n8171) );
  NAND2_X1 U10534 ( .A1(n8171), .A2(SI_24_), .ZN(n8186) );
  OAI21_X1 U10535 ( .B1(n8171), .B2(SI_24_), .A(n8186), .ZN(n8172) );
  NAND2_X1 U10536 ( .A1(n8173), .A2(n8172), .ZN(n8174) );
  NAND2_X1 U10537 ( .A1(n8187), .A2(n8174), .ZN(n11334) );
  INV_X1 U10538 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11333) );
  OR2_X1 U10539 ( .A1(n12013), .A2(n11333), .ZN(n8175) );
  INV_X1 U10540 ( .A(n8178), .ZN(n8177) );
  NAND2_X1 U10541 ( .A1(n8177), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n8191) );
  INV_X1 U10542 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n12855) );
  NAND2_X1 U10543 ( .A1(n8178), .A2(n12855), .ZN(n8179) );
  AND2_X1 U10544 ( .A1(n8191), .A2(n8179), .ZN(n13067) );
  NAND2_X1 U10545 ( .A1(n13067), .A2(n7997), .ZN(n8184) );
  INV_X1 U10546 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n13253) );
  NAND2_X1 U10547 ( .A1(n7832), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8181) );
  NAND2_X1 U10548 ( .A1(n8282), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8180) );
  OAI211_X1 U10549 ( .C1(n7773), .C2(n13253), .A(n8181), .B(n8180), .ZN(n8182)
         );
  INV_X1 U10550 ( .A(n8182), .ZN(n8183) );
  NAND2_X1 U10551 ( .A1(n8184), .A2(n8183), .ZN(n12921) );
  INV_X1 U10552 ( .A(n13058), .ZN(n13063) );
  NAND2_X1 U10553 ( .A1(n13066), .A2(n12827), .ZN(n8185) );
  MUX2_X1 U10554 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n8205), .Z(n8200) );
  XNOR2_X1 U10555 ( .A(n8200), .B(SI_25_), .ZN(n8201) );
  XNOR2_X1 U10556 ( .A(n8202), .B(n8201), .ZN(n11460) );
  NAND2_X1 U10557 ( .A1(n11460), .A2(n12011), .ZN(n8189) );
  INV_X1 U10558 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n11462) );
  OR2_X1 U10559 ( .A1(n12013), .A2(n11462), .ZN(n8188) );
  INV_X1 U10560 ( .A(n8191), .ZN(n8190) );
  NAND2_X1 U10561 ( .A1(n8190), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n8212) );
  INV_X1 U10562 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n12829) );
  NAND2_X1 U10563 ( .A1(n8191), .A2(n12829), .ZN(n8192) );
  NAND2_X1 U10564 ( .A1(n8212), .A2(n8192), .ZN(n13053) );
  INV_X1 U10565 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n13052) );
  NAND2_X1 U10566 ( .A1(n8281), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8194) );
  NAND2_X1 U10567 ( .A1(n8282), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8193) );
  OAI211_X1 U10568 ( .C1(n13052), .C2(n8262), .A(n8194), .B(n8193), .ZN(n8195)
         );
  INV_X1 U10569 ( .A(n8195), .ZN(n8196) );
  XNOR2_X1 U10570 ( .A(n13248), .B(n12890), .ZN(n12093) );
  OR2_X1 U10571 ( .A1(n13319), .A2(n12920), .ZN(n8198) );
  NAND2_X1 U10572 ( .A1(n8199), .A2(n8198), .ZN(n13029) );
  NAND2_X1 U10573 ( .A1(n8203), .A2(n11136), .ZN(n8204) );
  INV_X1 U10574 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14040) );
  INV_X1 U10575 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13358) );
  MUX2_X1 U10576 ( .A(n14040), .B(n13358), .S(n8205), .Z(n8206) );
  NAND2_X1 U10577 ( .A1(n8207), .A2(n8206), .ZN(n8208) );
  OR2_X1 U10578 ( .A1(n12013), .A2(n13358), .ZN(n8210) );
  INV_X1 U10579 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n12893) );
  NAND2_X1 U10580 ( .A1(n8212), .A2(n12893), .ZN(n8213) );
  NAND2_X1 U10581 ( .A1(n13034), .A2(n7997), .ZN(n8219) );
  INV_X1 U10582 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8216) );
  NAND2_X1 U10583 ( .A1(n12007), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8215) );
  NAND2_X1 U10584 ( .A1(n8282), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8214) );
  OAI211_X1 U10585 ( .C1(n8216), .C2(n8262), .A(n8215), .B(n8214), .ZN(n8217)
         );
  INV_X1 U10586 ( .A(n8217), .ZN(n8218) );
  XNOR2_X1 U10587 ( .A(n13238), .B(n12919), .ZN(n13037) );
  NAND2_X1 U10588 ( .A1(n13029), .A2(n13037), .ZN(n8221) );
  NAND2_X1 U10589 ( .A1(n13238), .A2(n12828), .ZN(n8220) );
  NAND2_X1 U10590 ( .A1(n8221), .A2(n8220), .ZN(n13015) );
  INV_X1 U10591 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n11831) );
  INV_X1 U10592 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13356) );
  MUX2_X1 U10593 ( .A(n11831), .B(n13356), .S(n8205), .Z(n8236) );
  INV_X1 U10594 ( .A(n8236), .ZN(n8239) );
  XNOR2_X1 U10595 ( .A(n8239), .B(SI_27_), .ZN(n8224) );
  NAND2_X1 U10596 ( .A1(n11830), .A2(n12011), .ZN(n8226) );
  OR2_X1 U10597 ( .A1(n12013), .A2(n13356), .ZN(n8225) );
  INV_X1 U10598 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n12794) );
  NAND2_X1 U10599 ( .A1(n8227), .A2(n12794), .ZN(n8228) );
  NAND2_X1 U10600 ( .A1(n11832), .A2(n8228), .ZN(n13023) );
  INV_X1 U10601 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n13022) );
  NAND2_X1 U10602 ( .A1(n8281), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8231) );
  NAND2_X1 U10603 ( .A1(n8282), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8230) );
  OAI211_X1 U10604 ( .C1(n13022), .C2(n8262), .A(n8231), .B(n8230), .ZN(n8232)
         );
  INV_X1 U10605 ( .A(n8232), .ZN(n8233) );
  OR2_X1 U10606 ( .A1(n13019), .A2(n12918), .ZN(n8235) );
  INV_X1 U10607 ( .A(SI_27_), .ZN(n11179) );
  NAND2_X1 U10608 ( .A1(n8236), .A2(n11179), .ZN(n8237) );
  NAND2_X1 U10609 ( .A1(n8239), .A2(SI_27_), .ZN(n8240) );
  MUX2_X1 U10610 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n8205), .Z(n8254) );
  XNOR2_X1 U10611 ( .A(n8254), .B(SI_28_), .ZN(n8252) );
  NAND2_X1 U10612 ( .A1(n13351), .A2(n12011), .ZN(n8243) );
  OR2_X1 U10613 ( .A1(n12013), .A2(n13354), .ZN(n8242) );
  XNOR2_X1 U10614 ( .A(n11832), .B(P2_REG3_REG_28__SCAN_IN), .ZN(n12165) );
  NAND2_X1 U10615 ( .A1(n12165), .A2(n7997), .ZN(n8249) );
  INV_X1 U10616 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8246) );
  NAND2_X1 U10617 ( .A1(n12007), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8245) );
  NAND2_X1 U10618 ( .A1(n12008), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8244) );
  OAI211_X1 U10619 ( .C1(n7792), .C2(n8246), .A(n8245), .B(n8244), .ZN(n8247)
         );
  INV_X1 U10620 ( .A(n8247), .ZN(n8248) );
  NAND2_X1 U10621 ( .A1(n13229), .A2(n12793), .ZN(n8250) );
  INV_X1 U10622 ( .A(n8254), .ZN(n8255) );
  INV_X1 U10623 ( .A(SI_28_), .ZN(n11818) );
  NAND2_X1 U10624 ( .A1(n8255), .A2(n11818), .ZN(n8256) );
  INV_X1 U10625 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14035) );
  INV_X1 U10626 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13349) );
  MUX2_X1 U10627 ( .A(n14035), .B(n13349), .S(n8205), .Z(n9484) );
  XNOR2_X1 U10628 ( .A(n9484), .B(SI_29_), .ZN(n9482) );
  NAND2_X1 U10629 ( .A1(n13347), .A2(n12011), .ZN(n8258) );
  OR2_X1 U10630 ( .A1(n12013), .A2(n13349), .ZN(n8257) );
  NAND3_X1 U10631 ( .A1(n8259), .A2(n7997), .A3(P2_REG3_REG_28__SCAN_IN), .ZN(
        n8266) );
  INV_X1 U10632 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8263) );
  NAND2_X1 U10633 ( .A1(n8281), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8261) );
  NAND2_X1 U10634 ( .A1(n8282), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8260) );
  OAI211_X1 U10635 ( .C1(n8263), .C2(n8262), .A(n8261), .B(n8260), .ZN(n8264)
         );
  INV_X1 U10636 ( .A(n8264), .ZN(n8265) );
  NAND2_X1 U10637 ( .A1(n8266), .A2(n8265), .ZN(n12916) );
  INV_X1 U10638 ( .A(n12916), .ZN(n8267) );
  OR2_X1 U10639 ( .A1(n12066), .A2(n8343), .ZN(n8280) );
  NAND2_X1 U10640 ( .A1(n8277), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8276) );
  MUX2_X1 U10641 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8276), .S(
        P2_IR_REG_22__SCAN_IN), .Z(n8278) );
  INV_X1 U10642 ( .A(n8360), .ZN(n8369) );
  NAND2_X2 U10643 ( .A1(n8278), .A2(n8369), .ZN(n12058) );
  NAND2_X1 U10644 ( .A1(n12105), .A2(n13195), .ZN(n8279) );
  NAND2_X1 U10645 ( .A1(n8281), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8285) );
  NAND2_X1 U10646 ( .A1(n7832), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8284) );
  NAND2_X1 U10647 ( .A1(n8282), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8283) );
  INV_X1 U10648 ( .A(P2_B_REG_SCAN_IN), .ZN(n8289) );
  OR2_X1 U10649 ( .A1(n8288), .A2(n8289), .ZN(n8290) );
  NAND2_X1 U10650 ( .A1(n12902), .A2(n8290), .ZN(n12990) );
  INV_X1 U10651 ( .A(n8287), .ZN(n8291) );
  NAND2_X1 U10652 ( .A1(n12917), .A2(n12901), .ZN(n8292) );
  OAI21_X1 U10653 ( .B1(n12018), .B2(n12990), .A(n8292), .ZN(n8293) );
  INV_X1 U10654 ( .A(n12068), .ZN(n8298) );
  AND2_X1 U10655 ( .A1(n11843), .A2(n14882), .ZN(n9915) );
  INV_X1 U10656 ( .A(n12069), .ZN(n8295) );
  NAND2_X1 U10657 ( .A1(n10044), .A2(n8295), .ZN(n8297) );
  INV_X1 U10658 ( .A(n11851), .ZN(n14834) );
  NAND2_X1 U10659 ( .A1(n9877), .A2(n14834), .ZN(n8296) );
  NAND2_X1 U10660 ( .A1(n8297), .A2(n8296), .ZN(n10265) );
  NAND2_X1 U10661 ( .A1(n8298), .A2(n10265), .ZN(n8302) );
  INV_X1 U10662 ( .A(n14891), .ZN(n8299) );
  NAND2_X1 U10663 ( .A1(n8300), .A2(n8299), .ZN(n8301) );
  NAND2_X1 U10664 ( .A1(n8302), .A2(n8301), .ZN(n10369) );
  NAND2_X1 U10665 ( .A1(n8303), .A2(n10378), .ZN(n8304) );
  NAND2_X1 U10666 ( .A1(n11876), .A2(n12940), .ZN(n8305) );
  NAND2_X1 U10667 ( .A1(n8306), .A2(n8305), .ZN(n10598) );
  OR2_X1 U10668 ( .A1(n10598), .A2(n12075), .ZN(n10599) );
  OR2_X1 U10669 ( .A1(n11884), .A2(n12939), .ZN(n8307) );
  NAND2_X2 U10670 ( .A1(n10599), .A2(n8307), .ZN(n10570) );
  XNOR2_X1 U10671 ( .A(n11890), .B(n12938), .ZN(n12076) );
  OR2_X1 U10672 ( .A1(n11890), .A2(n12938), .ZN(n8308) );
  NAND2_X1 U10673 ( .A1(n11895), .A2(n12937), .ZN(n8310) );
  OR2_X1 U10674 ( .A1(n11895), .A2(n12937), .ZN(n8309) );
  NAND2_X1 U10675 ( .A1(n8310), .A2(n8309), .ZN(n12078) );
  NAND2_X1 U10676 ( .A1(n10840), .A2(n12080), .ZN(n8312) );
  NAND2_X1 U10677 ( .A1(n11905), .A2(n12936), .ZN(n8311) );
  AND2_X1 U10678 ( .A1(n11910), .A2(n12935), .ZN(n8313) );
  NOR2_X1 U10679 ( .A1(n11919), .A2(n12934), .ZN(n8314) );
  NOR2_X1 U10680 ( .A1(n11934), .A2(n12932), .ZN(n8315) );
  NAND2_X1 U10681 ( .A1(n11934), .A2(n12932), .ZN(n8316) );
  AND2_X1 U10682 ( .A1(n14308), .A2(n12931), .ZN(n8318) );
  OR2_X1 U10683 ( .A1(n14308), .A2(n12931), .ZN(n8319) );
  NOR2_X1 U10684 ( .A1(n13336), .A2(n12930), .ZN(n8320) );
  NAND2_X1 U10685 ( .A1(n13199), .A2(n13198), .ZN(n13292) );
  NAND2_X1 U10686 ( .A1(n13294), .A2(n12929), .ZN(n8321) );
  NAND2_X1 U10687 ( .A1(n13292), .A2(n8321), .ZN(n13165) );
  OR2_X1 U10688 ( .A1(n13289), .A2(n12928), .ZN(n8322) );
  NAND2_X1 U10689 ( .A1(n13289), .A2(n12928), .ZN(n8323) );
  XNOR2_X1 U10690 ( .A(n13283), .B(n12927), .ZN(n13161) );
  OR2_X1 U10691 ( .A1(n13283), .A2(n12927), .ZN(n8324) );
  NAND2_X1 U10692 ( .A1(n13278), .A2(n12926), .ZN(n12064) );
  OR2_X1 U10693 ( .A1(n13278), .A2(n12926), .ZN(n12065) );
  NAND2_X1 U10694 ( .A1(n13273), .A2(n12925), .ZN(n8325) );
  NAND2_X1 U10695 ( .A1(n8326), .A2(n8325), .ZN(n13114) );
  XNOR2_X1 U10696 ( .A(n13270), .B(n12924), .ZN(n13112) );
  OR2_X2 U10697 ( .A1(n13114), .A2(n13112), .ZN(n8328) );
  OR2_X1 U10698 ( .A1(n13270), .A2(n12924), .ZN(n8327) );
  NAND2_X1 U10699 ( .A1(n13257), .A2(n12922), .ZN(n8330) );
  NAND2_X1 U10700 ( .A1(n8331), .A2(n8330), .ZN(n13064) );
  NAND2_X1 U10701 ( .A1(n13064), .A2(n13058), .ZN(n8333) );
  NAND2_X1 U10702 ( .A1(n13066), .A2(n12921), .ZN(n8332) );
  NAND2_X1 U10703 ( .A1(n8333), .A2(n8332), .ZN(n13046) );
  NAND2_X1 U10704 ( .A1(n13319), .A2(n12890), .ZN(n8334) );
  NAND2_X1 U10705 ( .A1(n13238), .A2(n12919), .ZN(n8335) );
  INV_X1 U10706 ( .A(n13021), .ZN(n8337) );
  NAND2_X1 U10707 ( .A1(n8337), .A2(n8336), .ZN(n13231) );
  OR2_X1 U10708 ( .A1(n13019), .A2(n12892), .ZN(n8338) );
  NAND2_X1 U10709 ( .A1(n13231), .A2(n8338), .ZN(n13002) );
  NAND2_X1 U10710 ( .A1(n13002), .A2(n13003), .ZN(n13001) );
  NAND2_X1 U10711 ( .A1(n13229), .A2(n12917), .ZN(n8339) );
  NAND2_X1 U10712 ( .A1(n13001), .A2(n8339), .ZN(n8341) );
  INV_X1 U10713 ( .A(n12096), .ZN(n8340) );
  NAND2_X1 U10714 ( .A1(n13195), .A2(n12058), .ZN(n11845) );
  NOR2_X1 U10715 ( .A1(n11845), .A2(n8342), .ZN(n14918) );
  INV_X1 U10716 ( .A(n14918), .ZN(n9916) );
  NAND2_X1 U10717 ( .A1(n11839), .A2(n14905), .ZN(n8346) );
  INV_X1 U10718 ( .A(n11884), .ZN(n10611) );
  NAND2_X1 U10719 ( .A1(n10606), .A2(n10611), .ZN(n10607) );
  NOR2_X1 U10720 ( .A1(n10575), .A2(n11895), .ZN(n10845) );
  INV_X1 U10721 ( .A(n11905), .ZN(n10939) );
  INV_X1 U10722 ( .A(n11910), .ZN(n14916) );
  NAND2_X1 U10723 ( .A1(n10968), .A2(n14916), .ZN(n11108) );
  OR2_X2 U10724 ( .A1(n11108), .A2(n11919), .ZN(n11168) );
  OR2_X2 U10725 ( .A1(n13190), .A2(n13294), .ZN(n13191) );
  INV_X1 U10726 ( .A(n13283), .ZN(n13157) );
  OR2_X2 U10727 ( .A1(n13257), .A2(n13095), .ZN(n13080) );
  AND2_X2 U10728 ( .A1(n13319), .A2(n13065), .ZN(n13051) );
  INV_X1 U10729 ( .A(n6684), .ZN(n8344) );
  AND2_X4 U10730 ( .A1(n14883), .A2(n12066), .ZN(n14313) );
  AOI21_X1 U10731 ( .B1(n12022), .B2(n8344), .A(n11181), .ZN(n8345) );
  NAND2_X1 U10732 ( .A1(n12995), .A2(n8345), .ZN(n11837) );
  NOR4_X1 U10733 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n8350) );
  NOR4_X1 U10734 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n8349) );
  NOR4_X1 U10735 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n8348) );
  NOR4_X1 U10736 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n8347) );
  NAND4_X1 U10737 ( .A1(n8350), .A2(n8349), .A3(n8348), .A4(n8347), .ZN(n8366)
         );
  NOR2_X1 U10738 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .ZN(
        n8354) );
  NOR4_X1 U10739 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n8353) );
  NOR4_X1 U10740 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n8352) );
  NOR4_X1 U10741 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n8351) );
  NAND4_X1 U10742 ( .A1(n8354), .A2(n8353), .A3(n8352), .A4(n8351), .ZN(n8365)
         );
  NAND2_X1 U10743 ( .A1(n8355), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8356) );
  NAND2_X1 U10744 ( .A1(n6791), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8357) );
  MUX2_X1 U10745 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8357), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8358) );
  NAND2_X1 U10746 ( .A1(n8358), .A2(n8355), .ZN(n11461) );
  NAND2_X1 U10747 ( .A1(n8360), .A2(n8359), .ZN(n8371) );
  NAND2_X1 U10748 ( .A1(n8371), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8362) );
  XNOR2_X1 U10749 ( .A(n11335), .B(P2_B_REG_SCAN_IN), .ZN(n8363) );
  NAND2_X1 U10750 ( .A1(n11461), .A2(n8363), .ZN(n8364) );
  OAI21_X1 U10751 ( .B1(n8366), .B2(n8365), .A(n14849), .ZN(n9806) );
  INV_X1 U10752 ( .A(n11461), .ZN(n8367) );
  NAND2_X1 U10753 ( .A1(n8373), .A2(n8367), .ZN(n8368) );
  NAND2_X1 U10754 ( .A1(n8369), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8370) );
  MUX2_X1 U10755 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8370), .S(
        P2_IR_REG_23__SCAN_IN), .Z(n8372) );
  NAND2_X1 U10756 ( .A1(n8372), .A2(n8371), .ZN(n11309) );
  NAND2_X1 U10757 ( .A1(n9643), .A2(n11309), .ZN(n9930) );
  NAND2_X1 U10758 ( .A1(n12066), .A2(n12983), .ZN(n12056) );
  NAND2_X1 U10759 ( .A1(n9816), .A2(n12056), .ZN(n9809) );
  NAND3_X1 U10760 ( .A1(n9806), .A2(n14881), .A3(n9809), .ZN(n10189) );
  INV_X1 U10761 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15552) );
  NAND2_X1 U10762 ( .A1(n14849), .A2(n15552), .ZN(n8375) );
  INV_X1 U10763 ( .A(n8373), .ZN(n13360) );
  NAND2_X1 U10764 ( .A1(n13360), .A2(n11461), .ZN(n8374) );
  NAND2_X1 U10765 ( .A1(n8375), .A2(n8374), .ZN(n14880) );
  INV_X1 U10766 ( .A(n14880), .ZN(n9805) );
  OR2_X1 U10767 ( .A1(n9813), .A2(n9805), .ZN(n8376) );
  INV_X1 U10768 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14878) );
  NAND2_X1 U10769 ( .A1(n14849), .A2(n14878), .ZN(n8378) );
  NAND2_X1 U10770 ( .A1(n11335), .A2(n13360), .ZN(n8377) );
  AND2_X1 U10771 ( .A1(n8378), .A2(n8377), .ZN(n10190) );
  OR2_X1 U10772 ( .A1(n14934), .A2(n8379), .ZN(n8380) );
  INV_X1 U10773 ( .A(n12056), .ZN(n12102) );
  INV_X1 U10774 ( .A(n14883), .ZN(n9812) );
  OR2_X1 U10775 ( .A1(n12102), .A2(n9812), .ZN(n14915) );
  INV_X1 U10776 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8381) );
  NAND2_X1 U10777 ( .A1(n8381), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8561) );
  INV_X1 U10778 ( .A(n8561), .ZN(n8382) );
  NAND2_X1 U10779 ( .A1(n8553), .A2(n8382), .ZN(n8384) );
  NAND2_X1 U10780 ( .A1(n6989), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8383) );
  NAND2_X1 U10781 ( .A1(n8384), .A2(n8383), .ZN(n8571) );
  NAND2_X1 U10782 ( .A1(n9600), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8386) );
  INV_X1 U10783 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9609) );
  NAND2_X1 U10784 ( .A1(n9609), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8385) );
  NAND2_X1 U10785 ( .A1(n9596), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8388) );
  NAND2_X1 U10786 ( .A1(n9607), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8387) );
  AND2_X1 U10787 ( .A1(n8388), .A2(n8387), .ZN(n8584) );
  NAND2_X1 U10788 ( .A1(n9599), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8390) );
  INV_X1 U10789 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9602) );
  NAND2_X1 U10790 ( .A1(n9602), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8389) );
  NAND2_X1 U10791 ( .A1(n8601), .A2(n8600), .ZN(n8391) );
  NAND2_X1 U10792 ( .A1(n8391), .A2(n8390), .ZN(n8613) );
  NAND2_X1 U10793 ( .A1(n9613), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8393) );
  NAND2_X1 U10794 ( .A1(n9614), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8392) );
  NAND2_X1 U10795 ( .A1(n9631), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8394) );
  NAND2_X1 U10796 ( .A1(n9630), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8395) );
  NAND2_X1 U10797 ( .A1(n9636), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8398) );
  NAND2_X1 U10798 ( .A1(n9635), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n8396) );
  INV_X1 U10799 ( .A(n8644), .ZN(n8397) );
  NAND2_X1 U10800 ( .A1(n9706), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8401) );
  NAND2_X1 U10801 ( .A1(n9705), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8400) );
  NAND2_X1 U10802 ( .A1(n9740), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8403) );
  NAND2_X1 U10803 ( .A1(n9743), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8402) );
  NAND2_X1 U10804 ( .A1(n8678), .A2(n8403), .ZN(n8693) );
  NAND2_X1 U10805 ( .A1(n9788), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8405) );
  NAND2_X1 U10806 ( .A1(n9792), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8404) );
  NAND2_X1 U10807 ( .A1(n9888), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8406) );
  XNOR2_X1 U10808 ( .A(n10043), .B(P1_DATAO_REG_12__SCAN_IN), .ZN(n8717) );
  INV_X1 U10809 ( .A(n8717), .ZN(n8407) );
  NAND2_X1 U10810 ( .A1(n8718), .A2(n8407), .ZN(n8409) );
  NAND2_X1 U10811 ( .A1(n10043), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8408) );
  NAND2_X1 U10812 ( .A1(n8736), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8413) );
  NAND2_X1 U10813 ( .A1(n8411), .A2(n8410), .ZN(n8412) );
  XNOR2_X1 U10814 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n8751) );
  INV_X1 U10815 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n8414) );
  NAND2_X1 U10816 ( .A1(n8414), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8415) );
  XNOR2_X1 U10817 ( .A(n10521), .B(P2_DATAO_REG_15__SCAN_IN), .ZN(n8767) );
  INV_X1 U10818 ( .A(n8767), .ZN(n8416) );
  XNOR2_X1 U10819 ( .A(n8418), .B(P1_DATAO_REG_16__SCAN_IN), .ZN(n8779) );
  INV_X1 U10820 ( .A(n8779), .ZN(n8417) );
  NAND2_X1 U10821 ( .A1(n8418), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8419) );
  XNOR2_X1 U10822 ( .A(n10524), .B(P2_DATAO_REG_17__SCAN_IN), .ZN(n8795) );
  INV_X1 U10823 ( .A(n8795), .ZN(n8421) );
  NAND2_X1 U10824 ( .A1(n15494), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8422) );
  XNOR2_X1 U10825 ( .A(n15387), .B(P2_DATAO_REG_18__SCAN_IN), .ZN(n8807) );
  INV_X1 U10826 ( .A(n8807), .ZN(n8424) );
  NAND2_X1 U10827 ( .A1(n10725), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8425) );
  XNOR2_X1 U10828 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .ZN(n8820) );
  INV_X1 U10829 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10923) );
  NAND2_X1 U10830 ( .A1(n10923), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8426) );
  XNOR2_X2 U10831 ( .A(n8427), .B(P1_DATAO_REG_20__SCAN_IN), .ZN(n8835) );
  NAND2_X1 U10832 ( .A1(n8427), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8428) );
  NAND2_X1 U10833 ( .A1(n11000), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8430) );
  INV_X1 U10834 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n10974) );
  NAND2_X1 U10835 ( .A1(n10974), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8429) );
  NAND2_X1 U10836 ( .A1(n8430), .A2(n8429), .ZN(n8845) );
  NAND2_X1 U10837 ( .A1(n11177), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8433) );
  INV_X1 U10838 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8431) );
  NAND2_X1 U10839 ( .A1(n8431), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8432) );
  NAND2_X1 U10840 ( .A1(n11311), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8435) );
  NAND2_X1 U10841 ( .A1(n11307), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8434) );
  INV_X1 U10842 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8436) );
  NAND2_X1 U10843 ( .A1(n8884), .A2(n8436), .ZN(n8439) );
  NOR2_X1 U10844 ( .A1(n11462), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8440) );
  NAND2_X1 U10845 ( .A1(n11462), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8441) );
  XNOR2_X1 U10846 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .ZN(n8906) );
  NAND2_X1 U10847 ( .A1(n13358), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8442) );
  AND2_X1 U10848 ( .A1(n13356), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8444) );
  NAND2_X1 U10849 ( .A1(n11831), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8445) );
  NOR2_X1 U10850 ( .A1(n13354), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8446) );
  NAND2_X1 U10851 ( .A1(n13354), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8447) );
  XNOR2_X1 U10852 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n11530) );
  XNOR2_X1 U10853 ( .A(n11532), .B(n11530), .ZN(n12782) );
  NOR2_X1 U10854 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_6__SCAN_IN), .ZN(
        n8450) );
  NOR2_X1 U10855 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n8449) );
  NOR2_X1 U10856 ( .A1(P3_IR_REG_7__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n8448) );
  NAND3_X1 U10857 ( .A1(n8719), .A2(n8617), .A3(n8453), .ZN(n8724) );
  NOR2_X1 U10858 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), 
        .ZN(n8460) );
  NOR2_X2 U10859 ( .A1(n8463), .A2(P3_IR_REG_28__SCAN_IN), .ZN(n8534) );
  INV_X1 U10860 ( .A(n8534), .ZN(n8531) );
  NAND2_X1 U10861 ( .A1(n8463), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8464) );
  NAND2_X2 U10862 ( .A1(n8531), .A2(n8465), .ZN(n11819) );
  NAND2_X1 U10863 ( .A1(n8466), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8468) );
  XNOR2_X2 U10864 ( .A(n8468), .B(n8467), .ZN(n8943) );
  NAND2_X4 U10865 ( .A1(n11819), .A2(n8943), .ZN(n9825) );
  NAND2_X2 U10866 ( .A1(n9825), .A2(n9042), .ZN(n8679) );
  NAND2_X1 U10867 ( .A1(n12782), .A2(n11549), .ZN(n8470) );
  INV_X1 U10868 ( .A(SI_29_), .ZN(n12786) );
  OR2_X1 U10869 ( .A1(n11550), .A2(n12786), .ZN(n8469) );
  NAND2_X1 U10870 ( .A1(n8470), .A2(n8469), .ZN(n8941) );
  INV_X1 U10871 ( .A(n8941), .ZN(n12494) );
  NAND2_X1 U10872 ( .A1(n8474), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8475) );
  NAND2_X1 U10873 ( .A1(n6735), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8476) );
  MUX2_X1 U10874 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8476), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8477) );
  NAND2_X1 U10875 ( .A1(n8477), .A2(n8474), .ZN(n11022) );
  NOR2_X1 U10876 ( .A1(n11022), .A2(n10959), .ZN(n8480) );
  XNOR2_X1 U10877 ( .A(n10959), .B(P3_B_REG_SCAN_IN), .ZN(n8481) );
  NAND2_X1 U10878 ( .A1(n8481), .A2(n11022), .ZN(n8482) );
  NOR2_X1 U10879 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .ZN(
        n8486) );
  NOR4_X1 U10880 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_2__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8485) );
  NOR4_X1 U10881 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n8484) );
  NOR4_X1 U10882 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_25__SCAN_IN), .A3(
        P3_D_REG_22__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n8483) );
  NAND4_X1 U10883 ( .A1(n8486), .A2(n8485), .A3(n8484), .A4(n8483), .ZN(n8492)
         );
  NOR4_X1 U10884 ( .A1(P3_D_REG_14__SCAN_IN), .A2(P3_D_REG_12__SCAN_IN), .A3(
        P3_D_REG_11__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n8490) );
  NOR4_X1 U10885 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_31__SCAN_IN), .ZN(n8489) );
  NOR4_X1 U10886 ( .A1(P3_D_REG_23__SCAN_IN), .A2(P3_D_REG_6__SCAN_IN), .A3(
        P3_D_REG_3__SCAN_IN), .A4(P3_D_REG_5__SCAN_IN), .ZN(n8488) );
  NOR4_X1 U10887 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_30__SCAN_IN), .A4(P3_D_REG_13__SCAN_IN), .ZN(n8487) );
  NAND4_X1 U10888 ( .A1(n8490), .A2(n8489), .A3(n8488), .A4(n8487), .ZN(n8491)
         );
  NOR2_X1 U10889 ( .A1(n8492), .A2(n8491), .ZN(n8493) );
  NOR2_X1 U10890 ( .A1(n11755), .A2(n9936), .ZN(n9577) );
  INV_X1 U10891 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n8495) );
  NAND2_X1 U10892 ( .A1(n9709), .A2(n8495), .ZN(n8498) );
  INV_X1 U10893 ( .A(n8496), .ZN(n11138) );
  NAND2_X1 U10894 ( .A1(n11138), .A2(n11022), .ZN(n8497) );
  NAND2_X1 U10895 ( .A1(n11138), .A2(n10959), .ZN(n8499) );
  NAND2_X1 U10896 ( .A1(n10279), .A2(n12774), .ZN(n9937) );
  INV_X1 U10897 ( .A(n10279), .ZN(n10277) );
  NAND2_X1 U10898 ( .A1(n10277), .A2(n7260), .ZN(n9581) );
  AND3_X1 U10899 ( .A1(n9577), .A2(n9937), .A3(n9581), .ZN(n10283) );
  NAND2_X1 U10900 ( .A1(n8501), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8502) );
  MUX2_X1 U10901 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8502), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n8504) );
  AND2_X4 U10902 ( .A1(n11756), .A2(n11566), .ZN(n11711) );
  NAND2_X1 U10903 ( .A1(n8506), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8508) );
  NAND2_X1 U10904 ( .A1(n8509), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8510) );
  NAND2_X1 U10905 ( .A1(n10326), .A2(n9966), .ZN(n11716) );
  NAND2_X1 U10906 ( .A1(n11711), .A2(n11716), .ZN(n9941) );
  AND2_X1 U10907 ( .A1(n11716), .A2(n9966), .ZN(n8511) );
  NAND2_X1 U10908 ( .A1(n11756), .A2(n8511), .ZN(n8973) );
  NAND2_X1 U10909 ( .A1(n11697), .A2(n8973), .ZN(n10278) );
  NAND2_X1 U10910 ( .A1(n9941), .A2(n10278), .ZN(n10276) );
  NAND2_X1 U10911 ( .A1(n11756), .A2(n12483), .ZN(n9579) );
  NAND2_X1 U10912 ( .A1(n9579), .A2(n11716), .ZN(n8512) );
  NAND2_X1 U10913 ( .A1(n11559), .A2(n10326), .ZN(n8969) );
  AOI22_X1 U10914 ( .A1(n8512), .A2(n11559), .B1(n8975), .B2(n8969), .ZN(n8513) );
  MUX2_X1 U10915 ( .A(n10276), .B(n8513), .S(n10277), .Z(n8514) );
  INV_X1 U10916 ( .A(n12721), .ZN(n8517) );
  INV_X1 U10917 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n8938) );
  NOR2_X1 U10918 ( .A1(n15202), .A2(n8938), .ZN(n8516) );
  NOR2_X1 U10919 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8605) );
  NAND2_X1 U10920 ( .A1(n8605), .A2(n15315), .ZN(n8623) );
  INV_X1 U10921 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n8518) );
  NAND2_X1 U10922 ( .A1(n8740), .A2(n8518), .ZN(n8760) );
  NOR2_X1 U10923 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(P3_REG3_REG_18__SCAN_IN), 
        .ZN(n8521) );
  INV_X1 U10924 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n15304) );
  INV_X1 U10925 ( .A(n8901), .ZN(n8527) );
  INV_X1 U10926 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n8526) );
  INV_X1 U10927 ( .A(n8924), .ZN(n8529) );
  INV_X1 U10928 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n8528) );
  NAND2_X1 U10929 ( .A1(n8529), .A2(n8528), .ZN(n8926) );
  NAND2_X1 U10930 ( .A1(n8926), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8530) );
  NAND2_X1 U10931 ( .A1(n12487), .A2(n8530), .ZN(n12509) );
  NAND2_X1 U10932 ( .A1(n8531), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8532) );
  MUX2_X1 U10933 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8532), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n8535) );
  INV_X1 U10934 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8533) );
  INV_X1 U10935 ( .A(n8536), .ZN(n12777) );
  INV_X1 U10936 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n12669) );
  NAND2_X1 U10937 ( .A1(n8654), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8540) );
  NAND2_X1 U10938 ( .A1(n11541), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8539) );
  OAI211_X1 U10939 ( .C1(n12669), .C2(n8949), .A(n8540), .B(n8539), .ZN(n8541)
         );
  AOI21_X1 U10940 ( .B1(n12509), .B2(n8934), .A(n8541), .ZN(n12231) );
  XNOR2_X1 U10941 ( .A(n13354), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n8542) );
  XNOR2_X1 U10942 ( .A(n8543), .B(n8542), .ZN(n11817) );
  NAND2_X1 U10943 ( .A1(n11817), .A2(n11549), .ZN(n8545) );
  OR2_X1 U10944 ( .A1(n11550), .A2(n11818), .ZN(n8544) );
  NAND2_X1 U10945 ( .A1(n8927), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8549) );
  NAND2_X1 U10946 ( .A1(n8578), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n8548) );
  NAND2_X1 U10947 ( .A1(n8565), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n8547) );
  NAND2_X1 U10948 ( .A1(n8579), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n8546) );
  INV_X1 U10949 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n8550) );
  INV_X1 U10950 ( .A(n8572), .ZN(n8552) );
  OR2_X1 U10951 ( .A1(n8611), .A2(n6891), .ZN(n8555) );
  XNOR2_X1 U10952 ( .A(n8553), .B(n8561), .ZN(n9591) );
  INV_X1 U10953 ( .A(n10028), .ZN(n8564) );
  NAND2_X1 U10954 ( .A1(n8578), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8559) );
  NAND2_X1 U10955 ( .A1(n8927), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8558) );
  NAND2_X1 U10956 ( .A1(n8565), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8557) );
  NAND2_X1 U10957 ( .A1(n8579), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8556) );
  NAND4_X1 U10958 ( .A1(n8559), .A2(n8558), .A3(n8557), .A4(n8556), .ZN(n12411) );
  INV_X1 U10959 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9023) );
  NAND2_X1 U10960 ( .A1(n9023), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8560) );
  AND2_X1 U10961 ( .A1(n8561), .A2(n8560), .ZN(n8563) );
  OAI21_X1 U10962 ( .B1(n8205), .B2(n8563), .A(n8562), .ZN(n12788) );
  MUX2_X1 U10963 ( .A(P3_IR_REG_0__SCAN_IN), .B(n12788), .S(n9825), .Z(n10286)
         );
  NAND2_X1 U10964 ( .A1(n12411), .A2(n10286), .ZN(n15116) );
  NAND2_X1 U10965 ( .A1(n10586), .A2(n15112), .ZN(n10588) );
  NAND2_X1 U10966 ( .A1(n15114), .A2(n10588), .ZN(n8576) );
  NAND2_X1 U10967 ( .A1(n8927), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8569) );
  NAND2_X1 U10968 ( .A1(n8578), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8568) );
  NAND2_X1 U10969 ( .A1(n8565), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8567) );
  NAND2_X1 U10970 ( .A1(n8579), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n8566) );
  XNOR2_X1 U10971 ( .A(n8571), .B(n8570), .ZN(n9620) );
  OR2_X1 U10972 ( .A1(n8679), .A2(n9620), .ZN(n8575) );
  XNOR2_X2 U10973 ( .A(n8573), .B(P3_IR_REG_2__SCAN_IN), .ZN(n9967) );
  OR2_X1 U10974 ( .A1(n9825), .A2(n9967), .ZN(n8574) );
  NAND2_X1 U10975 ( .A1(n15118), .A2(n10083), .ZN(n11568) );
  NAND2_X1 U10976 ( .A1(n11568), .A2(n11573), .ZN(n8956) );
  NAND2_X1 U10977 ( .A1(n8927), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8583) );
  INV_X1 U10978 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n8577) );
  NAND2_X1 U10979 ( .A1(n8578), .A2(n8577), .ZN(n8582) );
  NAND2_X1 U10980 ( .A1(n8565), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8581) );
  NAND2_X1 U10981 ( .A1(n8579), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n8580) );
  OR2_X1 U10982 ( .A1(n8611), .A2(SI_3_), .ZN(n8591) );
  OR2_X1 U10983 ( .A1(n8585), .A2(n8584), .ZN(n8586) );
  NAND2_X1 U10984 ( .A1(n8587), .A2(n8586), .ZN(n9624) );
  OR2_X1 U10985 ( .A1(n8679), .A2(n9624), .ZN(n8590) );
  NAND2_X1 U10986 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n6693), .ZN(n8588) );
  OR2_X1 U10987 ( .A1(n9825), .A2(n14956), .ZN(n8589) );
  NAND2_X1 U10988 ( .A1(n10587), .A2(n12258), .ZN(n11575) );
  INV_X1 U10989 ( .A(n12258), .ZN(n11578) );
  NAND2_X1 U10990 ( .A1(n11575), .A2(n11572), .ZN(n10384) );
  NAND2_X1 U10991 ( .A1(n15118), .A2(n10593), .ZN(n10385) );
  AND2_X1 U10992 ( .A1(n10384), .A2(n10385), .ZN(n8592) );
  NAND2_X1 U10993 ( .A1(n12407), .A2(n12258), .ZN(n8593) );
  NAND2_X1 U10994 ( .A1(n8828), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8597) );
  OR2_X1 U10995 ( .A1(n7691), .A2(n8605), .ZN(n10513) );
  NAND2_X1 U10996 ( .A1(n8578), .A2(n10513), .ZN(n8596) );
  NAND2_X1 U10997 ( .A1(n8670), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8595) );
  OR2_X1 U10998 ( .A1(n8617), .A2(n8598), .ZN(n8599) );
  XNOR2_X1 U10999 ( .A(n8601), .B(n8600), .ZN(n9616) );
  OR2_X1 U11000 ( .A1(n8679), .A2(n9616), .ZN(n8603) );
  OR2_X1 U11001 ( .A1(n11550), .A2(SI_4_), .ZN(n8602) );
  OAI211_X1 U11002 ( .C1(n10795), .C2(n9825), .A(n8603), .B(n8602), .ZN(n15147) );
  INV_X1 U11003 ( .A(n15147), .ZN(n10514) );
  NAND2_X1 U11004 ( .A1(n12406), .A2(n10514), .ZN(n8604) );
  NAND2_X1 U11005 ( .A1(n8828), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8610) );
  OR2_X1 U11006 ( .A1(n15315), .A2(n8605), .ZN(n8606) );
  NAND2_X1 U11007 ( .A1(n8623), .A2(n8606), .ZN(n10627) );
  NAND2_X1 U11008 ( .A1(n8578), .A2(n10627), .ZN(n8609) );
  NAND2_X1 U11009 ( .A1(n8670), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8608) );
  NAND2_X1 U11010 ( .A1(n8579), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8607) );
  OR2_X1 U11011 ( .A1(n11550), .A2(SI_5_), .ZN(n8621) );
  OR2_X1 U11012 ( .A1(n8613), .A2(n8612), .ZN(n8614) );
  NAND2_X1 U11013 ( .A1(n8615), .A2(n8614), .ZN(n9626) );
  OR2_X1 U11014 ( .A1(n8679), .A2(n9626), .ZN(n8620) );
  NAND2_X1 U11015 ( .A1(n8617), .A2(n8616), .ZN(n8629) );
  NAND2_X1 U11016 ( .A1(n8629), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8618) );
  OR2_X1 U11017 ( .A1(n9825), .A2(n14962), .ZN(n8619) );
  NAND2_X1 U11018 ( .A1(n10742), .A2(n10559), .ZN(n11586) );
  INV_X1 U11019 ( .A(n10559), .ZN(n10626) );
  NAND2_X1 U11020 ( .A1(n12405), .A2(n10626), .ZN(n11585) );
  NAND2_X1 U11021 ( .A1(n8828), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8628) );
  NAND2_X1 U11022 ( .A1(n8623), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8624) );
  NAND2_X1 U11023 ( .A1(n8638), .A2(n8624), .ZN(n10747) );
  NAND2_X1 U11024 ( .A1(n8934), .A2(n10747), .ZN(n8627) );
  NAND2_X1 U11025 ( .A1(n6640), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8626) );
  NAND2_X1 U11026 ( .A1(n11541), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8625) );
  AND4_X2 U11027 ( .A1(n8628), .A2(n8627), .A3(n8626), .A4(n8625), .ZN(n10785)
         );
  NAND2_X1 U11028 ( .A1(n8721), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8630) );
  XNOR2_X1 U11029 ( .A(n8630), .B(P3_IR_REG_6__SCAN_IN), .ZN(n14982) );
  INV_X1 U11030 ( .A(SI_6_), .ZN(n9597) );
  OR2_X1 U11031 ( .A1(n11550), .A2(n9597), .ZN(n8634) );
  XNOR2_X1 U11032 ( .A(n9630), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n8631) );
  XNOR2_X1 U11033 ( .A(n8632), .B(n8631), .ZN(n9598) );
  OR2_X1 U11034 ( .A1(n8679), .A2(n9598), .ZN(n8633) );
  OAI211_X1 U11035 ( .C1(n9825), .C2(n10812), .A(n8634), .B(n8633), .ZN(n15156) );
  INV_X1 U11036 ( .A(n15156), .ZN(n8635) );
  NAND2_X1 U11037 ( .A1(n12404), .A2(n8635), .ZN(n11590) );
  NAND2_X1 U11038 ( .A1(n11589), .A2(n11590), .ZN(n8958) );
  NAND2_X1 U11039 ( .A1(n10742), .A2(n10626), .ZN(n10705) );
  AND2_X1 U11040 ( .A1(n8958), .A2(n10705), .ZN(n8636) );
  NAND2_X1 U11041 ( .A1(n10706), .A2(n8636), .ZN(n10704) );
  NAND2_X1 U11042 ( .A1(n12404), .A2(n15156), .ZN(n8637) );
  NAND2_X1 U11043 ( .A1(n10704), .A2(n8637), .ZN(n10784) );
  AND2_X1 U11044 ( .A1(n8638), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8639) );
  OR2_X1 U11045 ( .A1(n8639), .A2(n8652), .ZN(n12185) );
  NAND2_X1 U11046 ( .A1(n8934), .A2(n12185), .ZN(n8643) );
  NAND2_X1 U11047 ( .A1(n8828), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8642) );
  NAND2_X1 U11048 ( .A1(n8654), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8641) );
  NAND2_X1 U11049 ( .A1(n11541), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n8640) );
  XNOR2_X1 U11050 ( .A(n8645), .B(n8644), .ZN(n9622) );
  OR2_X1 U11051 ( .A1(n8679), .A2(n9622), .ZN(n8649) );
  OR2_X1 U11052 ( .A1(n11550), .A2(SI_7_), .ZN(n8648) );
  OR2_X1 U11053 ( .A1(n8660), .A2(n8598), .ZN(n8646) );
  OR2_X1 U11054 ( .A1(n9825), .A2(n14993), .ZN(n8647) );
  NAND2_X1 U11055 ( .A1(n10948), .A2(n12184), .ZN(n11594) );
  INV_X1 U11056 ( .A(n12184), .ZN(n10791) );
  NAND2_X1 U11057 ( .A1(n12403), .A2(n10791), .ZN(n11595) );
  NAND2_X1 U11058 ( .A1(n11594), .A2(n11595), .ZN(n11142) );
  NAND2_X1 U11059 ( .A1(n10784), .A2(n11142), .ZN(n8651) );
  NAND2_X1 U11060 ( .A1(n12403), .A2(n12184), .ZN(n8650) );
  NOR2_X1 U11061 ( .A1(n8652), .A2(n12286), .ZN(n8653) );
  OR2_X1 U11062 ( .A1(n8668), .A2(n8653), .ZN(n12290) );
  NAND2_X1 U11063 ( .A1(n8934), .A2(n12290), .ZN(n8658) );
  NAND2_X1 U11064 ( .A1(n8828), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8657) );
  NAND2_X1 U11065 ( .A1(n8654), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8656) );
  NAND2_X1 U11066 ( .A1(n11541), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8655) );
  NAND2_X1 U11067 ( .A1(n8660), .A2(n8659), .ZN(n8680) );
  NAND2_X1 U11068 ( .A1(n8680), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8661) );
  OR2_X1 U11069 ( .A1(n8663), .A2(n8662), .ZN(n8664) );
  NAND2_X1 U11070 ( .A1(n8665), .A2(n8664), .ZN(n9593) );
  OR2_X1 U11071 ( .A1(n8679), .A2(n9593), .ZN(n8667) );
  INV_X1 U11072 ( .A(SI_8_), .ZN(n9592) );
  OR2_X1 U11073 ( .A1(n11550), .A2(n9592), .ZN(n8666) );
  OAI211_X1 U11074 ( .C1(n9825), .C2(n10808), .A(n8667), .B(n8666), .ZN(n11145) );
  NAND2_X1 U11075 ( .A1(n11146), .A2(n11145), .ZN(n11598) );
  INV_X1 U11076 ( .A(n11145), .ZN(n12287) );
  NAND2_X1 U11077 ( .A1(n12402), .A2(n12287), .ZN(n11599) );
  NAND2_X1 U11078 ( .A1(n8828), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8674) );
  OR2_X1 U11079 ( .A1(n8668), .A2(n11152), .ZN(n8669) );
  NAND2_X1 U11080 ( .A1(n8686), .A2(n8669), .ZN(n11155) );
  NAND2_X1 U11081 ( .A1(n8934), .A2(n11155), .ZN(n8673) );
  NAND2_X1 U11082 ( .A1(n8654), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8672) );
  NAND2_X1 U11083 ( .A1(n11541), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8671) );
  OR2_X1 U11084 ( .A1(n8676), .A2(n8675), .ZN(n8677) );
  AND2_X1 U11085 ( .A1(n8678), .A2(n8677), .ZN(n9618) );
  OR2_X1 U11086 ( .A1(n8679), .A2(n9618), .ZN(n8684) );
  OR2_X1 U11087 ( .A1(n11550), .A2(SI_9_), .ZN(n8683) );
  NAND2_X1 U11088 ( .A1(n8696), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8681) );
  XNOR2_X1 U11089 ( .A(n8681), .B(P3_IR_REG_9__SCAN_IN), .ZN(n12460) );
  OR2_X1 U11090 ( .A1(n9825), .A2(n12460), .ZN(n8682) );
  NAND2_X1 U11091 ( .A1(n11336), .A2(n11139), .ZN(n11603) );
  INV_X1 U11092 ( .A(n11139), .ZN(n11153) );
  NAND2_X1 U11093 ( .A1(n12401), .A2(n11153), .ZN(n11604) );
  NAND2_X1 U11094 ( .A1(n11603), .A2(n11604), .ZN(n11728) );
  NAND2_X1 U11095 ( .A1(n11146), .A2(n12287), .ZN(n10925) );
  AND2_X1 U11096 ( .A1(n11728), .A2(n10925), .ZN(n8685) );
  NAND2_X1 U11097 ( .A1(n8828), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8691) );
  NAND2_X1 U11098 ( .A1(n8686), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8687) );
  NAND2_X1 U11099 ( .A1(n8703), .A2(n8687), .ZN(n12247) );
  NAND2_X1 U11100 ( .A1(n8934), .A2(n12247), .ZN(n8690) );
  NAND2_X1 U11101 ( .A1(n8654), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8689) );
  NAND2_X1 U11102 ( .A1(n11541), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8688) );
  OR2_X1 U11103 ( .A1(n8693), .A2(n8692), .ZN(n8694) );
  NAND2_X1 U11104 ( .A1(n8695), .A2(n8694), .ZN(n9595) );
  NAND2_X1 U11105 ( .A1(n11549), .A2(n9595), .ZN(n8700) );
  NAND2_X1 U11106 ( .A1(n8711), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8698) );
  INV_X1 U11107 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8697) );
  OR2_X1 U11108 ( .A1(n9825), .A2(n12462), .ZN(n8699) );
  OAI211_X1 U11109 ( .C1(n8611), .C2(SI_10_), .A(n8700), .B(n8699), .ZN(n11609) );
  XNOR2_X1 U11110 ( .A(n12400), .B(n11609), .ZN(n11605) );
  NAND2_X1 U11111 ( .A1(n11027), .A2(n11605), .ZN(n8702) );
  INV_X1 U11112 ( .A(n11609), .ZN(n12251) );
  NAND2_X1 U11113 ( .A1(n12400), .A2(n12251), .ZN(n8701) );
  NAND2_X1 U11114 ( .A1(n8828), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8708) );
  NAND2_X1 U11115 ( .A1(n8703), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8704) );
  NAND2_X1 U11116 ( .A1(n8728), .A2(n8704), .ZN(n15590) );
  NAND2_X1 U11117 ( .A1(n8934), .A2(n15590), .ZN(n8707) );
  NAND2_X1 U11118 ( .A1(n8654), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8706) );
  NAND2_X1 U11119 ( .A1(n11541), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n8705) );
  XNOR2_X1 U11120 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n8709) );
  XNOR2_X1 U11121 ( .A(n8710), .B(n8709), .ZN(n9601) );
  NAND2_X1 U11122 ( .A1(n9601), .A2(n11549), .ZN(n8715) );
  OAI21_X1 U11123 ( .B1(n8711), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8713) );
  INV_X1 U11124 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8712) );
  XNOR2_X1 U11125 ( .A(n8713), .B(n8712), .ZN(n15041) );
  AOI22_X1 U11126 ( .A1(n8823), .A2(n15428), .B1(n8822), .B2(n15041), .ZN(
        n8714) );
  NAND2_X1 U11127 ( .A1(n12249), .A2(n14288), .ZN(n11615) );
  INV_X1 U11128 ( .A(n12249), .ZN(n12399) );
  NAND2_X1 U11129 ( .A1(n15594), .A2(n12399), .ZN(n11616) );
  NAND2_X1 U11130 ( .A1(n12249), .A2(n15594), .ZN(n8716) );
  XNOR2_X1 U11131 ( .A(n8718), .B(n8717), .ZN(n9628) );
  NAND2_X1 U11132 ( .A1(n9628), .A2(n11549), .ZN(n8727) );
  INV_X1 U11133 ( .A(n8719), .ZN(n8720) );
  OAI21_X1 U11134 ( .B1(n8721), .B2(n8720), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n8723) );
  MUX2_X1 U11135 ( .A(n8723), .B(P3_IR_REG_31__SCAN_IN), .S(n8722), .Z(n8725)
         );
  AOI22_X1 U11136 ( .A1(n8823), .A2(SI_12_), .B1(n8822), .B2(n12466), .ZN(
        n8726) );
  NAND2_X1 U11137 ( .A1(n8727), .A2(n8726), .ZN(n14274) );
  NOR2_X1 U11138 ( .A1(n8740), .A2(n7678), .ZN(n14269) );
  INV_X1 U11139 ( .A(n14269), .ZN(n8729) );
  NAND2_X1 U11140 ( .A1(n8934), .A2(n8729), .ZN(n8733) );
  NAND2_X1 U11141 ( .A1(n8828), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8732) );
  NAND2_X1 U11142 ( .A1(n8654), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8731) );
  NAND2_X1 U11143 ( .A1(n11541), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8730) );
  OR2_X1 U11144 ( .A1(n14274), .A2(n11430), .ZN(n11620) );
  NAND2_X1 U11145 ( .A1(n14274), .A2(n11430), .ZN(n11621) );
  INV_X1 U11146 ( .A(n11430), .ZN(n12398) );
  NAND2_X1 U11147 ( .A1(n14274), .A2(n12398), .ZN(n8735) );
  XNOR2_X1 U11148 ( .A(n8736), .B(n10091), .ZN(n9639) );
  NAND2_X1 U11149 ( .A1(n9639), .A2(n11549), .ZN(n8739) );
  XNOR2_X1 U11150 ( .A(n8737), .B(P3_IR_REG_13__SCAN_IN), .ZN(n15074) );
  AOI22_X1 U11151 ( .A1(n8823), .A2(SI_13_), .B1(n8822), .B2(n15074), .ZN(
        n8738) );
  NAND2_X1 U11152 ( .A1(n8739), .A2(n8738), .ZN(n11350) );
  NAND2_X1 U11153 ( .A1(n14255), .A2(n11350), .ZN(n8747) );
  INV_X1 U11154 ( .A(n8740), .ZN(n8741) );
  NAND2_X1 U11155 ( .A1(n8741), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8742) );
  AND2_X1 U11156 ( .A1(n8760), .A2(n8742), .ZN(n11348) );
  INV_X1 U11157 ( .A(n11348), .ZN(n14258) );
  NAND2_X1 U11158 ( .A1(n8934), .A2(n14258), .ZN(n8746) );
  NAND2_X1 U11159 ( .A1(n8828), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n8745) );
  NAND2_X1 U11160 ( .A1(n8654), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8744) );
  NAND2_X1 U11161 ( .A1(n11541), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n8743) );
  NAND2_X1 U11162 ( .A1(n8747), .A2(n11483), .ZN(n8750) );
  INV_X1 U11163 ( .A(n14255), .ZN(n8748) );
  INV_X1 U11164 ( .A(n11350), .ZN(n14261) );
  NAND2_X1 U11165 ( .A1(n8748), .A2(n14261), .ZN(n8749) );
  XNOR2_X1 U11166 ( .A(n8752), .B(n8751), .ZN(n9739) );
  NAND2_X1 U11167 ( .A1(n9739), .A2(n11549), .ZN(n8759) );
  INV_X1 U11168 ( .A(n8753), .ZN(n8755) );
  NAND2_X1 U11169 ( .A1(n8755), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8754) );
  MUX2_X1 U11170 ( .A(n8754), .B(P3_IR_REG_31__SCAN_IN), .S(n15342), .Z(n8757)
         );
  NOR2_X1 U11171 ( .A1(n8755), .A2(P3_IR_REG_14__SCAN_IN), .ZN(n8782) );
  INV_X1 U11172 ( .A(n8782), .ZN(n8756) );
  NAND2_X1 U11173 ( .A1(n8757), .A2(n8756), .ZN(n15100) );
  AOI22_X1 U11174 ( .A1(n8823), .A2(n9738), .B1(n8822), .B2(n15100), .ZN(n8758) );
  NAND2_X1 U11175 ( .A1(n8828), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8765) );
  NAND2_X1 U11176 ( .A1(n8760), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8761) );
  NAND2_X1 U11177 ( .A1(n8772), .A2(n8761), .ZN(n11454) );
  NAND2_X1 U11178 ( .A1(n8934), .A2(n11454), .ZN(n8764) );
  NAND2_X1 U11179 ( .A1(n6640), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8763) );
  NAND2_X1 U11180 ( .A1(n11541), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8762) );
  NAND2_X1 U11181 ( .A1(n11474), .A2(n11631), .ZN(n8766) );
  NAND2_X1 U11182 ( .A1(n11440), .A2(n8766), .ZN(n11371) );
  XNOR2_X1 U11183 ( .A(n8768), .B(n8767), .ZN(n9750) );
  NAND2_X1 U11184 ( .A1(n9750), .A2(n11549), .ZN(n8771) );
  OR2_X1 U11185 ( .A1(n8782), .A2(n8598), .ZN(n8769) );
  XNOR2_X1 U11186 ( .A(n8769), .B(P3_IR_REG_15__SCAN_IN), .ZN(n12473) );
  AOI22_X1 U11187 ( .A1(n8823), .A2(SI_15_), .B1(n8822), .B2(n12473), .ZN(
        n8770) );
  NAND2_X1 U11188 ( .A1(n8771), .A2(n8770), .ZN(n11499) );
  NAND2_X1 U11189 ( .A1(n8828), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n8777) );
  NAND2_X1 U11190 ( .A1(n8772), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8773) );
  NAND2_X1 U11191 ( .A1(n8788), .A2(n8773), .ZN(n11494) );
  NAND2_X1 U11192 ( .A1(n8934), .A2(n11494), .ZN(n8776) );
  NAND2_X1 U11193 ( .A1(n8654), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8775) );
  NAND2_X1 U11194 ( .A1(n11541), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n8774) );
  OR2_X1 U11195 ( .A1(n11499), .A2(n12192), .ZN(n11637) );
  NAND2_X1 U11196 ( .A1(n11499), .A2(n12192), .ZN(n11642) );
  NAND2_X1 U11197 ( .A1(n11637), .A2(n11642), .ZN(n11732) );
  INV_X1 U11198 ( .A(n12192), .ZN(n12396) );
  NAND2_X1 U11199 ( .A1(n11499), .A2(n12396), .ZN(n11506) );
  NAND2_X1 U11200 ( .A1(n11507), .A2(n11506), .ZN(n8794) );
  XNOR2_X1 U11201 ( .A(n8780), .B(n8779), .ZN(n9795) );
  NAND2_X1 U11202 ( .A1(n9795), .A2(n11549), .ZN(n8787) );
  NAND2_X1 U11203 ( .A1(n8782), .A2(n8781), .ZN(n8784) );
  NAND2_X1 U11204 ( .A1(n8784), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8783) );
  MUX2_X1 U11205 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8783), .S(
        P3_IR_REG_16__SCAN_IN), .Z(n8785) );
  NAND2_X1 U11206 ( .A1(n8785), .A2(n8797), .ZN(n14214) );
  INV_X1 U11207 ( .A(n14214), .ZN(n12447) );
  AOI22_X1 U11208 ( .A1(n8823), .A2(SI_16_), .B1(n8822), .B2(n12447), .ZN(
        n8786) );
  NAND2_X1 U11209 ( .A1(n8828), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n8793) );
  NAND2_X1 U11210 ( .A1(n8788), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8789) );
  NAND2_X1 U11211 ( .A1(n8813), .A2(n8789), .ZN(n12312) );
  NAND2_X1 U11212 ( .A1(n8934), .A2(n12312), .ZN(n8792) );
  NAND2_X1 U11213 ( .A1(n8654), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8791) );
  NAND2_X1 U11214 ( .A1(n11541), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n8790) );
  OR2_X1 U11215 ( .A1(n12317), .A2(n12326), .ZN(n11638) );
  NAND2_X1 U11216 ( .A1(n12317), .A2(n12326), .ZN(n11641) );
  NAND2_X1 U11217 ( .A1(n11638), .A2(n11641), .ZN(n8963) );
  NAND2_X1 U11218 ( .A1(n8794), .A2(n8963), .ZN(n11504) );
  INV_X1 U11219 ( .A(n12326), .ZN(n12395) );
  NAND2_X1 U11220 ( .A1(n12317), .A2(n12395), .ZN(n12646) );
  NAND2_X1 U11221 ( .A1(n11504), .A2(n12646), .ZN(n8805) );
  XNOR2_X1 U11222 ( .A(n8796), .B(n8795), .ZN(n9883) );
  NAND2_X1 U11223 ( .A1(n9883), .A2(n11549), .ZN(n8800) );
  NAND2_X1 U11224 ( .A1(n8797), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8798) );
  XNOR2_X1 U11225 ( .A(n8798), .B(P3_IR_REG_17__SCAN_IN), .ZN(n12478) );
  AOI22_X1 U11226 ( .A1(n8823), .A2(SI_17_), .B1(n8822), .B2(n12478), .ZN(
        n8799) );
  NAND2_X1 U11227 ( .A1(n8828), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8804) );
  XNOR2_X1 U11228 ( .A(n8813), .B(P3_REG3_REG_17__SCAN_IN), .ZN(n12654) );
  NAND2_X1 U11229 ( .A1(n8934), .A2(n12654), .ZN(n8803) );
  NAND2_X1 U11230 ( .A1(n6640), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8802) );
  NAND2_X1 U11231 ( .A1(n11541), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n8801) );
  OR2_X1 U11232 ( .A1(n12653), .A2(n12199), .ZN(n11655) );
  NAND2_X1 U11233 ( .A1(n12653), .A2(n12199), .ZN(n11650) );
  NAND2_X1 U11234 ( .A1(n11655), .A2(n11650), .ZN(n11651) );
  INV_X1 U11235 ( .A(n12199), .ZN(n12394) );
  NAND2_X1 U11236 ( .A1(n12653), .A2(n12394), .ZN(n8806) );
  XNOR2_X1 U11237 ( .A(n8808), .B(n8807), .ZN(n9913) );
  NAND2_X1 U11238 ( .A1(n9913), .A2(n11549), .ZN(n8812) );
  INV_X1 U11239 ( .A(n8471), .ZN(n8809) );
  NAND2_X1 U11240 ( .A1(n8809), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8810) );
  XNOR2_X1 U11241 ( .A(n8810), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12480) );
  AOI22_X1 U11242 ( .A1(n8823), .A2(SI_18_), .B1(n8822), .B2(n12480), .ZN(
        n8811) );
  NAND2_X1 U11243 ( .A1(n8828), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8818) );
  OAI21_X1 U11244 ( .B1(n8813), .B2(P3_REG3_REG_17__SCAN_IN), .A(
        P3_REG3_REG_18__SCAN_IN), .ZN(n8814) );
  NAND2_X1 U11245 ( .A1(n8814), .A2(n8826), .ZN(n12636) );
  NAND2_X1 U11246 ( .A1(n8934), .A2(n12636), .ZN(n8817) );
  NAND2_X1 U11247 ( .A1(n8654), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n8816) );
  NAND2_X1 U11248 ( .A1(n11541), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8815) );
  NAND2_X1 U11249 ( .A1(n12709), .A2(n12324), .ZN(n11653) );
  XNOR2_X1 U11250 ( .A(n8821), .B(n8820), .ZN(n9964) );
  NAND2_X1 U11251 ( .A1(n9964), .A2(n11549), .ZN(n8825) );
  AOI22_X1 U11252 ( .A1(n8823), .A2(n9965), .B1(n8822), .B2(n9966), .ZN(n8824)
         );
  NAND2_X1 U11253 ( .A1(n8826), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8827) );
  NAND2_X1 U11254 ( .A1(n8838), .A2(n8827), .ZN(n12622) );
  NAND2_X1 U11255 ( .A1(n12622), .A2(n8934), .ZN(n8833) );
  NAND2_X1 U11256 ( .A1(n8828), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n8832) );
  NAND2_X1 U11257 ( .A1(n8654), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8831) );
  NAND2_X1 U11258 ( .A1(n11541), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n8830) );
  NAND4_X1 U11259 ( .A1(n8833), .A2(n8832), .A3(n8831), .A4(n8830), .ZN(n12392) );
  NAND2_X1 U11260 ( .A1(n12759), .A2(n12392), .ZN(n8964) );
  NAND2_X1 U11261 ( .A1(n11660), .A2(n8964), .ZN(n12617) );
  INV_X1 U11262 ( .A(n12324), .ZN(n12393) );
  OR2_X1 U11263 ( .A1(n12709), .A2(n12393), .ZN(n12618) );
  AND2_X1 U11264 ( .A1(n12617), .A2(n12618), .ZN(n8834) );
  INV_X1 U11265 ( .A(n12392), .ZN(n12206) );
  OR2_X1 U11266 ( .A1(n12759), .A2(n12206), .ZN(n12605) );
  XNOR2_X1 U11267 ( .A(n8835), .B(n11827), .ZN(n10323) );
  NAND2_X1 U11268 ( .A1(n10323), .A2(n11549), .ZN(n8837) );
  OR2_X1 U11269 ( .A1(n8611), .A2(n10325), .ZN(n8836) );
  NAND2_X1 U11270 ( .A1(n8838), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8839) );
  NAND2_X1 U11271 ( .A1(n8849), .A2(n8839), .ZN(n12610) );
  NAND2_X1 U11272 ( .A1(n12610), .A2(n8934), .ZN(n8842) );
  AOI22_X1 U11273 ( .A1(n8828), .A2(P3_REG1_REG_20__SCAN_IN), .B1(n6640), .B2(
        P3_REG0_REG_20__SCAN_IN), .ZN(n8841) );
  NAND2_X1 U11274 ( .A1(n11541), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n8840) );
  NAND2_X1 U11275 ( .A1(n12343), .A2(n12210), .ZN(n11666) );
  NAND2_X1 U11276 ( .A1(n11665), .A2(n11666), .ZN(n12604) );
  NAND2_X1 U11277 ( .A1(n12343), .A2(n12391), .ZN(n8844) );
  XNOR2_X1 U11278 ( .A(n8846), .B(n8845), .ZN(n10432) );
  NAND2_X1 U11279 ( .A1(n10432), .A2(n11549), .ZN(n8848) );
  INV_X1 U11280 ( .A(SI_21_), .ZN(n10433) );
  OR2_X1 U11281 ( .A1(n11550), .A2(n10433), .ZN(n8847) );
  NAND2_X1 U11282 ( .A1(n8849), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8850) );
  NAND2_X1 U11283 ( .A1(n8861), .A2(n8850), .ZN(n12597) );
  NAND2_X1 U11284 ( .A1(n12597), .A2(n8934), .ZN(n8853) );
  AOI22_X1 U11285 ( .A1(n8828), .A2(P3_REG1_REG_21__SCAN_IN), .B1(n8654), .B2(
        P3_REG0_REG_21__SCAN_IN), .ZN(n8852) );
  NAND2_X1 U11286 ( .A1(n11541), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n8851) );
  NAND2_X1 U11287 ( .A1(n12596), .A2(n12354), .ZN(n11670) );
  INV_X1 U11288 ( .A(n12354), .ZN(n12390) );
  OR2_X1 U11289 ( .A1(n8855), .A2(n8854), .ZN(n8856) );
  NAND2_X1 U11290 ( .A1(n8857), .A2(n8856), .ZN(n10539) );
  NAND2_X1 U11291 ( .A1(n10539), .A2(n11549), .ZN(n8860) );
  OR2_X1 U11292 ( .A1(n11550), .A2(n8858), .ZN(n8859) );
  INV_X1 U11293 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n8865) );
  NAND2_X1 U11294 ( .A1(n8861), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8862) );
  NAND2_X1 U11295 ( .A1(n8873), .A2(n8862), .ZN(n12586) );
  NAND2_X1 U11296 ( .A1(n12586), .A2(n8934), .ZN(n8864) );
  AOI22_X1 U11297 ( .A1(n8828), .A2(P3_REG1_REG_22__SCAN_IN), .B1(n8654), .B2(
        P3_REG0_REG_22__SCAN_IN), .ZN(n8863) );
  OAI211_X1 U11298 ( .C1(n8594), .C2(n8865), .A(n8864), .B(n8863), .ZN(n12389)
         );
  NOR2_X1 U11299 ( .A1(n12361), .A2(n12389), .ZN(n8866) );
  INV_X1 U11300 ( .A(n12389), .ZN(n12568) );
  OR2_X1 U11301 ( .A1(n8868), .A2(n8867), .ZN(n8869) );
  NAND2_X1 U11302 ( .A1(n8870), .A2(n8869), .ZN(n10645) );
  NAND2_X1 U11303 ( .A1(n10645), .A2(n11549), .ZN(n8872) );
  OR2_X1 U11304 ( .A1(n8611), .A2(n10647), .ZN(n8871) );
  NAND2_X1 U11305 ( .A1(n8873), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8874) );
  NAND2_X1 U11306 ( .A1(n8887), .A2(n8874), .ZN(n12573) );
  NAND2_X1 U11307 ( .A1(n12573), .A2(n8934), .ZN(n8880) );
  INV_X1 U11308 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n8877) );
  NAND2_X1 U11309 ( .A1(n8828), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8876) );
  NAND2_X1 U11310 ( .A1(n8654), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8875) );
  OAI211_X1 U11311 ( .C1(n8877), .C2(n8594), .A(n8876), .B(n8875), .ZN(n8878)
         );
  INV_X1 U11312 ( .A(n8878), .ZN(n8879) );
  NAND2_X1 U11313 ( .A1(n12687), .A2(n12355), .ZN(n8881) );
  NAND2_X1 U11314 ( .A1(n11681), .A2(n8881), .ZN(n11675) );
  NAND2_X1 U11315 ( .A1(n12566), .A2(n11675), .ZN(n8883) );
  NAND2_X1 U11316 ( .A1(n12687), .A2(n12388), .ZN(n8882) );
  NAND2_X1 U11317 ( .A1(n8883), .A2(n8882), .ZN(n12553) );
  XNOR2_X1 U11318 ( .A(n8884), .B(P2_DATAO_REG_24__SCAN_IN), .ZN(n10956) );
  NAND2_X1 U11319 ( .A1(n10956), .A2(n11549), .ZN(n8886) );
  INV_X1 U11320 ( .A(SI_24_), .ZN(n10957) );
  OR2_X1 U11321 ( .A1(n11550), .A2(n10957), .ZN(n8885) );
  NAND2_X1 U11322 ( .A1(n8887), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8888) );
  NAND2_X1 U11323 ( .A1(n8901), .A2(n8888), .ZN(n12558) );
  NAND2_X1 U11324 ( .A1(n12558), .A2(n8934), .ZN(n8894) );
  INV_X1 U11325 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n8891) );
  NAND2_X1 U11326 ( .A1(n11541), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n8890) );
  NAND2_X1 U11327 ( .A1(n6640), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8889) );
  OAI211_X1 U11328 ( .C1(n8949), .C2(n8891), .A(n8890), .B(n8889), .ZN(n8892)
         );
  INV_X1 U11329 ( .A(n8892), .ZN(n8893) );
  AND2_X1 U11330 ( .A1(n12683), .A2(n12305), .ZN(n8895) );
  OR2_X1 U11331 ( .A1(n12683), .A2(n12305), .ZN(n8896) );
  XNOR2_X1 U11332 ( .A(n11462), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n8897) );
  XNOR2_X1 U11333 ( .A(n8898), .B(n8897), .ZN(n11020) );
  NAND2_X1 U11334 ( .A1(n11020), .A2(n11549), .ZN(n8900) );
  INV_X1 U11335 ( .A(SI_25_), .ZN(n11021) );
  OR2_X1 U11336 ( .A1(n11550), .A2(n11021), .ZN(n8899) );
  NAND2_X1 U11337 ( .A1(n8901), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8902) );
  NAND2_X1 U11338 ( .A1(n8910), .A2(n8902), .ZN(n12548) );
  INV_X1 U11339 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n12681) );
  NAND2_X1 U11340 ( .A1(n11541), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8904) );
  NAND2_X1 U11341 ( .A1(n6640), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8903) );
  OAI211_X1 U11342 ( .C1(n8949), .C2(n12681), .A(n8904), .B(n8903), .ZN(n8905)
         );
  AOI21_X1 U11343 ( .B1(n12548), .B2(n8934), .A(n8905), .ZN(n12227) );
  NAND2_X1 U11344 ( .A1(n12547), .A2(n12227), .ZN(n11692) );
  INV_X1 U11345 ( .A(n12227), .ZN(n12373) );
  XNOR2_X1 U11346 ( .A(n8907), .B(n8906), .ZN(n11135) );
  NAND2_X1 U11347 ( .A1(n11135), .A2(n11549), .ZN(n8909) );
  OR2_X1 U11348 ( .A1(n11550), .A2(n11136), .ZN(n8908) );
  NAND2_X1 U11349 ( .A1(n8910), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8911) );
  NAND2_X1 U11350 ( .A1(n8924), .A2(n8911), .ZN(n12531) );
  NAND2_X1 U11351 ( .A1(n12531), .A2(n8934), .ZN(n8917) );
  INV_X1 U11352 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n8914) );
  NAND2_X1 U11353 ( .A1(n11541), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8913) );
  NAND2_X1 U11354 ( .A1(n8654), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8912) );
  OAI211_X1 U11355 ( .C1(n8949), .C2(n8914), .A(n8913), .B(n8912), .ZN(n8915)
         );
  INV_X1 U11356 ( .A(n8915), .ZN(n8916) );
  OR2_X1 U11357 ( .A1(n12675), .A2(n12387), .ZN(n8919) );
  AND2_X1 U11358 ( .A1(n12675), .A2(n12387), .ZN(n8918) );
  XNOR2_X1 U11359 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n8920) );
  NAND2_X1 U11360 ( .A1(n11178), .A2(n11549), .ZN(n8923) );
  OR2_X1 U11361 ( .A1(n11550), .A2(n11179), .ZN(n8922) );
  NAND2_X1 U11362 ( .A1(n8924), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8925) );
  NAND2_X1 U11363 ( .A1(n8926), .A2(n8925), .ZN(n12525) );
  NAND2_X1 U11364 ( .A1(n12525), .A2(n8934), .ZN(n8932) );
  INV_X1 U11365 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n15398) );
  NAND2_X1 U11366 ( .A1(n8828), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8929) );
  NAND2_X1 U11367 ( .A1(n6640), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8928) );
  OAI211_X1 U11368 ( .C1(n15398), .C2(n8594), .A(n8929), .B(n8928), .ZN(n8930)
         );
  INV_X1 U11369 ( .A(n8930), .ZN(n8931) );
  OR2_X1 U11370 ( .A1(n12670), .A2(n12386), .ZN(n8933) );
  NAND2_X1 U11371 ( .A1(n12513), .A2(n12231), .ZN(n11702) );
  NAND2_X1 U11372 ( .A1(n11700), .A2(n11702), .ZN(n12500) );
  OAI21_X1 U11373 ( .B1(n12231), .B2(n12732), .A(n12499), .ZN(n8942) );
  INV_X1 U11374 ( .A(n12487), .ZN(n8935) );
  NAND2_X1 U11375 ( .A1(n8935), .A2(n8934), .ZN(n11546) );
  NAND2_X1 U11376 ( .A1(n8654), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8937) );
  NAND2_X1 U11377 ( .A1(n11541), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8936) );
  OAI211_X1 U11378 ( .C1(n8938), .C2(n8949), .A(n8937), .B(n8936), .ZN(n8939)
         );
  INV_X1 U11379 ( .A(n8939), .ZN(n8940) );
  OR2_X1 U11380 ( .A1(n8941), .A2(n12503), .ZN(n11707) );
  NAND2_X1 U11381 ( .A1(n8941), .A2(n12503), .ZN(n11708) );
  NAND2_X1 U11382 ( .A1(n11707), .A2(n11708), .ZN(n11743) );
  XNOR2_X1 U11383 ( .A(n8942), .B(n11743), .ZN(n8955) );
  INV_X1 U11384 ( .A(n10326), .ZN(n9578) );
  NAND2_X1 U11385 ( .A1(n11566), .A2(n9578), .ZN(n11558) );
  INV_X1 U11386 ( .A(P3_B_REG_SCAN_IN), .ZN(n8945) );
  INV_X1 U11387 ( .A(n11819), .ZN(n9826) );
  NAND2_X1 U11388 ( .A1(n9826), .A2(n11753), .ZN(n9833) );
  NAND2_X1 U11389 ( .A1(n9833), .A2(n9825), .ZN(n8944) );
  OAI21_X1 U11390 ( .B1(n11819), .B2(n8945), .A(n12375), .ZN(n12485) );
  INV_X1 U11391 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n8948) );
  NAND2_X1 U11392 ( .A1(n11541), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n8947) );
  NAND2_X1 U11393 ( .A1(n6640), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8946) );
  OAI211_X1 U11394 ( .C1(n8949), .C2(n8948), .A(n8947), .B(n8946), .ZN(n8950)
         );
  INV_X1 U11395 ( .A(n8950), .ZN(n8951) );
  NOR2_X1 U11396 ( .A1(n12485), .A2(n11554), .ZN(n8953) );
  NAND3_X1 U11397 ( .A1(n9833), .A2(n11711), .A3(n9825), .ZN(n15119) );
  NOR2_X1 U11398 ( .A1(n12231), .A2(n15119), .ZN(n8952) );
  INV_X1 U11399 ( .A(n10286), .ZN(n10056) );
  NAND2_X1 U11400 ( .A1(n15113), .A2(n11567), .ZN(n10031) );
  NAND2_X1 U11401 ( .A1(n10031), .A2(n11570), .ZN(n10585) );
  INV_X1 U11402 ( .A(n8956), .ZN(n11719) );
  INV_X1 U11403 ( .A(n10384), .ZN(n11723) );
  INV_X1 U11404 ( .A(n11729), .ZN(n11580) );
  NAND2_X1 U11405 ( .A1(n10504), .A2(n11580), .ZN(n10506) );
  INV_X1 U11406 ( .A(n12406), .ZN(n10562) );
  NAND2_X1 U11407 ( .A1(n10562), .A2(n10514), .ZN(n11582) );
  NAND2_X1 U11408 ( .A1(n10506), .A2(n11582), .ZN(n10617) );
  NAND2_X1 U11409 ( .A1(n10617), .A2(n11721), .ZN(n8957) );
  NAND2_X1 U11410 ( .A1(n8957), .A2(n11586), .ZN(n10702) );
  NAND2_X1 U11411 ( .A1(n10702), .A2(n11725), .ZN(n10701) );
  INV_X1 U11412 ( .A(n11142), .ZN(n11718) );
  INV_X1 U11413 ( .A(n11598), .ZN(n8959) );
  NAND2_X1 U11414 ( .A1(n8960), .A2(n11603), .ZN(n11024) );
  NAND2_X1 U11415 ( .A1(n12400), .A2(n11609), .ZN(n8961) );
  INV_X1 U11416 ( .A(n14290), .ZN(n11612) );
  NAND2_X1 U11417 ( .A1(n14273), .A2(n14272), .ZN(n8962) );
  AND2_X1 U11418 ( .A1(n11350), .A2(n11483), .ZN(n11625) );
  OR2_X1 U11419 ( .A1(n11350), .A2(n11483), .ZN(n11627) );
  INV_X1 U11420 ( .A(n11631), .ZN(n12397) );
  OR2_X1 U11421 ( .A1(n11474), .A2(n12397), .ZN(n11630) );
  INV_X1 U11422 ( .A(n11732), .ZN(n11441) );
  NAND2_X1 U11423 ( .A1(n11502), .A2(n11641), .ZN(n12645) );
  INV_X1 U11424 ( .A(n8964), .ZN(n11662) );
  NAND2_X1 U11425 ( .A1(n12591), .A2(n11670), .ZN(n8965) );
  NAND2_X1 U11426 ( .A1(n8965), .A2(n11669), .ZN(n12580) );
  NAND2_X1 U11427 ( .A1(n12361), .A2(n12568), .ZN(n11674) );
  NAND2_X1 U11428 ( .A1(n12580), .A2(n11674), .ZN(n8966) );
  OR2_X1 U11429 ( .A1(n12361), .A2(n12568), .ZN(n11673) );
  OR2_X1 U11430 ( .A1(n12683), .A2(n12569), .ZN(n11680) );
  NAND2_X1 U11431 ( .A1(n12683), .A2(n12569), .ZN(n11685) );
  NAND2_X1 U11432 ( .A1(n11680), .A2(n11685), .ZN(n11717) );
  INV_X1 U11433 ( .A(n11692), .ZN(n8967) );
  NOR2_X1 U11434 ( .A1(n12675), .A2(n12228), .ZN(n11694) );
  NAND2_X1 U11435 ( .A1(n12675), .A2(n12228), .ZN(n11691) );
  INV_X1 U11436 ( .A(n12518), .ZN(n12523) );
  NAND2_X1 U11437 ( .A1(n12524), .A2(n12523), .ZN(n12522) );
  NAND2_X1 U11438 ( .A1(n12670), .A2(n12502), .ZN(n11701) );
  NAND2_X1 U11439 ( .A1(n12522), .A2(n11701), .ZN(n12508) );
  INV_X1 U11440 ( .A(n11702), .ZN(n8968) );
  XNOR2_X1 U11441 ( .A(n11756), .B(n8969), .ZN(n8971) );
  NAND2_X1 U11442 ( .A1(n11559), .A2(n9966), .ZN(n8970) );
  NAND2_X1 U11443 ( .A1(n8971), .A2(n8970), .ZN(n9951) );
  INV_X1 U11444 ( .A(n11716), .ZN(n9950) );
  AND2_X1 U11445 ( .A1(n15146), .A2(n9950), .ZN(n8972) );
  NAND2_X1 U11446 ( .A1(n9951), .A2(n8972), .ZN(n8974) );
  NAND2_X1 U11447 ( .A1(n8974), .A2(n8973), .ZN(n11379) );
  NAND2_X1 U11448 ( .A1(n14924), .A2(n14892), .ZN(n13329) );
  NOR2_X1 U11449 ( .A1(n14924), .A2(n8980), .ZN(n8981) );
  NOR2_X1 U11450 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), 
        .ZN(n8987) );
  NOR2_X2 U11451 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n9197) );
  NOR2_X2 U11452 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n9196) );
  NOR2_X2 U11453 ( .A1(n9281), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n9294) );
  INV_X2 U11454 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9307) );
  INV_X1 U11455 ( .A(n8999), .ZN(n9555) );
  NAND2_X1 U11456 ( .A1(n8996), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8992) );
  MUX2_X1 U11457 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8992), .S(
        P1_IR_REG_21__SCAN_IN), .Z(n8993) );
  NAND2_X1 U11458 ( .A1(n8994), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8995) );
  INV_X1 U11459 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n8998) );
  XNOR2_X2 U11460 ( .A(n9000), .B(P1_IR_REG_22__SCAN_IN), .ZN(n10298) );
  NAND2_X1 U11461 ( .A1(n9001), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9002) );
  XNOR2_X2 U11462 ( .A(n9002), .B(P1_IR_REG_19__SCAN_IN), .ZN(n10878) );
  NAND2_X1 U11463 ( .A1(n10309), .A2(n9003), .ZN(n9497) );
  NAND4_X1 U11464 ( .A1(n9307), .A2(n9005), .A3(n9006), .A4(n9004), .ZN(n9008)
         );
  NAND2_X1 U11465 ( .A1(n9082), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n9021) );
  INV_X1 U11466 ( .A(n9017), .ZN(n11829) );
  NAND2_X1 U11467 ( .A1(n9057), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9020) );
  NAND2_X1 U11468 ( .A1(n9058), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9019) );
  NAND2_X1 U11469 ( .A1(n9085), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n9018) );
  INV_X1 U11470 ( .A(SI_0_), .ZN(n9022) );
  NOR2_X1 U11471 ( .A1(n8205), .A2(n9022), .ZN(n9024) );
  XNOR2_X1 U11472 ( .A(n9024), .B(n9023), .ZN(n14045) );
  INV_X1 U11473 ( .A(n9026), .ZN(n9027) );
  MUX2_X1 U11474 ( .A(n14044), .B(n14045), .S(n9043), .Z(n10365) );
  NAND2_X1 U11475 ( .A1(n10351), .A2(n10365), .ZN(n10302) );
  NAND2_X1 U11476 ( .A1(n10302), .A2(n10299), .ZN(n9031) );
  INV_X1 U11477 ( .A(n10365), .ZN(n10918) );
  NAND2_X1 U11478 ( .A1(n10017), .A2(n10918), .ZN(n9539) );
  NAND2_X1 U11479 ( .A1(n9031), .A2(n9539), .ZN(n9032) );
  NAND2_X1 U11480 ( .A1(n9057), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9037) );
  NAND2_X1 U11481 ( .A1(n9085), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n9036) );
  NAND2_X1 U11482 ( .A1(n9058), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9035) );
  NAND2_X1 U11483 ( .A1(n9082), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n9034) );
  NAND2_X1 U11484 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n14044), .ZN(n9038) );
  MUX2_X1 U11485 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9038), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n9041) );
  INV_X1 U11486 ( .A(n9039), .ZN(n9040) );
  INV_X1 U11487 ( .A(n10128), .ZN(n13602) );
  NAND2_X1 U11488 ( .A1(n9310), .A2(n13602), .ZN(n9047) );
  NAND2_X2 U11489 ( .A1(n9043), .A2(n8205), .ZN(n9486) );
  INV_X1 U11490 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n9605) );
  OR2_X1 U11491 ( .A1(n9486), .A2(n9605), .ZN(n9046) );
  CLKBUF_X2 U11492 ( .A(n6672), .Z(n12178) );
  NAND2_X1 U11493 ( .A1(n10152), .A2(n12178), .ZN(n10295) );
  NAND2_X1 U11494 ( .A1(n9082), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n9051) );
  NAND2_X1 U11495 ( .A1(n9058), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9050) );
  NAND2_X1 U11496 ( .A1(n9085), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n9048) );
  OR2_X1 U11497 ( .A1(n9486), .A2(n9609), .ZN(n9054) );
  OR2_X1 U11498 ( .A1(n9039), .A2(n8998), .ZN(n9052) );
  XNOR2_X1 U11499 ( .A(n9052), .B(P1_IR_REG_2__SCAN_IN), .ZN(n13620) );
  NAND2_X1 U11500 ( .A1(n9310), .A2(n13620), .ZN(n9053) );
  NAND2_X1 U11501 ( .A1(n10144), .A2(n14574), .ZN(n10885) );
  INV_X1 U11502 ( .A(n10144), .ZN(n13598) );
  NAND2_X1 U11503 ( .A1(n13598), .A2(n10313), .ZN(n9055) );
  NAND2_X1 U11504 ( .A1(n10885), .A2(n9055), .ZN(n10862) );
  OAI211_X1 U11505 ( .C1(n9069), .C2(n10295), .A(n10862), .B(n9056), .ZN(n9072) );
  NAND2_X1 U11506 ( .A1(n10144), .A2(n10313), .ZN(n10864) );
  INV_X1 U11507 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n11087) );
  NAND2_X1 U11508 ( .A1(n9082), .A2(n11087), .ZN(n9062) );
  NAND2_X1 U11509 ( .A1(n9057), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9061) );
  NAND2_X1 U11510 ( .A1(n9085), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9059) );
  OR2_X1 U11511 ( .A1(n9486), .A2(n9607), .ZN(n9065) );
  NAND3_X1 U11512 ( .A1(n9499), .A2(n14574), .A3(n13598), .ZN(n9066) );
  OAI211_X1 U11513 ( .C1(n10864), .C2(n9499), .A(n11090), .B(n9066), .ZN(n9067) );
  INV_X1 U11514 ( .A(n9067), .ZN(n9071) );
  NAND3_X1 U11515 ( .A1(n9072), .A2(n9071), .A3(n9070), .ZN(n9076) );
  NAND2_X1 U11516 ( .A1(n9499), .A2(n11088), .ZN(n9074) );
  INV_X1 U11517 ( .A(n11088), .ZN(n14612) );
  NAND2_X1 U11518 ( .A1(n9108), .A2(n14612), .ZN(n9073) );
  MUX2_X1 U11519 ( .A(n9074), .B(n9073), .S(n13597), .Z(n9075) );
  NAND2_X1 U11520 ( .A1(n9076), .A2(n9075), .ZN(n9092) );
  OR2_X1 U11521 ( .A1(n9485), .A2(n9603), .ZN(n9081) );
  OR2_X1 U11522 ( .A1(n9486), .A2(n9602), .ZN(n9080) );
  OR2_X1 U11523 ( .A1(n9077), .A2(n8998), .ZN(n9078) );
  XNOR2_X1 U11524 ( .A(n9078), .B(P1_IR_REG_4__SCAN_IN), .ZN(n13645) );
  NAND2_X1 U11525 ( .A1(n6935), .A2(n13645), .ZN(n9079) );
  INV_X2 U11526 ( .A(n9343), .ZN(n9454) );
  INV_X1 U11527 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n9083) );
  NAND2_X1 U11528 ( .A1(n11087), .A2(n9083), .ZN(n9084) );
  NAND2_X1 U11529 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n9102) );
  AND2_X1 U11530 ( .A1(n9084), .A2(n9102), .ZN(n11068) );
  NAND2_X1 U11531 ( .A1(n9454), .A2(n11068), .ZN(n9089) );
  NAND2_X1 U11532 ( .A1(n9492), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9088) );
  NAND2_X1 U11533 ( .A1(n9466), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n9087) );
  INV_X2 U11534 ( .A(n9491), .ZN(n9493) );
  NAND2_X1 U11535 ( .A1(n9493), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9086) );
  MUX2_X1 U11536 ( .A(n10889), .B(n11092), .S(n9499), .Z(n9091) );
  MUX2_X1 U11537 ( .A(n10867), .B(n11072), .S(n9499), .Z(n9090) );
  OAI21_X1 U11538 ( .B1(n9092), .B2(n9091), .A(n9090), .ZN(n9094) );
  NAND2_X1 U11539 ( .A1(n9092), .A2(n9091), .ZN(n9093) );
  NAND2_X1 U11540 ( .A1(n9096), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9098) );
  INV_X1 U11541 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9097) );
  XNOR2_X1 U11542 ( .A(n9098), .B(n9097), .ZN(n10133) );
  OR2_X1 U11543 ( .A1(n9485), .A2(n9615), .ZN(n9100) );
  OR2_X1 U11544 ( .A1(n9486), .A2(n9614), .ZN(n9099) );
  OAI211_X1 U11545 ( .C1(n9043), .C2(n10133), .A(n9100), .B(n9099), .ZN(n10899) );
  NOR2_X1 U11546 ( .A1(n9102), .A2(n9101), .ZN(n9116) );
  AND2_X1 U11547 ( .A1(n9102), .A2(n9101), .ZN(n9103) );
  NOR2_X1 U11548 ( .A1(n9116), .A2(n9103), .ZN(n10881) );
  NAND2_X1 U11549 ( .A1(n9454), .A2(n10881), .ZN(n9107) );
  NAND2_X1 U11550 ( .A1(n9492), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n9106) );
  NAND2_X1 U11551 ( .A1(n9493), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9105) );
  NAND2_X1 U11552 ( .A1(n9466), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n9104) );
  NAND4_X1 U11553 ( .A1(n9107), .A2(n9106), .A3(n9105), .A4(n9104), .ZN(n13596) );
  MUX2_X1 U11554 ( .A(n10899), .B(n13596), .S(n9473), .Z(n9110) );
  MUX2_X1 U11555 ( .A(n13596), .B(n10899), .S(n9473), .Z(n9109) );
  NOR2_X1 U11556 ( .A1(n9096), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n9113) );
  OR2_X1 U11557 ( .A1(n9113), .A2(n8998), .ZN(n9111) );
  MUX2_X1 U11558 ( .A(n9111), .B(P1_IR_REG_31__SCAN_IN), .S(n9112), .Z(n9114)
         );
  NAND2_X1 U11559 ( .A1(n9113), .A2(n9112), .ZN(n9200) );
  AND2_X1 U11560 ( .A1(n9114), .A2(n9200), .ZN(n10183) );
  AOI22_X1 U11561 ( .A1(n9136), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6935), .B2(
        n10183), .ZN(n9115) );
  NAND2_X1 U11562 ( .A1(n9492), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9121) );
  NAND2_X1 U11563 ( .A1(n9116), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9130) );
  OR2_X1 U11564 ( .A1(n9116), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9117) );
  AND2_X1 U11565 ( .A1(n9130), .A2(n9117), .ZN(n10672) );
  NAND2_X1 U11566 ( .A1(n9454), .A2(n10672), .ZN(n9120) );
  NAND2_X1 U11567 ( .A1(n9493), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n9119) );
  NAND2_X1 U11568 ( .A1(n9466), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n9118) );
  NAND4_X1 U11569 ( .A1(n9121), .A2(n9120), .A3(n9119), .A4(n9118), .ZN(n13595) );
  MUX2_X1 U11570 ( .A(n14631), .B(n13595), .S(n9499), .Z(n9125) );
  NAND2_X1 U11571 ( .A1(n9124), .A2(n9125), .ZN(n9123) );
  MUX2_X1 U11572 ( .A(n13595), .B(n14631), .S(n9499), .Z(n9122) );
  NAND2_X1 U11573 ( .A1(n9123), .A2(n9122), .ZN(n9129) );
  INV_X1 U11574 ( .A(n9124), .ZN(n9127) );
  INV_X1 U11575 ( .A(n9125), .ZN(n9126) );
  NAND2_X1 U11576 ( .A1(n9130), .A2(n10764), .ZN(n9131) );
  AND2_X1 U11577 ( .A1(n9159), .A2(n9131), .ZN(n14556) );
  NAND2_X1 U11578 ( .A1(n9454), .A2(n14556), .ZN(n9135) );
  NAND2_X1 U11579 ( .A1(n9492), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n9134) );
  NAND2_X1 U11580 ( .A1(n9466), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n9133) );
  NAND2_X1 U11581 ( .A1(n9493), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9132) );
  NAND4_X1 U11582 ( .A1(n9135), .A2(n9134), .A3(n9133), .A4(n9132), .ZN(n13594) );
  OR2_X1 U11583 ( .A1(n9637), .A2(n9485), .ZN(n9139) );
  NAND2_X1 U11584 ( .A1(n9200), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9137) );
  XNOR2_X1 U11585 ( .A(n9137), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10171) );
  AOI22_X1 U11586 ( .A1(n9507), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6935), .B2(
        n10171), .ZN(n9138) );
  NAND2_X1 U11587 ( .A1(n9139), .A2(n9138), .ZN(n14558) );
  MUX2_X1 U11588 ( .A(n13594), .B(n14558), .S(n9499), .Z(n9141) );
  MUX2_X1 U11589 ( .A(n14558), .B(n13594), .S(n9499), .Z(n9140) );
  OR2_X1 U11590 ( .A1(n9707), .A2(n9485), .ZN(n9145) );
  OR2_X1 U11591 ( .A1(n9200), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9143) );
  NAND2_X1 U11592 ( .A1(n9143), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9165) );
  XNOR2_X1 U11593 ( .A(n9165), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10222) );
  AOI22_X1 U11594 ( .A1(n9507), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6935), .B2(
        n10222), .ZN(n9144) );
  NAND2_X1 U11595 ( .A1(n9145), .A2(n9144), .ZN(n11198) );
  NAND2_X1 U11596 ( .A1(n9492), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9149) );
  XNOR2_X1 U11597 ( .A(n9159), .B(P1_REG3_REG_8__SCAN_IN), .ZN(n11124) );
  NAND2_X1 U11598 ( .A1(n9454), .A2(n11124), .ZN(n9148) );
  NAND2_X1 U11599 ( .A1(n9493), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9147) );
  NAND2_X1 U11600 ( .A1(n9466), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n9146) );
  OR2_X1 U11601 ( .A1(n11198), .A2(n14536), .ZN(n11205) );
  NAND2_X1 U11602 ( .A1(n11198), .A2(n14536), .ZN(n9541) );
  MUX2_X1 U11603 ( .A(n11205), .B(n9541), .S(n9499), .Z(n9150) );
  NAND2_X1 U11604 ( .A1(n9151), .A2(n9150), .ZN(n9155) );
  INV_X1 U11605 ( .A(n14536), .ZN(n13593) );
  MUX2_X1 U11606 ( .A(n13593), .B(n11198), .S(n9473), .Z(n9153) );
  NAND2_X1 U11607 ( .A1(n11198), .A2(n13593), .ZN(n9152) );
  NAND2_X1 U11608 ( .A1(n9153), .A2(n9152), .ZN(n9154) );
  NAND2_X1 U11609 ( .A1(n9155), .A2(n9154), .ZN(n9171) );
  NAND2_X1 U11610 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .ZN(n9156) );
  INV_X1 U11611 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n9158) );
  INV_X1 U11612 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n9157) );
  OAI21_X1 U11613 ( .B1(n9159), .B2(n9158), .A(n9157), .ZN(n9160) );
  AND2_X1 U11614 ( .A1(n9174), .A2(n9160), .ZN(n14540) );
  NAND2_X1 U11615 ( .A1(n9454), .A2(n14540), .ZN(n9164) );
  NAND2_X1 U11616 ( .A1(n9492), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n9163) );
  NAND2_X1 U11617 ( .A1(n9466), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n9162) );
  NAND2_X1 U11618 ( .A1(n9493), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9161) );
  OR2_X1 U11619 ( .A1(n9742), .A2(n9485), .ZN(n9168) );
  INV_X1 U11620 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n15401) );
  NAND2_X1 U11621 ( .A1(n9165), .A2(n15401), .ZN(n9166) );
  NAND2_X1 U11622 ( .A1(n9166), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9183) );
  XNOR2_X1 U11623 ( .A(n9183), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10208) );
  AOI22_X1 U11624 ( .A1(n9507), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6935), .B2(
        n10208), .ZN(n9167) );
  MUX2_X1 U11625 ( .A(n11207), .B(n14658), .S(n9499), .Z(n9170) );
  INV_X1 U11626 ( .A(n11207), .ZN(n13592) );
  MUX2_X1 U11627 ( .A(n13592), .B(n14541), .S(n9473), .Z(n9169) );
  OAI21_X1 U11628 ( .B1(n9171), .B2(n9170), .A(n9169), .ZN(n9173) );
  NAND2_X1 U11629 ( .A1(n9171), .A2(n9170), .ZN(n9172) );
  INV_X1 U11630 ( .A(n9190), .ZN(n9176) );
  NAND2_X1 U11631 ( .A1(n9174), .A2(n15558), .ZN(n9175) );
  NAND2_X1 U11632 ( .A1(n9176), .A2(n9175), .ZN(n14364) );
  INV_X1 U11633 ( .A(n14364), .ZN(n9177) );
  NAND2_X1 U11634 ( .A1(n9454), .A2(n9177), .ZN(n9181) );
  NAND2_X1 U11635 ( .A1(n9492), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n9180) );
  NAND2_X1 U11636 ( .A1(n9466), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n9179) );
  NAND2_X1 U11637 ( .A1(n9493), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n9178) );
  NAND4_X1 U11638 ( .A1(n9181), .A2(n9180), .A3(n9179), .A4(n9178), .ZN(n13591) );
  OR2_X1 U11639 ( .A1(n9791), .A2(n9485), .ZN(n9187) );
  INV_X1 U11640 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9182) );
  NAND2_X1 U11641 ( .A1(n9183), .A2(n9182), .ZN(n9184) );
  NAND2_X1 U11642 ( .A1(n9184), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9185) );
  XNOR2_X1 U11643 ( .A(n9185), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10424) );
  AOI22_X1 U11644 ( .A1(n9507), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6935), 
        .B2(n10424), .ZN(n9186) );
  MUX2_X1 U11645 ( .A(n13591), .B(n14357), .S(n9473), .Z(n9189) );
  MUX2_X1 U11646 ( .A(n13591), .B(n14357), .S(n9510), .Z(n9188) );
  OR2_X1 U11647 ( .A1(n9190), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9191) );
  NAND2_X1 U11648 ( .A1(n9190), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9213) );
  AND2_X1 U11649 ( .A1(n9191), .A2(n9213), .ZN(n11269) );
  NAND2_X1 U11650 ( .A1(n9454), .A2(n11269), .ZN(n9195) );
  NAND2_X1 U11651 ( .A1(n9492), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n9194) );
  NAND2_X1 U11652 ( .A1(n9493), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n9193) );
  NAND2_X1 U11653 ( .A1(n9466), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n9192) );
  NAND4_X1 U11654 ( .A1(n9195), .A2(n9194), .A3(n9193), .A4(n9192), .ZN(n13590) );
  NAND2_X1 U11655 ( .A1(n9885), .A2(n9488), .ZN(n9203) );
  INV_X1 U11656 ( .A(n9196), .ZN(n9199) );
  INV_X1 U11657 ( .A(n9197), .ZN(n9198) );
  NAND2_X1 U11658 ( .A1(n9219), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9201) );
  XNOR2_X1 U11659 ( .A(n9201), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10426) );
  AOI22_X1 U11660 ( .A1(n9507), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6935), 
        .B2(n10426), .ZN(n9202) );
  MUX2_X1 U11661 ( .A(n13590), .B(n11356), .S(n9510), .Z(n9207) );
  NAND2_X1 U11662 ( .A1(n9206), .A2(n9207), .ZN(n9205) );
  MUX2_X1 U11663 ( .A(n13590), .B(n11356), .S(n9473), .Z(n9204) );
  NAND2_X1 U11664 ( .A1(n9205), .A2(n9204), .ZN(n9211) );
  INV_X1 U11665 ( .A(n9206), .ZN(n9209) );
  INV_X1 U11666 ( .A(n9207), .ZN(n9208) );
  NAND2_X1 U11667 ( .A1(n9211), .A2(n9210), .ZN(n9225) );
  INV_X1 U11668 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n9212) );
  NAND2_X1 U11669 ( .A1(n9213), .A2(n9212), .ZN(n9214) );
  AND2_X1 U11670 ( .A1(n9230), .A2(n9214), .ZN(n11365) );
  NAND2_X1 U11671 ( .A1(n9454), .A2(n11365), .ZN(n9218) );
  NAND2_X1 U11672 ( .A1(n9492), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n9217) );
  NAND2_X1 U11673 ( .A1(n9466), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n9216) );
  NAND2_X1 U11674 ( .A1(n9493), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n9215) );
  NAND4_X1 U11675 ( .A1(n9218), .A2(n9217), .A3(n9216), .A4(n9215), .ZN(n13589) );
  NAND2_X1 U11676 ( .A1(n10040), .A2(n9488), .ZN(n9222) );
  NAND2_X1 U11677 ( .A1(n9220), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9236) );
  XNOR2_X1 U11678 ( .A(n9236), .B(P1_IR_REG_12__SCAN_IN), .ZN(n13671) );
  AOI22_X1 U11679 ( .A1(n9507), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6935), 
        .B2(n13671), .ZN(n9221) );
  MUX2_X1 U11680 ( .A(n13589), .B(n14156), .S(n9473), .Z(n9226) );
  NAND2_X1 U11681 ( .A1(n9225), .A2(n9226), .ZN(n9224) );
  MUX2_X1 U11682 ( .A(n13589), .B(n14156), .S(n9510), .Z(n9223) );
  INV_X1 U11683 ( .A(n9225), .ZN(n9228) );
  INV_X1 U11684 ( .A(n9226), .ZN(n9227) );
  AND2_X1 U11685 ( .A1(n9230), .A2(n9229), .ZN(n9231) );
  NOR2_X1 U11686 ( .A1(n9248), .A2(n9231), .ZN(n14168) );
  NAND2_X1 U11687 ( .A1(n9454), .A2(n14168), .ZN(n9235) );
  NAND2_X1 U11688 ( .A1(n9492), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n9234) );
  NAND2_X1 U11689 ( .A1(n9466), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n9233) );
  NAND2_X1 U11690 ( .A1(n9493), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9232) );
  NAND4_X1 U11691 ( .A1(n9235), .A2(n9234), .A3(n9233), .A4(n9232), .ZN(n13588) );
  NAND2_X1 U11692 ( .A1(n10059), .A2(n9488), .ZN(n9239) );
  INV_X1 U11693 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n15355) );
  NAND2_X1 U11694 ( .A1(n9236), .A2(n15355), .ZN(n9237) );
  NAND2_X1 U11695 ( .A1(n9237), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9243) );
  XNOR2_X1 U11696 ( .A(n9243), .B(P1_IR_REG_13__SCAN_IN), .ZN(n14449) );
  AOI22_X1 U11697 ( .A1(n9507), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6935), 
        .B2(n14449), .ZN(n9238) );
  MUX2_X1 U11698 ( .A(n13588), .B(n14169), .S(n9499), .Z(n9241) );
  MUX2_X1 U11699 ( .A(n13588), .B(n14169), .S(n9473), .Z(n9240) );
  NAND2_X1 U11700 ( .A1(n10367), .A2(n9488), .ZN(n9247) );
  NAND2_X1 U11701 ( .A1(n9243), .A2(n9242), .ZN(n9244) );
  NAND2_X1 U11702 ( .A1(n9244), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9245) );
  XNOR2_X1 U11703 ( .A(n9245), .B(P1_IR_REG_14__SCAN_IN), .ZN(n14453) );
  AOI22_X1 U11704 ( .A1(n9507), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6935), 
        .B2(n14453), .ZN(n9246) );
  NAND2_X1 U11705 ( .A1(n9248), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9260) );
  OR2_X1 U11706 ( .A1(n9248), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9249) );
  NAND2_X1 U11707 ( .A1(n9260), .A2(n9249), .ZN(n14347) );
  INV_X1 U11708 ( .A(n14347), .ZN(n11416) );
  NAND2_X1 U11709 ( .A1(n9454), .A2(n11416), .ZN(n9253) );
  NAND2_X1 U11710 ( .A1(n9492), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n9252) );
  NAND2_X1 U11711 ( .A1(n9493), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9251) );
  NAND2_X1 U11712 ( .A1(n9466), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n9250) );
  NAND2_X1 U11713 ( .A1(n14383), .A2(n13912), .ZN(n9266) );
  NAND2_X1 U11714 ( .A1(n10518), .A2(n9488), .ZN(n9258) );
  NAND2_X1 U11715 ( .A1(n9254), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9255) );
  XNOR2_X1 U11716 ( .A(n9255), .B(n8990), .ZN(n14478) );
  INV_X1 U11717 ( .A(n14478), .ZN(n9256) );
  AOI22_X1 U11718 ( .A1(n9507), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6935), 
        .B2(n9256), .ZN(n9257) );
  NAND2_X1 U11719 ( .A1(n9466), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n9265) );
  INV_X1 U11720 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9259) );
  NAND2_X1 U11721 ( .A1(n9260), .A2(n9259), .ZN(n9261) );
  AND2_X1 U11722 ( .A1(n9275), .A2(n9261), .ZN(n13921) );
  NAND2_X1 U11723 ( .A1(n9454), .A2(n13921), .ZN(n9264) );
  NAND2_X1 U11724 ( .A1(n9492), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n9263) );
  NAND2_X1 U11725 ( .A1(n9493), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n9262) );
  NAND2_X1 U11726 ( .A1(n14375), .A2(n13899), .ZN(n9536) );
  NAND2_X1 U11727 ( .A1(n9536), .A2(n9266), .ZN(n9268) );
  NAND2_X1 U11728 ( .A1(n11782), .A2(n11780), .ZN(n9267) );
  MUX2_X1 U11729 ( .A(n9268), .B(n9267), .S(n9510), .Z(n9269) );
  AOI21_X1 U11730 ( .B1(n9270), .B2(n11426), .A(n9269), .ZN(n9271) );
  INV_X1 U11731 ( .A(n9271), .ZN(n9273) );
  MUX2_X1 U11732 ( .A(n9536), .B(n11782), .S(n9473), .Z(n9272) );
  INV_X1 U11733 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9274) );
  AND2_X1 U11734 ( .A1(n9275), .A2(n9274), .ZN(n9276) );
  NOR2_X1 U11735 ( .A1(n9300), .A2(n9276), .ZN(n13900) );
  NAND2_X1 U11736 ( .A1(n9454), .A2(n13900), .ZN(n9280) );
  NAND2_X1 U11737 ( .A1(n9492), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9279) );
  NAND2_X1 U11738 ( .A1(n9466), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n9278) );
  NAND2_X1 U11739 ( .A1(n9493), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9277) );
  NAND4_X1 U11740 ( .A1(n9280), .A2(n9279), .A3(n9278), .A4(n9277), .ZN(n13914) );
  NAND2_X1 U11741 ( .A1(n10344), .A2(n9488), .ZN(n9284) );
  NAND2_X1 U11742 ( .A1(n9281), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9282) );
  XNOR2_X1 U11743 ( .A(n9282), .B(P1_IR_REG_16__SCAN_IN), .ZN(n14493) );
  AOI22_X1 U11744 ( .A1(n9507), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6935), 
        .B2(n14493), .ZN(n9283) );
  MUX2_X1 U11745 ( .A(n13914), .B(n14367), .S(n9510), .Z(n9321) );
  INV_X1 U11746 ( .A(n13914), .ZN(n13570) );
  INV_X1 U11747 ( .A(n14367), .ZN(n13515) );
  MUX2_X1 U11748 ( .A(n13570), .B(n13515), .S(n9473), .Z(n9285) );
  OAI21_X1 U11749 ( .B1(n9322), .B2(n9321), .A(n9285), .ZN(n9324) );
  NAND2_X1 U11750 ( .A1(n10920), .A2(n9488), .ZN(n9287) );
  AOI22_X1 U11751 ( .A1(n9507), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n10878), 
        .B2(n6935), .ZN(n9286) );
  NAND2_X2 U11752 ( .A1(n9287), .A2(n9286), .ZN(n13852) );
  INV_X1 U11753 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9288) );
  NAND2_X1 U11754 ( .A1(n9315), .A2(n9288), .ZN(n9289) );
  AND2_X1 U11755 ( .A1(n9341), .A2(n9289), .ZN(n13856) );
  NAND2_X1 U11756 ( .A1(n13856), .A2(n9454), .ZN(n9293) );
  NAND2_X1 U11757 ( .A1(n9466), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n9292) );
  NAND2_X1 U11758 ( .A1(n9493), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n9291) );
  NAND2_X1 U11759 ( .A1(n9492), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n9290) );
  NAND4_X1 U11760 ( .A1(n9293), .A2(n9292), .A3(n9291), .A4(n9290), .ZN(n13584) );
  XNOR2_X1 U11761 ( .A(n13852), .B(n13584), .ZN(n13850) );
  NAND2_X1 U11762 ( .A1(n10522), .A2(n9488), .ZN(n9299) );
  INV_X1 U11763 ( .A(n9295), .ZN(n9296) );
  NAND2_X1 U11764 ( .A1(n9296), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9297) );
  XNOR2_X1 U11765 ( .A(n9297), .B(P1_IR_REG_17__SCAN_IN), .ZN(n13676) );
  AOI22_X1 U11766 ( .A1(n9507), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6935), 
        .B2(n13676), .ZN(n9298) );
  NOR2_X1 U11767 ( .A1(n9300), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9301) );
  NOR2_X1 U11768 ( .A1(n9313), .A2(n9301), .ZN(n13890) );
  NAND2_X1 U11769 ( .A1(n9454), .A2(n13890), .ZN(n9305) );
  NAND2_X1 U11770 ( .A1(n9492), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9304) );
  NAND2_X1 U11771 ( .A1(n9466), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n9303) );
  NAND2_X1 U11772 ( .A1(n9493), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9302) );
  NAND4_X1 U11773 ( .A1(n9305), .A2(n9304), .A3(n9303), .A4(n9302), .ZN(n13585) );
  OR2_X1 U11774 ( .A1(n14015), .A2(n13585), .ZN(n11763) );
  NAND2_X1 U11775 ( .A1(n14015), .A2(n13585), .ZN(n11764) );
  NAND2_X1 U11776 ( .A1(n11763), .A2(n11764), .ZN(n13884) );
  NAND2_X1 U11777 ( .A1(n9306), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9308) );
  XNOR2_X1 U11778 ( .A(n9307), .B(n9308), .ZN(n14524) );
  INV_X1 U11779 ( .A(n14524), .ZN(n9309) );
  AOI22_X1 U11780 ( .A1(n9507), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6935), 
        .B2(n9309), .ZN(n9311) );
  OR2_X1 U11781 ( .A1(n9313), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9314) );
  AND2_X1 U11782 ( .A1(n9315), .A2(n9314), .ZN(n13876) );
  NAND2_X1 U11783 ( .A1(n9454), .A2(n13876), .ZN(n9319) );
  NAND2_X1 U11784 ( .A1(n9492), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9318) );
  NAND2_X1 U11785 ( .A1(n9466), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n9317) );
  NAND2_X1 U11786 ( .A1(n9493), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9316) );
  NAND4_X1 U11787 ( .A1(n9319), .A2(n9318), .A3(n9317), .A4(n9316), .ZN(n13853) );
  XNOR2_X1 U11788 ( .A(n14009), .B(n13853), .ZN(n9320) );
  NAND2_X1 U11789 ( .A1(n9324), .A2(n9323), .ZN(n9337) );
  INV_X1 U11790 ( .A(n13853), .ZN(n13406) );
  NAND2_X1 U11791 ( .A1(n9499), .A2(n13585), .ZN(n9326) );
  INV_X1 U11792 ( .A(n13585), .ZN(n13898) );
  NAND2_X1 U11793 ( .A1(n9473), .A2(n13898), .ZN(n9325) );
  MUX2_X1 U11794 ( .A(n9326), .B(n9325), .S(n14015), .Z(n9328) );
  NAND2_X1 U11795 ( .A1(n9328), .A2(n13406), .ZN(n9327) );
  OAI211_X1 U11796 ( .C1(n13406), .C2(n9499), .A(n13878), .B(n9327), .ZN(n9331) );
  NAND2_X1 U11797 ( .A1(n9328), .A2(n13853), .ZN(n9329) );
  OAI211_X1 U11798 ( .C1(n9473), .C2(n13853), .A(n9329), .B(n14009), .ZN(n9330) );
  NAND2_X1 U11799 ( .A1(n9331), .A2(n9330), .ZN(n9332) );
  NAND2_X1 U11800 ( .A1(n13850), .A2(n9332), .ZN(n9335) );
  INV_X1 U11801 ( .A(n13584), .ZN(n13872) );
  OR2_X1 U11802 ( .A1(n13852), .A2(n13872), .ZN(n9333) );
  NAND2_X1 U11803 ( .A1(n13852), .A2(n13872), .ZN(n11787) );
  MUX2_X1 U11804 ( .A(n9333), .B(n11787), .S(n9473), .Z(n9334) );
  AND2_X1 U11805 ( .A1(n9335), .A2(n9334), .ZN(n9336) );
  NAND2_X1 U11806 ( .A1(n9337), .A2(n9336), .ZN(n9351) );
  NAND2_X1 U11807 ( .A1(n9466), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n9339) );
  NAND2_X1 U11808 ( .A1(n9493), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n9338) );
  AND2_X1 U11809 ( .A1(n9339), .A2(n9338), .ZN(n9346) );
  INV_X1 U11810 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9340) );
  NAND2_X1 U11811 ( .A1(n9341), .A2(n9340), .ZN(n9342) );
  INV_X1 U11812 ( .A(n9354), .ZN(n9355) );
  NAND2_X1 U11813 ( .A1(n9342), .A2(n9355), .ZN(n13842) );
  OR2_X1 U11814 ( .A1(n9343), .A2(n13842), .ZN(n9345) );
  NAND2_X1 U11815 ( .A1(n9492), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n9344) );
  OR2_X1 U11816 ( .A1(n11826), .A2(n9485), .ZN(n9348) );
  NAND2_X1 U11817 ( .A1(n9507), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9347) );
  MUX2_X1 U11818 ( .A(n13827), .B(n13995), .S(n9510), .Z(n9350) );
  MUX2_X1 U11819 ( .A(n13855), .B(n13536), .S(n9473), .Z(n9349) );
  NAND2_X1 U11820 ( .A1(n9351), .A2(n9350), .ZN(n9352) );
  INV_X1 U11821 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n13492) );
  AOI21_X1 U11822 ( .B1(n13492), .B2(n9355), .A(n9365), .ZN(n13819) );
  NAND2_X1 U11823 ( .A1(n9454), .A2(n13819), .ZN(n9359) );
  NAND2_X1 U11824 ( .A1(n9492), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n9358) );
  NAND2_X1 U11825 ( .A1(n9466), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n9357) );
  NAND2_X1 U11826 ( .A1(n9493), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n9356) );
  NAND4_X1 U11827 ( .A1(n9359), .A2(n9358), .A3(n9357), .A4(n9356), .ZN(n13583) );
  OR2_X1 U11828 ( .A1(n10999), .A2(n9485), .ZN(n9361) );
  NAND2_X1 U11829 ( .A1(n9507), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9360) );
  MUX2_X1 U11830 ( .A(n13583), .B(n13990), .S(n9473), .Z(n9363) );
  MUX2_X1 U11831 ( .A(n13583), .B(n13990), .S(n9510), .Z(n9362) );
  INV_X1 U11832 ( .A(n9363), .ZN(n9364) );
  NAND2_X1 U11833 ( .A1(n9492), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n9370) );
  OAI21_X1 U11834 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n9365), .A(n9382), .ZN(
        n9366) );
  INV_X1 U11835 ( .A(n9366), .ZN(n13806) );
  NAND2_X1 U11836 ( .A1(n9454), .A2(n13806), .ZN(n9369) );
  NAND2_X1 U11837 ( .A1(n9493), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n9368) );
  NAND2_X1 U11838 ( .A1(n9466), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n9367) );
  NAND4_X1 U11839 ( .A1(n9370), .A2(n9369), .A3(n9368), .A4(n9367), .ZN(n13825) );
  OR2_X1 U11840 ( .A1(n9372), .A2(n9371), .ZN(n9373) );
  XNOR2_X1 U11841 ( .A(n9373), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14043) );
  MUX2_X1 U11842 ( .A(n13825), .B(n13812), .S(n9510), .Z(n9377) );
  NAND2_X1 U11843 ( .A1(n9376), .A2(n9377), .ZN(n9375) );
  MUX2_X1 U11844 ( .A(n13825), .B(n13812), .S(n9473), .Z(n9374) );
  NAND2_X1 U11845 ( .A1(n9375), .A2(n9374), .ZN(n9381) );
  INV_X1 U11846 ( .A(n9376), .ZN(n9379) );
  INV_X1 U11847 ( .A(n9377), .ZN(n9378) );
  NAND2_X1 U11848 ( .A1(n9381), .A2(n9380), .ZN(n9391) );
  INV_X1 U11849 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n15432) );
  AOI21_X1 U11850 ( .B1(n15432), .B2(n9382), .A(n9397), .ZN(n13791) );
  NAND2_X1 U11851 ( .A1(n9454), .A2(n13791), .ZN(n9386) );
  NAND2_X1 U11852 ( .A1(n9492), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n9385) );
  NAND2_X1 U11853 ( .A1(n9466), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n9384) );
  NAND2_X1 U11854 ( .A1(n9493), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n9383) );
  NAND4_X1 U11855 ( .A1(n9386), .A2(n9385), .A3(n9384), .A4(n9383), .ZN(n13582) );
  NAND2_X1 U11856 ( .A1(n11308), .A2(n9488), .ZN(n9388) );
  NAND2_X1 U11857 ( .A1(n9507), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n9387) );
  MUX2_X1 U11858 ( .A(n13582), .B(n13979), .S(n9473), .Z(n9392) );
  NAND2_X1 U11859 ( .A1(n9391), .A2(n9392), .ZN(n9390) );
  MUX2_X1 U11860 ( .A(n13582), .B(n13979), .S(n9510), .Z(n9389) );
  NAND2_X1 U11861 ( .A1(n9390), .A2(n9389), .ZN(n9396) );
  INV_X1 U11862 ( .A(n9391), .ZN(n9394) );
  INV_X1 U11863 ( .A(n9392), .ZN(n9393) );
  INV_X1 U11864 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n13525) );
  INV_X1 U11865 ( .A(n9397), .ZN(n9398) );
  NAND2_X1 U11866 ( .A1(n9397), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n9409) );
  AOI21_X1 U11867 ( .B1(n13525), .B2(n9398), .A(n9408), .ZN(n13778) );
  NAND2_X1 U11868 ( .A1(n9454), .A2(n13778), .ZN(n9402) );
  NAND2_X1 U11869 ( .A1(n9492), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n9401) );
  NAND2_X1 U11870 ( .A1(n9466), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n9400) );
  NAND2_X1 U11871 ( .A1(n9493), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n9399) );
  NAND4_X1 U11872 ( .A1(n9402), .A2(n9401), .A3(n9400), .A4(n9399), .ZN(n13581) );
  OR2_X1 U11873 ( .A1(n11334), .A2(n9485), .ZN(n9404) );
  NAND2_X1 U11874 ( .A1(n9507), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n9403) );
  MUX2_X1 U11875 ( .A(n13581), .B(n13973), .S(n9510), .Z(n9406) );
  MUX2_X1 U11876 ( .A(n13581), .B(n13973), .S(n9473), .Z(n9405) );
  INV_X1 U11877 ( .A(n9406), .ZN(n9407) );
  INV_X1 U11878 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n13502) );
  NAND2_X1 U11879 ( .A1(n9408), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n9424) );
  INV_X1 U11880 ( .A(n9424), .ZN(n9426) );
  AOI21_X1 U11881 ( .B1(n13502), .B2(n9409), .A(n9426), .ZN(n13760) );
  NAND2_X1 U11882 ( .A1(n9454), .A2(n13760), .ZN(n9413) );
  NAND2_X1 U11883 ( .A1(n9492), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n9412) );
  NAND2_X1 U11884 ( .A1(n9466), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n9411) );
  NAND2_X1 U11885 ( .A1(n9493), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n9410) );
  NAND4_X1 U11886 ( .A1(n9413), .A2(n9412), .A3(n9411), .A4(n9410), .ZN(n13736) );
  NAND2_X1 U11887 ( .A1(n11460), .A2(n9488), .ZN(n9415) );
  NAND2_X1 U11888 ( .A1(n9507), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n9414) );
  MUX2_X1 U11889 ( .A(n13736), .B(n13965), .S(n9473), .Z(n9419) );
  NAND2_X1 U11890 ( .A1(n9418), .A2(n9419), .ZN(n9417) );
  MUX2_X1 U11891 ( .A(n13736), .B(n13965), .S(n9510), .Z(n9416) );
  NAND2_X1 U11892 ( .A1(n9417), .A2(n9416), .ZN(n9423) );
  INV_X1 U11893 ( .A(n9418), .ZN(n9421) );
  INV_X1 U11894 ( .A(n9419), .ZN(n9420) );
  NAND2_X1 U11895 ( .A1(n9492), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n9431) );
  INV_X1 U11896 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9425) );
  NAND2_X1 U11897 ( .A1(n9425), .A2(n9424), .ZN(n9427) );
  NAND2_X1 U11898 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(n9426), .ZN(n9438) );
  AND2_X1 U11899 ( .A1(n9427), .A2(n9438), .ZN(n13740) );
  NAND2_X1 U11900 ( .A1(n9454), .A2(n13740), .ZN(n9430) );
  NAND2_X1 U11901 ( .A1(n9493), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n9429) );
  NAND2_X1 U11902 ( .A1(n9466), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n9428) );
  NAND2_X1 U11903 ( .A1(n9507), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9432) );
  MUX2_X1 U11904 ( .A(n13580), .B(n13957), .S(n9510), .Z(n9435) );
  MUX2_X1 U11905 ( .A(n13957), .B(n13580), .S(n9499), .Z(n9434) );
  INV_X1 U11906 ( .A(n9438), .ZN(n9436) );
  NAND2_X1 U11907 ( .A1(n9436), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n9465) );
  INV_X1 U11908 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9437) );
  NAND2_X1 U11909 ( .A1(n9438), .A2(n9437), .ZN(n9439) );
  NAND2_X1 U11910 ( .A1(n9454), .A2(n13723), .ZN(n9443) );
  NAND2_X1 U11911 ( .A1(n9492), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n9442) );
  NAND2_X1 U11912 ( .A1(n9466), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n9441) );
  NAND2_X1 U11913 ( .A1(n9493), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n9440) );
  NAND4_X1 U11914 ( .A1(n9443), .A2(n9442), .A3(n9441), .A4(n9440), .ZN(n13737) );
  NAND2_X1 U11915 ( .A1(n9507), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9444) );
  MUX2_X1 U11916 ( .A(n13737), .B(n13951), .S(n9473), .Z(n9449) );
  NAND2_X1 U11917 ( .A1(n9448), .A2(n9449), .ZN(n9447) );
  MUX2_X1 U11918 ( .A(n13737), .B(n13951), .S(n9499), .Z(n9446) );
  NAND2_X1 U11919 ( .A1(n9447), .A2(n9446), .ZN(n9453) );
  INV_X1 U11920 ( .A(n9448), .ZN(n9451) );
  INV_X1 U11921 ( .A(n9449), .ZN(n9450) );
  NAND2_X1 U11922 ( .A1(n9451), .A2(n9450), .ZN(n9452) );
  XNOR2_X1 U11923 ( .A(n9465), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n13710) );
  NAND2_X1 U11924 ( .A1(n9454), .A2(n13710), .ZN(n9458) );
  NAND2_X1 U11925 ( .A1(n9492), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n9457) );
  NAND2_X1 U11926 ( .A1(n9466), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n9456) );
  NAND2_X1 U11927 ( .A1(n9493), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n9455) );
  NAND4_X1 U11928 ( .A1(n9458), .A2(n9457), .A3(n9456), .A4(n9455), .ZN(n13579) );
  NAND2_X1 U11929 ( .A1(n13351), .A2(n9488), .ZN(n9460) );
  NAND2_X1 U11930 ( .A1(n9507), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9459) );
  MUX2_X1 U11931 ( .A(n13579), .B(n13943), .S(n9510), .Z(n9462) );
  MUX2_X1 U11932 ( .A(n13579), .B(n13943), .S(n9473), .Z(n9461) );
  INV_X1 U11933 ( .A(n9462), .ZN(n9463) );
  INV_X1 U11934 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9464) );
  NOR2_X1 U11935 ( .A1(n9465), .A2(n9464), .ZN(n11806) );
  NAND2_X1 U11936 ( .A1(n9454), .A2(n11806), .ZN(n9470) );
  NAND2_X1 U11937 ( .A1(n9492), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n9469) );
  NAND2_X1 U11938 ( .A1(n9466), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n9468) );
  NAND2_X1 U11939 ( .A1(n9493), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n9467) );
  NAND4_X1 U11940 ( .A1(n9470), .A2(n9469), .A3(n9468), .A4(n9467), .ZN(n13578) );
  NAND2_X1 U11941 ( .A1(n13347), .A2(n9488), .ZN(n9472) );
  NAND2_X1 U11942 ( .A1(n9507), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n9471) );
  MUX2_X1 U11943 ( .A(n13578), .B(n13941), .S(n9473), .Z(n9477) );
  NAND2_X1 U11944 ( .A1(n9476), .A2(n9477), .ZN(n9475) );
  MUX2_X1 U11945 ( .A(n13578), .B(n13941), .S(n9499), .Z(n9474) );
  NAND2_X1 U11946 ( .A1(n9475), .A2(n9474), .ZN(n9481) );
  INV_X1 U11947 ( .A(n9476), .ZN(n9479) );
  INV_X1 U11948 ( .A(n9477), .ZN(n9478) );
  NAND2_X1 U11949 ( .A1(n9479), .A2(n9478), .ZN(n9480) );
  NAND2_X1 U11950 ( .A1(n9481), .A2(n9480), .ZN(n9519) );
  MUX2_X1 U11951 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n8205), .Z(n9502) );
  XNOR2_X1 U11952 ( .A(n9502), .B(SI_30_), .ZN(n9503) );
  INV_X1 U11953 ( .A(n12012), .ZN(n13345) );
  INV_X1 U11954 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n11828) );
  INV_X1 U11955 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n15449) );
  NAND2_X1 U11956 ( .A1(n9492), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n9490) );
  NAND2_X1 U11957 ( .A1(n9466), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n9489) );
  OAI211_X1 U11958 ( .C1(n9491), .C2(n15449), .A(n9490), .B(n9489), .ZN(n13577) );
  NAND2_X1 U11959 ( .A1(n9492), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n9496) );
  NAND2_X1 U11960 ( .A1(n9493), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n9495) );
  NAND2_X1 U11961 ( .A1(n9466), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n9494) );
  AND3_X1 U11962 ( .A1(n9496), .A2(n9495), .A3(n9494), .ZN(n9516) );
  OAI22_X1 U11963 ( .A1(n9499), .A2(n9516), .B1(n10008), .B2(n9497), .ZN(n9498) );
  AOI22_X1 U11964 ( .A1(n13690), .A2(n9499), .B1(n13577), .B2(n9498), .ZN(
        n9513) );
  INV_X1 U11965 ( .A(n9516), .ZN(n13694) );
  INV_X1 U11966 ( .A(n11825), .ZN(n10879) );
  NAND2_X1 U11967 ( .A1(n10008), .A2(n10879), .ZN(n10308) );
  OAI21_X1 U11968 ( .B1(n13694), .B2(n10308), .A(n13577), .ZN(n9500) );
  MUX2_X1 U11969 ( .A(n13935), .B(n9500), .S(n9499), .Z(n9514) );
  INV_X1 U11970 ( .A(n9514), .ZN(n9501) );
  NOR2_X1 U11971 ( .A1(n9513), .A2(n9501), .ZN(n9522) );
  MUX2_X1 U11972 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n8205), .Z(n9505) );
  XNOR2_X1 U11973 ( .A(n9505), .B(SI_31_), .ZN(n9506) );
  NAND2_X1 U11974 ( .A1(n9507), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n9508) );
  NAND2_X1 U11975 ( .A1(n10013), .A2(n10878), .ZN(n10890) );
  NAND2_X1 U11976 ( .A1(n10298), .A2(n10008), .ZN(n10007) );
  OAI21_X1 U11977 ( .B1(n10879), .B2(n10298), .A(n10007), .ZN(n9512) );
  NAND2_X1 U11978 ( .A1(n10890), .A2(n9512), .ZN(n9528) );
  NAND2_X1 U11979 ( .A1(n7399), .A2(n10879), .ZN(n9552) );
  AND2_X1 U11980 ( .A1(n9528), .A2(n9552), .ZN(n9525) );
  NAND2_X1 U11981 ( .A1(n9526), .A2(n9525), .ZN(n9520) );
  INV_X1 U11982 ( .A(n9513), .ZN(n9515) );
  NOR2_X1 U11983 ( .A1(n9515), .A2(n9514), .ZN(n9524) );
  INV_X1 U11984 ( .A(n9521), .ZN(n9517) );
  NOR2_X1 U11985 ( .A1(n9524), .A2(n9517), .ZN(n9518) );
  INV_X1 U11986 ( .A(n9520), .ZN(n9523) );
  AOI22_X1 U11987 ( .A1(n9524), .A2(n9523), .B1(n9522), .B2(n9521), .ZN(n9530)
         );
  NAND2_X1 U11988 ( .A1(n9551), .A2(n9525), .ZN(n9527) );
  MUX2_X1 U11989 ( .A(n9528), .B(n9527), .S(n9526), .Z(n9529) );
  INV_X1 U11990 ( .A(n13578), .ZN(n13705) );
  XNOR2_X1 U11991 ( .A(n13941), .B(n13705), .ZN(n11800) );
  NAND2_X1 U11992 ( .A1(n13943), .A2(n13579), .ZN(n11779) );
  OR2_X1 U11993 ( .A1(n13943), .A2(n13579), .ZN(n9533) );
  NAND2_X1 U11994 ( .A1(n11779), .A2(n9533), .ZN(n13714) );
  NAND2_X1 U11995 ( .A1(n13951), .A2(n13704), .ZN(n11797) );
  OR2_X1 U11996 ( .A1(n13951), .A2(n13704), .ZN(n9534) );
  INV_X1 U11997 ( .A(n13736), .ZN(n9535) );
  XNOR2_X1 U11998 ( .A(n13965), .B(n9535), .ZN(n11794) );
  XNOR2_X1 U11999 ( .A(n13973), .B(n13581), .ZN(n13770) );
  XNOR2_X1 U12000 ( .A(n13536), .B(n13827), .ZN(n13832) );
  NAND2_X1 U12001 ( .A1(n14009), .A2(n13853), .ZN(n11765) );
  NAND2_X1 U12002 ( .A1(n11782), .A2(n9536), .ZN(n13923) );
  XNOR2_X1 U12003 ( .A(n14169), .B(n11415), .ZN(n14171) );
  INV_X1 U12004 ( .A(n13590), .ZN(n11355) );
  XNOR2_X1 U12005 ( .A(n11356), .B(n11355), .ZN(n11353) );
  INV_X1 U12006 ( .A(n13589), .ZN(n9537) );
  OR2_X1 U12007 ( .A1(n14156), .A2(n9537), .ZN(n11409) );
  NAND2_X1 U12008 ( .A1(n14156), .A2(n9537), .ZN(n9538) );
  NAND2_X1 U12009 ( .A1(n11409), .A2(n9538), .ZN(n11421) );
  XNOR2_X1 U12010 ( .A(n13596), .B(n10898), .ZN(n10893) );
  XNOR2_X1 U12011 ( .A(n13595), .B(n11127), .ZN(n11128) );
  INV_X1 U12012 ( .A(n10862), .ZN(n10307) );
  NAND2_X1 U12013 ( .A1(n10302), .A2(n9539), .ZN(n10915) );
  NOR2_X1 U12014 ( .A1(n10307), .A2(n10915), .ZN(n9540) );
  XNOR2_X2 U12015 ( .A(n10152), .B(n10976), .ZN(n10353) );
  XNOR2_X1 U12016 ( .A(n10867), .B(n11072), .ZN(n11074) );
  NAND4_X1 U12017 ( .A1(n9540), .A2(n11090), .A3(n10347), .A4(n11074), .ZN(
        n9542) );
  NAND2_X1 U12018 ( .A1(n11205), .A2(n9541), .ZN(n11196) );
  NOR4_X1 U12019 ( .A1(n10893), .A2(n11128), .A3(n9542), .A4(n11196), .ZN(
        n9543) );
  XNOR2_X1 U12020 ( .A(n14357), .B(n13591), .ZN(n11208) );
  XNOR2_X1 U12021 ( .A(n14541), .B(n13592), .ZN(n11199) );
  XNOR2_X1 U12022 ( .A(n14558), .B(n13594), .ZN(n14549) );
  NAND4_X1 U12023 ( .A1(n9543), .A2(n11208), .A3(n11199), .A4(n14549), .ZN(
        n9544) );
  NOR4_X1 U12024 ( .A1(n14171), .A2(n11353), .A3(n11421), .A4(n9544), .ZN(
        n9545) );
  XNOR2_X1 U12025 ( .A(n14367), .B(n13914), .ZN(n11783) );
  NAND4_X1 U12026 ( .A1(n13884), .A2(n11426), .A3(n9545), .A4(n11783), .ZN(
        n9546) );
  NOR4_X1 U12027 ( .A1(n13832), .A2(n11784), .A3(n13923), .A4(n9546), .ZN(
        n9547) );
  XNOR2_X1 U12028 ( .A(n13990), .B(n13583), .ZN(n13823) );
  NAND4_X1 U12029 ( .A1(n13770), .A2(n9547), .A3(n13850), .A4(n13823), .ZN(
        n9548) );
  INV_X1 U12030 ( .A(n13582), .ZN(n11791) );
  XNOR2_X1 U12031 ( .A(n13979), .B(n11791), .ZN(n13786) );
  XNOR2_X1 U12032 ( .A(n13983), .B(n13825), .ZN(n13808) );
  NOR4_X1 U12033 ( .A1(n11794), .A2(n9548), .A3(n13786), .A4(n13808), .ZN(
        n9549) );
  XNOR2_X1 U12034 ( .A(n13957), .B(n13580), .ZN(n13731) );
  NAND4_X1 U12035 ( .A1(n13714), .A2(n13728), .A3(n9549), .A4(n13731), .ZN(
        n9550) );
  INV_X1 U12036 ( .A(n9793), .ZN(n9558) );
  NAND2_X1 U12037 ( .A1(n9560), .A2(n9559), .ZN(n9575) );
  NAND2_X1 U12038 ( .A1(n9567), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9561) );
  NAND2_X1 U12039 ( .A1(n9562), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9563) );
  INV_X1 U12040 ( .A(n9564), .ZN(n9565) );
  NAND2_X1 U12041 ( .A1(n9565), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9566) );
  MUX2_X1 U12042 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9566), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n9568) );
  NAND2_X1 U12043 ( .A1(n11825), .A2(n13685), .ZN(n10009) );
  NAND2_X1 U12044 ( .A1(n10023), .A2(n10009), .ZN(n10450) );
  NAND2_X1 U12045 ( .A1(n10871), .A2(n10450), .ZN(n10293) );
  INV_X1 U12046 ( .A(n9571), .ZN(n13614) );
  NOR3_X1 U12047 ( .A1(n10293), .A2(n6641), .A3(n14537), .ZN(n9573) );
  OAI21_X1 U12048 ( .B1(n11305), .B2(n10298), .A(P1_B_REG_SCAN_IN), .ZN(n9572)
         );
  OR2_X1 U12049 ( .A1(n9573), .A2(n9572), .ZN(n9574) );
  NAND2_X1 U12050 ( .A1(n9575), .A2(n9574), .ZN(P1_U3242) );
  INV_X1 U12051 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n9585) );
  INV_X1 U12052 ( .A(n9937), .ZN(n9576) );
  NAND2_X1 U12053 ( .A1(n9577), .A2(n9576), .ZN(n9957) );
  NAND2_X1 U12054 ( .A1(n11711), .A2(n9950), .ZN(n11754) );
  OR2_X1 U12055 ( .A1(n9579), .A2(n11747), .ZN(n9938) );
  AND2_X1 U12056 ( .A1(n11754), .A2(n9938), .ZN(n9580) );
  OR2_X1 U12057 ( .A1(n9581), .A2(n9936), .ZN(n9947) );
  NAND2_X1 U12058 ( .A1(n9954), .A2(n9951), .ZN(n9582) );
  NAND2_X1 U12059 ( .A1(n11309), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9587) );
  NOR2_X1 U12060 ( .A1(n10451), .A2(P1_U3086), .ZN(n9588) );
  INV_X1 U12061 ( .A(n9589), .ZN(n9940) );
  AND2_X1 U12062 ( .A1(n8205), .A2(P2_U3088), .ZN(n13350) );
  INV_X2 U12063 ( .A(n13350), .ZN(n13359) );
  INV_X1 U12064 ( .A(n9659), .ZN(n9661) );
  NAND2_X1 U12065 ( .A1(n9661), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14695) );
  NOR2_X1 U12066 ( .A1(n8205), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13342) );
  NAND2_X1 U12067 ( .A1(n13342), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n9590) );
  OAI211_X1 U12068 ( .C1(n9606), .C2(n13359), .A(n14695), .B(n9590), .ZN(
        P2_U3326) );
  NAND2_X1 U12069 ( .A1(n8205), .A2(P3_U3151), .ZN(n12787) );
  NOR2_X2 U12070 ( .A1(n8205), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12775) );
  INV_X1 U12071 ( .A(n12775), .ZN(n12785) );
  OAI222_X1 U12072 ( .A1(P3_U3151), .A2(n9836), .B1(n12787), .B2(n6891), .C1(
        n12785), .C2(n9591), .ZN(P3_U3294) );
  OAI222_X1 U12073 ( .A1(n12785), .A2(n9593), .B1(n12787), .B2(n9592), .C1(
        n10808), .C2(P3_U3151), .ZN(P3_U3287) );
  INV_X1 U12074 ( .A(SI_10_), .ZN(n9594) );
  OAI222_X1 U12075 ( .A1(n12785), .A2(n9595), .B1(n12787), .B2(n9594), .C1(
        n15033), .C2(P3_U3151), .ZN(P3_U3285) );
  INV_X2 U12076 ( .A(n13342), .ZN(n13357) );
  OAI222_X1 U12077 ( .A1(n13357), .A2(n9596), .B1(n13359), .B2(n9608), .C1(
        n9686), .C2(P2_U3088), .ZN(P2_U3324) );
  OAI222_X1 U12078 ( .A1(n10812), .A2(P3_U3151), .B1(n12785), .B2(n9598), .C1(
        n9597), .C2(n12787), .ZN(P3_U3289) );
  OAI222_X1 U12079 ( .A1(n13357), .A2(n9599), .B1(n13359), .B2(n9603), .C1(
        n9687), .C2(P2_U3088), .ZN(P2_U3323) );
  OAI222_X1 U12080 ( .A1(P2_U3088), .A2(n14714), .B1(n13357), .B2(n9600), .C1(
        n13359), .C2(n9610), .ZN(P2_U3325) );
  OAI222_X1 U12081 ( .A1(n12785), .A2(n9601), .B1(n15041), .B2(P3_U3151), .C1(
        n12787), .C2(n15428), .ZN(P3_U3284) );
  INV_X1 U12082 ( .A(n13645), .ZN(n9604) );
  NOR2_X1 U12083 ( .A1(n8205), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11524) );
  INV_X2 U12084 ( .A(n11524), .ZN(n10724) );
  NAND2_X2 U12085 ( .A1(n8205), .A2(P1_U3086), .ZN(n14039) );
  OAI222_X1 U12086 ( .A1(P1_U3086), .A2(n9604), .B1(n10724), .B2(n9603), .C1(
        n9602), .C2(n14039), .ZN(P1_U3351) );
  OAI222_X1 U12087 ( .A1(P1_U3086), .A2(n10128), .B1(n10724), .B2(n9606), .C1(
        n9605), .C2(n14039), .ZN(P1_U3354) );
  OAI222_X1 U12088 ( .A1(P1_U3086), .A2(n13630), .B1(n10724), .B2(n9608), .C1(
        n9607), .C2(n14039), .ZN(P1_U3352) );
  INV_X1 U12089 ( .A(n13620), .ZN(n10130) );
  OAI222_X1 U12090 ( .A1(P1_U3086), .A2(n10130), .B1(n10724), .B2(n9610), .C1(
        n9609), .C2(n14039), .ZN(P1_U3353) );
  INV_X1 U12091 ( .A(n12773), .ZN(n9612) );
  NAND2_X1 U12092 ( .A1(n9612), .A2(n10279), .ZN(n9611) );
  OAI21_X1 U12093 ( .B1(n9612), .B2(n8495), .A(n9611), .ZN(P3_U3377) );
  OAI222_X1 U12094 ( .A1(n13357), .A2(n9613), .B1(n13359), .B2(n9615), .C1(
        n9695), .C2(P2_U3088), .ZN(P2_U3322) );
  OAI222_X1 U12095 ( .A1(P1_U3086), .A2(n10133), .B1(n10724), .B2(n9615), .C1(
        n9614), .C2(n14039), .ZN(P1_U3350) );
  INV_X1 U12096 ( .A(n12787), .ZN(n9882) );
  AOI222_X1 U12097 ( .A1(n9616), .A2(n12775), .B1(SI_4_), .B2(n9882), .C1(
        P3_STATE_REG_SCAN_IN), .C2(n10795), .ZN(n9617) );
  INV_X1 U12098 ( .A(n9617), .ZN(P3_U3291) );
  AOI222_X1 U12099 ( .A1(n9618), .A2(n12775), .B1(SI_9_), .B2(n9882), .C1(
        P3_STATE_REG_SCAN_IN), .C2(n12460), .ZN(n9619) );
  INV_X1 U12100 ( .A(n9619), .ZN(P3_U3286) );
  AOI222_X1 U12101 ( .A1(n9620), .A2(n12775), .B1(n9882), .B2(SI_2_), .C1(
        n9967), .C2(P3_STATE_REG_SCAN_IN), .ZN(n9621) );
  INV_X1 U12102 ( .A(n9621), .ZN(P3_U3293) );
  AOI222_X1 U12103 ( .A1(n9622), .A2(n12775), .B1(SI_7_), .B2(n9882), .C1(
        P3_STATE_REG_SCAN_IN), .C2(n14993), .ZN(n9623) );
  INV_X1 U12104 ( .A(n9623), .ZN(P3_U3288) );
  AOI222_X1 U12105 ( .A1(n9624), .A2(n12775), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n14956), .C1(SI_3_), .C2(n9882), .ZN(n9625) );
  INV_X1 U12106 ( .A(n9625), .ZN(P3_U3292) );
  AOI222_X1 U12107 ( .A1(n9626), .A2(n12775), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n14962), .C1(SI_5_), .C2(n9882), .ZN(n9627) );
  INV_X1 U12108 ( .A(n9627), .ZN(P3_U3290) );
  INV_X1 U12109 ( .A(n9628), .ZN(n9629) );
  INV_X1 U12110 ( .A(n12466), .ZN(n15063) );
  OAI222_X1 U12111 ( .A1(n12785), .A2(n9629), .B1(n15063), .B2(P3_U3151), .C1(
        n15490), .C2(n12787), .ZN(P3_U3283) );
  INV_X1 U12112 ( .A(n9769), .ZN(n14726) );
  OAI222_X1 U12113 ( .A1(n13357), .A2(n9630), .B1(n13359), .B2(n9632), .C1(
        n14726), .C2(P2_U3088), .ZN(P2_U3321) );
  INV_X1 U12114 ( .A(n10183), .ZN(n9633) );
  OAI222_X1 U12115 ( .A1(P1_U3086), .A2(n9633), .B1(n10724), .B2(n9632), .C1(
        n9631), .C2(n14039), .ZN(P1_U3349) );
  INV_X1 U12116 ( .A(n12951), .ZN(n9634) );
  OAI222_X1 U12117 ( .A1(n13357), .A2(n9635), .B1(n13359), .B2(n9637), .C1(
        n9634), .C2(P2_U3088), .ZN(P2_U3320) );
  INV_X1 U12118 ( .A(n10171), .ZN(n9638) );
  OAI222_X1 U12119 ( .A1(P1_U3086), .A2(n9638), .B1(n10724), .B2(n9637), .C1(
        n9636), .C2(n14039), .ZN(P1_U3348) );
  AOI222_X1 U12120 ( .A1(n9639), .A2(n12775), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15074), .C1(SI_13_), .C2(n9882), .ZN(n9640) );
  INV_X1 U12121 ( .A(n9640), .ZN(P3_U3282) );
  NAND2_X1 U12122 ( .A1(n9816), .A2(n11309), .ZN(n9641) );
  NAND2_X1 U12123 ( .A1(n9642), .A2(n9641), .ZN(n9646) );
  INV_X1 U12124 ( .A(n9643), .ZN(n9644) );
  NAND2_X1 U12125 ( .A1(n9644), .A2(n11309), .ZN(n9645) );
  NAND2_X1 U12126 ( .A1(n9646), .A2(n9645), .ZN(n9658) );
  NAND2_X1 U12127 ( .A1(n9658), .A2(n8287), .ZN(n14696) );
  INV_X1 U12128 ( .A(n14817), .ZN(n14825) );
  OR2_X1 U12129 ( .A1(n8287), .A2(P2_U3088), .ZN(n13352) );
  INV_X1 U12130 ( .A(n8288), .ZN(n12103) );
  NOR2_X1 U12131 ( .A1(n13352), .A2(n12103), .ZN(n9647) );
  NAND2_X1 U12132 ( .A1(n9658), .A2(n9647), .ZN(n14819) );
  INV_X1 U12133 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n15310) );
  MUX2_X1 U12134 ( .A(n15310), .B(P2_REG1_REG_4__SCAN_IN), .S(n9687), .Z(n9655) );
  XNOR2_X1 U12135 ( .A(n14714), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n14708) );
  XNOR2_X1 U12136 ( .A(n9659), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n14694) );
  AND2_X1 U12137 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n14693) );
  NAND2_X1 U12138 ( .A1(n14694), .A2(n14693), .ZN(n9649) );
  NAND2_X1 U12139 ( .A1(n9661), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9648) );
  NAND2_X1 U12140 ( .A1(n9649), .A2(n9648), .ZN(n14707) );
  NAND2_X1 U12141 ( .A1(n14708), .A2(n14707), .ZN(n14706) );
  INV_X1 U12142 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9650) );
  OR2_X1 U12143 ( .A1(n14714), .A2(n9650), .ZN(n9651) );
  NAND2_X1 U12144 ( .A1(n14706), .A2(n9651), .ZN(n9676) );
  XNOR2_X1 U12145 ( .A(n9686), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n9677) );
  NAND2_X1 U12146 ( .A1(n9676), .A2(n9677), .ZN(n9675) );
  INV_X1 U12147 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9652) );
  OR2_X1 U12148 ( .A1(n9686), .A2(n9652), .ZN(n9653) );
  NAND2_X1 U12149 ( .A1(n9675), .A2(n9653), .ZN(n9654) );
  NAND2_X1 U12150 ( .A1(n9654), .A2(n9655), .ZN(n9689) );
  OAI21_X1 U12151 ( .B1(n9655), .B2(n9654), .A(n9689), .ZN(n9656) );
  NAND2_X1 U12152 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n10110) );
  OAI21_X1 U12153 ( .B1(n14819), .B2(n9656), .A(n10110), .ZN(n9673) );
  NOR2_X1 U12154 ( .A1(n13352), .A2(n8288), .ZN(n9657) );
  INV_X1 U12155 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9663) );
  MUX2_X1 U12156 ( .A(n9663), .B(P2_REG2_REG_2__SCAN_IN), .S(n14714), .Z(
        n14717) );
  INV_X1 U12157 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9660) );
  MUX2_X1 U12158 ( .A(n9660), .B(P2_REG2_REG_1__SCAN_IN), .S(n9659), .Z(n14701) );
  AND2_X1 U12159 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n14702) );
  NAND2_X1 U12160 ( .A1(n14701), .A2(n14702), .ZN(n14700) );
  NAND2_X1 U12161 ( .A1(n9661), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9662) );
  NAND2_X1 U12162 ( .A1(n14700), .A2(n9662), .ZN(n14718) );
  NAND2_X1 U12163 ( .A1(n14717), .A2(n14718), .ZN(n14716) );
  OR2_X1 U12164 ( .A1(n14714), .A2(n9663), .ZN(n9679) );
  NAND2_X1 U12165 ( .A1(n14716), .A2(n9679), .ZN(n9665) );
  INV_X1 U12166 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10272) );
  MUX2_X1 U12167 ( .A(n10272), .B(P2_REG2_REG_3__SCAN_IN), .S(n9686), .Z(n9664) );
  NAND2_X1 U12168 ( .A1(n9665), .A2(n9664), .ZN(n9682) );
  OR2_X1 U12169 ( .A1(n9686), .A2(n10272), .ZN(n9670) );
  NAND2_X1 U12170 ( .A1(n9682), .A2(n9670), .ZN(n9668) );
  INV_X1 U12171 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n9666) );
  MUX2_X1 U12172 ( .A(n9666), .B(P2_REG2_REG_4__SCAN_IN), .S(n9687), .Z(n9667)
         );
  NAND2_X1 U12173 ( .A1(n9668), .A2(n9667), .ZN(n9698) );
  MUX2_X1 U12174 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n9666), .S(n9687), .Z(n9669)
         );
  NAND3_X1 U12175 ( .A1(n9682), .A2(n9670), .A3(n9669), .ZN(n9671) );
  AND3_X1 U12176 ( .A1(n14811), .A2(n9698), .A3(n9671), .ZN(n9672) );
  AOI211_X1 U12177 ( .C1(n14825), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n9673), .B(
        n9672), .ZN(n9674) );
  OAI21_X1 U12178 ( .B1(n9687), .B2(n14833), .A(n9674), .ZN(P2_U3218) );
  OAI21_X1 U12179 ( .B1(n9677), .B2(n9676), .A(n9675), .ZN(n9678) );
  OAI22_X1 U12180 ( .A1(n14819), .A2(n9678), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10270), .ZN(n9684) );
  MUX2_X1 U12181 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10272), .S(n9686), .Z(n9680) );
  NAND3_X1 U12182 ( .A1(n14716), .A2(n9680), .A3(n9679), .ZN(n9681) );
  AND3_X1 U12183 ( .A1(n14811), .A2(n9682), .A3(n9681), .ZN(n9683) );
  AOI211_X1 U12184 ( .C1(n14825), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n9684), .B(
        n9683), .ZN(n9685) );
  OAI21_X1 U12185 ( .B1(n9686), .B2(n14833), .A(n9685), .ZN(P2_U3217) );
  XNOR2_X1 U12186 ( .A(n9695), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n9691) );
  INV_X1 U12187 ( .A(n9687), .ZN(n9692) );
  NAND2_X1 U12188 ( .A1(n9692), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9688) );
  NAND2_X1 U12189 ( .A1(n9689), .A2(n9688), .ZN(n9690) );
  NAND2_X1 U12190 ( .A1(n9690), .A2(n9691), .ZN(n9755) );
  OAI21_X1 U12191 ( .B1(n9691), .B2(n9690), .A(n9755), .ZN(n9703) );
  INV_X1 U12192 ( .A(n14833), .ZN(n14809) );
  NOR2_X1 U12193 ( .A1(n7794), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10257) );
  NAND2_X1 U12194 ( .A1(n9692), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9697) );
  NAND2_X1 U12195 ( .A1(n9698), .A2(n9697), .ZN(n9694) );
  INV_X1 U12196 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10402) );
  MUX2_X1 U12197 ( .A(n10402), .B(P2_REG2_REG_5__SCAN_IN), .S(n9695), .Z(n9693) );
  NAND2_X1 U12198 ( .A1(n9694), .A2(n9693), .ZN(n9768) );
  MUX2_X1 U12199 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10402), .S(n9695), .Z(n9696) );
  NAND3_X1 U12200 ( .A1(n9698), .A2(n9697), .A3(n9696), .ZN(n9699) );
  AND3_X1 U12201 ( .A1(n14811), .A2(n9768), .A3(n9699), .ZN(n9700) );
  AOI211_X1 U12202 ( .C1(n14809), .C2(n9766), .A(n10257), .B(n9700), .ZN(n9702) );
  NAND2_X1 U12203 ( .A1(n14825), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n9701) );
  OAI211_X1 U12204 ( .C1(n14819), .C2(n9703), .A(n9702), .B(n9701), .ZN(
        P2_U3219) );
  INV_X1 U12205 ( .A(n14740), .ZN(n9704) );
  OAI222_X1 U12206 ( .A1(n13357), .A2(n9705), .B1(n13359), .B2(n9707), .C1(
        n9704), .C2(P2_U3088), .ZN(P2_U3319) );
  INV_X1 U12207 ( .A(n10222), .ZN(n9708) );
  OAI222_X1 U12208 ( .A1(P1_U3086), .A2(n9708), .B1(n10724), .B2(n9707), .C1(
        n9706), .C2(n14039), .ZN(P1_U3347) );
  NOR2_X1 U12209 ( .A1(n12773), .A2(n9709), .ZN(n9719) );
  CLKBUF_X1 U12210 ( .A(n9719), .Z(n9737) );
  INV_X1 U12211 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n9710) );
  NOR2_X1 U12212 ( .A1(n9737), .A2(n9710), .ZN(P3_U3251) );
  INV_X1 U12213 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n15444) );
  NOR2_X1 U12214 ( .A1(n9737), .A2(n15444), .ZN(P3_U3248) );
  INV_X1 U12215 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n9711) );
  NOR2_X1 U12216 ( .A1(n9737), .A2(n9711), .ZN(P3_U3247) );
  INV_X1 U12217 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n9712) );
  NOR2_X1 U12218 ( .A1(n9737), .A2(n9712), .ZN(P3_U3250) );
  INV_X1 U12219 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n9713) );
  NOR2_X1 U12220 ( .A1(n9737), .A2(n9713), .ZN(P3_U3249) );
  INV_X1 U12221 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n9714) );
  NOR2_X1 U12222 ( .A1(n9737), .A2(n9714), .ZN(P3_U3256) );
  INV_X1 U12223 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n9715) );
  NOR2_X1 U12224 ( .A1(n9737), .A2(n9715), .ZN(P3_U3255) );
  INV_X1 U12225 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n9716) );
  NOR2_X1 U12226 ( .A1(n9737), .A2(n9716), .ZN(P3_U3253) );
  INV_X1 U12227 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n9717) );
  NOR2_X1 U12228 ( .A1(n9737), .A2(n9717), .ZN(P3_U3252) );
  INV_X1 U12229 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n9718) );
  NOR2_X1 U12230 ( .A1(n9737), .A2(n9718), .ZN(P3_U3259) );
  INV_X1 U12231 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n9720) );
  NOR2_X1 U12232 ( .A1(n9737), .A2(n9720), .ZN(P3_U3260) );
  INV_X1 U12233 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n9721) );
  NOR2_X1 U12234 ( .A1(n9737), .A2(n9721), .ZN(P3_U3261) );
  INV_X1 U12235 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n9722) );
  NOR2_X1 U12236 ( .A1(n9719), .A2(n9722), .ZN(P3_U3262) );
  INV_X1 U12237 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n9723) );
  NOR2_X1 U12238 ( .A1(n9737), .A2(n9723), .ZN(P3_U3263) );
  INV_X1 U12239 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n9724) );
  NOR2_X1 U12240 ( .A1(n9737), .A2(n9724), .ZN(P3_U3246) );
  INV_X1 U12241 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n9725) );
  NOR2_X1 U12242 ( .A1(n9719), .A2(n9725), .ZN(P3_U3245) );
  INV_X1 U12243 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n9726) );
  NOR2_X1 U12244 ( .A1(n9719), .A2(n9726), .ZN(P3_U3244) );
  INV_X1 U12245 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n9727) );
  NOR2_X1 U12246 ( .A1(n9719), .A2(n9727), .ZN(P3_U3243) );
  INV_X1 U12247 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n9728) );
  NOR2_X1 U12248 ( .A1(n9719), .A2(n9728), .ZN(P3_U3242) );
  INV_X1 U12249 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n9729) );
  NOR2_X1 U12250 ( .A1(n9719), .A2(n9729), .ZN(P3_U3241) );
  INV_X1 U12251 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n15466) );
  NOR2_X1 U12252 ( .A1(n9719), .A2(n15466), .ZN(P3_U3240) );
  INV_X1 U12253 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n9730) );
  NOR2_X1 U12254 ( .A1(n9719), .A2(n9730), .ZN(P3_U3239) );
  INV_X1 U12255 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n9731) );
  NOR2_X1 U12256 ( .A1(n9719), .A2(n9731), .ZN(P3_U3238) );
  INV_X1 U12257 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n15349) );
  NOR2_X1 U12258 ( .A1(n9719), .A2(n15349), .ZN(P3_U3237) );
  INV_X1 U12259 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n9732) );
  NOR2_X1 U12260 ( .A1(n9719), .A2(n9732), .ZN(P3_U3236) );
  INV_X1 U12261 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n9733) );
  NOR2_X1 U12262 ( .A1(n9737), .A2(n9733), .ZN(P3_U3235) );
  INV_X1 U12263 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n9734) );
  NOR2_X1 U12264 ( .A1(n9737), .A2(n9734), .ZN(P3_U3234) );
  INV_X1 U12265 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n9735) );
  NOR2_X1 U12266 ( .A1(n9737), .A2(n9735), .ZN(P3_U3257) );
  INV_X1 U12267 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n15404) );
  NOR2_X1 U12268 ( .A1(n9737), .A2(n15404), .ZN(P3_U3258) );
  INV_X1 U12269 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n9736) );
  NOR2_X1 U12270 ( .A1(n9737), .A2(n9736), .ZN(P3_U3254) );
  OAI222_X1 U12271 ( .A1(n12785), .A2(n9739), .B1(n12787), .B2(n9738), .C1(
        n15100), .C2(P3_U3151), .ZN(P3_U3281) );
  INV_X1 U12272 ( .A(n10208), .ZN(n9741) );
  OAI222_X1 U12273 ( .A1(P1_U3086), .A2(n9741), .B1(n10724), .B2(n9742), .C1(
        n9740), .C2(n14039), .ZN(P1_U3346) );
  INV_X1 U12274 ( .A(n9776), .ZN(n14755) );
  OAI222_X1 U12275 ( .A1(n13357), .A2(n9743), .B1(n13359), .B2(n9742), .C1(
        n14755), .C2(P2_U3088), .ZN(P2_U3318) );
  NAND2_X1 U12276 ( .A1(n11463), .A2(P1_B_REG_SCAN_IN), .ZN(n9744) );
  MUX2_X1 U12277 ( .A(n9744), .B(P1_B_REG_SCAN_IN), .S(n11331), .Z(n9745) );
  NOR2_X1 U12278 ( .A1(n14038), .A2(P1_U3086), .ZN(n9746) );
  NAND2_X1 U12279 ( .A1(n9793), .A2(n9746), .ZN(n9748) );
  OAI22_X1 U12280 ( .A1(n14606), .A2(P1_D_REG_0__SCAN_IN), .B1(n11331), .B2(
        n9748), .ZN(n9747) );
  INV_X1 U12281 ( .A(n9747), .ZN(P1_U3445) );
  OAI22_X1 U12282 ( .A1(n14606), .A2(P1_D_REG_1__SCAN_IN), .B1(n9992), .B2(
        n9748), .ZN(n9749) );
  INV_X1 U12283 ( .A(n9749), .ZN(P1_U3446) );
  INV_X1 U12284 ( .A(n9750), .ZN(n9752) );
  INV_X1 U12285 ( .A(n12473), .ZN(n14198) );
  OAI222_X1 U12286 ( .A1(n12785), .A2(n9752), .B1(n12787), .B2(n9751), .C1(
        n14198), .C2(P3_U3151), .ZN(P3_U3280) );
  INV_X1 U12287 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9753) );
  MUX2_X1 U12288 ( .A(n9753), .B(P2_REG1_REG_10__SCAN_IN), .S(n10069), .Z(
        n9765) );
  NAND2_X1 U12289 ( .A1(n9766), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9754) );
  NAND2_X1 U12290 ( .A1(n9755), .A2(n9754), .ZN(n14722) );
  INV_X1 U12291 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9756) );
  MUX2_X1 U12292 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n9756), .S(n9769), .Z(n14723) );
  NAND2_X1 U12293 ( .A1(n14722), .A2(n14723), .ZN(n14721) );
  NAND2_X1 U12294 ( .A1(n9769), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9757) );
  NAND2_X1 U12295 ( .A1(n14721), .A2(n9757), .ZN(n12949) );
  INV_X1 U12296 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9758) );
  MUX2_X1 U12297 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n9758), .S(n12951), .Z(
        n12950) );
  NAND2_X1 U12298 ( .A1(n12949), .A2(n12950), .ZN(n12948) );
  NAND2_X1 U12299 ( .A1(n12951), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9759) );
  NAND2_X1 U12300 ( .A1(n12948), .A2(n9759), .ZN(n14736) );
  INV_X1 U12301 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n14930) );
  MUX2_X1 U12302 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n14930), .S(n14740), .Z(
        n14735) );
  NAND2_X1 U12303 ( .A1(n14736), .A2(n14735), .ZN(n14734) );
  NAND2_X1 U12304 ( .A1(n14740), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9760) );
  NAND2_X1 U12305 ( .A1(n14734), .A2(n9760), .ZN(n14748) );
  INV_X1 U12306 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9761) );
  MUX2_X1 U12307 ( .A(n9761), .B(P2_REG1_REG_9__SCAN_IN), .S(n9776), .Z(n14747) );
  OR2_X1 U12308 ( .A1(n14748), .A2(n14747), .ZN(n14750) );
  NAND2_X1 U12309 ( .A1(n14755), .A2(n9761), .ZN(n9762) );
  NAND2_X1 U12310 ( .A1(n14750), .A2(n9762), .ZN(n9764) );
  OR2_X1 U12311 ( .A1(n9764), .A2(n9765), .ZN(n10071) );
  INV_X1 U12312 ( .A(n10071), .ZN(n9763) );
  AOI211_X1 U12313 ( .C1(n9765), .C2(n9764), .A(n14819), .B(n9763), .ZN(n9786)
         );
  NAND2_X1 U12314 ( .A1(n9766), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9767) );
  NAND2_X1 U12315 ( .A1(n9768), .A2(n9767), .ZN(n14730) );
  INV_X1 U12316 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10605) );
  MUX2_X1 U12317 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10605), .S(n9769), .Z(
        n14729) );
  NAND2_X1 U12318 ( .A1(n14730), .A2(n14729), .ZN(n14728) );
  NAND2_X1 U12319 ( .A1(n9769), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n12953) );
  NAND2_X1 U12320 ( .A1(n14728), .A2(n12953), .ZN(n9772) );
  INV_X1 U12321 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n9770) );
  MUX2_X1 U12322 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n9770), .S(n12951), .Z(n9771) );
  NAND2_X1 U12323 ( .A1(n9772), .A2(n9771), .ZN(n12955) );
  NAND2_X1 U12324 ( .A1(n12951), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9773) );
  NAND2_X1 U12325 ( .A1(n12955), .A2(n9773), .ZN(n14743) );
  INV_X1 U12326 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n9774) );
  MUX2_X1 U12327 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n9774), .S(n14740), .Z(
        n14742) );
  NAND2_X1 U12328 ( .A1(n14743), .A2(n14742), .ZN(n14741) );
  NAND2_X1 U12329 ( .A1(n14740), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9775) );
  NAND2_X1 U12330 ( .A1(n14741), .A2(n9775), .ZN(n14752) );
  INV_X1 U12331 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n9777) );
  MUX2_X1 U12332 ( .A(n9777), .B(P2_REG2_REG_9__SCAN_IN), .S(n9776), .Z(n14751) );
  OR2_X1 U12333 ( .A1(n14752), .A2(n14751), .ZN(n14754) );
  NAND2_X1 U12334 ( .A1(n14755), .A2(n9777), .ZN(n9778) );
  NAND2_X1 U12335 ( .A1(n14754), .A2(n9778), .ZN(n9782) );
  INV_X1 U12336 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n9779) );
  MUX2_X1 U12337 ( .A(n9779), .B(P2_REG2_REG_10__SCAN_IN), .S(n10069), .Z(
        n9781) );
  INV_X1 U12338 ( .A(n14811), .ZN(n14829) );
  OR2_X1 U12339 ( .A1(n9782), .A2(n9781), .ZN(n10062) );
  INV_X1 U12340 ( .A(n10062), .ZN(n9780) );
  AOI211_X1 U12341 ( .C1(n9782), .C2(n9781), .A(n14829), .B(n9780), .ZN(n9785)
         );
  INV_X1 U12342 ( .A(n10069), .ZN(n9790) );
  AND2_X1 U12343 ( .A1(P2_U3088), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n10856) );
  AOI21_X1 U12344 ( .B1(n14825), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n10856), 
        .ZN(n9783) );
  OAI21_X1 U12345 ( .B1(n9790), .B2(n14833), .A(n9783), .ZN(n9784) );
  OR3_X1 U12346 ( .A1(n9786), .A2(n9785), .A3(n9784), .ZN(P2_U3224) );
  NAND2_X1 U12347 ( .A1(n12410), .A2(P3_DATAO_REG_13__SCAN_IN), .ZN(n9787) );
  OAI21_X1 U12348 ( .B1(n11483), .B2(n12410), .A(n9787), .ZN(P3_U3504) );
  INV_X1 U12349 ( .A(n10424), .ZN(n9789) );
  OAI222_X1 U12350 ( .A1(P1_U3086), .A2(n9789), .B1(n10724), .B2(n9791), .C1(
        n9788), .C2(n14039), .ZN(P1_U3345) );
  OAI222_X1 U12351 ( .A1(n13357), .A2(n9792), .B1(n13359), .B2(n9791), .C1(
        n9790), .C2(P2_U3088), .ZN(P2_U3317) );
  OR2_X1 U12352 ( .A1(n9559), .A2(n10871), .ZN(n9799) );
  NAND2_X1 U12353 ( .A1(n10023), .A2(n9793), .ZN(n9794) );
  NAND2_X1 U12354 ( .A1(n9794), .A2(n9043), .ZN(n9797) );
  INV_X1 U12355 ( .A(n14529), .ZN(n10418) );
  NOR2_X1 U12356 ( .A1(n10418), .A2(P1_U4016), .ZN(P1_U3085) );
  AOI222_X1 U12357 ( .A1(n9795), .A2(n12775), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12447), .C1(SI_16_), .C2(n9882), .ZN(n9796) );
  INV_X1 U12358 ( .A(n9796), .ZN(P3_U3279) );
  INV_X1 U12359 ( .A(n9797), .ZN(n9798) );
  AND2_X1 U12360 ( .A1(n9799), .A2(n9798), .ZN(n10139) );
  INV_X1 U12361 ( .A(n6641), .ZN(n9801) );
  INV_X1 U12362 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9800) );
  AOI21_X1 U12363 ( .B1(n9801), .B2(n9800), .A(n9571), .ZN(n13617) );
  OAI21_X1 U12364 ( .B1(n9801), .B2(P1_REG1_REG_0__SCAN_IN), .A(n13617), .ZN(
        n9802) );
  XNOR2_X1 U12365 ( .A(n9802), .B(n14044), .ZN(n9803) );
  AOI22_X1 U12366 ( .A1(n10139), .A2(n9803), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n9804) );
  OAI21_X1 U12367 ( .B1(n14529), .B2(n7546), .A(n9804), .ZN(P1_U3243) );
  NAND2_X1 U12368 ( .A1(n9806), .A2(n9805), .ZN(n9811) );
  INV_X1 U12369 ( .A(n9813), .ZN(n9807) );
  OAI21_X1 U12370 ( .B1(n9811), .B2(n9808), .A(n9807), .ZN(n9810) );
  NAND2_X1 U12371 ( .A1(n9810), .A2(n9809), .ZN(n9931) );
  INV_X1 U12372 ( .A(n14881), .ZN(n14879) );
  NOR2_X1 U12373 ( .A1(n9931), .A2(n14879), .ZN(n9907) );
  INV_X1 U12374 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10196) );
  NAND2_X1 U12375 ( .A1(n14881), .A2(n10190), .ZN(n14877) );
  NOR2_X1 U12376 ( .A1(n9811), .A2(n14877), .ZN(n9819) );
  NOR2_X1 U12377 ( .A1(n9812), .A2(n12066), .ZN(n10199) );
  NAND2_X1 U12378 ( .A1(n9819), .A2(n10199), .ZN(n9814) );
  INV_X1 U12379 ( .A(n12900), .ZN(n12913) );
  AND2_X1 U12380 ( .A1(n9819), .A2(n12102), .ZN(n12897) );
  INV_X1 U12381 ( .A(n12902), .ZN(n12891) );
  NOR2_X1 U12382 ( .A1(n9815), .A2(n12891), .ZN(n10193) );
  AOI22_X1 U12383 ( .A1(n12913), .A2(n14882), .B1(n12897), .B2(n10193), .ZN(
        n9823) );
  NAND2_X1 U12384 ( .A1(n14882), .A2(n14313), .ZN(n9871) );
  NAND2_X1 U12385 ( .A1(n11843), .A2(n7214), .ZN(n11846) );
  NOR2_X1 U12386 ( .A1(n11846), .A2(n14313), .ZN(n9820) );
  INV_X1 U12387 ( .A(n9816), .ZN(n9817) );
  AND2_X1 U12388 ( .A1(n9817), .A2(n14915), .ZN(n9818) );
  OAI21_X1 U12389 ( .B1(n9821), .B2(n9820), .A(n12887), .ZN(n9822) );
  OAI211_X1 U12390 ( .C1(n9907), .C2(n10196), .A(n9823), .B(n9822), .ZN(
        P2_U3204) );
  NAND2_X1 U12391 ( .A1(P3_U3897), .A2(n11819), .ZN(n15082) );
  INV_X4 U12392 ( .A(n11753), .ZN(n12452) );
  MUX2_X1 U12393 ( .A(P3_REG2_REG_0__SCAN_IN), .B(P3_REG1_REG_0__SCAN_IN), .S(
        n8943), .Z(n14939) );
  NOR2_X1 U12394 ( .A1(n14939), .A2(n6827), .ZN(n14937) );
  MUX2_X1 U12395 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n8943), .Z(n9846) );
  XOR2_X1 U12396 ( .A(n9836), .B(n9846), .Z(n9849) );
  XOR2_X1 U12397 ( .A(n14937), .B(n9849), .Z(n9845) );
  INV_X1 U12398 ( .A(n9836), .ZN(n9848) );
  NAND2_X1 U12399 ( .A1(n11711), .A2(n9939), .ZN(n9824) );
  AND2_X1 U12400 ( .A1(n9825), .A2(n9824), .ZN(n9827) );
  OR2_X1 U12401 ( .A1(n9939), .A2(P3_U3151), .ZN(n11759) );
  NAND2_X1 U12402 ( .A1(n11755), .A2(n11759), .ZN(n9828) );
  MUX2_X1 U12403 ( .A(n9835), .B(P3_U3897), .S(n9826), .Z(n15016) );
  INV_X1 U12404 ( .A(n9827), .ZN(n9829) );
  AOI22_X1 U12405 ( .A1(n15025), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n9842) );
  INV_X1 U12406 ( .A(n15095), .ZN(n14966) );
  INV_X1 U12407 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10055) );
  NAND2_X1 U12408 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n14936), .ZN(n9830) );
  NAND2_X1 U12409 ( .A1(n9831), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n9853) );
  OAI21_X1 U12410 ( .B1(n9831), .B2(P3_REG1_REG_1__SCAN_IN), .A(n9853), .ZN(
        n9832) );
  NAND2_X1 U12411 ( .A1(n14966), .A2(n9832), .ZN(n9841) );
  INV_X1 U12412 ( .A(n9833), .ZN(n9834) );
  INV_X1 U12413 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n15429) );
  NOR2_X1 U12414 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n15429), .ZN(n14935) );
  OAI21_X1 U12415 ( .B1(n9836), .B2(n14935), .A(n7687), .ZN(n9837) );
  INV_X1 U12416 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n15130) );
  OR2_X1 U12417 ( .A1(n9837), .A2(n15130), .ZN(n9859) );
  NAND2_X1 U12418 ( .A1(n9837), .A2(n15130), .ZN(n9838) );
  NAND2_X1 U12419 ( .A1(n9859), .A2(n9838), .ZN(n9839) );
  NAND2_X1 U12420 ( .A1(n14998), .A2(n9839), .ZN(n9840) );
  NAND3_X1 U12421 ( .A1(n9842), .A2(n9841), .A3(n9840), .ZN(n9843) );
  AOI21_X1 U12422 ( .B1(n9848), .B2(n15016), .A(n9843), .ZN(n9844) );
  OAI21_X1 U12423 ( .B1(n15082), .B2(n9845), .A(n9844), .ZN(P3_U3183) );
  MUX2_X1 U12424 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n12452), .Z(n9968) );
  XOR2_X1 U12425 ( .A(n9967), .B(n9968), .Z(n9969) );
  INV_X1 U12426 ( .A(n9846), .ZN(n9847) );
  AOI22_X1 U12427 ( .A1(n9849), .A2(n14937), .B1(n9848), .B2(n9847), .ZN(n9970) );
  XOR2_X1 U12428 ( .A(n9969), .B(n9970), .Z(n9869) );
  AOI22_X1 U12429 ( .A1(n15025), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n9866) );
  INV_X1 U12430 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n15186) );
  OR2_X1 U12431 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n9851), .ZN(n9852) );
  OAI21_X1 U12432 ( .B1(n9856), .B2(n9855), .A(n9854), .ZN(n9857) );
  NAND2_X1 U12433 ( .A1(n14966), .A2(n9857), .ZN(n9865) );
  OAI21_X1 U12434 ( .B1(n9967), .B2(P3_REG2_REG_2__SCAN_IN), .A(n9858), .ZN(
        n9862) );
  NAND2_X1 U12435 ( .A1(n9859), .A2(n7687), .ZN(n9861) );
  INV_X1 U12436 ( .A(n9979), .ZN(n9860) );
  OAI21_X1 U12437 ( .B1(n9862), .B2(n9861), .A(n9860), .ZN(n9863) );
  NAND2_X1 U12438 ( .A1(n14998), .A2(n9863), .ZN(n9864) );
  NAND3_X1 U12439 ( .A1(n9866), .A2(n9865), .A3(n9864), .ZN(n9867) );
  AOI21_X1 U12440 ( .B1(n9967), .B2(n15016), .A(n9867), .ZN(n9868) );
  OAI21_X1 U12441 ( .B1(n9869), .B2(n15082), .A(n9868), .ZN(P3_U3184) );
  INV_X1 U12442 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n9881) );
  XNOR2_X1 U12443 ( .A(n11854), .B(n10532), .ZN(n9895) );
  NAND2_X1 U12444 ( .A1(n12944), .A2(n11181), .ZN(n9896) );
  XNOR2_X1 U12445 ( .A(n9895), .B(n9896), .ZN(n9875) );
  OR2_X1 U12446 ( .A1(n14882), .A2(n9889), .ZN(n9872) );
  AND2_X1 U12447 ( .A1(n9872), .A2(n9871), .ZN(n9873) );
  NAND2_X1 U12448 ( .A1(n9874), .A2(n9875), .ZN(n9899) );
  OAI21_X1 U12449 ( .B1(n9875), .B2(n9874), .A(n9899), .ZN(n9876) );
  NAND2_X1 U12450 ( .A1(n9876), .A2(n12887), .ZN(n9880) );
  OAI22_X1 U12451 ( .A1(n9878), .A2(n12889), .B1(n9877), .B2(n12891), .ZN(
        n9918) );
  AOI22_X1 U12452 ( .A1(n12913), .A2(n9920), .B1(n9918), .B2(n12897), .ZN(
        n9879) );
  OAI211_X1 U12453 ( .C1(n9907), .C2(n9881), .A(n9880), .B(n9879), .ZN(
        P2_U3194) );
  AOI222_X1 U12454 ( .A1(n9883), .A2(n12775), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12478), .C1(SI_17_), .C2(n9882), .ZN(n9884) );
  INV_X1 U12455 ( .A(n9884), .ZN(P3_U3278) );
  INV_X1 U12456 ( .A(n9885), .ZN(n9887) );
  INV_X1 U12457 ( .A(n10426), .ZN(n14431) );
  OAI222_X1 U12458 ( .A1(n14039), .A2(n9886), .B1(n10724), .B2(n9887), .C1(
        P1_U3086), .C2(n14431), .ZN(P1_U3344) );
  INV_X1 U12459 ( .A(n10073), .ZN(n14771) );
  OAI222_X1 U12460 ( .A1(n13357), .A2(n9888), .B1(n13359), .B2(n9887), .C1(
        P2_U3088), .C2(n14771), .ZN(P2_U3316) );
  INV_X1 U12461 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n14709) );
  XNOR2_X1 U12462 ( .A(n11851), .B(n9889), .ZN(n9890) );
  NAND2_X1 U12463 ( .A1(n12943), .A2(n12126), .ZN(n9891) );
  NAND2_X1 U12464 ( .A1(n9890), .A2(n9891), .ZN(n9925) );
  INV_X1 U12465 ( .A(n9890), .ZN(n9893) );
  INV_X1 U12466 ( .A(n9891), .ZN(n9892) );
  NAND2_X1 U12467 ( .A1(n9893), .A2(n9892), .ZN(n9894) );
  AND2_X1 U12468 ( .A1(n9925), .A2(n9894), .ZN(n9901) );
  INV_X1 U12469 ( .A(n9895), .ZN(n9897) );
  NAND2_X1 U12470 ( .A1(n9897), .A2(n9896), .ZN(n9898) );
  NAND2_X1 U12471 ( .A1(n9899), .A2(n9898), .ZN(n9900) );
  OAI21_X1 U12472 ( .B1(n9901), .B2(n9900), .A(n9926), .ZN(n9902) );
  NAND2_X1 U12473 ( .A1(n9902), .A2(n12887), .ZN(n9906) );
  NAND2_X1 U12474 ( .A1(n12942), .A2(n12902), .ZN(n9904) );
  NAND2_X1 U12475 ( .A1(n12944), .A2(n12901), .ZN(n9903) );
  NAND2_X1 U12476 ( .A1(n9904), .A2(n9903), .ZN(n10046) );
  AOI22_X1 U12477 ( .A1(n12913), .A2(n11851), .B1(n12897), .B2(n10046), .ZN(
        n9905) );
  OAI211_X1 U12478 ( .C1(n9907), .C2(n14709), .A(n9906), .B(n9905), .ZN(
        P2_U3209) );
  INV_X1 U12479 ( .A(n12411), .ZN(n15120) );
  NOR2_X1 U12480 ( .A1(n15120), .A2(n10286), .ZN(n11560) );
  NOR2_X1 U12481 ( .A1(n11560), .A2(n15113), .ZN(n11722) );
  INV_X1 U12482 ( .A(n11754), .ZN(n9946) );
  NOR3_X1 U12483 ( .A1(n11722), .A2(n9946), .A3(n15157), .ZN(n9909) );
  AOI21_X1 U12484 ( .B1(n12375), .B2(n12409), .A(n9909), .ZN(n10284) );
  INV_X1 U12485 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n9910) );
  OAI22_X1 U12486 ( .A1(n10056), .A2(n12771), .B1(n15181), .B2(n9910), .ZN(
        n9911) );
  INV_X1 U12487 ( .A(n9911), .ZN(n9912) );
  OAI21_X1 U12488 ( .B1(n10284), .B2(n15183), .A(n9912), .ZN(P3_U3390) );
  INV_X1 U12489 ( .A(n9913), .ZN(n9914) );
  OAI222_X1 U12490 ( .A1(n12785), .A2(n9914), .B1(n12787), .B2(n15288), .C1(
        n14243), .C2(P3_U3151), .ZN(P3_U3277) );
  XOR2_X1 U12491 ( .A(n9915), .B(n12067), .Z(n10496) );
  AOI21_X1 U12492 ( .B1(n9870), .B2(n9916), .A(n10496), .ZN(n9923) );
  XNOR2_X1 U12493 ( .A(n9917), .B(n12067), .ZN(n9919) );
  AOI21_X1 U12494 ( .B1(n9919), .B2(n14304), .A(n9918), .ZN(n10503) );
  NAND2_X1 U12495 ( .A1(n9920), .A2(n14882), .ZN(n9921) );
  NAND3_X1 U12496 ( .A1(n10049), .A2(n14313), .A3(n9921), .ZN(n10497) );
  OAI211_X1 U12497 ( .C1(n7215), .C2(n14915), .A(n10503), .B(n10497), .ZN(
        n9922) );
  NOR2_X1 U12498 ( .A1(n9923), .A2(n9922), .ZN(n14889) );
  NAND2_X1 U12499 ( .A1(n14932), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9924) );
  OAI21_X1 U12500 ( .B1(n14889), .B2(n14932), .A(n9924), .ZN(P2_U3500) );
  NAND2_X1 U12501 ( .A1(n12942), .A2(n12126), .ZN(n10095) );
  XNOR2_X1 U12502 ( .A(n10092), .B(n10093), .ZN(n9935) );
  NAND2_X1 U12503 ( .A1(n12941), .A2(n12902), .ZN(n9928) );
  NAND2_X1 U12504 ( .A1(n12943), .A2(n12901), .ZN(n9927) );
  AND2_X1 U12505 ( .A1(n9928), .A2(n9927), .ZN(n10268) );
  INV_X1 U12506 ( .A(n10268), .ZN(n9929) );
  AOI22_X1 U12507 ( .A1(n12913), .A2(n14891), .B1(n12897), .B2(n9929), .ZN(
        n9934) );
  OR2_X1 U12508 ( .A1(n9931), .A2(n9930), .ZN(n9932) );
  NAND2_X1 U12509 ( .A1(n9932), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12894) );
  MUX2_X1 U12510 ( .A(P2_STATE_REG_SCAN_IN), .B(n12894), .S(n10270), .Z(n9933)
         );
  OAI211_X1 U12511 ( .C1(n9935), .C2(n12908), .A(n9934), .B(n9933), .ZN(
        P2_U3190) );
  OAI21_X1 U12512 ( .B1(n9937), .B2(n9936), .A(n9951), .ZN(n9944) );
  INV_X1 U12513 ( .A(n9938), .ZN(n9953) );
  NAND2_X1 U12514 ( .A1(n9947), .A2(n9953), .ZN(n9943) );
  AND3_X1 U12515 ( .A1(n9941), .A2(n9940), .A3(n9939), .ZN(n9942) );
  NAND3_X1 U12516 ( .A1(n9944), .A2(n9943), .A3(n9942), .ZN(n9945) );
  NAND2_X1 U12517 ( .A1(n9945), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9949) );
  INV_X1 U12518 ( .A(n11755), .ZN(n9959) );
  NAND3_X1 U12519 ( .A1(n9947), .A2(n9946), .A3(n9959), .ZN(n9948) );
  INV_X1 U12520 ( .A(n12376), .ZN(n12358) );
  NAND2_X1 U12521 ( .A1(n12358), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10086) );
  INV_X1 U12522 ( .A(n10086), .ZN(n10039) );
  INV_X1 U12523 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n9963) );
  NAND2_X1 U12524 ( .A1(n9954), .A2(n9950), .ZN(n12378) );
  OR2_X1 U12525 ( .A1(n12378), .A2(n15117), .ZN(n12278) );
  NAND2_X1 U12526 ( .A1(n9951), .A2(n15146), .ZN(n9952) );
  OR2_X1 U12527 ( .A1(n9957), .A2(n9952), .ZN(n9956) );
  NAND2_X1 U12528 ( .A1(n9954), .A2(n9953), .ZN(n9955) );
  AND2_X2 U12529 ( .A1(n9956), .A2(n9955), .ZN(n12382) );
  OR2_X1 U12530 ( .A1(n9957), .A2(n15146), .ZN(n9960) );
  NOR2_X1 U12531 ( .A1(n15146), .A2(n15126), .ZN(n9958) );
  OAI22_X1 U12532 ( .A1(n11722), .A2(n12382), .B1(n10056), .B2(n12352), .ZN(
        n9961) );
  AOI21_X1 U12533 ( .B1(n12289), .B2(n12409), .A(n9961), .ZN(n9962) );
  OAI21_X1 U12534 ( .B1(n10039), .B2(n9963), .A(n9962), .ZN(P3_U3172) );
  OAI222_X1 U12535 ( .A1(P3_U3151), .A2(n9966), .B1(n12787), .B2(n9965), .C1(
        n12785), .C2(n9964), .ZN(P3_U3276) );
  MUX2_X1 U12536 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12452), .Z(n10815) );
  XOR2_X1 U12537 ( .A(n10795), .B(n10815), .Z(n10816) );
  INV_X1 U12538 ( .A(n9967), .ZN(n9980) );
  OAI22_X1 U12539 ( .A1(n9970), .A2(n9969), .B1(n9968), .B2(n9980), .ZN(n14951) );
  MUX2_X1 U12540 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n12452), .Z(n9971) );
  XNOR2_X1 U12541 ( .A(n9971), .B(n14956), .ZN(n14952) );
  INV_X1 U12542 ( .A(n9971), .ZN(n9972) );
  XOR2_X1 U12543 ( .A(n10816), .B(n10817), .Z(n9991) );
  INV_X1 U12544 ( .A(n15025), .ZN(n15098) );
  INV_X1 U12545 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n9978) );
  INV_X1 U12546 ( .A(n14956), .ZN(n9983) );
  INV_X1 U12547 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n15566) );
  INV_X1 U12548 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n15189) );
  MUX2_X1 U12549 ( .A(n15189), .B(P3_REG1_REG_4__SCAN_IN), .S(n10795), .Z(
        n9975) );
  NOR3_X1 U12550 ( .A1(n9974), .A2(n9975), .A3(n14947), .ZN(n9976) );
  OAI21_X1 U12551 ( .B1(n10805), .B2(n9976), .A(n14966), .ZN(n9977) );
  NAND2_X1 U12552 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n10445) );
  OAI211_X1 U12553 ( .C1(n15098), .C2(n9978), .A(n9977), .B(n10445), .ZN(n9989) );
  INV_X1 U12554 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n14945) );
  AOI21_X1 U12555 ( .B1(P3_REG2_REG_2__SCAN_IN), .B2(n9980), .A(n9979), .ZN(
        n9981) );
  INV_X1 U12556 ( .A(n9981), .ZN(n9984) );
  INV_X1 U12557 ( .A(n9986), .ZN(n9982) );
  OAI21_X1 U12558 ( .B1(n9984), .B2(n9983), .A(n9982), .ZN(n14946) );
  MUX2_X1 U12559 ( .A(n7392), .B(P3_REG2_REG_4__SCAN_IN), .S(n10795), .Z(n9985) );
  OR3_X1 U12560 ( .A1(n9986), .A2(n9985), .A3(n14944), .ZN(n9987) );
  AOI21_X1 U12561 ( .B1(n10796), .B2(n9987), .A(n15110), .ZN(n9988) );
  AOI211_X1 U12562 ( .C1(n15016), .C2(n10795), .A(n9989), .B(n9988), .ZN(n9990) );
  OAI21_X1 U12563 ( .B1(n9991), .B2(n15082), .A(n9990), .ZN(P3_U3186) );
  OAI22_X1 U12564 ( .A1(n10003), .A2(P1_D_REG_1__SCAN_IN), .B1(n14038), .B2(
        n9992), .ZN(n10290) );
  NOR4_X1 U12565 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n10001) );
  NOR4_X1 U12566 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n10000) );
  INV_X1 U12567 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n15283) );
  INV_X1 U12568 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n15567) );
  INV_X1 U12569 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n15416) );
  INV_X1 U12570 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n15458) );
  NAND4_X1 U12571 ( .A1(n15283), .A2(n15567), .A3(n15416), .A4(n15458), .ZN(
        n9998) );
  NOR4_X1 U12572 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n9996) );
  NOR4_X1 U12573 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n9995) );
  NOR4_X1 U12574 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9994) );
  NOR4_X1 U12575 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n9993) );
  NAND4_X1 U12576 ( .A1(n9996), .A2(n9995), .A3(n9994), .A4(n9993), .ZN(n9997)
         );
  NOR4_X1 U12577 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        n9998), .A4(n9997), .ZN(n9999) );
  AND3_X1 U12578 ( .A1(n10001), .A2(n10000), .A3(n9999), .ZN(n10002) );
  NOR2_X1 U12579 ( .A1(n10003), .A2(n10002), .ZN(n10289) );
  NOR2_X1 U12580 ( .A1(n10290), .A2(n10289), .ZN(n10875) );
  INV_X1 U12581 ( .A(n10003), .ZN(n10006) );
  INV_X1 U12582 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10005) );
  NOR2_X1 U12583 ( .A1(n14038), .A2(n11331), .ZN(n10004) );
  NAND2_X1 U12584 ( .A1(n10875), .A2(n10318), .ZN(n10022) );
  INV_X1 U12585 ( .A(n10022), .ZN(n10011) );
  AND2_X1 U12586 ( .A1(n10871), .A2(n10007), .ZN(n10010) );
  NAND2_X1 U12587 ( .A1(n10012), .A2(n11825), .ZN(n10021) );
  INV_X1 U12588 ( .A(n10451), .ZN(n10018) );
  AOI22_X1 U12589 ( .A1(n10014), .A2(n10365), .B1(n10018), .B2(n14044), .ZN(
        n10015) );
  INV_X1 U12590 ( .A(n10351), .ZN(n10017) );
  NAND2_X1 U12591 ( .A1(n10017), .A2(n10014), .ZN(n10020) );
  AOI22_X1 U12592 ( .A1(n10365), .A2(n6643), .B1(n10018), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n10019) );
  NAND2_X1 U12593 ( .A1(n10020), .A2(n10019), .ZN(n10149) );
  XNOR2_X1 U12594 ( .A(n10147), .B(n10149), .ZN(n13612) );
  NAND2_X1 U12595 ( .A1(n10873), .A2(n10022), .ZN(n10452) );
  AND2_X1 U12596 ( .A1(n10452), .A2(n10871), .ZN(n11017) );
  INV_X1 U12597 ( .A(n10293), .ZN(n10876) );
  NAND2_X1 U12598 ( .A1(n10452), .A2(n10876), .ZN(n10161) );
  INV_X1 U12599 ( .A(n10161), .ZN(n12174) );
  INV_X1 U12600 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10911) );
  OR2_X1 U12601 ( .A1(n10022), .A2(n10293), .ZN(n13546) );
  OR2_X1 U12602 ( .A1(n13546), .A2(n14539), .ZN(n13571) );
  OAI22_X1 U12603 ( .A1(n12174), .A2(n10911), .B1(n13571), .B2(n10152), .ZN(
        n10024) );
  AOI21_X1 U12604 ( .B1(n10365), .B2(n14358), .A(n10024), .ZN(n10025) );
  OAI21_X1 U12605 ( .B1(n13564), .B2(n13612), .A(n10025), .ZN(P1_U3232) );
  INV_X1 U12606 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10038) );
  NAND2_X1 U12607 ( .A1(n11559), .A2(n12483), .ZN(n10026) );
  NAND2_X1 U12608 ( .A1(n10026), .A2(n10326), .ZN(n10027) );
  NAND3_X1 U12609 ( .A1(n12409), .A2(n12220), .A3(n10028), .ZN(n10029) );
  NAND2_X1 U12610 ( .A1(n15116), .A2(n12220), .ZN(n10030) );
  NAND2_X1 U12611 ( .A1(n10031), .A2(n10030), .ZN(n10032) );
  INV_X1 U12612 ( .A(n15113), .ZN(n11565) );
  NAND3_X1 U12613 ( .A1(n11565), .A2(n6960), .A3(n12273), .ZN(n10033) );
  INV_X1 U12614 ( .A(n12382), .ZN(n12282) );
  NAND2_X1 U12615 ( .A1(n10034), .A2(n12282), .ZN(n10037) );
  NOR2_X1 U12616 ( .A1(n12378), .A2(n15119), .ZN(n12291) );
  OAI22_X1 U12617 ( .A1(n15112), .A2(n12352), .B1(n15118), .B2(n12278), .ZN(
        n10035) );
  AOI21_X1 U12618 ( .B1(n12291), .B2(n12411), .A(n10035), .ZN(n10036) );
  OAI211_X1 U12619 ( .C1(n10039), .C2(n10038), .A(n10037), .B(n10036), .ZN(
        P3_U3162) );
  INV_X1 U12620 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10041) );
  INV_X1 U12621 ( .A(n10040), .ZN(n10042) );
  INV_X1 U12622 ( .A(n14786), .ZN(n10064) );
  OAI222_X1 U12623 ( .A1(n13357), .A2(n10041), .B1(n13359), .B2(n10042), .C1(
        n10064), .C2(P2_U3088), .ZN(P2_U3315) );
  INV_X1 U12624 ( .A(n13671), .ZN(n10422) );
  OAI222_X1 U12625 ( .A1(n14039), .A2(n10043), .B1(n10724), .B2(n10042), .C1(
        n10422), .C2(P1_U3086), .ZN(P1_U3343) );
  XNOR2_X1 U12626 ( .A(n10044), .B(n12069), .ZN(n14842) );
  XNOR2_X1 U12627 ( .A(n10045), .B(n12069), .ZN(n10047) );
  AOI21_X1 U12628 ( .B1(n10047), .B2(n14304), .A(n10046), .ZN(n14836) );
  INV_X1 U12629 ( .A(n10273), .ZN(n10048) );
  AOI21_X1 U12630 ( .B1(n11851), .B2(n10049), .A(n10048), .ZN(n14843) );
  AOI22_X1 U12631 ( .A1(n14843), .A2(n14313), .B1(n14892), .B2(n11851), .ZN(
        n10050) );
  OAI211_X1 U12632 ( .C1(n14842), .C2(n14895), .A(n14836), .B(n10050), .ZN(
        n10052) );
  NAND2_X1 U12633 ( .A1(n10052), .A2(n14934), .ZN(n10051) );
  OAI21_X1 U12634 ( .B1(n14934), .B2(n9650), .A(n10051), .ZN(P2_U3501) );
  INV_X1 U12635 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10054) );
  NAND2_X1 U12636 ( .A1(n10052), .A2(n14924), .ZN(n10053) );
  OAI21_X1 U12637 ( .B1(n14924), .B2(n10054), .A(n10053), .ZN(P2_U3436) );
  OAI22_X1 U12638 ( .A1(n12721), .A2(n10056), .B1(n15202), .B2(n10055), .ZN(
        n10057) );
  INV_X1 U12639 ( .A(n10057), .ZN(n10058) );
  OAI21_X1 U12640 ( .B1(n10284), .B2(n8976), .A(n10058), .ZN(P3_U3459) );
  INV_X1 U12641 ( .A(n10059), .ZN(n10090) );
  INV_X1 U12642 ( .A(n14039), .ZN(n11525) );
  AOI22_X1 U12643 ( .A1(n14449), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n11525), .ZN(n10060) );
  OAI21_X1 U12644 ( .B1(n10090), .B2(n10724), .A(n10060), .ZN(P1_U3342) );
  INV_X1 U12645 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n15385) );
  NAND2_X1 U12646 ( .A1(n10069), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n10061) );
  NAND2_X1 U12647 ( .A1(n10062), .A2(n10061), .ZN(n14762) );
  INV_X1 U12648 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10063) );
  MUX2_X1 U12649 ( .A(n10063), .B(P2_REG2_REG_11__SCAN_IN), .S(n10073), .Z(
        n14761) );
  NAND2_X1 U12650 ( .A1(n14771), .A2(n10063), .ZN(n14780) );
  MUX2_X1 U12651 ( .A(n15385), .B(P2_REG2_REG_12__SCAN_IN), .S(n14786), .Z(
        n14781) );
  AOI21_X1 U12652 ( .B1(n14782), .B2(n14780), .A(n14781), .ZN(n14779) );
  AOI21_X1 U12653 ( .B1(n15385), .B2(n10064), .A(n14779), .ZN(n10338) );
  INV_X1 U12654 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10065) );
  MUX2_X1 U12655 ( .A(n10065), .B(P2_REG2_REG_13__SCAN_IN), .S(n10335), .Z(
        n10336) );
  XNOR2_X1 U12656 ( .A(n10338), .B(n10336), .ZN(n10079) );
  INV_X1 U12657 ( .A(n10335), .ZN(n10089) );
  NOR2_X1 U12658 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11299), .ZN(n10066) );
  AOI21_X1 U12659 ( .B1(n14825), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n10066), 
        .ZN(n10067) );
  OAI21_X1 U12660 ( .B1(n10089), .B2(n14833), .A(n10067), .ZN(n10078) );
  INV_X1 U12661 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10068) );
  MUX2_X1 U12662 ( .A(n10068), .B(P2_REG1_REG_13__SCAN_IN), .S(n10335), .Z(
        n10076) );
  NAND2_X1 U12663 ( .A1(n10069), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10070) );
  NAND2_X1 U12664 ( .A1(n10071), .A2(n10070), .ZN(n14766) );
  INV_X1 U12665 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10072) );
  MUX2_X1 U12666 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n10072), .S(n10073), .Z(
        n14765) );
  AND2_X1 U12667 ( .A1(n14766), .A2(n14765), .ZN(n14768) );
  AOI21_X1 U12668 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n10073), .A(n14768), 
        .ZN(n14778) );
  INV_X1 U12669 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10074) );
  MUX2_X1 U12670 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n10074), .S(n14786), .Z(
        n14777) );
  NAND2_X1 U12671 ( .A1(n14778), .A2(n14777), .ZN(n14776) );
  OAI21_X1 U12672 ( .B1(n14786), .B2(P2_REG1_REG_12__SCAN_IN), .A(n14776), 
        .ZN(n10075) );
  NOR2_X1 U12673 ( .A1(n10075), .A2(n10076), .ZN(n10329) );
  AOI211_X1 U12674 ( .C1(n10076), .C2(n10075), .A(n14819), .B(n10329), .ZN(
        n10077) );
  AOI211_X1 U12675 ( .C1(n14811), .C2(n10079), .A(n10078), .B(n10077), .ZN(
        n10080) );
  INV_X1 U12676 ( .A(n10080), .ZN(P2_U3227) );
  XNOR2_X1 U12677 ( .A(n10083), .B(n12220), .ZN(n10435) );
  XNOR2_X1 U12678 ( .A(n10435), .B(n15118), .ZN(n10438) );
  NAND2_X1 U12679 ( .A1(n10082), .A2(n10081), .ZN(n10439) );
  XOR2_X1 U12680 ( .A(n10438), .B(n10439), .Z(n10088) );
  INV_X1 U12681 ( .A(n12291), .ZN(n12237) );
  AOI22_X1 U12682 ( .A1(n12407), .A2(n12289), .B1(n10083), .B2(n12380), .ZN(
        n10084) );
  OAI21_X1 U12683 ( .B1(n10586), .B2(n12237), .A(n10084), .ZN(n10085) );
  AOI21_X1 U12684 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(n10086), .A(n10085), .ZN(
        n10087) );
  OAI21_X1 U12685 ( .B1(n10088), .B2(n12382), .A(n10087), .ZN(P3_U3177) );
  OAI222_X1 U12686 ( .A1(n13357), .A2(n10091), .B1(n13359), .B2(n10090), .C1(
        n10089), .C2(P2_U3088), .ZN(P2_U3314) );
  INV_X1 U12687 ( .A(n10094), .ZN(n10097) );
  INV_X1 U12688 ( .A(n10095), .ZN(n10096) );
  XNOR2_X1 U12689 ( .A(n11870), .B(n9889), .ZN(n10099) );
  NAND2_X1 U12690 ( .A1(n12941), .A2(n12126), .ZN(n10100) );
  NAND2_X1 U12691 ( .A1(n10099), .A2(n10100), .ZN(n10250) );
  INV_X1 U12692 ( .A(n10099), .ZN(n10102) );
  INV_X1 U12693 ( .A(n10100), .ZN(n10101) );
  NAND2_X1 U12694 ( .A1(n10102), .A2(n10101), .ZN(n10103) );
  AND2_X1 U12695 ( .A1(n10250), .A2(n10103), .ZN(n10104) );
  NAND2_X1 U12696 ( .A1(n10105), .A2(n10104), .ZN(n10251) );
  OAI21_X1 U12697 ( .B1(n10105), .B2(n10104), .A(n10251), .ZN(n10106) );
  NAND2_X1 U12698 ( .A1(n10106), .A2(n12887), .ZN(n10114) );
  INV_X1 U12699 ( .A(n12894), .ZN(n12903) );
  NAND2_X1 U12700 ( .A1(n12940), .A2(n12902), .ZN(n10108) );
  NAND2_X1 U12701 ( .A1(n12942), .A2(n12901), .ZN(n10107) );
  AND2_X1 U12702 ( .A1(n10108), .A2(n10107), .ZN(n10374) );
  INV_X1 U12703 ( .A(n10374), .ZN(n10109) );
  NAND2_X1 U12704 ( .A1(n10109), .A2(n12897), .ZN(n10111) );
  OAI211_X1 U12705 ( .C1(n12900), .C2(n10378), .A(n10111), .B(n10110), .ZN(
        n10112) );
  AOI21_X1 U12706 ( .B1(n10488), .B2(n12903), .A(n10112), .ZN(n10113) );
  NAND2_X1 U12707 ( .A1(n10114), .A2(n10113), .ZN(P2_U3202) );
  INV_X1 U12708 ( .A(n10133), .ZN(n10235) );
  INV_X1 U12709 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10117) );
  INV_X1 U12710 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10116) );
  XNOR2_X1 U12711 ( .A(n10128), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n13607) );
  AND2_X1 U12712 ( .A1(n14044), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n13613) );
  NAND2_X1 U12713 ( .A1(n13607), .A2(n13613), .ZN(n13606) );
  NAND2_X1 U12714 ( .A1(n13602), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10115) );
  NAND2_X1 U12715 ( .A1(n13606), .A2(n10115), .ZN(n13622) );
  XNOR2_X1 U12716 ( .A(n13620), .B(n10116), .ZN(n13623) );
  NAND2_X1 U12717 ( .A1(n13622), .A2(n13623), .ZN(n13621) );
  OAI21_X1 U12718 ( .B1(n10116), .B2(n10130), .A(n13621), .ZN(n13634) );
  OAI21_X1 U12719 ( .B1(n13630), .B2(n10117), .A(n13633), .ZN(n13650) );
  INV_X1 U12720 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n11070) );
  MUX2_X1 U12721 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n11070), .S(n13645), .Z(
        n13651) );
  NAND2_X1 U12722 ( .A1(n13650), .A2(n13651), .ZN(n13649) );
  XNOR2_X1 U12723 ( .A(n10235), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n10239) );
  INV_X1 U12724 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10905) );
  MUX2_X1 U12725 ( .A(n10905), .B(P1_REG2_REG_6__SCAN_IN), .S(n10183), .Z(
        n10178) );
  NOR2_X1 U12726 ( .A1(n10179), .A2(n10178), .ZN(n10177) );
  INV_X1 U12727 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10118) );
  MUX2_X1 U12728 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n10118), .S(n10171), .Z(
        n10119) );
  INV_X1 U12729 ( .A(n10119), .ZN(n10166) );
  XNOR2_X1 U12730 ( .A(n10222), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n10226) );
  AOI21_X1 U12731 ( .B1(n10222), .B2(P1_REG2_REG_8__SCAN_IN), .A(n10225), .ZN(
        n10214) );
  INV_X1 U12732 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10120) );
  MUX2_X1 U12733 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n10120), .S(n10208), .Z(
        n10121) );
  INV_X1 U12734 ( .A(n10121), .ZN(n10213) );
  NOR2_X1 U12735 ( .A1(n10214), .A2(n10213), .ZN(n10212) );
  INV_X1 U12736 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10122) );
  MUX2_X1 U12737 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n10122), .S(n10424), .Z(
        n10123) );
  INV_X1 U12738 ( .A(n10123), .ZN(n10125) );
  NOR2_X1 U12739 ( .A1(n9571), .A2(n6641), .ZN(n10124) );
  INV_X1 U12740 ( .A(n14521), .ZN(n14487) );
  AOI211_X1 U12741 ( .C1(n10126), .C2(n10125), .A(n14487), .B(n10423), .ZN(
        n10143) );
  INV_X1 U12742 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10127) );
  MUX2_X1 U12743 ( .A(n10127), .B(P1_REG1_REG_10__SCAN_IN), .S(n10424), .Z(
        n10138) );
  INV_X1 U12744 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n14677) );
  MUX2_X1 U12745 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n14677), .S(n13645), .Z(
        n13648) );
  INV_X1 U12746 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10132) );
  MUX2_X1 U12747 ( .A(n10132), .B(P1_REG1_REG_3__SCAN_IN), .S(n13630), .Z(
        n13638) );
  INV_X1 U12748 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10131) );
  XNOR2_X1 U12749 ( .A(n10128), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n13605) );
  AND2_X1 U12750 ( .A1(n14044), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n13604) );
  NAND2_X1 U12751 ( .A1(n13605), .A2(n13604), .ZN(n13603) );
  NAND2_X1 U12752 ( .A1(n13602), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10129) );
  NAND2_X1 U12753 ( .A1(n13603), .A2(n10129), .ZN(n13625) );
  XNOR2_X1 U12754 ( .A(n13620), .B(n10131), .ZN(n13626) );
  NAND2_X1 U12755 ( .A1(n13625), .A2(n13626), .ZN(n13624) );
  OAI21_X1 U12756 ( .B1(n10131), .B2(n10130), .A(n13624), .ZN(n13637) );
  NAND2_X1 U12757 ( .A1(n13638), .A2(n13637), .ZN(n13636) );
  OAI21_X1 U12758 ( .B1(n13630), .B2(n10132), .A(n13636), .ZN(n13647) );
  XNOR2_X1 U12759 ( .A(n10133), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n10234) );
  NAND2_X1 U12760 ( .A1(n10233), .A2(n10234), .ZN(n10232) );
  OAI21_X1 U12761 ( .B1(n10235), .B2(P1_REG1_REG_5__SCAN_IN), .A(n10232), .ZN(
        n10181) );
  XNOR2_X1 U12762 ( .A(n10183), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n10182) );
  NOR2_X1 U12763 ( .A1(n10181), .A2(n10182), .ZN(n10180) );
  INV_X1 U12764 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10134) );
  MUX2_X1 U12765 ( .A(n10134), .B(P1_REG1_REG_7__SCAN_IN), .S(n10171), .Z(
        n10169) );
  NOR2_X1 U12766 ( .A1(n10170), .A2(n10169), .ZN(n10168) );
  AOI21_X1 U12767 ( .B1(n10171), .B2(P1_REG1_REG_7__SCAN_IN), .A(n10168), .ZN(
        n10221) );
  INV_X1 U12768 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10135) );
  MUX2_X1 U12769 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10135), .S(n10222), .Z(
        n10220) );
  NAND2_X1 U12770 ( .A1(n10221), .A2(n10220), .ZN(n10219) );
  INV_X1 U12771 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10136) );
  MUX2_X1 U12772 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10136), .S(n10208), .Z(
        n10207) );
  OAI21_X1 U12773 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n10208), .A(n10205), .ZN(
        n10137) );
  NAND2_X1 U12774 ( .A1(n10139), .A2(n6641), .ZN(n14483) );
  NOR2_X1 U12775 ( .A1(n10137), .A2(n10138), .ZN(n10414) );
  AOI211_X1 U12776 ( .C1(n10138), .C2(n10137), .A(n14483), .B(n10414), .ZN(
        n10142) );
  NAND2_X1 U12777 ( .A1(n10139), .A2(n9571), .ZN(n14525) );
  NAND2_X1 U12778 ( .A1(n14494), .A2(n10424), .ZN(n10140) );
  NAND2_X1 U12779 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n14348)
         );
  OAI211_X1 U12780 ( .C1(n14066), .C2(n14529), .A(n10140), .B(n14348), .ZN(
        n10141) );
  OR3_X1 U12781 ( .A1(n10143), .A2(n10142), .A3(n10141), .ZN(P1_U3253) );
  INV_X1 U12782 ( .A(n14358), .ZN(n13576) );
  NAND2_X1 U12783 ( .A1(n10298), .A2(n13685), .ZN(n10145) );
  AND2_X2 U12784 ( .A1(n10145), .A2(n10299), .ZN(n11318) );
  XNOR2_X1 U12785 ( .A(n10146), .B(n11318), .ZN(n10462) );
  OAI22_X1 U12786 ( .A1(n10144), .A2(n13405), .B1(n14574), .B2(n13407), .ZN(
        n10463) );
  XNOR2_X1 U12787 ( .A(n10462), .B(n10463), .ZN(n10159) );
  INV_X1 U12788 ( .A(n10147), .ZN(n10148) );
  INV_X1 U12789 ( .A(n10149), .ZN(n10150) );
  OAI22_X1 U12790 ( .A1(n10152), .A2(n13407), .B1(n6672), .B2(n13393), .ZN(
        n10153) );
  XNOR2_X1 U12791 ( .A(n10153), .B(n11318), .ZN(n10154) );
  OAI22_X1 U12792 ( .A1(n10152), .A2(n13405), .B1(n12178), .B2(n13407), .ZN(
        n10155) );
  XNOR2_X1 U12793 ( .A(n10155), .B(n10154), .ZN(n12170) );
  NAND2_X1 U12794 ( .A1(n12172), .A2(n12170), .ZN(n12171) );
  INV_X1 U12795 ( .A(n10154), .ZN(n10156) );
  OR2_X1 U12796 ( .A1(n10156), .A2(n10155), .ZN(n10157) );
  NAND2_X1 U12797 ( .A1(n10158), .A2(n10159), .ZN(n10466) );
  OAI21_X1 U12798 ( .B1(n10159), .B2(n10158), .A(n10466), .ZN(n10160) );
  NAND2_X1 U12799 ( .A1(n10160), .A2(n14350), .ZN(n10164) );
  AOI22_X1 U12800 ( .A1(n13599), .A2(n13854), .B1(n13913), .B2(n13597), .ZN(
        n10310) );
  INV_X1 U12801 ( .A(n10310), .ZN(n10162) );
  AOI22_X1 U12802 ( .A1(n10162), .A2(n14359), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n10161), .ZN(n10163) );
  OAI211_X1 U12803 ( .C1(n14574), .C2(n13576), .A(n10164), .B(n10163), .ZN(
        P1_U3237) );
  AOI211_X1 U12804 ( .C1(n10167), .C2(n10166), .A(n14487), .B(n10165), .ZN(
        n10176) );
  AOI211_X1 U12805 ( .C1(n10170), .C2(n10169), .A(n14483), .B(n10168), .ZN(
        n10175) );
  INV_X1 U12806 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n14060) );
  NAND2_X1 U12807 ( .A1(n14494), .A2(n10171), .ZN(n10173) );
  NAND2_X1 U12808 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n10172) );
  OAI211_X1 U12809 ( .C1(n14060), .C2(n14529), .A(n10173), .B(n10172), .ZN(
        n10174) );
  OR3_X1 U12810 ( .A1(n10176), .A2(n10175), .A3(n10174), .ZN(P1_U3250) );
  AOI211_X1 U12811 ( .C1(n10179), .C2(n10178), .A(n10177), .B(n14487), .ZN(
        n10188) );
  AOI211_X1 U12812 ( .C1(n10182), .C2(n10181), .A(n10180), .B(n14483), .ZN(
        n10187) );
  NAND2_X1 U12813 ( .A1(n14494), .A2(n10183), .ZN(n10185) );
  NAND2_X1 U12814 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n10184) );
  OAI211_X1 U12815 ( .C1(n14047), .C2(n14529), .A(n10185), .B(n10184), .ZN(
        n10186) );
  OR3_X1 U12816 ( .A1(n10188), .A2(n10187), .A3(n10186), .ZN(P1_U3249) );
  INV_X1 U12817 ( .A(n10189), .ZN(n10192) );
  NOR2_X1 U12818 ( .A1(n10190), .A2(n14880), .ZN(n10191) );
  NAND2_X1 U12819 ( .A1(n10192), .A2(n10191), .ZN(n10201) );
  NAND2_X1 U12820 ( .A1(n9870), .A2(n13171), .ZN(n10194) );
  AOI21_X1 U12821 ( .B1(n14884), .B2(n10194), .A(n10193), .ZN(n14886) );
  INV_X1 U12822 ( .A(n11842), .ZN(n10263) );
  OR2_X1 U12823 ( .A1(n13211), .A2(n10263), .ZN(n11115) );
  INV_X1 U12824 ( .A(n11115), .ZN(n14845) );
  INV_X1 U12825 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10197) );
  OAI22_X1 U12826 ( .A1(n14837), .A2(n10197), .B1(n10196), .B2(n13194), .ZN(
        n10198) );
  AOI21_X1 U12827 ( .B1(n14845), .B2(n14884), .A(n10198), .ZN(n10203) );
  INV_X1 U12828 ( .A(n10199), .ZN(n10200) );
  NOR2_X1 U12829 ( .A1(n13213), .A2(n11181), .ZN(n14844) );
  OAI21_X1 U12830 ( .B1(n14307), .B2(n14844), .A(n14882), .ZN(n10202) );
  OAI211_X1 U12831 ( .C1(n13211), .C2(n14886), .A(n10203), .B(n10202), .ZN(
        P2_U3265) );
  INV_X1 U12832 ( .A(P3_DATAO_REG_24__SCAN_IN), .ZN(n15445) );
  NAND2_X1 U12833 ( .A1(n12305), .A2(P3_U3897), .ZN(n10204) );
  OAI21_X1 U12834 ( .B1(P3_U3897), .B2(n15445), .A(n10204), .ZN(P3_U3515) );
  OAI21_X1 U12835 ( .B1(n10207), .B2(n10206), .A(n10205), .ZN(n10217) );
  INV_X1 U12836 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10211) );
  NAND2_X1 U12837 ( .A1(n14494), .A2(n10208), .ZN(n10210) );
  NAND2_X1 U12838 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n10209) );
  OAI211_X1 U12839 ( .C1(n10211), .C2(n14529), .A(n10210), .B(n10209), .ZN(
        n10216) );
  AOI211_X1 U12840 ( .C1(n10214), .C2(n10213), .A(n14487), .B(n10212), .ZN(
        n10215) );
  AOI211_X1 U12841 ( .C1(n14517), .C2(n10217), .A(n10216), .B(n10215), .ZN(
        n10218) );
  INV_X1 U12842 ( .A(n10218), .ZN(P1_U3252) );
  OAI21_X1 U12843 ( .B1(n10221), .B2(n10220), .A(n10219), .ZN(n10230) );
  INV_X1 U12844 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n14046) );
  NAND2_X1 U12845 ( .A1(n14494), .A2(n10222), .ZN(n10224) );
  NAND2_X1 U12846 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n10223) );
  OAI211_X1 U12847 ( .C1(n14046), .C2(n14529), .A(n10224), .B(n10223), .ZN(
        n10229) );
  AOI211_X1 U12848 ( .C1(n10227), .C2(n10226), .A(n14487), .B(n10225), .ZN(
        n10228) );
  AOI211_X1 U12849 ( .C1(n14517), .C2(n10230), .A(n10229), .B(n10228), .ZN(
        n10231) );
  INV_X1 U12850 ( .A(n10231), .ZN(P1_U3251) );
  OAI21_X1 U12851 ( .B1(n10234), .B2(n10233), .A(n10232), .ZN(n10243) );
  INV_X1 U12852 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14055) );
  NAND2_X1 U12853 ( .A1(n14494), .A2(n10235), .ZN(n10237) );
  NAND2_X1 U12854 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n10236) );
  OAI211_X1 U12855 ( .C1(n14055), .C2(n14529), .A(n10237), .B(n10236), .ZN(
        n10242) );
  AOI211_X1 U12856 ( .C1(n10240), .C2(n10239), .A(n10238), .B(n14487), .ZN(
        n10241) );
  AOI211_X1 U12857 ( .C1(n14517), .C2(n10243), .A(n10242), .B(n10241), .ZN(
        n10244) );
  INV_X1 U12858 ( .A(n10244), .ZN(P1_U3248) );
  XNOR2_X1 U12859 ( .A(n11876), .B(n9889), .ZN(n10245) );
  NAND2_X1 U12860 ( .A1(n12940), .A2(n12126), .ZN(n10246) );
  NAND2_X1 U12861 ( .A1(n10245), .A2(n10246), .ZN(n10476) );
  INV_X1 U12862 ( .A(n10245), .ZN(n10248) );
  INV_X1 U12863 ( .A(n10246), .ZN(n10247) );
  NAND2_X1 U12864 ( .A1(n10248), .A2(n10247), .ZN(n10249) );
  AND2_X1 U12865 ( .A1(n10476), .A2(n10249), .ZN(n10253) );
  NAND2_X1 U12866 ( .A1(n10251), .A2(n10250), .ZN(n10252) );
  NAND2_X1 U12867 ( .A1(n10252), .A2(n10253), .ZN(n10477) );
  OAI21_X1 U12868 ( .B1(n10253), .B2(n10252), .A(n10477), .ZN(n10254) );
  NAND2_X1 U12869 ( .A1(n10254), .A2(n12887), .ZN(n10262) );
  INV_X1 U12870 ( .A(n12897), .ZN(n12906) );
  NAND2_X1 U12871 ( .A1(n12939), .A2(n12902), .ZN(n10256) );
  NAND2_X1 U12872 ( .A1(n12941), .A2(n12901), .ZN(n10255) );
  NAND2_X1 U12873 ( .A1(n10256), .A2(n10255), .ZN(n10400) );
  INV_X1 U12874 ( .A(n10400), .ZN(n10259) );
  INV_X1 U12875 ( .A(n10257), .ZN(n10258) );
  OAI21_X1 U12876 ( .B1(n12906), .B2(n10259), .A(n10258), .ZN(n10260) );
  AOI21_X1 U12877 ( .B1(n10405), .B2(n12903), .A(n10260), .ZN(n10261) );
  OAI211_X1 U12878 ( .C1(n14901), .C2(n12900), .A(n10262), .B(n10261), .ZN(
        P2_U3199) );
  AND2_X1 U12879 ( .A1(n10263), .A2(n9870), .ZN(n10264) );
  XNOR2_X1 U12880 ( .A(n12068), .B(n10265), .ZN(n14894) );
  XNOR2_X1 U12881 ( .A(n12068), .B(n10266), .ZN(n10267) );
  NAND2_X1 U12882 ( .A1(n10267), .A2(n14304), .ZN(n10269) );
  NAND2_X1 U12883 ( .A1(n10269), .A2(n10268), .ZN(n14896) );
  AOI21_X1 U12884 ( .B1(n14841), .B2(n10270), .A(n14896), .ZN(n10271) );
  MUX2_X1 U12885 ( .A(n10272), .B(n10271), .S(n14837), .Z(n10275) );
  AOI211_X1 U12886 ( .C1(n14891), .C2(n10273), .A(n13049), .B(n10370), .ZN(
        n14890) );
  AOI22_X1 U12887 ( .A1(n14890), .A2(n14315), .B1(n14307), .B2(n14891), .ZN(
        n10274) );
  OAI211_X1 U12888 ( .C1(n13182), .C2(n14894), .A(n10275), .B(n10274), .ZN(
        P2_U3262) );
  NAND2_X1 U12889 ( .A1(n10277), .A2(n10276), .ZN(n10281) );
  NAND2_X1 U12890 ( .A1(n10279), .A2(n10278), .ZN(n10280) );
  NAND2_X1 U12891 ( .A1(n10283), .A2(n10282), .ZN(n10285) );
  INV_X1 U12892 ( .A(n15595), .ZN(n15131) );
  MUX2_X1 U12893 ( .A(n15429), .B(n10284), .S(n15131), .Z(n10288) );
  INV_X1 U12894 ( .A(n15593), .ZN(n12640) );
  AOI22_X1 U12895 ( .A1(n12640), .A2(n10286), .B1(n15591), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n10287) );
  NAND2_X1 U12896 ( .A1(n10288), .A2(n10287), .ZN(P3_U3233) );
  INV_X1 U12897 ( .A(n10289), .ZN(n10291) );
  NAND2_X1 U12898 ( .A1(n10291), .A2(n10290), .ZN(n10292) );
  NOR2_X1 U12899 ( .A1(n10293), .A2(n10292), .ZN(n10294) );
  AND2_X1 U12900 ( .A1(n10294), .A2(n10873), .ZN(n10319) );
  INV_X1 U12901 ( .A(n10318), .ZN(n10874) );
  INV_X1 U12902 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10317) );
  OR2_X1 U12903 ( .A1(n10351), .A2(n10918), .ZN(n10346) );
  OAI21_X1 U12904 ( .B1(n10296), .B2(n10307), .A(n10886), .ZN(n14576) );
  INV_X1 U12905 ( .A(n14576), .ZN(n10315) );
  NAND2_X1 U12906 ( .A1(n11825), .A2(n10878), .ZN(n10297) );
  INV_X1 U12907 ( .A(n10298), .ZN(n10300) );
  NOR2_X1 U12908 ( .A1(n10300), .A2(n10299), .ZN(n10301) );
  NOR2_X1 U12909 ( .A1(n10301), .A2(n11318), .ZN(n10914) );
  NAND2_X1 U12910 ( .A1(n10914), .A2(n13685), .ZN(n14551) );
  NAND2_X1 U12911 ( .A1(n10152), .A2(n10976), .ZN(n10305) );
  NAND2_X1 U12912 ( .A1(n10306), .A2(n10305), .ZN(n10863) );
  XNOR2_X1 U12913 ( .A(n10863), .B(n10307), .ZN(n10311) );
  OAI21_X1 U12914 ( .B1(n10311), .B2(n14666), .A(n10310), .ZN(n10312) );
  AOI21_X1 U12915 ( .B1(n14639), .B2(n14576), .A(n10312), .ZN(n14579) );
  NAND2_X1 U12916 ( .A1(n10918), .A2(n12178), .ZN(n10357) );
  AOI211_X1 U12917 ( .C1(n10313), .C2(n10357), .A(n13903), .B(n11086), .ZN(
        n14568) );
  AOI21_X1 U12918 ( .B1(n14632), .B2(n10313), .A(n14568), .ZN(n10314) );
  OAI211_X1 U12919 ( .C1(n10315), .C2(n14636), .A(n14579), .B(n10314), .ZN(
        n10320) );
  NAND2_X1 U12920 ( .A1(n10320), .A2(n14675), .ZN(n10316) );
  OAI21_X1 U12921 ( .B1(n14675), .B2(n10317), .A(n10316), .ZN(P1_U3465) );
  NAND2_X1 U12922 ( .A1(n10320), .A2(n14688), .ZN(n10321) );
  OAI21_X1 U12923 ( .B1(n14688), .B2(n10131), .A(n10321), .ZN(P1_U3530) );
  INV_X1 U12924 ( .A(P3_DATAO_REG_25__SCAN_IN), .ZN(n15407) );
  NAND2_X1 U12925 ( .A1(n12373), .A2(P3_U3897), .ZN(n10322) );
  OAI21_X1 U12926 ( .B1(P3_U3897), .B2(n15407), .A(n10322), .ZN(P3_U3516) );
  INV_X1 U12927 ( .A(n10323), .ZN(n10324) );
  OAI222_X1 U12928 ( .A1(P3_U3151), .A2(n10326), .B1(n12787), .B2(n10325), 
        .C1(n12785), .C2(n10324), .ZN(P3_U3275) );
  AND2_X1 U12929 ( .A1(P2_U3088), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n10327) );
  AOI21_X1 U12930 ( .B1(n14825), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n10327), 
        .ZN(n10328) );
  INV_X1 U12931 ( .A(n10328), .ZN(n10334) );
  AOI21_X1 U12932 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n10335), .A(n10329), 
        .ZN(n10332) );
  INV_X1 U12933 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n10330) );
  MUX2_X1 U12934 ( .A(n10330), .B(P2_REG1_REG_14__SCAN_IN), .S(n10732), .Z(
        n10331) );
  NOR2_X1 U12935 ( .A1(n10332), .A2(n10331), .ZN(n10731) );
  AOI211_X1 U12936 ( .C1(n10332), .C2(n10331), .A(n10731), .B(n14819), .ZN(
        n10333) );
  AOI211_X1 U12937 ( .C1(n14809), .C2(n10732), .A(n10334), .B(n10333), .ZN(
        n10343) );
  NAND2_X1 U12938 ( .A1(n10335), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n10340) );
  INV_X1 U12939 ( .A(n10336), .ZN(n10337) );
  NAND2_X1 U12940 ( .A1(n10338), .A2(n10337), .ZN(n10339) );
  NAND2_X1 U12941 ( .A1(n10340), .A2(n10339), .ZN(n10726) );
  XOR2_X1 U12942 ( .A(n10732), .B(n10726), .Z(n10341) );
  NAND2_X1 U12943 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n10341), .ZN(n10727) );
  OAI211_X1 U12944 ( .C1(n10341), .C2(P2_REG2_REG_14__SCAN_IN), .A(n14811), 
        .B(n10727), .ZN(n10342) );
  NAND2_X1 U12945 ( .A1(n10343), .A2(n10342), .ZN(P2_U3228) );
  INV_X1 U12946 ( .A(n10344), .ZN(n10396) );
  AOI22_X1 U12947 ( .A1(n14493), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n11525), .ZN(n10345) );
  OAI21_X1 U12948 ( .B1(n10396), .B2(n10724), .A(n10345), .ZN(P1_U3339) );
  INV_X1 U12949 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n15347) );
  INV_X1 U12950 ( .A(n10346), .ZN(n10348) );
  NAND2_X1 U12951 ( .A1(n10348), .A2(n10347), .ZN(n10349) );
  NAND2_X1 U12952 ( .A1(n10350), .A2(n10349), .ZN(n10981) );
  INV_X1 U12953 ( .A(n10981), .ZN(n10360) );
  NOR2_X1 U12954 ( .A1(n10144), .A2(n14539), .ZN(n10356) );
  OAI21_X1 U12955 ( .B1(n10353), .B2(n10351), .A(n14554), .ZN(n10354) );
  OAI21_X1 U12956 ( .B1(n10353), .B2(n10365), .A(n14554), .ZN(n10352) );
  AOI222_X1 U12957 ( .A1(n10354), .A2(n14537), .B1(n10353), .B2(n10304), .C1(
        n10352), .C2(n10351), .ZN(n10355) );
  AOI211_X1 U12958 ( .C1(n14639), .C2(n10981), .A(n10356), .B(n10355), .ZN(
        n10983) );
  OAI211_X1 U12959 ( .C1(n10918), .C2(n12178), .A(n14561), .B(n10357), .ZN(
        n10358) );
  INV_X1 U12960 ( .A(n10358), .ZN(n10975) );
  AOI21_X1 U12961 ( .B1(n14632), .B2(n10976), .A(n10975), .ZN(n10359) );
  OAI211_X1 U12962 ( .C1(n10360), .C2(n14636), .A(n10983), .B(n10359), .ZN(
        n14019) );
  NAND2_X1 U12963 ( .A1(n14019), .A2(n14675), .ZN(n10361) );
  OAI21_X1 U12964 ( .B1(n14675), .B2(n15347), .A(n10361), .ZN(P1_U3462) );
  OR2_X1 U12965 ( .A1(n10152), .A2(n14539), .ZN(n10912) );
  INV_X1 U12966 ( .A(n10912), .ZN(n10364) );
  INV_X1 U12967 ( .A(n10915), .ZN(n10362) );
  AOI21_X1 U12968 ( .B1(n14018), .B2(n14666), .A(n10362), .ZN(n10363) );
  AOI211_X1 U12969 ( .C1(n10365), .C2(n10012), .A(n10364), .B(n10363), .ZN(
        n14608) );
  NAND2_X1 U12970 ( .A1(n14686), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10366) );
  OAI21_X1 U12971 ( .B1(n14608), .B2(n14686), .A(n10366), .ZN(P1_U3528) );
  INV_X1 U12972 ( .A(n10367), .ZN(n10412) );
  AOI22_X1 U12973 ( .A1(n14453), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n11525), .ZN(n10368) );
  OAI21_X1 U12974 ( .B1(n10412), .B2(n10724), .A(n10368), .ZN(P1_U3341) );
  XNOR2_X1 U12975 ( .A(n10369), .B(n10372), .ZN(n10494) );
  OAI21_X1 U12976 ( .B1(n10370), .B2(n10378), .A(n14313), .ZN(n10371) );
  NOR2_X1 U12977 ( .A1(n10371), .A2(n10403), .ZN(n10487) );
  XNOR2_X1 U12978 ( .A(n10373), .B(n10372), .ZN(n10375) );
  OAI21_X1 U12979 ( .B1(n10375), .B2(n13171), .A(n10374), .ZN(n10491) );
  AOI211_X1 U12980 ( .C1(n10494), .C2(n14905), .A(n10487), .B(n10491), .ZN(
        n10381) );
  AOI22_X1 U12981 ( .A1(n13304), .A2(n11870), .B1(n14932), .B2(
        P2_REG1_REG_4__SCAN_IN), .ZN(n10376) );
  OAI21_X1 U12982 ( .B1(n10381), .B2(n14932), .A(n10376), .ZN(P2_U3503) );
  INV_X1 U12983 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10377) );
  OAI22_X1 U12984 ( .A1(n13329), .A2(n10378), .B1(n14924), .B2(n10377), .ZN(
        n10379) );
  INV_X1 U12985 ( .A(n10379), .ZN(n10380) );
  OAI21_X1 U12986 ( .B1(n10381), .B2(n14922), .A(n10380), .ZN(P2_U3442) );
  XNOR2_X1 U12987 ( .A(n10382), .B(n11723), .ZN(n15144) );
  INV_X1 U12988 ( .A(n15144), .ZN(n10395) );
  NOR2_X1 U12989 ( .A1(n15126), .A2(n11559), .ZN(n10383) );
  AOI21_X1 U12990 ( .B1(n10590), .B2(n10385), .A(n10384), .ZN(n10390) );
  NAND2_X1 U12991 ( .A1(n10386), .A2(n15122), .ZN(n10389) );
  NAND2_X1 U12992 ( .A1(n15144), .A2(n11379), .ZN(n10388) );
  AOI22_X1 U12993 ( .A1(n12408), .A2(n12374), .B1(n12375), .B2(n12406), .ZN(
        n10387) );
  OAI211_X1 U12994 ( .C1(n10390), .C2(n10389), .A(n10388), .B(n10387), .ZN(
        n15142) );
  MUX2_X1 U12995 ( .A(P3_REG2_REG_3__SCAN_IN), .B(n15142), .S(n15131), .Z(
        n10391) );
  INV_X1 U12996 ( .A(n10391), .ZN(n10394) );
  NOR2_X1 U12997 ( .A1(n11578), .A2(n15146), .ZN(n15143) );
  AOI22_X1 U12998 ( .A1(n14276), .A2(n15143), .B1(n15591), .B2(n8577), .ZN(
        n10393) );
  OAI211_X1 U12999 ( .C1(n10395), .C2(n12576), .A(n10394), .B(n10393), .ZN(
        P3_U3230) );
  OAI222_X1 U13000 ( .A1(P2_U3088), .A2(n14801), .B1(n13359), .B2(n10396), 
        .C1(n15311), .C2(n13357), .ZN(P2_U3311) );
  XNOR2_X1 U13001 ( .A(n10397), .B(n10398), .ZN(n14899) );
  XNOR2_X1 U13002 ( .A(n10399), .B(n10398), .ZN(n10401) );
  AOI21_X1 U13003 ( .B1(n10401), .B2(n14304), .A(n10400), .ZN(n14902) );
  MUX2_X1 U13004 ( .A(n10402), .B(n14902), .S(n14837), .Z(n10410) );
  OAI21_X1 U13005 ( .B1(n10403), .B2(n14901), .A(n14313), .ZN(n10404) );
  OR2_X1 U13006 ( .A1(n10606), .A2(n10404), .ZN(n14900) );
  INV_X1 U13007 ( .A(n14900), .ZN(n10408) );
  INV_X1 U13008 ( .A(n10405), .ZN(n10406) );
  OAI22_X1 U13009 ( .A1(n14835), .A2(n14901), .B1(n13194), .B2(n10406), .ZN(
        n10407) );
  AOI21_X1 U13010 ( .B1(n10408), .B2(n14315), .A(n10407), .ZN(n10409) );
  OAI211_X1 U13011 ( .C1(n13182), .C2(n14899), .A(n10410), .B(n10409), .ZN(
        P2_U3260) );
  INV_X1 U13012 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10413) );
  INV_X1 U13013 ( .A(n10732), .ZN(n10411) );
  OAI222_X1 U13014 ( .A1(n13357), .A2(n10413), .B1(n13359), .B2(n10412), .C1(
        n10411), .C2(P2_U3088), .ZN(P2_U3313) );
  INV_X1 U13015 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n15414) );
  AOI22_X1 U13016 ( .A1(n13671), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n15414), 
        .B2(n10422), .ZN(n10417) );
  INV_X1 U13017 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10415) );
  MUX2_X1 U13018 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10415), .S(n10426), .Z(
        n14429) );
  NAND2_X1 U13019 ( .A1(n14430), .A2(n14429), .ZN(n14428) );
  OAI21_X1 U13020 ( .B1(n10417), .B2(n10416), .A(n13670), .ZN(n10421) );
  NAND2_X1 U13021 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n11327)
         );
  NAND2_X1 U13022 ( .A1(n10418), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n10419) );
  OAI211_X1 U13023 ( .C1(n14525), .C2(n10422), .A(n11327), .B(n10419), .ZN(
        n10420) );
  AOI21_X1 U13024 ( .B1(n10421), .B2(n14517), .A(n10420), .ZN(n10431) );
  INV_X1 U13025 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n15491) );
  AOI22_X1 U13026 ( .A1(n13671), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n15491), 
        .B2(n10422), .ZN(n10428) );
  INV_X1 U13027 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10425) );
  MUX2_X1 U13028 ( .A(n10425), .B(P1_REG2_REG_11__SCAN_IN), .S(n10426), .Z(
        n14433) );
  AOI21_X1 U13029 ( .B1(n10426), .B2(P1_REG2_REG_11__SCAN_IN), .A(n14432), 
        .ZN(n10427) );
  NAND2_X1 U13030 ( .A1(n10428), .A2(n10427), .ZN(n13659) );
  OAI21_X1 U13031 ( .B1(n10428), .B2(n10427), .A(n13659), .ZN(n10429) );
  NAND2_X1 U13032 ( .A1(n10429), .A2(n14521), .ZN(n10430) );
  NAND2_X1 U13033 ( .A1(n10431), .A2(n10430), .ZN(P1_U3255) );
  INV_X1 U13034 ( .A(n10432), .ZN(n10434) );
  OAI222_X1 U13035 ( .A1(n11559), .A2(P3_U3151), .B1(n12785), .B2(n10434), 
        .C1(n10433), .C2(n12787), .ZN(P3_U3274) );
  XNOR2_X1 U13036 ( .A(n15147), .B(n12273), .ZN(n10560) );
  XNOR2_X1 U13037 ( .A(n10560), .B(n12406), .ZN(n10444) );
  INV_X1 U13038 ( .A(n10435), .ZN(n10436) );
  AND2_X1 U13039 ( .A1(n10436), .A2(n15118), .ZN(n10437) );
  XNOR2_X1 U13040 ( .A(n12258), .B(n12220), .ZN(n10440) );
  XNOR2_X1 U13041 ( .A(n10440), .B(n10587), .ZN(n12256) );
  NAND2_X1 U13042 ( .A1(n12257), .A2(n12256), .ZN(n12255) );
  NAND2_X1 U13043 ( .A1(n12407), .A2(n10440), .ZN(n10441) );
  NAND2_X1 U13044 ( .A1(n12255), .A2(n10441), .ZN(n10443) );
  INV_X1 U13045 ( .A(n10564), .ZN(n10442) );
  AOI21_X1 U13046 ( .B1(n10444), .B2(n10443), .A(n10442), .ZN(n10449) );
  OAI21_X1 U13047 ( .B1(n12352), .B2(n15147), .A(n10445), .ZN(n10446) );
  AOI21_X1 U13048 ( .B1(n12289), .B2(n12405), .A(n10446), .ZN(n10448) );
  AOI22_X1 U13049 ( .A1(n12407), .A2(n12291), .B1(n10513), .B2(n12376), .ZN(
        n10447) );
  OAI211_X1 U13050 ( .C1(n10449), .C2(n12382), .A(n10448), .B(n10447), .ZN(
        P3_U3170) );
  NAND3_X1 U13051 ( .A1(n10452), .A2(n10451), .A3(n10450), .ZN(n10453) );
  NAND2_X1 U13052 ( .A1(n10453), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10454) );
  NOR2_X1 U13053 ( .A1(n13546), .A2(n14537), .ZN(n13568) );
  INV_X1 U13054 ( .A(n13568), .ZN(n13493) );
  NAND2_X1 U13055 ( .A1(n14358), .A2(n11088), .ZN(n10457) );
  OAI22_X1 U13056 ( .A1(n13571), .A2(n11092), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11087), .ZN(n10455) );
  INV_X1 U13057 ( .A(n10455), .ZN(n10456) );
  OAI211_X1 U13058 ( .C1(n10144), .C2(n13493), .A(n10457), .B(n10456), .ZN(
        n10474) );
  NAND2_X1 U13059 ( .A1(n13597), .A2(n10014), .ZN(n10459) );
  INV_X2 U13060 ( .A(n13393), .ZN(n13475) );
  NAND2_X1 U13061 ( .A1(n11088), .A2(n13475), .ZN(n10458) );
  NAND2_X1 U13062 ( .A1(n10459), .A2(n10458), .ZN(n10460) );
  XNOR2_X1 U13063 ( .A(n10460), .B(n11318), .ZN(n10542) );
  INV_X2 U13064 ( .A(n13405), .ZN(n13478) );
  AND2_X1 U13065 ( .A1(n10014), .A2(n11088), .ZN(n10461) );
  AOI21_X1 U13066 ( .B1(n13478), .B2(n13597), .A(n10461), .ZN(n10543) );
  XNOR2_X1 U13067 ( .A(n10542), .B(n10543), .ZN(n10472) );
  INV_X1 U13068 ( .A(n10462), .ZN(n10464) );
  OR2_X1 U13069 ( .A1(n10464), .A2(n10463), .ZN(n10465) );
  INV_X1 U13070 ( .A(n10467), .ZN(n10469) );
  INV_X1 U13071 ( .A(n10470), .ZN(n10471) );
  AOI211_X1 U13072 ( .C1(n10472), .C2(n10467), .A(n13564), .B(n10471), .ZN(
        n10473) );
  AOI211_X1 U13073 ( .C1(n11087), .C2(n13573), .A(n10474), .B(n10473), .ZN(
        n10475) );
  INV_X1 U13074 ( .A(n10475), .ZN(P1_U3218) );
  XNOR2_X1 U13075 ( .A(n11884), .B(n9889), .ZN(n10525) );
  NAND2_X1 U13076 ( .A1(n12939), .A2(n12126), .ZN(n10526) );
  XNOR2_X1 U13077 ( .A(n10525), .B(n10526), .ZN(n10530) );
  NAND2_X1 U13078 ( .A1(n10477), .A2(n10476), .ZN(n10531) );
  XOR2_X1 U13079 ( .A(n10530), .B(n10531), .Z(n10485) );
  NOR2_X1 U13080 ( .A1(n12900), .A2(n10611), .ZN(n10484) );
  INV_X1 U13081 ( .A(n10478), .ZN(n10610) );
  NAND2_X1 U13082 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n14724) );
  NAND2_X1 U13083 ( .A1(n12938), .A2(n12902), .ZN(n10480) );
  NAND2_X1 U13084 ( .A1(n12940), .A2(n12901), .ZN(n10479) );
  AND2_X1 U13085 ( .A1(n10480), .A2(n10479), .ZN(n10602) );
  INV_X1 U13086 ( .A(n10602), .ZN(n10481) );
  NAND2_X1 U13087 ( .A1(n10481), .A2(n12897), .ZN(n10482) );
  OAI211_X1 U13088 ( .C1(n12894), .C2(n10610), .A(n14724), .B(n10482), .ZN(
        n10483) );
  AOI211_X1 U13089 ( .C1(n10485), .C2(n12887), .A(n10484), .B(n10483), .ZN(
        n10486) );
  INV_X1 U13090 ( .A(n10486), .ZN(P2_U3211) );
  INV_X1 U13091 ( .A(n10487), .ZN(n10490) );
  AOI22_X1 U13092 ( .A1(n14307), .A2(n11870), .B1(n14841), .B2(n10488), .ZN(
        n10489) );
  OAI21_X1 U13093 ( .B1(n10490), .B2(n13213), .A(n10489), .ZN(n10493) );
  MUX2_X1 U13094 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n10491), .S(n14837), .Z(
        n10492) );
  AOI211_X1 U13095 ( .C1(n14316), .C2(n10494), .A(n10493), .B(n10492), .ZN(
        n10495) );
  INV_X1 U13096 ( .A(n10495), .ZN(P2_U3261) );
  INV_X1 U13097 ( .A(n10496), .ZN(n10501) );
  NOR2_X1 U13098 ( .A1(n13213), .A2(n10497), .ZN(n10500) );
  AOI22_X1 U13099 ( .A1(n13216), .A2(P2_REG2_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(n14841), .ZN(n10498) );
  OAI21_X1 U13100 ( .B1(n14835), .B2(n7215), .A(n10498), .ZN(n10499) );
  AOI211_X1 U13101 ( .C1(n10501), .C2(n14316), .A(n10500), .B(n10499), .ZN(
        n10502) );
  OAI21_X1 U13102 ( .B1(n13211), .B2(n10503), .A(n10502), .ZN(P2_U3264) );
  OR2_X1 U13103 ( .A1(n10504), .A2(n11580), .ZN(n10505) );
  NAND2_X1 U13104 ( .A1(n10506), .A2(n10505), .ZN(n15150) );
  INV_X1 U13105 ( .A(n15150), .ZN(n10517) );
  XNOR2_X1 U13106 ( .A(n10507), .B(n11729), .ZN(n10511) );
  NAND2_X1 U13107 ( .A1(n15150), .A2(n11379), .ZN(n10510) );
  OAI22_X1 U13108 ( .A1(n10587), .A2(n15119), .B1(n10742), .B2(n15117), .ZN(
        n10508) );
  INV_X1 U13109 ( .A(n10508), .ZN(n10509) );
  OAI211_X1 U13110 ( .C1(n10511), .C2(n14264), .A(n10510), .B(n10509), .ZN(
        n15148) );
  MUX2_X1 U13111 ( .A(P3_REG2_REG_4__SCAN_IN), .B(n15148), .S(n15131), .Z(
        n10512) );
  INV_X1 U13112 ( .A(n10512), .ZN(n10516) );
  AOI22_X1 U13113 ( .A1(n12640), .A2(n10514), .B1(n15591), .B2(n10513), .ZN(
        n10515) );
  OAI211_X1 U13114 ( .C1(n10517), .C2(n12576), .A(n10516), .B(n10515), .ZN(
        P3_U3229) );
  INV_X1 U13115 ( .A(n10518), .ZN(n10520) );
  OAI222_X1 U13116 ( .A1(n14039), .A2(n10519), .B1(n10724), .B2(n10520), .C1(
        n14478), .C2(P1_U3086), .ZN(P1_U3340) );
  INV_X1 U13117 ( .A(n12970), .ZN(n12959) );
  OAI222_X1 U13118 ( .A1(n13357), .A2(n10521), .B1(n13359), .B2(n10520), .C1(
        n12959), .C2(P2_U3088), .ZN(P2_U3312) );
  INV_X1 U13119 ( .A(n10522), .ZN(n10523) );
  INV_X1 U13120 ( .A(n13676), .ZN(n14508) );
  OAI222_X1 U13121 ( .A1(n14039), .A2(n15494), .B1(n10724), .B2(n10523), .C1(
        n14508), .C2(P1_U3086), .ZN(P1_U3338) );
  INV_X1 U13122 ( .A(n14808), .ZN(n12973) );
  OAI222_X1 U13123 ( .A1(n13357), .A2(n10524), .B1(n13359), .B2(n10523), .C1(
        n12973), .C2(P2_U3088), .ZN(P2_U3310) );
  INV_X1 U13124 ( .A(n10525), .ZN(n10528) );
  INV_X1 U13125 ( .A(n10526), .ZN(n10527) );
  NAND2_X1 U13126 ( .A1(n10528), .A2(n10527), .ZN(n10529) );
  XNOR2_X1 U13127 ( .A(n11890), .B(n12154), .ZN(n10682) );
  NAND2_X1 U13128 ( .A1(n12938), .A2(n12126), .ZN(n10680) );
  XNOR2_X1 U13129 ( .A(n10682), .B(n10680), .ZN(n10684) );
  XNOR2_X1 U13130 ( .A(n10685), .B(n10684), .ZN(n10538) );
  NAND2_X1 U13131 ( .A1(n12937), .A2(n12902), .ZN(n10534) );
  NAND2_X1 U13132 ( .A1(n12939), .A2(n12901), .ZN(n10533) );
  AND2_X1 U13133 ( .A1(n10534), .A2(n10533), .ZN(n10573) );
  NAND2_X1 U13134 ( .A1(n12903), .A2(n10577), .ZN(n10535) );
  NAND2_X1 U13135 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n12945) );
  OAI211_X1 U13136 ( .C1(n10573), .C2(n12906), .A(n10535), .B(n12945), .ZN(
        n10536) );
  AOI21_X1 U13137 ( .B1(n11890), .B2(n12913), .A(n10536), .ZN(n10537) );
  OAI21_X1 U13138 ( .B1(n10538), .B2(n12908), .A(n10537), .ZN(P2_U3185) );
  INV_X1 U13139 ( .A(n10539), .ZN(n10541) );
  OAI22_X1 U13140 ( .A1(n11756), .A2(P3_U3151), .B1(SI_22_), .B2(n12787), .ZN(
        n10540) );
  AOI21_X1 U13141 ( .B1(n10541), .B2(n12775), .A(n10540), .ZN(P3_U3273) );
  INV_X1 U13142 ( .A(n10542), .ZN(n10545) );
  INV_X1 U13143 ( .A(n10543), .ZN(n10544) );
  NAND2_X1 U13144 ( .A1(n10545), .A2(n10544), .ZN(n10546) );
  OAI22_X1 U13145 ( .A1(n11092), .A2(n13405), .B1(n10889), .B2(n13407), .ZN(
        n10549) );
  INV_X1 U13146 ( .A(n10549), .ZN(n10548) );
  NAND2_X1 U13147 ( .A1(n10658), .A2(n10655), .ZN(n10552) );
  OAI22_X1 U13148 ( .A1(n11092), .A2(n13407), .B1(n10889), .B2(n6962), .ZN(
        n10551) );
  XNOR2_X1 U13149 ( .A(n10551), .B(n11318), .ZN(n10654) );
  XNOR2_X1 U13150 ( .A(n10552), .B(n10654), .ZN(n10558) );
  INV_X1 U13151 ( .A(n11017), .ZN(n10641) );
  NAND2_X1 U13152 ( .A1(n11072), .A2(n14632), .ZN(n14617) );
  NAND2_X1 U13153 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n13642) );
  NAND2_X1 U13154 ( .A1(n13597), .A2(n13854), .ZN(n10554) );
  NAND2_X1 U13155 ( .A1(n13596), .A2(n13913), .ZN(n10553) );
  NAND2_X1 U13156 ( .A1(n10554), .A2(n10553), .ZN(n11077) );
  NAND2_X1 U13157 ( .A1(n11077), .A2(n14359), .ZN(n10555) );
  OAI211_X1 U13158 ( .C1(n10641), .C2(n14617), .A(n13642), .B(n10555), .ZN(
        n10556) );
  AOI21_X1 U13159 ( .B1(n11068), .B2(n13573), .A(n10556), .ZN(n10557) );
  OAI21_X1 U13160 ( .B1(n10558), .B2(n13564), .A(n10557), .ZN(P1_U3230) );
  XNOR2_X1 U13161 ( .A(n10559), .B(n12220), .ZN(n10741) );
  XNOR2_X1 U13162 ( .A(n10741), .B(n10742), .ZN(n10739) );
  INV_X1 U13163 ( .A(n10560), .ZN(n10561) );
  NAND2_X1 U13164 ( .A1(n10562), .A2(n10561), .ZN(n10563) );
  XOR2_X1 U13165 ( .A(n10739), .B(n10740), .Z(n10568) );
  OAI22_X1 U13166 ( .A1(n12352), .A2(n10626), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15315), .ZN(n10565) );
  AOI21_X1 U13167 ( .B1(n12289), .B2(n12404), .A(n10565), .ZN(n10567) );
  AOI22_X1 U13168 ( .A1(n12291), .A2(n12406), .B1(n10627), .B2(n12376), .ZN(
        n10566) );
  OAI211_X1 U13169 ( .C1(n10568), .C2(n12382), .A(n10567), .B(n10566), .ZN(
        P3_U3167) );
  OAI21_X1 U13170 ( .B1(n10570), .B2(n10571), .A(n10569), .ZN(n10719) );
  INV_X1 U13171 ( .A(n10719), .ZN(n10583) );
  XNOR2_X1 U13172 ( .A(n10572), .B(n10571), .ZN(n10574) );
  OAI21_X1 U13173 ( .B1(n10574), .B2(n13171), .A(n10573), .ZN(n10717) );
  NAND2_X1 U13174 ( .A1(n10717), .A2(n14837), .ZN(n10582) );
  INV_X1 U13175 ( .A(n10575), .ZN(n10988) );
  AOI211_X1 U13176 ( .C1(n11890), .C2(n10607), .A(n13049), .B(n10988), .ZN(
        n10718) );
  INV_X1 U13177 ( .A(n11890), .ZN(n10576) );
  NOR2_X1 U13178 ( .A1(n10576), .A2(n14835), .ZN(n10580) );
  INV_X1 U13179 ( .A(n10577), .ZN(n10578) );
  OAI22_X1 U13180 ( .A1(n14837), .A2(n9770), .B1(n10578), .B2(n13194), .ZN(
        n10579) );
  AOI211_X1 U13181 ( .C1(n10718), .C2(n14315), .A(n10580), .B(n10579), .ZN(
        n10581) );
  OAI211_X1 U13182 ( .C1(n10583), .C2(n13182), .A(n10582), .B(n10581), .ZN(
        P2_U3258) );
  INV_X1 U13183 ( .A(n12576), .ZN(n15128) );
  OAI21_X1 U13184 ( .B1(n10585), .B2(n11719), .A(n10584), .ZN(n15140) );
  OAI22_X1 U13185 ( .A1(n10587), .A2(n15117), .B1(n10586), .B2(n15119), .ZN(
        n10592) );
  NAND3_X1 U13186 ( .A1(n15114), .A2(n11719), .A3(n10588), .ZN(n10589) );
  AOI21_X1 U13187 ( .B1(n10590), .B2(n10589), .A(n14264), .ZN(n10591) );
  AOI211_X1 U13188 ( .C1(n11379), .C2(n15140), .A(n10592), .B(n10591), .ZN(
        n15137) );
  NOR2_X1 U13189 ( .A1(n10593), .A2(n15146), .ZN(n15139) );
  AOI22_X1 U13190 ( .A1(n15139), .A2(n15126), .B1(P3_REG3_REG_2__SCAN_IN), 
        .B2(n15591), .ZN(n10594) );
  NAND2_X1 U13191 ( .A1(n15137), .A2(n10594), .ZN(n10595) );
  MUX2_X1 U13192 ( .A(P3_REG2_REG_2__SCAN_IN), .B(n10595), .S(n15131), .Z(
        n10596) );
  AOI21_X1 U13193 ( .B1(n15128), .B2(n15140), .A(n10596), .ZN(n10597) );
  INV_X1 U13194 ( .A(n10597), .ZN(P3_U3231) );
  INV_X1 U13195 ( .A(n10598), .ZN(n10600) );
  OAI21_X1 U13196 ( .B1(n10600), .B2(n7431), .A(n10599), .ZN(n10650) );
  INV_X1 U13197 ( .A(n10650), .ZN(n10615) );
  XOR2_X1 U13198 ( .A(n10601), .B(n12075), .Z(n10603) );
  OAI21_X1 U13199 ( .B1(n10603), .B2(n13171), .A(n10602), .ZN(n10648) );
  INV_X1 U13200 ( .A(n10648), .ZN(n10604) );
  MUX2_X1 U13201 ( .A(n10605), .B(n10604), .S(n14837), .Z(n10614) );
  INV_X1 U13202 ( .A(n10606), .ZN(n10609) );
  INV_X1 U13203 ( .A(n10607), .ZN(n10608) );
  AOI211_X1 U13204 ( .C1(n11884), .C2(n10609), .A(n13049), .B(n10608), .ZN(
        n10649) );
  OAI22_X1 U13205 ( .A1(n14835), .A2(n10611), .B1(n13194), .B2(n10610), .ZN(
        n10612) );
  AOI21_X1 U13206 ( .B1(n10649), .B2(n14315), .A(n10612), .ZN(n10613) );
  OAI211_X1 U13207 ( .C1(n13182), .C2(n10615), .A(n10614), .B(n10613), .ZN(
        P2_U3259) );
  NAND2_X1 U13208 ( .A1(n12410), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n10616) );
  OAI21_X1 U13209 ( .B1(n11554), .B2(n12410), .A(n10616), .ZN(P3_U3521) );
  XNOR2_X1 U13210 ( .A(n10617), .B(n11721), .ZN(n15155) );
  INV_X1 U13211 ( .A(n15155), .ZN(n10630) );
  INV_X1 U13212 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n10625) );
  NAND2_X1 U13213 ( .A1(n15155), .A2(n11379), .ZN(n10624) );
  NAND2_X1 U13214 ( .A1(n10618), .A2(n11721), .ZN(n10619) );
  NAND2_X1 U13215 ( .A1(n10706), .A2(n10619), .ZN(n10622) );
  NAND2_X1 U13216 ( .A1(n12406), .A2(n12374), .ZN(n10620) );
  OAI21_X1 U13217 ( .B1(n10785), .B2(n15117), .A(n10620), .ZN(n10621) );
  AOI21_X1 U13218 ( .B1(n10622), .B2(n15122), .A(n10621), .ZN(n10623) );
  AND2_X1 U13219 ( .A1(n10624), .A2(n10623), .ZN(n15152) );
  MUX2_X1 U13220 ( .A(n10625), .B(n15152), .S(n15131), .Z(n10629) );
  NOR2_X1 U13221 ( .A1(n10626), .A2(n15146), .ZN(n15154) );
  AOI22_X1 U13222 ( .A1(n14276), .A2(n15154), .B1(n15591), .B2(n10627), .ZN(
        n10628) );
  OAI211_X1 U13223 ( .C1(n10630), .C2(n12576), .A(n10629), .B(n10628), .ZN(
        P3_U3228) );
  INV_X1 U13224 ( .A(n10658), .ZN(n10631) );
  OAI21_X1 U13225 ( .B1(n10631), .B2(n10654), .A(n10655), .ZN(n10637) );
  NAND2_X1 U13226 ( .A1(n13596), .A2(n10014), .ZN(n10633) );
  NAND2_X1 U13227 ( .A1(n10899), .A2(n13475), .ZN(n10632) );
  NAND2_X1 U13228 ( .A1(n10633), .A2(n10632), .ZN(n10634) );
  XNOR2_X1 U13229 ( .A(n10634), .B(n11318), .ZN(n10659) );
  AND2_X1 U13230 ( .A1(n13445), .A2(n10899), .ZN(n10635) );
  AOI21_X1 U13231 ( .B1(n13478), .B2(n13596), .A(n10635), .ZN(n10656) );
  INV_X1 U13232 ( .A(n10656), .ZN(n10660) );
  XNOR2_X1 U13233 ( .A(n10659), .B(n10660), .ZN(n10636) );
  XNOR2_X1 U13234 ( .A(n10637), .B(n10636), .ZN(n10644) );
  NAND2_X1 U13235 ( .A1(n14632), .A2(n10899), .ZN(n14625) );
  OR2_X1 U13236 ( .A1(n11092), .A2(n14537), .ZN(n10639) );
  NAND2_X1 U13237 ( .A1(n13595), .A2(n13913), .ZN(n10638) );
  NAND2_X1 U13238 ( .A1(n10639), .A2(n10638), .ZN(n10869) );
  AOI22_X1 U13239 ( .A1(n10869), .A2(n14359), .B1(P1_REG3_REG_5__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10640) );
  OAI21_X1 U13240 ( .B1(n10641), .B2(n14625), .A(n10640), .ZN(n10642) );
  AOI21_X1 U13241 ( .B1(n10881), .B2(n13573), .A(n10642), .ZN(n10643) );
  OAI21_X1 U13242 ( .B1(n10644), .B2(n13564), .A(n10643), .ZN(P1_U3227) );
  NAND2_X1 U13243 ( .A1(n10645), .A2(n12775), .ZN(n10646) );
  OAI211_X1 U13244 ( .C1(n10647), .C2(n12787), .A(n10646), .B(n11759), .ZN(
        P3_U3272) );
  AOI211_X1 U13245 ( .C1(n14905), .C2(n10650), .A(n10649), .B(n10648), .ZN(
        n10653) );
  AOI22_X1 U13246 ( .A1(n8982), .A2(n11884), .B1(n14922), .B2(
        P2_REG0_REG_6__SCAN_IN), .ZN(n10651) );
  OAI21_X1 U13247 ( .B1(n10653), .B2(n14922), .A(n10651), .ZN(P2_U3448) );
  AOI22_X1 U13248 ( .A1(n13304), .A2(n11884), .B1(n14932), .B2(
        P2_REG1_REG_6__SCAN_IN), .ZN(n10652) );
  OAI21_X1 U13249 ( .B1(n10653), .B2(n14932), .A(n10652), .ZN(P2_U3505) );
  NAND2_X1 U13250 ( .A1(n10659), .A2(n10656), .ZN(n10657) );
  INV_X1 U13251 ( .A(n10659), .ZN(n10661) );
  NAND2_X1 U13252 ( .A1(n10661), .A2(n10660), .ZN(n10662) );
  NAND2_X1 U13253 ( .A1(n13595), .A2(n13445), .ZN(n10664) );
  NAND2_X1 U13254 ( .A1(n14631), .A2(n13475), .ZN(n10663) );
  NAND2_X1 U13255 ( .A1(n10664), .A2(n10663), .ZN(n10665) );
  XNOR2_X1 U13256 ( .A(n10665), .B(n11318), .ZN(n10669) );
  INV_X1 U13257 ( .A(n10669), .ZN(n10667) );
  AOI22_X1 U13258 ( .A1(n13478), .A2(n13595), .B1(n13445), .B2(n14631), .ZN(
        n10668) );
  INV_X1 U13259 ( .A(n10668), .ZN(n10666) );
  NAND2_X1 U13260 ( .A1(n10667), .A2(n10666), .ZN(n10753) );
  INV_X1 U13261 ( .A(n10753), .ZN(n10670) );
  AND2_X1 U13262 ( .A1(n10669), .A2(n10668), .ZN(n10752) );
  NOR2_X1 U13263 ( .A1(n10670), .A2(n10752), .ZN(n10671) );
  XNOR2_X1 U13264 ( .A(n10754), .B(n10671), .ZN(n10678) );
  INV_X1 U13265 ( .A(n10672), .ZN(n10907) );
  NAND2_X1 U13266 ( .A1(n13596), .A2(n13854), .ZN(n10674) );
  NAND2_X1 U13267 ( .A1(n13594), .A2(n13913), .ZN(n10673) );
  NAND2_X1 U13268 ( .A1(n10674), .A2(n10673), .ZN(n10903) );
  AOI22_X1 U13269 ( .A1(n10903), .A2(n14359), .B1(P1_REG3_REG_6__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10676) );
  NAND2_X1 U13270 ( .A1(n14358), .A2(n14631), .ZN(n10675) );
  OAI211_X1 U13271 ( .C1(n14365), .C2(n10907), .A(n10676), .B(n10675), .ZN(
        n10677) );
  AOI21_X1 U13272 ( .B1(n10678), .B2(n14350), .A(n10677), .ZN(n10679) );
  INV_X1 U13273 ( .A(n10679), .ZN(P1_U3239) );
  INV_X1 U13274 ( .A(n10680), .ZN(n10681) );
  AND2_X1 U13275 ( .A1(n10682), .A2(n10681), .ZN(n10683) );
  XNOR2_X1 U13276 ( .A(n11895), .B(n9889), .ZN(n10686) );
  NAND2_X1 U13277 ( .A1(n12937), .A2(n12126), .ZN(n10687) );
  NAND2_X1 U13278 ( .A1(n10686), .A2(n10687), .ZN(n10774) );
  INV_X1 U13279 ( .A(n10686), .ZN(n10689) );
  INV_X1 U13280 ( .A(n10687), .ZN(n10688) );
  NAND2_X1 U13281 ( .A1(n10689), .A2(n10688), .ZN(n10690) );
  AND2_X1 U13282 ( .A1(n10774), .A2(n10690), .ZN(n10691) );
  OAI21_X1 U13283 ( .B1(n10692), .B2(n10691), .A(n10775), .ZN(n10693) );
  NAND2_X1 U13284 ( .A1(n10693), .A2(n12887), .ZN(n10698) );
  AND2_X1 U13285 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n14739) );
  NAND2_X1 U13286 ( .A1(n12936), .A2(n12902), .ZN(n10695) );
  NAND2_X1 U13287 ( .A1(n12938), .A2(n12901), .ZN(n10694) );
  AND2_X1 U13288 ( .A1(n10695), .A2(n10694), .ZN(n10994) );
  NOR2_X1 U13289 ( .A1(n12906), .A2(n10994), .ZN(n10696) );
  AOI211_X1 U13290 ( .C1(n12903), .C2(n10989), .A(n14739), .B(n10696), .ZN(
        n10697) );
  OAI211_X1 U13291 ( .C1(n14909), .C2(n12900), .A(n10698), .B(n10697), .ZN(
        P2_U3193) );
  INV_X1 U13292 ( .A(P3_DATAO_REG_29__SCAN_IN), .ZN(n15390) );
  INV_X1 U13293 ( .A(n12503), .ZN(n10699) );
  NAND2_X1 U13294 ( .A1(n10699), .A2(P3_U3897), .ZN(n10700) );
  OAI21_X1 U13295 ( .B1(P3_U3897), .B2(n15390), .A(n10700), .ZN(P3_U3520) );
  OR2_X1 U13296 ( .A1(n10702), .A2(n11725), .ZN(n10703) );
  NAND2_X1 U13297 ( .A1(n10701), .A2(n10703), .ZN(n15158) );
  INV_X1 U13298 ( .A(n15158), .ZN(n10716) );
  INV_X1 U13299 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n10713) );
  AND2_X1 U13300 ( .A1(n10704), .A2(n15122), .ZN(n10710) );
  NAND2_X1 U13301 ( .A1(n10706), .A2(n10705), .ZN(n10707) );
  NAND2_X1 U13302 ( .A1(n10707), .A2(n11725), .ZN(n10709) );
  OAI22_X1 U13303 ( .A1(n10948), .A2(n15117), .B1(n10742), .B2(n15119), .ZN(
        n10708) );
  AOI21_X1 U13304 ( .B1(n10710), .B2(n10709), .A(n10708), .ZN(n10712) );
  NAND2_X1 U13305 ( .A1(n15158), .A2(n11379), .ZN(n10711) );
  AND2_X1 U13306 ( .A1(n10712), .A2(n10711), .ZN(n15160) );
  MUX2_X1 U13307 ( .A(n10713), .B(n15160), .S(n15131), .Z(n10715) );
  AOI22_X1 U13308 ( .A1(n12640), .A2(n15156), .B1(n15591), .B2(n10747), .ZN(
        n10714) );
  OAI211_X1 U13309 ( .C1(n10716), .C2(n12576), .A(n10715), .B(n10714), .ZN(
        P3_U3227) );
  AOI211_X1 U13310 ( .C1(n14905), .C2(n10719), .A(n10718), .B(n10717), .ZN(
        n10722) );
  AOI22_X1 U13311 ( .A1(n13304), .A2(n11890), .B1(n14932), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n10720) );
  OAI21_X1 U13312 ( .B1(n10722), .B2(n14932), .A(n10720), .ZN(P2_U3506) );
  AOI22_X1 U13313 ( .A1(n8982), .A2(n11890), .B1(n14922), .B2(
        P2_REG0_REG_7__SCAN_IN), .ZN(n10721) );
  OAI21_X1 U13314 ( .B1(n10722), .B2(n14922), .A(n10721), .ZN(P2_U3451) );
  INV_X1 U13315 ( .A(n12975), .ZN(n14832) );
  OAI222_X1 U13316 ( .A1(n13357), .A2(n15387), .B1(n13359), .B2(n10723), .C1(
        n14832), .C2(P2_U3088), .ZN(P2_U3309) );
  OAI222_X1 U13317 ( .A1(n14039), .A2(n10725), .B1(n10724), .B2(n10723), .C1(
        n14524), .C2(P1_U3086), .ZN(P1_U3337) );
  NAND2_X1 U13318 ( .A1(n10732), .A2(n10726), .ZN(n10728) );
  NAND2_X1 U13319 ( .A1(n10728), .A2(n10727), .ZN(n12969) );
  XNOR2_X1 U13320 ( .A(n12969), .B(n12959), .ZN(n10729) );
  NAND2_X1 U13321 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n10729), .ZN(n12971) );
  OAI211_X1 U13322 ( .C1(n10729), .C2(P2_REG2_REG_15__SCAN_IN), .A(n14811), 
        .B(n12971), .ZN(n10738) );
  INV_X1 U13323 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n10730) );
  NAND2_X1 U13324 ( .A1(P2_U3088), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n12904)
         );
  OAI21_X1 U13325 ( .B1(n14817), .B2(n10730), .A(n12904), .ZN(n10736) );
  AOI21_X1 U13326 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n10732), .A(n10731), 
        .ZN(n12960) );
  XNOR2_X1 U13327 ( .A(n12959), .B(n12960), .ZN(n10734) );
  INV_X1 U13328 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n10733) );
  NOR2_X1 U13329 ( .A1(n10733), .A2(n10734), .ZN(n12961) );
  AOI211_X1 U13330 ( .C1(n10734), .C2(n10733), .A(n12961), .B(n14819), .ZN(
        n10735) );
  AOI211_X1 U13331 ( .C1(n14809), .C2(n12970), .A(n10736), .B(n10735), .ZN(
        n10737) );
  NAND2_X1 U13332 ( .A1(n10738), .A2(n10737), .ZN(P2_U3229) );
  XNOR2_X1 U13333 ( .A(n15156), .B(n12273), .ZN(n11140) );
  XNOR2_X1 U13334 ( .A(n10785), .B(n11140), .ZN(n10746) );
  INV_X1 U13335 ( .A(n10741), .ZN(n10743) );
  NAND2_X1 U13336 ( .A1(n10743), .A2(n10742), .ZN(n10744) );
  AOI211_X1 U13337 ( .C1(n10746), .C2(n10745), .A(n12382), .B(n6793), .ZN(
        n10751) );
  AOI22_X1 U13338 ( .A1(n12405), .A2(n12291), .B1(n10747), .B2(n12376), .ZN(
        n10749) );
  AOI22_X1 U13339 ( .A1(n12380), .A2(n15156), .B1(P3_REG3_REG_6__SCAN_IN), 
        .B2(P3_U3151), .ZN(n10748) );
  OAI211_X1 U13340 ( .C1(n10948), .C2(n12278), .A(n10749), .B(n10748), .ZN(
        n10750) );
  OR2_X1 U13341 ( .A1(n10751), .A2(n10750), .ZN(P3_U3179) );
  INV_X1 U13342 ( .A(n14558), .ZN(n14642) );
  AOI21_X2 U13343 ( .B1(n10754), .B2(n10753), .A(n10752), .ZN(n10761) );
  NAND2_X1 U13344 ( .A1(n14558), .A2(n13475), .ZN(n10756) );
  NAND2_X1 U13345 ( .A1(n13594), .A2(n13445), .ZN(n10755) );
  NAND2_X1 U13346 ( .A1(n10756), .A2(n10755), .ZN(n10757) );
  XNOR2_X1 U13347 ( .A(n10757), .B(n11318), .ZN(n11004) );
  NAND2_X1 U13348 ( .A1(n14558), .A2(n13445), .ZN(n10759) );
  NAND2_X1 U13349 ( .A1(n13478), .A2(n13594), .ZN(n10758) );
  NAND2_X1 U13350 ( .A1(n10759), .A2(n10758), .ZN(n11005) );
  XNOR2_X1 U13351 ( .A(n11004), .B(n11005), .ZN(n10760) );
  OAI211_X1 U13352 ( .C1(n10761), .C2(n10760), .A(n11008), .B(n14350), .ZN(
        n10768) );
  OR2_X1 U13353 ( .A1(n14536), .A2(n14539), .ZN(n10763) );
  NAND2_X1 U13354 ( .A1(n13595), .A2(n13854), .ZN(n10762) );
  NAND2_X1 U13355 ( .A1(n10763), .A2(n10762), .ZN(n14552) );
  INV_X1 U13356 ( .A(n14552), .ZN(n10765) );
  OAI22_X1 U13357 ( .A1(n10765), .A2(n13546), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10764), .ZN(n10766) );
  AOI21_X1 U13358 ( .B1(n14556), .B2(n13573), .A(n10766), .ZN(n10767) );
  OAI211_X1 U13359 ( .C1(n14642), .C2(n13576), .A(n10768), .B(n10767), .ZN(
        P1_U3213) );
  XNOR2_X1 U13360 ( .A(n11905), .B(n9889), .ZN(n10769) );
  NAND2_X1 U13361 ( .A1(n12936), .A2(n12126), .ZN(n10770) );
  NAND2_X1 U13362 ( .A1(n10769), .A2(n10770), .ZN(n10852) );
  INV_X1 U13363 ( .A(n10769), .ZN(n10772) );
  INV_X1 U13364 ( .A(n10770), .ZN(n10771) );
  NAND2_X1 U13365 ( .A1(n10772), .A2(n10771), .ZN(n10773) );
  AND2_X1 U13366 ( .A1(n10852), .A2(n10773), .ZN(n10777) );
  NAND2_X1 U13367 ( .A1(n10776), .A2(n10777), .ZN(n10853) );
  OAI21_X1 U13368 ( .B1(n10777), .B2(n10776), .A(n10853), .ZN(n10778) );
  NAND2_X1 U13369 ( .A1(n10778), .A2(n12887), .ZN(n10781) );
  AOI22_X1 U13370 ( .A1(n12935), .A2(n12902), .B1(n12901), .B2(n12937), .ZN(
        n10843) );
  NAND2_X1 U13371 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n14759) );
  OAI21_X1 U13372 ( .B1(n10843), .B2(n12906), .A(n14759), .ZN(n10779) );
  AOI21_X1 U13373 ( .B1(n10846), .B2(n12903), .A(n10779), .ZN(n10780) );
  OAI211_X1 U13374 ( .C1(n10939), .C2(n12900), .A(n10781), .B(n10780), .ZN(
        P2_U3203) );
  OAI222_X1 U13375 ( .A1(n13357), .A2(n10782), .B1(P2_U3088), .B2(n12066), 
        .C1(n13359), .C2(n11826), .ZN(P2_U3307) );
  NAND3_X1 U13376 ( .A1(n10701), .A2(n11589), .A3(n11142), .ZN(n10783) );
  NAND2_X1 U13377 ( .A1(n10943), .A2(n10783), .ZN(n15164) );
  INV_X1 U13378 ( .A(n15164), .ZN(n10794) );
  XNOR2_X1 U13379 ( .A(n10784), .B(n11142), .ZN(n10789) );
  NAND2_X1 U13380 ( .A1(n15164), .A2(n11379), .ZN(n10788) );
  OAI22_X1 U13381 ( .A1(n11146), .A2(n15117), .B1(n10785), .B2(n15119), .ZN(
        n10786) );
  INV_X1 U13382 ( .A(n10786), .ZN(n10787) );
  OAI211_X1 U13383 ( .C1(n14264), .C2(n10789), .A(n10788), .B(n10787), .ZN(
        n15162) );
  MUX2_X1 U13384 ( .A(P3_REG2_REG_7__SCAN_IN), .B(n15162), .S(n15131), .Z(
        n10790) );
  INV_X1 U13385 ( .A(n10790), .ZN(n10793) );
  NOR2_X1 U13386 ( .A1(n10791), .A2(n15146), .ZN(n15163) );
  AOI22_X1 U13387 ( .A1(n14276), .A2(n15163), .B1(n15591), .B2(n12185), .ZN(
        n10792) );
  OAI211_X1 U13388 ( .C1(n10794), .C2(n12576), .A(n10793), .B(n10792), .ZN(
        P3_U3226) );
  INV_X1 U13389 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n10826) );
  INV_X1 U13390 ( .A(n10795), .ZN(n10814) );
  NOR2_X1 U13391 ( .A1(n10798), .A2(n10800), .ZN(n10799) );
  AOI22_X1 U13392 ( .A1(n14982), .A2(P3_REG2_REG_6__SCAN_IN), .B1(n10713), 
        .B2(n10812), .ZN(n14975) );
  NOR2_X1 U13393 ( .A1(n14993), .A2(n10801), .ZN(n10802) );
  INV_X1 U13394 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n15000) );
  INV_X1 U13395 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n10803) );
  AOI22_X1 U13396 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n15015), .B1(n10808), 
        .B2(n10803), .ZN(n15010) );
  AOI21_X1 U13397 ( .B1(n10826), .B2(n10804), .A(n12413), .ZN(n10839) );
  INV_X1 U13398 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n15199) );
  INV_X1 U13399 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15191) );
  INV_X1 U13400 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15193) );
  AOI22_X1 U13401 ( .A1(n14982), .A2(P3_REG1_REG_6__SCAN_IN), .B1(n15193), 
        .B2(n10812), .ZN(n14973) );
  INV_X1 U13402 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15195) );
  INV_X1 U13403 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15197) );
  AOI22_X1 U13404 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n15015), .B1(n10808), 
        .B2(n15197), .ZN(n15007) );
  XNOR2_X1 U13405 ( .A(n12459), .B(n12460), .ZN(n10809) );
  AOI21_X1 U13406 ( .B1(n15199), .B2(n10809), .A(n12461), .ZN(n10810) );
  NOR2_X1 U13407 ( .A1(n10810), .A2(n15095), .ZN(n10837) );
  MUX2_X1 U13408 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n12452), .Z(n10822) );
  XNOR2_X1 U13409 ( .A(n10822), .B(n15015), .ZN(n15013) );
  MUX2_X1 U13410 ( .A(n15000), .B(n15195), .S(n12452), .Z(n10811) );
  NAND2_X1 U13411 ( .A1(n10811), .A2(n14993), .ZN(n10821) );
  XOR2_X1 U13412 ( .A(n14993), .B(n10811), .Z(n14992) );
  MUX2_X1 U13413 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n12452), .Z(n10813) );
  OR2_X1 U13414 ( .A1(n10813), .A2(n10812), .ZN(n10820) );
  XNOR2_X1 U13415 ( .A(n10813), .B(n14982), .ZN(n14979) );
  MUX2_X1 U13416 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n12452), .Z(n10819) );
  INV_X1 U13417 ( .A(n14962), .ZN(n10818) );
  XNOR2_X1 U13418 ( .A(n10819), .B(n14962), .ZN(n14960) );
  OAI22_X1 U13419 ( .A1(n10817), .A2(n10816), .B1(n10815), .B2(n10814), .ZN(
        n14961) );
  NAND2_X1 U13420 ( .A1(n14960), .A2(n14961), .ZN(n14959) );
  OAI21_X1 U13421 ( .B1(n10819), .B2(n10818), .A(n14959), .ZN(n14980) );
  NAND2_X1 U13422 ( .A1(n14979), .A2(n14980), .ZN(n14978) );
  NAND2_X1 U13423 ( .A1(n10820), .A2(n14978), .ZN(n14991) );
  NAND2_X1 U13424 ( .A1(n14992), .A2(n14991), .ZN(n14990) );
  INV_X1 U13425 ( .A(n10822), .ZN(n10823) );
  NAND2_X1 U13426 ( .A1(n10823), .A2(n15015), .ZN(n10824) );
  NAND2_X1 U13427 ( .A1(n10825), .A2(n10824), .ZN(n12431) );
  MUX2_X1 U13428 ( .A(n10826), .B(n15199), .S(n12452), .Z(n10827) );
  AND2_X1 U13429 ( .A1(n10827), .A2(n12460), .ZN(n12430) );
  INV_X1 U13430 ( .A(n12430), .ZN(n10830) );
  INV_X1 U13431 ( .A(n10827), .ZN(n10829) );
  INV_X1 U13432 ( .A(n12460), .ZN(n10828) );
  NAND2_X1 U13433 ( .A1(n10829), .A2(n10828), .ZN(n12432) );
  NAND2_X1 U13434 ( .A1(n10830), .A2(n12432), .ZN(n10831) );
  XNOR2_X1 U13435 ( .A(n12431), .B(n10831), .ZN(n10835) );
  NAND2_X1 U13436 ( .A1(n15016), .A2(n12460), .ZN(n10834) );
  NOR2_X1 U13437 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11152), .ZN(n10832) );
  AOI21_X1 U13438 ( .B1(n15025), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n10832), .ZN(
        n10833) );
  OAI211_X1 U13439 ( .C1(n10835), .C2(n15082), .A(n10834), .B(n10833), .ZN(
        n10836) );
  NOR2_X1 U13440 ( .A1(n10837), .A2(n10836), .ZN(n10838) );
  OAI21_X1 U13441 ( .B1(n10839), .B2(n15110), .A(n10838), .ZN(P3_U3191) );
  XOR2_X1 U13442 ( .A(n12080), .B(n10840), .Z(n10936) );
  INV_X1 U13443 ( .A(n10936), .ZN(n10851) );
  INV_X1 U13444 ( .A(n12080), .ZN(n10842) );
  OAI211_X1 U13445 ( .C1(n6798), .C2(n10842), .A(n14304), .B(n10841), .ZN(
        n10844) );
  NAND2_X1 U13446 ( .A1(n10844), .A2(n10843), .ZN(n10934) );
  INV_X1 U13447 ( .A(n10845), .ZN(n10987) );
  AOI211_X1 U13448 ( .C1(n11905), .C2(n10987), .A(n13049), .B(n10968), .ZN(
        n10935) );
  NAND2_X1 U13449 ( .A1(n10935), .A2(n14315), .ZN(n10848) );
  AOI22_X1 U13450 ( .A1(n13216), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n10846), 
        .B2(n14841), .ZN(n10847) );
  OAI211_X1 U13451 ( .C1(n10939), .C2(n14835), .A(n10848), .B(n10847), .ZN(
        n10849) );
  AOI21_X1 U13452 ( .B1(n10934), .B2(n14837), .A(n10849), .ZN(n10850) );
  OAI21_X1 U13453 ( .B1(n10851), .B2(n13182), .A(n10850), .ZN(P2_U3256) );
  NAND2_X1 U13454 ( .A1(n10853), .A2(n10852), .ZN(n11043) );
  XNOR2_X1 U13455 ( .A(n11910), .B(n12154), .ZN(n11040) );
  NOR2_X1 U13456 ( .A1(n11909), .A2(n14313), .ZN(n11039) );
  XNOR2_X1 U13457 ( .A(n11040), .B(n11039), .ZN(n11042) );
  XNOR2_X1 U13458 ( .A(n11043), .B(n11042), .ZN(n10861) );
  INV_X1 U13459 ( .A(n10969), .ZN(n10858) );
  NAND2_X1 U13460 ( .A1(n12934), .A2(n12902), .ZN(n10855) );
  NAND2_X1 U13461 ( .A1(n12936), .A2(n12901), .ZN(n10854) );
  NAND2_X1 U13462 ( .A1(n10855), .A2(n10854), .ZN(n10964) );
  AOI21_X1 U13463 ( .B1(n12897), .B2(n10964), .A(n10856), .ZN(n10857) );
  OAI21_X1 U13464 ( .B1(n12894), .B2(n10858), .A(n10857), .ZN(n10859) );
  AOI21_X1 U13465 ( .B1(n11910), .B2(n12913), .A(n10859), .ZN(n10860) );
  OAI21_X1 U13466 ( .B1(n10861), .B2(n12908), .A(n10860), .ZN(P2_U3189) );
  NAND2_X1 U13467 ( .A1(n10863), .A2(n10862), .ZN(n10865) );
  NOR2_X1 U13468 ( .A1(n13597), .A2(n14612), .ZN(n10866) );
  XNOR2_X1 U13469 ( .A(n10897), .B(n10893), .ZN(n10870) );
  AOI21_X1 U13470 ( .B1(n10870), .B2(n14554), .A(n10869), .ZN(n14626) );
  INV_X1 U13471 ( .A(n10871), .ZN(n10872) );
  NAND3_X1 U13472 ( .A1(n10876), .A2(n10875), .A3(n10874), .ZN(n11808) );
  NAND2_X1 U13473 ( .A1(n11086), .A2(n14612), .ZN(n11085) );
  INV_X1 U13474 ( .A(n11066), .ZN(n10877) );
  OAI211_X1 U13475 ( .C1(n10898), .C2(n10877), .A(n10906), .B(n14561), .ZN(
        n14623) );
  INV_X1 U13476 ( .A(n14623), .ZN(n10884) );
  INV_X2 U13477 ( .A(n13902), .ZN(n14570) );
  NOR2_X2 U13478 ( .A1(n14570), .A2(n10878), .ZN(n14567) );
  NAND2_X1 U13479 ( .A1(n10012), .A2(n10879), .ZN(n10880) );
  NOR2_X2 U13480 ( .A1(n14570), .A2(n10880), .ZN(n14557) );
  AOI22_X1 U13481 ( .A1(n14570), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n10881), 
        .B2(n14569), .ZN(n10882) );
  OAI21_X1 U13482 ( .B1(n14573), .B2(n10898), .A(n10882), .ZN(n10883) );
  AOI21_X1 U13483 ( .B1(n10884), .B2(n14567), .A(n10883), .ZN(n10892) );
  INV_X1 U13484 ( .A(n11090), .ZN(n11081) );
  NAND2_X1 U13485 ( .A1(n11082), .A2(n11081), .ZN(n11084) );
  INV_X1 U13486 ( .A(n13597), .ZN(n10887) );
  NAND2_X1 U13487 ( .A1(n10887), .A2(n14612), .ZN(n10888) );
  XNOR2_X1 U13488 ( .A(n10894), .B(n10893), .ZN(n14628) );
  NOR2_X1 U13489 ( .A1(n14570), .A2(n10890), .ZN(n14577) );
  AOI21_X1 U13490 ( .B1(n14639), .B2(n13902), .A(n14577), .ZN(n13785) );
  NAND2_X1 U13491 ( .A1(n14628), .A2(n6805), .ZN(n10891) );
  OAI211_X1 U13492 ( .C1(n14626), .C2(n13930), .A(n10892), .B(n10891), .ZN(
        P1_U3288) );
  INV_X1 U13493 ( .A(n13596), .ZN(n10900) );
  NAND2_X1 U13494 ( .A1(n10900), .A2(n10898), .ZN(n10895) );
  NAND2_X1 U13495 ( .A1(n10896), .A2(n10895), .ZN(n11116) );
  XOR2_X1 U13496 ( .A(n11128), .B(n11116), .Z(n14635) );
  XNOR2_X1 U13497 ( .A(n11129), .B(n11128), .ZN(n10904) );
  AOI21_X1 U13498 ( .B1(n10904), .B2(n14554), .A(n10903), .ZN(n14634) );
  MUX2_X1 U13499 ( .A(n10905), .B(n14634), .S(n13902), .Z(n10910) );
  AOI211_X1 U13500 ( .C1(n14631), .C2(n10906), .A(n13903), .B(n14563), .ZN(
        n14630) );
  OAI22_X1 U13501 ( .A1(n14573), .A2(n11127), .B1(n10907), .B2(n13857), .ZN(
        n10908) );
  AOI21_X1 U13502 ( .B1(n14630), .B2(n14567), .A(n10908), .ZN(n10909) );
  OAI211_X1 U13503 ( .C1(n13785), .C2(n14635), .A(n10910), .B(n10909), .ZN(
        P1_U3287) );
  AOI21_X1 U13504 ( .B1(n14567), .B2(n10012), .A(n14557), .ZN(n10919) );
  OAI22_X1 U13505 ( .A1(n14570), .A2(n10912), .B1(n10911), .B2(n13857), .ZN(
        n10913) );
  AOI21_X1 U13506 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n13930), .A(n10913), .ZN(
        n10917) );
  NAND2_X1 U13507 ( .A1(n13902), .A2(n10914), .ZN(n13896) );
  NOR2_X1 U13508 ( .A1(n14570), .A2(n14666), .ZN(n13863) );
  OAI21_X1 U13509 ( .B1(n14175), .B2(n13863), .A(n10915), .ZN(n10916) );
  OAI211_X1 U13510 ( .C1(n10919), .C2(n10918), .A(n10917), .B(n10916), .ZN(
        P1_U3293) );
  INV_X1 U13511 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10921) );
  INV_X1 U13512 ( .A(n10920), .ZN(n10922) );
  OAI222_X1 U13513 ( .A1(n13357), .A2(n10921), .B1(n13359), .B2(n10922), .C1(
        n12983), .C2(P2_U3088), .ZN(P2_U3308) );
  OAI222_X1 U13514 ( .A1(n14039), .A2(n10923), .B1(n10724), .B2(n10922), .C1(
        P1_U3086), .C2(n13685), .ZN(P1_U3336) );
  XNOR2_X1 U13515 ( .A(n10924), .B(n11728), .ZN(n15171) );
  INV_X1 U13516 ( .A(n11379), .ZN(n15125) );
  AOI22_X1 U13517 ( .A1(n12402), .A2(n12374), .B1(n12375), .B2(n12400), .ZN(
        n10929) );
  AND2_X1 U13518 ( .A1(n10947), .A2(n10925), .ZN(n10927) );
  OAI211_X1 U13519 ( .C1(n10927), .C2(n11728), .A(n10926), .B(n15122), .ZN(
        n10928) );
  OAI211_X1 U13520 ( .C1(n15171), .C2(n15125), .A(n10929), .B(n10928), .ZN(
        n15172) );
  NAND2_X1 U13521 ( .A1(n15172), .A2(n12657), .ZN(n10933) );
  NOR2_X1 U13522 ( .A1(n11153), .A2(n15146), .ZN(n15173) );
  INV_X1 U13523 ( .A(n11155), .ZN(n10930) );
  OAI22_X1 U13524 ( .A1(n12657), .A2(n10826), .B1(n10930), .B2(n14270), .ZN(
        n10931) );
  AOI21_X1 U13525 ( .B1(n14276), .B2(n15173), .A(n10931), .ZN(n10932) );
  OAI211_X1 U13526 ( .C1(n15171), .C2(n12576), .A(n10933), .B(n10932), .ZN(
        P3_U3224) );
  AOI211_X1 U13527 ( .C1(n10936), .C2(n14905), .A(n10935), .B(n10934), .ZN(
        n10942) );
  AOI22_X1 U13528 ( .A1(n11905), .A2(n13304), .B1(n14932), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n10937) );
  OAI21_X1 U13529 ( .B1(n10942), .B2(n14932), .A(n10937), .ZN(P2_U3508) );
  INV_X1 U13530 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10938) );
  OAI22_X1 U13531 ( .A1(n10939), .A2(n13329), .B1(n14924), .B2(n10938), .ZN(
        n10940) );
  INV_X1 U13532 ( .A(n10940), .ZN(n10941) );
  OAI21_X1 U13533 ( .B1(n10942), .B2(n14922), .A(n10941), .ZN(P2_U3457) );
  NAND2_X1 U13534 ( .A1(n10943), .A2(n11594), .ZN(n10944) );
  XNOR2_X1 U13535 ( .A(n10944), .B(n11720), .ZN(n15169) );
  INV_X1 U13536 ( .A(n15169), .ZN(n10955) );
  NAND2_X1 U13537 ( .A1(n15169), .A2(n11379), .ZN(n10952) );
  NAND2_X1 U13538 ( .A1(n10945), .A2(n11720), .ZN(n10946) );
  NAND2_X1 U13539 ( .A1(n10947), .A2(n10946), .ZN(n10950) );
  OAI22_X1 U13540 ( .A1(n11336), .A2(n15117), .B1(n10948), .B2(n15119), .ZN(
        n10949) );
  AOI21_X1 U13541 ( .B1(n10950), .B2(n15122), .A(n10949), .ZN(n10951) );
  AND2_X1 U13542 ( .A1(n10952), .A2(n10951), .ZN(n15166) );
  MUX2_X1 U13543 ( .A(n10803), .B(n15166), .S(n15131), .Z(n10954) );
  NOR2_X1 U13544 ( .A1(n12287), .A2(n15146), .ZN(n15168) );
  AOI22_X1 U13545 ( .A1(n14276), .A2(n15168), .B1(n15591), .B2(n12290), .ZN(
        n10953) );
  OAI211_X1 U13546 ( .C1(n10955), .C2(n12576), .A(n10954), .B(n10953), .ZN(
        P3_U3225) );
  INV_X1 U13547 ( .A(n10956), .ZN(n10958) );
  OAI222_X1 U13548 ( .A1(P3_U3151), .A2(n10959), .B1(n12785), .B2(n10958), 
        .C1(n10957), .C2(n12787), .ZN(P3_U3271) );
  NAND2_X1 U13549 ( .A1(n11902), .A2(n10960), .ZN(n12081) );
  INV_X1 U13550 ( .A(n12081), .ZN(n10961) );
  XNOR2_X1 U13551 ( .A(n10962), .B(n10961), .ZN(n14919) );
  INV_X1 U13552 ( .A(n9870), .ZN(n11160) );
  NAND2_X1 U13553 ( .A1(n14919), .A2(n11160), .ZN(n10967) );
  XNOR2_X1 U13554 ( .A(n10963), .B(n12081), .ZN(n10965) );
  AOI21_X1 U13555 ( .B1(n10965), .B2(n14304), .A(n10964), .ZN(n10966) );
  AND2_X1 U13556 ( .A1(n10967), .A2(n10966), .ZN(n14921) );
  INV_X2 U13557 ( .A(n14837), .ZN(n13216) );
  OAI211_X1 U13558 ( .C1(n10968), .C2(n14916), .A(n14313), .B(n11108), .ZN(
        n14914) );
  AOI22_X1 U13559 ( .A1(n13216), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n10969), 
        .B2(n14841), .ZN(n10971) );
  NAND2_X1 U13560 ( .A1(n11910), .A2(n14307), .ZN(n10970) );
  OAI211_X1 U13561 ( .C1(n14914), .C2(n13213), .A(n10971), .B(n10970), .ZN(
        n10972) );
  AOI21_X1 U13562 ( .B1(n14919), .B2(n14845), .A(n10972), .ZN(n10973) );
  OAI21_X1 U13563 ( .B1(n14921), .B2(n13216), .A(n10973), .ZN(P2_U3255) );
  OAI222_X1 U13564 ( .A1(P1_U3086), .A2(n7399), .B1(n10724), .B2(n10999), .C1(
        n10974), .C2(n14039), .ZN(P1_U3334) );
  NAND2_X1 U13565 ( .A1(n14567), .A2(n10975), .ZN(n10979) );
  NAND2_X1 U13566 ( .A1(n14557), .A2(n10976), .ZN(n10978) );
  AOI22_X1 U13567 ( .A1(n14570), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n14569), .ZN(n10977) );
  NAND3_X1 U13568 ( .A1(n10979), .A2(n10978), .A3(n10977), .ZN(n10980) );
  AOI21_X1 U13569 ( .B1(n14577), .B2(n10981), .A(n10980), .ZN(n10982) );
  OAI21_X1 U13570 ( .B1(n10983), .B2(n13930), .A(n10982), .ZN(P1_U3292) );
  NAND2_X1 U13571 ( .A1(n10984), .A2(n12078), .ZN(n10985) );
  NAND2_X1 U13572 ( .A1(n10986), .A2(n10985), .ZN(n10995) );
  INV_X1 U13573 ( .A(n10995), .ZN(n14912) );
  OAI211_X1 U13574 ( .C1(n14909), .C2(n10988), .A(n10987), .B(n14313), .ZN(
        n14908) );
  AOI22_X1 U13575 ( .A1(n11895), .A2(n14307), .B1(n14841), .B2(n10989), .ZN(
        n10990) );
  OAI21_X1 U13576 ( .B1(n14908), .B2(n13213), .A(n10990), .ZN(n10997) );
  XNOR2_X1 U13577 ( .A(n10991), .B(n7510), .ZN(n10992) );
  NAND2_X1 U13578 ( .A1(n10992), .A2(n14304), .ZN(n10993) );
  OAI211_X1 U13579 ( .C1(n10995), .C2(n9870), .A(n10994), .B(n10993), .ZN(
        n14910) );
  MUX2_X1 U13580 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n14910), .S(n14837), .Z(
        n10996) );
  AOI211_X1 U13581 ( .C1(n14912), .C2(n14845), .A(n10997), .B(n10996), .ZN(
        n10998) );
  INV_X1 U13582 ( .A(n10998), .ZN(P2_U3257) );
  OAI222_X1 U13583 ( .A1(n13357), .A2(n11000), .B1(P2_U3088), .B2(n8343), .C1(
        n13359), .C2(n10999), .ZN(P2_U3306) );
  NAND2_X1 U13584 ( .A1(n11198), .A2(n13475), .ZN(n11002) );
  OR2_X1 U13585 ( .A1(n14536), .A2(n13407), .ZN(n11001) );
  NAND2_X1 U13586 ( .A1(n11002), .A2(n11001), .ZN(n11003) );
  XNOR2_X1 U13587 ( .A(n11003), .B(n11318), .ZN(n11052) );
  AOI22_X1 U13588 ( .A1(n11198), .A2(n13445), .B1(n13593), .B2(n13478), .ZN(
        n11051) );
  XNOR2_X1 U13589 ( .A(n11052), .B(n11051), .ZN(n11011) );
  INV_X1 U13590 ( .A(n11004), .ZN(n11006) );
  NAND2_X1 U13591 ( .A1(n11006), .A2(n11005), .ZN(n11007) );
  INV_X1 U13592 ( .A(n11011), .ZN(n11009) );
  INV_X1 U13593 ( .A(n11220), .ZN(n11053) );
  AOI21_X1 U13594 ( .B1(n11011), .B2(n11010), .A(n11053), .ZN(n11019) );
  INV_X1 U13595 ( .A(n11198), .ZN(n11123) );
  NOR2_X1 U13596 ( .A1(n11123), .A2(n14665), .ZN(n14649) );
  INV_X1 U13597 ( .A(n11124), .ZN(n11015) );
  OR2_X1 U13598 ( .A1(n11207), .A2(n14539), .ZN(n11013) );
  NAND2_X1 U13599 ( .A1(n13594), .A2(n13854), .ZN(n11012) );
  NAND2_X1 U13600 ( .A1(n11013), .A2(n11012), .ZN(n11131) );
  AOI22_X1 U13601 ( .A1(n11131), .A2(n14359), .B1(P1_REG3_REG_8__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11014) );
  OAI21_X1 U13602 ( .B1(n14365), .B2(n11015), .A(n11014), .ZN(n11016) );
  AOI21_X1 U13603 ( .B1(n11017), .B2(n14649), .A(n11016), .ZN(n11018) );
  OAI21_X1 U13604 ( .B1(n11019), .B2(n13564), .A(n11018), .ZN(P1_U3221) );
  INV_X1 U13605 ( .A(n11020), .ZN(n11023) );
  OAI222_X1 U13606 ( .A1(n12785), .A2(n11023), .B1(P3_U3151), .B2(n11022), 
        .C1(n11021), .C2(n12787), .ZN(P3_U3270) );
  INV_X1 U13607 ( .A(n11024), .ZN(n11026) );
  INV_X1 U13608 ( .A(n11605), .ZN(n11730) );
  OAI21_X1 U13609 ( .B1(n11026), .B2(n11730), .A(n11025), .ZN(n15176) );
  XNOR2_X1 U13610 ( .A(n11027), .B(n11730), .ZN(n11029) );
  OAI22_X1 U13611 ( .A1(n11336), .A2(n15119), .B1(n12249), .B2(n15117), .ZN(
        n11028) );
  AOI21_X1 U13612 ( .B1(n11029), .B2(n15122), .A(n11028), .ZN(n11030) );
  OAI21_X1 U13613 ( .B1(n15176), .B2(n15125), .A(n11030), .ZN(n15177) );
  NAND2_X1 U13614 ( .A1(n15177), .A2(n12657), .ZN(n11034) );
  NOR2_X1 U13615 ( .A1(n11609), .A2(n15146), .ZN(n15178) );
  INV_X1 U13616 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n12429) );
  INV_X1 U13617 ( .A(n12247), .ZN(n11031) );
  OAI22_X1 U13618 ( .A1(n12657), .A2(n12429), .B1(n11031), .B2(n14270), .ZN(
        n11032) );
  AOI21_X1 U13619 ( .B1(n14276), .B2(n15178), .A(n11032), .ZN(n11033) );
  OAI211_X1 U13620 ( .C1(n15176), .C2(n12576), .A(n11034), .B(n11033), .ZN(
        P3_U3223) );
  XNOR2_X1 U13621 ( .A(n11919), .B(n9889), .ZN(n11035) );
  NAND2_X1 U13622 ( .A1(n12934), .A2(n12126), .ZN(n11036) );
  NAND2_X1 U13623 ( .A1(n11035), .A2(n11036), .ZN(n11182) );
  INV_X1 U13624 ( .A(n11035), .ZN(n11038) );
  INV_X1 U13625 ( .A(n11036), .ZN(n11037) );
  NAND2_X1 U13626 ( .A1(n11038), .A2(n11037), .ZN(n11184) );
  NAND2_X1 U13627 ( .A1(n11182), .A2(n11184), .ZN(n11044) );
  NAND2_X1 U13628 ( .A1(n11040), .A2(n11039), .ZN(n11041) );
  OAI21_X1 U13629 ( .B1(n11043), .B2(n11042), .A(n11041), .ZN(n11183) );
  XOR2_X1 U13630 ( .A(n11044), .B(n11183), .Z(n11050) );
  INV_X1 U13631 ( .A(n11109), .ZN(n11047) );
  NAND2_X1 U13632 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n14773)
         );
  NAND2_X1 U13633 ( .A1(n12933), .A2(n12902), .ZN(n11045) );
  OAI21_X1 U13634 ( .B1(n11909), .B2(n12889), .A(n11045), .ZN(n11104) );
  NAND2_X1 U13635 ( .A1(n11104), .A2(n12897), .ZN(n11046) );
  OAI211_X1 U13636 ( .C1(n12894), .C2(n11047), .A(n14773), .B(n11046), .ZN(
        n11048) );
  AOI21_X1 U13637 ( .B1(n11919), .B2(n12913), .A(n11048), .ZN(n11049) );
  OAI21_X1 U13638 ( .B1(n11050), .B2(n12908), .A(n11049), .ZN(P2_U3208) );
  AND2_X1 U13639 ( .A1(n11052), .A2(n11051), .ZN(n11217) );
  NOR2_X1 U13640 ( .A1(n11053), .A2(n11217), .ZN(n11058) );
  OAI22_X1 U13641 ( .A1(n14658), .A2(n6962), .B1(n11207), .B2(n13407), .ZN(
        n11054) );
  XNOR2_X1 U13642 ( .A(n11054), .B(n11318), .ZN(n11221) );
  OR2_X1 U13643 ( .A1(n14658), .A2(n13407), .ZN(n11056) );
  OR2_X1 U13644 ( .A1(n11207), .A2(n13405), .ZN(n11055) );
  AND2_X1 U13645 ( .A1(n11056), .A2(n11055), .ZN(n11218) );
  INV_X1 U13646 ( .A(n11218), .ZN(n11222) );
  XNOR2_X1 U13647 ( .A(n11221), .B(n11222), .ZN(n11057) );
  XNOR2_X1 U13648 ( .A(n11058), .B(n11057), .ZN(n11064) );
  INV_X1 U13649 ( .A(n14540), .ZN(n11061) );
  AOI22_X1 U13650 ( .A1(n13568), .A2(n13593), .B1(P1_REG3_REG_9__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11060) );
  INV_X1 U13651 ( .A(n13571), .ZN(n11239) );
  NAND2_X1 U13652 ( .A1(n11239), .A2(n13591), .ZN(n11059) );
  OAI211_X1 U13653 ( .C1(n14365), .C2(n11061), .A(n11060), .B(n11059), .ZN(
        n11062) );
  AOI21_X1 U13654 ( .B1(n14358), .B2(n14541), .A(n11062), .ZN(n11063) );
  OAI21_X1 U13655 ( .B1(n11064), .B2(n13564), .A(n11063), .ZN(P1_U3231) );
  XOR2_X1 U13656 ( .A(n11074), .B(n11065), .Z(n14621) );
  AOI21_X1 U13657 ( .B1(n11085), .B2(n11072), .A(n13903), .ZN(n11067) );
  NAND2_X1 U13658 ( .A1(n11067), .A2(n11066), .ZN(n14616) );
  INV_X1 U13659 ( .A(n11068), .ZN(n11069) );
  OAI22_X1 U13660 ( .A1(n13902), .A2(n11070), .B1(n11069), .B2(n13857), .ZN(
        n11071) );
  AOI21_X1 U13661 ( .B1(n14557), .B2(n11072), .A(n11071), .ZN(n11073) );
  OAI21_X1 U13662 ( .B1(n13927), .B2(n14616), .A(n11073), .ZN(n11079) );
  INV_X1 U13663 ( .A(n11074), .ZN(n11075) );
  XNOR2_X1 U13664 ( .A(n6803), .B(n11075), .ZN(n11076) );
  NAND2_X1 U13665 ( .A1(n11076), .A2(n14554), .ZN(n14619) );
  INV_X1 U13666 ( .A(n11077), .ZN(n14618) );
  AOI21_X1 U13667 ( .B1(n14619), .B2(n14618), .A(n14570), .ZN(n11078) );
  AOI211_X1 U13668 ( .C1(n14621), .C2(n14175), .A(n11079), .B(n11078), .ZN(
        n11080) );
  INV_X1 U13669 ( .A(n11080), .ZN(P1_U3289) );
  OR2_X1 U13670 ( .A1(n11082), .A2(n11081), .ZN(n11083) );
  NAND2_X1 U13671 ( .A1(n11084), .A2(n11083), .ZN(n14609) );
  OAI211_X1 U13672 ( .C1(n11086), .C2(n14612), .A(n11085), .B(n14561), .ZN(
        n14610) );
  AOI22_X1 U13673 ( .A1(n14557), .A2(n11088), .B1(n14569), .B2(n11087), .ZN(
        n11089) );
  OAI21_X1 U13674 ( .B1(n13927), .B2(n14610), .A(n11089), .ZN(n11098) );
  NAND2_X1 U13675 ( .A1(n14609), .A2(n14639), .ZN(n11096) );
  XNOR2_X1 U13676 ( .A(n11091), .B(n11090), .ZN(n11094) );
  OAI22_X1 U13677 ( .A1(n10144), .A2(n14537), .B1(n11092), .B2(n14539), .ZN(
        n11093) );
  AOI21_X1 U13678 ( .B1(n11094), .B2(n14554), .A(n11093), .ZN(n11095) );
  NAND2_X1 U13679 ( .A1(n11096), .A2(n11095), .ZN(n14613) );
  MUX2_X1 U13680 ( .A(n14613), .B(P1_REG2_REG_3__SCAN_IN), .S(n13930), .Z(
        n11097) );
  AOI211_X1 U13681 ( .C1(n14577), .C2(n14609), .A(n11098), .B(n11097), .ZN(
        n11099) );
  INV_X1 U13682 ( .A(n11099), .ZN(P1_U3290) );
  XNOR2_X1 U13683 ( .A(n11100), .B(n11102), .ZN(n11276) );
  OAI21_X1 U13684 ( .B1(n11103), .B2(n11102), .A(n11101), .ZN(n11105) );
  AOI21_X1 U13685 ( .B1(n11105), .B2(n14304), .A(n11104), .ZN(n11106) );
  OAI21_X1 U13686 ( .B1(n11276), .B2(n9870), .A(n11106), .ZN(n11277) );
  NAND2_X1 U13687 ( .A1(n11277), .A2(n14837), .ZN(n11114) );
  INV_X1 U13688 ( .A(n11168), .ZN(n11107) );
  AOI211_X1 U13689 ( .C1(n11919), .C2(n11108), .A(n12126), .B(n11107), .ZN(
        n11278) );
  INV_X1 U13690 ( .A(n11919), .ZN(n11111) );
  AOI22_X1 U13691 ( .A1(n13216), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n11109), 
        .B2(n14841), .ZN(n11110) );
  OAI21_X1 U13692 ( .B1(n11111), .B2(n14835), .A(n11110), .ZN(n11112) );
  AOI21_X1 U13693 ( .B1(n11278), .B2(n14315), .A(n11112), .ZN(n11113) );
  OAI211_X1 U13694 ( .C1(n11276), .C2(n11115), .A(n11114), .B(n11113), .ZN(
        P2_U3254) );
  NAND2_X1 U13695 ( .A1(n11116), .A2(n11128), .ZN(n11119) );
  INV_X1 U13696 ( .A(n13595), .ZN(n11117) );
  NAND2_X1 U13697 ( .A1(n11117), .A2(n11127), .ZN(n11118) );
  INV_X1 U13698 ( .A(n14549), .ZN(n11120) );
  OR2_X1 U13699 ( .A1(n13594), .A2(n14558), .ZN(n11121) );
  XNOR2_X1 U13700 ( .A(n11197), .B(n11196), .ZN(n14655) );
  INV_X1 U13701 ( .A(n14543), .ZN(n11122) );
  OAI211_X1 U13702 ( .C1(n11123), .C2(n14560), .A(n11122), .B(n14561), .ZN(
        n14650) );
  AOI22_X1 U13703 ( .A1(n14570), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n11124), 
        .B2(n14569), .ZN(n11126) );
  NAND2_X1 U13704 ( .A1(n14557), .A2(n11198), .ZN(n11125) );
  OAI211_X1 U13705 ( .C1(n14650), .C2(n13927), .A(n11126), .B(n11125), .ZN(
        n11133) );
  INV_X1 U13706 ( .A(n11196), .ZN(n11130) );
  OAI211_X1 U13707 ( .C1(n6799), .C2(n11130), .A(n11206), .B(n14554), .ZN(
        n14653) );
  INV_X1 U13708 ( .A(n11131), .ZN(n14652) );
  AOI21_X1 U13709 ( .B1(n14653), .B2(n14652), .A(n13930), .ZN(n11132) );
  AOI211_X1 U13710 ( .C1(n14175), .C2(n14655), .A(n11133), .B(n11132), .ZN(
        n11134) );
  INV_X1 U13711 ( .A(n11134), .ZN(P1_U3285) );
  INV_X1 U13712 ( .A(n11135), .ZN(n11137) );
  OAI222_X1 U13713 ( .A1(P3_U3151), .A2(n11138), .B1(n12785), .B2(n11137), 
        .C1(n11136), .C2(n12787), .ZN(P3_U3269) );
  XNOR2_X1 U13714 ( .A(n11139), .B(n12273), .ZN(n11337) );
  XNOR2_X1 U13715 ( .A(n11337), .B(n11336), .ZN(n11151) );
  INV_X1 U13716 ( .A(n11140), .ZN(n11141) );
  XNOR2_X1 U13717 ( .A(n11142), .B(n12220), .ZN(n12182) );
  INV_X1 U13718 ( .A(n12182), .ZN(n11143) );
  NAND2_X1 U13719 ( .A1(n11143), .A2(n12403), .ZN(n11144) );
  XNOR2_X1 U13720 ( .A(n11145), .B(n12220), .ZN(n11147) );
  XNOR2_X1 U13721 ( .A(n11146), .B(n11147), .ZN(n12284) );
  NAND2_X1 U13722 ( .A1(n12285), .A2(n12284), .ZN(n12283) );
  NAND2_X1 U13723 ( .A1(n12402), .A2(n11147), .ZN(n11148) );
  NAND2_X1 U13724 ( .A1(n12283), .A2(n11148), .ZN(n11150) );
  INV_X1 U13725 ( .A(n11339), .ZN(n11149) );
  AOI21_X1 U13726 ( .B1(n11151), .B2(n11150), .A(n11149), .ZN(n11158) );
  OAI22_X1 U13727 ( .A1(n12352), .A2(n11153), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11152), .ZN(n11154) );
  AOI21_X1 U13728 ( .B1(n12289), .B2(n12400), .A(n11154), .ZN(n11157) );
  AOI22_X1 U13729 ( .A1(n12402), .A2(n12291), .B1(n11155), .B2(n12376), .ZN(
        n11156) );
  OAI211_X1 U13730 ( .C1(n11158), .C2(n12382), .A(n11157), .B(n11156), .ZN(
        P3_U3171) );
  XNOR2_X1 U13731 ( .A(n11159), .B(n7947), .ZN(n14333) );
  NAND2_X1 U13732 ( .A1(n14333), .A2(n11160), .ZN(n11167) );
  AOI21_X1 U13733 ( .B1(n11161), .B2(n12085), .A(n13171), .ZN(n11165) );
  NAND2_X1 U13734 ( .A1(n12932), .A2(n12902), .ZN(n11163) );
  NAND2_X1 U13735 ( .A1(n12934), .A2(n12901), .ZN(n11162) );
  NAND2_X1 U13736 ( .A1(n11163), .A2(n11162), .ZN(n11190) );
  AOI21_X1 U13737 ( .B1(n11165), .B2(n11164), .A(n11190), .ZN(n11166) );
  AND2_X1 U13738 ( .A1(n11167), .A2(n11166), .ZN(n14335) );
  NAND2_X1 U13739 ( .A1(n14329), .A2(n11168), .ZN(n11169) );
  NAND2_X1 U13740 ( .A1(n11169), .A2(n14313), .ZN(n11170) );
  OR2_X1 U13741 ( .A1(n11252), .A2(n11170), .ZN(n14331) );
  AOI22_X1 U13742 ( .A1(n13216), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n11189), 
        .B2(n14841), .ZN(n11172) );
  NAND2_X1 U13743 ( .A1(n14329), .A2(n14307), .ZN(n11171) );
  OAI211_X1 U13744 ( .C1(n14331), .C2(n13213), .A(n11172), .B(n11171), .ZN(
        n11173) );
  AOI21_X1 U13745 ( .B1(n14333), .B2(n14845), .A(n11173), .ZN(n11174) );
  OAI21_X1 U13746 ( .B1(n14335), .B2(n13216), .A(n11174), .ZN(P2_U3253) );
  INV_X1 U13747 ( .A(n11175), .ZN(n11176) );
  OAI222_X1 U13748 ( .A1(n13357), .A2(n11177), .B1(n13359), .B2(n11176), .C1(
        n12058), .C2(P2_U3088), .ZN(P2_U3305) );
  INV_X1 U13749 ( .A(n11178), .ZN(n11180) );
  OAI222_X1 U13750 ( .A1(n12452), .A2(P3_U3151), .B1(n12785), .B2(n11180), 
        .C1(n11179), .C2(n12787), .ZN(P3_U3268) );
  XNOR2_X1 U13751 ( .A(n14329), .B(n9889), .ZN(n11286) );
  NAND2_X1 U13752 ( .A1(n12933), .A2(n13049), .ZN(n11285) );
  XNOR2_X1 U13753 ( .A(n11286), .B(n11285), .ZN(n11188) );
  INV_X1 U13754 ( .A(n11288), .ZN(n11186) );
  AOI21_X1 U13755 ( .B1(n11188), .B2(n11187), .A(n11186), .ZN(n11195) );
  INV_X1 U13756 ( .A(n11189), .ZN(n11192) );
  NAND2_X1 U13757 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n14789)
         );
  NAND2_X1 U13758 ( .A1(n12897), .A2(n11190), .ZN(n11191) );
  OAI211_X1 U13759 ( .C1(n12894), .C2(n11192), .A(n14789), .B(n11191), .ZN(
        n11193) );
  AOI21_X1 U13760 ( .B1(n14329), .B2(n12913), .A(n11193), .ZN(n11194) );
  OAI21_X1 U13761 ( .B1(n11195), .B2(n12908), .A(n11194), .ZN(P2_U3196) );
  NAND2_X1 U13762 ( .A1(n14658), .A2(n11207), .ZN(n11200) );
  XNOR2_X1 U13763 ( .A(n11258), .B(n7189), .ZN(n14672) );
  NAND2_X1 U13764 ( .A1(n14543), .A2(n14658), .ZN(n14542) );
  OR2_X1 U13765 ( .A1(n14542), .A2(n14357), .ZN(n11267) );
  INV_X1 U13766 ( .A(n11267), .ZN(n11268) );
  AOI211_X1 U13767 ( .C1(n14357), .C2(n14542), .A(n13903), .B(n11268), .ZN(
        n11201) );
  AND2_X1 U13768 ( .A1(n13590), .A2(n13913), .ZN(n14360) );
  NOR2_X1 U13769 ( .A1(n11201), .A2(n14360), .ZN(n14664) );
  OR2_X1 U13770 ( .A1(n11207), .A2(n14537), .ZN(n14663) );
  OAI22_X1 U13771 ( .A1(n13930), .A2(n14663), .B1(n14364), .B2(n13857), .ZN(
        n11203) );
  NOR2_X1 U13772 ( .A1(n11260), .A2(n14573), .ZN(n11202) );
  AOI211_X1 U13773 ( .C1(n13930), .C2(P1_REG2_REG_10__SCAN_IN), .A(n11203), 
        .B(n11202), .ZN(n11204) );
  OAI21_X1 U13774 ( .B1(n14664), .B2(n13927), .A(n11204), .ZN(n11211) );
  NAND2_X1 U13775 ( .A1(n11206), .A2(n11205), .ZN(n14533) );
  NOR2_X1 U13776 ( .A1(n11209), .A2(n11208), .ZN(n14668) );
  INV_X1 U13777 ( .A(n11262), .ZN(n14667) );
  INV_X1 U13778 ( .A(n13863), .ZN(n13911) );
  NOR3_X1 U13779 ( .A1(n14668), .A2(n14667), .A3(n13911), .ZN(n11210) );
  AOI211_X1 U13780 ( .C1(n14672), .C2(n14175), .A(n11211), .B(n11210), .ZN(
        n11212) );
  INV_X1 U13781 ( .A(n11212), .ZN(P1_U3283) );
  NAND2_X1 U13782 ( .A1(n11356), .A2(n13475), .ZN(n11214) );
  NAND2_X1 U13783 ( .A1(n13590), .A2(n13445), .ZN(n11213) );
  NAND2_X1 U13784 ( .A1(n11214), .A2(n11213), .ZN(n11215) );
  XNOR2_X1 U13785 ( .A(n11215), .B(n11318), .ZN(n11313) );
  AND2_X1 U13786 ( .A1(n13478), .A2(n13590), .ZN(n11216) );
  AOI21_X1 U13787 ( .B1(n11356), .B2(n13445), .A(n11216), .ZN(n11312) );
  XNOR2_X1 U13788 ( .A(n11313), .B(n11312), .ZN(n11238) );
  AOI21_X1 U13789 ( .B1(n11221), .B2(n11218), .A(n11217), .ZN(n11219) );
  NAND2_X1 U13790 ( .A1(n11220), .A2(n11219), .ZN(n11225) );
  INV_X1 U13791 ( .A(n11221), .ZN(n11223) );
  NAND2_X1 U13792 ( .A1(n11223), .A2(n11222), .ZN(n11224) );
  NAND2_X1 U13793 ( .A1(n11225), .A2(n11224), .ZN(n14353) );
  NAND2_X1 U13794 ( .A1(n14357), .A2(n13475), .ZN(n11227) );
  NAND2_X1 U13795 ( .A1(n13591), .A2(n13445), .ZN(n11226) );
  NAND2_X1 U13796 ( .A1(n11227), .A2(n11226), .ZN(n11228) );
  XNOR2_X1 U13797 ( .A(n11228), .B(n13476), .ZN(n11232) );
  AND2_X1 U13798 ( .A1(n13478), .A2(n13591), .ZN(n11229) );
  AOI21_X1 U13799 ( .B1(n14357), .B2(n13445), .A(n11229), .ZN(n11230) );
  XNOR2_X1 U13800 ( .A(n11232), .B(n11230), .ZN(n14352) );
  NAND2_X1 U13801 ( .A1(n14353), .A2(n14352), .ZN(n14349) );
  INV_X1 U13802 ( .A(n11230), .ZN(n11231) );
  NAND2_X1 U13803 ( .A1(n11232), .A2(n11231), .ZN(n11233) );
  NAND2_X1 U13804 ( .A1(n14349), .A2(n11233), .ZN(n11237) );
  INV_X1 U13805 ( .A(n11237), .ZN(n11235) );
  INV_X1 U13806 ( .A(n11238), .ZN(n11234) );
  INV_X1 U13807 ( .A(n11315), .ZN(n11236) );
  AOI21_X1 U13808 ( .B1(n11238), .B2(n11237), .A(n11236), .ZN(n11244) );
  INV_X1 U13809 ( .A(n13591), .ZN(n14538) );
  NAND2_X1 U13810 ( .A1(n13573), .A2(n11269), .ZN(n11241) );
  AOI22_X1 U13811 ( .A1(n11239), .A2(n13589), .B1(P1_REG3_REG_11__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11240) );
  OAI211_X1 U13812 ( .C1(n14538), .C2(n13493), .A(n11241), .B(n11240), .ZN(
        n11242) );
  AOI21_X1 U13813 ( .B1(n11356), .B2(n14358), .A(n11242), .ZN(n11243) );
  OAI21_X1 U13814 ( .B1(n11244), .B2(n13564), .A(n11243), .ZN(P1_U3236) );
  XNOR2_X1 U13815 ( .A(n11934), .B(n11245), .ZN(n12084) );
  XNOR2_X1 U13816 ( .A(n11246), .B(n12084), .ZN(n11247) );
  NAND2_X1 U13817 ( .A1(n11247), .A2(n14304), .ZN(n11250) );
  NAND2_X1 U13818 ( .A1(n12931), .A2(n12902), .ZN(n11249) );
  NAND2_X1 U13819 ( .A1(n12933), .A2(n12901), .ZN(n11248) );
  AND2_X1 U13820 ( .A1(n11249), .A2(n11248), .ZN(n11300) );
  NAND2_X1 U13821 ( .A1(n11250), .A2(n11300), .ZN(n14326) );
  INV_X1 U13822 ( .A(n14326), .ZN(n11257) );
  XNOR2_X1 U13823 ( .A(n11251), .B(n12084), .ZN(n14328) );
  OAI211_X1 U13824 ( .C1(n14325), .C2(n11252), .A(n14313), .B(n14311), .ZN(
        n14324) );
  AOI22_X1 U13825 ( .A1(n13216), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n11302), 
        .B2(n14841), .ZN(n11254) );
  NAND2_X1 U13826 ( .A1(n11934), .A2(n14307), .ZN(n11253) );
  OAI211_X1 U13827 ( .C1(n14324), .C2(n13213), .A(n11254), .B(n11253), .ZN(
        n11255) );
  AOI21_X1 U13828 ( .B1(n14328), .B2(n14316), .A(n11255), .ZN(n11256) );
  OAI21_X1 U13829 ( .B1(n11257), .B2(n13216), .A(n11256), .ZN(P2_U3252) );
  OR2_X1 U13830 ( .A1(n14357), .A2(n13591), .ZN(n11259) );
  XNOR2_X1 U13831 ( .A(n11354), .B(n11353), .ZN(n14398) );
  INV_X1 U13832 ( .A(n14398), .ZN(n11275) );
  NAND2_X1 U13833 ( .A1(n11260), .A2(n13591), .ZN(n11261) );
  INV_X1 U13834 ( .A(n11353), .ZN(n11263) );
  OAI211_X1 U13835 ( .C1(n11264), .C2(n11263), .A(n11358), .B(n14554), .ZN(
        n11266) );
  AOI22_X1 U13836 ( .A1(n13854), .A2(n13591), .B1(n13589), .B2(n13913), .ZN(
        n11265) );
  NAND2_X1 U13837 ( .A1(n11266), .A2(n11265), .ZN(n14396) );
  INV_X1 U13838 ( .A(n11356), .ZN(n14395) );
  NOR2_X1 U13839 ( .A1(n11267), .A2(n11356), .ZN(n11363) );
  INV_X1 U13840 ( .A(n11363), .ZN(n11364) );
  OAI211_X1 U13841 ( .C1(n14395), .C2(n11268), .A(n11364), .B(n14561), .ZN(
        n14394) );
  INV_X1 U13842 ( .A(n11269), .ZN(n11270) );
  OAI22_X1 U13843 ( .A1(n13902), .A2(n10425), .B1(n11270), .B2(n13857), .ZN(
        n11271) );
  AOI21_X1 U13844 ( .B1(n11356), .B2(n14557), .A(n11271), .ZN(n11272) );
  OAI21_X1 U13845 ( .B1(n14394), .B2(n13927), .A(n11272), .ZN(n11273) );
  AOI21_X1 U13846 ( .B1(n14396), .B2(n13902), .A(n11273), .ZN(n11274) );
  OAI21_X1 U13847 ( .B1(n13896), .B2(n11275), .A(n11274), .ZN(P1_U3282) );
  INV_X1 U13848 ( .A(n11276), .ZN(n11279) );
  AOI211_X1 U13849 ( .C1(n11279), .C2(n14918), .A(n11278), .B(n11277), .ZN(
        n11284) );
  AOI22_X1 U13850 ( .A1(n11919), .A2(n13304), .B1(n14932), .B2(
        P2_REG1_REG_11__SCAN_IN), .ZN(n11280) );
  OAI21_X1 U13851 ( .B1(n11284), .B2(n14932), .A(n11280), .ZN(P2_U3510) );
  INV_X1 U13852 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n11281) );
  NOR2_X1 U13853 ( .A1(n14924), .A2(n11281), .ZN(n11282) );
  AOI21_X1 U13854 ( .B1(n11919), .B2(n8982), .A(n11282), .ZN(n11283) );
  OAI21_X1 U13855 ( .B1(n11284), .B2(n14922), .A(n11283), .ZN(P2_U3463) );
  NAND2_X1 U13856 ( .A1(n11286), .A2(n11285), .ZN(n11287) );
  NAND2_X1 U13857 ( .A1(n11288), .A2(n11287), .ZN(n11294) );
  XNOR2_X1 U13858 ( .A(n11934), .B(n12154), .ZN(n11289) );
  AND2_X1 U13859 ( .A1(n12932), .A2(n13049), .ZN(n11290) );
  NAND2_X1 U13860 ( .A1(n11289), .A2(n11290), .ZN(n11400) );
  INV_X1 U13861 ( .A(n11289), .ZN(n11292) );
  INV_X1 U13862 ( .A(n11290), .ZN(n11291) );
  NAND2_X1 U13863 ( .A1(n11292), .A2(n11291), .ZN(n11293) );
  NAND2_X1 U13864 ( .A1(n11400), .A2(n11293), .ZN(n11295) );
  AOI21_X1 U13865 ( .B1(n11294), .B2(n11295), .A(n12908), .ZN(n11298) );
  INV_X1 U13866 ( .A(n11294), .ZN(n11297) );
  INV_X1 U13867 ( .A(n11295), .ZN(n11296) );
  NAND2_X1 U13868 ( .A1(n11298), .A2(n11401), .ZN(n11304) );
  OAI22_X1 U13869 ( .A1(n12906), .A2(n11300), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11299), .ZN(n11301) );
  AOI21_X1 U13870 ( .B1(n11302), .B2(n12903), .A(n11301), .ZN(n11303) );
  OAI211_X1 U13871 ( .C1(n14325), .C2(n12900), .A(n11304), .B(n11303), .ZN(
        P2_U3206) );
  NAND2_X1 U13872 ( .A1(n11308), .A2(n11524), .ZN(n11306) );
  OAI211_X1 U13873 ( .C1(n11307), .C2(n14039), .A(n11306), .B(n11305), .ZN(
        P1_U3332) );
  NAND2_X1 U13874 ( .A1(n11308), .A2(n13350), .ZN(n11310) );
  OR2_X1 U13875 ( .A1(n11309), .A2(P2_U3088), .ZN(n12108) );
  OAI211_X1 U13876 ( .C1(n11311), .C2(n13357), .A(n11310), .B(n12108), .ZN(
        P2_U3304) );
  INV_X1 U13877 ( .A(n14156), .ZN(n11368) );
  NAND2_X1 U13878 ( .A1(n11313), .A2(n11312), .ZN(n11314) );
  NAND2_X1 U13879 ( .A1(n14156), .A2(n13475), .ZN(n11317) );
  NAND2_X1 U13880 ( .A1(n13589), .A2(n13445), .ZN(n11316) );
  NAND2_X1 U13881 ( .A1(n11317), .A2(n11316), .ZN(n11319) );
  XNOR2_X1 U13882 ( .A(n11319), .B(n11318), .ZN(n11383) );
  AND2_X1 U13883 ( .A1(n13478), .A2(n13589), .ZN(n11320) );
  AOI21_X1 U13884 ( .B1(n14156), .B2(n13445), .A(n11320), .ZN(n11384) );
  XNOR2_X1 U13885 ( .A(n11383), .B(n11384), .ZN(n11322) );
  AOI21_X1 U13886 ( .B1(n11321), .B2(n11322), .A(n13564), .ZN(n11324) );
  INV_X1 U13887 ( .A(n11322), .ZN(n11323) );
  NAND2_X1 U13888 ( .A1(n11324), .A2(n11388), .ZN(n11330) );
  NAND2_X1 U13889 ( .A1(n13590), .A2(n13854), .ZN(n11326) );
  NAND2_X1 U13890 ( .A1(n13588), .A2(n13913), .ZN(n11325) );
  AND2_X1 U13891 ( .A1(n11326), .A2(n11325), .ZN(n11361) );
  OAI21_X1 U13892 ( .B1(n11361), .B2(n13546), .A(n11327), .ZN(n11328) );
  AOI21_X1 U13893 ( .B1(n13573), .B2(n11365), .A(n11328), .ZN(n11329) );
  OAI211_X1 U13894 ( .C1(n11368), .C2(n13576), .A(n11330), .B(n11329), .ZN(
        P1_U3224) );
  AOI22_X1 U13895 ( .A1(n11331), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n11525), .ZN(n11332) );
  OAI21_X1 U13896 ( .B1(n11334), .B2(n10724), .A(n11332), .ZN(P1_U3331) );
  OAI222_X1 U13897 ( .A1(n11335), .A2(P2_U3088), .B1(n13359), .B2(n11334), 
        .C1(n11333), .C2(n13357), .ZN(P2_U3303) );
  NAND2_X1 U13898 ( .A1(n11337), .A2(n11336), .ZN(n11338) );
  XNOR2_X1 U13899 ( .A(n11609), .B(n12273), .ZN(n11340) );
  XNOR2_X1 U13900 ( .A(n11340), .B(n12400), .ZN(n12243) );
  XNOR2_X1 U13901 ( .A(n14288), .B(n12273), .ZN(n11475) );
  XNOR2_X1 U13902 ( .A(n14274), .B(n12220), .ZN(n11341) );
  NAND2_X1 U13903 ( .A1(n11341), .A2(n12398), .ZN(n11480) );
  OAI21_X1 U13904 ( .B1(n12249), .B2(n11475), .A(n11480), .ZN(n11345) );
  NAND3_X1 U13905 ( .A1(n11480), .A2(n12249), .A3(n11475), .ZN(n11343) );
  INV_X1 U13906 ( .A(n11341), .ZN(n11342) );
  NAND2_X1 U13907 ( .A1(n11342), .A2(n11430), .ZN(n11479) );
  AND2_X1 U13908 ( .A1(n11343), .A2(n11479), .ZN(n11344) );
  OAI21_X1 U13909 ( .B1(n11477), .B2(n11345), .A(n11344), .ZN(n11452) );
  XNOR2_X1 U13910 ( .A(n11350), .B(n12273), .ZN(n11451) );
  XNOR2_X1 U13911 ( .A(n11451), .B(n11483), .ZN(n11346) );
  XNOR2_X1 U13912 ( .A(n11452), .B(n11346), .ZN(n11352) );
  OAI22_X1 U13913 ( .A1(n11430), .A2(n15119), .B1(n11631), .B2(n15117), .ZN(
        n14256) );
  INV_X1 U13914 ( .A(n12378), .ZN(n12356) );
  AOI22_X1 U13915 ( .A1(n14256), .A2(n12356), .B1(P3_REG3_REG_13__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11347) );
  OAI21_X1 U13916 ( .B1(n11348), .B2(n12358), .A(n11347), .ZN(n11349) );
  AOI21_X1 U13917 ( .B1(n11350), .B2(n12380), .A(n11349), .ZN(n11351) );
  OAI21_X1 U13918 ( .B1(n11352), .B2(n12382), .A(n11351), .ZN(P3_U3174) );
  XNOR2_X1 U13919 ( .A(n11422), .B(n11359), .ZN(n14158) );
  NAND2_X1 U13920 ( .A1(n11360), .A2(n11359), .ZN(n11410) );
  OAI211_X1 U13921 ( .C1(n11360), .C2(n11359), .A(n11410), .B(n14554), .ZN(
        n11362) );
  NAND2_X1 U13922 ( .A1(n11362), .A2(n11361), .ZN(n14154) );
  AND2_X2 U13923 ( .A1(n11363), .A2(n11368), .ZN(n14173) );
  AOI211_X1 U13924 ( .C1(n14156), .C2(n11364), .A(n13903), .B(n14173), .ZN(
        n14155) );
  NAND2_X1 U13925 ( .A1(n14155), .A2(n14567), .ZN(n11367) );
  AOI22_X1 U13926 ( .A1(n14570), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n11365), 
        .B2(n14569), .ZN(n11366) );
  OAI211_X1 U13927 ( .C1(n11368), .C2(n14573), .A(n11367), .B(n11366), .ZN(
        n11369) );
  AOI21_X1 U13928 ( .B1(n14154), .B2(n13902), .A(n11369), .ZN(n11370) );
  OAI21_X1 U13929 ( .B1(n13785), .B2(n14158), .A(n11370), .ZN(P1_U3281) );
  AOI21_X1 U13930 ( .B1(n11372), .B2(n11371), .A(n14264), .ZN(n11374) );
  OR2_X1 U13931 ( .A1(n11483), .A2(n15119), .ZN(n11373) );
  OAI21_X1 U13932 ( .B1(n12192), .B2(n15117), .A(n11373), .ZN(n11453) );
  AOI21_X1 U13933 ( .B1(n11374), .B2(n11442), .A(n11453), .ZN(n11467) );
  INV_X1 U13934 ( .A(n11474), .ZN(n11632) );
  INV_X1 U13935 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n11376) );
  INV_X1 U13936 ( .A(n11454), .ZN(n11375) );
  OAI22_X1 U13937 ( .A1(n12657), .A2(n11376), .B1(n11375), .B2(n14270), .ZN(
        n11377) );
  AOI21_X1 U13938 ( .B1(n11632), .B2(n12640), .A(n11377), .ZN(n11382) );
  XNOR2_X1 U13939 ( .A(n11378), .B(n11735), .ZN(n11466) );
  NAND2_X1 U13940 ( .A1(n12657), .A2(n11379), .ZN(n11380) );
  NAND2_X1 U13941 ( .A1(n11466), .A2(n15600), .ZN(n11381) );
  OAI211_X1 U13942 ( .C1(n11467), .C2(n15595), .A(n11382), .B(n11381), .ZN(
        P3_U3219) );
  INV_X1 U13943 ( .A(n11383), .ZN(n11386) );
  INV_X1 U13944 ( .A(n11384), .ZN(n11385) );
  NAND2_X1 U13945 ( .A1(n11386), .A2(n11385), .ZN(n11387) );
  NAND2_X1 U13946 ( .A1(n14169), .A2(n13475), .ZN(n11390) );
  NAND2_X1 U13947 ( .A1(n13588), .A2(n13445), .ZN(n11389) );
  NAND2_X1 U13948 ( .A1(n11390), .A2(n11389), .ZN(n11391) );
  XNOR2_X1 U13949 ( .A(n11391), .B(n13476), .ZN(n13377) );
  AND2_X1 U13950 ( .A1(n13478), .A2(n13588), .ZN(n11392) );
  AOI21_X1 U13951 ( .B1(n14169), .B2(n13445), .A(n11392), .ZN(n13375) );
  XNOR2_X1 U13952 ( .A(n13377), .B(n13375), .ZN(n11393) );
  NAND2_X1 U13953 ( .A1(n11394), .A2(n11393), .ZN(n13379) );
  OAI211_X1 U13954 ( .C1(n11394), .C2(n11393), .A(n13379), .B(n14350), .ZN(
        n11399) );
  OR2_X1 U13955 ( .A1(n13912), .A2(n14539), .ZN(n11396) );
  NAND2_X1 U13956 ( .A1(n13589), .A2(n13854), .ZN(n11395) );
  AND2_X1 U13957 ( .A1(n11396), .A2(n11395), .ZN(n14166) );
  NAND2_X1 U13958 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n14450)
         );
  OAI21_X1 U13959 ( .B1(n14166), .B2(n13546), .A(n14450), .ZN(n11397) );
  AOI21_X1 U13960 ( .B1(n14168), .B2(n13573), .A(n11397), .ZN(n11398) );
  OAI211_X1 U13961 ( .C1(n14391), .C2(n13576), .A(n11399), .B(n11398), .ZN(
        P1_U3234) );
  XNOR2_X1 U13962 ( .A(n14308), .B(n12154), .ZN(n12109) );
  NAND2_X1 U13963 ( .A1(n12931), .A2(n13049), .ZN(n12110) );
  XNOR2_X1 U13964 ( .A(n12109), .B(n12110), .ZN(n11402) );
  OAI21_X1 U13965 ( .B1(n11403), .B2(n11402), .A(n12113), .ZN(n11404) );
  NAND2_X1 U13966 ( .A1(n11404), .A2(n12887), .ZN(n11408) );
  AOI22_X1 U13967 ( .A1(n12902), .A2(n12930), .B1(n12932), .B2(n12901), .ZN(
        n14302) );
  OAI22_X1 U13968 ( .A1(n12906), .A2(n14302), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11405), .ZN(n11406) );
  AOI21_X1 U13969 ( .B1(n14306), .B2(n12903), .A(n11406), .ZN(n11407) );
  OAI211_X1 U13970 ( .C1(n7218), .C2(n12900), .A(n11408), .B(n11407), .ZN(
        P2_U3187) );
  NAND2_X1 U13971 ( .A1(n11410), .A2(n11409), .ZN(n14165) );
  INV_X1 U13972 ( .A(n14171), .ZN(n14164) );
  NAND2_X1 U13973 ( .A1(n14165), .A2(n14164), .ZN(n14163) );
  NAND2_X1 U13974 ( .A1(n11412), .A2(n11426), .ZN(n11781) );
  OAI21_X1 U13975 ( .B1(n11412), .B2(n11426), .A(n11781), .ZN(n14387) );
  NAND2_X1 U13976 ( .A1(n14172), .A2(n14383), .ZN(n11413) );
  NAND2_X1 U13977 ( .A1(n11413), .A2(n14561), .ZN(n11414) );
  NOR2_X1 U13978 ( .A1(n6771), .A2(n11414), .ZN(n14381) );
  INV_X1 U13979 ( .A(n14383), .ZN(n11419) );
  OAI22_X1 U13980 ( .A1(n11415), .A2(n14537), .B1(n13899), .B2(n14539), .ZN(
        n14382) );
  AOI22_X1 U13981 ( .A1(n13902), .A2(n14382), .B1(n11416), .B2(n14569), .ZN(
        n11418) );
  NAND2_X1 U13982 ( .A1(n14570), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11417) );
  OAI211_X1 U13983 ( .C1(n11419), .C2(n14573), .A(n11418), .B(n11417), .ZN(
        n11420) );
  AOI21_X1 U13984 ( .B1(n14381), .B2(n14567), .A(n11420), .ZN(n11429) );
  NAND2_X1 U13985 ( .A1(n11422), .A2(n11421), .ZN(n11424) );
  OR2_X1 U13986 ( .A1(n14156), .A2(n13589), .ZN(n11423) );
  NAND2_X1 U13987 ( .A1(n11424), .A2(n11423), .ZN(n14170) );
  OR2_X1 U13988 ( .A1(n14169), .A2(n13588), .ZN(n11425) );
  NAND2_X1 U13989 ( .A1(n11427), .A2(n11426), .ZN(n14384) );
  NAND3_X1 U13990 ( .A1(n7679), .A2(n14384), .A3(n14175), .ZN(n11428) );
  OAI211_X1 U13991 ( .C1(n14387), .C2(n13911), .A(n11429), .B(n11428), .ZN(
        P1_U3279) );
  XOR2_X1 U13992 ( .A(n11475), .B(n11477), .Z(n11478) );
  XNOR2_X1 U13993 ( .A(n11478), .B(n12249), .ZN(n11437) );
  INV_X1 U13994 ( .A(n15590), .ZN(n11434) );
  OR2_X1 U13995 ( .A1(n11430), .A2(n15117), .ZN(n11432) );
  NAND2_X1 U13996 ( .A1(n12400), .A2(n12374), .ZN(n11431) );
  NAND2_X1 U13997 ( .A1(n11432), .A2(n11431), .ZN(n14292) );
  AOI22_X1 U13998 ( .A1(n14292), .A2(n12356), .B1(P3_REG3_REG_11__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11433) );
  OAI21_X1 U13999 ( .B1(n11434), .B2(n12358), .A(n11433), .ZN(n11435) );
  AOI21_X1 U14000 ( .B1(n14288), .B2(n12380), .A(n11435), .ZN(n11436) );
  OAI21_X1 U14001 ( .B1(n11437), .B2(n12382), .A(n11436), .ZN(P3_U3176) );
  OAI21_X1 U14002 ( .B1(n11439), .B2(n11441), .A(n11438), .ZN(n11517) );
  INV_X1 U14003 ( .A(n11517), .ZN(n11450) );
  NAND3_X1 U14004 ( .A1(n11442), .A2(n11441), .A3(n11440), .ZN(n11443) );
  NAND3_X1 U14005 ( .A1(n11507), .A2(n15122), .A3(n11443), .ZN(n11446) );
  OR2_X1 U14006 ( .A1(n11631), .A2(n15119), .ZN(n11444) );
  OAI21_X1 U14007 ( .B1(n12326), .B2(n15117), .A(n11444), .ZN(n11495) );
  INV_X1 U14008 ( .A(n11495), .ZN(n11445) );
  NAND2_X1 U14009 ( .A1(n11446), .A2(n11445), .ZN(n11516) );
  INV_X1 U14010 ( .A(n11499), .ZN(n11522) );
  AOI22_X1 U14011 ( .A1(n15595), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15591), 
        .B2(n11494), .ZN(n11447) );
  OAI21_X1 U14012 ( .B1(n11522), .B2(n15593), .A(n11447), .ZN(n11448) );
  AOI21_X1 U14013 ( .B1(n11516), .B2(n12657), .A(n11448), .ZN(n11449) );
  OAI21_X1 U14014 ( .B1(n11450), .B2(n12659), .A(n11449), .ZN(P3_U3218) );
  XNOR2_X1 U14015 ( .A(n11474), .B(n12273), .ZN(n11491) );
  XNOR2_X1 U14016 ( .A(n11491), .B(n11631), .ZN(n11489) );
  XOR2_X1 U14017 ( .A(n11489), .B(n11490), .Z(n11459) );
  AOI22_X1 U14018 ( .A1(n11453), .A2(n12356), .B1(P3_REG3_REG_14__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11456) );
  NAND2_X1 U14019 ( .A1(n12376), .A2(n11454), .ZN(n11455) );
  OAI211_X1 U14020 ( .C1(n11474), .C2(n12352), .A(n11456), .B(n11455), .ZN(
        n11457) );
  INV_X1 U14021 ( .A(n11457), .ZN(n11458) );
  OAI21_X1 U14022 ( .B1(n11459), .B2(n12382), .A(n11458), .ZN(P3_U3155) );
  INV_X1 U14023 ( .A(n11460), .ZN(n11464) );
  OAI222_X1 U14024 ( .A1(n13357), .A2(n11462), .B1(n13359), .B2(n11464), .C1(
        n11461), .C2(P2_U3088), .ZN(P2_U3302) );
  INV_X1 U14025 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n11465) );
  OAI222_X1 U14026 ( .A1(n14039), .A2(n11465), .B1(n10724), .B2(n11464), .C1(
        P1_U3086), .C2(n11463), .ZN(P1_U3330) );
  INV_X1 U14027 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n11469) );
  NAND2_X1 U14028 ( .A1(n11466), .A2(n14289), .ZN(n11468) );
  AND2_X1 U14029 ( .A1(n11468), .A2(n11467), .ZN(n11472) );
  MUX2_X1 U14030 ( .A(n11469), .B(n11472), .S(n15202), .Z(n11470) );
  OAI21_X1 U14031 ( .B1(n12721), .B2(n11474), .A(n11470), .ZN(P3_U3473) );
  INV_X1 U14032 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n11471) );
  MUX2_X1 U14033 ( .A(n11472), .B(n11471), .S(n15183), .Z(n11473) );
  OAI21_X1 U14034 ( .B1(n12771), .B2(n11474), .A(n11473), .ZN(P3_U3432) );
  INV_X1 U14035 ( .A(n11475), .ZN(n11476) );
  OAI22_X1 U14036 ( .A1(n11478), .A2(n12399), .B1(n11477), .B2(n11476), .ZN(
        n11482) );
  NAND2_X1 U14037 ( .A1(n11480), .A2(n11479), .ZN(n11481) );
  XNOR2_X1 U14038 ( .A(n11482), .B(n11481), .ZN(n11488) );
  OR2_X1 U14039 ( .A1(n11483), .A2(n15117), .ZN(n11484) );
  OAI21_X1 U14040 ( .B1(n12249), .B2(n15119), .A(n11484), .ZN(n14266) );
  AOI22_X1 U14041 ( .A1(n14266), .A2(n12356), .B1(P3_REG3_REG_12__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11485) );
  OAI21_X1 U14042 ( .B1(n14269), .B2(n12358), .A(n11485), .ZN(n11486) );
  AOI21_X1 U14043 ( .B1(n14274), .B2(n12380), .A(n11486), .ZN(n11487) );
  OAI21_X1 U14044 ( .B1(n11488), .B2(n12382), .A(n11487), .ZN(P3_U3164) );
  XNOR2_X1 U14045 ( .A(n11499), .B(n12273), .ZN(n12193) );
  XNOR2_X1 U14046 ( .A(n12193), .B(n12396), .ZN(n12190) );
  INV_X1 U14047 ( .A(n11491), .ZN(n11492) );
  NAND2_X1 U14048 ( .A1(n11492), .A2(n11631), .ZN(n11493) );
  XOR2_X1 U14049 ( .A(n12190), .B(n12191), .Z(n11501) );
  INV_X1 U14050 ( .A(n11494), .ZN(n11497) );
  NAND2_X1 U14051 ( .A1(n11495), .A2(n12356), .ZN(n11496) );
  NAND2_X1 U14052 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n14197)
         );
  OAI211_X1 U14053 ( .C1(n11497), .C2(n12358), .A(n11496), .B(n14197), .ZN(
        n11498) );
  AOI21_X1 U14054 ( .B1(n11499), .B2(n12380), .A(n11498), .ZN(n11500) );
  OAI21_X1 U14055 ( .B1(n11501), .B2(n12382), .A(n11500), .ZN(P3_U3181) );
  OAI21_X1 U14056 ( .B1(n11503), .B2(n11737), .A(n11502), .ZN(n12718) );
  INV_X1 U14057 ( .A(n12718), .ZN(n11515) );
  NAND3_X1 U14058 ( .A1(n11507), .A2(n11737), .A3(n11506), .ZN(n11508) );
  NAND3_X1 U14059 ( .A1(n11505), .A2(n15122), .A3(n11508), .ZN(n11511) );
  OR2_X1 U14060 ( .A1(n12199), .A2(n15117), .ZN(n11509) );
  OAI21_X1 U14061 ( .B1(n12192), .B2(n15119), .A(n11509), .ZN(n12313) );
  INV_X1 U14062 ( .A(n12313), .ZN(n11510) );
  NAND2_X1 U14063 ( .A1(n11511), .A2(n11510), .ZN(n12717) );
  INV_X1 U14064 ( .A(n12317), .ZN(n12772) );
  AOI22_X1 U14065 ( .A1(n15595), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15591), 
        .B2(n12312), .ZN(n11512) );
  OAI21_X1 U14066 ( .B1(n12772), .B2(n15593), .A(n11512), .ZN(n11513) );
  AOI21_X1 U14067 ( .B1(n12717), .B2(n12657), .A(n11513), .ZN(n11514) );
  OAI21_X1 U14068 ( .B1(n11515), .B2(n12659), .A(n11514), .ZN(P3_U3217) );
  INV_X1 U14069 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n11518) );
  AOI21_X1 U14070 ( .B1(n14289), .B2(n11517), .A(n11516), .ZN(n11520) );
  MUX2_X1 U14071 ( .A(n11518), .B(n11520), .S(n15181), .Z(n11519) );
  OAI21_X1 U14072 ( .B1(n11522), .B2(n12771), .A(n11519), .ZN(P3_U3435) );
  INV_X1 U14073 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n14194) );
  MUX2_X1 U14074 ( .A(n14194), .B(n11520), .S(n15202), .Z(n11521) );
  OAI21_X1 U14075 ( .B1(n11522), .B2(n12721), .A(n11521), .ZN(P3_U3474) );
  INV_X1 U14076 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n11523) );
  NAND3_X1 U14077 ( .A1(n11523), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n11528) );
  NAND2_X1 U14078 ( .A1(n13339), .A2(n11524), .ZN(n11527) );
  NAND2_X1 U14079 ( .A1(n11525), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n11526) );
  OAI211_X1 U14080 ( .C1(n9014), .C2(n11528), .A(n11527), .B(n11526), .ZN(
        P1_U3324) );
  INV_X1 U14081 ( .A(n11530), .ZN(n11531) );
  NAND2_X1 U14082 ( .A1(n14035), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n11533) );
  INV_X1 U14083 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n15399) );
  NAND2_X1 U14084 ( .A1(n15399), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n11536) );
  NAND2_X1 U14085 ( .A1(n11828), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n11535) );
  NAND2_X1 U14086 ( .A1(n11536), .A2(n11535), .ZN(n11547) );
  OAI21_X1 U14087 ( .B1(n11548), .B2(n11547), .A(n11536), .ZN(n11538) );
  XNOR2_X1 U14088 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n11537) );
  XNOR2_X1 U14089 ( .A(n11538), .B(n11537), .ZN(n12776) );
  NAND2_X1 U14090 ( .A1(n12776), .A2(n11549), .ZN(n11540) );
  INV_X1 U14091 ( .A(SI_31_), .ZN(n12781) );
  OR2_X1 U14092 ( .A1(n11550), .A2(n12781), .ZN(n11539) );
  NAND2_X1 U14093 ( .A1(n8828), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n11544) );
  NAND2_X1 U14094 ( .A1(n11541), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n11543) );
  NAND2_X1 U14095 ( .A1(n6640), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n11542) );
  AND3_X1 U14096 ( .A1(n11544), .A2(n11543), .A3(n11542), .ZN(n11545) );
  XNOR2_X1 U14097 ( .A(n11548), .B(n11547), .ZN(n11821) );
  NAND2_X1 U14098 ( .A1(n11821), .A2(n11549), .ZN(n11552) );
  INV_X1 U14099 ( .A(SI_30_), .ZN(n11824) );
  OR2_X1 U14100 ( .A1(n11550), .A2(n11824), .ZN(n11551) );
  NAND2_X1 U14101 ( .A1(n11552), .A2(n11551), .ZN(n12726) );
  NAND2_X1 U14102 ( .A1(n12726), .A2(n11554), .ZN(n11712) );
  NAND2_X1 U14103 ( .A1(n11713), .A2(n11712), .ZN(n11745) );
  INV_X1 U14104 ( .A(n12726), .ZN(n12665) );
  INV_X1 U14105 ( .A(n12486), .ZN(n12384) );
  OAI21_X1 U14106 ( .B1(n12665), .B2(n12384), .A(n11708), .ZN(n11553) );
  NOR2_X1 U14107 ( .A1(n11745), .A2(n11553), .ZN(n11557) );
  NAND2_X1 U14108 ( .A1(n12722), .A2(n12486), .ZN(n11556) );
  OR2_X1 U14109 ( .A1(n12726), .A2(n11554), .ZN(n11555) );
  NAND2_X1 U14110 ( .A1(n11556), .A2(n11555), .ZN(n11744) );
  INV_X1 U14111 ( .A(n11558), .ZN(n11752) );
  NOR2_X1 U14112 ( .A1(n12388), .A2(n11697), .ZN(n11679) );
  OAI21_X1 U14113 ( .B1(n11560), .B2(n11559), .A(n11697), .ZN(n11563) );
  INV_X1 U14114 ( .A(n11560), .ZN(n11561) );
  NAND3_X1 U14115 ( .A1(n11567), .A2(n11561), .A3(n11756), .ZN(n11562) );
  NAND2_X1 U14116 ( .A1(n11563), .A2(n11562), .ZN(n11564) );
  OAI211_X1 U14117 ( .C1(n11566), .C2(n11565), .A(n11564), .B(n11570), .ZN(
        n11571) );
  NAND3_X1 U14118 ( .A1(n11571), .A2(n11719), .A3(n11567), .ZN(n11569) );
  NAND3_X1 U14119 ( .A1(n11569), .A2(n11568), .A3(n11575), .ZN(n11577) );
  NAND3_X1 U14120 ( .A1(n11571), .A2(n11719), .A3(n11570), .ZN(n11574) );
  MUX2_X1 U14121 ( .A(n11577), .B(n11576), .S(n11711), .Z(n11581) );
  NAND3_X1 U14122 ( .A1(n12407), .A2(n11697), .A3(n11578), .ZN(n11579) );
  NAND2_X1 U14123 ( .A1(n12406), .A2(n15147), .ZN(n11583) );
  MUX2_X1 U14124 ( .A(n11583), .B(n11582), .S(n11697), .Z(n11584) );
  NAND2_X1 U14125 ( .A1(n11590), .A2(n11585), .ZN(n11588) );
  NAND2_X1 U14126 ( .A1(n11589), .A2(n11586), .ZN(n11587) );
  MUX2_X1 U14127 ( .A(n11588), .B(n11587), .S(n11711), .Z(n11592) );
  MUX2_X1 U14128 ( .A(n11590), .B(n11589), .S(n11697), .Z(n11591) );
  OAI211_X1 U14129 ( .C1(n11593), .C2(n11592), .A(n11718), .B(n11591), .ZN(
        n11597) );
  MUX2_X1 U14130 ( .A(n11595), .B(n11594), .S(n11711), .Z(n11596) );
  NAND3_X1 U14131 ( .A1(n11597), .A2(n11720), .A3(n11596), .ZN(n11602) );
  INV_X1 U14132 ( .A(n11728), .ZN(n11601) );
  MUX2_X1 U14133 ( .A(n11599), .B(n11598), .S(n11697), .Z(n11600) );
  NAND3_X1 U14134 ( .A1(n11602), .A2(n11601), .A3(n11600), .ZN(n11607) );
  MUX2_X1 U14135 ( .A(n11604), .B(n11603), .S(n11711), .Z(n11606) );
  AOI21_X1 U14136 ( .B1(n11607), .B2(n11606), .A(n11605), .ZN(n11614) );
  NOR2_X1 U14137 ( .A1(n12400), .A2(n11697), .ZN(n11611) );
  INV_X1 U14138 ( .A(n12400), .ZN(n11608) );
  NOR2_X1 U14139 ( .A1(n11608), .A2(n11711), .ZN(n11610) );
  MUX2_X1 U14140 ( .A(n11611), .B(n11610), .S(n11609), .Z(n11613) );
  NAND2_X1 U14141 ( .A1(n11621), .A2(n11615), .ZN(n11618) );
  NAND2_X1 U14142 ( .A1(n11620), .A2(n11616), .ZN(n11617) );
  MUX2_X1 U14143 ( .A(n11618), .B(n11617), .S(n11711), .Z(n11623) );
  INV_X1 U14144 ( .A(n11627), .ZN(n11619) );
  OR2_X1 U14145 ( .A1(n11619), .A2(n11625), .ZN(n11734) );
  INV_X1 U14146 ( .A(n11734), .ZN(n14260) );
  MUX2_X1 U14147 ( .A(n11621), .B(n11620), .S(n11697), .Z(n11622) );
  OAI211_X1 U14148 ( .C1(n11624), .C2(n11623), .A(n14260), .B(n11622), .ZN(
        n11629) );
  INV_X1 U14149 ( .A(n11625), .ZN(n11626) );
  MUX2_X1 U14150 ( .A(n11627), .B(n11626), .S(n11697), .Z(n11628) );
  AOI21_X1 U14151 ( .B1(n11629), .B2(n11628), .A(n11735), .ZN(n11636) );
  INV_X1 U14152 ( .A(n11630), .ZN(n11634) );
  NOR2_X1 U14153 ( .A1(n11632), .A2(n11631), .ZN(n11633) );
  MUX2_X1 U14154 ( .A(n11634), .B(n11633), .S(n11711), .Z(n11635) );
  NOR3_X1 U14155 ( .A1(n11636), .A2(n11635), .A3(n11732), .ZN(n11640) );
  AOI21_X1 U14156 ( .B1(n11638), .B2(n11637), .A(n11711), .ZN(n11639) );
  INV_X1 U14157 ( .A(n11641), .ZN(n11644) );
  INV_X1 U14158 ( .A(n11642), .ZN(n11643) );
  OAI21_X1 U14159 ( .B1(n11644), .B2(n11643), .A(n11711), .ZN(n11646) );
  NOR3_X1 U14160 ( .A1(n12317), .A2(n12326), .A3(n11697), .ZN(n11645) );
  AOI21_X1 U14161 ( .B1(n11647), .B2(n11646), .A(n11645), .ZN(n11652) );
  INV_X1 U14162 ( .A(n11648), .ZN(n11649) );
  NOR3_X1 U14163 ( .A1(n11662), .A2(n11649), .A3(n11697), .ZN(n11654) );
  OAI22_X1 U14164 ( .A1(n11652), .A2(n11651), .B1(n11654), .B2(n11650), .ZN(
        n11659) );
  NAND3_X1 U14165 ( .A1(n11660), .A2(n11697), .A3(n11653), .ZN(n11658) );
  INV_X1 U14166 ( .A(n11653), .ZN(n11656) );
  OAI21_X1 U14167 ( .B1(n11656), .B2(n11655), .A(n11654), .ZN(n11657) );
  AOI22_X1 U14168 ( .A1(n11659), .A2(n12633), .B1(n11658), .B2(n11657), .ZN(
        n11664) );
  INV_X1 U14169 ( .A(n11660), .ZN(n11661) );
  MUX2_X1 U14170 ( .A(n11662), .B(n11661), .S(n11711), .Z(n11663) );
  NOR2_X1 U14171 ( .A1(n11664), .A2(n11663), .ZN(n11668) );
  MUX2_X1 U14172 ( .A(n11666), .B(n11665), .S(n11697), .Z(n11667) );
  OAI211_X1 U14173 ( .C1(n11668), .C2(n12604), .A(n12593), .B(n11667), .ZN(
        n11672) );
  NAND2_X1 U14174 ( .A1(n11673), .A2(n11674), .ZN(n12579) );
  INV_X1 U14175 ( .A(n12579), .ZN(n12581) );
  MUX2_X1 U14176 ( .A(n11670), .B(n11669), .S(n11711), .Z(n11671) );
  NAND3_X1 U14177 ( .A1(n11672), .A2(n12581), .A3(n11671), .ZN(n11677) );
  MUX2_X1 U14178 ( .A(n11674), .B(n11673), .S(n11697), .Z(n11676) );
  AOI21_X1 U14179 ( .B1(n11677), .B2(n11676), .A(n11675), .ZN(n11678) );
  INV_X1 U14180 ( .A(n11680), .ZN(n11683) );
  INV_X1 U14181 ( .A(n11681), .ZN(n11682) );
  OAI21_X1 U14182 ( .B1(n11683), .B2(n11682), .A(n11685), .ZN(n11684) );
  MUX2_X1 U14183 ( .A(n11685), .B(n11684), .S(n11697), .Z(n11686) );
  OAI211_X1 U14184 ( .C1(n11687), .C2(n11717), .A(n12542), .B(n11686), .ZN(
        n11693) );
  INV_X1 U14185 ( .A(n11694), .ZN(n11688) );
  NAND2_X1 U14186 ( .A1(n11688), .A2(n11691), .ZN(n12535) );
  NOR2_X1 U14187 ( .A1(n12518), .A2(n12535), .ZN(n11741) );
  NAND3_X1 U14188 ( .A1(n11693), .A2(n11741), .A3(n11689), .ZN(n11690) );
  OAI21_X1 U14189 ( .B1(n12518), .B2(n11691), .A(n11690), .ZN(n11699) );
  NAND2_X1 U14190 ( .A1(n12523), .A2(n11694), .ZN(n11695) );
  OAI211_X1 U14191 ( .C1(n12502), .C2(n12670), .A(n11696), .B(n11695), .ZN(
        n11698) );
  MUX2_X1 U14192 ( .A(n11699), .B(n11698), .S(n11697), .Z(n11706) );
  INV_X1 U14193 ( .A(n11700), .ZN(n11704) );
  AOI21_X1 U14194 ( .B1(n11702), .B2(n11701), .A(n11704), .ZN(n11703) );
  MUX2_X1 U14195 ( .A(n11704), .B(n11703), .S(n11711), .Z(n11705) );
  INV_X1 U14196 ( .A(n11708), .ZN(n11709) );
  INV_X1 U14197 ( .A(n11713), .ZN(n11714) );
  NAND4_X1 U14198 ( .A1(n11721), .A2(n11720), .A3(n11719), .A4(n11718), .ZN(
        n11727) );
  INV_X1 U14199 ( .A(n6960), .ZN(n11724) );
  NAND4_X1 U14200 ( .A1(n11725), .A2(n11724), .A3(n11723), .A4(n11722), .ZN(
        n11726) );
  NOR4_X1 U14201 ( .A1(n11729), .A2(n11728), .A3(n11727), .A4(n11726), .ZN(
        n11731) );
  NAND4_X1 U14202 ( .A1(n11731), .A2(n14272), .A3(n11730), .A4(n14290), .ZN(
        n11733) );
  NOR4_X1 U14203 ( .A1(n11735), .A2(n11734), .A3(n11733), .A4(n11732), .ZN(
        n11736) );
  NAND4_X1 U14204 ( .A1(n12633), .A2(n12647), .A3(n11737), .A4(n11736), .ZN(
        n11738) );
  NOR4_X1 U14205 ( .A1(n12579), .A2(n12604), .A3(n12617), .A4(n11738), .ZN(
        n11739) );
  AND4_X1 U14206 ( .A1(n7374), .A2(n12593), .A3(n12567), .A4(n11739), .ZN(
        n11740) );
  NAND4_X1 U14207 ( .A1(n11741), .A2(n12507), .A3(n12542), .A4(n11740), .ZN(
        n11742) );
  XNOR2_X1 U14208 ( .A(n11746), .B(n12483), .ZN(n11748) );
  NOR4_X1 U14209 ( .A1(n11755), .A2(n11754), .A3(n11819), .A4(n11753), .ZN(
        n11758) );
  OAI21_X1 U14210 ( .B1(n11759), .B2(n11756), .A(P3_B_REG_SCAN_IN), .ZN(n11757) );
  INV_X1 U14211 ( .A(n13912), .ZN(n13587) );
  NAND2_X1 U14212 ( .A1(n14383), .A2(n13587), .ZN(n11760) );
  INV_X1 U14213 ( .A(n13899), .ZN(n13586) );
  OR2_X1 U14214 ( .A1(n14375), .A2(n13586), .ZN(n11761) );
  NAND2_X1 U14215 ( .A1(n14367), .A2(n13914), .ZN(n11762) );
  INV_X1 U14216 ( .A(n11765), .ZN(n11767) );
  INV_X1 U14217 ( .A(n13850), .ZN(n11786) );
  NAND2_X1 U14218 ( .A1(n13848), .A2(n11786), .ZN(n11769) );
  OR2_X1 U14219 ( .A1(n13852), .A2(n13584), .ZN(n11768) );
  INV_X1 U14220 ( .A(n13832), .ZN(n13840) );
  OR2_X1 U14221 ( .A1(n13995), .A2(n13827), .ZN(n11770) );
  OR2_X1 U14222 ( .A1(n13990), .A2(n13583), .ZN(n11771) );
  OR2_X1 U14223 ( .A1(n13812), .A2(n13825), .ZN(n11772) );
  NAND2_X1 U14224 ( .A1(n13979), .A2(n13582), .ZN(n11773) );
  OR2_X1 U14225 ( .A1(n13973), .A2(n13581), .ZN(n11774) );
  INV_X1 U14226 ( .A(n11794), .ZN(n13765) );
  NAND2_X1 U14227 ( .A1(n13965), .A2(n13736), .ZN(n11775) );
  INV_X1 U14228 ( .A(n13731), .ZN(n13746) );
  NAND2_X1 U14229 ( .A1(n13957), .A2(n13580), .ZN(n11776) );
  OR2_X1 U14230 ( .A1(n13951), .A2(n13737), .ZN(n11778) );
  NAND2_X1 U14231 ( .A1(n11781), .A2(n11780), .ZN(n13919) );
  INV_X1 U14232 ( .A(n14015), .ZN(n13893) );
  NAND2_X1 U14233 ( .A1(n13878), .A2(n13853), .ZN(n11785) );
  NAND2_X1 U14234 ( .A1(n13995), .A2(n13855), .ZN(n11788) );
  NAND2_X1 U14235 ( .A1(n13824), .A2(n13823), .ZN(n13822) );
  INV_X1 U14236 ( .A(n13990), .ZN(n13821) );
  NAND2_X1 U14237 ( .A1(n13821), .A2(n13583), .ZN(n11789) );
  NAND2_X1 U14238 ( .A1(n13822), .A2(n11789), .ZN(n13803) );
  INV_X1 U14239 ( .A(n13825), .ZN(n13790) );
  NAND2_X1 U14240 ( .A1(n13812), .A2(n13790), .ZN(n11790) );
  INV_X1 U14241 ( .A(n13786), .ZN(n13795) );
  NAND2_X1 U14242 ( .A1(n13979), .A2(n11791), .ZN(n11792) );
  INV_X1 U14243 ( .A(n13581), .ZN(n13789) );
  INV_X1 U14244 ( .A(n13965), .ZN(n11795) );
  INV_X1 U14245 ( .A(n13957), .ZN(n13743) );
  NOR2_X1 U14246 ( .A1(n13743), .A2(n13580), .ZN(n11796) );
  INV_X1 U14247 ( .A(n13580), .ZN(n13719) );
  NAND2_X1 U14248 ( .A1(n13709), .A2(n13579), .ZN(n11798) );
  INV_X1 U14249 ( .A(n11800), .ZN(n11801) );
  NAND2_X1 U14250 ( .A1(n13936), .A2(n13863), .ZN(n11816) );
  OR2_X2 U14251 ( .A1(n13888), .A2(n14009), .ZN(n13874) );
  NAND2_X1 U14252 ( .A1(n13851), .A2(n13995), .ZN(n13841) );
  INV_X1 U14253 ( .A(n13973), .ZN(n13781) );
  NAND2_X1 U14254 ( .A1(n13792), .A2(n13781), .ZN(n13776) );
  NOR2_X2 U14255 ( .A1(n13776), .A2(n13965), .ZN(n13759) );
  AOI21_X1 U14256 ( .B1(n13708), .B2(n13941), .A(n13903), .ZN(n11803) );
  NAND2_X1 U14257 ( .A1(n13941), .A2(n14557), .ZN(n11813) );
  NAND2_X1 U14258 ( .A1(n13579), .A2(n13854), .ZN(n13937) );
  INV_X1 U14259 ( .A(n13937), .ZN(n11810) );
  INV_X1 U14260 ( .A(P1_B_REG_SCAN_IN), .ZN(n11804) );
  NOR2_X1 U14261 ( .A1(n6641), .A2(n11804), .ZN(n11805) );
  NOR2_X1 U14262 ( .A1(n14539), .A2(n11805), .ZN(n13693) );
  NAND2_X1 U14263 ( .A1(n13693), .A2(n13577), .ZN(n13938) );
  INV_X1 U14264 ( .A(n11806), .ZN(n11807) );
  OAI22_X1 U14265 ( .A1(n11808), .A2(n13938), .B1(n13857), .B2(n11807), .ZN(
        n11809) );
  AOI21_X1 U14266 ( .B1(n13902), .B2(n11810), .A(n11809), .ZN(n11812) );
  NAND2_X1 U14267 ( .A1(n13930), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n11811) );
  NAND3_X1 U14268 ( .A1(n11813), .A2(n11812), .A3(n11811), .ZN(n11814) );
  AOI21_X1 U14269 ( .B1(n13939), .B2(n14567), .A(n11814), .ZN(n11815) );
  OAI211_X1 U14270 ( .C1(n13942), .C2(n13896), .A(n11816), .B(n11815), .ZN(
        P1_U3356) );
  INV_X1 U14271 ( .A(n11817), .ZN(n11820) );
  OAI222_X1 U14272 ( .A1(n12785), .A2(n11820), .B1(n11819), .B2(P3_U3151), 
        .C1(n11818), .C2(n12787), .ZN(P3_U3267) );
  INV_X1 U14273 ( .A(n11821), .ZN(n11823) );
  OAI222_X1 U14274 ( .A1(n12787), .A2(n11824), .B1(n12785), .B2(n11823), .C1(
        P3_U3151), .C2(n11822), .ZN(P3_U3265) );
  OAI222_X1 U14275 ( .A1(n14039), .A2(n11827), .B1(n10724), .B2(n11826), .C1(
        n11825), .C2(P1_U3086), .ZN(P1_U3335) );
  OAI222_X1 U14276 ( .A1(P1_U3086), .A2(n11829), .B1(n14039), .B2(n11828), 
        .C1(n10724), .C2(n13345), .ZN(P1_U3325) );
  INV_X1 U14277 ( .A(n11830), .ZN(n13355) );
  OAI222_X1 U14278 ( .A1(n14039), .A2(n11831), .B1(n10724), .B2(n13355), .C1(
        P1_U3086), .C2(n6641), .ZN(P1_U3328) );
  INV_X1 U14279 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n12166) );
  NOR3_X1 U14280 ( .A1(n11832), .A2(n13194), .A3(n12166), .ZN(n11835) );
  NOR2_X1 U14281 ( .A1(n11833), .A2(n14835), .ZN(n11834) );
  AOI211_X1 U14282 ( .C1(n13216), .C2(P2_REG2_REG_29__SCAN_IN), .A(n11835), 
        .B(n11834), .ZN(n11836) );
  OAI21_X1 U14283 ( .B1(n11837), .B2(n13213), .A(n11836), .ZN(n11838) );
  AOI21_X1 U14284 ( .B1(n11839), .B2(n14316), .A(n11838), .ZN(n11840) );
  OAI21_X1 U14285 ( .B1(n11841), .B2(n13216), .A(n11840), .ZN(P2_U3236) );
  NAND2_X1 U14286 ( .A1(n11843), .A2(n12051), .ZN(n11844) );
  INV_X1 U14287 ( .A(n10195), .ZN(n12059) );
  NAND3_X1 U14288 ( .A1(n11846), .A2(n12059), .A3(n11845), .ZN(n11847) );
  NAND2_X1 U14289 ( .A1(n12944), .A2(n12031), .ZN(n11850) );
  NAND2_X1 U14290 ( .A1(n11854), .A2(n12051), .ZN(n11849) );
  NAND2_X1 U14291 ( .A1(n11850), .A2(n11849), .ZN(n11856) );
  NAND2_X1 U14292 ( .A1(n12943), .A2(n12031), .ZN(n11853) );
  NAND2_X1 U14293 ( .A1(n11853), .A2(n11852), .ZN(n11858) );
  AOI22_X1 U14294 ( .A1(n12944), .A2(n12051), .B1(n12031), .B2(n11854), .ZN(
        n11855) );
  AOI21_X1 U14295 ( .B1(n11857), .B2(n11856), .A(n11855), .ZN(n11862) );
  INV_X1 U14296 ( .A(n11858), .ZN(n11861) );
  INV_X1 U14297 ( .A(n11859), .ZN(n11860) );
  NAND2_X1 U14298 ( .A1(n12942), .A2(n12031), .ZN(n11865) );
  NAND2_X1 U14299 ( .A1(n14891), .A2(n6986), .ZN(n11864) );
  AOI22_X1 U14300 ( .A1(n12942), .A2(n12051), .B1(n12031), .B2(n14891), .ZN(
        n11866) );
  NAND2_X1 U14301 ( .A1(n12941), .A2(n6986), .ZN(n11869) );
  NAND2_X1 U14302 ( .A1(n11870), .A2(n12031), .ZN(n11868) );
  NAND2_X1 U14303 ( .A1(n11869), .A2(n11868), .ZN(n11872) );
  NAND2_X1 U14304 ( .A1(n11876), .A2(n6986), .ZN(n11875) );
  NAND2_X1 U14305 ( .A1(n12940), .A2(n12031), .ZN(n11874) );
  NAND2_X1 U14306 ( .A1(n11876), .A2(n12031), .ZN(n11878) );
  NAND2_X1 U14307 ( .A1(n12940), .A2(n6986), .ZN(n11877) );
  NAND2_X1 U14308 ( .A1(n11878), .A2(n11877), .ZN(n11879) );
  NAND2_X1 U14309 ( .A1(n11884), .A2(n12031), .ZN(n11883) );
  NAND2_X1 U14310 ( .A1(n12939), .A2(n6986), .ZN(n11882) );
  NAND2_X1 U14311 ( .A1(n11884), .A2(n6986), .ZN(n11885) );
  NAND2_X1 U14312 ( .A1(n11890), .A2(n6986), .ZN(n11889) );
  NAND2_X1 U14313 ( .A1(n12938), .A2(n12031), .ZN(n11888) );
  NAND2_X1 U14314 ( .A1(n11889), .A2(n11888), .ZN(n11892) );
  AOI22_X1 U14315 ( .A1(n11890), .A2(n12031), .B1(n12938), .B2(n12051), .ZN(
        n11891) );
  NAND2_X1 U14316 ( .A1(n11895), .A2(n12031), .ZN(n11894) );
  NAND2_X1 U14317 ( .A1(n12937), .A2(n6986), .ZN(n11893) );
  NAND2_X1 U14318 ( .A1(n11894), .A2(n11893), .ZN(n11898) );
  AOI22_X1 U14319 ( .A1(n11895), .A2(n12051), .B1(n12031), .B2(n12937), .ZN(
        n11896) );
  AOI21_X1 U14320 ( .B1(n11899), .B2(n11898), .A(n11896), .ZN(n11897) );
  NAND2_X1 U14321 ( .A1(n11905), .A2(n6986), .ZN(n11901) );
  NAND2_X1 U14322 ( .A1(n12936), .A2(n12031), .ZN(n11900) );
  NAND2_X1 U14323 ( .A1(n11901), .A2(n11900), .ZN(n11913) );
  NAND2_X1 U14324 ( .A1(n11902), .A2(n12031), .ZN(n11904) );
  NAND2_X1 U14325 ( .A1(n12935), .A2(n6986), .ZN(n11903) );
  OAI211_X1 U14326 ( .C1(n12031), .C2(n11910), .A(n11904), .B(n11903), .ZN(
        n11915) );
  NAND2_X1 U14327 ( .A1(n11905), .A2(n12031), .ZN(n11906) );
  OAI21_X1 U14328 ( .B1(n11907), .B2(n12031), .A(n11906), .ZN(n11908) );
  OR3_X1 U14329 ( .A1(n11910), .A2(n11909), .A3(n12031), .ZN(n11912) );
  NAND3_X1 U14330 ( .A1(n11910), .A2(n11909), .A3(n12031), .ZN(n11911) );
  AND2_X1 U14331 ( .A1(n11912), .A2(n11911), .ZN(n11917) );
  INV_X1 U14332 ( .A(n11913), .ZN(n11914) );
  NAND2_X1 U14333 ( .A1(n11915), .A2(n11914), .ZN(n11916) );
  AND2_X1 U14334 ( .A1(n12934), .A2(n12031), .ZN(n11918) );
  AOI21_X1 U14335 ( .B1(n11919), .B2(n6986), .A(n11918), .ZN(n11923) );
  NAND2_X1 U14336 ( .A1(n11919), .A2(n12031), .ZN(n11920) );
  OAI21_X1 U14337 ( .B1(n11921), .B2(n12031), .A(n11920), .ZN(n11922) );
  OAI21_X1 U14338 ( .B1(n11924), .B2(n11923), .A(n11922), .ZN(n11926) );
  NAND2_X1 U14339 ( .A1(n11924), .A2(n11923), .ZN(n11925) );
  NAND2_X1 U14340 ( .A1(n14329), .A2(n12031), .ZN(n11928) );
  NAND2_X1 U14341 ( .A1(n12933), .A2(n6986), .ZN(n11927) );
  NAND2_X1 U14342 ( .A1(n11928), .A2(n11927), .ZN(n11930) );
  AOI22_X1 U14343 ( .A1(n14329), .A2(n6986), .B1(n12031), .B2(n12933), .ZN(
        n11929) );
  NAND2_X1 U14344 ( .A1(n11934), .A2(n6986), .ZN(n11933) );
  NAND2_X1 U14345 ( .A1(n12932), .A2(n12031), .ZN(n11932) );
  AOI22_X1 U14346 ( .A1(n11934), .A2(n12031), .B1(n12932), .B2(n12051), .ZN(
        n11935) );
  NAND2_X1 U14347 ( .A1(n14308), .A2(n12031), .ZN(n11937) );
  NAND2_X1 U14348 ( .A1(n12931), .A2(n6986), .ZN(n11936) );
  AOI22_X1 U14349 ( .A1(n14308), .A2(n12051), .B1(n12031), .B2(n12931), .ZN(
        n11938) );
  NAND2_X1 U14350 ( .A1(n13336), .A2(n6986), .ZN(n11941) );
  NAND2_X1 U14351 ( .A1(n12930), .A2(n12031), .ZN(n11940) );
  NAND2_X1 U14352 ( .A1(n11941), .A2(n11940), .ZN(n11947) );
  NAND2_X1 U14353 ( .A1(n13336), .A2(n12031), .ZN(n11942) );
  NAND2_X1 U14354 ( .A1(n11945), .A2(n11944), .ZN(n11946) );
  NAND2_X1 U14355 ( .A1(n13294), .A2(n12031), .ZN(n11950) );
  NAND2_X1 U14356 ( .A1(n12929), .A2(n6986), .ZN(n11949) );
  NAND2_X1 U14357 ( .A1(n11950), .A2(n11949), .ZN(n11952) );
  AOI22_X1 U14358 ( .A1(n13294), .A2(n6986), .B1(n12031), .B2(n12929), .ZN(
        n11951) );
  NAND2_X1 U14359 ( .A1(n13289), .A2(n12051), .ZN(n11954) );
  NAND2_X1 U14360 ( .A1(n12928), .A2(n12031), .ZN(n11953) );
  AOI22_X1 U14361 ( .A1(n13289), .A2(n12031), .B1(n12928), .B2(n12051), .ZN(
        n11955) );
  INV_X1 U14362 ( .A(n11955), .ZN(n11956) );
  NAND2_X1 U14363 ( .A1(n13283), .A2(n12031), .ZN(n11959) );
  NAND2_X1 U14364 ( .A1(n12927), .A2(n6986), .ZN(n11958) );
  NAND2_X1 U14365 ( .A1(n11959), .A2(n11958), .ZN(n11965) );
  NAND2_X1 U14366 ( .A1(n13283), .A2(n6986), .ZN(n11961) );
  NAND2_X1 U14367 ( .A1(n12927), .A2(n12031), .ZN(n11960) );
  NAND2_X1 U14368 ( .A1(n11961), .A2(n11960), .ZN(n11962) );
  NAND2_X1 U14369 ( .A1(n11963), .A2(n11962), .ZN(n11969) );
  INV_X1 U14370 ( .A(n11964), .ZN(n11967) );
  INV_X1 U14371 ( .A(n11965), .ZN(n11966) );
  NAND2_X1 U14372 ( .A1(n11967), .A2(n11966), .ZN(n11968) );
  NAND2_X1 U14373 ( .A1(n13278), .A2(n12051), .ZN(n11971) );
  NAND2_X1 U14374 ( .A1(n12926), .A2(n12031), .ZN(n11970) );
  NAND2_X1 U14375 ( .A1(n13278), .A2(n12031), .ZN(n11972) );
  NAND2_X1 U14376 ( .A1(n13273), .A2(n12031), .ZN(n11976) );
  NAND2_X1 U14377 ( .A1(n12925), .A2(n12051), .ZN(n11975) );
  NAND2_X1 U14378 ( .A1(n13273), .A2(n6986), .ZN(n11977) );
  OAI21_X1 U14379 ( .B1(n12810), .B2(n12051), .A(n11977), .ZN(n11978) );
  NAND2_X1 U14380 ( .A1(n13270), .A2(n12051), .ZN(n11980) );
  NAND2_X1 U14381 ( .A1(n12924), .A2(n12031), .ZN(n11979) );
  NAND2_X1 U14382 ( .A1(n13270), .A2(n12031), .ZN(n11981) );
  NAND2_X1 U14383 ( .A1(n13262), .A2(n12031), .ZN(n11985) );
  NAND2_X1 U14384 ( .A1(n12923), .A2(n6986), .ZN(n11984) );
  NAND2_X1 U14385 ( .A1(n11985), .A2(n11984), .ZN(n11988) );
  AOI22_X1 U14386 ( .A1(n13262), .A2(n12051), .B1(n12031), .B2(n12923), .ZN(
        n11986) );
  NAND2_X1 U14387 ( .A1(n13257), .A2(n6986), .ZN(n11991) );
  NAND2_X1 U14388 ( .A1(n12922), .A2(n12031), .ZN(n11990) );
  NAND2_X1 U14389 ( .A1(n11991), .A2(n11990), .ZN(n11993) );
  AOI22_X1 U14390 ( .A1(n13257), .A2(n12031), .B1(n12922), .B2(n12051), .ZN(
        n11992) );
  NAND2_X1 U14391 ( .A1(n13066), .A2(n12031), .ZN(n11995) );
  NAND2_X1 U14392 ( .A1(n12921), .A2(n12051), .ZN(n11994) );
  AOI22_X1 U14393 ( .A1(n13066), .A2(n6986), .B1(n12031), .B2(n12921), .ZN(
        n11996) );
  OAI22_X1 U14394 ( .A1(n13319), .A2(n12031), .B1(n12890), .B2(n12051), .ZN(
        n12000) );
  AOI22_X1 U14395 ( .A1(n13248), .A2(n12031), .B1(n12920), .B2(n6986), .ZN(
        n11997) );
  INV_X1 U14396 ( .A(n11998), .ZN(n12004) );
  INV_X1 U14397 ( .A(n11999), .ZN(n12002) );
  INV_X1 U14398 ( .A(n12000), .ZN(n12001) );
  AOI22_X1 U14399 ( .A1(n13238), .A2(n12031), .B1(n12919), .B2(n12051), .ZN(
        n12033) );
  OAI22_X1 U14400 ( .A1(n13036), .A2(n12031), .B1(n12828), .B2(n12051), .ZN(
        n12032) );
  AOI21_X1 U14401 ( .B1(n12004), .B2(n12003), .A(n7686), .ZN(n12035) );
  INV_X1 U14402 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n12005) );
  OR2_X1 U14403 ( .A1(n12013), .A2(n12005), .ZN(n12006) );
  INV_X1 U14404 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n15447) );
  NAND2_X1 U14405 ( .A1(n12007), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n12010) );
  NAND2_X1 U14406 ( .A1(n12008), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n12009) );
  OAI211_X1 U14407 ( .C1(n7792), .C2(n15447), .A(n12010), .B(n12009), .ZN(
        n12992) );
  XNOR2_X1 U14408 ( .A(n12989), .B(n12992), .ZN(n12041) );
  OR2_X1 U14409 ( .A1(n12013), .A2(n15399), .ZN(n12014) );
  OAI211_X1 U14410 ( .C1(n8342), .C2(n12058), .A(n12098), .B(n12056), .ZN(
        n12015) );
  AOI21_X1 U14411 ( .B1(n12992), .B2(n6986), .A(n12015), .ZN(n12016) );
  NOR2_X1 U14412 ( .A1(n12016), .A2(n12018), .ZN(n12017) );
  AOI21_X1 U14413 ( .B1(n13224), .B2(n12031), .A(n12017), .ZN(n12037) );
  NAND2_X1 U14414 ( .A1(n13224), .A2(n6986), .ZN(n12020) );
  INV_X1 U14415 ( .A(n12018), .ZN(n12915) );
  NAND2_X1 U14416 ( .A1(n12915), .A2(n12031), .ZN(n12019) );
  NAND2_X1 U14417 ( .A1(n12020), .A2(n12019), .ZN(n12036) );
  AND2_X1 U14418 ( .A1(n12916), .A2(n6986), .ZN(n12021) );
  AOI21_X1 U14419 ( .B1(n12022), .B2(n12031), .A(n12021), .ZN(n12043) );
  NAND2_X1 U14420 ( .A1(n12022), .A2(n6986), .ZN(n12024) );
  NAND2_X1 U14421 ( .A1(n12916), .A2(n12031), .ZN(n12023) );
  NAND2_X1 U14422 ( .A1(n12024), .A2(n12023), .ZN(n12042) );
  OAI22_X1 U14423 ( .A1(n12037), .A2(n12036), .B1(n12043), .B2(n12042), .ZN(
        n12025) );
  AND2_X1 U14424 ( .A1(n12917), .A2(n12031), .ZN(n12026) );
  AOI21_X1 U14425 ( .B1(n13229), .B2(n6986), .A(n12026), .ZN(n12045) );
  NAND2_X1 U14426 ( .A1(n13229), .A2(n12031), .ZN(n12029) );
  NAND2_X1 U14427 ( .A1(n12917), .A2(n6986), .ZN(n12028) );
  NAND2_X1 U14428 ( .A1(n12029), .A2(n12028), .ZN(n12044) );
  NAND2_X1 U14429 ( .A1(n12045), .A2(n12044), .ZN(n12030) );
  OAI22_X1 U14430 ( .A1(n13019), .A2(n12031), .B1(n12892), .B2(n12051), .ZN(
        n12039) );
  AOI22_X1 U14431 ( .A1(n13232), .A2(n12031), .B1(n12918), .B2(n6986), .ZN(
        n12040) );
  OAI22_X1 U14432 ( .A1(n12039), .A2(n12040), .B1(n12033), .B2(n12032), .ZN(
        n12034) );
  INV_X1 U14433 ( .A(n12041), .ZN(n12097) );
  INV_X1 U14434 ( .A(n12042), .ZN(n12047) );
  INV_X1 U14435 ( .A(n12043), .ZN(n12046) );
  OAI22_X1 U14436 ( .A1(n12047), .A2(n12046), .B1(n12045), .B2(n12044), .ZN(
        n12049) );
  INV_X1 U14437 ( .A(n12992), .ZN(n12052) );
  NAND3_X1 U14438 ( .A1(n12989), .A2(n12052), .A3(n12051), .ZN(n12054) );
  NAND3_X1 U14439 ( .A1(n13308), .A2(n12031), .A3(n12992), .ZN(n12053) );
  OAI21_X1 U14440 ( .B1(n8343), .B2(n13195), .A(n12056), .ZN(n12057) );
  AOI21_X1 U14441 ( .B1(n12059), .B2(n12058), .A(n12057), .ZN(n12060) );
  INV_X1 U14442 ( .A(n12060), .ZN(n12063) );
  MUX2_X1 U14443 ( .A(n12105), .B(n12098), .S(n8342), .Z(n12061) );
  NAND2_X1 U14444 ( .A1(n12061), .A2(n13195), .ZN(n12062) );
  NOR2_X1 U14445 ( .A1(n14884), .A2(n12066), .ZN(n12072) );
  AND2_X1 U14446 ( .A1(n12068), .A2(n12067), .ZN(n12071) );
  NAND4_X1 U14447 ( .A1(n12072), .A2(n12071), .A3(n12070), .A4(n12069), .ZN(
        n12074) );
  NOR2_X1 U14448 ( .A1(n12074), .A2(n12073), .ZN(n12077) );
  NAND4_X1 U14449 ( .A1(n12078), .A2(n12077), .A3(n12076), .A4(n12075), .ZN(
        n12079) );
  OR4_X1 U14450 ( .A1(n12082), .A2(n12081), .A3(n12080), .A4(n12079), .ZN(
        n12083) );
  OR4_X1 U14451 ( .A1(n13198), .A2(n12085), .A3(n12084), .A4(n12083), .ZN(
        n12086) );
  NOR2_X1 U14452 ( .A1(n13167), .A2(n12086), .ZN(n12087) );
  XNOR2_X1 U14453 ( .A(n14308), .B(n12931), .ZN(n14309) );
  NAND3_X1 U14454 ( .A1(n13161), .A2(n12087), .A3(n14309), .ZN(n12088) );
  NOR4_X1 U14455 ( .A1(n13136), .A2(n12089), .A3(n13208), .A4(n12088), .ZN(
        n12090) );
  NAND3_X1 U14456 ( .A1(n12091), .A2(n12090), .A3(n13112), .ZN(n12092) );
  NOR4_X1 U14457 ( .A1(n12093), .A2(n13074), .A3(n13058), .A4(n12092), .ZN(
        n12094) );
  NOR3_X1 U14458 ( .A1(n12099), .A2(n12098), .A3(n12108), .ZN(n12100) );
  NAND4_X1 U14459 ( .A1(n14881), .A2(n12103), .A3(n12102), .A4(n12901), .ZN(
        n12104) );
  OAI211_X1 U14460 ( .C1(n12105), .C2(n12108), .A(n12104), .B(P2_B_REG_SCAN_IN), .ZN(n12106) );
  XNOR2_X1 U14461 ( .A(n13283), .B(n12154), .ZN(n12120) );
  NAND2_X1 U14462 ( .A1(n12927), .A2(n12126), .ZN(n12121) );
  XNOR2_X1 U14463 ( .A(n13289), .B(n9889), .ZN(n12119) );
  NAND2_X1 U14464 ( .A1(n12928), .A2(n12126), .ZN(n12118) );
  INV_X1 U14465 ( .A(n12109), .ZN(n12111) );
  NAND2_X1 U14466 ( .A1(n12111), .A2(n12110), .ZN(n12112) );
  XOR2_X1 U14467 ( .A(n12154), .B(n13336), .Z(n12114) );
  NAND2_X1 U14468 ( .A1(n12930), .A2(n13049), .ZN(n12909) );
  XNOR2_X1 U14469 ( .A(n13294), .B(n12154), .ZN(n12115) );
  NAND2_X1 U14470 ( .A1(n12929), .A2(n13049), .ZN(n12116) );
  XNOR2_X1 U14471 ( .A(n12115), .B(n12116), .ZN(n12833) );
  INV_X1 U14472 ( .A(n12115), .ZN(n12117) );
  NAND2_X1 U14473 ( .A1(n12117), .A2(n12116), .ZN(n12842) );
  XNOR2_X1 U14474 ( .A(n12119), .B(n12118), .ZN(n12843) );
  XNOR2_X1 U14475 ( .A(n12120), .B(n12121), .ZN(n12878) );
  XNOR2_X1 U14476 ( .A(n13278), .B(n9889), .ZN(n12123) );
  NAND2_X1 U14477 ( .A1(n12926), .A2(n13049), .ZN(n12122) );
  NOR2_X1 U14478 ( .A1(n12123), .A2(n12122), .ZN(n12806) );
  XNOR2_X1 U14479 ( .A(n13273), .B(n12154), .ZN(n12125) );
  AND2_X1 U14480 ( .A1(n12925), .A2(n13049), .ZN(n12124) );
  NAND2_X1 U14481 ( .A1(n12125), .A2(n12124), .ZN(n12860) );
  XNOR2_X1 U14482 ( .A(n13270), .B(n12154), .ZN(n12127) );
  NAND2_X1 U14483 ( .A1(n12924), .A2(n12126), .ZN(n12128) );
  XNOR2_X1 U14484 ( .A(n12127), .B(n12128), .ZN(n12816) );
  INV_X1 U14485 ( .A(n12128), .ZN(n12129) );
  XNOR2_X1 U14486 ( .A(n13262), .B(n12154), .ZN(n12131) );
  NAND2_X1 U14487 ( .A1(n12923), .A2(n13049), .ZN(n12872) );
  NOR2_X2 U14488 ( .A1(n12873), .A2(n12872), .ZN(n12871) );
  AND2_X1 U14489 ( .A1(n12132), .A2(n12131), .ZN(n12133) );
  NOR2_X2 U14490 ( .A1(n12871), .A2(n12133), .ZN(n12134) );
  XNOR2_X1 U14491 ( .A(n13257), .B(n12154), .ZN(n12135) );
  XNOR2_X1 U14492 ( .A(n12134), .B(n12135), .ZN(n12800) );
  NOR2_X1 U14493 ( .A1(n12854), .A2(n14313), .ZN(n12799) );
  NAND2_X1 U14494 ( .A1(n12800), .A2(n12799), .ZN(n12798) );
  XNOR2_X1 U14495 ( .A(n13066), .B(n9889), .ZN(n12139) );
  NAND2_X1 U14496 ( .A1(n12921), .A2(n13049), .ZN(n12138) );
  NOR2_X1 U14497 ( .A1(n12139), .A2(n12138), .ZN(n12140) );
  AOI21_X1 U14498 ( .B1(n12139), .B2(n12138), .A(n12140), .ZN(n12852) );
  INV_X1 U14499 ( .A(n12140), .ZN(n12141) );
  XNOR2_X1 U14500 ( .A(n13319), .B(n12154), .ZN(n12143) );
  NAND2_X1 U14501 ( .A1(n12920), .A2(n13049), .ZN(n12142) );
  NOR2_X1 U14502 ( .A1(n12143), .A2(n12142), .ZN(n12144) );
  AOI21_X1 U14503 ( .B1(n12143), .B2(n12142), .A(n12144), .ZN(n12826) );
  INV_X1 U14504 ( .A(n12144), .ZN(n12145) );
  XNOR2_X1 U14505 ( .A(n13238), .B(n12154), .ZN(n12146) );
  NAND2_X1 U14506 ( .A1(n12919), .A2(n13049), .ZN(n12147) );
  XNOR2_X1 U14507 ( .A(n12146), .B(n12147), .ZN(n12885) );
  INV_X1 U14508 ( .A(n12146), .ZN(n12148) );
  INV_X1 U14509 ( .A(n12790), .ZN(n12152) );
  XNOR2_X1 U14510 ( .A(n13019), .B(n9889), .ZN(n12150) );
  NOR2_X1 U14511 ( .A1(n12892), .A2(n14313), .ZN(n12149) );
  NAND2_X1 U14512 ( .A1(n12150), .A2(n12149), .ZN(n12153) );
  OAI21_X1 U14513 ( .B1(n12150), .B2(n12149), .A(n12153), .ZN(n12789) );
  NAND2_X1 U14514 ( .A1(n12152), .A2(n12151), .ZN(n12791) );
  NAND2_X1 U14515 ( .A1(n12791), .A2(n12153), .ZN(n12163) );
  NAND2_X1 U14516 ( .A1(n12917), .A2(n13049), .ZN(n12155) );
  XNOR2_X1 U14517 ( .A(n12155), .B(n12154), .ZN(n12158) );
  NOR3_X1 U14518 ( .A1(n7221), .A2(n12913), .A3(n12158), .ZN(n12156) );
  AOI21_X1 U14519 ( .B1(n7221), .B2(n12158), .A(n12156), .ZN(n12162) );
  NAND3_X1 U14520 ( .A1(n13229), .A2(n12900), .A3(n12158), .ZN(n12157) );
  OAI21_X1 U14521 ( .B1(n13229), .B2(n12158), .A(n12157), .ZN(n12159) );
  NAND2_X1 U14522 ( .A1(n12163), .A2(n12159), .ZN(n12161) );
  OAI21_X1 U14523 ( .B1(n7221), .B2(n12900), .A(n12908), .ZN(n12160) );
  OAI211_X1 U14524 ( .C1(n12163), .C2(n12162), .A(n12161), .B(n12160), .ZN(
        n12169) );
  NAND2_X1 U14525 ( .A1(n12916), .A2(n12902), .ZN(n12164) );
  OAI21_X1 U14526 ( .B1(n12892), .B2(n12889), .A(n12164), .ZN(n13005) );
  INV_X1 U14527 ( .A(n12165), .ZN(n13010) );
  OAI22_X1 U14528 ( .A1(n13010), .A2(n12894), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12166), .ZN(n12167) );
  AOI21_X1 U14529 ( .B1(n13005), .B2(n12897), .A(n12167), .ZN(n12168) );
  NAND2_X1 U14530 ( .A1(n12169), .A2(n12168), .ZN(P2_U3192) );
  OAI21_X1 U14531 ( .B1(n12170), .B2(n12172), .A(n12171), .ZN(n12173) );
  NAND2_X1 U14532 ( .A1(n12173), .A2(n14350), .ZN(n12177) );
  INV_X1 U14533 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n13600) );
  OAI22_X1 U14534 ( .A1(n12174), .A2(n13600), .B1(n13571), .B2(n10144), .ZN(
        n12175) );
  AOI21_X1 U14535 ( .B1(n13568), .B2(n10017), .A(n12175), .ZN(n12176) );
  OAI211_X1 U14536 ( .C1(n12178), .C2(n13576), .A(n12177), .B(n12176), .ZN(
        P1_U3222) );
  INV_X1 U14537 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n12180) );
  INV_X1 U14538 ( .A(n13351), .ZN(n12179) );
  OAI222_X1 U14539 ( .A1(n14039), .A2(n12180), .B1(n10724), .B2(n12179), .C1(
        P1_U3086), .C2(n9571), .ZN(P1_U3327) );
  OAI211_X1 U14540 ( .C1(n12183), .C2(n12182), .A(n12181), .B(n12282), .ZN(
        n12189) );
  AOI22_X1 U14541 ( .A1(n12380), .A2(n12184), .B1(P3_REG3_REG_7__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12188) );
  AOI22_X1 U14542 ( .A1(n12404), .A2(n12291), .B1(n12185), .B2(n12376), .ZN(
        n12187) );
  NAND2_X1 U14543 ( .A1(n12402), .A2(n12289), .ZN(n12186) );
  NAND4_X1 U14544 ( .A1(n12189), .A2(n12188), .A3(n12187), .A4(n12186), .ZN(
        P3_U3153) );
  XNOR2_X1 U14545 ( .A(n12670), .B(n12273), .ZN(n12270) );
  XNOR2_X1 U14546 ( .A(n12270), .B(n12386), .ZN(n12271) );
  NAND2_X1 U14547 ( .A1(n12193), .A2(n12192), .ZN(n12194) );
  XNOR2_X1 U14548 ( .A(n12317), .B(n12273), .ZN(n12195) );
  XNOR2_X1 U14549 ( .A(n12195), .B(n12395), .ZN(n12311) );
  NAND2_X1 U14550 ( .A1(n12310), .A2(n12311), .ZN(n12197) );
  NAND2_X1 U14551 ( .A1(n12195), .A2(n12326), .ZN(n12196) );
  XNOR2_X1 U14552 ( .A(n12653), .B(n12220), .ZN(n12198) );
  NAND2_X1 U14553 ( .A1(n12198), .A2(n12394), .ZN(n12320) );
  INV_X1 U14554 ( .A(n12198), .ZN(n12200) );
  NAND2_X1 U14555 ( .A1(n12200), .A2(n12199), .ZN(n12321) );
  XNOR2_X1 U14556 ( .A(n12709), .B(n12220), .ZN(n12364) );
  NAND2_X1 U14557 ( .A1(n12364), .A2(n12393), .ZN(n12201) );
  INV_X1 U14558 ( .A(n12364), .ZN(n12202) );
  NAND2_X1 U14559 ( .A1(n12202), .A2(n12324), .ZN(n12203) );
  NAND2_X1 U14560 ( .A1(n12204), .A2(n12203), .ZN(n12263) );
  XNOR2_X1 U14561 ( .A(n12759), .B(n12273), .ZN(n12205) );
  XNOR2_X1 U14562 ( .A(n12205), .B(n12206), .ZN(n12264) );
  NAND2_X1 U14563 ( .A1(n12263), .A2(n12264), .ZN(n12209) );
  INV_X1 U14564 ( .A(n12205), .ZN(n12207) );
  NAND2_X1 U14565 ( .A1(n12207), .A2(n12206), .ZN(n12208) );
  XNOR2_X1 U14566 ( .A(n12343), .B(n12273), .ZN(n12211) );
  XNOR2_X1 U14567 ( .A(n12211), .B(n12210), .ZN(n12344) );
  INV_X1 U14568 ( .A(n12211), .ZN(n12212) );
  NAND2_X1 U14569 ( .A1(n12212), .A2(n12391), .ZN(n12213) );
  XNOR2_X1 U14570 ( .A(n12596), .B(n12273), .ZN(n12214) );
  XNOR2_X1 U14571 ( .A(n12214), .B(n12354), .ZN(n12298) );
  NAND2_X1 U14572 ( .A1(n12214), .A2(n12354), .ZN(n12215) );
  XNOR2_X1 U14573 ( .A(n12361), .B(n12220), .ZN(n12216) );
  INV_X1 U14574 ( .A(n12216), .ZN(n12217) );
  AND2_X1 U14575 ( .A1(n12218), .A2(n12217), .ZN(n12219) );
  XNOR2_X1 U14576 ( .A(n12683), .B(n12273), .ZN(n12335) );
  XNOR2_X1 U14577 ( .A(n12687), .B(n12220), .ZN(n12332) );
  INV_X1 U14578 ( .A(n12332), .ZN(n12221) );
  OAI22_X1 U14579 ( .A1(n12335), .A2(n12569), .B1(n12355), .B2(n12221), .ZN(
        n12225) );
  OAI21_X1 U14580 ( .B1(n12332), .B2(n12388), .A(n12305), .ZN(n12223) );
  NOR2_X1 U14581 ( .A1(n12305), .A2(n12388), .ZN(n12222) );
  AOI22_X1 U14582 ( .A1(n12335), .A2(n12223), .B1(n12222), .B2(n12221), .ZN(
        n12224) );
  XNOR2_X1 U14583 ( .A(n12547), .B(n12273), .ZN(n12226) );
  XNOR2_X1 U14584 ( .A(n12226), .B(n12373), .ZN(n12304) );
  XNOR2_X1 U14585 ( .A(n12675), .B(n12273), .ZN(n12229) );
  XNOR2_X1 U14586 ( .A(n12229), .B(n12228), .ZN(n12372) );
  INV_X1 U14587 ( .A(n12229), .ZN(n12230) );
  XOR2_X1 U14588 ( .A(n12271), .B(n12272), .Z(n12235) );
  INV_X1 U14589 ( .A(n12231), .ZN(n12385) );
  AOI22_X1 U14590 ( .A1(n12385), .A2(n12375), .B1(n12374), .B2(n12387), .ZN(
        n12519) );
  AOI22_X1 U14591 ( .A1(n12525), .A2(n12376), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12232) );
  OAI21_X1 U14592 ( .B1(n12519), .B2(n12378), .A(n12232), .ZN(n12233) );
  AOI21_X1 U14593 ( .B1(n12670), .B2(n12380), .A(n12233), .ZN(n12234) );
  OAI21_X1 U14594 ( .B1(n12235), .B2(n12382), .A(n12234), .ZN(P3_U3154) );
  XNOR2_X1 U14595 ( .A(n12333), .B(n12332), .ZN(n12334) );
  XNOR2_X1 U14596 ( .A(n12334), .B(n12355), .ZN(n12242) );
  INV_X1 U14597 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n12236) );
  OAI22_X1 U14598 ( .A1(n12568), .A2(n12237), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12236), .ZN(n12240) );
  INV_X1 U14599 ( .A(n12573), .ZN(n12238) );
  OAI22_X1 U14600 ( .A1(n12569), .A2(n12278), .B1(n12238), .B2(n12358), .ZN(
        n12239) );
  AOI211_X1 U14601 ( .C1(n12687), .C2(n12380), .A(n12240), .B(n12239), .ZN(
        n12241) );
  OAI21_X1 U14602 ( .B1(n12242), .B2(n12382), .A(n12241), .ZN(P3_U3156) );
  AOI21_X1 U14603 ( .B1(n12244), .B2(n12243), .A(n12382), .ZN(n12246) );
  NAND2_X1 U14604 ( .A1(n12246), .A2(n12245), .ZN(n12254) );
  AOI22_X1 U14605 ( .A1(n12401), .A2(n12291), .B1(n12247), .B2(n12376), .ZN(
        n12253) );
  INV_X1 U14606 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n12248) );
  OAI22_X1 U14607 ( .A1(n12249), .A2(n12278), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12248), .ZN(n12250) );
  AOI21_X1 U14608 ( .B1(n12251), .B2(n12380), .A(n12250), .ZN(n12252) );
  NAND3_X1 U14609 ( .A1(n12254), .A2(n12253), .A3(n12252), .ZN(P3_U3157) );
  OAI211_X1 U14610 ( .C1(n12257), .C2(n12256), .A(n12255), .B(n12282), .ZN(
        n12262) );
  AOI22_X1 U14611 ( .A1(n12380), .A2(n12258), .B1(P3_REG3_REG_3__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12261) );
  AOI22_X1 U14612 ( .A1(n12408), .A2(n12291), .B1(n8577), .B2(n12376), .ZN(
        n12260) );
  NAND2_X1 U14613 ( .A1(n12289), .A2(n12406), .ZN(n12259) );
  NAND4_X1 U14614 ( .A1(n12262), .A2(n12261), .A3(n12260), .A4(n12259), .ZN(
        P3_U3158) );
  XOR2_X1 U14615 ( .A(n12264), .B(n12263), .Z(n12269) );
  AOI22_X1 U14616 ( .A1(n12391), .A2(n12375), .B1(n12374), .B2(n12393), .ZN(
        n12619) );
  INV_X1 U14617 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n12265) );
  OAI22_X1 U14618 ( .A1(n12619), .A2(n12378), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12265), .ZN(n12267) );
  NOR2_X1 U14619 ( .A1(n12759), .A2(n12352), .ZN(n12266) );
  AOI211_X1 U14620 ( .C1(n12622), .C2(n12376), .A(n12267), .B(n12266), .ZN(
        n12268) );
  OAI21_X1 U14621 ( .B1(n12269), .B2(n12382), .A(n12268), .ZN(P3_U3159) );
  XNOR2_X1 U14622 ( .A(n12507), .B(n12273), .ZN(n12274) );
  XNOR2_X1 U14623 ( .A(n12275), .B(n12274), .ZN(n12281) );
  AOI22_X1 U14624 ( .A1(n12509), .A2(n12376), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12277) );
  NAND2_X1 U14625 ( .A1(n12386), .A2(n12291), .ZN(n12276) );
  OAI211_X1 U14626 ( .C1(n12503), .C2(n12278), .A(n12277), .B(n12276), .ZN(
        n12279) );
  AOI21_X1 U14627 ( .B1(n12513), .B2(n12380), .A(n12279), .ZN(n12280) );
  OAI21_X1 U14628 ( .B1(n12281), .B2(n12382), .A(n12280), .ZN(P3_U3160) );
  OAI211_X1 U14629 ( .C1(n12285), .C2(n12284), .A(n12283), .B(n12282), .ZN(
        n12294) );
  OAI22_X1 U14630 ( .A1(n12352), .A2(n12287), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12286), .ZN(n12288) );
  AOI21_X1 U14631 ( .B1(n12289), .B2(n12401), .A(n12288), .ZN(n12293) );
  AOI22_X1 U14632 ( .A1(n12403), .A2(n12291), .B1(n12290), .B2(n12376), .ZN(
        n12292) );
  NAND3_X1 U14633 ( .A1(n12294), .A2(n12293), .A3(n12292), .ZN(P3_U3161) );
  INV_X1 U14634 ( .A(n12295), .ZN(n12296) );
  AOI21_X1 U14635 ( .B1(n12298), .B2(n12297), .A(n12296), .ZN(n12302) );
  AOI22_X1 U14636 ( .A1(n12389), .A2(n12375), .B1(n12391), .B2(n12374), .ZN(
        n12594) );
  OAI22_X1 U14637 ( .A1(n12594), .A2(n12378), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15313), .ZN(n12299) );
  AOI21_X1 U14638 ( .B1(n12597), .B2(n12376), .A(n12299), .ZN(n12301) );
  NAND2_X1 U14639 ( .A1(n12596), .A2(n12380), .ZN(n12300) );
  OAI211_X1 U14640 ( .C1(n12302), .C2(n12382), .A(n12301), .B(n12300), .ZN(
        P3_U3163) );
  XOR2_X1 U14641 ( .A(n12304), .B(n12303), .Z(n12309) );
  AOI22_X1 U14642 ( .A1(n12387), .A2(n12375), .B1(n12374), .B2(n12305), .ZN(
        n12545) );
  AOI22_X1 U14643 ( .A1(n12548), .A2(n12376), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12306) );
  OAI21_X1 U14644 ( .B1(n12545), .B2(n12378), .A(n12306), .ZN(n12307) );
  AOI21_X1 U14645 ( .B1(n12547), .B2(n12380), .A(n12307), .ZN(n12308) );
  OAI21_X1 U14646 ( .B1(n12309), .B2(n12382), .A(n12308), .ZN(P3_U3165) );
  XOR2_X1 U14647 ( .A(n12311), .B(n12310), .Z(n12319) );
  INV_X1 U14648 ( .A(n12312), .ZN(n12315) );
  AOI22_X1 U14649 ( .A1(n12313), .A2(n12356), .B1(P3_REG3_REG_16__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12314) );
  OAI21_X1 U14650 ( .B1(n12315), .B2(n12358), .A(n12314), .ZN(n12316) );
  AOI21_X1 U14651 ( .B1(n12317), .B2(n12380), .A(n12316), .ZN(n12318) );
  OAI21_X1 U14652 ( .B1(n12319), .B2(n12382), .A(n12318), .ZN(P3_U3166) );
  NAND2_X1 U14653 ( .A1(n12321), .A2(n12320), .ZN(n12322) );
  XNOR2_X1 U14654 ( .A(n12323), .B(n12322), .ZN(n12331) );
  INV_X1 U14655 ( .A(n12654), .ZN(n12328) );
  OR2_X1 U14656 ( .A1(n12324), .A2(n15117), .ZN(n12325) );
  OAI21_X1 U14657 ( .B1(n12326), .B2(n15119), .A(n12325), .ZN(n12650) );
  NAND2_X1 U14658 ( .A1(n12650), .A2(n12356), .ZN(n12327) );
  NAND2_X1 U14659 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n14230)
         );
  OAI211_X1 U14660 ( .C1(n12358), .C2(n12328), .A(n12327), .B(n14230), .ZN(
        n12329) );
  AOI21_X1 U14661 ( .B1(n12653), .B2(n12380), .A(n12329), .ZN(n12330) );
  OAI21_X1 U14662 ( .B1(n12331), .B2(n12382), .A(n12330), .ZN(P3_U3168) );
  OAI22_X1 U14663 ( .A1(n12334), .A2(n12388), .B1(n12333), .B2(n12332), .ZN(
        n12337) );
  XNOR2_X1 U14664 ( .A(n12335), .B(n12569), .ZN(n12336) );
  XNOR2_X1 U14665 ( .A(n12337), .B(n12336), .ZN(n12342) );
  AOI22_X1 U14666 ( .A1(n12373), .A2(n12375), .B1(n12374), .B2(n12388), .ZN(
        n12554) );
  AOI22_X1 U14667 ( .A1(n12558), .A2(n12376), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12339) );
  OAI21_X1 U14668 ( .B1(n12554), .B2(n12378), .A(n12339), .ZN(n12340) );
  AOI21_X1 U14669 ( .B1(n12683), .B2(n12380), .A(n12340), .ZN(n12341) );
  OAI21_X1 U14670 ( .B1(n12342), .B2(n12382), .A(n12341), .ZN(P3_U3169) );
  AOI21_X1 U14671 ( .B1(n12345), .B2(n12344), .A(n12382), .ZN(n12347) );
  NAND2_X1 U14672 ( .A1(n12347), .A2(n12346), .ZN(n12351) );
  AOI22_X1 U14673 ( .A1(n12390), .A2(n12375), .B1(n12374), .B2(n12392), .ZN(
        n12608) );
  OAI22_X1 U14674 ( .A1(n12608), .A2(n12378), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12348), .ZN(n12349) );
  AOI21_X1 U14675 ( .B1(n12610), .B2(n12376), .A(n12349), .ZN(n12350) );
  OAI211_X1 U14676 ( .C1(n12755), .C2(n12352), .A(n12351), .B(n12350), .ZN(
        P3_U3173) );
  XNOR2_X1 U14677 ( .A(n12353), .B(n12389), .ZN(n12363) );
  INV_X1 U14678 ( .A(n12586), .ZN(n12359) );
  OAI22_X1 U14679 ( .A1(n12355), .A2(n15117), .B1(n12354), .B2(n15119), .ZN(
        n12583) );
  AOI22_X1 U14680 ( .A1(n12583), .A2(n12356), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12357) );
  OAI21_X1 U14681 ( .B1(n12359), .B2(n12358), .A(n12357), .ZN(n12360) );
  AOI21_X1 U14682 ( .B1(n12361), .B2(n12380), .A(n12360), .ZN(n12362) );
  OAI21_X1 U14683 ( .B1(n12363), .B2(n12382), .A(n12362), .ZN(P3_U3175) );
  XNOR2_X1 U14684 ( .A(n12364), .B(n12393), .ZN(n12365) );
  XNOR2_X1 U14685 ( .A(n12366), .B(n12365), .ZN(n12370) );
  AOI22_X1 U14686 ( .A1(n12394), .A2(n12374), .B1(n12375), .B2(n12392), .ZN(
        n12634) );
  NAND2_X1 U14687 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n14242)
         );
  NAND2_X1 U14688 ( .A1(n12376), .A2(n12636), .ZN(n12367) );
  OAI211_X1 U14689 ( .C1(n12634), .C2(n12378), .A(n14242), .B(n12367), .ZN(
        n12368) );
  AOI21_X1 U14690 ( .B1(n12709), .B2(n12380), .A(n12368), .ZN(n12369) );
  OAI21_X1 U14691 ( .B1(n12370), .B2(n12382), .A(n12369), .ZN(P3_U3178) );
  XOR2_X1 U14692 ( .A(n12372), .B(n12371), .Z(n12383) );
  AOI22_X1 U14693 ( .A1(n12386), .A2(n12375), .B1(n12374), .B2(n12373), .ZN(
        n12537) );
  AOI22_X1 U14694 ( .A1(n12531), .A2(n12376), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12377) );
  OAI21_X1 U14695 ( .B1(n12537), .B2(n12378), .A(n12377), .ZN(n12379) );
  AOI21_X1 U14696 ( .B1(n12675), .B2(n12380), .A(n12379), .ZN(n12381) );
  OAI21_X1 U14697 ( .B1(n12383), .B2(n12382), .A(n12381), .ZN(P3_U3180) );
  MUX2_X1 U14698 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12384), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U14699 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12385), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14700 ( .A(n12386), .B(P3_DATAO_REG_27__SCAN_IN), .S(n12410), .Z(
        P3_U3518) );
  MUX2_X1 U14701 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n12387), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U14702 ( .A(n12388), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12410), .Z(
        P3_U3514) );
  MUX2_X1 U14703 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12389), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U14704 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12390), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14705 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12391), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14706 ( .A(n12392), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12410), .Z(
        P3_U3510) );
  MUX2_X1 U14707 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12393), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14708 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n12394), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14709 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n12395), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14710 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n12396), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U14711 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n12397), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U14712 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12398), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14713 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n12399), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U14714 ( .A(n12400), .B(P3_DATAO_REG_10__SCAN_IN), .S(n12410), .Z(
        P3_U3501) );
  MUX2_X1 U14715 ( .A(n12401), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12410), .Z(
        P3_U3500) );
  MUX2_X1 U14716 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12402), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U14717 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12403), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14718 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12404), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14719 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12405), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U14720 ( .A(n12406), .B(P3_DATAO_REG_4__SCAN_IN), .S(n12410), .Z(
        P3_U3495) );
  MUX2_X1 U14721 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n12407), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U14722 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n12408), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U14723 ( .A(n12409), .B(P3_DATAO_REG_1__SCAN_IN), .S(n12410), .Z(
        P3_U3492) );
  MUX2_X1 U14724 ( .A(n12411), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12410), .Z(
        P3_U3491) );
  NOR2_X1 U14725 ( .A1(n12460), .A2(n12412), .ZN(n12414) );
  AOI22_X1 U14726 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n12462), .B1(n15033), 
        .B2(n12429), .ZN(n15024) );
  NOR2_X1 U14727 ( .A1(n12464), .A2(n12415), .ZN(n12416) );
  INV_X1 U14728 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n15329) );
  NOR2_X1 U14729 ( .A1(n12416), .A2(n15038), .ZN(n15057) );
  INV_X1 U14730 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12417) );
  MUX2_X1 U14731 ( .A(P3_REG2_REG_12__SCAN_IN), .B(n12417), .S(n12466), .Z(
        n15056) );
  NAND2_X1 U14732 ( .A1(n15063), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n12418) );
  INV_X1 U14733 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n15557) );
  NAND2_X1 U14734 ( .A1(n15100), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12442) );
  OAI21_X1 U14735 ( .B1(n15100), .B2(P3_REG2_REG_14__SCAN_IN), .A(n12442), 
        .ZN(n15090) );
  NOR2_X1 U14736 ( .A1(n15091), .A2(n15090), .ZN(n15089) );
  INV_X1 U14737 ( .A(n12442), .ZN(n12420) );
  INV_X1 U14738 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n14192) );
  NAND2_X1 U14739 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n14214), .ZN(n12422) );
  OAI21_X1 U14740 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(n14214), .A(n12422), 
        .ZN(n14209) );
  NOR2_X1 U14741 ( .A1(n12478), .A2(n12423), .ZN(n12424) );
  INV_X1 U14742 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n14225) );
  NAND2_X1 U14743 ( .A1(P3_REG2_REG_18__SCAN_IN), .A2(n14243), .ZN(n12425) );
  OAI21_X1 U14744 ( .B1(P3_REG2_REG_18__SCAN_IN), .B2(n14243), .A(n12425), 
        .ZN(n14241) );
  AOI21_X1 U14745 ( .B1(P3_REG2_REG_18__SCAN_IN), .B2(n14243), .A(n14240), 
        .ZN(n12426) );
  XNOR2_X1 U14746 ( .A(n12483), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12453) );
  XNOR2_X1 U14747 ( .A(n12426), .B(n12453), .ZN(n12484) );
  MUX2_X1 U14748 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12452), .Z(n14248) );
  MUX2_X1 U14749 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12452), .Z(n12448) );
  INV_X1 U14750 ( .A(n12478), .ZN(n14231) );
  NAND2_X1 U14751 ( .A1(n12448), .A2(n14231), .ZN(n12449) );
  MUX2_X1 U14752 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12452), .Z(n12427) );
  INV_X1 U14753 ( .A(n12427), .ZN(n12440) );
  XOR2_X1 U14754 ( .A(n15074), .B(n12427), .Z(n15081) );
  MUX2_X1 U14755 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12452), .Z(n12438) );
  NAND2_X1 U14756 ( .A1(n12438), .A2(n15063), .ZN(n12439) );
  MUX2_X1 U14757 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12452), .Z(n12436) );
  INV_X1 U14758 ( .A(n12436), .ZN(n12437) );
  INV_X1 U14759 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n12428) );
  MUX2_X1 U14760 ( .A(n12429), .B(n12428), .S(n12452), .Z(n12434) );
  AND2_X1 U14761 ( .A1(n12434), .A2(n12462), .ZN(n12435) );
  INV_X1 U14762 ( .A(n12435), .ZN(n12433) );
  OAI21_X1 U14763 ( .B1(n12462), .B2(n12434), .A(n12433), .ZN(n15028) );
  NOR2_X1 U14764 ( .A1(n15027), .A2(n15028), .ZN(n15026) );
  NOR2_X1 U14765 ( .A1(n12435), .A2(n15026), .ZN(n15046) );
  XNOR2_X1 U14766 ( .A(n12436), .B(n15041), .ZN(n15047) );
  NOR2_X1 U14767 ( .A1(n15046), .A2(n15047), .ZN(n15045) );
  XNOR2_X1 U14768 ( .A(n12438), .B(n12466), .ZN(n15067) );
  NAND2_X1 U14769 ( .A1(n15068), .A2(n15067), .ZN(n15066) );
  NAND2_X1 U14770 ( .A1(n12439), .A2(n15066), .ZN(n15080) );
  NOR2_X1 U14771 ( .A1(n15081), .A2(n15080), .ZN(n15079) );
  INV_X1 U14772 ( .A(n15090), .ZN(n12441) );
  NAND2_X1 U14773 ( .A1(n15100), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12472) );
  OAI21_X1 U14774 ( .B1(n15100), .B2(P3_REG1_REG_14__SCAN_IN), .A(n12472), 
        .ZN(n15093) );
  MUX2_X1 U14775 ( .A(n12441), .B(n12471), .S(n12452), .Z(n15106) );
  NAND2_X1 U14776 ( .A1(n15107), .A2(n15106), .ZN(n15105) );
  MUX2_X1 U14777 ( .A(n12442), .B(n12472), .S(n12452), .Z(n12443) );
  NAND2_X1 U14778 ( .A1(n15105), .A2(n12443), .ZN(n12444) );
  XNOR2_X1 U14779 ( .A(n12444), .B(n14198), .ZN(n14203) );
  MUX2_X1 U14780 ( .A(n14192), .B(n14194), .S(n12452), .Z(n14202) );
  MUX2_X1 U14781 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n12452), .Z(n12445) );
  XNOR2_X1 U14782 ( .A(n12445), .B(n14214), .ZN(n14218) );
  INV_X1 U14783 ( .A(n12445), .ZN(n12446) );
  XNOR2_X1 U14784 ( .A(n12448), .B(n12478), .ZN(n14235) );
  NAND2_X1 U14785 ( .A1(n14236), .A2(n14235), .ZN(n14234) );
  NAND2_X1 U14786 ( .A1(n12449), .A2(n14234), .ZN(n12450) );
  XNOR2_X1 U14787 ( .A(n14243), .B(n12450), .ZN(n14249) );
  NOR2_X1 U14788 ( .A1(n14248), .A2(n14249), .ZN(n14247) );
  NOR2_X1 U14789 ( .A1(n14243), .A2(n12450), .ZN(n12451) );
  XNOR2_X1 U14790 ( .A(n12483), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12481) );
  MUX2_X1 U14791 ( .A(n12453), .B(n12481), .S(n12452), .Z(n12454) );
  XNOR2_X1 U14792 ( .A(n12455), .B(n12454), .ZN(n12458) );
  NAND2_X1 U14793 ( .A1(P3_REG3_REG_19__SCAN_IN), .A2(P3_U3151), .ZN(n12457)
         );
  NAND2_X1 U14794 ( .A1(n15025), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12456) );
  OAI211_X1 U14795 ( .C1(n12458), .C2(n15082), .A(n12457), .B(n12456), .ZN(
        n12482) );
  INV_X1 U14796 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n14227) );
  INV_X1 U14797 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n15078) );
  INV_X1 U14798 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n15044) );
  AOI22_X1 U14799 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n12462), .B1(n15033), 
        .B2(n12428), .ZN(n15030) );
  NOR2_X1 U14800 ( .A1(n12464), .A2(n12463), .ZN(n12465) );
  INV_X1 U14801 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n12467) );
  MUX2_X1 U14802 ( .A(P3_REG1_REG_12__SCAN_IN), .B(n12467), .S(n12466), .Z(
        n15058) );
  NAND2_X1 U14803 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n14214), .ZN(n12475) );
  OAI21_X1 U14804 ( .B1(P3_REG1_REG_16__SCAN_IN), .B2(n14214), .A(n12475), 
        .ZN(n14211) );
  XNOR2_X1 U14805 ( .A(n12477), .B(n12478), .ZN(n14228) );
  NOR2_X1 U14806 ( .A1(n12478), .A2(n12477), .ZN(n12479) );
  INV_X1 U14807 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12712) );
  AOI22_X1 U14808 ( .A1(P3_REG1_REG_18__SCAN_IN), .A2(n12480), .B1(n14243), 
        .B2(n12712), .ZN(n14245) );
  INV_X1 U14809 ( .A(n12722), .ZN(n12662) );
  NOR2_X1 U14810 ( .A1(n12486), .A2(n12485), .ZN(n12723) );
  NOR2_X1 U14811 ( .A1(n12487), .A2(n14270), .ZN(n12492) );
  AOI21_X1 U14812 ( .B1(n12723), .B2(n15131), .A(n12492), .ZN(n12490) );
  NAND2_X1 U14813 ( .A1(n15595), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12488) );
  OAI211_X1 U14814 ( .C1(n12662), .C2(n15593), .A(n12490), .B(n12488), .ZN(
        P3_U3202) );
  NAND2_X1 U14815 ( .A1(n15595), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n12489) );
  OAI211_X1 U14816 ( .C1(n12665), .C2(n15593), .A(n12490), .B(n12489), .ZN(
        P3_U3203) );
  INV_X1 U14817 ( .A(n12491), .ZN(n12498) );
  AOI21_X1 U14818 ( .B1(n15595), .B2(P3_REG2_REG_29__SCAN_IN), .A(n12492), 
        .ZN(n12493) );
  OAI21_X1 U14819 ( .B1(n12494), .B2(n15593), .A(n12493), .ZN(n12495) );
  AOI21_X1 U14820 ( .B1(n12496), .B2(n15600), .A(n12495), .ZN(n12497) );
  OAI21_X1 U14821 ( .B1(n12498), .B2(n15595), .A(n12497), .ZN(P3_U3204) );
  OAI211_X1 U14822 ( .C1(n12501), .C2(n12500), .A(n12499), .B(n15122), .ZN(
        n12506) );
  OAI22_X1 U14823 ( .A1(n12503), .A2(n15117), .B1(n12502), .B2(n15119), .ZN(
        n12504) );
  INV_X1 U14824 ( .A(n12504), .ZN(n12505) );
  XNOR2_X1 U14825 ( .A(n12508), .B(n12507), .ZN(n12666) );
  NAND2_X1 U14826 ( .A1(n12666), .A2(n15600), .ZN(n12515) );
  INV_X1 U14827 ( .A(n12509), .ZN(n12511) );
  INV_X1 U14828 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n12510) );
  OAI22_X1 U14829 ( .A1(n12511), .A2(n14270), .B1(n15131), .B2(n12510), .ZN(
        n12512) );
  AOI21_X1 U14830 ( .B1(n12513), .B2(n12640), .A(n12512), .ZN(n12514) );
  OAI211_X1 U14831 ( .C1(n12667), .C2(n15595), .A(n12515), .B(n12514), .ZN(
        P3_U3205) );
  OAI21_X1 U14832 ( .B1(n12518), .B2(n12517), .A(n12516), .ZN(n12521) );
  INV_X1 U14833 ( .A(n12519), .ZN(n12520) );
  AOI21_X1 U14834 ( .B1(n12521), .B2(n15122), .A(n12520), .ZN(n12672) );
  OAI21_X1 U14835 ( .B1(n12524), .B2(n12523), .A(n12522), .ZN(n12671) );
  INV_X1 U14836 ( .A(n12670), .ZN(n12527) );
  AOI22_X1 U14837 ( .A1(n12525), .A2(n15591), .B1(n15595), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12526) );
  OAI21_X1 U14838 ( .B1(n12527), .B2(n15593), .A(n12526), .ZN(n12528) );
  AOI21_X1 U14839 ( .B1(n12671), .B2(n15600), .A(n12528), .ZN(n12529) );
  OAI21_X1 U14840 ( .B1(n15595), .B2(n12672), .A(n12529), .ZN(P3_U3206) );
  XOR2_X1 U14841 ( .A(n12535), .B(n12530), .Z(n12678) );
  INV_X1 U14842 ( .A(n12531), .ZN(n12533) );
  INV_X1 U14843 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n12532) );
  OAI22_X1 U14844 ( .A1(n12533), .A2(n14270), .B1(n15131), .B2(n12532), .ZN(
        n12534) );
  AOI21_X1 U14845 ( .B1(n12675), .B2(n12640), .A(n12534), .ZN(n12540) );
  XNOR2_X1 U14846 ( .A(n12536), .B(n12535), .ZN(n12538) );
  OAI21_X1 U14847 ( .B1(n12538), .B2(n14264), .A(n12537), .ZN(n12674) );
  NAND2_X1 U14848 ( .A1(n12674), .A2(n12657), .ZN(n12539) );
  OAI211_X1 U14849 ( .C1(n12678), .C2(n12659), .A(n12540), .B(n12539), .ZN(
        P3_U3207) );
  XOR2_X1 U14850 ( .A(n12542), .B(n12541), .Z(n12546) );
  OAI211_X1 U14851 ( .C1(n6730), .C2(n7601), .A(n15122), .B(n12543), .ZN(
        n12544) );
  OAI211_X1 U14852 ( .C1(n12546), .C2(n15125), .A(n12545), .B(n12544), .ZN(
        n12679) );
  INV_X1 U14853 ( .A(n12679), .ZN(n12552) );
  INV_X1 U14854 ( .A(n12546), .ZN(n12680) );
  INV_X1 U14855 ( .A(n12547), .ZN(n12738) );
  AOI22_X1 U14856 ( .A1(n12548), .A2(n15591), .B1(n15595), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n12549) );
  OAI21_X1 U14857 ( .B1(n12738), .B2(n15593), .A(n12549), .ZN(n12550) );
  AOI21_X1 U14858 ( .B1(n12680), .B2(n15128), .A(n12550), .ZN(n12551) );
  OAI21_X1 U14859 ( .B1(n12552), .B2(n15595), .A(n12551), .ZN(P3_U3208) );
  XNOR2_X1 U14860 ( .A(n12553), .B(n7374), .ZN(n12556) );
  INV_X1 U14861 ( .A(n12554), .ZN(n12555) );
  AOI21_X1 U14862 ( .B1(n12556), .B2(n15122), .A(n12555), .ZN(n12685) );
  OAI21_X1 U14863 ( .B1(n6709), .B2(n7374), .A(n12557), .ZN(n12684) );
  INV_X1 U14864 ( .A(n12683), .ZN(n12560) );
  AOI22_X1 U14865 ( .A1(n12558), .A2(n15591), .B1(n15595), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n12559) );
  OAI21_X1 U14866 ( .B1(n12560), .B2(n15593), .A(n12559), .ZN(n12561) );
  AOI21_X1 U14867 ( .B1(n12684), .B2(n15600), .A(n12561), .ZN(n12562) );
  OAI21_X1 U14868 ( .B1(n15595), .B2(n12685), .A(n12562), .ZN(P3_U3209) );
  OR2_X1 U14869 ( .A1(n12563), .A2(n12567), .ZN(n12564) );
  NAND2_X1 U14870 ( .A1(n12565), .A2(n12564), .ZN(n12688) );
  XNOR2_X1 U14871 ( .A(n12566), .B(n12567), .ZN(n12571) );
  OAI22_X1 U14872 ( .A1(n12569), .A2(n15117), .B1(n12568), .B2(n15119), .ZN(
        n12570) );
  AOI21_X1 U14873 ( .B1(n12571), .B2(n15122), .A(n12570), .ZN(n12572) );
  OAI21_X1 U14874 ( .B1(n12688), .B2(n15125), .A(n12572), .ZN(n12689) );
  AOI22_X1 U14875 ( .A1(n12573), .A2(n15591), .B1(n15595), .B2(
        P3_REG2_REG_23__SCAN_IN), .ZN(n12575) );
  NAND2_X1 U14876 ( .A1(n12687), .A2(n12640), .ZN(n12574) );
  OAI211_X1 U14877 ( .C1(n12688), .C2(n12576), .A(n12575), .B(n12574), .ZN(
        n12577) );
  AOI21_X1 U14878 ( .B1(n12689), .B2(n12657), .A(n12577), .ZN(n12578) );
  INV_X1 U14879 ( .A(n12578), .ZN(P3_U3210) );
  XNOR2_X1 U14880 ( .A(n12580), .B(n12579), .ZN(n12694) );
  INV_X1 U14881 ( .A(n12694), .ZN(n12590) );
  XNOR2_X1 U14882 ( .A(n12582), .B(n12581), .ZN(n12585) );
  INV_X1 U14883 ( .A(n12583), .ZN(n12584) );
  OAI21_X1 U14884 ( .B1(n12585), .B2(n14264), .A(n12584), .ZN(n12693) );
  AOI22_X1 U14885 ( .A1(n15595), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n12586), 
        .B2(n15591), .ZN(n12587) );
  OAI21_X1 U14886 ( .B1(n12747), .B2(n15593), .A(n12587), .ZN(n12588) );
  AOI21_X1 U14887 ( .B1(n12693), .B2(n12657), .A(n12588), .ZN(n12589) );
  OAI21_X1 U14888 ( .B1(n12590), .B2(n12659), .A(n12589), .ZN(P3_U3211) );
  XOR2_X1 U14889 ( .A(n12593), .B(n12591), .Z(n12698) );
  INV_X1 U14890 ( .A(n12698), .ZN(n12601) );
  AOI21_X1 U14891 ( .B1(n12593), .B2(n12592), .A(n6715), .ZN(n12595) );
  OAI21_X1 U14892 ( .B1(n12595), .B2(n14264), .A(n12594), .ZN(n12697) );
  INV_X1 U14893 ( .A(n12596), .ZN(n12751) );
  AOI22_X1 U14894 ( .A1(n15595), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n15591), 
        .B2(n12597), .ZN(n12598) );
  OAI21_X1 U14895 ( .B1(n12751), .B2(n15593), .A(n12598), .ZN(n12599) );
  AOI21_X1 U14896 ( .B1(n12697), .B2(n12657), .A(n12599), .ZN(n12600) );
  OAI21_X1 U14897 ( .B1(n12601), .B2(n12659), .A(n12600), .ZN(P3_U3212) );
  AOI21_X1 U14898 ( .B1(n12604), .B2(n12602), .A(n6781), .ZN(n12702) );
  INV_X1 U14899 ( .A(n12702), .ZN(n12614) );
  NAND3_X1 U14900 ( .A1(n12616), .A2(n7109), .A3(n12605), .ZN(n12606) );
  NAND3_X1 U14901 ( .A1(n12607), .A2(n15122), .A3(n12606), .ZN(n12609) );
  NAND2_X1 U14902 ( .A1(n12609), .A2(n12608), .ZN(n12701) );
  AOI22_X1 U14903 ( .A1(n15595), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n15591), 
        .B2(n12610), .ZN(n12611) );
  OAI21_X1 U14904 ( .B1(n12755), .B2(n15593), .A(n12611), .ZN(n12612) );
  AOI21_X1 U14905 ( .B1(n12701), .B2(n12657), .A(n12612), .ZN(n12613) );
  OAI21_X1 U14906 ( .B1(n12614), .B2(n12659), .A(n12613), .ZN(P3_U3213) );
  XNOR2_X1 U14907 ( .A(n12615), .B(n12617), .ZN(n12706) );
  INV_X1 U14908 ( .A(n12706), .ZN(n12626) );
  NAND2_X1 U14909 ( .A1(n12616), .A2(n15122), .ZN(n12621) );
  AOI21_X1 U14910 ( .B1(n12630), .B2(n12618), .A(n12617), .ZN(n12620) );
  OAI21_X1 U14911 ( .B1(n12621), .B2(n12620), .A(n12619), .ZN(n12705) );
  AOI22_X1 U14912 ( .A1(n15595), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n15591), 
        .B2(n12622), .ZN(n12623) );
  OAI21_X1 U14913 ( .B1(n12759), .B2(n15593), .A(n12623), .ZN(n12624) );
  AOI21_X1 U14914 ( .B1(n12705), .B2(n12657), .A(n12624), .ZN(n12625) );
  OAI21_X1 U14915 ( .B1(n12626), .B2(n12659), .A(n12625), .ZN(P3_U3214) );
  NAND2_X1 U14916 ( .A1(n12627), .A2(n8819), .ZN(n12628) );
  INV_X1 U14917 ( .A(n12711), .ZN(n12643) );
  INV_X1 U14918 ( .A(n12630), .ZN(n12631) );
  AOI21_X1 U14919 ( .B1(n12633), .B2(n12632), .A(n12631), .ZN(n12635) );
  OAI21_X1 U14920 ( .B1(n12635), .B2(n14264), .A(n12634), .ZN(n12710) );
  NAND2_X1 U14921 ( .A1(n12710), .A2(n12657), .ZN(n12642) );
  INV_X1 U14922 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12638) );
  INV_X1 U14923 ( .A(n12636), .ZN(n12637) );
  OAI22_X1 U14924 ( .A1(n12657), .A2(n12638), .B1(n12637), .B2(n14270), .ZN(
        n12639) );
  AOI21_X1 U14925 ( .B1(n12709), .B2(n12640), .A(n12639), .ZN(n12641) );
  OAI211_X1 U14926 ( .C1(n12659), .C2(n12643), .A(n12642), .B(n12641), .ZN(
        P3_U3215) );
  OAI21_X1 U14927 ( .B1(n12645), .B2(n12647), .A(n12644), .ZN(n12715) );
  INV_X1 U14928 ( .A(n12715), .ZN(n12660) );
  NAND3_X1 U14929 ( .A1(n11505), .A2(n12647), .A3(n12646), .ZN(n12648) );
  NAND3_X1 U14930 ( .A1(n12649), .A2(n15122), .A3(n12648), .ZN(n12652) );
  INV_X1 U14931 ( .A(n12650), .ZN(n12651) );
  NAND2_X1 U14932 ( .A1(n12652), .A2(n12651), .ZN(n12714) );
  INV_X1 U14933 ( .A(n12653), .ZN(n12767) );
  AOI22_X1 U14934 ( .A1(n15595), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n12654), 
        .B2(n15591), .ZN(n12655) );
  OAI21_X1 U14935 ( .B1(n12767), .B2(n15593), .A(n12655), .ZN(n12656) );
  AOI21_X1 U14936 ( .B1(n12714), .B2(n12657), .A(n12656), .ZN(n12658) );
  OAI21_X1 U14937 ( .B1(n12660), .B2(n12659), .A(n12658), .ZN(P3_U3216) );
  NAND2_X1 U14938 ( .A1(n12723), .A2(n15202), .ZN(n12663) );
  NAND2_X1 U14939 ( .A1(n8976), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12661) );
  OAI211_X1 U14940 ( .C1(n12662), .C2(n12721), .A(n12663), .B(n12661), .ZN(
        P3_U3490) );
  NAND2_X1 U14941 ( .A1(n8976), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n12664) );
  OAI211_X1 U14942 ( .C1(n12665), .C2(n12721), .A(n12664), .B(n12663), .ZN(
        P3_U3489) );
  NAND2_X1 U14943 ( .A1(n12666), .A2(n14289), .ZN(n12668) );
  AOI22_X1 U14944 ( .A1(n12671), .A2(n14289), .B1(n15157), .B2(n12670), .ZN(
        n12673) );
  NAND2_X1 U14945 ( .A1(n12673), .A2(n12672), .ZN(n12733) );
  MUX2_X1 U14946 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n12733), .S(n15202), .Z(
        P3_U3486) );
  INV_X1 U14947 ( .A(n14289), .ZN(n12677) );
  AOI21_X1 U14948 ( .B1(n15157), .B2(n12675), .A(n12674), .ZN(n12676) );
  OAI21_X1 U14949 ( .B1(n12678), .B2(n12677), .A(n12676), .ZN(n12734) );
  MUX2_X1 U14950 ( .A(P3_REG1_REG_26__SCAN_IN), .B(n12734), .S(n15202), .Z(
        P3_U3485) );
  AOI21_X1 U14951 ( .B1(n15179), .B2(n12680), .A(n12679), .ZN(n12735) );
  MUX2_X1 U14952 ( .A(n12681), .B(n12735), .S(n15202), .Z(n12682) );
  OAI21_X1 U14953 ( .B1(n12738), .B2(n12721), .A(n12682), .ZN(P3_U3484) );
  AOI22_X1 U14954 ( .A1(n12684), .A2(n14289), .B1(n15157), .B2(n12683), .ZN(
        n12686) );
  NAND2_X1 U14955 ( .A1(n12686), .A2(n12685), .ZN(n12739) );
  MUX2_X1 U14956 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n12739), .S(n15202), .Z(
        P3_U3483) );
  INV_X1 U14957 ( .A(n12687), .ZN(n12743) );
  INV_X1 U14958 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n12691) );
  INV_X1 U14959 ( .A(n12688), .ZN(n12690) );
  AOI21_X1 U14960 ( .B1(n15179), .B2(n12690), .A(n12689), .ZN(n12740) );
  MUX2_X1 U14961 ( .A(n12691), .B(n12740), .S(n15202), .Z(n12692) );
  OAI21_X1 U14962 ( .B1(n12743), .B2(n12721), .A(n12692), .ZN(P3_U3482) );
  INV_X1 U14963 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12695) );
  AOI21_X1 U14964 ( .B1(n14289), .B2(n12694), .A(n12693), .ZN(n12744) );
  MUX2_X1 U14965 ( .A(n12695), .B(n12744), .S(n15202), .Z(n12696) );
  OAI21_X1 U14966 ( .B1(n12747), .B2(n12721), .A(n12696), .ZN(P3_U3481) );
  INV_X1 U14967 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12699) );
  AOI21_X1 U14968 ( .B1(n14289), .B2(n12698), .A(n12697), .ZN(n12748) );
  MUX2_X1 U14969 ( .A(n12699), .B(n12748), .S(n15202), .Z(n12700) );
  OAI21_X1 U14970 ( .B1(n12751), .B2(n12721), .A(n12700), .ZN(P3_U3480) );
  INV_X1 U14971 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n12703) );
  AOI21_X1 U14972 ( .B1(n12702), .B2(n14289), .A(n12701), .ZN(n12752) );
  MUX2_X1 U14973 ( .A(n12703), .B(n12752), .S(n15202), .Z(n12704) );
  OAI21_X1 U14974 ( .B1(n12755), .B2(n12721), .A(n12704), .ZN(P3_U3479) );
  INV_X1 U14975 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12707) );
  AOI21_X1 U14976 ( .B1(n14289), .B2(n12706), .A(n12705), .ZN(n12756) );
  MUX2_X1 U14977 ( .A(n12707), .B(n12756), .S(n15202), .Z(n12708) );
  OAI21_X1 U14978 ( .B1(n12721), .B2(n12759), .A(n12708), .ZN(P3_U3478) );
  INV_X1 U14979 ( .A(n12709), .ZN(n12763) );
  AOI21_X1 U14980 ( .B1(n12711), .B2(n14289), .A(n12710), .ZN(n12760) );
  MUX2_X1 U14981 ( .A(n12712), .B(n12760), .S(n15202), .Z(n12713) );
  OAI21_X1 U14982 ( .B1(n12763), .B2(n12721), .A(n12713), .ZN(P3_U3477) );
  AOI21_X1 U14983 ( .B1(n12715), .B2(n14289), .A(n12714), .ZN(n12764) );
  MUX2_X1 U14984 ( .A(n14227), .B(n12764), .S(n15202), .Z(n12716) );
  OAI21_X1 U14985 ( .B1(n12767), .B2(n12721), .A(n12716), .ZN(P3_U3476) );
  INV_X1 U14986 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12719) );
  AOI21_X1 U14987 ( .B1(n14289), .B2(n12718), .A(n12717), .ZN(n12768) );
  MUX2_X1 U14988 ( .A(n12719), .B(n12768), .S(n15202), .Z(n12720) );
  OAI21_X1 U14989 ( .B1(n12772), .B2(n12721), .A(n12720), .ZN(P3_U3475) );
  INV_X1 U14990 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n12725) );
  NAND2_X1 U14991 ( .A1(n12722), .A2(n9586), .ZN(n12724) );
  NAND2_X1 U14992 ( .A1(n12723), .A2(n15181), .ZN(n12727) );
  OAI211_X1 U14993 ( .C1(n12725), .C2(n15181), .A(n12724), .B(n12727), .ZN(
        P3_U3458) );
  INV_X1 U14994 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n12729) );
  NAND2_X1 U14995 ( .A1(n12726), .A2(n9586), .ZN(n12728) );
  OAI211_X1 U14996 ( .C1(n12729), .C2(n15181), .A(n12728), .B(n12727), .ZN(
        P3_U3457) );
  INV_X1 U14997 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n12731) );
  MUX2_X1 U14998 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n12733), .S(n15181), .Z(
        P3_U3454) );
  MUX2_X1 U14999 ( .A(P3_REG0_REG_26__SCAN_IN), .B(n12734), .S(n15181), .Z(
        P3_U3453) );
  INV_X1 U15000 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n12736) );
  MUX2_X1 U15001 ( .A(n12736), .B(n12735), .S(n15181), .Z(n12737) );
  OAI21_X1 U15002 ( .B1(n12738), .B2(n12771), .A(n12737), .ZN(P3_U3452) );
  MUX2_X1 U15003 ( .A(P3_REG0_REG_24__SCAN_IN), .B(n12739), .S(n15181), .Z(
        P3_U3451) );
  INV_X1 U15004 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n12741) );
  MUX2_X1 U15005 ( .A(n12741), .B(n12740), .S(n15181), .Z(n12742) );
  OAI21_X1 U15006 ( .B1(n12743), .B2(n12771), .A(n12742), .ZN(P3_U3450) );
  INV_X1 U15007 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n12745) );
  MUX2_X1 U15008 ( .A(n12745), .B(n12744), .S(n15181), .Z(n12746) );
  OAI21_X1 U15009 ( .B1(n12747), .B2(n12771), .A(n12746), .ZN(P3_U3449) );
  INV_X1 U15010 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12749) );
  MUX2_X1 U15011 ( .A(n12749), .B(n12748), .S(n15181), .Z(n12750) );
  OAI21_X1 U15012 ( .B1(n12751), .B2(n12771), .A(n12750), .ZN(P3_U3448) );
  INV_X1 U15013 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n12753) );
  MUX2_X1 U15014 ( .A(n12753), .B(n12752), .S(n15181), .Z(n12754) );
  OAI21_X1 U15015 ( .B1(n12755), .B2(n12771), .A(n12754), .ZN(P3_U3447) );
  INV_X1 U15016 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n12757) );
  MUX2_X1 U15017 ( .A(n12757), .B(n12756), .S(n15181), .Z(n12758) );
  OAI21_X1 U15018 ( .B1(n12771), .B2(n12759), .A(n12758), .ZN(P3_U3446) );
  INV_X1 U15019 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n12761) );
  MUX2_X1 U15020 ( .A(n12761), .B(n12760), .S(n15181), .Z(n12762) );
  OAI21_X1 U15021 ( .B1(n12763), .B2(n12771), .A(n12762), .ZN(P3_U3444) );
  INV_X1 U15022 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n12765) );
  MUX2_X1 U15023 ( .A(n12765), .B(n12764), .S(n15181), .Z(n12766) );
  OAI21_X1 U15024 ( .B1(n12767), .B2(n12771), .A(n12766), .ZN(P3_U3441) );
  INV_X1 U15025 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n12769) );
  MUX2_X1 U15026 ( .A(n12769), .B(n12768), .S(n15181), .Z(n12770) );
  OAI21_X1 U15027 ( .B1(n12772), .B2(n12771), .A(n12770), .ZN(P3_U3438) );
  MUX2_X1 U15028 ( .A(n12774), .B(P3_D_REG_0__SCAN_IN), .S(n12773), .Z(
        P3_U3376) );
  NAND2_X1 U15029 ( .A1(n12776), .A2(n12775), .ZN(n12780) );
  NAND4_X1 U15030 ( .A1(n8536), .A2(P3_STATE_REG_SCAN_IN), .A3(
        P3_IR_REG_31__SCAN_IN), .A4(n12778), .ZN(n12779) );
  OAI211_X1 U15031 ( .C1(n12781), .C2(n12787), .A(n12780), .B(n12779), .ZN(
        P3_U3264) );
  INV_X1 U15032 ( .A(n12782), .ZN(n12784) );
  OAI222_X1 U15033 ( .A1(n12787), .A2(n12786), .B1(n12785), .B2(n12784), .C1(
        P3_U3151), .C2(n12783), .ZN(P3_U3266) );
  MUX2_X1 U15034 ( .A(n12788), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  AOI21_X1 U15035 ( .B1(n12790), .B2(n12789), .A(n12908), .ZN(n12792) );
  NAND2_X1 U15036 ( .A1(n12792), .A2(n12791), .ZN(n12797) );
  OAI22_X1 U15037 ( .A1(n12793), .A2(n12891), .B1(n12828), .B2(n12889), .ZN(
        n13016) );
  OAI22_X1 U15038 ( .A1(n13023), .A2(n12894), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12794), .ZN(n12795) );
  AOI21_X1 U15039 ( .B1(n13016), .B2(n12897), .A(n12795), .ZN(n12796) );
  OAI211_X1 U15040 ( .C1(n13019), .C2(n12900), .A(n12797), .B(n12796), .ZN(
        P2_U3186) );
  INV_X1 U15041 ( .A(n13257), .ZN(n13083) );
  OAI211_X1 U15042 ( .C1(n12800), .C2(n12799), .A(n12798), .B(n12887), .ZN(
        n12805) );
  OAI22_X1 U15043 ( .A1(n12827), .A2(n12891), .B1(n12801), .B2(n12889), .ZN(
        n13076) );
  OAI22_X1 U15044 ( .A1(n13078), .A2(n12894), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12802), .ZN(n12803) );
  AOI21_X1 U15045 ( .B1(n13076), .B2(n12897), .A(n12803), .ZN(n12804) );
  OAI211_X1 U15046 ( .C1(n13083), .C2(n12900), .A(n12805), .B(n12804), .ZN(
        P2_U3188) );
  NOR2_X1 U15047 ( .A1(n12806), .A2(n6772), .ZN(n12807) );
  XNOR2_X1 U15048 ( .A(n12808), .B(n12807), .ZN(n12814) );
  OAI22_X1 U15049 ( .A1(n12810), .A2(n12891), .B1(n12809), .B2(n12889), .ZN(
        n13134) );
  NAND2_X1 U15050 ( .A1(n13134), .A2(n12897), .ZN(n12811) );
  NAND2_X1 U15051 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n12986)
         );
  OAI211_X1 U15052 ( .C1(n12894), .C2(n13140), .A(n12811), .B(n12986), .ZN(
        n12812) );
  AOI21_X1 U15053 ( .B1(n13278), .B2(n12913), .A(n12812), .ZN(n12813) );
  OAI21_X1 U15054 ( .B1(n12814), .B2(n12908), .A(n12813), .ZN(P2_U3191) );
  OAI211_X1 U15055 ( .C1(n12817), .C2(n12816), .A(n12815), .B(n12887), .ZN(
        n12823) );
  NAND2_X1 U15056 ( .A1(n12923), .A2(n12902), .ZN(n12819) );
  NAND2_X1 U15057 ( .A1(n12925), .A2(n12901), .ZN(n12818) );
  NAND2_X1 U15058 ( .A1(n12819), .A2(n12818), .ZN(n13105) );
  OAI22_X1 U15059 ( .A1(n13107), .A2(n12894), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12820), .ZN(n12821) );
  AOI21_X1 U15060 ( .B1(n13105), .B2(n12897), .A(n12821), .ZN(n12822) );
  OAI211_X1 U15061 ( .C1(n13330), .C2(n12900), .A(n12823), .B(n12822), .ZN(
        P2_U3195) );
  OAI211_X1 U15062 ( .C1(n12824), .C2(n12826), .A(n12825), .B(n12887), .ZN(
        n12832) );
  OAI22_X1 U15063 ( .A1(n12828), .A2(n12891), .B1(n12827), .B2(n12889), .ZN(
        n13043) );
  OAI22_X1 U15064 ( .A1(n13053), .A2(n12894), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12829), .ZN(n12830) );
  AOI21_X1 U15065 ( .B1(n13043), .B2(n12897), .A(n12830), .ZN(n12831) );
  OAI211_X1 U15066 ( .C1(n13319), .C2(n12900), .A(n12832), .B(n12831), .ZN(
        P2_U3197) );
  INV_X1 U15067 ( .A(n13294), .ZN(n12841) );
  OAI21_X1 U15068 ( .B1(n12834), .B2(n12833), .A(n12844), .ZN(n12835) );
  NAND2_X1 U15069 ( .A1(n12835), .A2(n12887), .ZN(n12840) );
  INV_X1 U15070 ( .A(n13193), .ZN(n12838) );
  AOI22_X1 U15071 ( .A1(n12928), .A2(n12902), .B1(n12901), .B2(n12930), .ZN(
        n13187) );
  OAI22_X1 U15072 ( .A1(n12906), .A2(n13187), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12836), .ZN(n12837) );
  AOI21_X1 U15073 ( .B1(n12838), .B2(n12903), .A(n12837), .ZN(n12839) );
  OAI211_X1 U15074 ( .C1(n12841), .C2(n12900), .A(n12840), .B(n12839), .ZN(
        P2_U3198) );
  INV_X1 U15075 ( .A(n13289), .ZN(n13179) );
  AND3_X1 U15076 ( .A1(n12844), .A2(n12843), .A3(n12842), .ZN(n12845) );
  OAI21_X1 U15077 ( .B1(n12846), .B2(n12845), .A(n12887), .ZN(n12850) );
  INV_X1 U15078 ( .A(n12847), .ZN(n13176) );
  AOI22_X1 U15079 ( .A1(n12927), .A2(n12902), .B1(n12901), .B2(n12929), .ZN(
        n13170) );
  OAI22_X1 U15080 ( .A1(n13170), .A2(n12906), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14802), .ZN(n12848) );
  AOI21_X1 U15081 ( .B1(n13176), .B2(n12903), .A(n12848), .ZN(n12849) );
  OAI211_X1 U15082 ( .C1(n13179), .C2(n12900), .A(n12850), .B(n12849), .ZN(
        P2_U3200) );
  OAI211_X1 U15083 ( .C1(n12853), .C2(n12852), .A(n12851), .B(n12887), .ZN(
        n12859) );
  OAI22_X1 U15084 ( .A1(n12890), .A2(n12891), .B1(n12854), .B2(n12889), .ZN(
        n13060) );
  INV_X1 U15085 ( .A(n13067), .ZN(n12856) );
  OAI22_X1 U15086 ( .A1(n12856), .A2(n12894), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12855), .ZN(n12857) );
  AOI21_X1 U15087 ( .B1(n13060), .B2(n12897), .A(n12857), .ZN(n12858) );
  OAI211_X1 U15088 ( .C1(n13323), .C2(n12900), .A(n12859), .B(n12858), .ZN(
        P2_U3201) );
  NAND2_X1 U15089 ( .A1(n6788), .A2(n12860), .ZN(n12861) );
  XNOR2_X1 U15090 ( .A(n12862), .B(n12861), .ZN(n12868) );
  AND2_X1 U15091 ( .A1(n12926), .A2(n12901), .ZN(n12863) );
  AOI21_X1 U15092 ( .B1(n12924), .B2(n12902), .A(n12863), .ZN(n13121) );
  OAI22_X1 U15093 ( .A1(n13121), .A2(n12906), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12864), .ZN(n12865) );
  AOI21_X1 U15094 ( .B1(n13127), .B2(n12903), .A(n12865), .ZN(n12867) );
  NAND2_X1 U15095 ( .A1(n13273), .A2(n12913), .ZN(n12866) );
  OAI211_X1 U15096 ( .C1(n12868), .C2(n12908), .A(n12867), .B(n12866), .ZN(
        P2_U3205) );
  AND2_X1 U15097 ( .A1(n12924), .A2(n12901), .ZN(n12869) );
  AOI21_X1 U15098 ( .B1(n12922), .B2(n12902), .A(n12869), .ZN(n13088) );
  AOI22_X1 U15099 ( .A1(n13097), .A2(n12903), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12870) );
  OAI21_X1 U15100 ( .B1(n13088), .B2(n12906), .A(n12870), .ZN(n12875) );
  AOI211_X1 U15101 ( .C1(n12873), .C2(n12872), .A(n12908), .B(n12871), .ZN(
        n12874) );
  AOI211_X1 U15102 ( .C1(n13262), .C2(n12913), .A(n12875), .B(n12874), .ZN(
        n12876) );
  INV_X1 U15103 ( .A(n12876), .ZN(P2_U3207) );
  OAI211_X1 U15104 ( .C1(n12879), .C2(n12878), .A(n12877), .B(n12887), .ZN(
        n12883) );
  INV_X1 U15105 ( .A(n12880), .ZN(n13155) );
  AOI22_X1 U15106 ( .A1(n12926), .A2(n12902), .B1(n12901), .B2(n12928), .ZN(
        n13149) );
  OAI22_X1 U15107 ( .A1(n13149), .A2(n12906), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14818), .ZN(n12881) );
  AOI21_X1 U15108 ( .B1(n13155), .B2(n12903), .A(n12881), .ZN(n12882) );
  OAI211_X1 U15109 ( .C1(n13157), .C2(n12900), .A(n12883), .B(n12882), .ZN(
        P2_U3210) );
  OAI21_X1 U15110 ( .B1(n12886), .B2(n12885), .A(n12884), .ZN(n12888) );
  NAND2_X1 U15111 ( .A1(n12888), .A2(n12887), .ZN(n12899) );
  OAI22_X1 U15112 ( .A1(n12892), .A2(n12891), .B1(n12890), .B2(n12889), .ZN(
        n13030) );
  INV_X1 U15113 ( .A(n13034), .ZN(n12895) );
  OAI22_X1 U15114 ( .A1(n12895), .A2(n12894), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12893), .ZN(n12896) );
  AOI21_X1 U15115 ( .B1(n13030), .B2(n12897), .A(n12896), .ZN(n12898) );
  OAI211_X1 U15116 ( .C1(n13036), .C2(n12900), .A(n12899), .B(n12898), .ZN(
        P2_U3212) );
  AOI22_X1 U15117 ( .A1(n12929), .A2(n12902), .B1(n12931), .B2(n12901), .ZN(
        n13300) );
  NAND2_X1 U15118 ( .A1(n12903), .A2(n13207), .ZN(n12905) );
  OAI211_X1 U15119 ( .C1(n13300), .C2(n12906), .A(n12905), .B(n12904), .ZN(
        n12912) );
  AOI211_X1 U15120 ( .C1(n12910), .C2(n12909), .A(n12908), .B(n12907), .ZN(
        n12911) );
  AOI211_X1 U15121 ( .C1(n13336), .C2(n12913), .A(n12912), .B(n12911), .ZN(
        n12914) );
  INV_X1 U15122 ( .A(n12914), .ZN(P2_U3213) );
  MUX2_X1 U15123 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n12992), .S(n6642), .Z(
        P2_U3562) );
  MUX2_X1 U15124 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n12915), .S(n6642), .Z(
        P2_U3561) );
  MUX2_X1 U15125 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n12916), .S(n6642), .Z(
        P2_U3560) );
  MUX2_X1 U15126 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n12917), .S(P2_U3947), .Z(
        P2_U3559) );
  MUX2_X1 U15127 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n12918), .S(P2_U3947), .Z(
        P2_U3558) );
  MUX2_X1 U15128 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n12919), .S(P2_U3947), .Z(
        P2_U3557) );
  MUX2_X1 U15129 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n12920), .S(P2_U3947), .Z(
        P2_U3556) );
  MUX2_X1 U15130 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n12921), .S(P2_U3947), .Z(
        P2_U3555) );
  MUX2_X1 U15131 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n12922), .S(P2_U3947), .Z(
        P2_U3554) );
  MUX2_X1 U15132 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n12923), .S(n6642), .Z(
        P2_U3553) );
  MUX2_X1 U15133 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n12924), .S(n6642), .Z(
        P2_U3552) );
  MUX2_X1 U15134 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n12925), .S(n6642), .Z(
        P2_U3551) );
  MUX2_X1 U15135 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n12926), .S(n6642), .Z(
        P2_U3550) );
  MUX2_X1 U15136 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n12927), .S(n6642), .Z(
        P2_U3549) );
  MUX2_X1 U15137 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n12928), .S(n6642), .Z(
        P2_U3548) );
  MUX2_X1 U15138 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n12929), .S(n6642), .Z(
        P2_U3547) );
  MUX2_X1 U15139 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n12930), .S(n6642), .Z(
        P2_U3546) );
  MUX2_X1 U15140 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n12931), .S(n6642), .Z(
        P2_U3545) );
  MUX2_X1 U15141 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n12932), .S(n6642), .Z(
        P2_U3544) );
  MUX2_X1 U15142 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n12933), .S(n6642), .Z(
        P2_U3543) );
  MUX2_X1 U15143 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n12934), .S(n6642), .Z(
        P2_U3542) );
  MUX2_X1 U15144 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n12935), .S(n6642), .Z(
        P2_U3541) );
  MUX2_X1 U15145 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n12936), .S(n6642), .Z(
        P2_U3540) );
  MUX2_X1 U15146 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n12937), .S(n6642), .Z(
        P2_U3539) );
  MUX2_X1 U15147 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n12938), .S(n6642), .Z(
        P2_U3538) );
  MUX2_X1 U15148 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n12939), .S(n6642), .Z(
        P2_U3537) );
  MUX2_X1 U15149 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n12940), .S(n6642), .Z(
        P2_U3536) );
  MUX2_X1 U15150 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n12941), .S(n6642), .Z(
        P2_U3535) );
  MUX2_X1 U15151 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n12942), .S(n6642), .Z(
        P2_U3534) );
  MUX2_X1 U15152 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n12943), .S(n6642), .Z(
        P2_U3533) );
  MUX2_X1 U15153 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n12944), .S(n6642), .Z(
        P2_U3532) );
  MUX2_X1 U15154 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n11843), .S(n6642), .Z(
        P2_U3531) );
  INV_X1 U15155 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n12946) );
  OAI21_X1 U15156 ( .B1(n14817), .B2(n12946), .A(n12945), .ZN(n12947) );
  AOI21_X1 U15157 ( .B1(n12951), .B2(n14809), .A(n12947), .ZN(n12958) );
  INV_X1 U15158 ( .A(n14819), .ZN(n14787) );
  OAI211_X1 U15159 ( .C1(n12950), .C2(n12949), .A(n14787), .B(n12948), .ZN(
        n12957) );
  MUX2_X1 U15160 ( .A(n9770), .B(P2_REG2_REG_7__SCAN_IN), .S(n12951), .Z(
        n12952) );
  NAND3_X1 U15161 ( .A1(n14728), .A2(n12953), .A3(n12952), .ZN(n12954) );
  NAND3_X1 U15162 ( .A1(n12955), .A2(n14811), .A3(n12954), .ZN(n12956) );
  NAND3_X1 U15163 ( .A1(n12958), .A2(n12957), .A3(n12956), .ZN(P2_U3221) );
  INV_X1 U15164 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n14821) );
  INV_X1 U15165 ( .A(n14801), .ZN(n12963) );
  NOR2_X1 U15166 ( .A1(n12960), .A2(n12959), .ZN(n12962) );
  NOR2_X1 U15167 ( .A1(n12962), .A2(n12961), .ZN(n14793) );
  XOR2_X1 U15168 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n14801), .Z(n14792) );
  NOR2_X1 U15169 ( .A1(n14793), .A2(n14792), .ZN(n14791) );
  AOI21_X1 U15170 ( .B1(n12963), .B2(P2_REG1_REG_16__SCAN_IN), .A(n14791), 
        .ZN(n14805) );
  XNOR2_X1 U15171 ( .A(n14808), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n14804) );
  NOR2_X1 U15172 ( .A1(n14805), .A2(n14804), .ZN(n14803) );
  AOI21_X1 U15173 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n14808), .A(n14803), 
        .ZN(n12964) );
  XNOR2_X1 U15174 ( .A(n14832), .B(n12964), .ZN(n14822) );
  NOR2_X1 U15175 ( .A1(n14821), .A2(n14822), .ZN(n14820) );
  NOR2_X1 U15176 ( .A1(n12964), .A2(n14832), .ZN(n12965) );
  NOR2_X1 U15177 ( .A1(n14820), .A2(n12965), .ZN(n12966) );
  XOR2_X1 U15178 ( .A(n12966), .B(n15340), .Z(n12982) );
  NOR2_X1 U15179 ( .A1(n12973), .A2(n12967), .ZN(n12968) );
  AOI21_X1 U15180 ( .B1(n12967), .B2(n12973), .A(n12968), .ZN(n14812) );
  XNOR2_X1 U15181 ( .A(n14801), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n14797) );
  NAND2_X1 U15182 ( .A1(n12970), .A2(n12969), .ZN(n12972) );
  NAND2_X1 U15183 ( .A1(n12972), .A2(n12971), .ZN(n14798) );
  NAND2_X1 U15184 ( .A1(n14797), .A2(n14798), .ZN(n14796) );
  OAI21_X1 U15185 ( .B1(n14801), .B2(n15405), .A(n14796), .ZN(n14813) );
  NAND2_X1 U15186 ( .A1(n14812), .A2(n14813), .ZN(n14810) );
  OAI21_X1 U15187 ( .B1(n12967), .B2(n12973), .A(n14810), .ZN(n12974) );
  XNOR2_X1 U15188 ( .A(n12975), .B(n12974), .ZN(n14827) );
  NOR2_X1 U15189 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n14827), .ZN(n14826) );
  NOR2_X1 U15190 ( .A1(n12975), .A2(n12974), .ZN(n12976) );
  NOR2_X1 U15191 ( .A1(n14826), .A2(n12976), .ZN(n12977) );
  XOR2_X1 U15192 ( .A(n12977), .B(P2_REG2_REG_19__SCAN_IN), .Z(n12981) );
  INV_X1 U15193 ( .A(n12981), .ZN(n12978) );
  NAND2_X1 U15194 ( .A1(n12978), .A2(n14811), .ZN(n12979) );
  OAI211_X1 U15195 ( .C1(n12982), .C2(n14819), .A(n14833), .B(n12979), .ZN(
        n12980) );
  INV_X1 U15196 ( .A(n12980), .ZN(n12985) );
  AOI22_X1 U15197 ( .A1(n12982), .A2(n14787), .B1(n14811), .B2(n12981), .ZN(
        n12984) );
  MUX2_X1 U15198 ( .A(n12985), .B(n12984), .S(n12983), .Z(n12987) );
  OAI211_X1 U15199 ( .C1(n12988), .C2(n14817), .A(n12987), .B(n12986), .ZN(
        P2_U3233) );
  NOR2_X1 U15200 ( .A1(n12995), .A2(n13224), .ZN(n12997) );
  XNOR2_X1 U15201 ( .A(n12997), .B(n12989), .ZN(n13219) );
  NAND2_X1 U15202 ( .A1(n13219), .A2(n14844), .ZN(n12994) );
  INV_X1 U15203 ( .A(n12990), .ZN(n12991) );
  AND2_X1 U15204 ( .A1(n12992), .A2(n12991), .ZN(n13218) );
  INV_X1 U15205 ( .A(n13218), .ZN(n13222) );
  NOR2_X1 U15206 ( .A1(n13211), .A2(n13222), .ZN(n12999) );
  AOI21_X1 U15207 ( .B1(n13211), .B2(P2_REG2_REG_31__SCAN_IN), .A(n12999), 
        .ZN(n12993) );
  OAI211_X1 U15208 ( .C1(n13308), .C2(n14835), .A(n12994), .B(n12993), .ZN(
        P2_U3234) );
  AND2_X1 U15209 ( .A1(n13224), .A2(n12995), .ZN(n12996) );
  NOR2_X1 U15210 ( .A1(n13312), .A2(n14835), .ZN(n12998) );
  AOI211_X1 U15211 ( .C1(n13211), .C2(P2_REG2_REG_30__SCAN_IN), .A(n12999), 
        .B(n12998), .ZN(n13000) );
  OAI21_X1 U15212 ( .B1(n13213), .B2(n13223), .A(n13000), .ZN(P2_U3235) );
  OAI21_X1 U15213 ( .B1(n13002), .B2(n13003), .A(n13001), .ZN(n13228) );
  AOI21_X1 U15214 ( .B1(n13004), .B2(n13003), .A(n13171), .ZN(n13007) );
  AOI21_X1 U15215 ( .B1(n13007), .B2(n13006), .A(n13005), .ZN(n13227) );
  INV_X1 U15216 ( .A(n13227), .ZN(n13012) );
  NAND2_X1 U15217 ( .A1(n13229), .A2(n13018), .ZN(n13008) );
  NAND2_X1 U15218 ( .A1(n13008), .A2(n14313), .ZN(n13009) );
  OR2_X1 U15219 ( .A1(n6684), .A2(n13009), .ZN(n13226) );
  OAI22_X1 U15220 ( .A1(n13226), .A2(n13195), .B1(n13010), .B2(n13194), .ZN(
        n13011) );
  OAI21_X1 U15221 ( .B1(n13012), .B2(n13011), .A(n14837), .ZN(n13014) );
  AOI22_X1 U15222 ( .A1(n13229), .A2(n14307), .B1(n13211), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n13013) );
  OAI211_X1 U15223 ( .C1(n13182), .C2(n13228), .A(n13014), .B(n13013), .ZN(
        P2_U3237) );
  XNOR2_X1 U15224 ( .A(n13015), .B(n13020), .ZN(n13017) );
  AOI21_X1 U15225 ( .B1(n13017), .B2(n14304), .A(n13016), .ZN(n13235) );
  OAI211_X1 U15226 ( .C1(n13019), .C2(n13032), .A(n14313), .B(n13018), .ZN(
        n13234) );
  NAND2_X1 U15227 ( .A1(n13021), .A2(n13020), .ZN(n13230) );
  NAND3_X1 U15228 ( .A1(n13231), .A2(n13230), .A3(n14316), .ZN(n13026) );
  OAI22_X1 U15229 ( .A1(n13023), .A2(n13194), .B1(n13022), .B2(n14837), .ZN(
        n13024) );
  AOI21_X1 U15230 ( .B1(n13232), .B2(n14307), .A(n13024), .ZN(n13025) );
  OAI211_X1 U15231 ( .C1(n13234), .C2(n13213), .A(n13026), .B(n13025), .ZN(
        n13027) );
  INV_X1 U15232 ( .A(n13027), .ZN(n13028) );
  OAI21_X1 U15233 ( .B1(n13235), .B2(n13216), .A(n13028), .ZN(P2_U3238) );
  XNOR2_X1 U15234 ( .A(n13029), .B(n13037), .ZN(n13031) );
  AOI21_X1 U15235 ( .B1(n13031), .B2(n14304), .A(n13030), .ZN(n13240) );
  OAI21_X1 U15236 ( .B1(n13036), .B2(n13051), .A(n14313), .ZN(n13033) );
  NOR2_X1 U15237 ( .A1(n13033), .A2(n13032), .ZN(n13237) );
  AOI22_X1 U15238 ( .A1(n13034), .A2(n14841), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n13216), .ZN(n13035) );
  OAI21_X1 U15239 ( .B1(n13036), .B2(n14835), .A(n13035), .ZN(n13040) );
  XNOR2_X1 U15240 ( .A(n13038), .B(n13037), .ZN(n13241) );
  NOR2_X1 U15241 ( .A1(n13241), .A2(n13182), .ZN(n13039) );
  AOI211_X1 U15242 ( .C1(n13237), .C2(n14315), .A(n13040), .B(n13039), .ZN(
        n13041) );
  OAI21_X1 U15243 ( .B1(n13211), .B2(n13240), .A(n13041), .ZN(P2_U3239) );
  XNOR2_X1 U15244 ( .A(n13042), .B(n13045), .ZN(n13044) );
  AOI21_X1 U15245 ( .B1(n13044), .B2(n14304), .A(n13043), .ZN(n13245) );
  NAND2_X1 U15246 ( .A1(n13046), .A2(n13045), .ZN(n13047) );
  NAND2_X1 U15247 ( .A1(n13048), .A2(n13047), .ZN(n13244) );
  NOR2_X1 U15248 ( .A1(n13319), .A2(n13065), .ZN(n13050) );
  OR3_X1 U15249 ( .A1(n13051), .A2(n13050), .A3(n13049), .ZN(n13242) );
  OAI22_X1 U15250 ( .A1(n13053), .A2(n13194), .B1(n13052), .B2(n14837), .ZN(
        n13054) );
  AOI21_X1 U15251 ( .B1(n13248), .B2(n14307), .A(n13054), .ZN(n13055) );
  OAI21_X1 U15252 ( .B1(n13242), .B2(n13213), .A(n13055), .ZN(n13056) );
  AOI21_X1 U15253 ( .B1(n13244), .B2(n14316), .A(n13056), .ZN(n13057) );
  OAI21_X1 U15254 ( .B1(n13245), .B2(n13216), .A(n13057), .ZN(P2_U3240) );
  XNOR2_X1 U15255 ( .A(n13059), .B(n13058), .ZN(n13062) );
  INV_X1 U15256 ( .A(n13060), .ZN(n13061) );
  OAI21_X1 U15257 ( .B1(n13062), .B2(n13171), .A(n13061), .ZN(n13250) );
  INV_X1 U15258 ( .A(n13250), .ZN(n13072) );
  XNOR2_X1 U15259 ( .A(n13064), .B(n13063), .ZN(n13252) );
  AOI211_X1 U15260 ( .C1(n13066), .C2(n13080), .A(n13049), .B(n13065), .ZN(
        n13251) );
  NAND2_X1 U15261 ( .A1(n13251), .A2(n14315), .ZN(n13069) );
  AOI22_X1 U15262 ( .A1(n13067), .A2(n14841), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n13216), .ZN(n13068) );
  OAI211_X1 U15263 ( .C1(n13323), .C2(n14835), .A(n13069), .B(n13068), .ZN(
        n13070) );
  AOI21_X1 U15264 ( .B1(n13252), .B2(n14316), .A(n13070), .ZN(n13071) );
  OAI21_X1 U15265 ( .B1(n13072), .B2(n13216), .A(n13071), .ZN(P2_U3241) );
  XNOR2_X1 U15266 ( .A(n13073), .B(n13074), .ZN(n13260) );
  OAI21_X1 U15267 ( .B1(n6677), .B2(n8167), .A(n13075), .ZN(n13077) );
  AOI21_X1 U15268 ( .B1(n13077), .B2(n14304), .A(n13076), .ZN(n13259) );
  OAI21_X1 U15269 ( .B1(n13078), .B2(n13194), .A(n13259), .ZN(n13079) );
  NAND2_X1 U15270 ( .A1(n13079), .A2(n14837), .ZN(n13086) );
  INV_X1 U15271 ( .A(n13080), .ZN(n13081) );
  AOI211_X1 U15272 ( .C1(n13257), .C2(n13095), .A(n13049), .B(n13081), .ZN(
        n13256) );
  OAI22_X1 U15273 ( .A1(n13083), .A2(n14835), .B1(n14837), .B2(n13082), .ZN(
        n13084) );
  AOI21_X1 U15274 ( .B1(n13256), .B2(n14315), .A(n13084), .ZN(n13085) );
  OAI211_X1 U15275 ( .C1(n13260), .C2(n13182), .A(n13086), .B(n13085), .ZN(
        P2_U3242) );
  AOI21_X1 U15276 ( .B1(n13087), .B2(n13094), .A(n13171), .ZN(n13091) );
  INV_X1 U15277 ( .A(n13088), .ZN(n13089) );
  AOI21_X1 U15278 ( .B1(n13091), .B2(n13090), .A(n13089), .ZN(n13264) );
  OAI21_X1 U15279 ( .B1(n13092), .B2(n13094), .A(n13093), .ZN(n13265) );
  INV_X1 U15280 ( .A(n13265), .ZN(n13102) );
  INV_X1 U15281 ( .A(n13262), .ZN(n13100) );
  AOI21_X1 U15282 ( .B1(n13262), .B2(n13109), .A(n13049), .ZN(n13096) );
  AND2_X1 U15283 ( .A1(n13096), .A2(n13095), .ZN(n13261) );
  NAND2_X1 U15284 ( .A1(n13261), .A2(n14315), .ZN(n13099) );
  AOI22_X1 U15285 ( .A1(n13097), .A2(n14841), .B1(P2_REG2_REG_22__SCAN_IN), 
        .B2(n13216), .ZN(n13098) );
  OAI211_X1 U15286 ( .C1(n13100), .C2(n14835), .A(n13099), .B(n13098), .ZN(
        n13101) );
  AOI21_X1 U15287 ( .B1(n13102), .B2(n14316), .A(n13101), .ZN(n13103) );
  OAI21_X1 U15288 ( .B1(n13211), .B2(n13264), .A(n13103), .ZN(P2_U3243) );
  XNOR2_X1 U15289 ( .A(n13104), .B(n13112), .ZN(n13106) );
  AOI21_X1 U15290 ( .B1(n13106), .B2(n14304), .A(n13105), .ZN(n13267) );
  INV_X1 U15291 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n13108) );
  OAI22_X1 U15292 ( .A1(n13108), .A2(n14837), .B1(n13107), .B2(n13194), .ZN(
        n13111) );
  OAI211_X1 U15293 ( .C1(n13126), .C2(n13330), .A(n14313), .B(n13109), .ZN(
        n13266) );
  NOR2_X1 U15294 ( .A1(n13266), .A2(n13213), .ZN(n13110) );
  AOI211_X1 U15295 ( .C1(n14307), .C2(n13270), .A(n13111), .B(n13110), .ZN(
        n13116) );
  INV_X1 U15296 ( .A(n13112), .ZN(n13113) );
  XNOR2_X1 U15297 ( .A(n13114), .B(n13113), .ZN(n13268) );
  OR2_X1 U15298 ( .A1(n13268), .A2(n13182), .ZN(n13115) );
  OAI211_X1 U15299 ( .C1(n13267), .C2(n13216), .A(n13116), .B(n13115), .ZN(
        P2_U3244) );
  XNOR2_X1 U15300 ( .A(n13117), .B(n13120), .ZN(n13276) );
  OAI21_X1 U15301 ( .B1(n13120), .B2(n13119), .A(n13118), .ZN(n13123) );
  INV_X1 U15302 ( .A(n13121), .ZN(n13122) );
  AOI21_X1 U15303 ( .B1(n13123), .B2(n14304), .A(n13122), .ZN(n13275) );
  INV_X1 U15304 ( .A(n13275), .ZN(n13131) );
  NAND2_X1 U15305 ( .A1(n13138), .A2(n13273), .ZN(n13124) );
  NAND2_X1 U15306 ( .A1(n13124), .A2(n14313), .ZN(n13125) );
  NOR2_X1 U15307 ( .A1(n13126), .A2(n13125), .ZN(n13272) );
  NAND2_X1 U15308 ( .A1(n13272), .A2(n14315), .ZN(n13129) );
  AOI22_X1 U15309 ( .A1(P2_REG2_REG_20__SCAN_IN), .A2(n13216), .B1(n13127), 
        .B2(n14841), .ZN(n13128) );
  OAI211_X1 U15310 ( .C1(n7229), .C2(n14835), .A(n13129), .B(n13128), .ZN(
        n13130) );
  AOI21_X1 U15311 ( .B1(n13131), .B2(n14837), .A(n13130), .ZN(n13132) );
  OAI21_X1 U15312 ( .B1(n13276), .B2(n13182), .A(n13132), .ZN(P2_U3245) );
  XNOR2_X1 U15313 ( .A(n13133), .B(n13136), .ZN(n13135) );
  AOI21_X1 U15314 ( .B1(n13135), .B2(n14304), .A(n13134), .ZN(n13280) );
  XOR2_X1 U15315 ( .A(n13137), .B(n13136), .Z(n13281) );
  INV_X1 U15316 ( .A(n13281), .ZN(n13146) );
  INV_X1 U15317 ( .A(n13278), .ZN(n13144) );
  AOI21_X1 U15318 ( .B1(n13152), .B2(n13278), .A(n13049), .ZN(n13139) );
  AND2_X1 U15319 ( .A1(n13139), .A2(n13138), .ZN(n13277) );
  NAND2_X1 U15320 ( .A1(n13277), .A2(n14315), .ZN(n13143) );
  INV_X1 U15321 ( .A(n13140), .ZN(n13141) );
  AOI22_X1 U15322 ( .A1(n13216), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13141), 
        .B2(n14841), .ZN(n13142) );
  OAI211_X1 U15323 ( .C1(n13144), .C2(n14835), .A(n13143), .B(n13142), .ZN(
        n13145) );
  AOI21_X1 U15324 ( .B1(n13146), .B2(n14316), .A(n13145), .ZN(n13147) );
  OAI21_X1 U15325 ( .B1(n13211), .B2(n13280), .A(n13147), .ZN(P2_U3246) );
  XNOR2_X1 U15326 ( .A(n13148), .B(n13161), .ZN(n13151) );
  INV_X1 U15327 ( .A(n13149), .ZN(n13150) );
  AOI21_X1 U15328 ( .B1(n13151), .B2(n14304), .A(n13150), .ZN(n13285) );
  INV_X1 U15329 ( .A(n13175), .ZN(n13154) );
  INV_X1 U15330 ( .A(n13152), .ZN(n13153) );
  AOI211_X1 U15331 ( .C1(n13283), .C2(n13154), .A(n13049), .B(n13153), .ZN(
        n13282) );
  AOI22_X1 U15332 ( .A1(n13216), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13155), 
        .B2(n14841), .ZN(n13156) );
  OAI21_X1 U15333 ( .B1(n13157), .B2(n14835), .A(n13156), .ZN(n13163) );
  INV_X1 U15334 ( .A(n13158), .ZN(n13159) );
  AOI21_X1 U15335 ( .B1(n13161), .B2(n13160), .A(n13159), .ZN(n13286) );
  NOR2_X1 U15336 ( .A1(n13286), .A2(n13182), .ZN(n13162) );
  AOI211_X1 U15337 ( .C1(n13282), .C2(n14315), .A(n13163), .B(n13162), .ZN(
        n13164) );
  OAI21_X1 U15338 ( .B1(n13211), .B2(n13285), .A(n13164), .ZN(P2_U3247) );
  XNOR2_X1 U15339 ( .A(n13165), .B(n13167), .ZN(n13291) );
  NAND3_X1 U15340 ( .A1(n13184), .A2(n13167), .A3(n13166), .ZN(n13168) );
  AND2_X1 U15341 ( .A1(n13169), .A2(n13168), .ZN(n13172) );
  OAI21_X1 U15342 ( .B1(n13172), .B2(n13171), .A(n13170), .ZN(n13287) );
  NAND2_X1 U15343 ( .A1(n13191), .A2(n13289), .ZN(n13173) );
  NAND2_X1 U15344 ( .A1(n13173), .A2(n14313), .ZN(n13174) );
  NOR2_X1 U15345 ( .A1(n13175), .A2(n13174), .ZN(n13288) );
  NAND2_X1 U15346 ( .A1(n13288), .A2(n14315), .ZN(n13178) );
  AOI22_X1 U15347 ( .A1(n13216), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n13176), 
        .B2(n14841), .ZN(n13177) );
  OAI211_X1 U15348 ( .C1(n13179), .C2(n14835), .A(n13178), .B(n13177), .ZN(
        n13180) );
  AOI21_X1 U15349 ( .B1(n13287), .B2(n14837), .A(n13180), .ZN(n13181) );
  OAI21_X1 U15350 ( .B1(n13291), .B2(n13182), .A(n13181), .ZN(P2_U3248) );
  INV_X1 U15351 ( .A(n13183), .ZN(n13186) );
  INV_X1 U15352 ( .A(n13198), .ZN(n13185) );
  OAI21_X1 U15353 ( .B1(n13186), .B2(n13185), .A(n13184), .ZN(n13189) );
  INV_X1 U15354 ( .A(n13187), .ZN(n13188) );
  AOI21_X1 U15355 ( .B1(n13189), .B2(n14304), .A(n13188), .ZN(n13297) );
  INV_X1 U15356 ( .A(n13297), .ZN(n13197) );
  AOI21_X1 U15357 ( .B1(n13190), .B2(n13294), .A(n11181), .ZN(n13192) );
  NAND2_X1 U15358 ( .A1(n13192), .A2(n13191), .ZN(n13296) );
  OAI22_X1 U15359 ( .A1(n13296), .A2(n13195), .B1(n13194), .B2(n13193), .ZN(
        n13196) );
  OAI21_X1 U15360 ( .B1(n13197), .B2(n13196), .A(n14837), .ZN(n13202) );
  AOI22_X1 U15361 ( .A1(n13294), .A2(n14307), .B1(P2_REG2_REG_16__SCAN_IN), 
        .B2(n13216), .ZN(n13201) );
  OR2_X1 U15362 ( .A1(n13199), .A2(n13198), .ZN(n13293) );
  NAND3_X1 U15363 ( .A1(n13293), .A2(n13292), .A3(n14316), .ZN(n13200) );
  NAND3_X1 U15364 ( .A1(n13202), .A2(n13201), .A3(n13200), .ZN(P2_U3249) );
  INV_X1 U15365 ( .A(n13300), .ZN(n13206) );
  XNOR2_X1 U15366 ( .A(n13203), .B(n13208), .ZN(n13204) );
  NAND2_X1 U15367 ( .A1(n13204), .A2(n14304), .ZN(n13301) );
  INV_X1 U15368 ( .A(n13301), .ZN(n13205) );
  AOI211_X1 U15369 ( .C1(n14841), .C2(n13207), .A(n13206), .B(n13205), .ZN(
        n13217) );
  XNOR2_X1 U15370 ( .A(n13209), .B(n13208), .ZN(n13303) );
  XOR2_X1 U15371 ( .A(n14312), .B(n13336), .Z(n13210) );
  NAND2_X1 U15372 ( .A1(n13210), .A2(n14313), .ZN(n13299) );
  AOI22_X1 U15373 ( .A1(n13336), .A2(n14307), .B1(n13211), .B2(
        P2_REG2_REG_15__SCAN_IN), .ZN(n13212) );
  OAI21_X1 U15374 ( .B1(n13299), .B2(n13213), .A(n13212), .ZN(n13214) );
  AOI21_X1 U15375 ( .B1(n13303), .B2(n14316), .A(n13214), .ZN(n13215) );
  OAI21_X1 U15376 ( .B1(n13217), .B2(n13216), .A(n13215), .ZN(P2_U3250) );
  INV_X1 U15377 ( .A(n13304), .ZN(n13255) );
  INV_X1 U15378 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n13220) );
  AOI21_X1 U15379 ( .B1(n13219), .B2(n14313), .A(n13218), .ZN(n13306) );
  MUX2_X1 U15380 ( .A(n13220), .B(n13306), .S(n14934), .Z(n13221) );
  OAI21_X1 U15381 ( .B1(n13308), .B2(n13255), .A(n13221), .ZN(P2_U3530) );
  INV_X1 U15382 ( .A(n13225), .ZN(P2_U3529) );
  NAND3_X1 U15383 ( .A1(n13231), .A2(n14905), .A3(n13230), .ZN(n13236) );
  NAND2_X1 U15384 ( .A1(n13232), .A2(n14892), .ZN(n13233) );
  NAND4_X1 U15385 ( .A1(n13236), .A2(n13235), .A3(n13234), .A4(n13233), .ZN(
        n13314) );
  MUX2_X1 U15386 ( .A(n13314), .B(P2_REG1_REG_27__SCAN_IN), .S(n14932), .Z(
        P2_U3526) );
  AOI21_X1 U15387 ( .B1(n14892), .B2(n13238), .A(n13237), .ZN(n13239) );
  OAI211_X1 U15388 ( .C1(n13241), .C2(n14895), .A(n13240), .B(n13239), .ZN(
        n13315) );
  MUX2_X1 U15389 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13315), .S(n14934), .Z(
        P2_U3525) );
  INV_X1 U15390 ( .A(n13242), .ZN(n13243) );
  AOI21_X1 U15391 ( .B1(n13244), .B2(n14905), .A(n13243), .ZN(n13246) );
  NAND2_X1 U15392 ( .A1(n13246), .A2(n13245), .ZN(n13316) );
  MUX2_X1 U15393 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13316), .S(n14934), .Z(
        n13247) );
  AOI21_X1 U15394 ( .B1(n13304), .B2(n13248), .A(n13247), .ZN(n13249) );
  INV_X1 U15395 ( .A(n13249), .ZN(P2_U3524) );
  AOI211_X1 U15396 ( .C1(n14905), .C2(n13252), .A(n13251), .B(n13250), .ZN(
        n13320) );
  MUX2_X1 U15397 ( .A(n13253), .B(n13320), .S(n14934), .Z(n13254) );
  OAI21_X1 U15398 ( .B1(n13323), .B2(n13255), .A(n13254), .ZN(P2_U3523) );
  AOI21_X1 U15399 ( .B1(n14892), .B2(n13257), .A(n13256), .ZN(n13258) );
  OAI211_X1 U15400 ( .C1(n14895), .C2(n13260), .A(n13259), .B(n13258), .ZN(
        n13324) );
  MUX2_X1 U15401 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13324), .S(n14934), .Z(
        P2_U3522) );
  AOI21_X1 U15402 ( .B1(n14892), .B2(n13262), .A(n13261), .ZN(n13263) );
  OAI211_X1 U15403 ( .C1(n13265), .C2(n14895), .A(n13264), .B(n13263), .ZN(
        n13325) );
  MUX2_X1 U15404 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13325), .S(n14934), .Z(
        P2_U3521) );
  OAI211_X1 U15405 ( .C1(n13268), .C2(n14895), .A(n13267), .B(n13266), .ZN(
        n13326) );
  MUX2_X1 U15406 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13326), .S(n14934), .Z(
        n13269) );
  AOI21_X1 U15407 ( .B1(n13304), .B2(n13270), .A(n13269), .ZN(n13271) );
  INV_X1 U15408 ( .A(n13271), .ZN(P2_U3520) );
  AOI21_X1 U15409 ( .B1(n14892), .B2(n13273), .A(n13272), .ZN(n13274) );
  OAI211_X1 U15410 ( .C1(n14895), .C2(n13276), .A(n13275), .B(n13274), .ZN(
        n13331) );
  MUX2_X1 U15411 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13331), .S(n14934), .Z(
        P2_U3519) );
  AOI21_X1 U15412 ( .B1(n14892), .B2(n13278), .A(n13277), .ZN(n13279) );
  OAI211_X1 U15413 ( .C1(n13281), .C2(n14895), .A(n13280), .B(n13279), .ZN(
        n13332) );
  MUX2_X1 U15414 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13332), .S(n14934), .Z(
        P2_U3518) );
  AOI21_X1 U15415 ( .B1(n14892), .B2(n13283), .A(n13282), .ZN(n13284) );
  OAI211_X1 U15416 ( .C1(n13286), .C2(n14895), .A(n13285), .B(n13284), .ZN(
        n13333) );
  MUX2_X1 U15417 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13333), .S(n14934), .Z(
        P2_U3517) );
  AOI211_X1 U15418 ( .C1(n14892), .C2(n13289), .A(n13288), .B(n13287), .ZN(
        n13290) );
  OAI21_X1 U15419 ( .B1(n14895), .B2(n13291), .A(n13290), .ZN(n13334) );
  MUX2_X1 U15420 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13334), .S(n14934), .Z(
        P2_U3516) );
  NAND3_X1 U15421 ( .A1(n13293), .A2(n14905), .A3(n13292), .ZN(n13298) );
  NAND2_X1 U15422 ( .A1(n13294), .A2(n14892), .ZN(n13295) );
  NAND4_X1 U15423 ( .A1(n13298), .A2(n13297), .A3(n13296), .A4(n13295), .ZN(
        n13335) );
  MUX2_X1 U15424 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13335), .S(n14934), .Z(
        P2_U3515) );
  NAND3_X1 U15425 ( .A1(n13301), .A2(n13300), .A3(n13299), .ZN(n13302) );
  AOI21_X1 U15426 ( .B1(n13303), .B2(n14905), .A(n13302), .ZN(n13338) );
  AOI22_X1 U15427 ( .A1(n13336), .A2(n13304), .B1(P2_REG1_REG_15__SCAN_IN), 
        .B2(n14932), .ZN(n13305) );
  OAI21_X1 U15428 ( .B1(n13338), .B2(n14932), .A(n13305), .ZN(P2_U3514) );
  MUX2_X1 U15429 ( .A(n15447), .B(n13306), .S(n14924), .Z(n13307) );
  OAI21_X1 U15430 ( .B1(n13308), .B2(n13329), .A(n13307), .ZN(P2_U3498) );
  MUX2_X1 U15431 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13309), .S(n14924), .Z(
        n13310) );
  INV_X1 U15432 ( .A(n13310), .ZN(n13311) );
  OAI21_X1 U15433 ( .B1(n13312), .B2(n13329), .A(n13311), .ZN(P2_U3497) );
  MUX2_X1 U15434 ( .A(n13314), .B(P2_REG0_REG_27__SCAN_IN), .S(n14922), .Z(
        P2_U3494) );
  MUX2_X1 U15435 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13315), .S(n14924), .Z(
        P2_U3493) );
  MUX2_X1 U15436 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13316), .S(n14924), .Z(
        n13317) );
  INV_X1 U15437 ( .A(n13317), .ZN(n13318) );
  OAI21_X1 U15438 ( .B1(n13319), .B2(n13329), .A(n13318), .ZN(P2_U3492) );
  INV_X1 U15439 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n13321) );
  MUX2_X1 U15440 ( .A(n13321), .B(n13320), .S(n14924), .Z(n13322) );
  OAI21_X1 U15441 ( .B1(n13323), .B2(n13329), .A(n13322), .ZN(P2_U3491) );
  MUX2_X1 U15442 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13324), .S(n14924), .Z(
        P2_U3490) );
  MUX2_X1 U15443 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13325), .S(n14924), .Z(
        P2_U3489) );
  MUX2_X1 U15444 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13326), .S(n14924), .Z(
        n13327) );
  INV_X1 U15445 ( .A(n13327), .ZN(n13328) );
  OAI21_X1 U15446 ( .B1(n13330), .B2(n13329), .A(n13328), .ZN(P2_U3488) );
  MUX2_X1 U15447 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13331), .S(n14924), .Z(
        P2_U3487) );
  MUX2_X1 U15448 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13332), .S(n14924), .Z(
        P2_U3486) );
  MUX2_X1 U15449 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13333), .S(n14924), .Z(
        P2_U3484) );
  MUX2_X1 U15450 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13334), .S(n14924), .Z(
        P2_U3481) );
  MUX2_X1 U15451 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13335), .S(n14924), .Z(
        P2_U3478) );
  AOI22_X1 U15452 ( .A1(n13336), .A2(n8982), .B1(P2_REG0_REG_15__SCAN_IN), 
        .B2(n14922), .ZN(n13337) );
  OAI21_X1 U15453 ( .B1(n13338), .B2(n14922), .A(n13337), .ZN(P2_U3475) );
  INV_X1 U15454 ( .A(n13339), .ZN(n13344) );
  INV_X1 U15455 ( .A(n7710), .ZN(n13340) );
  NOR4_X1 U15456 ( .A1(n13340), .A2(P2_IR_REG_30__SCAN_IN), .A3(n8268), .A4(
        P2_U3088), .ZN(n13341) );
  AOI21_X1 U15457 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n13342), .A(n13341), 
        .ZN(n13343) );
  OAI21_X1 U15458 ( .B1(n13344), .B2(n13359), .A(n13343), .ZN(P2_U3296) );
  OAI222_X1 U15459 ( .A1(n13357), .A2(n15399), .B1(P2_U3088), .B2(n13346), 
        .C1(n13359), .C2(n13345), .ZN(P2_U3297) );
  INV_X1 U15460 ( .A(n13347), .ZN(n14036) );
  OAI222_X1 U15461 ( .A1(n13357), .A2(n13349), .B1(P2_U3088), .B2(n13348), 
        .C1(n13359), .C2(n14036), .ZN(P2_U3298) );
  NAND2_X1 U15462 ( .A1(n13351), .A2(n13350), .ZN(n13353) );
  OAI211_X1 U15463 ( .C1(n13357), .C2(n13354), .A(n13353), .B(n13352), .ZN(
        P2_U3299) );
  OAI222_X1 U15464 ( .A1(n13357), .A2(n13356), .B1(n13359), .B2(n13355), .C1(
        P2_U3088), .C2(n8288), .ZN(P2_U3300) );
  OAI222_X1 U15465 ( .A1(n13360), .A2(P2_U3088), .B1(n13359), .B2(n14041), 
        .C1(n13358), .C2(n13357), .ZN(P2_U3301) );
  MUX2_X1 U15466 ( .A(n13361), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  AOI22_X1 U15467 ( .A1(n13951), .A2(n13445), .B1(n13478), .B2(n13737), .ZN(
        n13471) );
  NAND2_X1 U15468 ( .A1(n13951), .A2(n13475), .ZN(n13363) );
  NAND2_X1 U15469 ( .A1(n13737), .A2(n13445), .ZN(n13362) );
  NAND2_X1 U15470 ( .A1(n13363), .A2(n13362), .ZN(n13364) );
  XNOR2_X1 U15471 ( .A(n13364), .B(n13476), .ZN(n13473) );
  XOR2_X1 U15472 ( .A(n13471), .B(n13473), .Z(n13474) );
  AND2_X1 U15473 ( .A1(n13478), .A2(n13825), .ZN(n13365) );
  AOI21_X1 U15474 ( .B1(n13812), .B2(n13445), .A(n13365), .ZN(n13425) );
  AOI22_X1 U15475 ( .A1(n13812), .A2(n13475), .B1(n13445), .B2(n13825), .ZN(
        n13366) );
  XNOR2_X1 U15476 ( .A(n13366), .B(n13476), .ZN(n13424) );
  AOI22_X1 U15477 ( .A1(n13990), .A2(n13445), .B1(n13478), .B2(n13583), .ZN(
        n13421) );
  INV_X1 U15478 ( .A(n13421), .ZN(n13423) );
  AOI22_X1 U15479 ( .A1(n13990), .A2(n13475), .B1(n13445), .B2(n13583), .ZN(
        n13367) );
  XNOR2_X1 U15480 ( .A(n13367), .B(n13476), .ZN(n13420) );
  INV_X1 U15481 ( .A(n13420), .ZN(n13422) );
  OR2_X1 U15482 ( .A1(n13995), .A2(n13407), .ZN(n13369) );
  NAND2_X1 U15483 ( .A1(n13855), .A2(n13478), .ZN(n13368) );
  NAND2_X1 U15484 ( .A1(n13369), .A2(n13368), .ZN(n13419) );
  OAI22_X1 U15485 ( .A1(n13995), .A2(n6962), .B1(n13827), .B2(n13407), .ZN(
        n13370) );
  XNOR2_X1 U15486 ( .A(n13370), .B(n13476), .ZN(n13418) );
  AND2_X1 U15487 ( .A1(n13478), .A2(n13584), .ZN(n13371) );
  AOI21_X1 U15488 ( .B1(n13852), .B2(n13445), .A(n13371), .ZN(n13417) );
  NAND2_X1 U15489 ( .A1(n13852), .A2(n13475), .ZN(n13373) );
  NAND2_X1 U15490 ( .A1(n13584), .A2(n13445), .ZN(n13372) );
  NAND2_X1 U15491 ( .A1(n13373), .A2(n13372), .ZN(n13374) );
  XNOR2_X1 U15492 ( .A(n13374), .B(n13476), .ZN(n13415) );
  INV_X1 U15493 ( .A(n13415), .ZN(n13416) );
  INV_X1 U15494 ( .A(n13375), .ZN(n13376) );
  NAND2_X1 U15495 ( .A1(n13377), .A2(n13376), .ZN(n13378) );
  NAND2_X1 U15496 ( .A1(n14383), .A2(n13475), .ZN(n13381) );
  OR2_X1 U15497 ( .A1(n13912), .A2(n13407), .ZN(n13380) );
  NAND2_X1 U15498 ( .A1(n13381), .A2(n13380), .ZN(n13382) );
  XNOR2_X1 U15499 ( .A(n13382), .B(n13476), .ZN(n13384) );
  NOR2_X1 U15500 ( .A1(n13912), .A2(n13405), .ZN(n13383) );
  AOI21_X1 U15501 ( .B1(n14383), .B2(n13445), .A(n13383), .ZN(n13385) );
  XNOR2_X1 U15502 ( .A(n13384), .B(n13385), .ZN(n14344) );
  INV_X1 U15503 ( .A(n13384), .ZN(n13386) );
  NAND2_X1 U15504 ( .A1(n13386), .A2(n13385), .ZN(n13387) );
  INV_X1 U15505 ( .A(n13390), .ZN(n13392) );
  OAI22_X1 U15506 ( .A1(n13925), .A2(n6962), .B1(n13899), .B2(n13407), .ZN(
        n13388) );
  XOR2_X1 U15507 ( .A(n13476), .B(n13388), .Z(n13389) );
  INV_X1 U15508 ( .A(n13389), .ZN(n13391) );
  AOI22_X1 U15509 ( .A1(n14375), .A2(n13445), .B1(n13478), .B2(n13586), .ZN(
        n13565) );
  OAI22_X1 U15510 ( .A1(n13515), .A2(n13407), .B1(n13570), .B2(n13405), .ZN(
        n13395) );
  OAI22_X1 U15511 ( .A1(n13515), .A2(n6962), .B1(n13570), .B2(n13407), .ZN(
        n13394) );
  XNOR2_X1 U15512 ( .A(n13394), .B(n13476), .ZN(n13396) );
  XOR2_X1 U15513 ( .A(n13395), .B(n13396), .Z(n13509) );
  OR2_X1 U15514 ( .A1(n13396), .A2(n13395), .ZN(n13397) );
  NAND2_X1 U15515 ( .A1(n14015), .A2(n13475), .ZN(n13399) );
  NAND2_X1 U15516 ( .A1(n13585), .A2(n13445), .ZN(n13398) );
  NAND2_X1 U15517 ( .A1(n13399), .A2(n13398), .ZN(n13400) );
  XNOR2_X1 U15518 ( .A(n13400), .B(n13476), .ZN(n13403) );
  AOI22_X1 U15519 ( .A1(n14015), .A2(n13445), .B1(n13478), .B2(n13585), .ZN(
        n13401) );
  XNOR2_X1 U15520 ( .A(n13403), .B(n13401), .ZN(n13518) );
  INV_X1 U15521 ( .A(n13401), .ZN(n13402) );
  OR2_X1 U15522 ( .A1(n13403), .A2(n13402), .ZN(n13404) );
  OAI22_X1 U15523 ( .A1(n13878), .A2(n13407), .B1(n13406), .B2(n13405), .ZN(
        n13411) );
  NAND2_X1 U15524 ( .A1(n14009), .A2(n13475), .ZN(n13409) );
  NAND2_X1 U15525 ( .A1(n13853), .A2(n13445), .ZN(n13408) );
  NAND2_X1 U15526 ( .A1(n13409), .A2(n13408), .ZN(n13410) );
  XNOR2_X1 U15527 ( .A(n13410), .B(n13476), .ZN(n13412) );
  XOR2_X1 U15528 ( .A(n13411), .B(n13412), .Z(n13551) );
  INV_X1 U15529 ( .A(n13411), .ZN(n13414) );
  INV_X1 U15530 ( .A(n13412), .ZN(n13413) );
  XNOR2_X1 U15531 ( .A(n13415), .B(n13417), .ZN(n13465) );
  OAI21_X1 U15532 ( .B1(n13417), .B2(n13416), .A(n13464), .ZN(n13531) );
  XOR2_X1 U15533 ( .A(n13419), .B(n13418), .Z(n13530) );
  XOR2_X1 U15534 ( .A(n13421), .B(n13420), .Z(n13490) );
  XOR2_X1 U15535 ( .A(n13425), .B(n13424), .Z(n13542) );
  NAND2_X1 U15536 ( .A1(n13979), .A2(n13475), .ZN(n13427) );
  NAND2_X1 U15537 ( .A1(n13582), .A2(n13445), .ZN(n13426) );
  NAND2_X1 U15538 ( .A1(n13427), .A2(n13426), .ZN(n13428) );
  XNOR2_X1 U15539 ( .A(n13428), .B(n13476), .ZN(n13429) );
  AOI22_X1 U15540 ( .A1(n13979), .A2(n13445), .B1(n13478), .B2(n13582), .ZN(
        n13430) );
  XNOR2_X1 U15541 ( .A(n13429), .B(n13430), .ZN(n13458) );
  INV_X1 U15542 ( .A(n13429), .ZN(n13431) );
  AOI22_X1 U15543 ( .A1(n13973), .A2(n13445), .B1(n13478), .B2(n13581), .ZN(
        n13435) );
  NAND2_X1 U15544 ( .A1(n13973), .A2(n13475), .ZN(n13433) );
  NAND2_X1 U15545 ( .A1(n13581), .A2(n13445), .ZN(n13432) );
  NAND2_X1 U15546 ( .A1(n13433), .A2(n13432), .ZN(n13434) );
  XNOR2_X1 U15547 ( .A(n13434), .B(n13476), .ZN(n13437) );
  XOR2_X1 U15548 ( .A(n13435), .B(n13437), .Z(n13524) );
  INV_X1 U15549 ( .A(n13435), .ZN(n13436) );
  NAND2_X1 U15550 ( .A1(n13965), .A2(n13475), .ZN(n13439) );
  NAND2_X1 U15551 ( .A1(n13736), .A2(n13445), .ZN(n13438) );
  NAND2_X1 U15552 ( .A1(n13439), .A2(n13438), .ZN(n13440) );
  XNOR2_X1 U15553 ( .A(n13440), .B(n13476), .ZN(n13443) );
  AOI22_X1 U15554 ( .A1(n13965), .A2(n13445), .B1(n13478), .B2(n13736), .ZN(
        n13441) );
  XNOR2_X1 U15555 ( .A(n13443), .B(n13441), .ZN(n13499) );
  INV_X1 U15556 ( .A(n13441), .ZN(n13442) );
  OR2_X1 U15557 ( .A1(n13443), .A2(n13442), .ZN(n13444) );
  NAND2_X1 U15558 ( .A1(n13957), .A2(n13475), .ZN(n13447) );
  NAND2_X1 U15559 ( .A1(n13580), .A2(n13445), .ZN(n13446) );
  NAND2_X1 U15560 ( .A1(n13447), .A2(n13446), .ZN(n13448) );
  XNOR2_X1 U15561 ( .A(n13448), .B(n13476), .ZN(n13449) );
  AOI22_X1 U15562 ( .A1(n13957), .A2(n13445), .B1(n13478), .B2(n13580), .ZN(
        n13450) );
  XNOR2_X1 U15563 ( .A(n13449), .B(n13450), .ZN(n13557) );
  INV_X1 U15564 ( .A(n13449), .ZN(n13451) );
  INV_X1 U15565 ( .A(n13579), .ZN(n13720) );
  NAND2_X1 U15566 ( .A1(n13573), .A2(n13723), .ZN(n13453) );
  AOI22_X1 U15567 ( .A1(n13568), .A2(n13580), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13452) );
  OAI211_X1 U15568 ( .C1(n13720), .C2(n13571), .A(n13453), .B(n13452), .ZN(
        n13454) );
  AOI21_X1 U15569 ( .B1(n13951), .B2(n14358), .A(n13454), .ZN(n13455) );
  OAI21_X1 U15570 ( .B1(n13456), .B2(n13564), .A(n13455), .ZN(P1_U3214) );
  XOR2_X1 U15571 ( .A(n13458), .B(n13457), .Z(n13463) );
  NAND2_X1 U15572 ( .A1(n13573), .A2(n13791), .ZN(n13460) );
  AOI22_X1 U15573 ( .A1(n13568), .A2(n13825), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13459) );
  OAI211_X1 U15574 ( .C1(n13789), .C2(n13571), .A(n13460), .B(n13459), .ZN(
        n13461) );
  AOI21_X1 U15575 ( .B1(n13979), .B2(n14358), .A(n13461), .ZN(n13462) );
  OAI21_X1 U15576 ( .B1(n13463), .B2(n13564), .A(n13462), .ZN(P1_U3216) );
  INV_X1 U15577 ( .A(n13852), .ZN(n14001) );
  OAI211_X1 U15578 ( .C1(n13466), .C2(n13465), .A(n13464), .B(n14350), .ZN(
        n13470) );
  NAND2_X1 U15579 ( .A1(n13568), .A2(n13853), .ZN(n13467) );
  NAND2_X1 U15580 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13688)
         );
  OAI211_X1 U15581 ( .C1(n13571), .C2(n13827), .A(n13467), .B(n13688), .ZN(
        n13468) );
  AOI21_X1 U15582 ( .B1(n13573), .B2(n13856), .A(n13468), .ZN(n13469) );
  OAI211_X1 U15583 ( .C1(n14001), .C2(n13576), .A(n13470), .B(n13469), .ZN(
        P1_U3219) );
  INV_X1 U15584 ( .A(n13471), .ZN(n13472) );
  AOI22_X1 U15585 ( .A1(n13943), .A2(n13475), .B1(n13445), .B2(n13579), .ZN(
        n13477) );
  XNOR2_X1 U15586 ( .A(n13477), .B(n13476), .ZN(n13480) );
  AOI22_X1 U15587 ( .A1(n13943), .A2(n13445), .B1(n13478), .B2(n13579), .ZN(
        n13479) );
  XNOR2_X1 U15588 ( .A(n13480), .B(n13479), .ZN(n13481) );
  XNOR2_X1 U15589 ( .A(n13482), .B(n13481), .ZN(n13487) );
  NAND2_X1 U15590 ( .A1(n13573), .A2(n13710), .ZN(n13484) );
  AOI22_X1 U15591 ( .A1(n13568), .A2(n13737), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13483) );
  OAI211_X1 U15592 ( .C1(n13705), .C2(n13571), .A(n13484), .B(n13483), .ZN(
        n13485) );
  AOI21_X1 U15593 ( .B1(n13943), .B2(n14358), .A(n13485), .ZN(n13486) );
  OAI21_X1 U15594 ( .B1(n13487), .B2(n13564), .A(n13486), .ZN(P1_U3220) );
  OAI21_X1 U15595 ( .B1(n13490), .B2(n13489), .A(n13488), .ZN(n13491) );
  NAND2_X1 U15596 ( .A1(n13491), .A2(n14350), .ZN(n13497) );
  OAI22_X1 U15597 ( .A1(n13571), .A2(n13790), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13492), .ZN(n13495) );
  NOR2_X1 U15598 ( .A1(n13493), .A2(n13827), .ZN(n13494) );
  AOI211_X1 U15599 ( .C1(n13819), .C2(n13573), .A(n13495), .B(n13494), .ZN(
        n13496) );
  OAI211_X1 U15600 ( .C1(n13821), .C2(n13576), .A(n13497), .B(n13496), .ZN(
        P1_U3223) );
  XOR2_X1 U15601 ( .A(n13499), .B(n13498), .Z(n13506) );
  NAND2_X1 U15602 ( .A1(n13581), .A2(n13854), .ZN(n13501) );
  NAND2_X1 U15603 ( .A1(n13580), .A2(n13913), .ZN(n13500) );
  AND2_X1 U15604 ( .A1(n13501), .A2(n13500), .ZN(n13754) );
  OAI22_X1 U15605 ( .A1(n13754), .A2(n13546), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13502), .ZN(n13503) );
  AOI21_X1 U15606 ( .B1(n13573), .B2(n13760), .A(n13503), .ZN(n13505) );
  NAND2_X1 U15607 ( .A1(n13965), .A2(n14358), .ZN(n13504) );
  OAI211_X1 U15608 ( .C1(n13506), .C2(n13564), .A(n13505), .B(n13504), .ZN(
        P1_U3225) );
  OAI21_X1 U15609 ( .B1(n13509), .B2(n13508), .A(n13507), .ZN(n13510) );
  NAND2_X1 U15610 ( .A1(n13510), .A2(n14350), .ZN(n13514) );
  NAND2_X1 U15611 ( .A1(n13568), .A2(n13586), .ZN(n13511) );
  NAND2_X1 U15612 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14495)
         );
  OAI211_X1 U15613 ( .C1(n13571), .C2(n13898), .A(n13511), .B(n14495), .ZN(
        n13512) );
  AOI21_X1 U15614 ( .B1(n13573), .B2(n13900), .A(n13512), .ZN(n13513) );
  OAI211_X1 U15615 ( .C1(n13515), .C2(n13576), .A(n13514), .B(n13513), .ZN(
        P1_U3226) );
  OAI21_X1 U15616 ( .B1(n13518), .B2(n13517), .A(n13516), .ZN(n13519) );
  NAND2_X1 U15617 ( .A1(n13519), .A2(n14350), .ZN(n13522) );
  AOI22_X1 U15618 ( .A1(n13913), .A2(n13853), .B1(n13914), .B2(n13854), .ZN(
        n13886) );
  NAND2_X1 U15619 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14510)
         );
  OAI21_X1 U15620 ( .B1(n13886), .B2(n13546), .A(n14510), .ZN(n13520) );
  AOI21_X1 U15621 ( .B1(n13573), .B2(n13890), .A(n13520), .ZN(n13521) );
  OAI211_X1 U15622 ( .C1(n13893), .C2(n13576), .A(n13522), .B(n13521), .ZN(
        P1_U3228) );
  XOR2_X1 U15623 ( .A(n13524), .B(n13523), .Z(n13529) );
  AOI22_X1 U15624 ( .A1(n13913), .A2(n13736), .B1(n13582), .B2(n13854), .ZN(
        n13777) );
  OAI22_X1 U15625 ( .A1(n13777), .A2(n13546), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13525), .ZN(n13526) );
  AOI21_X1 U15626 ( .B1(n13573), .B2(n13778), .A(n13526), .ZN(n13528) );
  NAND2_X1 U15627 ( .A1(n13973), .A2(n14358), .ZN(n13527) );
  OAI211_X1 U15628 ( .C1(n13529), .C2(n13564), .A(n13528), .B(n13527), .ZN(
        P1_U3229) );
  OAI21_X1 U15629 ( .B1(n13531), .B2(n13530), .A(n14350), .ZN(n13539) );
  NAND2_X1 U15630 ( .A1(n13584), .A2(n13854), .ZN(n13533) );
  NAND2_X1 U15631 ( .A1(n13583), .A2(n13913), .ZN(n13532) );
  NAND2_X1 U15632 ( .A1(n13533), .A2(n13532), .ZN(n13834) );
  AOI22_X1 U15633 ( .A1(n13834), .A2(n14359), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13534) );
  OAI21_X1 U15634 ( .B1(n14365), .B2(n13842), .A(n13534), .ZN(n13535) );
  AOI21_X1 U15635 ( .B1(n13536), .B2(n14358), .A(n13535), .ZN(n13537) );
  OAI21_X1 U15636 ( .B1(n13539), .B2(n13538), .A(n13537), .ZN(P1_U3233) );
  OAI21_X1 U15637 ( .B1(n13542), .B2(n13541), .A(n13540), .ZN(n13543) );
  NAND2_X1 U15638 ( .A1(n13543), .A2(n14350), .ZN(n13549) );
  NAND2_X1 U15639 ( .A1(n13583), .A2(n13854), .ZN(n13545) );
  NAND2_X1 U15640 ( .A1(n13582), .A2(n13913), .ZN(n13544) );
  AND2_X1 U15641 ( .A1(n13545), .A2(n13544), .ZN(n13804) );
  INV_X1 U15642 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n15476) );
  OAI22_X1 U15643 ( .A1(n13804), .A2(n13546), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15476), .ZN(n13547) );
  AOI21_X1 U15644 ( .B1(n13573), .B2(n13806), .A(n13547), .ZN(n13548) );
  OAI211_X1 U15645 ( .C1(n13576), .C2(n13983), .A(n13549), .B(n13548), .ZN(
        P1_U3235) );
  XOR2_X1 U15646 ( .A(n13551), .B(n13550), .Z(n13556) );
  NAND2_X1 U15647 ( .A1(n13568), .A2(n13585), .ZN(n13552) );
  NAND2_X1 U15648 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14527)
         );
  OAI211_X1 U15649 ( .C1(n13571), .C2(n13872), .A(n13552), .B(n14527), .ZN(
        n13554) );
  NOR2_X1 U15650 ( .A1(n13878), .A2(n13576), .ZN(n13553) );
  AOI211_X1 U15651 ( .C1(n13876), .C2(n13573), .A(n13554), .B(n13553), .ZN(
        n13555) );
  OAI21_X1 U15652 ( .B1(n13556), .B2(n13564), .A(n13555), .ZN(P1_U3238) );
  NAND2_X1 U15653 ( .A1(n13573), .A2(n13740), .ZN(n13559) );
  AOI22_X1 U15654 ( .A1(n13568), .A2(n13736), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13558) );
  OAI211_X1 U15655 ( .C1(n13704), .C2(n13571), .A(n13559), .B(n13558), .ZN(
        n13560) );
  AOI21_X1 U15656 ( .B1(n13957), .B2(n14358), .A(n13560), .ZN(n13561) );
  OAI21_X1 U15657 ( .B1(n13562), .B2(n13564), .A(n13561), .ZN(P1_U3240) );
  AOI211_X1 U15658 ( .C1(n13566), .C2(n13565), .A(n13564), .B(n13563), .ZN(
        n13567) );
  INV_X1 U15659 ( .A(n13567), .ZN(n13575) );
  NAND2_X1 U15660 ( .A1(n13568), .A2(n13587), .ZN(n13569) );
  NAND2_X1 U15661 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14480)
         );
  OAI211_X1 U15662 ( .C1(n13571), .C2(n13570), .A(n13569), .B(n14480), .ZN(
        n13572) );
  AOI21_X1 U15663 ( .B1(n13573), .B2(n13921), .A(n13572), .ZN(n13574) );
  OAI211_X1 U15664 ( .C1(n13925), .C2(n13576), .A(n13575), .B(n13574), .ZN(
        P1_U3241) );
  MUX2_X1 U15665 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n13694), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U15666 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n13577), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U15667 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13578), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U15668 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n13579), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U15669 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n13737), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15670 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n13580), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15671 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n13736), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15672 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n13581), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15673 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n13582), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U15674 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n13825), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U15675 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n13583), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U15676 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n13855), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U15677 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n13584), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U15678 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n13853), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U15679 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n13585), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U15680 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n13914), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U15681 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n13586), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U15682 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n13587), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U15683 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n13588), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U15684 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n13589), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U15685 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n13590), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U15686 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n13591), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U15687 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n13592), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U15688 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n13593), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U15689 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n13594), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U15690 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n13595), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U15691 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n13596), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U15692 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n10867), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U15693 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n13597), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U15694 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n13598), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U15695 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n13599), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U15696 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n10017), .S(P1_U4016), .Z(
        P1_U3560) );
  OAI22_X1 U15697 ( .A1(n14529), .A2(n7545), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13600), .ZN(n13601) );
  AOI21_X1 U15698 ( .B1(n14494), .B2(n13602), .A(n13601), .ZN(n13610) );
  OAI211_X1 U15699 ( .C1(n13605), .C2(n13604), .A(n14517), .B(n13603), .ZN(
        n13609) );
  OAI211_X1 U15700 ( .C1(n13607), .C2(n13613), .A(n14521), .B(n13606), .ZN(
        n13608) );
  NAND3_X1 U15701 ( .A1(n13610), .A2(n13609), .A3(n13608), .ZN(P1_U3244) );
  MUX2_X1 U15702 ( .A(n13613), .B(n13612), .S(n6641), .Z(n13615) );
  NAND2_X1 U15703 ( .A1(n13615), .A2(n13614), .ZN(n13616) );
  OAI211_X1 U15704 ( .C1(n14044), .C2(n13617), .A(n13616), .B(P1_U4016), .ZN(
        n13655) );
  INV_X1 U15705 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n13618) );
  OAI22_X1 U15706 ( .A1(n14529), .A2(n7012), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13618), .ZN(n13619) );
  AOI21_X1 U15707 ( .B1(n14494), .B2(n13620), .A(n13619), .ZN(n13629) );
  OAI211_X1 U15708 ( .C1(n13623), .C2(n13622), .A(n14521), .B(n13621), .ZN(
        n13628) );
  OAI211_X1 U15709 ( .C1(n13626), .C2(n13625), .A(n14517), .B(n13624), .ZN(
        n13627) );
  NAND4_X1 U15710 ( .A1(n13655), .A2(n13629), .A3(n13628), .A4(n13627), .ZN(
        P1_U3245) );
  NAND2_X1 U15711 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n13631) );
  OAI21_X1 U15712 ( .B1(n14529), .B2(n14049), .A(n13631), .ZN(n13632) );
  AOI21_X1 U15713 ( .B1(n14494), .B2(n7286), .A(n13632), .ZN(n13641) );
  OAI211_X1 U15714 ( .C1(n13635), .C2(n13634), .A(n14521), .B(n13633), .ZN(
        n13640) );
  OAI211_X1 U15715 ( .C1(n13638), .C2(n13637), .A(n14517), .B(n13636), .ZN(
        n13639) );
  NAND3_X1 U15716 ( .A1(n13641), .A2(n13640), .A3(n13639), .ZN(P1_U3246) );
  INV_X1 U15717 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n13643) );
  OAI21_X1 U15718 ( .B1(n14529), .B2(n13643), .A(n13642), .ZN(n13644) );
  AOI21_X1 U15719 ( .B1(n14494), .B2(n13645), .A(n13644), .ZN(n13654) );
  OAI211_X1 U15720 ( .C1(n13648), .C2(n13647), .A(n14517), .B(n13646), .ZN(
        n13653) );
  OAI211_X1 U15721 ( .C1(n13651), .C2(n13650), .A(n14521), .B(n13649), .ZN(
        n13652) );
  NAND4_X1 U15722 ( .A1(n13655), .A2(n13654), .A3(n13653), .A4(n13652), .ZN(
        P1_U3247) );
  INV_X1 U15723 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n15332) );
  NOR2_X1 U15724 ( .A1(n14493), .A2(n15332), .ZN(n13656) );
  AOI21_X1 U15725 ( .B1(n15332), .B2(n14493), .A(n13656), .ZN(n14489) );
  INV_X1 U15726 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n13657) );
  MUX2_X1 U15727 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n13657), .S(n14449), .Z(
        n13658) );
  INV_X1 U15728 ( .A(n13658), .ZN(n14445) );
  OAI21_X1 U15729 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n13671), .A(n13659), 
        .ZN(n14446) );
  NOR2_X1 U15730 ( .A1(n14445), .A2(n14446), .ZN(n14444) );
  INV_X1 U15731 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n13660) );
  MUX2_X1 U15732 ( .A(n13660), .B(P1_REG2_REG_14__SCAN_IN), .S(n14453), .Z(
        n14460) );
  NAND2_X1 U15733 ( .A1(n13661), .A2(n14478), .ZN(n13663) );
  XNOR2_X1 U15734 ( .A(n14478), .B(n13662), .ZN(n14474) );
  INV_X1 U15735 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n14473) );
  NAND2_X1 U15736 ( .A1(n14474), .A2(n14473), .ZN(n14472) );
  NAND2_X1 U15737 ( .A1(n13663), .A2(n14472), .ZN(n14490) );
  INV_X1 U15738 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n13664) );
  MUX2_X1 U15739 ( .A(n13664), .B(P1_REG2_REG_17__SCAN_IN), .S(n13676), .Z(
        n14504) );
  NOR2_X1 U15740 ( .A1(n13665), .A2(n14524), .ZN(n13666) );
  INV_X1 U15741 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n15327) );
  XNOR2_X1 U15742 ( .A(n14524), .B(n13665), .ZN(n14519) );
  NOR2_X1 U15743 ( .A1(n15327), .A2(n14519), .ZN(n14518) );
  NOR2_X1 U15744 ( .A1(n13666), .A2(n14518), .ZN(n13667) );
  XNOR2_X1 U15745 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n13667), .ZN(n13684) );
  INV_X1 U15746 ( .A(n13684), .ZN(n13682) );
  INV_X1 U15747 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n14514) );
  INV_X1 U15748 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n14373) );
  NOR2_X1 U15749 ( .A1(n14493), .A2(n14373), .ZN(n13668) );
  AOI21_X1 U15750 ( .B1(n14493), .B2(n14373), .A(n13668), .ZN(n14485) );
  INV_X1 U15751 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n13669) );
  MUX2_X1 U15752 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n13669), .S(n14453), .Z(
        n14456) );
  OAI21_X1 U15753 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n13671), .A(n13670), 
        .ZN(n14443) );
  INV_X1 U15754 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n13672) );
  MUX2_X1 U15755 ( .A(n13672), .B(P1_REG1_REG_13__SCAN_IN), .S(n14449), .Z(
        n14442) );
  NOR2_X1 U15756 ( .A1(n14443), .A2(n14442), .ZN(n14441) );
  NAND2_X1 U15757 ( .A1(n14456), .A2(n14455), .ZN(n14454) );
  OAI21_X1 U15758 ( .B1(n14453), .B2(P1_REG1_REG_14__SCAN_IN), .A(n14454), 
        .ZN(n13673) );
  NAND2_X1 U15759 ( .A1(n14478), .A2(n13673), .ZN(n13675) );
  INV_X1 U15760 ( .A(n13673), .ZN(n13674) );
  INV_X1 U15761 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n15488) );
  NAND2_X1 U15762 ( .A1(n14470), .A2(n15488), .ZN(n14469) );
  NAND2_X1 U15763 ( .A1(n13675), .A2(n14469), .ZN(n14486) );
  NOR2_X1 U15764 ( .A1(n14485), .A2(n14486), .ZN(n14484) );
  XNOR2_X1 U15765 ( .A(n13676), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n14500) );
  NOR2_X1 U15766 ( .A1(n14499), .A2(n14500), .ZN(n14498) );
  XNOR2_X1 U15767 ( .A(n14524), .B(n13677), .ZN(n14515) );
  NOR2_X1 U15768 ( .A1(n14514), .A2(n14515), .ZN(n14513) );
  NOR2_X1 U15769 ( .A1(n13677), .A2(n14524), .ZN(n13678) );
  NOR2_X1 U15770 ( .A1(n14513), .A2(n13678), .ZN(n13680) );
  INV_X1 U15771 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n13679) );
  XOR2_X1 U15772 ( .A(n13680), .B(n13679), .Z(n13683) );
  OAI21_X1 U15773 ( .B1(n13683), .B2(n14483), .A(n14525), .ZN(n13681) );
  AOI21_X1 U15774 ( .B1(n13682), .B2(n14521), .A(n13681), .ZN(n13687) );
  AOI22_X1 U15775 ( .A1(n13684), .A2(n14521), .B1(n14517), .B2(n13683), .ZN(
        n13686) );
  MUX2_X1 U15776 ( .A(n13687), .B(n13686), .S(n13685), .Z(n13689) );
  OAI211_X1 U15777 ( .C1(n7718), .C2(n14529), .A(n13689), .B(n13688), .ZN(
        P1_U3262) );
  NOR2_X1 U15778 ( .A1(n13690), .A2(n13698), .ZN(n13691) );
  XNOR2_X1 U15779 ( .A(n13691), .B(n13695), .ZN(n13692) );
  NAND2_X1 U15780 ( .A1(n13692), .A2(n14561), .ZN(n13932) );
  NAND2_X1 U15781 ( .A1(n13694), .A2(n13693), .ZN(n13933) );
  NOR2_X1 U15782 ( .A1(n14570), .A2(n13933), .ZN(n13701) );
  NOR2_X1 U15783 ( .A1(n6998), .A2(n14573), .ZN(n13696) );
  AOI211_X1 U15784 ( .C1(n14570), .C2(P1_REG2_REG_31__SCAN_IN), .A(n13701), 
        .B(n13696), .ZN(n13697) );
  OAI21_X1 U15785 ( .B1(n13932), .B2(n13927), .A(n13697), .ZN(P1_U3263) );
  XNOR2_X1 U15786 ( .A(n13935), .B(n13698), .ZN(n13699) );
  NAND2_X1 U15787 ( .A1(n13699), .A2(n14561), .ZN(n13934) );
  NOR2_X1 U15788 ( .A1(n13935), .A2(n14573), .ZN(n13700) );
  AOI211_X1 U15789 ( .C1(n14570), .C2(P1_REG2_REG_30__SCAN_IN), .A(n13701), 
        .B(n13700), .ZN(n13702) );
  OAI21_X1 U15790 ( .B1(n13927), .B2(n13934), .A(n13702), .ZN(P1_U3264) );
  XNOR2_X1 U15791 ( .A(n13703), .B(n13714), .ZN(n13707) );
  OAI22_X1 U15792 ( .A1(n13705), .A2(n14539), .B1(n13704), .B2(n14537), .ZN(
        n13706) );
  OAI211_X1 U15793 ( .C1(n13709), .C2(n6676), .A(n14561), .B(n13708), .ZN(
        n13946) );
  AOI22_X1 U15794 ( .A1(n14570), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n13710), 
        .B2(n14569), .ZN(n13712) );
  NAND2_X1 U15795 ( .A1(n13943), .A2(n14557), .ZN(n13711) );
  OAI211_X1 U15796 ( .C1(n13946), .C2(n13927), .A(n13712), .B(n13711), .ZN(
        n13713) );
  INV_X1 U15797 ( .A(n13713), .ZN(n13717) );
  NAND2_X1 U15798 ( .A1(n13715), .A2(n13714), .ZN(n13944) );
  NAND3_X1 U15799 ( .A1(n13945), .A2(n13944), .A3(n14175), .ZN(n13716) );
  OAI211_X1 U15800 ( .C1(n13949), .C2(n13930), .A(n13717), .B(n13716), .ZN(
        P1_U3265) );
  OAI21_X1 U15801 ( .B1(n6708), .B2(n13728), .A(n13718), .ZN(n13722) );
  OAI22_X1 U15802 ( .A1(n13720), .A2(n14539), .B1(n13719), .B2(n14537), .ZN(
        n13721) );
  AOI21_X1 U15803 ( .B1(n13722), .B2(n14554), .A(n13721), .ZN(n13953) );
  AOI211_X1 U15804 ( .C1(n13951), .C2(n13735), .A(n13903), .B(n6676), .ZN(
        n13950) );
  INV_X1 U15805 ( .A(n13951), .ZN(n13725) );
  AOI22_X1 U15806 ( .A1(n13930), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n13723), 
        .B2(n14569), .ZN(n13724) );
  OAI21_X1 U15807 ( .B1(n13725), .B2(n14573), .A(n13724), .ZN(n13729) );
  AOI211_X1 U15808 ( .C1(n13950), .C2(n14567), .A(n13729), .B(n6667), .ZN(
        n13730) );
  OAI21_X1 U15809 ( .B1(n13953), .B2(n13930), .A(n13730), .ZN(P1_U3266) );
  XNOR2_X1 U15810 ( .A(n13732), .B(n13731), .ZN(n13955) );
  INV_X1 U15811 ( .A(n13955), .ZN(n13750) );
  INV_X1 U15812 ( .A(n13759), .ZN(n13733) );
  AOI21_X1 U15813 ( .B1(n13957), .B2(n13733), .A(n13903), .ZN(n13734) );
  NAND2_X1 U15814 ( .A1(n13735), .A2(n13734), .ZN(n13960) );
  INV_X1 U15815 ( .A(n13960), .ZN(n13745) );
  NAND2_X1 U15816 ( .A1(n13736), .A2(n13854), .ZN(n13739) );
  NAND2_X1 U15817 ( .A1(n13737), .A2(n13913), .ZN(n13738) );
  NAND2_X1 U15818 ( .A1(n13739), .A2(n13738), .ZN(n13956) );
  AOI22_X1 U15819 ( .A1(n13902), .A2(n13956), .B1(n13740), .B2(n14569), .ZN(
        n13742) );
  NAND2_X1 U15820 ( .A1(n14570), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n13741) );
  OAI211_X1 U15821 ( .C1(n13743), .C2(n14573), .A(n13742), .B(n13741), .ZN(
        n13744) );
  AOI21_X1 U15822 ( .B1(n13745), .B2(n14567), .A(n13744), .ZN(n13749) );
  OR2_X1 U15823 ( .A1(n13747), .A2(n13746), .ZN(n13959) );
  NAND3_X1 U15824 ( .A1(n13959), .A2(n13958), .A3(n14175), .ZN(n13748) );
  OAI211_X1 U15825 ( .C1(n13750), .C2(n13911), .A(n13749), .B(n13748), .ZN(
        P1_U3267) );
  INV_X1 U15826 ( .A(n13751), .ZN(n13753) );
  OAI21_X1 U15827 ( .B1(n13753), .B2(n13765), .A(n13752), .ZN(n13756) );
  INV_X1 U15828 ( .A(n13754), .ZN(n13755) );
  AOI21_X1 U15829 ( .B1(n13756), .B2(n14554), .A(n13755), .ZN(n13969) );
  NAND2_X1 U15830 ( .A1(n13776), .A2(n13965), .ZN(n13757) );
  NAND2_X1 U15831 ( .A1(n13757), .A2(n14561), .ZN(n13758) );
  NOR2_X1 U15832 ( .A1(n13759), .A2(n13758), .ZN(n13964) );
  NAND2_X1 U15833 ( .A1(n13965), .A2(n14557), .ZN(n13762) );
  AOI22_X1 U15834 ( .A1(n14570), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n13760), 
        .B2(n14569), .ZN(n13761) );
  NAND2_X1 U15835 ( .A1(n13762), .A2(n13761), .ZN(n13763) );
  AOI21_X1 U15836 ( .B1(n13964), .B2(n14567), .A(n13763), .ZN(n13768) );
  NAND2_X1 U15837 ( .A1(n13766), .A2(n13765), .ZN(n13966) );
  NAND3_X1 U15838 ( .A1(n13764), .A2(n13966), .A3(n14175), .ZN(n13767) );
  OAI211_X1 U15839 ( .C1(n13969), .C2(n13930), .A(n13768), .B(n13767), .ZN(
        P1_U3268) );
  XNOR2_X1 U15840 ( .A(n13769), .B(n13770), .ZN(n13976) );
  NAND2_X1 U15841 ( .A1(n13773), .A2(n13772), .ZN(n13970) );
  NAND3_X1 U15842 ( .A1(n13771), .A2(n13970), .A3(n13863), .ZN(n13784) );
  AOI21_X1 U15843 ( .B1(n13774), .B2(n13973), .A(n13903), .ZN(n13775) );
  AND2_X1 U15844 ( .A1(n13776), .A2(n13775), .ZN(n13971) );
  INV_X1 U15845 ( .A(n13777), .ZN(n13972) );
  AOI22_X1 U15846 ( .A1(n13902), .A2(n13972), .B1(n13778), .B2(n14569), .ZN(
        n13780) );
  NAND2_X1 U15847 ( .A1(n14570), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n13779) );
  OAI211_X1 U15848 ( .C1(n13781), .C2(n14573), .A(n13780), .B(n13779), .ZN(
        n13782) );
  AOI21_X1 U15849 ( .B1(n13971), .B2(n14567), .A(n13782), .ZN(n13783) );
  OAI211_X1 U15850 ( .C1(n13785), .C2(n13976), .A(n13784), .B(n13783), .ZN(
        P1_U3269) );
  XNOR2_X1 U15851 ( .A(n13787), .B(n13786), .ZN(n13788) );
  OAI222_X1 U15852 ( .A1(n14537), .A2(n13790), .B1(n14539), .B2(n13789), .C1(
        n14666), .C2(n13788), .ZN(n13977) );
  AOI21_X1 U15853 ( .B1(n13791), .B2(n14569), .A(n13977), .ZN(n13800) );
  AOI211_X1 U15854 ( .C1(n13979), .C2(n13810), .A(n13903), .B(n13792), .ZN(
        n13978) );
  INV_X1 U15855 ( .A(n13979), .ZN(n13794) );
  INV_X1 U15856 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n13793) );
  OAI22_X1 U15857 ( .A1(n13794), .A2(n14573), .B1(n13793), .B2(n13902), .ZN(
        n13798) );
  XNOR2_X1 U15858 ( .A(n13796), .B(n13795), .ZN(n13981) );
  NOR2_X1 U15859 ( .A1(n13981), .A2(n13896), .ZN(n13797) );
  AOI211_X1 U15860 ( .C1(n13978), .C2(n14567), .A(n13798), .B(n13797), .ZN(
        n13799) );
  OAI21_X1 U15861 ( .B1(n13800), .B2(n13930), .A(n13799), .ZN(P1_U3270) );
  INV_X1 U15862 ( .A(n13801), .ZN(n13802) );
  AOI21_X1 U15863 ( .B1(n13808), .B2(n13803), .A(n13802), .ZN(n13805) );
  OAI21_X1 U15864 ( .B1(n13805), .B2(n14666), .A(n13804), .ZN(n13984) );
  AOI21_X1 U15865 ( .B1(n13806), .B2(n14569), .A(n13984), .ZN(n13816) );
  OAI21_X1 U15866 ( .B1(n13809), .B2(n13808), .A(n13807), .ZN(n13986) );
  AOI21_X1 U15867 ( .B1(n13812), .B2(n13818), .A(n13903), .ZN(n13811) );
  NAND2_X1 U15868 ( .A1(n13811), .A2(n13810), .ZN(n13982) );
  AOI22_X1 U15869 ( .A1(n13812), .A2(n14557), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n13930), .ZN(n13813) );
  OAI21_X1 U15870 ( .B1(n13982), .B2(n13927), .A(n13813), .ZN(n13814) );
  AOI21_X1 U15871 ( .B1(n13986), .B2(n14175), .A(n13814), .ZN(n13815) );
  OAI21_X1 U15872 ( .B1(n13816), .B2(n13930), .A(n13815), .ZN(P1_U3271) );
  XOR2_X1 U15873 ( .A(n13817), .B(n13823), .Z(n13993) );
  AOI211_X1 U15874 ( .C1(n13990), .C2(n13841), .A(n13903), .B(n7296), .ZN(
        n13988) );
  AOI22_X1 U15875 ( .A1(n13930), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n13819), 
        .B2(n14569), .ZN(n13820) );
  OAI21_X1 U15876 ( .B1(n13821), .B2(n14573), .A(n13820), .ZN(n13830) );
  OAI211_X1 U15877 ( .C1(n13824), .C2(n13823), .A(n14554), .B(n13822), .ZN(
        n13992) );
  NAND2_X1 U15878 ( .A1(n13825), .A2(n13913), .ZN(n13826) );
  OAI21_X1 U15879 ( .B1(n13827), .B2(n14537), .A(n13826), .ZN(n13989) );
  INV_X1 U15880 ( .A(n13989), .ZN(n13828) );
  AOI21_X1 U15881 ( .B1(n13992), .B2(n13828), .A(n14570), .ZN(n13829) );
  AOI211_X1 U15882 ( .C1(n13988), .C2(n14567), .A(n13830), .B(n13829), .ZN(
        n13831) );
  OAI21_X1 U15883 ( .B1(n13993), .B2(n13896), .A(n13831), .ZN(P1_U3272) );
  AOI21_X1 U15884 ( .B1(n13833), .B2(n13832), .A(n14666), .ZN(n13836) );
  AOI21_X1 U15885 ( .B1(n13836), .B2(n13835), .A(n13834), .ZN(n13999) );
  INV_X1 U15886 ( .A(n13837), .ZN(n13838) );
  AOI21_X1 U15887 ( .B1(n13840), .B2(n13839), .A(n13838), .ZN(n13997) );
  OAI211_X1 U15888 ( .C1(n13851), .C2(n13995), .A(n14561), .B(n13841), .ZN(
        n13994) );
  NOR2_X1 U15889 ( .A1(n13994), .A2(n13927), .ZN(n13846) );
  INV_X1 U15890 ( .A(n13842), .ZN(n13843) );
  AOI22_X1 U15891 ( .A1(n13930), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n13843), 
        .B2(n14569), .ZN(n13844) );
  OAI21_X1 U15892 ( .B1(n13995), .B2(n14573), .A(n13844), .ZN(n13845) );
  AOI211_X1 U15893 ( .C1(n13997), .C2(n14175), .A(n13846), .B(n13845), .ZN(
        n13847) );
  OAI21_X1 U15894 ( .B1(n13999), .B2(n13930), .A(n13847), .ZN(P1_U3273) );
  XNOR2_X1 U15895 ( .A(n13848), .B(n13850), .ZN(n14006) );
  OAI21_X1 U15896 ( .B1(n6784), .B2(n13850), .A(n13849), .ZN(n14004) );
  AOI211_X1 U15897 ( .C1(n13852), .C2(n13874), .A(n13903), .B(n13851), .ZN(
        n14003) );
  NAND2_X1 U15898 ( .A1(n14003), .A2(n14567), .ZN(n13861) );
  AOI22_X1 U15899 ( .A1(n13855), .A2(n13913), .B1(n13854), .B2(n13853), .ZN(
        n14000) );
  INV_X1 U15900 ( .A(n13856), .ZN(n13858) );
  OAI22_X1 U15901 ( .A1(n14000), .A2(n13930), .B1(n13858), .B2(n13857), .ZN(
        n13859) );
  AOI21_X1 U15902 ( .B1(P1_REG2_REG_19__SCAN_IN), .B2(n14570), .A(n13859), 
        .ZN(n13860) );
  OAI211_X1 U15903 ( .C1(n14001), .C2(n14573), .A(n13861), .B(n13860), .ZN(
        n13862) );
  AOI21_X1 U15904 ( .B1(n14004), .B2(n13863), .A(n13862), .ZN(n13864) );
  OAI21_X1 U15905 ( .B1(n13896), .B2(n14006), .A(n13864), .ZN(P1_U3274) );
  XNOR2_X1 U15906 ( .A(n13865), .B(n13867), .ZN(n13871) );
  INV_X1 U15907 ( .A(n13871), .ZN(n14012) );
  INV_X1 U15908 ( .A(n14577), .ZN(n13882) );
  OAI211_X1 U15909 ( .C1(n13868), .C2(n13867), .A(n13866), .B(n14554), .ZN(
        n13869) );
  OAI21_X1 U15910 ( .B1(n13898), .B2(n14537), .A(n13869), .ZN(n13870) );
  AOI21_X1 U15911 ( .B1(n14639), .B2(n13871), .A(n13870), .ZN(n14011) );
  INV_X1 U15912 ( .A(n14011), .ZN(n13873) );
  NOR2_X1 U15913 ( .A1(n13872), .A2(n14539), .ZN(n14008) );
  OAI21_X1 U15914 ( .B1(n13873), .B2(n14008), .A(n13902), .ZN(n13881) );
  INV_X1 U15915 ( .A(n13874), .ZN(n13875) );
  AOI211_X1 U15916 ( .C1(n14009), .C2(n13888), .A(n13903), .B(n13875), .ZN(
        n14007) );
  AOI22_X1 U15917 ( .A1(n14570), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n13876), 
        .B2(n14569), .ZN(n13877) );
  OAI21_X1 U15918 ( .B1(n13878), .B2(n14573), .A(n13877), .ZN(n13879) );
  AOI21_X1 U15919 ( .B1(n14007), .B2(n14567), .A(n13879), .ZN(n13880) );
  OAI211_X1 U15920 ( .C1(n14012), .C2(n13882), .A(n13881), .B(n13880), .ZN(
        P1_U3275) );
  XNOR2_X1 U15921 ( .A(n13883), .B(n7346), .ZN(n14017) );
  XNOR2_X1 U15922 ( .A(n13885), .B(n7346), .ZN(n13887) );
  OAI21_X1 U15923 ( .B1(n13887), .B2(n14666), .A(n13886), .ZN(n14013) );
  AOI21_X1 U15924 ( .B1(n13904), .B2(n14015), .A(n13903), .ZN(n13889) );
  AND2_X1 U15925 ( .A1(n13889), .A2(n13888), .ZN(n14014) );
  NAND2_X1 U15926 ( .A1(n14014), .A2(n14567), .ZN(n13892) );
  AOI22_X1 U15927 ( .A1(n13930), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n13890), 
        .B2(n14569), .ZN(n13891) );
  OAI211_X1 U15928 ( .C1(n13893), .C2(n14573), .A(n13892), .B(n13891), .ZN(
        n13894) );
  AOI21_X1 U15929 ( .B1(n14013), .B2(n13902), .A(n13894), .ZN(n13895) );
  OAI21_X1 U15930 ( .B1(n14017), .B2(n13896), .A(n13895), .ZN(P1_U3276) );
  AOI21_X1 U15931 ( .B1(n7359), .B2(n13897), .A(n6778), .ZN(n14370) );
  OAI22_X1 U15932 ( .A1(n13899), .A2(n14537), .B1(n13898), .B2(n14539), .ZN(
        n14366) );
  AOI22_X1 U15933 ( .A1(n13902), .A2(n14366), .B1(n13900), .B2(n14569), .ZN(
        n13901) );
  OAI21_X1 U15934 ( .B1(n15332), .B2(n13902), .A(n13901), .ZN(n13907) );
  AOI21_X1 U15935 ( .B1(n13924), .B2(n14367), .A(n13903), .ZN(n13905) );
  NAND2_X1 U15936 ( .A1(n13905), .A2(n13904), .ZN(n14368) );
  NOR2_X1 U15937 ( .A1(n14368), .A2(n13927), .ZN(n13906) );
  AOI211_X1 U15938 ( .C1(n14557), .C2(n14367), .A(n13907), .B(n13906), .ZN(
        n13910) );
  XNOR2_X1 U15939 ( .A(n13908), .B(n7359), .ZN(n14372) );
  NAND2_X1 U15940 ( .A1(n14372), .A2(n14175), .ZN(n13909) );
  OAI211_X1 U15941 ( .C1(n14370), .C2(n13911), .A(n13910), .B(n13909), .ZN(
        P1_U3277) );
  OR2_X1 U15942 ( .A1(n13912), .A2(n14537), .ZN(n13916) );
  NAND2_X1 U15943 ( .A1(n13914), .A2(n13913), .ZN(n13915) );
  NAND2_X1 U15944 ( .A1(n13916), .A2(n13915), .ZN(n14374) );
  OAI211_X1 U15945 ( .C1(n13919), .C2(n13918), .A(n13917), .B(n14554), .ZN(
        n14378) );
  INV_X1 U15946 ( .A(n14378), .ZN(n13920) );
  AOI211_X1 U15947 ( .C1(n14569), .C2(n13921), .A(n14374), .B(n13920), .ZN(
        n13931) );
  OAI21_X1 U15948 ( .B1(n7685), .B2(n13923), .A(n13922), .ZN(n14380) );
  OAI211_X1 U15949 ( .C1(n13925), .C2(n6771), .A(n14561), .B(n13924), .ZN(
        n14376) );
  AOI22_X1 U15950 ( .A1(n14375), .A2(n14557), .B1(n13930), .B2(
        P1_REG2_REG_15__SCAN_IN), .ZN(n13926) );
  OAI21_X1 U15951 ( .B1(n14376), .B2(n13927), .A(n13926), .ZN(n13928) );
  AOI21_X1 U15952 ( .B1(n14380), .B2(n14175), .A(n13928), .ZN(n13929) );
  OAI21_X1 U15953 ( .B1(n13931), .B2(n13930), .A(n13929), .ZN(P1_U3278) );
  OAI211_X1 U15954 ( .C1(n6998), .C2(n14665), .A(n13932), .B(n13933), .ZN(
        n14020) );
  MUX2_X1 U15955 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14020), .S(n14688), .Z(
        P1_U3559) );
  OAI211_X1 U15956 ( .C1(n13935), .C2(n14665), .A(n13934), .B(n13933), .ZN(
        n14021) );
  MUX2_X1 U15957 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14021), .S(n14688), .Z(
        P1_U3558) );
  NAND2_X1 U15958 ( .A1(n13938), .A2(n13937), .ZN(n13940) );
  MUX2_X1 U15959 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14022), .S(n14688), .Z(
        P1_U3557) );
  NAND2_X1 U15960 ( .A1(n13943), .A2(n14632), .ZN(n13948) );
  NAND3_X1 U15961 ( .A1(n13945), .A2(n14671), .A3(n13944), .ZN(n13947) );
  NAND4_X1 U15962 ( .A1(n13949), .A2(n13948), .A3(n13947), .A4(n13946), .ZN(
        n14023) );
  MUX2_X1 U15963 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14023), .S(n14688), .Z(
        P1_U3556) );
  AOI21_X1 U15964 ( .B1(n14632), .B2(n13951), .A(n13950), .ZN(n13952) );
  OAI211_X1 U15965 ( .C1(n14018), .C2(n13954), .A(n13953), .B(n13952), .ZN(
        n14024) );
  MUX2_X1 U15966 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14024), .S(n14688), .Z(
        P1_U3555) );
  NAND2_X1 U15967 ( .A1(n13955), .A2(n14554), .ZN(n13963) );
  AOI21_X1 U15968 ( .B1(n13957), .B2(n14632), .A(n13956), .ZN(n13962) );
  NAND3_X1 U15969 ( .A1(n13959), .A2(n13958), .A3(n14671), .ZN(n13961) );
  NAND4_X1 U15970 ( .A1(n13963), .A2(n13962), .A3(n13961), .A4(n13960), .ZN(
        n14025) );
  MUX2_X1 U15971 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14025), .S(n14688), .Z(
        P1_U3554) );
  AOI21_X1 U15972 ( .B1(n14632), .B2(n13965), .A(n13964), .ZN(n13968) );
  NAND3_X1 U15973 ( .A1(n13764), .A2(n13966), .A3(n14671), .ZN(n13967) );
  NAND3_X1 U15974 ( .A1(n13969), .A2(n13968), .A3(n13967), .ZN(n14026) );
  MUX2_X1 U15975 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14026), .S(n14688), .Z(
        P1_U3553) );
  NAND3_X1 U15976 ( .A1(n13771), .A2(n13970), .A3(n14554), .ZN(n13975) );
  AOI211_X1 U15977 ( .C1(n14632), .C2(n13973), .A(n13972), .B(n13971), .ZN(
        n13974) );
  OAI211_X1 U15978 ( .C1(n14018), .C2(n13976), .A(n13975), .B(n13974), .ZN(
        n14027) );
  MUX2_X1 U15979 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14027), .S(n14688), .Z(
        P1_U3552) );
  AOI211_X1 U15980 ( .C1(n14632), .C2(n13979), .A(n13978), .B(n13977), .ZN(
        n13980) );
  OAI21_X1 U15981 ( .B1(n14018), .B2(n13981), .A(n13980), .ZN(n14028) );
  MUX2_X1 U15982 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14028), .S(n14688), .Z(
        P1_U3551) );
  OAI21_X1 U15983 ( .B1(n14665), .B2(n13983), .A(n13982), .ZN(n13985) );
  AOI211_X1 U15984 ( .C1(n14671), .C2(n13986), .A(n13985), .B(n13984), .ZN(
        n13987) );
  INV_X1 U15985 ( .A(n13987), .ZN(n14029) );
  MUX2_X1 U15986 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14029), .S(n14688), .Z(
        P1_U3550) );
  AOI211_X1 U15987 ( .C1(n14632), .C2(n13990), .A(n13989), .B(n13988), .ZN(
        n13991) );
  OAI211_X1 U15988 ( .C1(n14018), .C2(n13993), .A(n13992), .B(n13991), .ZN(
        n14030) );
  MUX2_X1 U15989 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14030), .S(n14688), .Z(
        P1_U3549) );
  OAI21_X1 U15990 ( .B1(n13995), .B2(n14665), .A(n13994), .ZN(n13996) );
  AOI21_X1 U15991 ( .B1(n13997), .B2(n14671), .A(n13996), .ZN(n13998) );
  NAND2_X1 U15992 ( .A1(n13999), .A2(n13998), .ZN(n14031) );
  MUX2_X1 U15993 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14031), .S(n14688), .Z(
        P1_U3548) );
  OAI21_X1 U15994 ( .B1(n14001), .B2(n14665), .A(n14000), .ZN(n14002) );
  AOI211_X1 U15995 ( .C1(n14004), .C2(n14554), .A(n14003), .B(n14002), .ZN(
        n14005) );
  OAI21_X1 U15996 ( .B1(n14018), .B2(n14006), .A(n14005), .ZN(n14032) );
  MUX2_X1 U15997 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14032), .S(n14688), .Z(
        P1_U3547) );
  AOI211_X1 U15998 ( .C1(n14632), .C2(n14009), .A(n14008), .B(n14007), .ZN(
        n14010) );
  OAI211_X1 U15999 ( .C1(n14012), .C2(n14636), .A(n14011), .B(n14010), .ZN(
        n14033) );
  MUX2_X1 U16000 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14033), .S(n14688), .Z(
        P1_U3546) );
  AOI211_X1 U16001 ( .C1(n14632), .C2(n14015), .A(n14014), .B(n14013), .ZN(
        n14016) );
  OAI21_X1 U16002 ( .B1(n14018), .B2(n14017), .A(n14016), .ZN(n14034) );
  MUX2_X1 U16003 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14034), .S(n14688), .Z(
        P1_U3545) );
  MUX2_X1 U16004 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n14019), .S(n14688), .Z(
        P1_U3529) );
  MUX2_X1 U16005 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14020), .S(n14675), .Z(
        P1_U3527) );
  MUX2_X1 U16006 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14021), .S(n14675), .Z(
        P1_U3526) );
  MUX2_X1 U16007 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14023), .S(n14675), .Z(
        P1_U3524) );
  MUX2_X1 U16008 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14024), .S(n14675), .Z(
        P1_U3523) );
  MUX2_X1 U16009 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14025), .S(n14675), .Z(
        P1_U3522) );
  MUX2_X1 U16010 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14026), .S(n14675), .Z(
        P1_U3521) );
  MUX2_X1 U16011 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14027), .S(n14675), .Z(
        P1_U3520) );
  MUX2_X1 U16012 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14028), .S(n14675), .Z(
        P1_U3519) );
  MUX2_X1 U16013 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14029), .S(n14675), .Z(
        P1_U3518) );
  MUX2_X1 U16014 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14030), .S(n14675), .Z(
        P1_U3517) );
  MUX2_X1 U16015 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14031), .S(n14675), .Z(
        P1_U3516) );
  MUX2_X1 U16016 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14032), .S(n14675), .Z(
        P1_U3515) );
  MUX2_X1 U16017 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14033), .S(n14675), .Z(
        P1_U3513) );
  MUX2_X1 U16018 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14034), .S(n14675), .Z(
        P1_U3510) );
  OAI222_X1 U16019 ( .A1(n14037), .A2(P1_U3086), .B1(n10724), .B2(n14036), 
        .C1(n14035), .C2(n14039), .ZN(P1_U3326) );
  INV_X1 U16020 ( .A(n14038), .ZN(n14042) );
  OAI222_X1 U16021 ( .A1(P1_U3086), .A2(n14042), .B1(n10724), .B2(n14041), 
        .C1(n14040), .C2(n14039), .ZN(P1_U3329) );
  MUX2_X1 U16022 ( .A(n10298), .B(n14043), .S(P1_U3086), .Z(P1_U3333) );
  MUX2_X1 U16023 ( .A(n14045), .B(n14044), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3355) );
  INV_X1 U16024 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n15402) );
  INV_X1 U16025 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n14117) );
  INV_X1 U16026 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n14452) );
  INV_X1 U16027 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n15062) );
  XOR2_X1 U16028 ( .A(n15062), .B(P1_ADDR_REG_12__SCAN_IN), .Z(n14114) );
  XOR2_X1 U16029 ( .A(n15040), .B(P1_ADDR_REG_11__SCAN_IN), .Z(n14112) );
  XOR2_X1 U16030 ( .A(n15282), .B(P1_ADDR_REG_9__SCAN_IN), .Z(n14105) );
  XNOR2_X1 U16031 ( .A(n15366), .B(n14046), .ZN(n14099) );
  XNOR2_X1 U16032 ( .A(n14047), .B(n14989), .ZN(n14094) );
  NAND2_X1 U16033 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n14048), .ZN(n14051) );
  NAND2_X1 U16034 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n14052), .ZN(n14053) );
  NAND2_X1 U16035 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n14054), .ZN(n14057) );
  NAND2_X1 U16036 ( .A1(n14057), .A2(n14056), .ZN(n14095) );
  NAND2_X1 U16037 ( .A1(n14094), .A2(n14095), .ZN(n14058) );
  NAND2_X1 U16038 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n14059), .ZN(n14062) );
  NAND2_X1 U16039 ( .A1(n14097), .A2(n14060), .ZN(n14061) );
  NAND2_X1 U16040 ( .A1(n14062), .A2(n14061), .ZN(n14100) );
  NAND2_X1 U16041 ( .A1(n14099), .A2(n14100), .ZN(n14063) );
  NAND2_X1 U16042 ( .A1(n14105), .A2(n14104), .ZN(n14064) );
  NAND2_X1 U16043 ( .A1(n14066), .A2(n14065), .ZN(n14068) );
  XOR2_X1 U16044 ( .A(n14066), .B(n14065), .Z(n14108) );
  NAND2_X1 U16045 ( .A1(P3_ADDR_REG_10__SCAN_IN), .A2(n14108), .ZN(n14067) );
  NAND2_X1 U16046 ( .A1(n14068), .A2(n14067), .ZN(n14111) );
  NAND2_X1 U16047 ( .A1(n14112), .A2(n14111), .ZN(n14069) );
  NAND2_X1 U16048 ( .A1(n14114), .A2(n14113), .ZN(n14070) );
  INV_X1 U16049 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n15075) );
  NAND2_X1 U16050 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n15075), .ZN(n14071) );
  AOI22_X1 U16051 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n14452), .B1(n14073), 
        .B2(n14071), .ZN(n14072) );
  INV_X1 U16052 ( .A(n14072), .ZN(n14119) );
  INV_X1 U16053 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n15099) );
  XNOR2_X1 U16054 ( .A(n15099), .B(P1_ADDR_REG_14__SCAN_IN), .ZN(n14118) );
  XOR2_X1 U16055 ( .A(n14119), .B(n14118), .Z(n14419) );
  INV_X1 U16056 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n15485) );
  XOR2_X1 U16057 ( .A(n15075), .B(P1_ADDR_REG_13__SCAN_IN), .Z(n14074) );
  XNOR2_X1 U16058 ( .A(n14074), .B(n14073), .ZN(n14415) );
  NOR2_X1 U16059 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n14087), .ZN(n14089) );
  INV_X1 U16060 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n14084) );
  XNOR2_X1 U16061 ( .A(n14076), .B(n14075), .ZN(n14141) );
  XNOR2_X1 U16062 ( .A(n14077), .B(n14078), .ZN(n14080) );
  NAND2_X1 U16063 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14080), .ZN(n14082) );
  AOI21_X1 U16064 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n14079), .A(n14078), .ZN(
        n15604) );
  INV_X1 U16065 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15603) );
  NOR2_X1 U16066 ( .A1(n15604), .A2(n15603), .ZN(n15616) );
  NAND2_X1 U16067 ( .A1(n14082), .A2(n14081), .ZN(n14142) );
  NAND2_X1 U16068 ( .A1(n14141), .A2(n14142), .ZN(n14083) );
  NOR2_X1 U16069 ( .A1(n14141), .A2(n14142), .ZN(n14140) );
  XOR2_X1 U16070 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n14085), .Z(n15612) );
  NOR2_X1 U16071 ( .A1(n15611), .A2(n15612), .ZN(n14086) );
  INV_X1 U16072 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15613) );
  NAND2_X1 U16073 ( .A1(n15611), .A2(n15612), .ZN(n15610) );
  OAI21_X1 U16074 ( .B1(n14086), .B2(n15613), .A(n15610), .ZN(n15606) );
  XNOR2_X1 U16075 ( .A(P2_ADDR_REG_4__SCAN_IN), .B(n14087), .ZN(n15605) );
  NOR2_X1 U16076 ( .A1(n15606), .A2(n15605), .ZN(n14088) );
  NAND2_X1 U16077 ( .A1(n14093), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14096) );
  INV_X1 U16078 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n14733) );
  XNOR2_X1 U16079 ( .A(n14095), .B(n14094), .ZN(n14144) );
  XOR2_X1 U16080 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n14097), .Z(n15609) );
  XNOR2_X1 U16081 ( .A(n14100), .B(n14099), .ZN(n14102) );
  NAND2_X1 U16082 ( .A1(n14101), .A2(n14102), .ZN(n14103) );
  XNOR2_X1 U16083 ( .A(n14105), .B(n14104), .ZN(n14148) );
  NOR2_X1 U16084 ( .A1(n14149), .A2(n14148), .ZN(n14106) );
  INV_X1 U16085 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n15462) );
  NAND2_X1 U16086 ( .A1(n14149), .A2(n14148), .ZN(n14147) );
  XOR2_X1 U16087 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(n14108), .Z(n14109) );
  XNOR2_X1 U16088 ( .A(n14112), .B(n14111), .ZN(n14411) );
  INV_X1 U16089 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n14775) );
  XNOR2_X1 U16090 ( .A(n14114), .B(n14113), .ZN(n14115) );
  NOR2_X1 U16091 ( .A1(n14415), .A2(n14416), .ZN(n14414) );
  INV_X1 U16092 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14482) );
  XOR2_X1 U16093 ( .A(n14482), .B(P3_ADDR_REG_15__SCAN_IN), .Z(n14121) );
  NOR2_X1 U16094 ( .A1(n14119), .A2(n14118), .ZN(n14120) );
  AOI21_X1 U16095 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n15099), .A(n14120), 
        .ZN(n14125) );
  XNOR2_X1 U16096 ( .A(n14121), .B(n14125), .ZN(n14123) );
  NOR2_X1 U16097 ( .A1(n14122), .A2(n14123), .ZN(n14423) );
  INV_X1 U16098 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14129) );
  XOR2_X1 U16099 ( .A(n14129), .B(P1_ADDR_REG_16__SCAN_IN), .Z(n14127) );
  OR2_X1 U16100 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n14482), .ZN(n14126) );
  AOI22_X1 U16101 ( .A1(n14126), .A2(n14125), .B1(n14482), .B2(
        P3_ADDR_REG_15__SCAN_IN), .ZN(n14131) );
  XOR2_X1 U16102 ( .A(n14127), .B(n14131), .Z(n14128) );
  INV_X1 U16103 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n14512) );
  INV_X1 U16104 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n14497) );
  NAND2_X1 U16105 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n14497), .ZN(n14130) );
  AOI22_X1 U16106 ( .A1(n14131), .A2(n14130), .B1(P1_ADDR_REG_16__SCAN_IN), 
        .B2(n14129), .ZN(n14133) );
  XOR2_X1 U16107 ( .A(n14512), .B(n14133), .Z(n14134) );
  XOR2_X1 U16108 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n14134), .Z(n14132) );
  INV_X1 U16109 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n14530) );
  INV_X1 U16110 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n14181) );
  AND2_X1 U16111 ( .A1(n14512), .A2(n14133), .ZN(n14136) );
  AND2_X1 U16112 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n14134), .ZN(n14135) );
  NOR2_X1 U16113 ( .A1(n14136), .A2(n14135), .ZN(n14183) );
  XNOR2_X1 U16114 ( .A(n14181), .B(n14183), .ZN(n14137) );
  XOR2_X1 U16115 ( .A(n14530), .B(n14137), .Z(n14187) );
  XOR2_X1 U16116 ( .A(n15402), .B(n14189), .Z(SUB_1596_U62) );
  AOI21_X1 U16117 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14138) );
  OAI21_X1 U16118 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14138), 
        .ZN(U28) );
  INV_X1 U16119 ( .A(P2_RD_REG_SCAN_IN), .ZN(n14139) );
  INV_X1 U16120 ( .A(P3_RD_REG_SCAN_IN), .ZN(n15350) );
  OAI221_X1 U16121 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .C1(
        n14139), .C2(n7476), .A(n15350), .ZN(U29) );
  AOI21_X1 U16122 ( .B1(n14142), .B2(n14141), .A(n14140), .ZN(n14143) );
  XOR2_X1 U16123 ( .A(n14143), .B(P2_ADDR_REG_2__SCAN_IN), .Z(SUB_1596_U61) );
  XOR2_X1 U16124 ( .A(n14145), .B(n14144), .Z(SUB_1596_U57) );
  XOR2_X1 U16125 ( .A(n14146), .B(P2_ADDR_REG_8__SCAN_IN), .Z(SUB_1596_U55) );
  OAI21_X1 U16126 ( .B1(n14149), .B2(n14148), .A(n14147), .ZN(n14150) );
  XOR2_X1 U16127 ( .A(n14150), .B(n15462), .Z(SUB_1596_U54) );
  NOR2_X1 U16128 ( .A1(n14152), .A2(n14151), .ZN(n14153) );
  XOR2_X1 U16129 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n14153), .Z(SUB_1596_U70)
         );
  INV_X1 U16130 ( .A(n14158), .ZN(n14160) );
  AOI211_X1 U16131 ( .C1(n14632), .C2(n14156), .A(n14155), .B(n14154), .ZN(
        n14157) );
  OAI21_X1 U16132 ( .B1(n14158), .B2(n14636), .A(n14157), .ZN(n14159) );
  AOI21_X1 U16133 ( .B1(n14639), .B2(n14160), .A(n14159), .ZN(n14162) );
  INV_X1 U16134 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14161) );
  AOI22_X1 U16135 ( .A1(n14675), .A2(n14162), .B1(n14161), .B2(n14673), .ZN(
        P1_U3495) );
  AOI22_X1 U16136 ( .A1(n14688), .A2(n14162), .B1(n15414), .B2(n14686), .ZN(
        P1_U3540) );
  OAI211_X1 U16137 ( .C1(n14165), .C2(n14164), .A(n14163), .B(n14554), .ZN(
        n14167) );
  AOI222_X1 U16138 ( .A1(n14169), .A2(n14557), .B1(n14168), .B2(n14569), .C1(
        P1_REG2_REG_13__SCAN_IN), .C2(n14570), .ZN(n14177) );
  XNOR2_X1 U16139 ( .A(n14170), .B(n14171), .ZN(n14393) );
  OAI211_X1 U16140 ( .C1(n14173), .C2(n14391), .A(n14561), .B(n14172), .ZN(
        n14389) );
  INV_X1 U16141 ( .A(n14389), .ZN(n14174) );
  AOI22_X1 U16142 ( .A1(n14393), .A2(n14175), .B1(n14567), .B2(n14174), .ZN(
        n14176) );
  OAI211_X1 U16143 ( .C1(n13930), .C2(n14390), .A(n14177), .B(n14176), .ZN(
        P1_U3280) );
  INV_X1 U16144 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n14816) );
  NOR2_X1 U16145 ( .A1(n14179), .A2(n14178), .ZN(n14180) );
  XNOR2_X1 U16146 ( .A(n14816), .B(n14180), .ZN(SUB_1596_U63) );
  NAND2_X1 U16147 ( .A1(P3_ADDR_REG_18__SCAN_IN), .A2(n14530), .ZN(n14182) );
  AOI22_X1 U16148 ( .A1(n14183), .A2(n14182), .B1(P1_ADDR_REG_18__SCAN_IN), 
        .B2(n14181), .ZN(n14185) );
  XNOR2_X1 U16149 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n14184) );
  XNOR2_X1 U16150 ( .A(n14185), .B(n14184), .ZN(n14186) );
  AOI21_X1 U16151 ( .B1(n14192), .B2(n14191), .A(n14190), .ZN(n14207) );
  AOI21_X1 U16152 ( .B1(n14195), .B2(n14194), .A(n14193), .ZN(n14196) );
  NOR2_X1 U16153 ( .A1(n14196), .A2(n15095), .ZN(n14200) );
  OAI21_X1 U16154 ( .B1(n15101), .B2(n14198), .A(n14197), .ZN(n14199) );
  AOI211_X1 U16155 ( .C1(P3_ADDR_REG_15__SCAN_IN), .C2(n15025), .A(n14200), 
        .B(n14199), .ZN(n14206) );
  AOI211_X1 U16156 ( .C1(n14203), .C2(n14202), .A(n15082), .B(n14201), .ZN(
        n14204) );
  INV_X1 U16157 ( .A(n14204), .ZN(n14205) );
  OAI211_X1 U16158 ( .C1(n14207), .C2(n15110), .A(n14206), .B(n14205), .ZN(
        P3_U3197) );
  AOI21_X1 U16159 ( .B1(n6704), .B2(n14209), .A(n14208), .ZN(n14222) );
  AOI21_X1 U16160 ( .B1(n6705), .B2(n14211), .A(n14210), .ZN(n14212) );
  NOR2_X1 U16161 ( .A1(n14212), .A2(n15095), .ZN(n14216) );
  NAND2_X1 U16162 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(P3_U3151), .ZN(n14213)
         );
  OAI21_X1 U16163 ( .B1(n15101), .B2(n14214), .A(n14213), .ZN(n14215) );
  AOI211_X1 U16164 ( .C1(n15025), .C2(P3_ADDR_REG_16__SCAN_IN), .A(n14216), 
        .B(n14215), .ZN(n14221) );
  XOR2_X1 U16165 ( .A(n14218), .B(n14217), .Z(n14219) );
  NAND2_X1 U16166 ( .A1(n14219), .A2(n15104), .ZN(n14220) );
  OAI211_X1 U16167 ( .C1(n14222), .C2(n15110), .A(n14221), .B(n14220), .ZN(
        P3_U3198) );
  AOI21_X1 U16168 ( .B1(n14225), .B2(n14224), .A(n14223), .ZN(n14239) );
  AOI21_X1 U16169 ( .B1(n14228), .B2(n14227), .A(n14226), .ZN(n14229) );
  NOR2_X1 U16170 ( .A1(n14229), .A2(n15095), .ZN(n14233) );
  OAI21_X1 U16171 ( .B1(n15101), .B2(n14231), .A(n14230), .ZN(n14232) );
  AOI211_X1 U16172 ( .C1(n15025), .C2(P3_ADDR_REG_17__SCAN_IN), .A(n14233), 
        .B(n14232), .ZN(n14238) );
  OAI211_X1 U16173 ( .C1(n14236), .C2(n14235), .A(n14234), .B(n15104), .ZN(
        n14237) );
  OAI211_X1 U16174 ( .C1(n14239), .C2(n15110), .A(n14238), .B(n14237), .ZN(
        P3_U3199) );
  AOI21_X1 U16175 ( .B1(n6706), .B2(n14241), .A(n14240), .ZN(n14254) );
  OAI21_X1 U16176 ( .B1(n15101), .B2(n14243), .A(n14242), .ZN(n14253) );
  AOI21_X1 U16177 ( .B1(n14246), .B2(n14245), .A(n14244), .ZN(n14251) );
  AOI21_X1 U16178 ( .B1(n14249), .B2(n14248), .A(n14247), .ZN(n14250) );
  OAI22_X1 U16179 ( .A1(n14251), .A2(n15095), .B1(n14250), .B2(n15082), .ZN(
        n14252) );
  XNOR2_X1 U16180 ( .A(n14255), .B(n14260), .ZN(n14257) );
  AOI21_X1 U16181 ( .B1(n14257), .B2(n15122), .A(n14256), .ZN(n14279) );
  AOI22_X1 U16182 ( .A1(n15595), .A2(P3_REG2_REG_13__SCAN_IN), .B1(n15591), 
        .B2(n14258), .ZN(n14263) );
  XNOR2_X1 U16183 ( .A(n14259), .B(n14260), .ZN(n14282) );
  NOR2_X1 U16184 ( .A1(n14261), .A2(n15146), .ZN(n14281) );
  AOI22_X1 U16185 ( .A1(n14282), .A2(n15600), .B1(n14281), .B2(n14276), .ZN(
        n14262) );
  OAI211_X1 U16186 ( .C1(n15595), .C2(n14279), .A(n14263), .B(n14262), .ZN(
        P3_U3220) );
  AOI21_X1 U16187 ( .B1(n14265), .B2(n14272), .A(n14264), .ZN(n14268) );
  AOI21_X1 U16188 ( .B1(n14268), .B2(n14267), .A(n14266), .ZN(n14283) );
  OAI22_X1 U16189 ( .A1(n15131), .A2(n12417), .B1(n14270), .B2(n14269), .ZN(
        n14271) );
  INV_X1 U16190 ( .A(n14271), .ZN(n14278) );
  XNOR2_X1 U16191 ( .A(n14273), .B(n14272), .ZN(n14286) );
  INV_X1 U16192 ( .A(n14274), .ZN(n14275) );
  NOR2_X1 U16193 ( .A1(n14275), .A2(n15146), .ZN(n14285) );
  AOI22_X1 U16194 ( .A1(n14286), .A2(n15600), .B1(n14285), .B2(n14276), .ZN(
        n14277) );
  OAI211_X1 U16195 ( .C1(n15595), .C2(n14283), .A(n14278), .B(n14277), .ZN(
        P3_U3221) );
  INV_X1 U16196 ( .A(n14279), .ZN(n14280) );
  AOI211_X1 U16197 ( .C1(n14282), .C2(n14289), .A(n14281), .B(n14280), .ZN(
        n14295) );
  AOI22_X1 U16198 ( .A1(n15202), .A2(n14295), .B1(n15078), .B2(n8976), .ZN(
        P3_U3472) );
  INV_X1 U16199 ( .A(n14283), .ZN(n14284) );
  AOI211_X1 U16200 ( .C1(n14286), .C2(n14289), .A(n14285), .B(n14284), .ZN(
        n14297) );
  AOI22_X1 U16201 ( .A1(n15202), .A2(n14297), .B1(n12467), .B2(n8976), .ZN(
        P3_U3471) );
  OAI21_X1 U16202 ( .B1(n6792), .B2(n14290), .A(n14287), .ZN(n15599) );
  AOI22_X1 U16203 ( .A1(n15599), .A2(n14289), .B1(n14288), .B2(n15157), .ZN(
        n14294) );
  XNOR2_X1 U16204 ( .A(n14291), .B(n14290), .ZN(n14293) );
  AOI21_X1 U16205 ( .B1(n14293), .B2(n15122), .A(n14292), .ZN(n15596) );
  AND2_X1 U16206 ( .A1(n14294), .A2(n15596), .ZN(n14299) );
  AOI22_X1 U16207 ( .A1(n15202), .A2(n14299), .B1(n15044), .B2(n8976), .ZN(
        P3_U3470) );
  INV_X1 U16208 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14296) );
  AOI22_X1 U16209 ( .A1(n15183), .A2(n14296), .B1(n14295), .B2(n15181), .ZN(
        P3_U3429) );
  INV_X1 U16210 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14298) );
  AOI22_X1 U16211 ( .A1(n15183), .A2(n14298), .B1(n14297), .B2(n15181), .ZN(
        P3_U3426) );
  INV_X1 U16212 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14300) );
  AOI22_X1 U16213 ( .A1(n15183), .A2(n14300), .B1(n14299), .B2(n15181), .ZN(
        P3_U3423) );
  XNOR2_X1 U16214 ( .A(n14301), .B(n14309), .ZN(n14305) );
  INV_X1 U16215 ( .A(n14302), .ZN(n14303) );
  AOI21_X1 U16216 ( .B1(n14305), .B2(n14304), .A(n14303), .ZN(n14320) );
  AOI222_X1 U16217 ( .A1(n14308), .A2(n14307), .B1(P2_REG2_REG_14__SCAN_IN), 
        .B2(n13216), .C1(n14841), .C2(n14306), .ZN(n14318) );
  XNOR2_X1 U16218 ( .A(n14310), .B(n14309), .ZN(n14323) );
  OAI211_X1 U16219 ( .C1(n7218), .C2(n7219), .A(n14313), .B(n14312), .ZN(
        n14319) );
  INV_X1 U16220 ( .A(n14319), .ZN(n14314) );
  AOI22_X1 U16221 ( .A1(n14323), .A2(n14316), .B1(n14315), .B2(n14314), .ZN(
        n14317) );
  OAI211_X1 U16222 ( .C1(n13216), .C2(n14320), .A(n14318), .B(n14317), .ZN(
        P2_U3251) );
  OAI21_X1 U16223 ( .B1(n7218), .B2(n14915), .A(n14319), .ZN(n14322) );
  INV_X1 U16224 ( .A(n14320), .ZN(n14321) );
  AOI211_X1 U16225 ( .C1(n14905), .C2(n14323), .A(n14322), .B(n14321), .ZN(
        n14337) );
  AOI22_X1 U16226 ( .A1(n14934), .A2(n14337), .B1(n10330), .B2(n14932), .ZN(
        P2_U3513) );
  OAI21_X1 U16227 ( .B1(n14325), .B2(n14915), .A(n14324), .ZN(n14327) );
  AOI211_X1 U16228 ( .C1(n14328), .C2(n14905), .A(n14327), .B(n14326), .ZN(
        n14339) );
  AOI22_X1 U16229 ( .A1(n14934), .A2(n14339), .B1(n10068), .B2(n14932), .ZN(
        P2_U3512) );
  NAND2_X1 U16230 ( .A1(n14329), .A2(n14892), .ZN(n14330) );
  NAND2_X1 U16231 ( .A1(n14331), .A2(n14330), .ZN(n14332) );
  AOI21_X1 U16232 ( .B1(n14333), .B2(n14918), .A(n14332), .ZN(n14334) );
  AOI22_X1 U16233 ( .A1(n14934), .A2(n14341), .B1(n10074), .B2(n14932), .ZN(
        P2_U3511) );
  INV_X1 U16234 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n14336) );
  AOI22_X1 U16235 ( .A1(n14924), .A2(n14337), .B1(n14336), .B2(n14922), .ZN(
        P2_U3472) );
  INV_X1 U16236 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n14338) );
  AOI22_X1 U16237 ( .A1(n14924), .A2(n14339), .B1(n14338), .B2(n14922), .ZN(
        P2_U3469) );
  INV_X1 U16238 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14340) );
  AOI22_X1 U16239 ( .A1(n14924), .A2(n14341), .B1(n14340), .B2(n14922), .ZN(
        P2_U3466) );
  OAI21_X1 U16240 ( .B1(n14344), .B2(n14343), .A(n14342), .ZN(n14345) );
  AOI222_X1 U16241 ( .A1(n14382), .A2(n14359), .B1(n14345), .B2(n14350), .C1(
        n14383), .C2(n14358), .ZN(n14346) );
  NAND2_X1 U16242 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14466)
         );
  OAI211_X1 U16243 ( .C1(n14365), .C2(n14347), .A(n14346), .B(n14466), .ZN(
        P1_U3215) );
  INV_X1 U16244 ( .A(n14348), .ZN(n14356) );
  OAI211_X1 U16245 ( .C1(n14353), .C2(n14352), .A(n14351), .B(n14350), .ZN(
        n14354) );
  INV_X1 U16246 ( .A(n14354), .ZN(n14355) );
  AOI211_X1 U16247 ( .C1(n14358), .C2(n14357), .A(n14356), .B(n14355), .ZN(
        n14363) );
  INV_X1 U16248 ( .A(n14663), .ZN(n14361) );
  OAI21_X1 U16249 ( .B1(n14361), .B2(n14360), .A(n14359), .ZN(n14362) );
  OAI211_X1 U16250 ( .C1(n14365), .C2(n14364), .A(n14363), .B(n14362), .ZN(
        P1_U3217) );
  AOI21_X1 U16251 ( .B1(n14367), .B2(n14632), .A(n14366), .ZN(n14369) );
  OAI211_X1 U16252 ( .C1(n14370), .C2(n14666), .A(n14369), .B(n14368), .ZN(
        n14371) );
  AOI21_X1 U16253 ( .B1(n14372), .B2(n14671), .A(n14371), .ZN(n14400) );
  AOI22_X1 U16254 ( .A1(n14688), .A2(n14400), .B1(n14373), .B2(n14686), .ZN(
        P1_U3544) );
  AOI21_X1 U16255 ( .B1(n14375), .B2(n14632), .A(n14374), .ZN(n14377) );
  NAND3_X1 U16256 ( .A1(n14378), .A2(n14377), .A3(n14376), .ZN(n14379) );
  AOI21_X1 U16257 ( .B1(n14671), .B2(n14380), .A(n14379), .ZN(n14402) );
  AOI22_X1 U16258 ( .A1(n14688), .A2(n14402), .B1(n15488), .B2(n14686), .ZN(
        P1_U3543) );
  AOI211_X1 U16259 ( .C1(n14632), .C2(n14383), .A(n14382), .B(n14381), .ZN(
        n14386) );
  NAND3_X1 U16260 ( .A1(n7679), .A2(n14384), .A3(n14671), .ZN(n14385) );
  OAI211_X1 U16261 ( .C1(n14387), .C2(n14666), .A(n14386), .B(n14385), .ZN(
        n14388) );
  INV_X1 U16262 ( .A(n14388), .ZN(n14404) );
  AOI22_X1 U16263 ( .A1(n14688), .A2(n14404), .B1(n13669), .B2(n14686), .ZN(
        P1_U3542) );
  OAI211_X1 U16264 ( .C1(n14391), .C2(n14665), .A(n14390), .B(n14389), .ZN(
        n14392) );
  AOI21_X1 U16265 ( .B1(n14393), .B2(n14671), .A(n14392), .ZN(n14406) );
  AOI22_X1 U16266 ( .A1(n14688), .A2(n14406), .B1(n13672), .B2(n14686), .ZN(
        P1_U3541) );
  OAI21_X1 U16267 ( .B1(n14395), .B2(n14665), .A(n14394), .ZN(n14397) );
  AOI211_X1 U16268 ( .C1(n14398), .C2(n14671), .A(n14397), .B(n14396), .ZN(
        n14408) );
  AOI22_X1 U16269 ( .A1(n14688), .A2(n14408), .B1(n10415), .B2(n14686), .ZN(
        P1_U3539) );
  INV_X1 U16270 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n14399) );
  AOI22_X1 U16271 ( .A1(n14675), .A2(n14400), .B1(n14399), .B2(n14673), .ZN(
        P1_U3507) );
  INV_X1 U16272 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n14401) );
  AOI22_X1 U16273 ( .A1(n14675), .A2(n14402), .B1(n14401), .B2(n14673), .ZN(
        P1_U3504) );
  INV_X1 U16274 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14403) );
  AOI22_X1 U16275 ( .A1(n14675), .A2(n14404), .B1(n14403), .B2(n14673), .ZN(
        P1_U3501) );
  INV_X1 U16276 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n14405) );
  AOI22_X1 U16277 ( .A1(n14675), .A2(n14406), .B1(n14405), .B2(n14673), .ZN(
        P1_U3498) );
  INV_X1 U16278 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14407) );
  AOI22_X1 U16279 ( .A1(n14675), .A2(n14408), .B1(n14407), .B2(n14673), .ZN(
        P1_U3492) );
  OAI21_X1 U16280 ( .B1(n14411), .B2(n14410), .A(n14409), .ZN(n14412) );
  XOR2_X1 U16281 ( .A(n14412), .B(n14775), .Z(SUB_1596_U69) );
  INV_X1 U16282 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n15450) );
  XOR2_X1 U16283 ( .A(n15450), .B(n14413), .Z(SUB_1596_U68) );
  AOI21_X1 U16284 ( .B1(n14416), .B2(n14415), .A(n14414), .ZN(n14417) );
  XOR2_X1 U16285 ( .A(n14417), .B(P2_ADDR_REG_13__SCAN_IN), .Z(SUB_1596_U67)
         );
  AOI21_X1 U16286 ( .B1(n14420), .B2(n14419), .A(n14418), .ZN(n14421) );
  XOR2_X1 U16287 ( .A(n14421), .B(P2_ADDR_REG_14__SCAN_IN), .Z(SUB_1596_U66)
         );
  NOR2_X1 U16288 ( .A1(n14423), .A2(n14422), .ZN(n14424) );
  XOR2_X1 U16289 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n14424), .Z(SUB_1596_U65)
         );
  NOR2_X1 U16290 ( .A1(n14426), .A2(n14425), .ZN(n14427) );
  XOR2_X1 U16291 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n14427), .Z(SUB_1596_U64)
         );
  INV_X1 U16292 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n14440) );
  OAI21_X1 U16293 ( .B1(n14430), .B2(n14429), .A(n14428), .ZN(n14437) );
  NOR2_X1 U16294 ( .A1(n14525), .A2(n14431), .ZN(n14436) );
  AOI211_X1 U16295 ( .C1(n14434), .C2(n14433), .A(n14487), .B(n14432), .ZN(
        n14435) );
  AOI211_X1 U16296 ( .C1(n14517), .C2(n14437), .A(n14436), .B(n14435), .ZN(
        n14439) );
  NAND2_X1 U16297 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14438)
         );
  OAI211_X1 U16298 ( .C1(n14440), .C2(n14529), .A(n14439), .B(n14438), .ZN(
        P1_U3254) );
  AOI211_X1 U16299 ( .C1(n14443), .C2(n14442), .A(n14441), .B(n14483), .ZN(
        n14448) );
  AOI211_X1 U16300 ( .C1(n14446), .C2(n14445), .A(n14444), .B(n14487), .ZN(
        n14447) );
  AOI211_X1 U16301 ( .C1(n14494), .C2(n14449), .A(n14448), .B(n14447), .ZN(
        n14451) );
  OAI211_X1 U16302 ( .C1(n14452), .C2(n14529), .A(n14451), .B(n14450), .ZN(
        P1_U3256) );
  INV_X1 U16303 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14468) );
  INV_X1 U16304 ( .A(n14453), .ZN(n14464) );
  OAI21_X1 U16305 ( .B1(n14456), .B2(n14455), .A(n14454), .ZN(n14457) );
  NAND2_X1 U16306 ( .A1(n14517), .A2(n14457), .ZN(n14463) );
  AOI21_X1 U16307 ( .B1(n14460), .B2(n14459), .A(n14458), .ZN(n14461) );
  NAND2_X1 U16308 ( .A1(n14521), .A2(n14461), .ZN(n14462) );
  OAI211_X1 U16309 ( .C1(n14525), .C2(n14464), .A(n14463), .B(n14462), .ZN(
        n14465) );
  INV_X1 U16310 ( .A(n14465), .ZN(n14467) );
  OAI211_X1 U16311 ( .C1(n14468), .C2(n14529), .A(n14467), .B(n14466), .ZN(
        P1_U3257) );
  OAI21_X1 U16312 ( .B1(n14470), .B2(n15488), .A(n14469), .ZN(n14471) );
  NAND2_X1 U16313 ( .A1(n14517), .A2(n14471), .ZN(n14477) );
  OAI21_X1 U16314 ( .B1(n14474), .B2(n14473), .A(n14472), .ZN(n14475) );
  NAND2_X1 U16315 ( .A1(n14521), .A2(n14475), .ZN(n14476) );
  OAI211_X1 U16316 ( .C1(n14525), .C2(n14478), .A(n14477), .B(n14476), .ZN(
        n14479) );
  INV_X1 U16317 ( .A(n14479), .ZN(n14481) );
  OAI211_X1 U16318 ( .C1(n14482), .C2(n14529), .A(n14481), .B(n14480), .ZN(
        P1_U3258) );
  AOI211_X1 U16319 ( .C1(n14486), .C2(n14485), .A(n14484), .B(n14483), .ZN(
        n14492) );
  AOI211_X1 U16320 ( .C1(n14490), .C2(n14489), .A(n14488), .B(n14487), .ZN(
        n14491) );
  AOI211_X1 U16321 ( .C1(n14494), .C2(n14493), .A(n14492), .B(n14491), .ZN(
        n14496) );
  OAI211_X1 U16322 ( .C1(n14497), .C2(n14529), .A(n14496), .B(n14495), .ZN(
        P1_U3259) );
  AOI21_X1 U16323 ( .B1(n14500), .B2(n14499), .A(n14498), .ZN(n14501) );
  NAND2_X1 U16324 ( .A1(n14517), .A2(n14501), .ZN(n14507) );
  AOI21_X1 U16325 ( .B1(n14504), .B2(n14503), .A(n14502), .ZN(n14505) );
  NAND2_X1 U16326 ( .A1(n14521), .A2(n14505), .ZN(n14506) );
  OAI211_X1 U16327 ( .C1(n14525), .C2(n14508), .A(n14507), .B(n14506), .ZN(
        n14509) );
  INV_X1 U16328 ( .A(n14509), .ZN(n14511) );
  OAI211_X1 U16329 ( .C1(n14512), .C2(n14529), .A(n14511), .B(n14510), .ZN(
        P1_U3260) );
  AOI21_X1 U16330 ( .B1(n14515), .B2(n14514), .A(n14513), .ZN(n14516) );
  NAND2_X1 U16331 ( .A1(n14517), .A2(n14516), .ZN(n14523) );
  AOI21_X1 U16332 ( .B1(n14519), .B2(n15327), .A(n14518), .ZN(n14520) );
  NAND2_X1 U16333 ( .A1(n14521), .A2(n14520), .ZN(n14522) );
  OAI211_X1 U16334 ( .C1(n14525), .C2(n14524), .A(n14523), .B(n14522), .ZN(
        n14526) );
  INV_X1 U16335 ( .A(n14526), .ZN(n14528) );
  OAI211_X1 U16336 ( .C1(n14530), .C2(n14529), .A(n14528), .B(n14527), .ZN(
        P1_U3261) );
  XNOR2_X1 U16337 ( .A(n14531), .B(n14534), .ZN(n14661) );
  AOI21_X1 U16338 ( .B1(n14534), .B2(n14533), .A(n14532), .ZN(n14535) );
  OAI222_X1 U16339 ( .A1(n14539), .A2(n14538), .B1(n14537), .B2(n14536), .C1(
        n14666), .C2(n14535), .ZN(n14659) );
  AOI21_X1 U16340 ( .B1(n14639), .B2(n14661), .A(n14659), .ZN(n14547) );
  AOI222_X1 U16341 ( .A1(n14541), .A2(n14557), .B1(n14540), .B2(n14569), .C1(
        P1_REG2_REG_9__SCAN_IN), .C2(n14570), .ZN(n14546) );
  OAI211_X1 U16342 ( .C1(n14543), .C2(n14658), .A(n14561), .B(n14542), .ZN(
        n14657) );
  INV_X1 U16343 ( .A(n14657), .ZN(n14544) );
  AOI22_X1 U16344 ( .A1(n14661), .A2(n14577), .B1(n14567), .B2(n14544), .ZN(
        n14545) );
  OAI211_X1 U16345 ( .C1(n14570), .C2(n14547), .A(n14546), .B(n14545), .ZN(
        P1_U3284) );
  XNOR2_X1 U16346 ( .A(n14548), .B(n14549), .ZN(n14555) );
  XNOR2_X1 U16347 ( .A(n14550), .B(n14549), .ZN(n14559) );
  NOR2_X1 U16348 ( .A1(n14559), .A2(n14551), .ZN(n14553) );
  AOI211_X1 U16349 ( .C1(n14555), .C2(n14554), .A(n14553), .B(n14552), .ZN(
        n14643) );
  AOI222_X1 U16350 ( .A1(n14558), .A2(n14557), .B1(n14556), .B2(n14569), .C1(
        P1_REG2_REG_7__SCAN_IN), .C2(n14570), .ZN(n14566) );
  INV_X1 U16351 ( .A(n14559), .ZN(n14646) );
  INV_X1 U16352 ( .A(n14560), .ZN(n14562) );
  OAI211_X1 U16353 ( .C1(n14642), .C2(n14563), .A(n14562), .B(n14561), .ZN(
        n14641) );
  INV_X1 U16354 ( .A(n14641), .ZN(n14564) );
  AOI22_X1 U16355 ( .A1(n14646), .A2(n14577), .B1(n14567), .B2(n14564), .ZN(
        n14565) );
  OAI211_X1 U16356 ( .C1(n13930), .C2(n14643), .A(n14566), .B(n14565), .ZN(
        P1_U3286) );
  NAND2_X1 U16357 ( .A1(n14568), .A2(n14567), .ZN(n14572) );
  AOI22_X1 U16358 ( .A1(n14570), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n14569), .ZN(n14571) );
  OAI211_X1 U16359 ( .C1(n14574), .C2(n14573), .A(n14572), .B(n14571), .ZN(
        n14575) );
  AOI21_X1 U16360 ( .B1(n14577), .B2(n14576), .A(n14575), .ZN(n14578) );
  OAI21_X1 U16361 ( .B1(n14570), .B2(n14579), .A(n14578), .ZN(P1_U3291) );
  INV_X1 U16362 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n14580) );
  NOR2_X1 U16363 ( .A1(n14606), .A2(n14580), .ZN(P1_U3294) );
  NOR2_X1 U16364 ( .A1(n14606), .A2(n15567), .ZN(P1_U3295) );
  INV_X1 U16365 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n14581) );
  NOR2_X1 U16366 ( .A1(n14606), .A2(n14581), .ZN(P1_U3296) );
  INV_X1 U16367 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n14582) );
  NOR2_X1 U16368 ( .A1(n14606), .A2(n14582), .ZN(P1_U3297) );
  INV_X1 U16369 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n14583) );
  NOR2_X1 U16370 ( .A1(n14606), .A2(n14583), .ZN(P1_U3298) );
  INV_X1 U16371 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n14584) );
  NOR2_X1 U16372 ( .A1(n14606), .A2(n14584), .ZN(P1_U3299) );
  INV_X1 U16373 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n14585) );
  NOR2_X1 U16374 ( .A1(n14606), .A2(n14585), .ZN(P1_U3300) );
  INV_X1 U16375 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n14586) );
  NOR2_X1 U16376 ( .A1(n14606), .A2(n14586), .ZN(P1_U3301) );
  INV_X1 U16377 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n14587) );
  NOR2_X1 U16378 ( .A1(n14606), .A2(n14587), .ZN(P1_U3302) );
  INV_X1 U16379 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n14588) );
  NOR2_X1 U16380 ( .A1(n14606), .A2(n14588), .ZN(P1_U3303) );
  INV_X1 U16381 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n14589) );
  NOR2_X1 U16382 ( .A1(n14606), .A2(n14589), .ZN(P1_U3304) );
  INV_X1 U16383 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n14590) );
  NOR2_X1 U16384 ( .A1(n14606), .A2(n14590), .ZN(P1_U3305) );
  INV_X1 U16385 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n14591) );
  NOR2_X1 U16386 ( .A1(n14606), .A2(n14591), .ZN(P1_U3306) );
  INV_X1 U16387 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n14592) );
  NOR2_X1 U16388 ( .A1(n14606), .A2(n14592), .ZN(P1_U3307) );
  NOR2_X1 U16389 ( .A1(n14606), .A2(n15416), .ZN(P1_U3308) );
  INV_X1 U16390 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n14593) );
  NOR2_X1 U16391 ( .A1(n14606), .A2(n14593), .ZN(P1_U3309) );
  INV_X1 U16392 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n14594) );
  NOR2_X1 U16393 ( .A1(n14606), .A2(n14594), .ZN(P1_U3310) );
  INV_X1 U16394 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n14595) );
  NOR2_X1 U16395 ( .A1(n14606), .A2(n14595), .ZN(P1_U3311) );
  INV_X1 U16396 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n14596) );
  NOR2_X1 U16397 ( .A1(n14606), .A2(n14596), .ZN(P1_U3312) );
  INV_X1 U16398 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n14597) );
  NOR2_X1 U16399 ( .A1(n14606), .A2(n14597), .ZN(P1_U3313) );
  INV_X1 U16400 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n14598) );
  NOR2_X1 U16401 ( .A1(n14606), .A2(n14598), .ZN(P1_U3314) );
  INV_X1 U16402 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n14599) );
  NOR2_X1 U16403 ( .A1(n14606), .A2(n14599), .ZN(P1_U3315) );
  INV_X1 U16404 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n14600) );
  NOR2_X1 U16405 ( .A1(n14606), .A2(n14600), .ZN(P1_U3316) );
  INV_X1 U16406 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n14601) );
  NOR2_X1 U16407 ( .A1(n14606), .A2(n14601), .ZN(P1_U3317) );
  INV_X1 U16408 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n14602) );
  NOR2_X1 U16409 ( .A1(n14606), .A2(n14602), .ZN(P1_U3318) );
  INV_X1 U16410 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n14603) );
  NOR2_X1 U16411 ( .A1(n14606), .A2(n14603), .ZN(P1_U3319) );
  NOR2_X1 U16412 ( .A1(n14606), .A2(n15458), .ZN(P1_U3320) );
  NOR2_X1 U16413 ( .A1(n14606), .A2(n15283), .ZN(P1_U3321) );
  INV_X1 U16414 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n14604) );
  NOR2_X1 U16415 ( .A1(n14606), .A2(n14604), .ZN(P1_U3322) );
  INV_X1 U16416 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n14605) );
  NOR2_X1 U16417 ( .A1(n14606), .A2(n14605), .ZN(P1_U3323) );
  INV_X1 U16418 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n14607) );
  AOI22_X1 U16419 ( .A1(n14675), .A2(n14608), .B1(n14607), .B2(n14673), .ZN(
        P1_U3459) );
  INV_X1 U16420 ( .A(n14636), .ZN(n14647) );
  NAND2_X1 U16421 ( .A1(n14609), .A2(n14647), .ZN(n14611) );
  OAI211_X1 U16422 ( .C1(n14612), .C2(n14665), .A(n14611), .B(n14610), .ZN(
        n14614) );
  NOR2_X1 U16423 ( .A1(n14614), .A2(n14613), .ZN(n14676) );
  INV_X1 U16424 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n14615) );
  AOI22_X1 U16425 ( .A1(n14675), .A2(n14676), .B1(n14615), .B2(n14673), .ZN(
        P1_U3468) );
  NAND4_X1 U16426 ( .A1(n14619), .A2(n14618), .A3(n14617), .A4(n14616), .ZN(
        n14620) );
  AOI21_X1 U16427 ( .B1(n14621), .B2(n14671), .A(n14620), .ZN(n14678) );
  INV_X1 U16428 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n14622) );
  AOI22_X1 U16429 ( .A1(n14675), .A2(n14678), .B1(n14622), .B2(n14673), .ZN(
        P1_U3471) );
  NAND2_X1 U16430 ( .A1(n14628), .A2(n14639), .ZN(n14624) );
  NAND4_X1 U16431 ( .A1(n14626), .A2(n14625), .A3(n14624), .A4(n14623), .ZN(
        n14627) );
  AOI21_X1 U16432 ( .B1(n14647), .B2(n14628), .A(n14627), .ZN(n14680) );
  INV_X1 U16433 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n14629) );
  AOI22_X1 U16434 ( .A1(n14675), .A2(n14680), .B1(n14629), .B2(n14673), .ZN(
        P1_U3474) );
  INV_X1 U16435 ( .A(n14635), .ZN(n14638) );
  AOI21_X1 U16436 ( .B1(n14632), .B2(n14631), .A(n14630), .ZN(n14633) );
  OAI211_X1 U16437 ( .C1(n14636), .C2(n14635), .A(n14634), .B(n14633), .ZN(
        n14637) );
  AOI21_X1 U16438 ( .B1(n14639), .B2(n14638), .A(n14637), .ZN(n14682) );
  INV_X1 U16439 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n14640) );
  AOI22_X1 U16440 ( .A1(n14675), .A2(n14682), .B1(n14640), .B2(n14673), .ZN(
        P1_U3477) );
  OAI21_X1 U16441 ( .B1(n14642), .B2(n14665), .A(n14641), .ZN(n14645) );
  INV_X1 U16442 ( .A(n14643), .ZN(n14644) );
  AOI211_X1 U16443 ( .C1(n14647), .C2(n14646), .A(n14645), .B(n14644), .ZN(
        n14683) );
  INV_X1 U16444 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n14648) );
  AOI22_X1 U16445 ( .A1(n14675), .A2(n14683), .B1(n14648), .B2(n14673), .ZN(
        P1_U3480) );
  INV_X1 U16446 ( .A(n14649), .ZN(n14651) );
  NAND4_X1 U16447 ( .A1(n14653), .A2(n14652), .A3(n14651), .A4(n14650), .ZN(
        n14654) );
  AOI21_X1 U16448 ( .B1(n14671), .B2(n14655), .A(n14654), .ZN(n14684) );
  INV_X1 U16449 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14656) );
  AOI22_X1 U16450 ( .A1(n14675), .A2(n14684), .B1(n14656), .B2(n14673), .ZN(
        P1_U3483) );
  OAI21_X1 U16451 ( .B1(n14658), .B2(n14665), .A(n14657), .ZN(n14660) );
  AOI211_X1 U16452 ( .C1(n14661), .C2(n14671), .A(n14660), .B(n14659), .ZN(
        n14685) );
  INV_X1 U16453 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n14662) );
  AOI22_X1 U16454 ( .A1(n14675), .A2(n14685), .B1(n14662), .B2(n14673), .ZN(
        P1_U3486) );
  OAI211_X1 U16455 ( .C1(n11260), .C2(n14665), .A(n14664), .B(n14663), .ZN(
        n14670) );
  NOR3_X1 U16456 ( .A1(n14668), .A2(n14667), .A3(n14666), .ZN(n14669) );
  AOI211_X1 U16457 ( .C1(n14672), .C2(n14671), .A(n14670), .B(n14669), .ZN(
        n14687) );
  INV_X1 U16458 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n14674) );
  AOI22_X1 U16459 ( .A1(n14675), .A2(n14687), .B1(n14674), .B2(n14673), .ZN(
        P1_U3489) );
  AOI22_X1 U16460 ( .A1(n14688), .A2(n14676), .B1(n10132), .B2(n14686), .ZN(
        P1_U3531) );
  AOI22_X1 U16461 ( .A1(n14688), .A2(n14678), .B1(n14677), .B2(n14686), .ZN(
        P1_U3532) );
  INV_X1 U16462 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n14679) );
  AOI22_X1 U16463 ( .A1(n14688), .A2(n14680), .B1(n14679), .B2(n14686), .ZN(
        P1_U3533) );
  INV_X1 U16464 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n14681) );
  AOI22_X1 U16465 ( .A1(n14688), .A2(n14682), .B1(n14681), .B2(n14686), .ZN(
        P1_U3534) );
  AOI22_X1 U16466 ( .A1(n14688), .A2(n14683), .B1(n10134), .B2(n14686), .ZN(
        P1_U3535) );
  AOI22_X1 U16467 ( .A1(n14688), .A2(n14684), .B1(n10135), .B2(n14686), .ZN(
        P1_U3536) );
  AOI22_X1 U16468 ( .A1(n14688), .A2(n14685), .B1(n10136), .B2(n14686), .ZN(
        P1_U3537) );
  AOI22_X1 U16469 ( .A1(n14688), .A2(n14687), .B1(n10127), .B2(n14686), .ZN(
        P1_U3538) );
  NOR2_X1 U16470 ( .A1(n14825), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U16471 ( .A1(n14787), .A2(P2_REG1_REG_0__SCAN_IN), .B1(n14811), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n14692) );
  AOI22_X1 U16472 ( .A1(n14825), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n14691) );
  OAI22_X1 U16473 ( .A1(n14829), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n14819), .ZN(n14689) );
  OAI21_X1 U16474 ( .B1(n14809), .B2(n14689), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n14690) );
  OAI211_X1 U16475 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n14692), .A(n14691), .B(
        n14690), .ZN(P2_U3214) );
  AOI22_X1 U16476 ( .A1(n14825), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n14705) );
  XNOR2_X1 U16477 ( .A(n14694), .B(n14693), .ZN(n14698) );
  OR2_X1 U16478 ( .A1(n14696), .A2(n14695), .ZN(n14697) );
  OAI21_X1 U16479 ( .B1(n14819), .B2(n14698), .A(n14697), .ZN(n14699) );
  INV_X1 U16480 ( .A(n14699), .ZN(n14704) );
  OAI211_X1 U16481 ( .C1(n14702), .C2(n14701), .A(n14811), .B(n14700), .ZN(
        n14703) );
  NAND3_X1 U16482 ( .A1(n14705), .A2(n14704), .A3(n14703), .ZN(P2_U3215) );
  OAI21_X1 U16483 ( .B1(n14708), .B2(n14707), .A(n14706), .ZN(n14710) );
  OAI22_X1 U16484 ( .A1(n14819), .A2(n14710), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14709), .ZN(n14711) );
  INV_X1 U16485 ( .A(n14711), .ZN(n14713) );
  NAND2_X1 U16486 ( .A1(n14825), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n14712) );
  OAI211_X1 U16487 ( .C1(n14833), .C2(n14714), .A(n14713), .B(n14712), .ZN(
        n14715) );
  INV_X1 U16488 ( .A(n14715), .ZN(n14720) );
  OAI211_X1 U16489 ( .C1(n14718), .C2(n14717), .A(n14811), .B(n14716), .ZN(
        n14719) );
  NAND2_X1 U16490 ( .A1(n14720), .A2(n14719), .ZN(P2_U3216) );
  OAI211_X1 U16491 ( .C1(n14723), .C2(n14722), .A(n14787), .B(n14721), .ZN(
        n14725) );
  OAI211_X1 U16492 ( .C1(n14833), .C2(n14726), .A(n14725), .B(n14724), .ZN(
        n14727) );
  INV_X1 U16493 ( .A(n14727), .ZN(n14732) );
  OAI211_X1 U16494 ( .C1(n14730), .C2(n14729), .A(n14811), .B(n14728), .ZN(
        n14731) );
  OAI211_X1 U16495 ( .C1(n14817), .C2(n14733), .A(n14732), .B(n14731), .ZN(
        P2_U3220) );
  INV_X1 U16496 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n14746) );
  OAI211_X1 U16497 ( .C1(n14736), .C2(n14735), .A(n14734), .B(n14787), .ZN(
        n14737) );
  INV_X1 U16498 ( .A(n14737), .ZN(n14738) );
  AOI211_X1 U16499 ( .C1(n14809), .C2(n14740), .A(n14739), .B(n14738), .ZN(
        n14745) );
  OAI211_X1 U16500 ( .C1(n14743), .C2(n14742), .A(n14741), .B(n14811), .ZN(
        n14744) );
  OAI211_X1 U16501 ( .C1(n14817), .C2(n14746), .A(n14745), .B(n14744), .ZN(
        P2_U3222) );
  NAND2_X1 U16502 ( .A1(n14748), .A2(n14747), .ZN(n14749) );
  AOI21_X1 U16503 ( .B1(n14750), .B2(n14749), .A(n14819), .ZN(n14758) );
  NAND2_X1 U16504 ( .A1(n14752), .A2(n14751), .ZN(n14753) );
  AOI21_X1 U16505 ( .B1(n14754), .B2(n14753), .A(n14829), .ZN(n14757) );
  NOR2_X1 U16506 ( .A1(n14833), .A2(n14755), .ZN(n14756) );
  NOR3_X1 U16507 ( .A1(n14758), .A2(n14757), .A3(n14756), .ZN(n14760) );
  OAI211_X1 U16508 ( .C1(n15462), .C2(n14817), .A(n14760), .B(n14759), .ZN(
        P2_U3223) );
  NAND2_X1 U16509 ( .A1(n14762), .A2(n14761), .ZN(n14763) );
  NAND2_X1 U16510 ( .A1(n14782), .A2(n14763), .ZN(n14764) );
  NAND2_X1 U16511 ( .A1(n14764), .A2(n14811), .ZN(n14770) );
  NOR2_X1 U16512 ( .A1(n14766), .A2(n14765), .ZN(n14767) );
  OR3_X1 U16513 ( .A1(n14768), .A2(n14767), .A3(n14819), .ZN(n14769) );
  OAI211_X1 U16514 ( .C1(n14833), .C2(n14771), .A(n14770), .B(n14769), .ZN(
        n14772) );
  INV_X1 U16515 ( .A(n14772), .ZN(n14774) );
  OAI211_X1 U16516 ( .C1(n14775), .C2(n14817), .A(n14774), .B(n14773), .ZN(
        P2_U3225) );
  OAI21_X1 U16517 ( .B1(n14778), .B2(n14777), .A(n14776), .ZN(n14788) );
  INV_X1 U16518 ( .A(n14779), .ZN(n14784) );
  NAND3_X1 U16519 ( .A1(n14782), .A2(n14781), .A3(n14780), .ZN(n14783) );
  NAND2_X1 U16520 ( .A1(n14784), .A2(n14783), .ZN(n14785) );
  AOI222_X1 U16521 ( .A1(n14788), .A2(n14787), .B1(n14786), .B2(n14809), .C1(
        n14785), .C2(n14811), .ZN(n14790) );
  OAI211_X1 U16522 ( .C1(n15450), .C2(n14817), .A(n14790), .B(n14789), .ZN(
        P2_U3226) );
  AND2_X1 U16523 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n14795) );
  AOI211_X1 U16524 ( .C1(n14793), .C2(n14792), .A(n14791), .B(n14819), .ZN(
        n14794) );
  AOI211_X1 U16525 ( .C1(P2_ADDR_REG_16__SCAN_IN), .C2(n14825), .A(n14795), 
        .B(n14794), .ZN(n14800) );
  OAI211_X1 U16526 ( .C1(n14798), .C2(n14797), .A(n14811), .B(n14796), .ZN(
        n14799) );
  OAI211_X1 U16527 ( .C1(n14833), .C2(n14801), .A(n14800), .B(n14799), .ZN(
        P2_U3230) );
  NOR2_X1 U16528 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n14802), .ZN(n14807) );
  AOI211_X1 U16529 ( .C1(n14805), .C2(n14804), .A(n14803), .B(n14819), .ZN(
        n14806) );
  AOI211_X1 U16530 ( .C1(n14809), .C2(n14808), .A(n14807), .B(n14806), .ZN(
        n14815) );
  OAI211_X1 U16531 ( .C1(n14813), .C2(n14812), .A(n14811), .B(n14810), .ZN(
        n14814) );
  OAI211_X1 U16532 ( .C1(n14817), .C2(n14816), .A(n14815), .B(n14814), .ZN(
        P2_U3231) );
  NOR2_X1 U16533 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n14818), .ZN(n14824) );
  AOI211_X1 U16534 ( .C1(n14822), .C2(n14821), .A(n14820), .B(n14819), .ZN(
        n14823) );
  AOI211_X1 U16535 ( .C1(P2_ADDR_REG_18__SCAN_IN), .C2(n14825), .A(n14824), 
        .B(n14823), .ZN(n14831) );
  AOI21_X1 U16536 ( .B1(n14827), .B2(P2_REG2_REG_18__SCAN_IN), .A(n14826), 
        .ZN(n14828) );
  OR2_X1 U16537 ( .A1(n14829), .A2(n14828), .ZN(n14830) );
  OAI211_X1 U16538 ( .C1(n14833), .C2(n14832), .A(n14831), .B(n14830), .ZN(
        P2_U3232) );
  NOR2_X1 U16539 ( .A1(n14835), .A2(n14834), .ZN(n14840) );
  OAI21_X1 U16540 ( .B1(n9870), .B2(n14842), .A(n14836), .ZN(n14838) );
  MUX2_X1 U16541 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n14838), .S(n14837), .Z(
        n14839) );
  AOI211_X1 U16542 ( .C1(n14841), .C2(P2_REG3_REG_2__SCAN_IN), .A(n14840), .B(
        n14839), .ZN(n14848) );
  INV_X1 U16543 ( .A(n14842), .ZN(n14846) );
  AOI22_X1 U16544 ( .A1(n14846), .A2(n14845), .B1(n14844), .B2(n14843), .ZN(
        n14847) );
  NAND2_X1 U16545 ( .A1(n14848), .A2(n14847), .ZN(P2_U3263) );
  INV_X1 U16546 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n14850) );
  NOR2_X1 U16547 ( .A1(n14876), .A2(n14850), .ZN(P2_U3266) );
  INV_X1 U16548 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n15461) );
  NOR2_X1 U16549 ( .A1(n14876), .A2(n15461), .ZN(P2_U3267) );
  INV_X1 U16550 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n15426) );
  NOR2_X1 U16551 ( .A1(n14876), .A2(n15426), .ZN(P2_U3268) );
  INV_X1 U16552 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n14851) );
  NOR2_X1 U16553 ( .A1(n14872), .A2(n14851), .ZN(P2_U3269) );
  INV_X1 U16554 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n14852) );
  NOR2_X1 U16555 ( .A1(n14872), .A2(n14852), .ZN(P2_U3270) );
  INV_X1 U16556 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n14853) );
  NOR2_X1 U16557 ( .A1(n14872), .A2(n14853), .ZN(P2_U3271) );
  INV_X1 U16558 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n14854) );
  NOR2_X1 U16559 ( .A1(n14872), .A2(n14854), .ZN(P2_U3272) );
  INV_X1 U16560 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n14855) );
  NOR2_X1 U16561 ( .A1(n14872), .A2(n14855), .ZN(P2_U3273) );
  INV_X1 U16562 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n14856) );
  NOR2_X1 U16563 ( .A1(n14872), .A2(n14856), .ZN(P2_U3274) );
  INV_X1 U16564 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n14857) );
  NOR2_X1 U16565 ( .A1(n14872), .A2(n14857), .ZN(P2_U3275) );
  INV_X1 U16566 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n14858) );
  NOR2_X1 U16567 ( .A1(n14872), .A2(n14858), .ZN(P2_U3276) );
  INV_X1 U16568 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n14859) );
  NOR2_X1 U16569 ( .A1(n14872), .A2(n14859), .ZN(P2_U3277) );
  INV_X1 U16570 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n14860) );
  NOR2_X1 U16571 ( .A1(n14876), .A2(n14860), .ZN(P2_U3278) );
  INV_X1 U16572 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n14861) );
  NOR2_X1 U16573 ( .A1(n14876), .A2(n14861), .ZN(P2_U3279) );
  INV_X1 U16574 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n15341) );
  NOR2_X1 U16575 ( .A1(n14876), .A2(n15341), .ZN(P2_U3280) );
  INV_X1 U16576 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n14862) );
  NOR2_X1 U16577 ( .A1(n14876), .A2(n14862), .ZN(P2_U3281) );
  INV_X1 U16578 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n15459) );
  NOR2_X1 U16579 ( .A1(n14876), .A2(n15459), .ZN(P2_U3282) );
  INV_X1 U16580 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n14863) );
  NOR2_X1 U16581 ( .A1(n14876), .A2(n14863), .ZN(P2_U3283) );
  INV_X1 U16582 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n14864) );
  NOR2_X1 U16583 ( .A1(n14876), .A2(n14864), .ZN(P2_U3284) );
  INV_X1 U16584 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n14865) );
  NOR2_X1 U16585 ( .A1(n14876), .A2(n14865), .ZN(P2_U3285) );
  INV_X1 U16586 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n14866) );
  NOR2_X1 U16587 ( .A1(n14876), .A2(n14866), .ZN(P2_U3286) );
  INV_X1 U16588 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n14867) );
  NOR2_X1 U16589 ( .A1(n14876), .A2(n14867), .ZN(P2_U3287) );
  INV_X1 U16590 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n14868) );
  NOR2_X1 U16591 ( .A1(n14876), .A2(n14868), .ZN(P2_U3288) );
  INV_X1 U16592 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n14869) );
  NOR2_X1 U16593 ( .A1(n14876), .A2(n14869), .ZN(P2_U3289) );
  INV_X1 U16594 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n14870) );
  NOR2_X1 U16595 ( .A1(n14872), .A2(n14870), .ZN(P2_U3290) );
  INV_X1 U16596 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n15554) );
  NOR2_X1 U16597 ( .A1(n14876), .A2(n15554), .ZN(P2_U3291) );
  INV_X1 U16598 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n14871) );
  NOR2_X1 U16599 ( .A1(n14872), .A2(n14871), .ZN(P2_U3292) );
  INV_X1 U16600 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n14873) );
  NOR2_X1 U16601 ( .A1(n14876), .A2(n14873), .ZN(P2_U3293) );
  INV_X1 U16602 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n14874) );
  NOR2_X1 U16603 ( .A1(n14876), .A2(n14874), .ZN(P2_U3294) );
  INV_X1 U16604 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n14875) );
  NOR2_X1 U16605 ( .A1(n14876), .A2(n14875), .ZN(P2_U3295) );
  OAI21_X1 U16606 ( .B1(n14881), .B2(n14878), .A(n14877), .ZN(P2_U3416) );
  AOI22_X1 U16607 ( .A1(n14881), .A2(n14880), .B1(n15552), .B2(n14879), .ZN(
        P2_U3417) );
  AOI22_X1 U16608 ( .A1(n14884), .A2(n14918), .B1(n14883), .B2(n14882), .ZN(
        n14885) );
  AND2_X1 U16609 ( .A1(n14886), .A2(n14885), .ZN(n14926) );
  INV_X1 U16610 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n14887) );
  AOI22_X1 U16611 ( .A1(n14924), .A2(n14926), .B1(n14887), .B2(n14922), .ZN(
        P2_U3430) );
  INV_X1 U16612 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n14888) );
  AOI22_X1 U16613 ( .A1(n14924), .A2(n14889), .B1(n14888), .B2(n14922), .ZN(
        P2_U3433) );
  AOI21_X1 U16614 ( .B1(n14892), .B2(n14891), .A(n14890), .ZN(n14893) );
  OAI21_X1 U16615 ( .B1(n14895), .B2(n14894), .A(n14893), .ZN(n14897) );
  NOR2_X1 U16616 ( .A1(n14897), .A2(n14896), .ZN(n14927) );
  INV_X1 U16617 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n14898) );
  AOI22_X1 U16618 ( .A1(n14924), .A2(n14927), .B1(n14898), .B2(n14922), .ZN(
        P2_U3439) );
  INV_X1 U16619 ( .A(n14899), .ZN(n14906) );
  OAI21_X1 U16620 ( .B1(n14901), .B2(n14915), .A(n14900), .ZN(n14904) );
  INV_X1 U16621 ( .A(n14902), .ZN(n14903) );
  AOI211_X1 U16622 ( .C1(n14906), .C2(n14905), .A(n14904), .B(n14903), .ZN(
        n14929) );
  INV_X1 U16623 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n14907) );
  AOI22_X1 U16624 ( .A1(n14924), .A2(n14929), .B1(n14907), .B2(n14922), .ZN(
        P2_U3445) );
  OAI21_X1 U16625 ( .B1(n14909), .B2(n14915), .A(n14908), .ZN(n14911) );
  AOI211_X1 U16626 ( .C1(n14918), .C2(n14912), .A(n14911), .B(n14910), .ZN(
        n14931) );
  INV_X1 U16627 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n14913) );
  AOI22_X1 U16628 ( .A1(n14924), .A2(n14931), .B1(n14913), .B2(n14922), .ZN(
        P2_U3454) );
  OAI21_X1 U16629 ( .B1(n14916), .B2(n14915), .A(n14914), .ZN(n14917) );
  AOI21_X1 U16630 ( .B1(n14919), .B2(n14918), .A(n14917), .ZN(n14920) );
  AND2_X1 U16631 ( .A1(n14921), .A2(n14920), .ZN(n14933) );
  INV_X1 U16632 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n14923) );
  AOI22_X1 U16633 ( .A1(n14924), .A2(n14933), .B1(n14923), .B2(n14922), .ZN(
        P2_U3460) );
  INV_X1 U16634 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n14925) );
  AOI22_X1 U16635 ( .A1(n14934), .A2(n14926), .B1(n14925), .B2(n14932), .ZN(
        P2_U3499) );
  AOI22_X1 U16636 ( .A1(n14934), .A2(n14927), .B1(n9652), .B2(n14932), .ZN(
        P2_U3502) );
  INV_X1 U16637 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n14928) );
  AOI22_X1 U16638 ( .A1(n14934), .A2(n14929), .B1(n14928), .B2(n14932), .ZN(
        P2_U3504) );
  AOI22_X1 U16639 ( .A1(n14934), .A2(n14931), .B1(n14930), .B2(n14932), .ZN(
        P2_U3507) );
  AOI22_X1 U16640 ( .A1(n14934), .A2(n14933), .B1(n9753), .B2(n14932), .ZN(
        P2_U3509) );
  NOR2_X1 U16641 ( .A1(P3_U3897), .A2(n15025), .ZN(P3_U3150) );
  AOI22_X1 U16642 ( .A1(n14966), .A2(n14936), .B1(n14998), .B2(n14935), .ZN(
        n14943) );
  AOI22_X1 U16643 ( .A1(P3_ADDR_REG_0__SCAN_IN), .A2(n15025), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n14942) );
  NAND3_X1 U16644 ( .A1(n15110), .A2(n15095), .A3(n15082), .ZN(n14938) );
  AOI22_X1 U16645 ( .A1(n14938), .A2(n14937), .B1(P3_IR_REG_0__SCAN_IN), .B2(
        n15016), .ZN(n14941) );
  NAND3_X1 U16646 ( .A1(n15104), .A2(n14939), .A3(n6827), .ZN(n14940) );
  NAND4_X1 U16647 ( .A1(n14943), .A2(n14942), .A3(n14941), .A4(n14940), .ZN(
        P3_U3182) );
  AOI21_X1 U16648 ( .B1(n14946), .B2(n14945), .A(n14944), .ZN(n14950) );
  AOI21_X1 U16649 ( .B1(n14948), .B2(n15566), .A(n14947), .ZN(n14949) );
  OAI22_X1 U16650 ( .A1(n15110), .A2(n14950), .B1(n14949), .B2(n15095), .ZN(
        n14955) );
  XOR2_X1 U16651 ( .A(n14952), .B(n14951), .Z(n14953) );
  NOR2_X1 U16652 ( .A1(n14953), .A2(n15082), .ZN(n14954) );
  AOI211_X1 U16653 ( .C1(n15016), .C2(n14956), .A(n14955), .B(n14954), .ZN(
        n14958) );
  NAND2_X1 U16654 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_U3151), .ZN(n14957) );
  OAI211_X1 U16655 ( .C1(n15493), .C2(n15098), .A(n14958), .B(n14957), .ZN(
        P3_U3185) );
  AOI22_X1 U16656 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n15025), .B1(
        P3_REG3_REG_5__SCAN_IN), .B2(P3_U3151), .ZN(n14971) );
  OAI21_X1 U16657 ( .B1(n14961), .B2(n14960), .A(n14959), .ZN(n14963) );
  AOI22_X1 U16658 ( .A1(n14963), .A2(n15104), .B1(n14962), .B2(n15016), .ZN(
        n14970) );
  OAI221_X1 U16659 ( .B1(n14965), .B2(n10625), .C1(n14965), .C2(n14964), .A(
        n14998), .ZN(n14969) );
  XOR2_X1 U16660 ( .A(n6801), .B(n15191), .Z(n14967) );
  NAND2_X1 U16661 ( .A1(n14967), .A2(n14966), .ZN(n14968) );
  NAND4_X1 U16662 ( .A1(n14971), .A2(n14970), .A3(n14969), .A4(n14968), .ZN(
        P3_U3187) );
  AOI21_X1 U16663 ( .B1(n6690), .B2(n14973), .A(n14972), .ZN(n14985) );
  AOI21_X1 U16664 ( .B1(n14976), .B2(n14975), .A(n14974), .ZN(n14977) );
  OR2_X1 U16665 ( .A1(n14977), .A2(n15110), .ZN(n14984) );
  OAI21_X1 U16666 ( .B1(n14980), .B2(n14979), .A(n14978), .ZN(n14981) );
  AOI22_X1 U16667 ( .A1(n15016), .A2(n14982), .B1(n14981), .B2(n15104), .ZN(
        n14983) );
  OAI211_X1 U16668 ( .C1(n14985), .C2(n15095), .A(n14984), .B(n14983), .ZN(
        n14986) );
  INV_X1 U16669 ( .A(n14986), .ZN(n14988) );
  NAND2_X1 U16670 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P3_U3151), .ZN(n14987) );
  OAI211_X1 U16671 ( .C1(n14989), .C2(n15098), .A(n14988), .B(n14987), .ZN(
        P3_U3188) );
  AOI22_X1 U16672 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n15025), .B1(
        P3_REG3_REG_7__SCAN_IN), .B2(P3_U3151), .ZN(n15005) );
  OAI21_X1 U16673 ( .B1(n14992), .B2(n14991), .A(n14990), .ZN(n14994) );
  AOI22_X1 U16674 ( .A1(n14994), .A2(n15104), .B1(n14993), .B2(n15016), .ZN(
        n15004) );
  AOI21_X1 U16675 ( .B1(n14996), .B2(n15195), .A(n14995), .ZN(n14997) );
  OR2_X1 U16676 ( .A1(n14997), .A2(n15095), .ZN(n15003) );
  OAI221_X1 U16677 ( .B1(n15001), .B2(n15000), .C1(n15001), .C2(n14999), .A(
        n14998), .ZN(n15002) );
  NAND4_X1 U16678 ( .A1(n15005), .A2(n15004), .A3(n15003), .A4(n15002), .ZN(
        P3_U3189) );
  AOI21_X1 U16679 ( .B1(n15008), .B2(n15007), .A(n15006), .ZN(n15019) );
  AOI21_X1 U16680 ( .B1(n6795), .B2(n15010), .A(n15009), .ZN(n15011) );
  OR2_X1 U16681 ( .A1(n15011), .A2(n15110), .ZN(n15018) );
  XNOR2_X1 U16682 ( .A(n15013), .B(n15012), .ZN(n15014) );
  AOI22_X1 U16683 ( .A1(n15016), .A2(n15015), .B1(n15014), .B2(n15104), .ZN(
        n15017) );
  OAI211_X1 U16684 ( .C1(n15019), .C2(n15095), .A(n15018), .B(n15017), .ZN(
        n15020) );
  INV_X1 U16685 ( .A(n15020), .ZN(n15022) );
  NAND2_X1 U16686 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_U3151), .ZN(n15021) );
  OAI211_X1 U16687 ( .C1(n15366), .C2(n15098), .A(n15022), .B(n15021), .ZN(
        P3_U3190) );
  AOI21_X1 U16688 ( .B1(n6794), .B2(n15024), .A(n15023), .ZN(n15037) );
  AOI22_X1 U16689 ( .A1(P3_ADDR_REG_10__SCAN_IN), .A2(n15025), .B1(
        P3_REG3_REG_10__SCAN_IN), .B2(P3_U3151), .ZN(n15036) );
  AOI21_X1 U16690 ( .B1(n15028), .B2(n15027), .A(n15026), .ZN(n15032) );
  AOI21_X1 U16691 ( .B1(n6800), .B2(n15030), .A(n15029), .ZN(n15031) );
  OAI222_X1 U16692 ( .A1(n15101), .A2(n15033), .B1(n15082), .B2(n15032), .C1(
        n15095), .C2(n15031), .ZN(n15034) );
  INV_X1 U16693 ( .A(n15034), .ZN(n15035) );
  OAI211_X1 U16694 ( .C1(n15037), .C2(n15110), .A(n15036), .B(n15035), .ZN(
        P3_U3192) );
  AOI21_X1 U16695 ( .B1(n15329), .B2(n15039), .A(n15038), .ZN(n15053) );
  OAI22_X1 U16696 ( .A1(n15101), .A2(n15041), .B1(n15040), .B2(n15098), .ZN(
        n15051) );
  AOI21_X1 U16697 ( .B1(n15044), .B2(n15043), .A(n15042), .ZN(n15049) );
  AOI21_X1 U16698 ( .B1(n15047), .B2(n15046), .A(n15045), .ZN(n15048) );
  OAI22_X1 U16699 ( .A1(n15049), .A2(n15095), .B1(n15048), .B2(n15082), .ZN(
        n15050) );
  AOI211_X1 U16700 ( .C1(P3_REG3_REG_11__SCAN_IN), .C2(P3_U3151), .A(n15051), 
        .B(n15050), .ZN(n15052) );
  OAI21_X1 U16701 ( .B1(n15053), .B2(n15110), .A(n15052), .ZN(P3_U3193) );
  INV_X1 U16702 ( .A(n15054), .ZN(n15055) );
  AOI21_X1 U16703 ( .B1(n15057), .B2(n15056), .A(n15055), .ZN(n15071) );
  NAND2_X1 U16704 ( .A1(n15059), .A2(n15058), .ZN(n15060) );
  AOI21_X1 U16705 ( .B1(n15061), .B2(n15060), .A(n15095), .ZN(n15065) );
  OAI22_X1 U16706 ( .A1(n15101), .A2(n15063), .B1(n15062), .B2(n15098), .ZN(
        n15064) );
  AOI211_X1 U16707 ( .C1(P3_REG3_REG_12__SCAN_IN), .C2(P3_U3151), .A(n15065), 
        .B(n15064), .ZN(n15070) );
  OAI211_X1 U16708 ( .C1(n15068), .C2(n15067), .A(n15066), .B(n15104), .ZN(
        n15069) );
  OAI211_X1 U16709 ( .C1(n15071), .C2(n15110), .A(n15070), .B(n15069), .ZN(
        P3_U3194) );
  AOI21_X1 U16710 ( .B1(n15557), .B2(n15073), .A(n15072), .ZN(n15088) );
  OAI22_X1 U16711 ( .A1(n15101), .A2(n12468), .B1(n15075), .B2(n15098), .ZN(
        n15086) );
  AOI21_X1 U16712 ( .B1(n15078), .B2(n15077), .A(n15076), .ZN(n15084) );
  AOI21_X1 U16713 ( .B1(n15081), .B2(n15080), .A(n15079), .ZN(n15083) );
  OAI22_X1 U16714 ( .A1(n15084), .A2(n15095), .B1(n15083), .B2(n15082), .ZN(
        n15085) );
  AOI211_X1 U16715 ( .C1(P3_REG3_REG_13__SCAN_IN), .C2(P3_U3151), .A(n15086), 
        .B(n15085), .ZN(n15087) );
  OAI21_X1 U16716 ( .B1(n15088), .B2(n15110), .A(n15087), .ZN(P3_U3195) );
  AOI21_X1 U16717 ( .B1(n15091), .B2(n15090), .A(n15089), .ZN(n15111) );
  INV_X1 U16718 ( .A(n15092), .ZN(n15094) );
  NAND2_X1 U16719 ( .A1(n15094), .A2(n15093), .ZN(n15096) );
  AOI21_X1 U16720 ( .B1(n15097), .B2(n15096), .A(n15095), .ZN(n15103) );
  OAI22_X1 U16721 ( .A1(n15101), .A2(n15100), .B1(n15099), .B2(n15098), .ZN(
        n15102) );
  AOI211_X1 U16722 ( .C1(P3_REG3_REG_14__SCAN_IN), .C2(P3_U3151), .A(n15103), 
        .B(n15102), .ZN(n15109) );
  OAI211_X1 U16723 ( .C1(n15107), .C2(n15106), .A(n15105), .B(n15104), .ZN(
        n15108) );
  OAI211_X1 U16724 ( .C1(n15111), .C2(n15110), .A(n15109), .B(n15108), .ZN(
        P3_U3196) );
  NOR2_X1 U16725 ( .A1(n15112), .A2(n15146), .ZN(n15134) );
  XNOR2_X1 U16726 ( .A(n6960), .B(n15113), .ZN(n15127) );
  OAI21_X1 U16727 ( .B1(n15116), .B2(n6960), .A(n15114), .ZN(n15123) );
  OAI22_X1 U16728 ( .A1(n15120), .A2(n15119), .B1(n15118), .B2(n15117), .ZN(
        n15121) );
  AOI21_X1 U16729 ( .B1(n15123), .B2(n15122), .A(n15121), .ZN(n15124) );
  OAI21_X1 U16730 ( .B1(n15127), .B2(n15125), .A(n15124), .ZN(n15133) );
  AOI21_X1 U16731 ( .B1(n15134), .B2(n15126), .A(n15133), .ZN(n15132) );
  INV_X1 U16732 ( .A(n15127), .ZN(n15135) );
  AOI22_X1 U16733 ( .A1(n15135), .A2(n15128), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n15591), .ZN(n15129) );
  OAI221_X1 U16734 ( .B1(n15595), .B2(n15132), .C1(n15131), .C2(n15130), .A(
        n15129), .ZN(P3_U3232) );
  INV_X1 U16735 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15136) );
  AOI211_X1 U16736 ( .C1(n15179), .C2(n15135), .A(n15134), .B(n15133), .ZN(
        n15185) );
  AOI22_X1 U16737 ( .A1(n15183), .A2(n15136), .B1(n15185), .B2(n15181), .ZN(
        P3_U3393) );
  INV_X1 U16738 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15141) );
  INV_X1 U16739 ( .A(n15137), .ZN(n15138) );
  AOI211_X1 U16740 ( .C1(n15179), .C2(n15140), .A(n15139), .B(n15138), .ZN(
        n15187) );
  AOI22_X1 U16741 ( .A1(n15183), .A2(n15141), .B1(n15187), .B2(n15181), .ZN(
        P3_U3396) );
  INV_X1 U16742 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15145) );
  AOI211_X1 U16743 ( .C1(n15144), .C2(n15179), .A(n15143), .B(n15142), .ZN(
        n15188) );
  AOI22_X1 U16744 ( .A1(n15183), .A2(n15145), .B1(n15188), .B2(n15181), .ZN(
        P3_U3399) );
  INV_X1 U16745 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15151) );
  NOR2_X1 U16746 ( .A1(n15147), .A2(n15146), .ZN(n15149) );
  AOI211_X1 U16747 ( .C1(n15179), .C2(n15150), .A(n15149), .B(n15148), .ZN(
        n15190) );
  AOI22_X1 U16748 ( .A1(n15183), .A2(n15151), .B1(n15190), .B2(n15181), .ZN(
        P3_U3402) );
  INV_X1 U16749 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15555) );
  INV_X1 U16750 ( .A(n15152), .ZN(n15153) );
  AOI211_X1 U16751 ( .C1(n15155), .C2(n15179), .A(n15154), .B(n15153), .ZN(
        n15192) );
  AOI22_X1 U16752 ( .A1(n15183), .A2(n15555), .B1(n15192), .B2(n15181), .ZN(
        P3_U3405) );
  INV_X1 U16753 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15161) );
  AOI22_X1 U16754 ( .A1(n15158), .A2(n15179), .B1(n15157), .B2(n15156), .ZN(
        n15159) );
  AND2_X1 U16755 ( .A1(n15160), .A2(n15159), .ZN(n15194) );
  AOI22_X1 U16756 ( .A1(n15183), .A2(n15161), .B1(n15194), .B2(n15181), .ZN(
        P3_U3408) );
  INV_X1 U16757 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15165) );
  AOI211_X1 U16758 ( .C1(n15179), .C2(n15164), .A(n15163), .B(n15162), .ZN(
        n15196) );
  AOI22_X1 U16759 ( .A1(n15183), .A2(n15165), .B1(n15196), .B2(n15181), .ZN(
        P3_U3411) );
  INV_X1 U16760 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15170) );
  INV_X1 U16761 ( .A(n15166), .ZN(n15167) );
  AOI211_X1 U16762 ( .C1(n15169), .C2(n15179), .A(n15168), .B(n15167), .ZN(
        n15198) );
  AOI22_X1 U16763 ( .A1(n15183), .A2(n15170), .B1(n15198), .B2(n15181), .ZN(
        P3_U3414) );
  INV_X1 U16764 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15175) );
  INV_X1 U16765 ( .A(n15171), .ZN(n15174) );
  AOI211_X1 U16766 ( .C1(n15174), .C2(n15179), .A(n15173), .B(n15172), .ZN(
        n15200) );
  AOI22_X1 U16767 ( .A1(n15183), .A2(n15175), .B1(n15200), .B2(n15181), .ZN(
        P3_U3417) );
  INV_X1 U16768 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15182) );
  INV_X1 U16769 ( .A(n15176), .ZN(n15180) );
  AOI211_X1 U16770 ( .C1(n15180), .C2(n15179), .A(n15178), .B(n15177), .ZN(
        n15201) );
  AOI22_X1 U16771 ( .A1(n15183), .A2(n15182), .B1(n15201), .B2(n15181), .ZN(
        P3_U3420) );
  INV_X1 U16772 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n15184) );
  AOI22_X1 U16773 ( .A1(n15202), .A2(n15185), .B1(n15184), .B2(n8976), .ZN(
        P3_U3460) );
  AOI22_X1 U16774 ( .A1(n15202), .A2(n15187), .B1(n15186), .B2(n8976), .ZN(
        P3_U3461) );
  AOI22_X1 U16775 ( .A1(n15202), .A2(n15188), .B1(n15566), .B2(n8976), .ZN(
        P3_U3462) );
  AOI22_X1 U16776 ( .A1(n15202), .A2(n15190), .B1(n15189), .B2(n8976), .ZN(
        P3_U3463) );
  AOI22_X1 U16777 ( .A1(n15202), .A2(n15192), .B1(n15191), .B2(n8976), .ZN(
        P3_U3464) );
  AOI22_X1 U16778 ( .A1(n15202), .A2(n15194), .B1(n15193), .B2(n8976), .ZN(
        P3_U3465) );
  AOI22_X1 U16779 ( .A1(n15202), .A2(n15196), .B1(n15195), .B2(n8976), .ZN(
        P3_U3466) );
  AOI22_X1 U16780 ( .A1(n15202), .A2(n15198), .B1(n15197), .B2(n8976), .ZN(
        P3_U3467) );
  AOI22_X1 U16781 ( .A1(n15202), .A2(n15200), .B1(n15199), .B2(n8976), .ZN(
        P3_U3468) );
  AOI22_X1 U16782 ( .A1(n15202), .A2(n15201), .B1(n12428), .B2(n8976), .ZN(
        P3_U3469) );
  AOI22_X1 U16783 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(keyinput228), .B1(
        P3_D_REG_2__SCAN_IN), .B2(keyinput245), .ZN(n15203) );
  OAI221_X1 U16784 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(keyinput228), .C1(
        P3_D_REG_2__SCAN_IN), .C2(keyinput245), .A(n15203), .ZN(n15210) );
  AOI22_X1 U16785 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(keyinput201), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(keyinput165), .ZN(n15204) );
  OAI221_X1 U16786 ( .B1(P1_REG3_REG_10__SCAN_IN), .B2(keyinput201), .C1(
        P2_DATAO_REG_20__SCAN_IN), .C2(keyinput165), .A(n15204), .ZN(n15209)
         );
  AOI22_X1 U16787 ( .A1(P1_D_REG_17__SCAN_IN), .A2(keyinput227), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(keyinput219), .ZN(n15205) );
  OAI221_X1 U16788 ( .B1(P1_D_REG_17__SCAN_IN), .B2(keyinput227), .C1(
        P1_DATAO_REG_19__SCAN_IN), .C2(keyinput219), .A(n15205), .ZN(n15208)
         );
  AOI22_X1 U16789 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(keyinput237), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(keyinput139), .ZN(n15206) );
  OAI221_X1 U16790 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(keyinput237), .C1(
        P2_REG3_REG_0__SCAN_IN), .C2(keyinput139), .A(n15206), .ZN(n15207) );
  NOR4_X1 U16791 ( .A1(n15210), .A2(n15209), .A3(n15208), .A4(n15207), .ZN(
        n15238) );
  AOI22_X1 U16792 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(keyinput217), .B1(SI_26_), .B2(keyinput200), .ZN(n15211) );
  OAI221_X1 U16793 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(keyinput217), .C1(
        SI_26_), .C2(keyinput200), .A(n15211), .ZN(n15218) );
  AOI22_X1 U16794 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(keyinput252), .B1(
        P2_IR_REG_23__SCAN_IN), .B2(keyinput173), .ZN(n15212) );
  OAI221_X1 U16795 ( .B1(P2_REG1_REG_18__SCAN_IN), .B2(keyinput252), .C1(
        P2_IR_REG_23__SCAN_IN), .C2(keyinput173), .A(n15212), .ZN(n15217) );
  AOI22_X1 U16796 ( .A1(P2_D_REG_15__SCAN_IN), .A2(keyinput159), .B1(
        P3_IR_REG_22__SCAN_IN), .B2(keyinput185), .ZN(n15213) );
  OAI221_X1 U16797 ( .B1(P2_D_REG_15__SCAN_IN), .B2(keyinput159), .C1(
        P3_IR_REG_22__SCAN_IN), .C2(keyinput185), .A(n15213), .ZN(n15216) );
  AOI22_X1 U16798 ( .A1(P2_D_REG_31__SCAN_IN), .A2(keyinput176), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(keyinput150), .ZN(n15214) );
  OAI221_X1 U16799 ( .B1(P2_D_REG_31__SCAN_IN), .B2(keyinput176), .C1(
        P2_DATAO_REG_15__SCAN_IN), .C2(keyinput150), .A(n15214), .ZN(n15215)
         );
  NOR4_X1 U16800 ( .A1(n15218), .A2(n15217), .A3(n15216), .A4(n15215), .ZN(
        n15237) );
  AOI22_X1 U16801 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(keyinput178), .B1(
        P3_D_REG_1__SCAN_IN), .B2(keyinput229), .ZN(n15219) );
  OAI221_X1 U16802 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(keyinput178), .C1(
        P3_D_REG_1__SCAN_IN), .C2(keyinput229), .A(n15219), .ZN(n15226) );
  AOI22_X1 U16803 ( .A1(P3_DATAO_REG_24__SCAN_IN), .A2(keyinput255), .B1(
        P2_REG2_REG_7__SCAN_IN), .B2(keyinput164), .ZN(n15220) );
  OAI221_X1 U16804 ( .B1(P3_DATAO_REG_24__SCAN_IN), .B2(keyinput255), .C1(
        P2_REG2_REG_7__SCAN_IN), .C2(keyinput164), .A(n15220), .ZN(n15225) );
  AOI22_X1 U16805 ( .A1(P3_REG1_REG_3__SCAN_IN), .A2(keyinput130), .B1(
        P3_D_REG_17__SCAN_IN), .B2(keyinput207), .ZN(n15221) );
  OAI221_X1 U16806 ( .B1(P3_REG1_REG_3__SCAN_IN), .B2(keyinput130), .C1(
        P3_D_REG_17__SCAN_IN), .C2(keyinput207), .A(n15221), .ZN(n15224) );
  AOI22_X1 U16807 ( .A1(P3_DATAO_REG_29__SCAN_IN), .A2(keyinput149), .B1(
        P2_WR_REG_SCAN_IN), .B2(keyinput187), .ZN(n15222) );
  OAI221_X1 U16808 ( .B1(P3_DATAO_REG_29__SCAN_IN), .B2(keyinput149), .C1(
        P2_WR_REG_SCAN_IN), .C2(keyinput187), .A(n15222), .ZN(n15223) );
  NOR4_X1 U16809 ( .A1(n15226), .A2(n15225), .A3(n15224), .A4(n15223), .ZN(
        n15236) );
  AOI22_X1 U16810 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(keyinput166), .B1(
        P2_D_REG_29__SCAN_IN), .B2(keyinput158), .ZN(n15227) );
  OAI221_X1 U16811 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(keyinput166), .C1(
        P2_D_REG_29__SCAN_IN), .C2(keyinput158), .A(n15227), .ZN(n15234) );
  AOI22_X1 U16812 ( .A1(P3_REG2_REG_27__SCAN_IN), .A2(keyinput218), .B1(
        P3_D_REG_25__SCAN_IN), .B2(keyinput135), .ZN(n15228) );
  OAI221_X1 U16813 ( .B1(P3_REG2_REG_27__SCAN_IN), .B2(keyinput218), .C1(
        P3_D_REG_25__SCAN_IN), .C2(keyinput135), .A(n15228), .ZN(n15233) );
  AOI22_X1 U16814 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(keyinput195), .B1(
        P1_IR_REG_3__SCAN_IN), .B2(keyinput157), .ZN(n15229) );
  OAI221_X1 U16815 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(keyinput195), .C1(
        P1_IR_REG_3__SCAN_IN), .C2(keyinput157), .A(n15229), .ZN(n15232) );
  AOI22_X1 U16816 ( .A1(P1_REG1_REG_24__SCAN_IN), .A2(keyinput193), .B1(
        P2_D_REG_30__SCAN_IN), .B2(keyinput239), .ZN(n15230) );
  OAI221_X1 U16817 ( .B1(P1_REG1_REG_24__SCAN_IN), .B2(keyinput193), .C1(
        P2_D_REG_30__SCAN_IN), .C2(keyinput239), .A(n15230), .ZN(n15231) );
  NOR4_X1 U16818 ( .A1(n15234), .A2(n15233), .A3(n15232), .A4(n15231), .ZN(
        n15235) );
  NAND4_X1 U16819 ( .A1(n15238), .A2(n15237), .A3(n15236), .A4(n15235), .ZN(
        n15382) );
  AOI22_X1 U16820 ( .A1(P3_DATAO_REG_25__SCAN_IN), .A2(keyinput137), .B1(
        P2_REG0_REG_6__SCAN_IN), .B2(keyinput240), .ZN(n15239) );
  OAI221_X1 U16821 ( .B1(P3_DATAO_REG_25__SCAN_IN), .B2(keyinput137), .C1(
        P2_REG0_REG_6__SCAN_IN), .C2(keyinput240), .A(n15239), .ZN(n15246) );
  AOI22_X1 U16822 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(keyinput206), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(keyinput212), .ZN(n15240) );
  OAI221_X1 U16823 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(keyinput206), .C1(
        P2_DATAO_REG_24__SCAN_IN), .C2(keyinput212), .A(n15240), .ZN(n15245)
         );
  AOI22_X1 U16824 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(keyinput251), .B1(
        P2_REG0_REG_28__SCAN_IN), .B2(keyinput197), .ZN(n15241) );
  OAI221_X1 U16825 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(keyinput251), .C1(
        P2_REG0_REG_28__SCAN_IN), .C2(keyinput197), .A(n15241), .ZN(n15244) );
  AOI22_X1 U16826 ( .A1(P2_D_REG_1__SCAN_IN), .A2(keyinput177), .B1(
        P3_REG2_REG_23__SCAN_IN), .B2(keyinput191), .ZN(n15242) );
  OAI221_X1 U16827 ( .B1(P2_D_REG_1__SCAN_IN), .B2(keyinput177), .C1(
        P3_REG2_REG_23__SCAN_IN), .C2(keyinput191), .A(n15242), .ZN(n15243) );
  NOR4_X1 U16828 ( .A1(n15246), .A2(n15245), .A3(n15244), .A4(n15243), .ZN(
        n15275) );
  AOI22_X1 U16829 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(keyinput171), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(keyinput225), .ZN(n15247) );
  OAI221_X1 U16830 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(keyinput171), .C1(
        P2_DATAO_REG_17__SCAN_IN), .C2(keyinput225), .A(n15247), .ZN(n15254)
         );
  AOI22_X1 U16831 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(keyinput144), .B1(
        P1_IR_REG_20__SCAN_IN), .B2(keyinput128), .ZN(n15248) );
  OAI221_X1 U16832 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(keyinput144), .C1(
        P1_IR_REG_20__SCAN_IN), .C2(keyinput128), .A(n15248), .ZN(n15253) );
  AOI22_X1 U16833 ( .A1(P2_REG2_REG_21__SCAN_IN), .A2(keyinput155), .B1(
        P3_REG0_REG_21__SCAN_IN), .B2(keyinput162), .ZN(n15249) );
  OAI221_X1 U16834 ( .B1(P2_REG2_REG_21__SCAN_IN), .B2(keyinput155), .C1(
        P3_REG0_REG_21__SCAN_IN), .C2(keyinput162), .A(n15249), .ZN(n15252) );
  AOI22_X1 U16835 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(keyinput133), .B1(
        P3_IR_REG_2__SCAN_IN), .B2(keyinput249), .ZN(n15250) );
  OAI221_X1 U16836 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(keyinput133), .C1(
        P3_IR_REG_2__SCAN_IN), .C2(keyinput249), .A(n15250), .ZN(n15251) );
  NOR4_X1 U16837 ( .A1(n15254), .A2(n15253), .A3(n15252), .A4(n15251), .ZN(
        n15274) );
  AOI22_X1 U16838 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(keyinput142), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(keyinput241), .ZN(n15255) );
  OAI221_X1 U16839 ( .B1(P1_IR_REG_28__SCAN_IN), .B2(keyinput142), .C1(
        P3_REG3_REG_1__SCAN_IN), .C2(keyinput241), .A(n15255), .ZN(n15262) );
  AOI22_X1 U16840 ( .A1(P1_D_REG_30__SCAN_IN), .A2(keyinput175), .B1(
        P3_D_REG_15__SCAN_IN), .B2(keyinput132), .ZN(n15256) );
  OAI221_X1 U16841 ( .B1(P1_D_REG_30__SCAN_IN), .B2(keyinput175), .C1(
        P3_D_REG_15__SCAN_IN), .C2(keyinput132), .A(n15256), .ZN(n15261) );
  AOI22_X1 U16842 ( .A1(SI_12_), .A2(keyinput188), .B1(P3_IR_REG_15__SCAN_IN), 
        .B2(keyinput209), .ZN(n15257) );
  OAI221_X1 U16843 ( .B1(SI_12_), .B2(keyinput188), .C1(P3_IR_REG_15__SCAN_IN), 
        .C2(keyinput209), .A(n15257), .ZN(n15260) );
  AOI22_X1 U16844 ( .A1(P1_REG1_REG_17__SCAN_IN), .A2(keyinput180), .B1(
        P3_REG2_REG_18__SCAN_IN), .B2(keyinput168), .ZN(n15258) );
  OAI221_X1 U16845 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(keyinput180), .C1(
        P3_REG2_REG_18__SCAN_IN), .C2(keyinput168), .A(n15258), .ZN(n15259) );
  NOR4_X1 U16846 ( .A1(n15262), .A2(n15261), .A3(n15260), .A4(n15259), .ZN(
        n15273) );
  AOI22_X1 U16847 ( .A1(n15554), .A2(keyinput131), .B1(keyinput181), .B2(
        n15462), .ZN(n15263) );
  OAI221_X1 U16848 ( .B1(n15554), .B2(keyinput131), .C1(n15462), .C2(
        keyinput181), .A(n15263), .ZN(n15271) );
  AOI22_X1 U16849 ( .A1(P3_REG0_REG_12__SCAN_IN), .A2(keyinput223), .B1(
        P3_IR_REG_8__SCAN_IN), .B2(keyinput186), .ZN(n15264) );
  OAI221_X1 U16850 ( .B1(P3_REG0_REG_12__SCAN_IN), .B2(keyinput223), .C1(
        P3_IR_REG_8__SCAN_IN), .C2(keyinput186), .A(n15264), .ZN(n15270) );
  XNOR2_X1 U16851 ( .A(P1_REG3_REG_2__SCAN_IN), .B(keyinput174), .ZN(n15268)
         );
  XNOR2_X1 U16852 ( .A(P3_REG1_REG_24__SCAN_IN), .B(keyinput136), .ZN(n15267)
         );
  XNOR2_X1 U16853 ( .A(P2_REG1_REG_24__SCAN_IN), .B(keyinput160), .ZN(n15266)
         );
  XNOR2_X1 U16854 ( .A(P2_IR_REG_10__SCAN_IN), .B(keyinput246), .ZN(n15265) );
  NAND4_X1 U16855 ( .A1(n15268), .A2(n15267), .A3(n15266), .A4(n15265), .ZN(
        n15269) );
  NOR3_X1 U16856 ( .A1(n15271), .A2(n15270), .A3(n15269), .ZN(n15272) );
  NAND4_X1 U16857 ( .A1(n15275), .A2(n15274), .A3(n15273), .A4(n15272), .ZN(
        n15381) );
  AOI22_X1 U16858 ( .A1(n15432), .A2(keyinput248), .B1(keyinput204), .B2(
        n10905), .ZN(n15276) );
  OAI221_X1 U16859 ( .B1(n15432), .B2(keyinput248), .C1(n10905), .C2(
        keyinput204), .A(n15276), .ZN(n15280) );
  INV_X1 U16860 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n15431) );
  AOI22_X1 U16861 ( .A1(n15401), .A2(keyinput138), .B1(n15431), .B2(
        keyinput134), .ZN(n15277) );
  OAI221_X1 U16862 ( .B1(n15401), .B2(keyinput138), .C1(n15431), .C2(
        keyinput134), .A(n15277), .ZN(n15279) );
  XOR2_X1 U16863 ( .A(P2_IR_REG_4__SCAN_IN), .B(keyinput224), .Z(n15278) );
  OR3_X1 U16864 ( .A1(n15280), .A2(n15279), .A3(n15278), .ZN(n15286) );
  AOI22_X1 U16865 ( .A1(n15429), .A2(keyinput222), .B1(keyinput148), .B2(
        n15282), .ZN(n15281) );
  OAI221_X1 U16866 ( .B1(n15429), .B2(keyinput222), .C1(n15282), .C2(
        keyinput148), .A(n15281), .ZN(n15285) );
  XNOR2_X1 U16867 ( .A(n15283), .B(keyinput216), .ZN(n15284) );
  NOR3_X1 U16868 ( .A1(n15286), .A2(n15285), .A3(n15284), .ZN(n15325) );
  AOI22_X1 U16869 ( .A1(n15288), .A2(keyinput147), .B1(keyinput170), .B2(
        n12428), .ZN(n15287) );
  OAI221_X1 U16870 ( .B1(n15288), .B2(keyinput147), .C1(n12428), .C2(
        keyinput170), .A(n15287), .ZN(n15298) );
  INV_X1 U16871 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n15290) );
  AOI22_X1 U16872 ( .A1(n15450), .A2(keyinput231), .B1(n15290), .B2(
        keyinput129), .ZN(n15289) );
  OAI221_X1 U16873 ( .B1(n15450), .B2(keyinput231), .C1(n15290), .C2(
        keyinput129), .A(n15289), .ZN(n15297) );
  INV_X1 U16874 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n15292) );
  AOI22_X1 U16875 ( .A1(n15428), .A2(keyinput236), .B1(keyinput211), .B2(
        n15292), .ZN(n15291) );
  OAI221_X1 U16876 ( .B1(n15428), .B2(keyinput236), .C1(n15292), .C2(
        keyinput211), .A(n15291), .ZN(n15296) );
  XOR2_X1 U16877 ( .A(n7794), .B(keyinput172), .Z(n15294) );
  XNOR2_X1 U16878 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput250), .ZN(n15293) );
  NAND2_X1 U16879 ( .A1(n15294), .A2(n15293), .ZN(n15295) );
  NOR4_X1 U16880 ( .A1(n15298), .A2(n15297), .A3(n15296), .A4(n15295), .ZN(
        n15324) );
  INV_X1 U16881 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n15300) );
  AOI22_X1 U16882 ( .A1(n15300), .A2(keyinput230), .B1(n15487), .B2(
        keyinput220), .ZN(n15299) );
  OAI221_X1 U16883 ( .B1(n15300), .B2(keyinput230), .C1(n15487), .C2(
        keyinput220), .A(n15299), .ZN(n15308) );
  INV_X1 U16884 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n15389) );
  AOI22_X1 U16885 ( .A1(n15389), .A2(keyinput226), .B1(keyinput169), .B2(
        n15402), .ZN(n15301) );
  OAI221_X1 U16886 ( .B1(n15389), .B2(keyinput226), .C1(n15402), .C2(
        keyinput169), .A(n15301), .ZN(n15307) );
  INV_X1 U16887 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n15384) );
  INV_X1 U16888 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n15413) );
  AOI22_X1 U16889 ( .A1(n15384), .A2(keyinput221), .B1(n15413), .B2(
        keyinput146), .ZN(n15302) );
  OAI221_X1 U16890 ( .B1(n15384), .B2(keyinput221), .C1(n15413), .C2(
        keyinput146), .A(n15302), .ZN(n15306) );
  INV_X1 U16891 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n15472) );
  AOI22_X1 U16892 ( .A1(n15472), .A2(keyinput210), .B1(n15304), .B2(
        keyinput199), .ZN(n15303) );
  OAI221_X1 U16893 ( .B1(n15472), .B2(keyinput210), .C1(n15304), .C2(
        keyinput199), .A(n15303), .ZN(n15305) );
  NOR4_X1 U16894 ( .A1(n15308), .A2(n15307), .A3(n15306), .A4(n15305), .ZN(
        n15323) );
  AOI22_X1 U16895 ( .A1(n15311), .A2(keyinput213), .B1(keyinput161), .B2(
        n15310), .ZN(n15309) );
  OAI221_X1 U16896 ( .B1(n15311), .B2(keyinput213), .C1(n15310), .C2(
        keyinput161), .A(n15309), .ZN(n15321) );
  AOI22_X1 U16897 ( .A1(n15313), .A2(keyinput167), .B1(keyinput247), .B2(
        n15555), .ZN(n15312) );
  OAI221_X1 U16898 ( .B1(n15313), .B2(keyinput167), .C1(n15555), .C2(
        keyinput247), .A(n15312), .ZN(n15320) );
  AOI22_X1 U16899 ( .A1(n15315), .A2(keyinput163), .B1(keyinput243), .B2(n8216), .ZN(n15314) );
  OAI221_X1 U16900 ( .B1(n15315), .B2(keyinput163), .C1(n8216), .C2(
        keyinput243), .A(n15314), .ZN(n15319) );
  XNOR2_X1 U16901 ( .A(P3_IR_REG_12__SCAN_IN), .B(keyinput235), .ZN(n15317) );
  XNOR2_X1 U16902 ( .A(P2_REG0_REG_21__SCAN_IN), .B(keyinput153), .ZN(n15316)
         );
  NAND2_X1 U16903 ( .A1(n15317), .A2(n15316), .ZN(n15318) );
  NOR4_X1 U16904 ( .A1(n15321), .A2(n15320), .A3(n15319), .A4(n15318), .ZN(
        n15322) );
  NAND4_X1 U16905 ( .A1(n15325), .A2(n15324), .A3(n15323), .A4(n15322), .ZN(
        n15380) );
  AOI22_X1 U16906 ( .A1(n15399), .A2(keyinput184), .B1(keyinput253), .B2(
        n15327), .ZN(n15326) );
  OAI221_X1 U16907 ( .B1(n15399), .B2(keyinput184), .C1(n15327), .C2(
        keyinput253), .A(n15326), .ZN(n15338) );
  AOI22_X1 U16908 ( .A1(n15330), .A2(keyinput202), .B1(keyinput238), .B2(
        n15329), .ZN(n15328) );
  OAI221_X1 U16909 ( .B1(n15330), .B2(keyinput202), .C1(n15329), .C2(
        keyinput238), .A(n15328), .ZN(n15337) );
  AOI22_X1 U16910 ( .A1(n15449), .A2(keyinput145), .B1(n15332), .B2(
        keyinput189), .ZN(n15331) );
  OAI221_X1 U16911 ( .B1(n15449), .B2(keyinput145), .C1(n15332), .C2(
        keyinput189), .A(n15331), .ZN(n15336) );
  XNOR2_X1 U16912 ( .A(P3_REG1_REG_31__SCAN_IN), .B(keyinput152), .ZN(n15334)
         );
  XNOR2_X1 U16913 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(keyinput154), .ZN(n15333)
         );
  NAND2_X1 U16914 ( .A1(n15334), .A2(n15333), .ZN(n15335) );
  NOR4_X1 U16915 ( .A1(n15338), .A2(n15337), .A3(n15336), .A4(n15335), .ZN(
        n15378) );
  AOI22_X1 U16916 ( .A1(n15404), .A2(keyinput194), .B1(keyinput214), .B2(
        n15340), .ZN(n15339) );
  OAI221_X1 U16917 ( .B1(n15404), .B2(keyinput194), .C1(n15340), .C2(
        keyinput214), .A(n15339), .ZN(n15345) );
  XNOR2_X1 U16918 ( .A(n15341), .B(keyinput205), .ZN(n15344) );
  XNOR2_X1 U16919 ( .A(n15342), .B(keyinput183), .ZN(n15343) );
  OR3_X1 U16920 ( .A1(n15345), .A2(n15344), .A3(n15343), .ZN(n15353) );
  AOI22_X1 U16921 ( .A1(n15387), .A2(keyinput232), .B1(keyinput190), .B2(
        n15347), .ZN(n15346) );
  OAI221_X1 U16922 ( .B1(n15387), .B2(keyinput232), .C1(n15347), .C2(
        keyinput190), .A(n15346), .ZN(n15352) );
  AOI22_X1 U16923 ( .A1(n15350), .A2(keyinput242), .B1(n15349), .B2(
        keyinput140), .ZN(n15348) );
  OAI221_X1 U16924 ( .B1(n15350), .B2(keyinput242), .C1(n15349), .C2(
        keyinput140), .A(n15348), .ZN(n15351) );
  NOR3_X1 U16925 ( .A1(n15353), .A2(n15352), .A3(n15351), .ZN(n15377) );
  AOI22_X1 U16926 ( .A1(n15355), .A2(keyinput234), .B1(keyinput182), .B2(
        n15493), .ZN(n15354) );
  OAI221_X1 U16927 ( .B1(n15355), .B2(keyinput234), .C1(n15493), .C2(
        keyinput182), .A(n15354), .ZN(n15363) );
  INV_X1 U16928 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n15475) );
  AOI22_X1 U16929 ( .A1(n15447), .A2(keyinput141), .B1(n15475), .B2(
        keyinput208), .ZN(n15356) );
  OAI221_X1 U16930 ( .B1(n15447), .B2(keyinput141), .C1(n15475), .C2(
        keyinput208), .A(n15356), .ZN(n15362) );
  XOR2_X1 U16931 ( .A(n15557), .B(keyinput179), .Z(n15360) );
  XNOR2_X1 U16932 ( .A(P2_IR_REG_21__SCAN_IN), .B(keyinput143), .ZN(n15359) );
  XNOR2_X1 U16933 ( .A(P2_IR_REG_19__SCAN_IN), .B(keyinput203), .ZN(n15358) );
  XNOR2_X1 U16934 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(keyinput192), .ZN(n15357)
         );
  NAND4_X1 U16935 ( .A1(n15360), .A2(n15359), .A3(n15358), .A4(n15357), .ZN(
        n15361) );
  NOR3_X1 U16936 ( .A1(n15363), .A2(n15362), .A3(n15361), .ZN(n15376) );
  AOI22_X1 U16937 ( .A1(n11087), .A2(keyinput198), .B1(n15458), .B2(
        keyinput156), .ZN(n15364) );
  OAI221_X1 U16938 ( .B1(n11087), .B2(keyinput198), .C1(n15458), .C2(
        keyinput156), .A(n15364), .ZN(n15374) );
  AOI22_X1 U16939 ( .A1(n15366), .A2(keyinput196), .B1(n10134), .B2(
        keyinput254), .ZN(n15365) );
  OAI221_X1 U16940 ( .B1(n15366), .B2(keyinput196), .C1(n10134), .C2(
        keyinput254), .A(n15365), .ZN(n15373) );
  INV_X1 U16941 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n15368) );
  AOI22_X1 U16942 ( .A1(n15368), .A2(keyinput215), .B1(n8361), .B2(keyinput151), .ZN(n15367) );
  OAI221_X1 U16943 ( .B1(n15368), .B2(keyinput215), .C1(n8361), .C2(
        keyinput151), .A(n15367), .ZN(n15372) );
  XNOR2_X1 U16944 ( .A(P3_REG1_REG_25__SCAN_IN), .B(keyinput244), .ZN(n15370)
         );
  XNOR2_X1 U16945 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput233), .ZN(n15369) );
  NAND2_X1 U16946 ( .A1(n15370), .A2(n15369), .ZN(n15371) );
  NOR4_X1 U16947 ( .A1(n15374), .A2(n15373), .A3(n15372), .A4(n15371), .ZN(
        n15375) );
  NAND4_X1 U16948 ( .A1(n15378), .A2(n15377), .A3(n15376), .A4(n15375), .ZN(
        n15379) );
  NOR4_X1 U16949 ( .A1(n15382), .A2(n15381), .A3(n15380), .A4(n15379), .ZN(
        n15589) );
  AOI22_X1 U16950 ( .A1(n15385), .A2(keyinput50), .B1(keyinput93), .B2(n15384), 
        .ZN(n15383) );
  OAI221_X1 U16951 ( .B1(n15385), .B2(keyinput50), .C1(n15384), .C2(keyinput93), .A(n15383), .ZN(n15396) );
  AOI22_X1 U16952 ( .A1(n15387), .A2(keyinput104), .B1(keyinput23), .B2(n8361), 
        .ZN(n15386) );
  OAI221_X1 U16953 ( .B1(n15387), .B2(keyinput104), .C1(n8361), .C2(keyinput23), .A(n15386), .ZN(n15395) );
  AOI22_X1 U16954 ( .A1(n15390), .A2(keyinput21), .B1(n15389), .B2(keyinput98), 
        .ZN(n15388) );
  OAI221_X1 U16955 ( .B1(n15390), .B2(keyinput21), .C1(n15389), .C2(keyinput98), .A(n15388), .ZN(n15394) );
  XNOR2_X1 U16956 ( .A(P1_REG3_REG_2__SCAN_IN), .B(keyinput46), .ZN(n15392) );
  XNOR2_X1 U16957 ( .A(P1_REG0_REG_22__SCAN_IN), .B(keyinput102), .ZN(n15391)
         );
  NAND2_X1 U16958 ( .A1(n15392), .A2(n15391), .ZN(n15393) );
  NOR4_X1 U16959 ( .A1(n15396), .A2(n15395), .A3(n15394), .A4(n15393), .ZN(
        n15442) );
  AOI22_X1 U16960 ( .A1(n15399), .A2(keyinput56), .B1(n15398), .B2(keyinput90), 
        .ZN(n15397) );
  OAI221_X1 U16961 ( .B1(n15399), .B2(keyinput56), .C1(n15398), .C2(keyinput90), .A(n15397), .ZN(n15411) );
  AOI22_X1 U16962 ( .A1(n15402), .A2(keyinput41), .B1(n15401), .B2(keyinput10), 
        .ZN(n15400) );
  OAI221_X1 U16963 ( .B1(n15402), .B2(keyinput41), .C1(n15401), .C2(keyinput10), .A(n15400), .ZN(n15410) );
  AOI22_X1 U16964 ( .A1(n15405), .A2(keyinput100), .B1(n15404), .B2(keyinput66), .ZN(n15403) );
  OAI221_X1 U16965 ( .B1(n15405), .B2(keyinput100), .C1(n15404), .C2(
        keyinput66), .A(n15403), .ZN(n15409) );
  AOI22_X1 U16966 ( .A1(n15407), .A2(keyinput9), .B1(n8495), .B2(keyinput101), 
        .ZN(n15406) );
  OAI221_X1 U16967 ( .B1(n15407), .B2(keyinput9), .C1(n8495), .C2(keyinput101), 
        .A(n15406), .ZN(n15408) );
  NOR4_X1 U16968 ( .A1(n15411), .A2(n15410), .A3(n15409), .A4(n15408), .ZN(
        n15441) );
  AOI22_X1 U16969 ( .A1(n15414), .A2(keyinput109), .B1(n15413), .B2(keyinput18), .ZN(n15412) );
  OAI221_X1 U16970 ( .B1(n15414), .B2(keyinput109), .C1(n15413), .C2(
        keyinput18), .A(n15412), .ZN(n15424) );
  INV_X1 U16971 ( .A(P2_WR_REG_SCAN_IN), .ZN(n15417) );
  AOI22_X1 U16972 ( .A1(n15417), .A2(keyinput59), .B1(n15416), .B2(keyinput99), 
        .ZN(n15415) );
  OAI221_X1 U16973 ( .B1(n15417), .B2(keyinput59), .C1(n15416), .C2(keyinput99), .A(n15415), .ZN(n15423) );
  XNOR2_X1 U16974 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput0), .ZN(n15421) );
  XNOR2_X1 U16975 ( .A(P3_REG1_REG_25__SCAN_IN), .B(keyinput116), .ZN(n15420)
         );
  XNOR2_X1 U16976 ( .A(P2_IR_REG_19__SCAN_IN), .B(keyinput75), .ZN(n15419) );
  XNOR2_X1 U16977 ( .A(keyinput36), .B(P2_REG2_REG_7__SCAN_IN), .ZN(n15418) );
  NAND4_X1 U16978 ( .A1(n15421), .A2(n15420), .A3(n15419), .A4(n15418), .ZN(
        n15422) );
  NOR3_X1 U16979 ( .A1(n15424), .A2(n15423), .A3(n15422), .ZN(n15440) );
  AOI22_X1 U16980 ( .A1(n12638), .A2(keyinput40), .B1(keyinput30), .B2(n15426), 
        .ZN(n15425) );
  OAI221_X1 U16981 ( .B1(n12638), .B2(keyinput40), .C1(n15426), .C2(keyinput30), .A(n15425), .ZN(n15438) );
  AOI22_X1 U16982 ( .A1(n15429), .A2(keyinput94), .B1(n15428), .B2(keyinput108), .ZN(n15427) );
  OAI221_X1 U16983 ( .B1(n15429), .B2(keyinput94), .C1(n15428), .C2(
        keyinput108), .A(n15427), .ZN(n15437) );
  AOI22_X1 U16984 ( .A1(n15432), .A2(keyinput120), .B1(n15431), .B2(keyinput6), 
        .ZN(n15430) );
  OAI221_X1 U16985 ( .B1(n15432), .B2(keyinput120), .C1(n15431), .C2(keyinput6), .A(n15430), .ZN(n15436) );
  XNOR2_X1 U16986 ( .A(P2_IR_REG_4__SCAN_IN), .B(keyinput96), .ZN(n15434) );
  XNOR2_X1 U16987 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput105), .ZN(n15433) );
  NAND2_X1 U16988 ( .A1(n15434), .A2(n15433), .ZN(n15435) );
  NOR4_X1 U16989 ( .A1(n15438), .A2(n15437), .A3(n15436), .A4(n15435), .ZN(
        n15439) );
  NAND4_X1 U16990 ( .A1(n15442), .A2(n15441), .A3(n15440), .A4(n15439), .ZN(
        n15588) );
  AOI22_X1 U16991 ( .A1(n15445), .A2(keyinput127), .B1(n15444), .B2(keyinput79), .ZN(n15443) );
  OAI221_X1 U16992 ( .B1(n15445), .B2(keyinput127), .C1(n15444), .C2(
        keyinput79), .A(n15443), .ZN(n15456) );
  AOI22_X1 U16993 ( .A1(n15447), .A2(keyinput13), .B1(n13664), .B2(keyinput78), 
        .ZN(n15446) );
  OAI221_X1 U16994 ( .B1(n15447), .B2(keyinput13), .C1(n13664), .C2(keyinput78), .A(n15446), .ZN(n15455) );
  AOI22_X1 U16995 ( .A1(n15450), .A2(keyinput103), .B1(n15449), .B2(keyinput17), .ZN(n15448) );
  OAI221_X1 U16996 ( .B1(n15450), .B2(keyinput103), .C1(n15449), .C2(
        keyinput17), .A(n15448), .ZN(n15454) );
  XNOR2_X1 U16997 ( .A(P3_REG1_REG_31__SCAN_IN), .B(keyinput24), .ZN(n15452)
         );
  XNOR2_X1 U16998 ( .A(P3_IR_REG_14__SCAN_IN), .B(keyinput55), .ZN(n15451) );
  NAND2_X1 U16999 ( .A1(n15452), .A2(n15451), .ZN(n15453) );
  NOR4_X1 U17000 ( .A1(n15456), .A2(n15455), .A3(n15454), .A4(n15453), .ZN(
        n15502) );
  AOI22_X1 U17001 ( .A1(n15459), .A2(keyinput31), .B1(keyinput28), .B2(n15458), 
        .ZN(n15457) );
  OAI221_X1 U17002 ( .B1(n15459), .B2(keyinput31), .C1(n15458), .C2(keyinput28), .A(n15457), .ZN(n15470) );
  AOI22_X1 U17003 ( .A1(n15462), .A2(keyinput53), .B1(n15461), .B2(keyinput111), .ZN(n15460) );
  OAI221_X1 U17004 ( .B1(n15462), .B2(keyinput53), .C1(n15461), .C2(
        keyinput111), .A(n15460), .ZN(n15469) );
  XNOR2_X1 U17005 ( .A(P3_IR_REG_15__SCAN_IN), .B(keyinput81), .ZN(n15465) );
  XNOR2_X1 U17006 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput14), .ZN(n15464) );
  XNOR2_X1 U17007 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput43), .ZN(n15463) );
  NAND3_X1 U17008 ( .A1(n15465), .A2(n15464), .A3(n15463), .ZN(n15468) );
  XNOR2_X1 U17009 ( .A(n15466), .B(keyinput7), .ZN(n15467) );
  NOR4_X1 U17010 ( .A1(n15470), .A2(n15469), .A3(n15468), .A4(n15467), .ZN(
        n15501) );
  AOI22_X1 U17011 ( .A1(n15473), .A2(keyinput25), .B1(keyinput82), .B2(n15472), 
        .ZN(n15471) );
  OAI221_X1 U17012 ( .B1(n15473), .B2(keyinput25), .C1(n15472), .C2(keyinput82), .A(n15471), .ZN(n15483) );
  AOI22_X1 U17013 ( .A1(n15476), .A2(keyinput67), .B1(n15475), .B2(keyinput80), 
        .ZN(n15474) );
  OAI221_X1 U17014 ( .B1(n15476), .B2(keyinput67), .C1(n15475), .C2(keyinput80), .A(n15474), .ZN(n15482) );
  XNOR2_X1 U17015 ( .A(P2_IR_REG_10__SCAN_IN), .B(keyinput118), .ZN(n15480) );
  XNOR2_X1 U17016 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput29), .ZN(n15479) );
  XNOR2_X1 U17017 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput22), .ZN(n15478)
         );
  XNOR2_X1 U17018 ( .A(keyinput112), .B(P2_REG0_REG_6__SCAN_IN), .ZN(n15477)
         );
  NAND4_X1 U17019 ( .A1(n15480), .A2(n15479), .A3(n15478), .A4(n15477), .ZN(
        n15481) );
  NOR3_X1 U17020 ( .A1(n15483), .A2(n15482), .A3(n15481), .ZN(n15500) );
  AOI22_X1 U17021 ( .A1(n15485), .A2(keyinput5), .B1(n7794), .B2(keyinput44), 
        .ZN(n15484) );
  OAI221_X1 U17022 ( .B1(n15485), .B2(keyinput5), .C1(n7794), .C2(keyinput44), 
        .A(n15484), .ZN(n15498) );
  AOI22_X1 U17023 ( .A1(n15488), .A2(keyinput89), .B1(n15487), .B2(keyinput92), 
        .ZN(n15486) );
  OAI221_X1 U17024 ( .B1(n15488), .B2(keyinput89), .C1(n15487), .C2(keyinput92), .A(n15486), .ZN(n15497) );
  AOI22_X1 U17025 ( .A1(n15491), .A2(keyinput38), .B1(n15490), .B2(keyinput60), 
        .ZN(n15489) );
  OAI221_X1 U17026 ( .B1(n15491), .B2(keyinput38), .C1(n15490), .C2(keyinput60), .A(n15489), .ZN(n15496) );
  AOI22_X1 U17027 ( .A1(n15494), .A2(keyinput97), .B1(keyinput54), .B2(n15493), 
        .ZN(n15492) );
  OAI221_X1 U17028 ( .B1(n15494), .B2(keyinput97), .C1(n15493), .C2(keyinput54), .A(n15492), .ZN(n15495) );
  NOR4_X1 U17029 ( .A1(n15498), .A2(n15497), .A3(n15496), .A4(n15495), .ZN(
        n15499) );
  NAND4_X1 U17030 ( .A1(n15502), .A2(n15501), .A3(n15500), .A4(n15499), .ZN(
        n15587) );
  AOI22_X1 U17031 ( .A1(P2_REG1_REG_4__SCAN_IN), .A2(keyinput33), .B1(
        P3_IR_REG_12__SCAN_IN), .B2(keyinput107), .ZN(n15503) );
  OAI221_X1 U17032 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(keyinput33), .C1(
        P3_IR_REG_12__SCAN_IN), .C2(keyinput107), .A(n15503), .ZN(n15510) );
  AOI22_X1 U17033 ( .A1(P1_REG1_REG_24__SCAN_IN), .A2(keyinput65), .B1(
        P1_REG0_REG_29__SCAN_IN), .B2(keyinput83), .ZN(n15504) );
  OAI221_X1 U17034 ( .B1(P1_REG1_REG_24__SCAN_IN), .B2(keyinput65), .C1(
        P1_REG0_REG_29__SCAN_IN), .C2(keyinput83), .A(n15504), .ZN(n15509) );
  AOI22_X1 U17035 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(keyinput91), .B1(
        P3_REG3_REG_5__SCAN_IN), .B2(keyinput35), .ZN(n15505) );
  OAI221_X1 U17036 ( .B1(P1_DATAO_REG_19__SCAN_IN), .B2(keyinput91), .C1(
        P3_REG3_REG_5__SCAN_IN), .C2(keyinput35), .A(n15505), .ZN(n15508) );
  AOI22_X1 U17037 ( .A1(P3_RD_REG_SCAN_IN), .A2(keyinput114), .B1(
        P2_REG1_REG_24__SCAN_IN), .B2(keyinput32), .ZN(n15506) );
  OAI221_X1 U17038 ( .B1(P3_RD_REG_SCAN_IN), .B2(keyinput114), .C1(
        P2_REG1_REG_24__SCAN_IN), .C2(keyinput32), .A(n15506), .ZN(n15507) );
  NOR4_X1 U17039 ( .A1(n15510), .A2(n15509), .A3(n15508), .A4(n15507), .ZN(
        n15585) );
  AOI22_X1 U17040 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(keyinput70), .B1(
        P1_IR_REG_25__SCAN_IN), .B2(keyinput122), .ZN(n15511) );
  OAI221_X1 U17041 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(keyinput70), .C1(
        P1_IR_REG_25__SCAN_IN), .C2(keyinput122), .A(n15511), .ZN(n15518) );
  AOI22_X1 U17042 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput11), .B1(
        P2_REG1_REG_18__SCAN_IN), .B2(keyinput124), .ZN(n15512) );
  OAI221_X1 U17043 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput11), .C1(
        P2_REG1_REG_18__SCAN_IN), .C2(keyinput124), .A(n15512), .ZN(n15517) );
  AOI22_X1 U17044 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(keyinput106), .B1(
        P3_REG0_REG_21__SCAN_IN), .B2(keyinput34), .ZN(n15513) );
  OAI221_X1 U17045 ( .B1(P1_IR_REG_12__SCAN_IN), .B2(keyinput106), .C1(
        P3_REG0_REG_21__SCAN_IN), .C2(keyinput34), .A(n15513), .ZN(n15516) );
  AOI22_X1 U17046 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(keyinput16), .B1(
        P1_REG2_REG_6__SCAN_IN), .B2(keyinput76), .ZN(n15514) );
  OAI221_X1 U17047 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(keyinput16), .C1(
        P1_REG2_REG_6__SCAN_IN), .C2(keyinput76), .A(n15514), .ZN(n15515) );
  NOR4_X1 U17048 ( .A1(n15518), .A2(n15517), .A3(n15516), .A4(n15515), .ZN(
        n15584) );
  OAI22_X1 U17049 ( .A1(P3_REG1_REG_24__SCAN_IN), .A2(keyinput8), .B1(
        P3_REG0_REG_12__SCAN_IN), .B2(keyinput95), .ZN(n15519) );
  AOI221_X1 U17050 ( .B1(P3_REG1_REG_24__SCAN_IN), .B2(keyinput8), .C1(
        keyinput95), .C2(P3_REG0_REG_12__SCAN_IN), .A(n15519), .ZN(n15526) );
  OAI22_X1 U17051 ( .A1(P3_REG3_REG_1__SCAN_IN), .A2(keyinput113), .B1(
        P1_ADDR_REG_3__SCAN_IN), .B2(keyinput123), .ZN(n15520) );
  AOI221_X1 U17052 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(keyinput113), .C1(
        keyinput123), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n15520), .ZN(n15525) );
  OAI22_X1 U17053 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(keyinput26), .B1(
        P2_D_REG_17__SCAN_IN), .B2(keyinput77), .ZN(n15521) );
  AOI221_X1 U17054 ( .B1(P1_DATAO_REG_8__SCAN_IN), .B2(keyinput26), .C1(
        keyinput77), .C2(P2_D_REG_17__SCAN_IN), .A(n15521), .ZN(n15524) );
  OAI22_X1 U17055 ( .A1(P3_D_REG_15__SCAN_IN), .A2(keyinput4), .B1(
        P2_REG0_REG_28__SCAN_IN), .B2(keyinput69), .ZN(n15522) );
  AOI221_X1 U17056 ( .B1(P3_D_REG_15__SCAN_IN), .B2(keyinput4), .C1(keyinput69), .C2(P2_REG0_REG_28__SCAN_IN), .A(n15522), .ZN(n15523) );
  NAND4_X1 U17057 ( .A1(n15526), .A2(n15525), .A3(n15524), .A4(n15523), .ZN(
        n15582) );
  OAI22_X1 U17058 ( .A1(P3_IR_REG_23__SCAN_IN), .A2(keyinput74), .B1(
        P1_REG1_REG_17__SCAN_IN), .B2(keyinput52), .ZN(n15527) );
  AOI221_X1 U17059 ( .B1(P3_IR_REG_23__SCAN_IN), .B2(keyinput74), .C1(
        keyinput52), .C2(P1_REG1_REG_17__SCAN_IN), .A(n15527), .ZN(n15534) );
  OAI22_X1 U17060 ( .A1(P1_REG0_REG_1__SCAN_IN), .A2(keyinput62), .B1(
        P3_ADDR_REG_8__SCAN_IN), .B2(keyinput68), .ZN(n15528) );
  AOI221_X1 U17061 ( .B1(P1_REG0_REG_1__SCAN_IN), .B2(keyinput62), .C1(
        keyinput68), .C2(P3_ADDR_REG_8__SCAN_IN), .A(n15528), .ZN(n15533) );
  OAI22_X1 U17062 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(keyinput85), .B1(
        keyinput1), .B2(P1_REG0_REG_21__SCAN_IN), .ZN(n15529) );
  AOI221_X1 U17063 ( .B1(P1_DATAO_REG_16__SCAN_IN), .B2(keyinput85), .C1(
        P1_REG0_REG_21__SCAN_IN), .C2(keyinput1), .A(n15529), .ZN(n15532) );
  OAI22_X1 U17064 ( .A1(P2_REG1_REG_19__SCAN_IN), .A2(keyinput86), .B1(
        keyinput20), .B2(P3_ADDR_REG_9__SCAN_IN), .ZN(n15530) );
  AOI221_X1 U17065 ( .B1(P2_REG1_REG_19__SCAN_IN), .B2(keyinput86), .C1(
        P3_ADDR_REG_9__SCAN_IN), .C2(keyinput20), .A(n15530), .ZN(n15531) );
  NAND4_X1 U17066 ( .A1(n15534), .A2(n15533), .A3(n15532), .A4(n15531), .ZN(
        n15581) );
  AOI22_X1 U17067 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(keyinput121), .B1(
        P3_IR_REG_8__SCAN_IN), .B2(keyinput58), .ZN(n15535) );
  OAI221_X1 U17068 ( .B1(P3_IR_REG_2__SCAN_IN), .B2(keyinput121), .C1(
        P3_IR_REG_8__SCAN_IN), .C2(keyinput58), .A(n15535), .ZN(n15542) );
  AOI22_X1 U17069 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(keyinput61), .B1(
        P3_REG3_REG_21__SCAN_IN), .B2(keyinput39), .ZN(n15536) );
  OAI221_X1 U17070 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(keyinput61), .C1(
        P3_REG3_REG_21__SCAN_IN), .C2(keyinput39), .A(n15536), .ZN(n15541) );
  AOI22_X1 U17071 ( .A1(P3_REG2_REG_23__SCAN_IN), .A2(keyinput63), .B1(
        P3_REG1_REG_10__SCAN_IN), .B2(keyinput42), .ZN(n15537) );
  OAI221_X1 U17072 ( .B1(P3_REG2_REG_23__SCAN_IN), .B2(keyinput63), .C1(
        P3_REG1_REG_10__SCAN_IN), .C2(keyinput42), .A(n15537), .ZN(n15540) );
  AOI22_X1 U17073 ( .A1(P2_REG2_REG_26__SCAN_IN), .A2(keyinput115), .B1(
        P2_D_REG_31__SCAN_IN), .B2(keyinput48), .ZN(n15538) );
  OAI221_X1 U17074 ( .B1(P2_REG2_REG_26__SCAN_IN), .B2(keyinput115), .C1(
        P2_D_REG_31__SCAN_IN), .C2(keyinput48), .A(n15538), .ZN(n15539) );
  NOR4_X1 U17075 ( .A1(n15542), .A2(n15541), .A3(n15540), .A4(n15539), .ZN(
        n15579) );
  AOI22_X1 U17076 ( .A1(P1_D_REG_4__SCAN_IN), .A2(keyinput88), .B1(
        P3_D_REG_28__SCAN_IN), .B2(keyinput12), .ZN(n15543) );
  OAI221_X1 U17077 ( .B1(P1_D_REG_4__SCAN_IN), .B2(keyinput88), .C1(
        P3_D_REG_28__SCAN_IN), .C2(keyinput12), .A(n15543), .ZN(n15550) );
  AOI22_X1 U17078 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(keyinput125), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(keyinput84), .ZN(n15544) );
  OAI221_X1 U17079 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(keyinput125), .C1(
        P2_DATAO_REG_24__SCAN_IN), .C2(keyinput84), .A(n15544), .ZN(n15549) );
  AOI22_X1 U17080 ( .A1(SI_26_), .A2(keyinput72), .B1(P3_IR_REG_22__SCAN_IN), 
        .B2(keyinput57), .ZN(n15545) );
  OAI221_X1 U17081 ( .B1(SI_26_), .B2(keyinput72), .C1(P3_IR_REG_22__SCAN_IN), 
        .C2(keyinput57), .A(n15545), .ZN(n15548) );
  AOI22_X1 U17082 ( .A1(P3_REG2_REG_11__SCAN_IN), .A2(keyinput110), .B1(SI_18_), .B2(keyinput19), .ZN(n15546) );
  OAI221_X1 U17083 ( .B1(P3_REG2_REG_11__SCAN_IN), .B2(keyinput110), .C1(
        SI_18_), .C2(keyinput19), .A(n15546), .ZN(n15547) );
  NOR4_X1 U17084 ( .A1(n15550), .A2(n15549), .A3(n15548), .A4(n15547), .ZN(
        n15578) );
  AOI22_X1 U17085 ( .A1(n15552), .A2(keyinput49), .B1(keyinput126), .B2(n10134), .ZN(n15551) );
  OAI221_X1 U17086 ( .B1(n15552), .B2(keyinput49), .C1(n10134), .C2(
        keyinput126), .A(n15551), .ZN(n15564) );
  AOI22_X1 U17087 ( .A1(n15555), .A2(keyinput119), .B1(keyinput3), .B2(n15554), 
        .ZN(n15553) );
  OAI221_X1 U17088 ( .B1(n15555), .B2(keyinput119), .C1(n15554), .C2(keyinput3), .A(n15553), .ZN(n15563) );
  AOI22_X1 U17089 ( .A1(n15558), .A2(keyinput73), .B1(n15557), .B2(keyinput51), 
        .ZN(n15556) );
  OAI221_X1 U17090 ( .B1(n15558), .B2(keyinput73), .C1(n15557), .C2(keyinput51), .A(n15556), .ZN(n15562) );
  XNOR2_X1 U17091 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(keyinput64), .ZN(n15560)
         );
  XNOR2_X1 U17092 ( .A(P2_IR_REG_23__SCAN_IN), .B(keyinput45), .ZN(n15559) );
  NAND2_X1 U17093 ( .A1(n15560), .A2(n15559), .ZN(n15561) );
  NOR4_X1 U17094 ( .A1(n15564), .A2(n15563), .A3(n15562), .A4(n15561), .ZN(
        n15577) );
  AOI22_X1 U17095 ( .A1(n15567), .A2(keyinput47), .B1(n15566), .B2(keyinput2), 
        .ZN(n15565) );
  OAI221_X1 U17096 ( .B1(n15567), .B2(keyinput47), .C1(n15566), .C2(keyinput2), 
        .A(n15565), .ZN(n15575) );
  AOI22_X1 U17097 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(keyinput37), .B1(
        P3_D_REG_2__SCAN_IN), .B2(keyinput117), .ZN(n15568) );
  OAI221_X1 U17098 ( .B1(P2_DATAO_REG_20__SCAN_IN), .B2(keyinput37), .C1(
        P3_D_REG_2__SCAN_IN), .C2(keyinput117), .A(n15568), .ZN(n15574) );
  AOI22_X1 U17099 ( .A1(P1_REG1_REG_25__SCAN_IN), .A2(keyinput87), .B1(
        P3_REG3_REG_24__SCAN_IN), .B2(keyinput71), .ZN(n15569) );
  OAI221_X1 U17100 ( .B1(P1_REG1_REG_25__SCAN_IN), .B2(keyinput87), .C1(
        P3_REG3_REG_24__SCAN_IN), .C2(keyinput71), .A(n15569), .ZN(n15573) );
  XOR2_X1 U17101 ( .A(n13108), .B(keyinput27), .Z(n15571) );
  XNOR2_X1 U17102 ( .A(P2_IR_REG_21__SCAN_IN), .B(keyinput15), .ZN(n15570) );
  NAND2_X1 U17103 ( .A1(n15571), .A2(n15570), .ZN(n15572) );
  NOR4_X1 U17104 ( .A1(n15575), .A2(n15574), .A3(n15573), .A4(n15572), .ZN(
        n15576) );
  NAND4_X1 U17105 ( .A1(n15579), .A2(n15578), .A3(n15577), .A4(n15576), .ZN(
        n15580) );
  NOR3_X1 U17106 ( .A1(n15582), .A2(n15581), .A3(n15580), .ZN(n15583) );
  NAND3_X1 U17107 ( .A1(n15585), .A2(n15584), .A3(n15583), .ZN(n15586) );
  NOR4_X1 U17108 ( .A1(n15589), .A2(n15588), .A3(n15587), .A4(n15586), .ZN(
        n15602) );
  AOI22_X1 U17109 ( .A1(n15595), .A2(P3_REG2_REG_11__SCAN_IN), .B1(n15591), 
        .B2(n15590), .ZN(n15592) );
  OAI21_X1 U17110 ( .B1(n15594), .B2(n15593), .A(n15592), .ZN(n15598) );
  NOR2_X1 U17111 ( .A1(n15596), .A2(n15595), .ZN(n15597) );
  AOI211_X1 U17112 ( .C1(n15600), .C2(n15599), .A(n15598), .B(n15597), .ZN(
        n15601) );
  XNOR2_X1 U17113 ( .A(n15602), .B(n15601), .ZN(P3_U3222) );
  AOI21_X1 U17114 ( .B1(n15604), .B2(n15603), .A(n15616), .ZN(SUB_1596_U53) );
  XNOR2_X1 U17115 ( .A(n15605), .B(n15606), .ZN(SUB_1596_U59) );
  XNOR2_X1 U17116 ( .A(n15607), .B(P2_ADDR_REG_5__SCAN_IN), .ZN(SUB_1596_U58)
         );
  XNOR2_X1 U17117 ( .A(n15608), .B(n15609), .ZN(SUB_1596_U56) );
  OAI21_X1 U17118 ( .B1(n15612), .B2(n15611), .A(n15610), .ZN(n15614) );
  XOR2_X1 U17119 ( .A(n15614), .B(n15613), .Z(SUB_1596_U60) );
  XOR2_X1 U17120 ( .A(n15616), .B(n15615), .Z(SUB_1596_U5) );
  CLKBUF_X2 U7392 ( .A(n12027), .Z(n12051) );
  CLKBUF_X1 U7400 ( .A(n8565), .Z(n8670) );
  NAND3_X1 U7423 ( .A1(n8750), .A2(n8749), .A3(n11735), .ZN(n11442) );
endmodule

