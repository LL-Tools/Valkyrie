

module b21_C_AntiSAT_k_256_7 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, 
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, 
        keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, 
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, 
        keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, 
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, 
        keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, 
        keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, 
        keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, 
        keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, 
        keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, 
        keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, 
        keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, 
        keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, 
        keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, 
        keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, 
        keyinput180, keyinput181, keyinput182, keyinput183, keyinput184, 
        keyinput185, keyinput186, keyinput187, keyinput188, keyinput189, 
        keyinput190, keyinput191, keyinput192, keyinput193, keyinput194, 
        keyinput195, keyinput196, keyinput197, keyinput198, keyinput199, 
        keyinput200, keyinput201, keyinput202, keyinput203, keyinput204, 
        keyinput205, keyinput206, keyinput207, keyinput208, keyinput209, 
        keyinput210, keyinput211, keyinput212, keyinput213, keyinput214, 
        keyinput215, keyinput216, keyinput217, keyinput218, keyinput219, 
        keyinput220, keyinput221, keyinput222, keyinput223, keyinput224, 
        keyinput225, keyinput226, keyinput227, keyinput228, keyinput229, 
        keyinput230, keyinput231, keyinput232, keyinput233, keyinput234, 
        keyinput235, keyinput236, keyinput237, keyinput238, keyinput239, 
        keyinput240, keyinput241, keyinput242, keyinput243, keyinput244, 
        keyinput245, keyinput246, keyinput247, keyinput248, keyinput249, 
        keyinput250, keyinput251, keyinput252, keyinput253, keyinput254, 
        keyinput255, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, 
        ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, 
        ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, 
        ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, 
        ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, 
        P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, 
        P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, 
        P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, 
        P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, 
        P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, 
        P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, 
        P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, 
        P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, 
        P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, 
        P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, 
        P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, 
        P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, 
        P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, 
        P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, 
        P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, 
        P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, 
        P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, 
        P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, 
        P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, 
        P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, 
        P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, 
        P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, 
        P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, 
        P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, 
        P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, 
        P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, 
        P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, 
        P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, 
        P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, 
        P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, 
        P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, 
        P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, 
        P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, 
        P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, 
        P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, 
        P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, 
        P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10593;

  INV_X1 U5002 ( .A(n7014), .ZN(n6820) );
  OR2_X1 U5003 ( .A1(n7100), .A2(n6715), .ZN(n7172) );
  CLKBUF_X2 U5004 ( .A(n6163), .Z(n6131) );
  AND2_X1 U5005 ( .A1(n8883), .A2(n8474), .ZN(n6163) );
  XNOR2_X1 U5006 ( .A(n5852), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5865) );
  AND2_X1 U5007 ( .A1(n5830), .A2(n4908), .ZN(n4774) );
  AND2_X1 U5008 ( .A1(n5102), .A2(n5057), .ZN(n5103) );
  INV_X2 U5009 ( .A(n7173), .ZN(n6676) );
  INV_X1 U5010 ( .A(n8879), .ZN(n7272) );
  AND2_X1 U5011 ( .A1(n5833), .A2(n4743), .ZN(n4742) );
  INV_X1 U5012 ( .A(n8938), .ZN(n7521) );
  NAND2_X1 U5013 ( .A1(n9541), .A2(n9522), .ZN(n8938) );
  INV_X1 U5014 ( .A(n7013), .ZN(n5311) );
  INV_X1 U5015 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9696) );
  INV_X1 U5016 ( .A(n6160), .ZN(n6173) );
  INV_X2 U5017 ( .A(n4502), .ZN(n6244) );
  INV_X1 U5018 ( .A(n6410), .ZN(n4733) );
  AND2_X1 U5019 ( .A1(n8883), .A2(n5865), .ZN(n6164) );
  NAND2_X1 U5020 ( .A1(n6458), .A2(n6457), .ZN(n6160) );
  AND2_X1 U5021 ( .A1(n8867), .A2(n9928), .ZN(n9912) );
  INV_X1 U5022 ( .A(n6180), .ZN(n10373) );
  NAND2_X1 U5023 ( .A1(n5310), .A2(n5309), .ZN(n10505) );
  AOI21_X1 U5024 ( .B1(n8515), .B2(n8514), .A(n9912), .ZN(n8869) );
  NAND2_X1 U5025 ( .A1(n7920), .A2(n7919), .ZN(n8149) );
  XNOR2_X1 U5026 ( .A(n5851), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5854) );
  CLKBUF_X3 U5027 ( .A(n5175), .Z(n6889) );
  INV_X1 U5028 ( .A(n5109), .ZN(n8476) );
  INV_X1 U5029 ( .A(n5155), .ZN(n8931) );
  AND3_X1 U5030 ( .A1(n4547), .A2(n4582), .A3(n8872), .ZN(n4497) );
  NAND2_X2 U5031 ( .A1(n7836), .A2(n7837), .ZN(n8078) );
  NOR2_X4 U5032 ( .A1(n8233), .A2(n8332), .ZN(n8317) );
  OR2_X2 U5033 ( .A1(n5150), .A2(n9696), .ZN(n5147) );
  AOI21_X2 U5034 ( .B1(n5213), .B2(n5212), .A(n5070), .ZN(n5235) );
  OAI21_X2 U5035 ( .B1(n9262), .B2(n9626), .A(n6778), .ZN(n9494) );
  XNOR2_X2 U5036 ( .A(n6467), .B(n6466), .ZN(n7951) );
  AOI22_X2 U5037 ( .A1(n10026), .A2(n8483), .B1(n8482), .B2(n10032), .ZN(
        n10013) );
  BUF_X4 U5038 ( .A(n5279), .Z(n4498) );
  NAND2_X1 U5039 ( .A1(n8478), .A2(n8476), .ZN(n5279) );
  OAI21_X1 U5040 ( .B1(n9920), .B2(n9919), .A(n9918), .ZN(n10066) );
  INV_X2 U5041 ( .A(n10349), .ZN(n10048) );
  INV_X4 U5042 ( .A(n5576), .ZN(n5661) );
  NAND2_X1 U5043 ( .A1(n8877), .A2(n6180), .ZN(n6417) );
  INV_X1 U5044 ( .A(n7173), .ZN(n6660) );
  INV_X4 U5045 ( .A(n6678), .ZN(n6476) );
  INV_X2 U5046 ( .A(n4498), .ZN(n5189) );
  INV_X1 U5047 ( .A(n9902), .ZN(n7367) );
  OAI21_X1 U5048 ( .B1(n4736), .B2(n4735), .A(n4734), .ZN(n6407) );
  OAI21_X1 U5049 ( .B1(n4698), .B2(n9122), .A(n8942), .ZN(n4697) );
  OR2_X1 U5050 ( .A1(n10063), .A2(n4767), .ZN(n10138) );
  NAND2_X1 U5051 ( .A1(n6399), .A2(n4737), .ZN(n6405) );
  AOI21_X1 U5052 ( .B1(n9117), .B2(n4700), .A(n4699), .ZN(n4698) );
  OR2_X1 U5053 ( .A1(n10066), .A2(n10412), .ZN(n4769) );
  NAND2_X1 U5054 ( .A1(n9375), .A2(n6784), .ZN(n9366) );
  AND2_X1 U5055 ( .A1(n4859), .A2(n4857), .ZN(n9239) );
  AOI21_X1 U5056 ( .B1(n9200), .B2(n9199), .A(n5072), .ZN(n9191) );
  AND2_X1 U5057 ( .A1(n4614), .A2(n4613), .ZN(n5671) );
  NOR2_X1 U5058 ( .A1(n10064), .A2(n4551), .ZN(n4768) );
  OR2_X1 U5059 ( .A1(n8923), .A2(n4505), .ZN(n8925) );
  AND2_X1 U5060 ( .A1(n9407), .A2(n9656), .ZN(n4516) );
  NAND2_X1 U5061 ( .A1(n6243), .A2(n6242), .ZN(n8923) );
  OR3_X1 U5062 ( .A1(n9407), .A2(n9406), .A3(n10520), .ZN(n9588) );
  OAI21_X1 U5063 ( .B1(n6249), .B2(n6241), .A(n6240), .ZN(n6242) );
  OR2_X1 U5064 ( .A1(n6251), .A2(n6249), .ZN(n6243) );
  NAND2_X1 U5065 ( .A1(n5740), .A2(n5739), .ZN(n9372) );
  NAND2_X1 U5066 ( .A1(n10051), .A2(n8496), .ZN(n10034) );
  NAND2_X1 U5067 ( .A1(n6195), .A2(n6194), .ZN(n10079) );
  NAND2_X1 U5068 ( .A1(n10052), .A2(n10053), .ZN(n10051) );
  NAND2_X1 U5069 ( .A1(n6806), .A2(n6805), .ZN(n9557) );
  NAND2_X1 U5070 ( .A1(n5893), .A2(n5892), .ZN(n10092) );
  XNOR2_X1 U5071 ( .A(n5650), .B(n5649), .ZN(n7844) );
  NAND2_X1 U5072 ( .A1(n5903), .A2(n5902), .ZN(n10098) );
  NAND2_X1 U5073 ( .A1(n5615), .A2(n5614), .ZN(n9486) );
  OR2_X1 U5074 ( .A1(n5644), .A2(n5643), .ZN(n5658) );
  OR2_X1 U5075 ( .A1(n5422), .A2(n7994), .ZN(n5424) );
  AND2_X1 U5076 ( .A1(n9043), .A2(n9045), .ZN(n8956) );
  NAND2_X1 U5077 ( .A1(n5976), .A2(n5975), .ZN(n10122) );
  NAND2_X1 U5078 ( .A1(n6001), .A2(n6000), .ZN(n10270) );
  NAND2_X1 U5079 ( .A1(n9041), .A2(n9039), .ZN(n8953) );
  OAI211_X1 U5080 ( .C1(n4619), .C2(n5661), .A(n4616), .B(n4615), .ZN(n8047)
         );
  AND2_X1 U5081 ( .A1(n10327), .A2(n10415), .ZN(n10329) );
  NAND2_X1 U5082 ( .A1(n4619), .A2(n5388), .ZN(n6765) );
  NAND2_X1 U5083 ( .A1(n6027), .A2(n6026), .ZN(n10237) );
  AND2_X1 U5084 ( .A1(n10334), .A2(n7400), .ZN(n7320) );
  AND2_X1 U5085 ( .A1(n7178), .A2(n7337), .ZN(n7242) );
  INV_X2 U5086 ( .A(n9540), .ZN(n4499) );
  AND2_X1 U5087 ( .A1(n7069), .A2(n7073), .ZN(n8875) );
  NOR2_X1 U5089 ( .A1(n7291), .A2(n6179), .ZN(n7178) );
  AND3_X1 U5090 ( .A1(n5294), .A2(n5293), .A3(n5292), .ZN(n7633) );
  INV_X1 U5091 ( .A(n7244), .ZN(n10391) );
  NAND2_X1 U5092 ( .A1(n4923), .A2(n4921), .ZN(n5349) );
  AND2_X1 U5093 ( .A1(n9009), .A2(n9011), .ZN(n7467) );
  NOR2_X1 U5094 ( .A1(n7225), .A2(n7205), .ZN(n7219) );
  AND3_X1 U5095 ( .A1(n5179), .A2(n5178), .A3(n5177), .ZN(n10482) );
  NAND2_X1 U5096 ( .A1(n4648), .A2(n5260), .ZN(n5286) );
  NAND4_X2 U5097 ( .A1(n5168), .A2(n5167), .A3(n5166), .A4(n5165), .ZN(n9279)
         );
  AND4_X1 U5098 ( .A1(n6099), .A2(n6098), .A3(n6097), .A4(n6096), .ZN(n8877)
         );
  NAND2_X1 U5099 ( .A1(n7803), .A2(n9902), .ZN(n6717) );
  NAND2_X1 U5100 ( .A1(n5238), .A2(n5237), .ZN(n5257) );
  CLKBUF_X2 U5101 ( .A(n6174), .Z(n4502) );
  AND2_X2 U5102 ( .A1(n5110), .A2(n8476), .ZN(n7013) );
  INV_X2 U5103 ( .A(n6487), .ZN(n6731) );
  INV_X2 U5104 ( .A(n5437), .ZN(n4504) );
  NAND2_X2 U5105 ( .A1(n5106), .A2(n5109), .ZN(n5792) );
  XNOR2_X1 U5106 ( .A(n4636), .B(P1_IR_REG_22__SCAN_IN), .ZN(n6470) );
  XNOR2_X1 U5107 ( .A(n5108), .B(n5107), .ZN(n8478) );
  NOR2_X1 U5108 ( .A1(n8883), .A2(n5865), .ZN(n6162) );
  NAND2_X1 U5109 ( .A1(n5152), .A2(n5151), .ZN(n9129) );
  NAND2_X1 U5110 ( .A1(n6294), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4636) );
  OAI21_X1 U5111 ( .B1(n5172), .B2(n4917), .A(n5174), .ZN(n5197) );
  NAND2_X1 U5112 ( .A1(n5850), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5852) );
  NAND2_X1 U5113 ( .A1(n10153), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5851) );
  XNOR2_X1 U5114 ( .A(n5923), .B(P1_IR_REG_19__SCAN_IN), .ZN(n9902) );
  AND2_X1 U5115 ( .A1(n5290), .A2(n5047), .ZN(n5758) );
  INV_X1 U5116 ( .A(n5844), .ZN(n5843) );
  NAND2_X1 U5117 ( .A1(n4775), .A2(n5921), .ZN(n5844) );
  AND2_X1 U5118 ( .A1(n4532), .A2(n4785), .ZN(n5047) );
  AND2_X1 U5119 ( .A1(n5829), .A2(n5828), .ZN(n4773) );
  AND4_X1 U5120 ( .A1(n5933), .A2(n5997), .A3(n5983), .A4(n6023), .ZN(n5830)
         );
  AND4_X1 U5121 ( .A1(n6115), .A2(n5824), .A3(n5823), .A4(n5822), .ZN(n5829)
         );
  AND2_X1 U5122 ( .A1(n5100), .A2(n5101), .ZN(n4784) );
  INV_X1 U5123 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n6115) );
  INV_X1 U5124 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5997) );
  NOR2_X1 U5125 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5831) );
  NOR2_X1 U5126 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n5840) );
  OR2_X1 U5127 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n5842) );
  NOR3_X1 U5128 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .A3(
        P1_IR_REG_21__SCAN_IN), .ZN(n5835) );
  NOR2_X2 U5129 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5176) );
  NOR2_X1 U5130 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5031) );
  INV_X4 U5131 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U5132 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5141) );
  INV_X1 U5133 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5462) );
  NOR2_X1 U5134 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n6101) );
  INV_X4 U5135 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  XNOR2_X2 U5136 ( .A(n9327), .B(n9332), .ZN(n9314) );
  AND2_X2 U5137 ( .A1(n9312), .A2(n4877), .ZN(n9327) );
  NAND4_X2 U5138 ( .A1(n6147), .A2(n6146), .A3(n6145), .A4(n6144), .ZN(n6410)
         );
  NOR3_X2 U5139 ( .A1(n9501), .A2(n9439), .A3(n4788), .ZN(n4786) );
  INV_X1 U5140 ( .A(n6458), .ZN(n4500) );
  INV_X1 U5141 ( .A(n4500), .ZN(n4501) );
  OAI22_X2 U5142 ( .A1(n8310), .A2(n4650), .B1(n4533), .B2(n4649), .ZN(n8481)
         );
  OAI22_X4 U5143 ( .A1(n8151), .A2(n4981), .B1(n8229), .B2(n4985), .ZN(n8310)
         );
  XNOR2_X2 U5144 ( .A(n5147), .B(n5146), .ZN(n5799) );
  AND2_X1 U5145 ( .A1(n7723), .A2(n6889), .ZN(n4503) );
  XNOR2_X2 U5146 ( .A(n5838), .B(P1_IR_REG_27__SCAN_IN), .ZN(n6457) );
  NOR3_X4 U5147 ( .A1(n10014), .A2(n4914), .A3(n10072), .ZN(n4564) );
  OR2_X4 U5148 ( .A1(n10027), .A2(n10092), .ZN(n10014) );
  INV_X1 U5149 ( .A(n5436), .ZN(n4505) );
  INV_X1 U5150 ( .A(n5437), .ZN(n5436) );
  NAND2_X1 U5151 ( .A1(n7723), .A2(n5199), .ZN(n5437) );
  OR2_X1 U5152 ( .A1(n5476), .A2(n4850), .ZN(n4849) );
  OR2_X1 U5153 ( .A1(n9402), .A2(n9391), .ZN(n9381) );
  AND2_X1 U5154 ( .A1(n4820), .A2(n5528), .ZN(n4819) );
  NAND2_X1 U5155 ( .A1(n5516), .A2(n5492), .ZN(n4820) );
  AOI21_X1 U5156 ( .B1(n4660), .B2(n4663), .A(n4535), .ZN(n4658) );
  AND2_X1 U5157 ( .A1(n9026), .A2(n9028), .ZN(n4683) );
  INV_X1 U5158 ( .A(n9701), .ZN(n5011) );
  INV_X1 U5159 ( .A(n8047), .ZN(n5394) );
  OR2_X1 U5160 ( .A1(n8361), .A2(n8303), .ZN(n9061) );
  OR2_X1 U5161 ( .A1(n8917), .A2(n8249), .ZN(n9056) );
  OR2_X1 U5162 ( .A1(n9279), .A2(n7457), .ZN(n9008) );
  OR2_X1 U5163 ( .A1(n6668), .A2(n6667), .ZN(n6670) );
  NAND2_X1 U5164 ( .A1(n6664), .A2(n5011), .ZN(n5009) );
  AND2_X1 U5165 ( .A1(n6670), .A2(n5009), .ZN(n5008) );
  NAND2_X1 U5166 ( .A1(n10243), .A2(n4759), .ZN(n7764) );
  AND2_X1 U5167 ( .A1(n7761), .A2(n7760), .ZN(n4759) );
  INV_X1 U5168 ( .A(n7320), .ZN(n7315) );
  NAND2_X1 U5169 ( .A1(n10270), .A2(n7928), .ZN(n7924) );
  AND2_X1 U5170 ( .A1(n4962), .A2(n4776), .ZN(n4775) );
  NOR2_X1 U5171 ( .A1(n5841), .A2(n5842), .ZN(n4776) );
  NAND2_X1 U5172 ( .A1(n4797), .A2(n5610), .ZN(n5631) );
  NAND2_X1 U5173 ( .A1(n5612), .A2(n5611), .ZN(n4797) );
  AND2_X1 U5174 ( .A1(n5609), .A2(n5608), .ZN(n5611) );
  AND2_X1 U5175 ( .A1(n5529), .A2(n5496), .ZN(n5528) );
  NAND2_X1 U5176 ( .A1(n5489), .A2(n5488), .ZN(n5492) );
  NAND2_X1 U5177 ( .A1(n5487), .A2(n5486), .ZN(n5517) );
  NAND2_X1 U5178 ( .A1(n4809), .A2(n4807), .ZN(n5487) );
  OAI21_X1 U5179 ( .B1(P1_ADDR_REG_19__SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        n5141), .ZN(n4645) );
  NAND2_X1 U5180 ( .A1(n4647), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4646) );
  NAND2_X1 U5181 ( .A1(n5421), .A2(n4622), .ZN(n7996) );
  INV_X1 U5182 ( .A(n5420), .ZN(n4622) );
  OR2_X1 U5183 ( .A1(n5665), .A2(n5664), .ZN(n5685) );
  AND2_X1 U5184 ( .A1(n4848), .A2(n5527), .ZN(n4847) );
  NAND2_X1 U5185 ( .A1(n4517), .A2(n4850), .ZN(n4848) );
  NOR2_X1 U5186 ( .A1(n8093), .A2(n4872), .ZN(n8182) );
  AND2_X1 U5187 ( .A1(n7708), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4872) );
  NOR2_X1 U5188 ( .A1(n7707), .A2(n4598), .ZN(n8186) );
  AND2_X1 U5189 ( .A1(n7708), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4598) );
  NAND2_X1 U5190 ( .A1(n9299), .A2(n4562), .ZN(n9317) );
  NAND2_X1 U5191 ( .A1(n9106), .A2(n6785), .ZN(n9365) );
  AND2_X1 U5192 ( .A1(n4927), .A2(n6783), .ZN(n4926) );
  NAND2_X1 U5193 ( .A1(n9403), .A2(n4928), .ZN(n4927) );
  INV_X1 U5194 ( .A(n6782), .ZN(n4928) );
  INV_X1 U5195 ( .A(n9403), .ZN(n4929) );
  NAND2_X1 U5196 ( .A1(n9381), .A2(n9380), .ZN(n9403) );
  NAND2_X1 U5197 ( .A1(n6815), .A2(n6814), .ZN(n9379) );
  OR2_X1 U5198 ( .A1(n6813), .A2(n6812), .ZN(n6814) );
  OR2_X1 U5199 ( .A1(n9439), .A2(n9257), .ZN(n6781) );
  NAND2_X1 U5200 ( .A1(n8976), .A2(n8975), .ZN(n9425) );
  NAND2_X1 U5201 ( .A1(n6776), .A2(n6775), .ZN(n9512) );
  INV_X2 U5202 ( .A(n7723), .ZN(n7009) );
  OR2_X1 U5203 ( .A1(n5103), .A2(n9696), .ZN(n5105) );
  AND2_X1 U5204 ( .A1(n5290), .A2(n5116), .ZN(n4864) );
  NAND2_X1 U5205 ( .A1(n5029), .A2(n5028), .ZN(n5027) );
  INV_X1 U5206 ( .A(n6689), .ZN(n5029) );
  NAND2_X1 U5207 ( .A1(n5007), .A2(n6670), .ZN(n5006) );
  INV_X1 U5208 ( .A(n9752), .ZN(n5007) );
  NOR2_X1 U5209 ( .A1(n7056), .A2(n4890), .ZN(n6948) );
  AND2_X1 U5210 ( .A1(n7052), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4890) );
  NAND2_X1 U5211 ( .A1(n4574), .A2(n4573), .ZN(n4896) );
  INV_X1 U5212 ( .A(n7195), .ZN(n4573) );
  NOR2_X1 U5213 ( .A1(n8016), .A2(n7923), .ZN(n8279) );
  NAND2_X1 U5214 ( .A1(n4563), .A2(n9926), .ZN(n8489) );
  NOR2_X1 U5215 ( .A1(n4979), .A2(n4975), .ZN(n4974) );
  INV_X1 U5216 ( .A(n4977), .ZN(n4975) );
  NAND2_X1 U5217 ( .A1(n4973), .A2(n4972), .ZN(n4971) );
  NAND2_X1 U5218 ( .A1(n4980), .A2(n8487), .ZN(n4972) );
  INV_X1 U5219 ( .A(n4979), .ZN(n4973) );
  INV_X1 U5220 ( .A(n4655), .ZN(n4649) );
  NAND2_X1 U5221 ( .A1(n4653), .A2(n4655), .ZN(n4650) );
  OR2_X1 U5222 ( .A1(n10122), .A2(n8226), .ZN(n8223) );
  INV_X1 U5223 ( .A(n4982), .ZN(n8229) );
  NAND2_X1 U5224 ( .A1(n10122), .A2(n9818), .ZN(n4985) );
  AOI21_X1 U5225 ( .B1(n4957), .B2(n4959), .A(n4528), .ZN(n4955) );
  NAND2_X1 U5226 ( .A1(n5988), .A2(n5987), .ZN(n10129) );
  NAND2_X1 U5227 ( .A1(n6459), .A2(n5837), .ZN(n5838) );
  NAND2_X1 U5228 ( .A1(n7530), .A2(n5252), .ZN(n7532) );
  NAND2_X1 U5229 ( .A1(n4691), .A2(n4690), .ZN(n4689) );
  AND2_X1 U5230 ( .A1(n9013), .A2(n9014), .ZN(n4690) );
  OAI21_X1 U5231 ( .B1(n9004), .B2(n9005), .A(n9003), .ZN(n4691) );
  AOI21_X1 U5232 ( .B1(n6306), .B2(n6305), .A(n6426), .ZN(n6307) );
  NOR2_X1 U5233 ( .A1(n6373), .A2(n7401), .ZN(n4730) );
  AOI21_X1 U5234 ( .B1(n9027), .B2(n4682), .A(n4681), .ZN(n9042) );
  AND2_X1 U5235 ( .A1(n9038), .A2(n4683), .ZN(n4682) );
  NAND2_X1 U5236 ( .A1(n4728), .A2(n4725), .ZN(n6318) );
  AOI21_X1 U5237 ( .B1(n4707), .B2(n4705), .A(n4704), .ZN(n4703) );
  NAND2_X1 U5238 ( .A1(n9053), .A2(n9054), .ZN(n4704) );
  AOI21_X1 U5239 ( .B1(n9048), .B2(n4706), .A(n9055), .ZN(n4705) );
  NAND2_X1 U5240 ( .A1(n9047), .A2(n9111), .ZN(n4707) );
  NOR2_X1 U5241 ( .A1(n4721), .A2(n4720), .ZN(n4719) );
  AOI21_X1 U5242 ( .B1(n4721), .B2(n8455), .A(n4718), .ZN(n4717) );
  NOR2_X1 U5243 ( .A1(n9816), .A2(n6717), .ZN(n4720) );
  NAND2_X1 U5244 ( .A1(n4679), .A2(n4676), .ZN(n9083) );
  OAI21_X1 U5245 ( .B1(n4680), .B2(n9077), .A(n9111), .ZN(n4679) );
  AOI21_X1 U5246 ( .B1(n9079), .B2(n9082), .A(n5051), .ZN(n4680) );
  NAND2_X1 U5247 ( .A1(n9275), .A2(n7539), .ZN(n8987) );
  OAI21_X1 U5248 ( .B1(n6357), .B2(n6356), .A(n4747), .ZN(n4746) );
  AND2_X1 U5249 ( .A1(n8498), .A2(n6355), .ZN(n4747) );
  NAND2_X1 U5250 ( .A1(n4713), .A2(n4710), .ZN(n4709) );
  AOI21_X1 U5251 ( .B1(n9084), .B2(n4711), .A(n9446), .ZN(n4710) );
  NAND2_X1 U5252 ( .A1(n4714), .A2(n9111), .ZN(n4713) );
  NOR2_X1 U5253 ( .A1(n4712), .A2(n9111), .ZN(n4711) );
  NAND2_X1 U5254 ( .A1(n9097), .A2(n9419), .ZN(n4708) );
  INV_X1 U5255 ( .A(n6643), .ZN(n5004) );
  OR2_X1 U5256 ( .A1(n9913), .A2(n6266), .ZN(n6290) );
  INV_X1 U5257 ( .A(n5692), .ZN(n4827) );
  NAND2_X1 U5258 ( .A1(n5377), .A2(SI_11_), .ZN(n5378) );
  NAND2_X1 U5259 ( .A1(n7996), .A2(n5415), .ZN(n5422) );
  INV_X1 U5260 ( .A(n5388), .ZN(n4618) );
  INV_X1 U5261 ( .A(n4860), .ZN(n4858) );
  NAND2_X1 U5262 ( .A1(n9113), .A2(n6818), .ZN(n5036) );
  NAND2_X1 U5263 ( .A1(n4538), .A2(n9113), .ZN(n5035) );
  AOI21_X1 U5264 ( .B1(n5035), .B2(n5036), .A(n8930), .ZN(n5033) );
  OR2_X1 U5265 ( .A1(n6834), .A2(n7185), .ZN(n9112) );
  OR2_X1 U5266 ( .A1(n9427), .A2(n9244), .ZN(n8976) );
  NAND2_X1 U5267 ( .A1(n4949), .A2(n4951), .ZN(n4946) );
  OR2_X1 U5268 ( .A1(n9468), .A2(n9259), .ZN(n4945) );
  NOR2_X1 U5269 ( .A1(n4950), .A2(n9463), .ZN(n4948) );
  NOR2_X1 U5270 ( .A1(n9054), .A2(n4934), .ZN(n4932) );
  OR2_X1 U5271 ( .A1(n6765), .A2(n8051), .ZN(n9043) );
  OR2_X1 U5272 ( .A1(n7957), .A2(n7992), .ZN(n9041) );
  OR2_X1 U5273 ( .A1(n8040), .A2(n8895), .ZN(n9032) );
  AND2_X1 U5274 ( .A1(n7508), .A2(n6794), .ZN(n6795) );
  OR2_X1 U5275 ( .A1(n9273), .A2(n7633), .ZN(n9018) );
  INV_X1 U5276 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5101) );
  AND2_X1 U5277 ( .A1(n5758), .A2(n5100), .ZN(n5102) );
  INV_X1 U5278 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5438) );
  INV_X1 U5279 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5384) );
  INV_X1 U5280 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5459) );
  AOI21_X1 U5281 ( .B1(n7350), .B2(n4992), .A(n4991), .ZN(n4990) );
  INV_X1 U5282 ( .A(n6545), .ZN(n4991) );
  NAND2_X1 U5283 ( .A1(n7148), .A2(n4632), .ZN(n4631) );
  NOR2_X1 U5284 ( .A1(n6535), .A2(n4633), .ZN(n4632) );
  INV_X1 U5285 ( .A(n6519), .ZN(n4633) );
  AOI21_X1 U5286 ( .B1(n9813), .B2(n9909), .A(n10262), .ZN(n6397) );
  OR2_X1 U5287 ( .A1(n10067), .A2(n9926), .ZN(n9923) );
  OR2_X1 U5288 ( .A1(n10072), .A2(n9974), .ZN(n6268) );
  AND2_X1 U5289 ( .A1(n10084), .A2(n10007), .ZN(n4979) );
  AND2_X1 U5290 ( .A1(n4906), .A2(n9722), .ZN(n4905) );
  NAND2_X1 U5291 ( .A1(n10112), .A2(n9815), .ZN(n4655) );
  NOR2_X1 U5292 ( .A1(n10112), .A2(n10119), .ZN(n4906) );
  OAI211_X1 U5293 ( .C1(n7765), .C2(n4762), .A(n4761), .B(n6332), .ZN(n4760)
         );
  NAND2_X1 U5294 ( .A1(n4765), .A2(n4766), .ZN(n4761) );
  NAND2_X1 U5295 ( .A1(n4763), .A2(n4766), .ZN(n4762) );
  NAND2_X1 U5296 ( .A1(n9829), .A2(n7166), .ZN(n7126) );
  NAND2_X1 U5297 ( .A1(n7319), .A2(n4526), .ZN(n10335) );
  OAI21_X1 U5298 ( .B1(n5658), .B2(n4826), .A(n4822), .ZN(n5709) );
  AOI21_X1 U5299 ( .B1(n4825), .B2(n4824), .A(n4823), .ZN(n4822) );
  INV_X1 U5300 ( .A(n5691), .ZN(n4823) );
  INV_X1 U5301 ( .A(n4831), .ZN(n4824) );
  INV_X1 U5302 ( .A(n5835), .ZN(n4963) );
  NAND2_X1 U5303 ( .A1(n4798), .A2(n5593), .ZN(n5612) );
  INV_X1 U5304 ( .A(n5591), .ZN(n4798) );
  INV_X1 U5305 ( .A(n4817), .ZN(n4816) );
  OAI21_X1 U5306 ( .B1(n4819), .B2(n4818), .A(n5549), .ZN(n4817) );
  NAND2_X1 U5307 ( .A1(n5492), .A2(n5491), .ZN(n5516) );
  NAND2_X1 U5308 ( .A1(n4666), .A2(n4664), .ZN(n4809) );
  AND2_X1 U5309 ( .A1(n4665), .A2(n4810), .ZN(n4664) );
  AND2_X1 U5310 ( .A1(n4811), .A2(n5067), .ZN(n4810) );
  NAND2_X1 U5311 ( .A1(n4583), .A2(n5378), .ZN(n5432) );
  NAND2_X1 U5312 ( .A1(n5375), .A2(n4670), .ZN(n4583) );
  NAND2_X1 U5313 ( .A1(n5430), .A2(n5383), .ZN(n5431) );
  XNOR2_X1 U5314 ( .A(n5376), .B(SI_11_), .ZN(n5398) );
  AOI21_X1 U5315 ( .B1(n5349), .B2(n5348), .A(n4673), .ZN(n5373) );
  INV_X1 U5316 ( .A(n5350), .ZN(n4673) );
  NAND2_X1 U5317 ( .A1(n5299), .A2(n5298), .ZN(n4923) );
  INV_X1 U5318 ( .A(n5297), .ZN(n5298) );
  XNOR2_X1 U5319 ( .A(n5300), .B(SI_7_), .ZN(n5297) );
  XNOR2_X1 U5320 ( .A(n5287), .B(SI_6_), .ZN(n5284) );
  XNOR2_X1 U5321 ( .A(n5236), .B(SI_4_), .ZN(n5233) );
  NAND2_X1 U5322 ( .A1(n7558), .A2(n5274), .ZN(n7646) );
  NOR2_X1 U5323 ( .A1(n5733), .A2(n4855), .ZN(n4854) );
  NAND2_X1 U5324 ( .A1(n4612), .A2(n4611), .ZN(n9149) );
  NOR2_X1 U5325 ( .A1(n5642), .A2(n4509), .ZN(n4611) );
  AND2_X1 U5326 ( .A1(n4842), .A2(n4843), .ZN(n4841) );
  AND2_X1 U5327 ( .A1(n5415), .A2(n5397), .ZN(n5421) );
  NAND2_X1 U5328 ( .A1(n7558), .A2(n4866), .ZN(n7782) );
  NOR2_X1 U5329 ( .A1(n5323), .A2(n4867), .ZN(n4866) );
  INV_X1 U5330 ( .A(n5274), .ZN(n4867) );
  INV_X1 U5331 ( .A(n5587), .ZN(n4846) );
  AOI21_X1 U5332 ( .B1(n9179), .B2(n9178), .A(n5628), .ZN(n5641) );
  XNOR2_X1 U5333 ( .A(n5576), .B(n10474), .ZN(n7584) );
  AND2_X1 U5334 ( .A1(n4847), .A2(n5545), .ZN(n4620) );
  NAND2_X1 U5335 ( .A1(n4836), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5751) );
  NAND2_X1 U5336 ( .A1(n5118), .A2(n4835), .ZN(n4836) );
  AND2_X1 U5337 ( .A1(n5119), .A2(n5117), .ZN(n4835) );
  AND2_X1 U5338 ( .A1(n5727), .A2(n5726), .ZN(n9243) );
  AND3_X1 U5339 ( .A1(n5669), .A2(n5668), .A3(n5667), .ZN(n9155) );
  AND3_X1 U5340 ( .A1(n5134), .A2(n5133), .A3(n5132), .ZN(n9181) );
  AND4_X1 U5341 ( .A1(n5474), .A2(n5473), .A3(n5472), .A4(n5471), .ZN(n8249)
         );
  OR2_X1 U5342 ( .A1(n4498), .A2(n5190), .ZN(n5192) );
  OR2_X1 U5343 ( .A1(n8186), .A2(n8185), .ZN(n4597) );
  NAND2_X1 U5344 ( .A1(n4597), .A2(n4596), .ZN(n4595) );
  NAND2_X1 U5345 ( .A1(n7709), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4596) );
  OR2_X1 U5346 ( .A1(n7883), .A2(n7882), .ZN(n4584) );
  NAND2_X1 U5347 ( .A1(n8122), .A2(n8123), .ZN(n8121) );
  NAND2_X1 U5348 ( .A1(n4600), .A2(n4599), .ZN(n7717) );
  INV_X1 U5349 ( .A(n7857), .ZN(n4599) );
  NAND2_X1 U5350 ( .A1(n7859), .A2(n7858), .ZN(n4600) );
  NAND2_X1 U5351 ( .A1(n4602), .A2(n4601), .ZN(n7859) );
  INV_X1 U5352 ( .A(n7871), .ZN(n4601) );
  INV_X1 U5353 ( .A(n7872), .ZN(n4602) );
  INV_X1 U5354 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5400) );
  NAND2_X1 U5355 ( .A1(n7834), .A2(n4868), .ZN(n7836) );
  OR2_X1 U5356 ( .A1(n7835), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4868) );
  OR2_X1 U5357 ( .A1(n7722), .A2(n7721), .ZN(n4606) );
  AND2_X1 U5358 ( .A1(n4608), .A2(n4607), .ZN(n9299) );
  NAND2_X1 U5359 ( .A1(n9296), .A2(n8383), .ZN(n4607) );
  NOR2_X1 U5360 ( .A1(n8930), .A2(n4792), .ZN(n4790) );
  NAND2_X1 U5361 ( .A1(n9112), .A2(n9113), .ZN(n8921) );
  NAND2_X1 U5362 ( .A1(n4925), .A2(n4924), .ZN(n9375) );
  AOI21_X1 U5363 ( .B1(n4926), .B2(n4929), .A(n9099), .ZN(n4924) );
  OR2_X1 U5364 ( .A1(n9439), .A2(n9155), .ZN(n9417) );
  NOR2_X2 U5365 ( .A1(n9438), .A2(n9427), .ZN(n9414) );
  NOR2_X1 U5366 ( .A1(n9450), .A2(n6780), .ZN(n9437) );
  INV_X1 U5367 ( .A(n9452), .ZN(n9446) );
  OR2_X1 U5368 ( .A1(n9468), .A2(n9181), .ZN(n8980) );
  XNOR2_X1 U5369 ( .A(n9159), .B(n9258), .ZN(n9452) );
  OAI21_X1 U5370 ( .B1(n5049), .B2(n5050), .A(n8981), .ZN(n5048) );
  INV_X1 U5371 ( .A(n6810), .ZN(n5049) );
  NAND2_X1 U5372 ( .A1(n9497), .A2(n4952), .ZN(n4951) );
  INV_X1 U5373 ( .A(n6779), .ZN(n4952) );
  AND2_X1 U5374 ( .A1(n8980), .A2(n8983), .ZN(n9463) );
  OR2_X1 U5375 ( .A1(n9494), .A2(n9495), .ZN(n4953) );
  NAND2_X1 U5376 ( .A1(n5083), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5617) );
  INV_X1 U5377 ( .A(n5577), .ZN(n5083) );
  OR2_X1 U5378 ( .A1(n9559), .A2(n8341), .ZN(n9527) );
  NAND2_X1 U5379 ( .A1(n4938), .A2(n4937), .ZN(n9534) );
  AOI21_X1 U5380 ( .B1(n4939), .B2(n9063), .A(n4507), .ZN(n4937) );
  NAND2_X1 U5381 ( .A1(n5081), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5557) );
  AND2_X1 U5382 ( .A1(n9554), .A2(n4540), .ZN(n4939) );
  OR2_X1 U5383 ( .A1(n8423), .A2(n9063), .ZN(n4941) );
  AND2_X1 U5384 ( .A1(n9063), .A2(n9061), .ZN(n5055) );
  NAND2_X1 U5385 ( .A1(n8353), .A2(n9061), .ZN(n8416) );
  NAND2_X1 U5386 ( .A1(n8354), .A2(n9059), .ZN(n8353) );
  NAND2_X1 U5387 ( .A1(n8263), .A2(n5056), .ZN(n8165) );
  AND2_X1 U5388 ( .A1(n9054), .A2(n6804), .ZN(n5056) );
  AND2_X1 U5389 ( .A1(n9056), .A2(n9057), .ZN(n9054) );
  OR2_X1 U5390 ( .A1(n8261), .A2(n9055), .ZN(n8263) );
  OR2_X1 U5391 ( .A1(n5336), .A2(n5335), .ZN(n5359) );
  AND2_X1 U5392 ( .A1(n9033), .A2(n9028), .ZN(n8951) );
  OR2_X1 U5393 ( .A1(n9274), .A2(n10501), .ZN(n9017) );
  OR2_X1 U5394 ( .A1(n9276), .A2(n10494), .ZN(n8997) );
  NAND2_X1 U5395 ( .A1(n9276), .A2(n10494), .ZN(n7443) );
  AND2_X1 U5396 ( .A1(n10467), .A2(n8942), .ZN(n9541) );
  AND2_X1 U5397 ( .A1(n5801), .A2(n5800), .ZN(n9245) );
  NAND2_X1 U5398 ( .A1(n5436), .A2(n6148), .ZN(n5163) );
  OR2_X1 U5399 ( .A1(n9281), .A2(n7655), .ZN(n7498) );
  NAND2_X1 U5400 ( .A1(n8927), .A2(n8926), .ZN(n9340) );
  INV_X1 U5401 ( .A(n9541), .ZN(n10520) );
  NAND2_X1 U5402 ( .A1(n9695), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5108) );
  INV_X1 U5403 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n4865) );
  INV_X1 U5404 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4610) );
  NAND2_X1 U5405 ( .A1(n5199), .A2(n5144), .ZN(n5159) );
  AND2_X1 U5406 ( .A1(n5006), .A2(n4642), .ZN(n4641) );
  INV_X1 U5407 ( .A(n9733), .ZN(n4642) );
  XNOR2_X1 U5408 ( .A(n6489), .B(n6660), .ZN(n7067) );
  AND2_X1 U5409 ( .A1(n5010), .A2(n5008), .ZN(n4640) );
  NAND2_X1 U5410 ( .A1(n9741), .A2(n9742), .ZN(n9740) );
  AND2_X1 U5411 ( .A1(n6670), .A2(n6669), .ZN(n9752) );
  NAND2_X1 U5412 ( .A1(n5010), .A2(n5009), .ZN(n9754) );
  INV_X1 U5413 ( .A(n4644), .ZN(n9753) );
  AND2_X1 U5414 ( .A1(n6480), .A2(n6479), .ZN(n7045) );
  OR2_X1 U5415 ( .A1(n6574), .A2(n4629), .ZN(n4628) );
  INV_X1 U5416 ( .A(n6578), .ZN(n4629) );
  NAND2_X1 U5417 ( .A1(n5001), .A2(n4999), .ZN(n9773) );
  AOI21_X1 U5418 ( .B1(n5002), .B2(n5005), .A(n5000), .ZN(n4999) );
  INV_X1 U5419 ( .A(n6656), .ZN(n5000) );
  OR2_X1 U5420 ( .A1(n6657), .A2(n6656), .ZN(n9774) );
  NAND2_X1 U5421 ( .A1(n4994), .A2(n4995), .ZN(n7665) );
  INV_X1 U5422 ( .A(n4996), .ZN(n4995) );
  OAI21_X1 U5423 ( .B1(n6561), .B2(n4997), .A(n7638), .ZN(n4996) );
  NOR2_X1 U5424 ( .A1(n6120), .A2(n8817), .ZN(n6108) );
  NOR2_X1 U5425 ( .A1(n7057), .A2(n7058), .ZN(n7056) );
  XNOR2_X1 U5426 ( .A(n6915), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n6947) );
  OR2_X1 U5427 ( .A1(n6948), .A2(n6947), .ZN(n4889) );
  OR2_X1 U5428 ( .A1(n10315), .A2(n10316), .ZN(n4894) );
  AND2_X1 U5429 ( .A1(n4894), .A2(n4893), .ZN(n6963) );
  NAND2_X1 U5430 ( .A1(n10311), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4893) );
  NAND2_X1 U5431 ( .A1(n4572), .A2(n4571), .ZN(n4892) );
  INV_X1 U5432 ( .A(n6962), .ZN(n4571) );
  INV_X1 U5433 ( .A(n6963), .ZN(n4572) );
  OR2_X1 U5434 ( .A1(n7193), .A2(n4897), .ZN(n4574) );
  NOR2_X1 U5435 ( .A1(n7192), .A2(n4898), .ZN(n4897) );
  INV_X1 U5436 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n4898) );
  NAND2_X1 U5437 ( .A1(n4567), .A2(n4556), .ZN(n7433) );
  OR2_X1 U5438 ( .A1(n7429), .A2(n7430), .ZN(n4567) );
  OR2_X1 U5439 ( .A1(n7433), .A2(n7432), .ZN(n4902) );
  NOR2_X1 U5440 ( .A1(n8280), .A2(n8279), .ZN(n9833) );
  OR2_X1 U5441 ( .A1(n9837), .A2(n9836), .ZN(n4569) );
  AND2_X1 U5442 ( .A1(n6255), .A2(n6844), .ZN(n6263) );
  NAND2_X1 U5443 ( .A1(n5849), .A2(n5848), .ZN(n8515) );
  NOR2_X1 U5444 ( .A1(n10065), .A2(n9938), .ZN(n9928) );
  NAND2_X1 U5445 ( .A1(n4564), .A2(n4563), .ZN(n9938) );
  OR2_X1 U5446 ( .A1(n10072), .A2(n9814), .ZN(n8488) );
  OR2_X1 U5447 ( .A1(n10079), .A2(n9990), .ZN(n9959) );
  NAND2_X1 U5448 ( .A1(n9970), .A2(n8502), .ZN(n9960) );
  NOR2_X1 U5449 ( .A1(n8486), .A2(n4978), .ZN(n4977) );
  INV_X1 U5450 ( .A(n5062), .ZN(n4978) );
  AOI21_X1 U5451 ( .B1(n6353), .B2(n4754), .A(n4753), .ZN(n4752) );
  INV_X1 U5452 ( .A(n8498), .ZN(n4753) );
  INV_X1 U5453 ( .A(n10035), .ZN(n4754) );
  OR2_X1 U5454 ( .A1(n10034), .A2(n6190), .ZN(n4748) );
  NAND2_X1 U5455 ( .A1(n4751), .A2(n4749), .ZN(n10004) );
  AND2_X1 U5456 ( .A1(n4750), .A2(n10005), .ZN(n4749) );
  NAND2_X1 U5457 ( .A1(n10034), .A2(n4752), .ZN(n4751) );
  NAND2_X1 U5458 ( .A1(n4752), .A2(n6190), .ZN(n4750) );
  OR2_X1 U5459 ( .A1(n10018), .A2(n9728), .ZN(n5062) );
  OR2_X1 U5460 ( .A1(n10092), .A2(n10037), .ZN(n8484) );
  AND2_X1 U5461 ( .A1(n8500), .A2(n6269), .ZN(n10005) );
  NAND2_X1 U5462 ( .A1(n10034), .A2(n10035), .ZN(n10033) );
  NAND2_X1 U5463 ( .A1(n4576), .A2(n8454), .ZN(n8457) );
  NAND2_X1 U5464 ( .A1(n4578), .A2(n4577), .ZN(n4576) );
  OR2_X1 U5465 ( .A1(n8408), .A2(n8407), .ZN(n4578) );
  NAND2_X1 U5466 ( .A1(n4579), .A2(n8311), .ZN(n8408) );
  NAND2_X1 U5467 ( .A1(n4760), .A2(n4580), .ZN(n4579) );
  INV_X1 U5468 ( .A(n8312), .ZN(n4580) );
  AND2_X1 U5469 ( .A1(n8332), .A2(n9817), .ZN(n4984) );
  NAND2_X1 U5470 ( .A1(n4982), .A2(n4983), .ZN(n4981) );
  INV_X1 U5471 ( .A(n8150), .ZN(n4983) );
  INV_X1 U5472 ( .A(n4967), .ZN(n4966) );
  OAI22_X1 U5473 ( .A1(n4968), .A2(n7315), .B1(n9824), .B2(n7547), .ZN(n4967)
         );
  INV_X1 U5474 ( .A(n7316), .ZN(n4970) );
  NAND2_X1 U5475 ( .A1(n7238), .A2(n4530), .ZN(n7260) );
  NAND2_X1 U5476 ( .A1(n7219), .A2(n7272), .ZN(n7289) );
  INV_X1 U5477 ( .A(n7215), .ZN(n7211) );
  NAND2_X1 U5478 ( .A1(n8515), .A2(n10133), .ZN(n4916) );
  INV_X1 U5479 ( .A(n7924), .ZN(n7925) );
  XNOR2_X1 U5480 ( .A(n5709), .B(n5708), .ZN(n8177) );
  XNOR2_X1 U5481 ( .A(n5693), .B(n5692), .ZN(n8090) );
  NAND2_X1 U5482 ( .A1(n4828), .A2(n4829), .ZN(n5693) );
  NAND2_X1 U5483 ( .A1(n5658), .A2(n4831), .ZN(n4828) );
  XNOR2_X1 U5484 ( .A(n4570), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6915) );
  NAND2_X1 U5485 ( .A1(n6171), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4570) );
  AND2_X1 U5486 ( .A1(n6172), .A2(n6171), .ZN(n7052) );
  AND2_X1 U5487 ( .A1(n5748), .A2(n5747), .ZN(n9145) );
  NAND2_X1 U5488 ( .A1(n7596), .A2(n5188), .ZN(n7417) );
  XNOR2_X1 U5489 ( .A(n5169), .B(n7584), .ZN(n7371) );
  AND2_X1 U5490 ( .A1(n7657), .A2(n5157), .ZN(n7372) );
  NAND2_X1 U5491 ( .A1(n5500), .A2(n5499), .ZN(n9066) );
  AND2_X1 U5492 ( .A1(n9211), .A2(n5232), .ZN(n7530) );
  NAND2_X1 U5493 ( .A1(n5600), .A2(n5599), .ZN(n9503) );
  NAND2_X1 U5494 ( .A1(n4696), .A2(n4694), .ZN(n9127) );
  NAND2_X1 U5495 ( .A1(n4697), .A2(n9126), .ZN(n4696) );
  NAND2_X1 U5496 ( .A1(n4695), .A2(n9125), .ZN(n4694) );
  OR2_X1 U5497 ( .A1(n10450), .A2(n5803), .ZN(n9130) );
  XNOR2_X1 U5498 ( .A(n5751), .B(P2_IR_REG_22__SCAN_IN), .ZN(n9131) );
  OR2_X1 U5499 ( .A1(n7833), .A2(n7832), .ZN(n4604) );
  AND2_X1 U5500 ( .A1(n4606), .A2(n4605), .ZN(n7833) );
  NAND2_X1 U5501 ( .A1(n7831), .A2(n5443), .ZN(n4605) );
  OR2_X1 U5502 ( .A1(n8386), .A2(n8385), .ZN(n4608) );
  OAI21_X1 U5503 ( .B1(n9336), .B2(n10444), .A(n4593), .ZN(n4592) );
  NAND2_X1 U5504 ( .A1(n4588), .A2(n4587), .ZN(n4586) );
  NAND2_X1 U5505 ( .A1(n9336), .A2(n10439), .ZN(n4588) );
  NAND2_X1 U5506 ( .A1(n9401), .A2(n9403), .ZN(n9400) );
  NAND2_X1 U5507 ( .A1(n9424), .A2(n6782), .ZN(n9401) );
  OAI21_X1 U5508 ( .B1(n9405), .B2(n9553), .A(n9404), .ZN(n9589) );
  CLKBUF_X1 U5509 ( .A(n5153), .Z(n9522) );
  AND2_X1 U5510 ( .A1(n5023), .A2(n4548), .ZN(n5021) );
  AOI21_X1 U5511 ( .B1(n5026), .B2(n5027), .A(n9795), .ZN(n5023) );
  NAND2_X1 U5512 ( .A1(n5027), .A2(n5028), .ZN(n5024) );
  INV_X1 U5513 ( .A(n6730), .ZN(n5020) );
  NAND2_X1 U5514 ( .A1(n4643), .A2(n4641), .ZN(n9732) );
  AND4_X1 U5515 ( .A1(n5884), .A2(n5883), .A3(n5882), .A4(n5881), .ZN(n9973)
         );
  AND4_X1 U5516 ( .A1(n5930), .A2(n5929), .A3(n5928), .A4(n5927), .ZN(n9789)
         );
  NAND2_X1 U5517 ( .A1(n4520), .A2(n10292), .ZN(n10291) );
  AND2_X1 U5518 ( .A1(n6855), .A2(n6854), .ZN(n7193) );
  XNOR2_X1 U5519 ( .A(n9833), .B(n9832), .ZN(n8282) );
  AOI21_X1 U5520 ( .B1(n9894), .B2(n4886), .A(n9902), .ZN(n4885) );
  OR2_X1 U5521 ( .A1(n9898), .A2(n9895), .ZN(n4886) );
  OAI21_X1 U5522 ( .B1(n9901), .B2(n9900), .A(n4883), .ZN(n4882) );
  NOR2_X1 U5523 ( .A1(n4511), .A2(n10310), .ZN(n4883) );
  XNOR2_X1 U5524 ( .A(n8508), .B(n8492), .ZN(n8513) );
  AOI22_X1 U5525 ( .A1(n8490), .A2(n10054), .B1(n9908), .B2(n9813), .ZN(n8511)
         );
  NAND2_X1 U5526 ( .A1(n9918), .A2(n8491), .ZN(n8493) );
  NAND2_X1 U5527 ( .A1(n10065), .A2(n8490), .ZN(n8491) );
  NAND2_X1 U5528 ( .A1(n4772), .A2(n4770), .ZN(n10063) );
  AOI21_X1 U5529 ( .B1(n9964), .B2(n10054), .A(n4771), .ZN(n4770) );
  OAI21_X1 U5530 ( .B1(n9925), .B2(n9924), .A(n10343), .ZN(n4772) );
  NOR2_X1 U5531 ( .A1(n9927), .A2(n10338), .ZN(n4771) );
  NAND2_X1 U5532 ( .A1(n4741), .A2(n6301), .ZN(n4740) );
  OR2_X1 U5533 ( .A1(n7164), .A2(n6422), .ZN(n4741) );
  NAND2_X1 U5534 ( .A1(n4688), .A2(n4686), .ZN(n9022) );
  NOR2_X1 U5535 ( .A1(n9016), .A2(n4687), .ZN(n4686) );
  OR2_X1 U5536 ( .A1(n6309), .A2(n6717), .ZN(n4731) );
  AND2_X1 U5537 ( .A1(n4726), .A2(n6314), .ZN(n4725) );
  NOR2_X1 U5538 ( .A1(n7762), .A2(n4727), .ZN(n4726) );
  INV_X1 U5539 ( .A(n6313), .ZN(n4727) );
  NAND2_X1 U5540 ( .A1(n9042), .A2(n4684), .ZN(n9040) );
  NOR2_X1 U5541 ( .A1(n4685), .A2(n5045), .ZN(n4684) );
  INV_X1 U5542 ( .A(n9045), .ZN(n4685) );
  NOR2_X1 U5543 ( .A1(n4722), .A2(n6717), .ZN(n4718) );
  NOR2_X1 U5544 ( .A1(n4724), .A2(n4723), .ZN(n4722) );
  INV_X1 U5545 ( .A(n8454), .ZN(n4724) );
  NOR2_X1 U5546 ( .A1(n9750), .A2(n9816), .ZN(n4723) );
  AOI21_X1 U5547 ( .B1(n4577), .B2(n10119), .A(n6373), .ZN(n4721) );
  OAI21_X1 U5548 ( .B1(n4703), .B2(n4702), .A(n9062), .ZN(n9064) );
  NAND2_X1 U5549 ( .A1(n9059), .A2(n9058), .ZN(n4702) );
  AOI21_X1 U5550 ( .B1(n9079), .B2(n9078), .A(n4678), .ZN(n4677) );
  INV_X1 U5551 ( .A(n9082), .ZN(n4678) );
  AOI21_X1 U5552 ( .B1(n6345), .B2(n4715), .A(n6344), .ZN(n6350) );
  INV_X1 U5553 ( .A(n4716), .ZN(n4715) );
  INV_X1 U5554 ( .A(n9089), .ZN(n4712) );
  NAND2_X1 U5555 ( .A1(n9090), .A2(n9089), .ZN(n4714) );
  INV_X1 U5556 ( .A(n9083), .ZN(n9088) );
  NAND2_X1 U5557 ( .A1(n7443), .A2(n8987), .ZN(n8985) );
  OAI211_X1 U5558 ( .C1(n6359), .C2(n6373), .A(n6361), .B(n4745), .ZN(n6379)
         );
  INV_X1 U5559 ( .A(n5378), .ZN(n4669) );
  AOI21_X1 U5560 ( .B1(n4709), .B2(n9095), .A(n4708), .ZN(n9100) );
  INV_X1 U5561 ( .A(n8985), .ZN(n8989) );
  NOR2_X1 U5562 ( .A1(n9372), .A2(n9393), .ZN(n4794) );
  NAND2_X1 U5563 ( .A1(n4672), .A2(n9817), .ZN(n6336) );
  NOR2_X1 U5564 ( .A1(n10084), .A2(n10087), .ZN(n4915) );
  AOI21_X1 U5565 ( .B1(n5738), .B2(n4804), .A(n4803), .ZN(n4802) );
  OAI21_X1 U5566 ( .B1(n4805), .B2(n5815), .A(n6229), .ZN(n4803) );
  NOR2_X1 U5567 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5825) );
  NAND2_X1 U5568 ( .A1(n5547), .A2(n5529), .ZN(n4818) );
  NOR2_X1 U5569 ( .A1(n4818), .A2(n4814), .ZN(n4813) );
  INV_X1 U5570 ( .A(n5492), .ZN(n4814) );
  NOR2_X1 U5571 ( .A1(n5482), .A2(n4808), .ZN(n4807) );
  INV_X1 U5572 ( .A(n5458), .ZN(n4808) );
  NAND2_X1 U5573 ( .A1(n5431), .A2(n5430), .ZN(n4811) );
  INV_X1 U5574 ( .A(n4668), .ZN(n4667) );
  OAI21_X1 U5575 ( .B1(n4670), .B2(n4669), .A(n5430), .ZN(n4668) );
  NAND2_X1 U5576 ( .A1(n4667), .A2(n4669), .ZN(n4665) );
  NOR2_X1 U5577 ( .A1(n5379), .A2(n4671), .ZN(n4670) );
  INV_X1 U5578 ( .A(n5374), .ZN(n4671) );
  INV_X1 U5579 ( .A(n5398), .ZN(n5379) );
  INV_X1 U5580 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4575) );
  INV_X1 U5581 ( .A(n5480), .ZN(n4850) );
  NAND2_X1 U5582 ( .A1(n9189), .A2(n9188), .ZN(n4861) );
  INV_X1 U5583 ( .A(n9123), .ZN(n4699) );
  NOR2_X1 U5584 ( .A1(n8970), .A2(n4701), .ZN(n4700) );
  NAND2_X1 U5585 ( .A1(n9115), .A2(n9114), .ZN(n4701) );
  OR2_X1 U5586 ( .A1(n5355), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5386) );
  NAND2_X1 U5587 ( .A1(n9459), .A2(n5042), .ZN(n5041) );
  NOR2_X1 U5588 ( .A1(n9446), .A2(n5043), .ZN(n5042) );
  INV_X1 U5589 ( .A(n8980), .ZN(n5043) );
  NAND2_X1 U5590 ( .A1(n9672), .A2(n4789), .ZN(n4788) );
  NOR2_X1 U5591 ( .A1(n9468), .A2(n9486), .ZN(n4789) );
  OR2_X1 U5592 ( .A1(n9503), .A2(n9180), .ZN(n9478) );
  NOR2_X1 U5593 ( .A1(n9497), .A2(n5051), .ZN(n5050) );
  NAND2_X1 U5594 ( .A1(n5080), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5511) );
  OR2_X1 U5595 ( .A1(n5469), .A2(n5468), .ZN(n5509) );
  OR2_X1 U5596 ( .A1(n8956), .A2(n7964), .ZN(n6772) );
  NOR2_X1 U5597 ( .A1(n6765), .A2(n7957), .ZN(n4781) );
  NOR2_X1 U5598 ( .A1(n6798), .A2(n7737), .ZN(n6799) );
  NOR2_X1 U5599 ( .A1(n7571), .A2(n7581), .ZN(n7513) );
  OR2_X1 U5600 ( .A1(n9520), .A2(n9503), .ZN(n9501) );
  OR2_X1 U5601 ( .A1(n9519), .A2(n9626), .ZN(n9520) );
  NOR2_X1 U5602 ( .A1(n9560), .A2(n9559), .ZN(n9542) );
  AND2_X1 U5603 ( .A1(n8034), .A2(n10512), .ZN(n8036) );
  AND2_X1 U5604 ( .A1(n10471), .A2(n10482), .ZN(n7472) );
  AND2_X1 U5605 ( .A1(n5118), .A2(n5117), .ZN(n5123) );
  OR2_X1 U5606 ( .A1(n5306), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5355) );
  AND4_X1 U5607 ( .A1(n5176), .A2(n5031), .A3(n5086), .A4(n4837), .ZN(n5261)
         );
  INV_X1 U5608 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n4837) );
  INV_X1 U5609 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5086) );
  INV_X1 U5610 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4609) );
  AND2_X1 U5611 ( .A1(n5003), .A2(n6651), .ZN(n5002) );
  NAND2_X1 U5612 ( .A1(n9725), .A2(n5004), .ZN(n5003) );
  INV_X1 U5613 ( .A(n9725), .ZN(n5005) );
  INV_X1 U5614 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5832) );
  AND2_X1 U5615 ( .A1(n4900), .A2(n4899), .ZN(n8278) );
  NAND2_X1 U5616 ( .A1(n8015), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4899) );
  OR2_X1 U5617 ( .A1(n8515), .A2(n9927), .ZN(n6390) );
  NAND2_X1 U5618 ( .A1(n10065), .A2(n9945), .ZN(n8506) );
  OR2_X1 U5619 ( .A1(n10065), .A2(n9945), .ZN(n6380) );
  NAND2_X1 U5620 ( .A1(n9980), .A2(n4915), .ZN(n4914) );
  AOI21_X1 U5621 ( .B1(n4662), .B2(n4971), .A(n4661), .ZN(n4660) );
  INV_X1 U5622 ( .A(n9971), .ZN(n4661) );
  INV_X1 U5623 ( .A(n4974), .ZN(n4662) );
  INV_X1 U5624 ( .A(n4971), .ZN(n4663) );
  OR2_X1 U5625 ( .A1(n10092), .A2(n9728), .ZN(n8498) );
  NAND2_X1 U5626 ( .A1(n4653), .A2(n8401), .ZN(n4652) );
  OR2_X1 U5627 ( .A1(n10108), .A2(n9789), .ZN(n6346) );
  NAND2_X1 U5628 ( .A1(n8332), .A2(n8316), .ZN(n8311) );
  NAND2_X1 U5629 ( .A1(n6336), .A2(n8311), .ZN(n4982) );
  NAND2_X1 U5630 ( .A1(n8144), .A2(n7924), .ZN(n4765) );
  INV_X1 U5631 ( .A(n8143), .ZN(n4766) );
  OR2_X1 U5632 ( .A1(n4960), .A2(n4959), .ZN(n4958) );
  INV_X1 U5633 ( .A(n7755), .ZN(n4959) );
  NOR2_X1 U5634 ( .A1(n10238), .A2(n10237), .ZN(n4910) );
  OR2_X1 U5635 ( .A1(n7399), .A2(n4969), .ZN(n4968) );
  INV_X1 U5636 ( .A(n7397), .ZN(n4969) );
  INV_X1 U5637 ( .A(n4968), .ZN(n4965) );
  NOR2_X1 U5638 ( .A1(n10014), .A2(n4913), .ZN(n9991) );
  INV_X1 U5639 ( .A(n4915), .ZN(n4913) );
  INV_X1 U5640 ( .A(n6719), .ZN(n6715) );
  NAND2_X1 U5641 ( .A1(n10243), .A2(n7760), .ZN(n10246) );
  INV_X1 U5642 ( .A(n4830), .ZN(n4829) );
  OAI21_X1 U5643 ( .B1(n5673), .B2(n5655), .A(n5677), .ZN(n4830) );
  NOR2_X1 U5644 ( .A1(n4832), .A2(n5673), .ZN(n4831) );
  INV_X1 U5645 ( .A(n5657), .ZN(n4832) );
  NAND2_X1 U5646 ( .A1(n5921), .A2(n5834), .ZN(n6257) );
  INV_X1 U5647 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5983) );
  NOR2_X1 U5648 ( .A1(n5326), .A2(n4922), .ZN(n4921) );
  INV_X1 U5649 ( .A(n5301), .ZN(n4922) );
  NAND2_X1 U5650 ( .A1(n5329), .A2(SI_9_), .ZN(n5350) );
  OAI21_X1 U5651 ( .B1(n6889), .B2(n5215), .A(n5214), .ZN(n5236) );
  NAND2_X1 U5652 ( .A1(n6889), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5214) );
  XNOR2_X1 U5653 ( .A(n5198), .B(SI_2_), .ZN(n5195) );
  INV_X1 U5654 ( .A(n5173), .ZN(n4917) );
  NOR2_X1 U5655 ( .A1(n6101), .A2(n6113), .ZN(n6170) );
  XNOR2_X1 U5656 ( .A(n4656), .B(SI_1_), .ZN(n5172) );
  NAND2_X1 U5657 ( .A1(n8048), .A2(n4517), .ZN(n4621) );
  OR2_X1 U5658 ( .A1(n5445), .A2(n5444), .ZN(n5469) );
  INV_X1 U5659 ( .A(n5422), .ZN(n5425) );
  NAND2_X1 U5660 ( .A1(n5576), .A2(n4618), .ZN(n4615) );
  NAND2_X1 U5661 ( .A1(n4619), .A2(n4617), .ZN(n4616) );
  NOR2_X1 U5662 ( .A1(n5576), .A2(n4618), .ZN(n4617) );
  INV_X1 U5663 ( .A(n5618), .ZN(n5085) );
  NAND2_X1 U5664 ( .A1(n5690), .A2(n4862), .ZN(n4860) );
  NAND2_X1 U5665 ( .A1(n8920), .A2(n5480), .ZN(n8295) );
  NOR2_X1 U5666 ( .A1(n9343), .A2(n8931), .ZN(n5038) );
  INV_X1 U5667 ( .A(n5035), .ZN(n5034) );
  NOR2_X1 U5668 ( .A1(n9644), .A2(n9343), .ZN(n9121) );
  XNOR2_X1 U5669 ( .A(n4799), .B(n9522), .ZN(n8966) );
  NAND2_X1 U5670 ( .A1(n8973), .A2(n4800), .ZN(n4799) );
  NOR2_X1 U5671 ( .A1(n9121), .A2(n4801), .ZN(n4800) );
  NAND2_X1 U5672 ( .A1(n4522), .A2(n9116), .ZN(n4801) );
  INV_X1 U5673 ( .A(n4697), .ZN(n4695) );
  AND3_X1 U5674 ( .A1(n5689), .A2(n5688), .A3(n5687), .ZN(n9244) );
  AND4_X1 U5675 ( .A1(n5582), .A2(n5581), .A3(n5580), .A4(n5579), .ZN(n8464)
         );
  AND4_X1 U5676 ( .A1(n5515), .A2(n5514), .A3(n5513), .A4(n5512), .ZN(n8303)
         );
  AND4_X1 U5677 ( .A1(n5393), .A2(n5392), .A3(n5391), .A4(n5390), .ZN(n8051)
         );
  AND4_X1 U5678 ( .A1(n5414), .A2(n5413), .A3(n5412), .A4(n5411), .ZN(n7992)
         );
  NAND2_X1 U5679 ( .A1(n4584), .A2(n4554), .ZN(n8122) );
  OR2_X1 U5680 ( .A1(n8107), .A2(n8106), .ZN(n4874) );
  AND2_X1 U5681 ( .A1(n4874), .A2(n4873), .ZN(n9283) );
  NAND2_X1 U5682 ( .A1(n7698), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4873) );
  AND2_X1 U5683 ( .A1(n4604), .A2(n4603), .ZN(n8379) );
  NAND2_X1 U5684 ( .A1(n8086), .A2(n5467), .ZN(n4603) );
  NAND2_X1 U5685 ( .A1(n9313), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4877) );
  OR2_X1 U5686 ( .A1(n5742), .A2(n5741), .ZN(n9353) );
  INV_X1 U5687 ( .A(n9436), .ZN(n9432) );
  AND2_X1 U5688 ( .A1(n5041), .A2(n4518), .ZN(n9416) );
  NAND2_X1 U5689 ( .A1(n9417), .A2(n9096), .ZN(n9436) );
  NAND2_X1 U5690 ( .A1(n4947), .A2(n4943), .ZN(n9451) );
  INV_X1 U5691 ( .A(n4944), .ZN(n4943) );
  OAI21_X1 U5692 ( .B1(n4946), .B2(n9463), .A(n4945), .ZN(n4944) );
  NOR2_X1 U5693 ( .A1(n9501), .A2(n9486), .ZN(n9485) );
  NOR2_X1 U5694 ( .A1(n9501), .A2(n4787), .ZN(n9466) );
  INV_X1 U5695 ( .A(n4789), .ZN(n4787) );
  NAND2_X1 U5696 ( .A1(n9516), .A2(n9515), .ZN(n5052) );
  AND2_X1 U5697 ( .A1(n5575), .A2(n5574), .ZN(n6777) );
  AND2_X1 U5698 ( .A1(n9076), .A2(n9080), .ZN(n9515) );
  NAND2_X1 U5699 ( .A1(n9557), .A2(n6808), .ZN(n9529) );
  OR2_X1 U5700 ( .A1(n5557), .A2(n5082), .ZN(n5577) );
  AOI21_X1 U5701 ( .B1(n5055), .B2(n8351), .A(n4537), .ZN(n5053) );
  INV_X1 U5702 ( .A(n5055), .ZN(n5054) );
  OR2_X1 U5703 ( .A1(n8358), .A2(n9066), .ZN(n9560) );
  NAND2_X1 U5704 ( .A1(n4931), .A2(n4930), .ZN(n8352) );
  AOI21_X1 U5705 ( .B1(n4932), .B2(n4935), .A(n4534), .ZN(n4930) );
  AND2_X1 U5706 ( .A1(n8036), .A2(n4777), .ZN(n8357) );
  NOR2_X1 U5707 ( .A1(n8917), .A2(n4779), .ZN(n4777) );
  NAND2_X1 U5708 ( .A1(n8036), .A2(n4781), .ZN(n8268) );
  NAND2_X1 U5709 ( .A1(n5046), .A2(n5044), .ZN(n7967) );
  NOR2_X1 U5710 ( .A1(n6803), .A2(n5045), .ZN(n5044) );
  NAND2_X1 U5711 ( .A1(n4920), .A2(n4919), .ZN(n7964) );
  INV_X1 U5712 ( .A(n6770), .ZN(n4919) );
  NAND2_X1 U5713 ( .A1(n7907), .A2(n8953), .ZN(n4920) );
  OR2_X1 U5714 ( .A1(n8022), .A2(n6769), .ZN(n7907) );
  AND2_X1 U5715 ( .A1(n8025), .A2(n8021), .ZN(n8022) );
  NOR2_X1 U5716 ( .A1(n4514), .A2(n8898), .ZN(n8034) );
  NAND2_X1 U5717 ( .A1(n7513), .A2(n7633), .ZN(n7744) );
  AND2_X1 U5718 ( .A1(n9017), .A2(n9014), .ZN(n8945) );
  NAND2_X1 U5719 ( .A1(n4796), .A2(n4795), .ZN(n7571) );
  NOR2_X1 U5720 ( .A1(n9214), .A2(n7524), .ZN(n4795) );
  INV_X1 U5721 ( .A(n7618), .ZN(n4796) );
  AND2_X1 U5722 ( .A1(n7383), .A2(n8996), .ZN(n7614) );
  NAND2_X1 U5723 ( .A1(n8997), .A2(n7443), .ZN(n8940) );
  NAND2_X1 U5724 ( .A1(n8996), .A2(n8988), .ZN(n8943) );
  NAND2_X1 U5725 ( .A1(n7466), .A2(n7467), .ZN(n7465) );
  NAND2_X1 U5726 ( .A1(n5660), .A2(n5659), .ZN(n9439) );
  NAND2_X1 U5727 ( .A1(n5521), .A2(n5520), .ZN(n8361) );
  AND3_X1 U5728 ( .A1(n5265), .A2(n5264), .A3(n5263), .ZN(n10501) );
  AND3_X1 U5729 ( .A1(n5222), .A2(n5221), .A3(n5220), .ZN(n10494) );
  NOR2_X1 U5730 ( .A1(n10474), .A2(n10466), .ZN(n10471) );
  AND2_X1 U5731 ( .A1(n8902), .A2(n8931), .ZN(n10467) );
  AND2_X1 U5732 ( .A1(n5761), .A2(n5776), .ZN(n10451) );
  NOR2_X1 U5733 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(n5058), .ZN(n5057) );
  NAND2_X1 U5734 ( .A1(n5101), .A2(n5059), .ZN(n5058) );
  AND2_X1 U5735 ( .A1(n4784), .A2(n5059), .ZN(n4783) );
  OR2_X1 U5736 ( .A1(n5123), .A2(n9696), .ZN(n5128) );
  AND2_X1 U5737 ( .A1(n5094), .A2(n5088), .ZN(n4785) );
  XNOR2_X1 U5738 ( .A(n5160), .B(P2_IR_REG_1__SCAN_IN), .ZN(n7704) );
  OR2_X1 U5739 ( .A1(n5906), .A2(n5895), .ZN(n5897) );
  NAND2_X1 U5740 ( .A1(n4988), .A2(n4987), .ZN(n7486) );
  AOI21_X1 U5741 ( .B1(n4990), .B2(n4993), .A(n4536), .ZN(n4987) );
  AND2_X1 U5742 ( .A1(n7350), .A2(n6534), .ZN(n4630) );
  NAND2_X1 U5743 ( .A1(n7043), .A2(n6486), .ZN(n7068) );
  NAND2_X1 U5744 ( .A1(n5015), .A2(n5014), .ZN(n4635) );
  NOR2_X1 U5745 ( .A1(n4521), .A2(n5016), .ZN(n5014) );
  NAND2_X1 U5746 ( .A1(n9740), .A2(n5030), .ZN(n9783) );
  AND2_X1 U5747 ( .A1(n6623), .A2(n6620), .ZN(n5030) );
  NAND2_X1 U5748 ( .A1(n4639), .A2(n4637), .ZN(n9797) );
  OR2_X1 U5749 ( .A1(n4641), .A2(n4638), .ZN(n4637) );
  INV_X1 U5750 ( .A(n4738), .ZN(n4737) );
  OAI21_X1 U5751 ( .B1(n6398), .B2(n6397), .A(n6396), .ZN(n6399) );
  OAI21_X1 U5752 ( .B1(n6400), .B2(n6717), .A(n6404), .ZN(n4738) );
  NOR2_X1 U5753 ( .A1(n6405), .A2(n7100), .ZN(n4736) );
  NAND2_X1 U5754 ( .A1(n6402), .A2(n7367), .ZN(n4734) );
  AND4_X1 U5755 ( .A1(n6042), .A2(n6041), .A3(n6040), .A4(n6039), .ZN(n10339)
         );
  XNOR2_X1 U5756 ( .A(n6890), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n6934) );
  INV_X1 U5757 ( .A(n6849), .ZN(n7057) );
  INV_X1 U5758 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n8817) );
  AND2_X1 U5759 ( .A1(n4892), .A2(n4891), .ZN(n6981) );
  NAND2_X1 U5760 ( .A1(n6850), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4891) );
  NAND2_X1 U5761 ( .A1(n6981), .A2(n6980), .ZN(n6979) );
  AND2_X1 U5762 ( .A1(n7027), .A2(n6851), .ZN(n6855) );
  NAND2_X1 U5763 ( .A1(n4896), .A2(n4895), .ZN(n7429) );
  NAND2_X1 U5764 ( .A1(n7305), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4895) );
  OR2_X1 U5765 ( .A1(n6022), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n6010) );
  NAND2_X1 U5766 ( .A1(n4566), .A2(n4565), .ZN(n4900) );
  INV_X1 U5767 ( .A(n7607), .ZN(n4565) );
  NAND2_X1 U5768 ( .A1(n4902), .A2(n4901), .ZN(n4566) );
  NAND2_X1 U5769 ( .A1(n7606), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4901) );
  XNOR2_X1 U5770 ( .A(n8278), .B(n8284), .ZN(n8016) );
  AND2_X1 U5771 ( .A1(n4569), .A2(n4568), .ZN(n9861) );
  NAND2_X1 U5772 ( .A1(n9858), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4568) );
  NOR2_X1 U5773 ( .A1(n9861), .A2(n9860), .ZN(n9876) );
  NAND2_X1 U5774 ( .A1(n6246), .A2(n6245), .ZN(n9913) );
  OR2_X1 U5775 ( .A1(n8923), .A2(n6177), .ZN(n6246) );
  AND2_X1 U5776 ( .A1(n6380), .A2(n8506), .ZN(n9922) );
  NAND2_X1 U5777 ( .A1(n9923), .A2(n6295), .ZN(n9943) );
  NAND2_X1 U5778 ( .A1(n6268), .A2(n6267), .ZN(n9961) );
  NOR2_X1 U5779 ( .A1(n9984), .A2(n8501), .ZN(n9970) );
  AND4_X1 U5780 ( .A1(n6220), .A2(n6219), .A3(n6218), .A4(n6217), .ZN(n9974)
         );
  NOR2_X1 U5781 ( .A1(n9985), .A2(n9986), .ZN(n9984) );
  NOR2_X1 U5782 ( .A1(n10014), .A2(n10087), .ZN(n10000) );
  NAND2_X1 U5783 ( .A1(n8495), .A2(n8494), .ZN(n10052) );
  NOR2_X1 U5784 ( .A1(n10102), .A2(n4904), .ZN(n4903) );
  INV_X1 U5785 ( .A(n4905), .ZN(n4904) );
  AND2_X1 U5786 ( .A1(n6346), .A2(n8494), .ZN(n8480) );
  NAND2_X1 U5787 ( .A1(n8317), .A2(n9750), .ZN(n8404) );
  NAND2_X1 U5788 ( .A1(n8317), .A2(n4906), .ZN(n8452) );
  INV_X1 U5789 ( .A(n5977), .ZN(n5965) );
  INV_X1 U5790 ( .A(n4760), .ZN(n8313) );
  OR2_X1 U5791 ( .A1(n8151), .A2(n8150), .ZN(n4986) );
  OR2_X1 U5792 ( .A1(n8156), .A2(n10122), .ZN(n8233) );
  AND2_X1 U5793 ( .A1(n8223), .A2(n6332), .ZN(n8150) );
  INV_X1 U5794 ( .A(n4764), .ZN(n8222) );
  OAI21_X1 U5795 ( .B1(n7926), .B2(n4765), .A(n4766), .ZN(n4764) );
  NAND2_X1 U5796 ( .A1(n7921), .A2(n7984), .ZN(n8156) );
  NOR2_X1 U5797 ( .A1(n7820), .A2(n10270), .ZN(n7921) );
  NOR2_X1 U5798 ( .A1(n7765), .A2(n7917), .ZN(n7926) );
  NAND2_X1 U5799 ( .A1(n4910), .A2(n4909), .ZN(n7820) );
  AND4_X1 U5800 ( .A1(n6008), .A2(n6007), .A3(n6006), .A4(n6005), .ZN(n7928)
         );
  INV_X1 U5801 ( .A(n4910), .ZN(n10240) );
  AND2_X1 U5802 ( .A1(n6053), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6038) );
  NAND2_X1 U5803 ( .A1(n7404), .A2(n7403), .ZN(n7758) );
  AND2_X1 U5804 ( .A1(n6091), .A2(n6090), .ZN(n7312) );
  AND4_X1 U5805 ( .A1(n6112), .A2(n6111), .A3(n6110), .A4(n6109), .ZN(n7258)
         );
  AND4_X1 U5806 ( .A1(n6135), .A2(n6134), .A3(n6133), .A4(n6132), .ZN(n7284)
         );
  OR2_X1 U5807 ( .A1(n6177), .A2(n6891), .ZN(n6150) );
  OR2_X1 U5808 ( .A1(n6174), .A2(n6892), .ZN(n6151) );
  NAND2_X1 U5809 ( .A1(n7215), .A2(n7214), .ZN(n7213) );
  AND2_X1 U5810 ( .A1(n4732), .A2(n7205), .ZN(n7214) );
  AND4_X1 U5811 ( .A1(n6168), .A2(n6167), .A3(n6166), .A4(n6165), .ZN(n7285)
         );
  NAND2_X1 U5812 ( .A1(n8256), .A2(n6117), .ZN(n6207) );
  NAND2_X1 U5813 ( .A1(n6213), .A2(n6212), .ZN(n10072) );
  NAND2_X1 U5814 ( .A1(n8177), .A2(n6117), .ZN(n6213) );
  AND2_X1 U5815 ( .A1(n7141), .A2(n6715), .ZN(n10133) );
  NAND2_X1 U5816 ( .A1(n7398), .A2(n7397), .ZN(n10326) );
  INV_X1 U5817 ( .A(n7205), .ZN(n7221) );
  XNOR2_X1 U5818 ( .A(n6254), .B(n6253), .ZN(n9694) );
  XNOR2_X1 U5819 ( .A(n6232), .B(n5821), .ZN(n8472) );
  XNOR2_X1 U5820 ( .A(n5816), .B(n5815), .ZN(n8347) );
  XNOR2_X1 U5821 ( .A(n5736), .B(n5735), .ZN(n8256) );
  XNOR2_X1 U5822 ( .A(n6460), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6697) );
  INV_X1 U5823 ( .A(n5842), .ZN(n4743) );
  INV_X1 U5824 ( .A(n5631), .ZN(n5629) );
  XNOR2_X1 U5825 ( .A(n5598), .B(n5597), .ZN(n7537) );
  NAND2_X1 U5826 ( .A1(n4815), .A2(n5529), .ZN(n5550) );
  NAND2_X1 U5827 ( .A1(n4821), .A2(n4819), .ZN(n4815) );
  NAND2_X1 U5828 ( .A1(n5517), .A2(n5492), .ZN(n4821) );
  XNOR2_X1 U5829 ( .A(n4674), .B(n5528), .ZN(n7162) );
  OAI21_X1 U5830 ( .B1(n5517), .B2(n5516), .A(n5492), .ZN(n4674) );
  NAND2_X1 U5831 ( .A1(n4809), .A2(n5458), .ZN(n5483) );
  OAI21_X1 U5832 ( .B1(n5432), .B2(n5431), .A(n5430), .ZN(n5457) );
  INV_X1 U5833 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U5834 ( .A1(n5375), .A2(n5374), .ZN(n5399) );
  XNOR2_X1 U5835 ( .A(n5373), .B(n5065), .ZN(n6975) );
  OR3_X1 U5836 ( .A1(n6061), .A2(P1_IR_REG_7__SCAN_IN), .A3(
        P1_IR_REG_8__SCAN_IN), .ZN(n6043) );
  NAND2_X1 U5837 ( .A1(n4923), .A2(n5301), .ZN(n5325) );
  XNOR2_X1 U5838 ( .A(n5258), .B(SI_5_), .ZN(n5256) );
  XNOR2_X1 U5839 ( .A(n4887), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6890) );
  NAND2_X1 U5840 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4887) );
  NOR2_X1 U5841 ( .A1(n4506), .A2(n4853), .ZN(n4852) );
  NAND2_X1 U5842 ( .A1(n9191), .A2(n4854), .ZN(n4851) );
  INV_X1 U5843 ( .A(n9137), .ZN(n4853) );
  NAND2_X1 U5844 ( .A1(n8048), .A2(n5476), .ZN(n8920) );
  NAND2_X1 U5845 ( .A1(n5652), .A2(n5651), .ZN(n9159) );
  AND4_X1 U5846 ( .A1(n5342), .A2(n5341), .A3(n5340), .A4(n5339), .ZN(n7808)
         );
  NAND2_X1 U5847 ( .A1(n4840), .A2(n4838), .ZN(n9179) );
  AND2_X1 U5848 ( .A1(n4839), .A2(n5607), .ZN(n4838) );
  NAND2_X1 U5849 ( .A1(n5563), .A2(n4841), .ZN(n4840) );
  INV_X1 U5850 ( .A(n5421), .ZN(n7990) );
  NAND2_X1 U5851 ( .A1(n4621), .A2(n4847), .ZN(n8438) );
  NAND2_X1 U5852 ( .A1(n7782), .A2(n5345), .ZN(n8901) );
  AND4_X1 U5853 ( .A1(n5365), .A2(n5364), .A3(n5363), .A4(n5362), .ZN(n8895)
         );
  NAND2_X1 U5854 ( .A1(n8938), .A2(n4863), .ZN(n7657) );
  INV_X1 U5855 ( .A(n7452), .ZN(n4863) );
  OAI21_X1 U5856 ( .B1(n5563), .B2(n4846), .A(n4843), .ZN(n8462) );
  NOR2_X1 U5857 ( .A1(n9240), .A2(n7521), .ZN(n9235) );
  NAND2_X1 U5858 ( .A1(n5184), .A2(n7586), .ZN(n7596) );
  NAND2_X1 U5859 ( .A1(n5563), .A2(n8336), .ZN(n8338) );
  NAND2_X1 U5860 ( .A1(n7532), .A2(n4525), .ZN(n7558) );
  AND2_X1 U5861 ( .A1(n7532), .A2(n7529), .ZN(n7560) );
  INV_X1 U5862 ( .A(n9239), .ZN(n4624) );
  NAND2_X1 U5863 ( .A1(n9241), .A2(n9242), .ZN(n4623) );
  NAND2_X1 U5864 ( .A1(n4859), .A2(n4860), .ZN(n9241) );
  AND2_X1 U5865 ( .A1(n5721), .A2(n5701), .ZN(n9408) );
  INV_X1 U5866 ( .A(n10593), .ZN(n9252) );
  NAND4_X1 U5867 ( .A1(n5318), .A2(n5317), .A3(n5316), .A4(n5315), .ZN(n9272)
         );
  NAND4_X1 U5868 ( .A1(n5283), .A2(n5282), .A3(n5281), .A4(n5280), .ZN(n9273)
         );
  NAND4_X1 U5869 ( .A1(n5251), .A2(n5250), .A3(n5249), .A4(n5248), .ZN(n9275)
         );
  NAND2_X1 U5870 ( .A1(n5224), .A2(n4692), .ZN(n9276) );
  OR2_X1 U5871 ( .A1(n4498), .A2(n5223), .ZN(n5224) );
  NOR2_X1 U5872 ( .A1(n4524), .A2(n4693), .ZN(n4692) );
  NAND2_X1 U5873 ( .A1(n5225), .A2(n5226), .ZN(n4693) );
  NAND4_X1 U5874 ( .A1(n5194), .A2(n5193), .A3(n5192), .A4(n5191), .ZN(n9277)
         );
  NAND4_X2 U5875 ( .A1(n5183), .A2(n5182), .A3(n5181), .A4(n5180), .ZN(n9278)
         );
  OR2_X1 U5876 ( .A1(n7014), .A2(n7705), .ZN(n5165) );
  NAND4_X1 U5877 ( .A1(n5140), .A2(n5139), .A3(n5138), .A4(n5137), .ZN(n9281)
         );
  OR2_X1 U5878 ( .A1(n7014), .A2(n5136), .ZN(n5137) );
  XNOR2_X1 U5879 ( .A(n4879), .B(n4878), .ZN(n10164) );
  INV_X1 U5880 ( .A(n4871), .ZN(n8180) );
  INV_X1 U5881 ( .A(n4597), .ZN(n8184) );
  NOR2_X1 U5882 ( .A1(n8213), .A2(n8212), .ZN(n8211) );
  AND2_X1 U5883 ( .A1(n4871), .A2(n4870), .ZN(n8213) );
  NAND2_X1 U5884 ( .A1(n7709), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4870) );
  INV_X1 U5885 ( .A(n4595), .ZN(n8206) );
  NAND2_X1 U5886 ( .A1(n4595), .A2(n4594), .ZN(n7710) );
  INV_X1 U5887 ( .A(n8205), .ZN(n4594) );
  INV_X1 U5888 ( .A(n4584), .ZN(n7881) );
  OR2_X1 U5889 ( .A1(n7887), .A2(n7886), .ZN(n7888) );
  NOR2_X1 U5890 ( .A1(n8119), .A2(n8118), .ZN(n8117) );
  AND2_X1 U5891 ( .A1(n7888), .A2(n4876), .ZN(n8119) );
  NAND2_X1 U5892 ( .A1(n7712), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4876) );
  INV_X1 U5893 ( .A(n7859), .ZN(n7870) );
  INV_X1 U5894 ( .A(n7717), .ZN(n7861) );
  AND2_X1 U5895 ( .A1(n7864), .A2(n4875), .ZN(n8107) );
  NAND2_X1 U5896 ( .A1(n7716), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4875) );
  INV_X1 U5897 ( .A(n4874), .ZN(n8105) );
  NOR2_X1 U5898 ( .A1(n8198), .A2(n4869), .ZN(n7696) );
  AND2_X1 U5899 ( .A1(n8203), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4869) );
  NAND2_X1 U5900 ( .A1(n7696), .A2(n7695), .ZN(n7834) );
  INV_X1 U5901 ( .A(n4606), .ZN(n7830) );
  INV_X1 U5902 ( .A(n9317), .ZN(n9315) );
  OR2_X1 U5903 ( .A1(n9305), .A2(n9306), .ZN(n9312) );
  INV_X1 U5904 ( .A(n9339), .ZN(n10441) );
  OAI21_X1 U5905 ( .B1(n9339), .B2(n5141), .A(n9338), .ZN(n4590) );
  NOR2_X1 U5906 ( .A1(n9341), .A2(n10520), .ZN(n9570) );
  OAI21_X1 U5907 ( .B1(n6824), .B2(n9553), .A(n6823), .ZN(n9358) );
  AOI21_X1 U5908 ( .B1(n9363), .B2(n9532), .A(n9362), .ZN(n9578) );
  OAI21_X1 U5909 ( .B1(n9424), .B2(n4929), .A(n4926), .ZN(n9376) );
  NAND2_X1 U5910 ( .A1(n5699), .A2(n5698), .ZN(n9402) );
  NAND2_X1 U5911 ( .A1(n5683), .A2(n5682), .ZN(n9427) );
  NAND2_X1 U5912 ( .A1(n9459), .A2(n8980), .ZN(n9447) );
  NAND2_X1 U5913 ( .A1(n4942), .A2(n4949), .ZN(n9464) );
  OR2_X1 U5914 ( .A1(n9494), .A2(n4951), .ZN(n4942) );
  AND2_X1 U5915 ( .A1(n4953), .A2(n4515), .ZN(n9476) );
  INV_X1 U5916 ( .A(n6777), .ZN(n9626) );
  NAND2_X1 U5917 ( .A1(n4941), .A2(n4939), .ZN(n9548) );
  NAND2_X1 U5918 ( .A1(n8353), .A2(n5055), .ZN(n8418) );
  AND2_X1 U5919 ( .A1(n8263), .A2(n6804), .ZN(n8166) );
  NAND2_X1 U5920 ( .A1(n8258), .A2(n4933), .ZN(n8170) );
  INV_X1 U5921 ( .A(n10501), .ZN(n7581) );
  AND3_X1 U5922 ( .A1(n5204), .A2(n5203), .A3(n5202), .ZN(n10489) );
  OR2_X1 U5923 ( .A1(n10450), .A2(n6827), .ZN(n9537) );
  NAND2_X1 U5924 ( .A1(n6826), .A2(n4918), .ZN(n6838) );
  AND2_X1 U5925 ( .A1(n6825), .A2(n10541), .ZN(n4918) );
  INV_X1 U5926 ( .A(n9340), .ZN(n9644) );
  INV_X1 U5927 ( .A(n9372), .ZN(n9652) );
  AOI211_X1 U5928 ( .C1(n9591), .C2(n10524), .A(n9590), .B(n9589), .ZN(n9657)
         );
  INV_X1 U5929 ( .A(n9427), .ZN(n9664) );
  INV_X1 U5930 ( .A(n9159), .ZN(n9672) );
  AND2_X1 U5931 ( .A1(n5554), .A2(n5553), .ZN(n9689) );
  INV_X1 U5932 ( .A(n7524), .ZN(n7539) );
  NAND2_X1 U5933 ( .A1(n10528), .A2(n10475), .ZN(n9692) );
  AND2_X1 U5934 ( .A1(n7008), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10465) );
  INV_X1 U5935 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5107) );
  NOR2_X1 U5936 ( .A1(n5199), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9698) );
  NAND2_X1 U5937 ( .A1(n5199), .A2(SI_0_), .ZN(n5143) );
  AND4_X1 U5938 ( .A1(n6073), .A2(n6072), .A3(n6071), .A4(n6070), .ZN(n10341)
         );
  NAND2_X1 U5939 ( .A1(n7348), .A2(n7349), .ZN(n4989) );
  AND4_X1 U5940 ( .A1(n5982), .A2(n5981), .A3(n5980), .A4(n5979), .ZN(n8226)
         );
  AOI21_X1 U5941 ( .B1(n6665), .B2(n9774), .A(n6664), .ZN(n9702) );
  NAND2_X1 U5942 ( .A1(n7546), .A2(n6562), .ZN(n7637) );
  NOR2_X1 U5943 ( .A1(n9797), .A2(n5027), .ZN(n6741) );
  NAND2_X1 U5944 ( .A1(n9724), .A2(n9725), .ZN(n9723) );
  NAND2_X1 U5945 ( .A1(n9765), .A2(n6643), .ZN(n9724) );
  NAND2_X1 U5946 ( .A1(n4643), .A2(n5006), .ZN(n9734) );
  NAND2_X1 U5947 ( .A1(n4635), .A2(n6603), .ZN(n8327) );
  AND4_X1 U5948 ( .A1(n5944), .A2(n5943), .A3(n5942), .A4(n5941), .ZN(n9745)
         );
  OAI21_X1 U5949 ( .B1(n9754), .B2(n9753), .A(n9752), .ZN(n9751) );
  AND4_X1 U5950 ( .A1(n6124), .A2(n6123), .A3(n6122), .A4(n6121), .ZN(n7155)
         );
  NAND2_X1 U5951 ( .A1(n4998), .A2(n6561), .ZN(n7546) );
  INV_X1 U5952 ( .A(n7543), .ZN(n4998) );
  AOI21_X1 U5953 ( .B1(n4519), .B2(n4629), .A(n4626), .ZN(n4625) );
  INV_X1 U5954 ( .A(n7792), .ZN(n4626) );
  AND4_X1 U5955 ( .A1(n6021), .A2(n6020), .A3(n6019), .A4(n6018), .ZN(n10248)
         );
  NAND2_X1 U5956 ( .A1(n7665), .A2(n6574), .ZN(n7666) );
  OAI211_X1 U5957 ( .C1(n6910), .C2(n6177), .A(n6176), .B(n6175), .ZN(n8879)
         );
  OR2_X1 U5958 ( .A1(n4502), .A2(n6893), .ZN(n6175) );
  NAND2_X1 U5959 ( .A1(n5937), .A2(n5936), .ZN(n10112) );
  AND4_X1 U5960 ( .A1(n6203), .A2(n6202), .A3(n6201), .A4(n6200), .ZN(n9990)
         );
  AND2_X1 U5961 ( .A1(n5015), .A2(n5013), .ZN(n8072) );
  INV_X1 U5962 ( .A(n5016), .ZN(n5013) );
  INV_X1 U5963 ( .A(n7284), .ZN(n9829) );
  INV_X1 U5964 ( .A(n4889), .ZN(n6946) );
  NAND2_X1 U5965 ( .A1(n6915), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4888) );
  INV_X1 U5966 ( .A(n4894), .ZN(n10314) );
  INV_X1 U5967 ( .A(n4892), .ZN(n6961) );
  INV_X1 U5968 ( .A(n4574), .ZN(n7196) );
  INV_X1 U5969 ( .A(n4896), .ZN(n7304) );
  INV_X1 U5970 ( .A(n4902), .ZN(n7605) );
  INV_X1 U5971 ( .A(n4900), .ZN(n8014) );
  INV_X1 U5972 ( .A(n4566), .ZN(n7608) );
  NOR2_X1 U5973 ( .A1(n9834), .A2(n9835), .ZN(n9837) );
  INV_X1 U5974 ( .A(n4569), .ZN(n9857) );
  AND2_X1 U5975 ( .A1(n5874), .A2(n5873), .ZN(n9929) );
  INV_X1 U5976 ( .A(n10079), .ZN(n9980) );
  NAND2_X1 U5977 ( .A1(n4659), .A2(n4971), .ZN(n9969) );
  NAND2_X1 U5978 ( .A1(n8485), .A2(n4974), .ZN(n4659) );
  AOI21_X1 U5979 ( .B1(n8485), .B2(n4977), .A(n4976), .ZN(n9983) );
  NAND2_X1 U5980 ( .A1(n4748), .A2(n4752), .ZN(n10006) );
  NAND2_X1 U5981 ( .A1(n8485), .A2(n5062), .ZN(n9999) );
  NAND2_X1 U5982 ( .A1(n10033), .A2(n8497), .ZN(n10020) );
  INV_X1 U5983 ( .A(n4578), .ZN(n8456) );
  NAND2_X1 U5984 ( .A1(n4651), .A2(n4653), .ZN(n8451) );
  NAND2_X1 U5985 ( .A1(n8310), .A2(n4654), .ZN(n4651) );
  NOR2_X1 U5986 ( .A1(n8310), .A2(n4984), .ZN(n8402) );
  NAND2_X1 U5987 ( .A1(n4956), .A2(n7755), .ZN(n7816) );
  NAND2_X1 U5988 ( .A1(n7754), .A2(n4960), .ZN(n4956) );
  AND2_X1 U5989 ( .A1(n7238), .A2(n7237), .ZN(n7241) );
  INV_X2 U5990 ( .A(n10436), .ZN(n10438) );
  NAND2_X1 U5991 ( .A1(n8863), .A2(n10401), .ZN(n4582) );
  NAND2_X1 U5992 ( .A1(n4769), .A2(n4768), .ZN(n4767) );
  NOR2_X1 U5993 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n5012) );
  NAND2_X1 U5994 ( .A1(n6464), .A2(n6452), .ZN(n6465) );
  INV_X1 U5995 ( .A(n6470), .ZN(n7803) );
  INV_X1 U5996 ( .A(n7140), .ZN(n7557) );
  INV_X1 U5997 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6921) );
  OAI21_X1 U5998 ( .B1(n5199), .B2(n6157), .A(n6156), .ZN(n6159) );
  NOR2_X1 U5999 ( .A1(n9128), .A2(n9127), .ZN(n9135) );
  INV_X1 U6000 ( .A(n4604), .ZN(n8085) );
  INV_X1 U6001 ( .A(n4608), .ZN(n9295) );
  INV_X1 U6002 ( .A(n4590), .ZN(n4589) );
  NAND2_X1 U6003 ( .A1(n4586), .A2(n9522), .ZN(n4585) );
  NAND2_X1 U6004 ( .A1(n4592), .A2(n9565), .ZN(n4591) );
  NOR2_X1 U6005 ( .A1(n5020), .A2(n4552), .ZN(n5019) );
  NAND2_X1 U6006 ( .A1(n5023), .A2(n5024), .ZN(n5022) );
  INV_X1 U6007 ( .A(n9905), .ZN(n4880) );
  NAND2_X1 U6008 ( .A1(n4882), .A2(n9902), .ZN(n4881) );
  INV_X1 U6009 ( .A(n4885), .ZN(n4884) );
  AND2_X2 U6010 ( .A1(n5156), .A2(n7389), .ZN(n5576) );
  NAND2_X2 U6011 ( .A1(n6478), .A2(n7131), .ZN(n6487) );
  NOR3_X1 U6012 ( .A1(n5733), .A2(n4855), .A3(n4857), .ZN(n4506) );
  AND2_X1 U6013 ( .A1(n4940), .A2(n8341), .ZN(n4507) );
  AOI21_X1 U6014 ( .B1(n5587), .B2(n4845), .A(n4844), .ZN(n4843) );
  INV_X2 U6015 ( .A(n5894), .ZN(n6004) );
  INV_X1 U6016 ( .A(n6173), .ZN(n6844) );
  INV_X1 U6017 ( .A(n9055), .ZN(n4935) );
  NAND2_X1 U6018 ( .A1(n5833), .A2(n5832), .ZN(n5931) );
  NAND2_X1 U6019 ( .A1(n4634), .A2(n4542), .ZN(n4508) );
  XOR2_X1 U6020 ( .A(n9159), .B(n5661), .Z(n4509) );
  NAND2_X1 U6021 ( .A1(n5947), .A2(n5946), .ZN(n10119) );
  AND2_X1 U6022 ( .A1(n6825), .A2(n10528), .ZN(n4510) );
  AND2_X1 U6023 ( .A1(n9898), .A2(n10319), .ZN(n4511) );
  OR2_X1 U6024 ( .A1(n9501), .A2(n4788), .ZN(n4512) );
  NAND2_X1 U6025 ( .A1(n5466), .A2(n5465), .ZN(n8917) );
  INV_X1 U6026 ( .A(n4857), .ZN(n4856) );
  NOR2_X1 U6027 ( .A1(n9242), .A2(n4858), .ZN(n4857) );
  NOR2_X1 U6028 ( .A1(n4856), .A2(n4861), .ZN(n4855) );
  AOI21_X1 U6029 ( .B1(n4654), .B2(n4984), .A(n4550), .ZN(n4653) );
  INV_X1 U6030 ( .A(n4792), .ZN(n4791) );
  NAND2_X1 U6031 ( .A1(n4794), .A2(n4793), .ZN(n4792) );
  INV_X1 U6032 ( .A(n5026), .ZN(n5025) );
  OAI21_X1 U6033 ( .B1(n5073), .B2(n6690), .A(n6689), .ZN(n5026) );
  OR2_X1 U6034 ( .A1(n9680), .A2(n6809), .ZN(n4513) );
  INV_X1 U6035 ( .A(n9170), .ZN(n4844) );
  NOR2_X1 U6036 ( .A1(n9236), .A2(n4553), .ZN(n9229) );
  AND4_X1 U6037 ( .A1(n5540), .A2(n5539), .A3(n5538), .A4(n5537), .ZN(n8341)
         );
  NAND2_X1 U6038 ( .A1(n6279), .A2(n7924), .ZN(n7917) );
  INV_X1 U6039 ( .A(n7917), .ZN(n4763) );
  INV_X1 U6040 ( .A(n5815), .ZN(n4806) );
  AND2_X2 U6041 ( .A1(n7723), .A2(n6889), .ZN(n5240) );
  OR2_X1 U6042 ( .A1(n7744), .A2(n10505), .ZN(n4514) );
  NAND2_X1 U6043 ( .A1(n6160), .A2(n5199), .ZN(n6174) );
  AND3_X1 U6044 ( .A1(n6151), .A2(n6150), .A3(n6149), .ZN(n7222) );
  NAND2_X1 U6045 ( .A1(n9503), .A2(n9261), .ZN(n4515) );
  INV_X1 U6046 ( .A(n5073), .ZN(n4638) );
  NAND2_X1 U6047 ( .A1(n5290), .A2(n5088), .ZN(n5306) );
  NAND2_X1 U6048 ( .A1(n6160), .A2(n6889), .ZN(n6177) );
  NAND2_X1 U6049 ( .A1(n6697), .A2(n6468), .ZN(n6478) );
  AND2_X2 U6050 ( .A1(n5865), .A2(n5854), .ZN(n6143) );
  OR2_X1 U6051 ( .A1(n9372), .A2(n9145), .ZN(n9106) );
  AND2_X1 U6052 ( .A1(n5522), .A2(n4849), .ZN(n4517) );
  NAND2_X1 U6053 ( .A1(n9159), .A2(n9091), .ZN(n4518) );
  INV_X1 U6054 ( .A(n9080), .ZN(n5051) );
  AND2_X1 U6055 ( .A1(n4628), .A2(n7791), .ZN(n4519) );
  XNOR2_X1 U6056 ( .A(n9393), .B(n9243), .ZN(n9382) );
  INV_X1 U6057 ( .A(n7318), .ZN(n4757) );
  AND2_X1 U6058 ( .A1(n4889), .A2(n4888), .ZN(n4520) );
  AND3_X1 U6059 ( .A1(n5163), .A2(n5162), .A3(n5161), .ZN(n7457) );
  INV_X1 U6060 ( .A(n7457), .ZN(n10474) );
  INV_X1 U6061 ( .A(n8492), .ZN(n8507) );
  AND2_X1 U6062 ( .A1(n6390), .A2(n6443), .ZN(n8492) );
  NAND2_X1 U6063 ( .A1(n5442), .A2(n5441), .ZN(n10220) );
  INV_X1 U6064 ( .A(n10220), .ZN(n4780) );
  AND2_X1 U6065 ( .A1(n8070), .A2(n6601), .ZN(n4521) );
  AND3_X1 U6066 ( .A1(n9108), .A2(n8965), .A3(n9099), .ZN(n4522) );
  INV_X1 U6067 ( .A(n8455), .ZN(n4577) );
  NAND2_X1 U6068 ( .A1(n4744), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6459) );
  AND2_X1 U6069 ( .A1(n5073), .A2(n5008), .ZN(n4523) );
  NAND2_X1 U6070 ( .A1(n5052), .A2(n9080), .ZN(n9496) );
  XNOR2_X1 U6071 ( .A(n8493), .B(n8492), .ZN(n8863) );
  AND2_X1 U6072 ( .A1(n6820), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4524) );
  INV_X1 U6073 ( .A(n4564), .ZN(n9955) );
  NAND2_X1 U6074 ( .A1(n7957), .A2(n7992), .ZN(n9039) );
  INV_X1 U6075 ( .A(n9039), .ZN(n5045) );
  NAND2_X1 U6076 ( .A1(n5031), .A2(n5176), .ZN(n5216) );
  NAND2_X1 U6077 ( .A1(n5912), .A2(n5911), .ZN(n10102) );
  INV_X1 U6078 ( .A(n8401), .ZN(n4654) );
  AND2_X1 U6079 ( .A1(n5880), .A2(n5879), .ZN(n9996) );
  INV_X1 U6080 ( .A(n9996), .ZN(n10084) );
  AND2_X1 U6081 ( .A1(n7529), .A2(n7559), .ZN(n4525) );
  INV_X1 U6082 ( .A(n9468), .ZN(n9676) );
  NAND2_X1 U6083 ( .A1(n5639), .A2(n5638), .ZN(n9468) );
  NOR2_X1 U6084 ( .A1(n7401), .A2(n4757), .ZN(n4526) );
  INV_X1 U6085 ( .A(n9393), .ZN(n9656) );
  NAND2_X1 U6086 ( .A1(n5718), .A2(n5717), .ZN(n9393) );
  INV_X1 U6087 ( .A(n4912), .ZN(n9975) );
  NOR2_X1 U6088 ( .A1(n10014), .A2(n4914), .ZN(n4912) );
  AND2_X1 U6089 ( .A1(n5207), .A2(n5188), .ZN(n4527) );
  AND2_X1 U6090 ( .A1(n10132), .A2(n9821), .ZN(n4528) );
  NAND3_X1 U6091 ( .A1(n4610), .A2(n4878), .A3(n4609), .ZN(n4529) );
  AND2_X1 U6092 ( .A1(n7240), .A2(n7237), .ZN(n4530) );
  INV_X1 U6093 ( .A(n8497), .ZN(n4755) );
  INV_X1 U6094 ( .A(n4950), .ZN(n4949) );
  NAND2_X1 U6095 ( .A1(n4531), .A2(n4513), .ZN(n4950) );
  NAND2_X1 U6096 ( .A1(n9648), .A2(n9253), .ZN(n9116) );
  INV_X1 U6097 ( .A(n9116), .ZN(n8970) );
  OR2_X1 U6098 ( .A1(n6779), .A2(n4515), .ZN(n4531) );
  INV_X1 U6099 ( .A(n4934), .ZN(n4933) );
  NOR2_X1 U6100 ( .A1(n4780), .A2(n9049), .ZN(n4934) );
  AND4_X1 U6101 ( .A1(n5099), .A2(n5098), .A3(n5097), .A4(n5096), .ZN(n4532)
         );
  AND2_X1 U6102 ( .A1(n4652), .A2(n8450), .ZN(n4533) );
  NOR2_X1 U6103 ( .A1(n8917), .A2(n9267), .ZN(n4534) );
  AND2_X1 U6104 ( .A1(n9980), .A2(n9990), .ZN(n4535) );
  INV_X1 U6105 ( .A(n4779), .ZN(n4778) );
  NAND2_X1 U6106 ( .A1(n4780), .A2(n4781), .ZN(n4779) );
  NAND2_X1 U6107 ( .A1(n6547), .A2(n6546), .ZN(n4536) );
  INV_X1 U6108 ( .A(n8930), .ZN(n9648) );
  NAND2_X1 U6109 ( .A1(n8925), .A2(n8924), .ZN(n8930) );
  AND2_X1 U6110 ( .A1(n9478), .A2(n9085), .ZN(n9495) );
  NAND2_X1 U6111 ( .A1(n5871), .A2(n5870), .ZN(n10065) );
  AND2_X1 U6112 ( .A1(n9066), .A2(n9065), .ZN(n4537) );
  NAND2_X1 U6113 ( .A1(n5052), .A2(n5050), .ZN(n9477) );
  INV_X1 U6114 ( .A(n4980), .ZN(n4976) );
  NAND2_X1 U6115 ( .A1(n10003), .A2(n9989), .ZN(n4980) );
  NAND2_X1 U6116 ( .A1(n9108), .A2(n9106), .ZN(n4538) );
  AND2_X1 U6117 ( .A1(n4785), .A2(n4865), .ZN(n4539) );
  NAND2_X1 U6118 ( .A1(n5926), .A2(n5925), .ZN(n10108) );
  NAND2_X1 U6119 ( .A1(n9066), .A2(n9265), .ZN(n4540) );
  AND2_X1 U6120 ( .A1(n6810), .A2(n9515), .ZN(n4541) );
  AND2_X1 U6121 ( .A1(n4990), .A2(n4536), .ZN(n4542) );
  INV_X1 U6122 ( .A(n7350), .ZN(n4993) );
  OR2_X1 U6123 ( .A1(n9030), .A2(n9029), .ZN(n4543) );
  INV_X1 U6124 ( .A(n6562), .ZN(n4997) );
  AND2_X1 U6125 ( .A1(n5758), .A2(n4783), .ZN(n5150) );
  AND2_X1 U6126 ( .A1(n6611), .A2(n6603), .ZN(n4544) );
  AND2_X1 U6127 ( .A1(n6311), .A2(n7757), .ZN(n4545) );
  AND2_X1 U6128 ( .A1(n6811), .A2(n4518), .ZN(n4546) );
  AND2_X1 U6129 ( .A1(n4675), .A2(n4916), .ZN(n4547) );
  OR2_X1 U6130 ( .A1(n5025), .A2(n4638), .ZN(n4548) );
  INV_X1 U6131 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5059) );
  INV_X1 U6132 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4878) );
  NAND2_X1 U6133 ( .A1(n5347), .A2(n5305), .ZN(n5326) );
  CLKBUF_X3 U6134 ( .A(n6162), .Z(n6095) );
  NAND2_X1 U6135 ( .A1(n6788), .A2(n6787), .ZN(n6834) );
  INV_X1 U6136 ( .A(n6834), .ZN(n4793) );
  OR2_X1 U6137 ( .A1(n6773), .A2(n6774), .ZN(n4936) );
  INV_X1 U6138 ( .A(n9926), .ZN(n9964) );
  AND4_X1 U6139 ( .A1(n6211), .A2(n6210), .A3(n6209), .A4(n6208), .ZN(n9926)
         );
  INV_X1 U6140 ( .A(n4826), .ZN(n4825) );
  NAND2_X1 U6141 ( .A1(n4829), .A2(n4827), .ZN(n4826) );
  NAND2_X1 U6142 ( .A1(n6207), .A2(n6206), .ZN(n10067) );
  INV_X1 U6143 ( .A(n10067), .ZN(n4563) );
  NAND2_X1 U6144 ( .A1(n7666), .A2(n6578), .ZN(n7793) );
  NAND2_X1 U6145 ( .A1(n4627), .A2(n4625), .ZN(n7846) );
  AND3_X1 U6146 ( .A1(n6745), .A2(n9802), .A3(n6744), .ZN(n4549) );
  AND2_X1 U6147 ( .A1(n10119), .A2(n9816), .ZN(n4550) );
  OR2_X1 U6148 ( .A1(n4936), .A2(n4935), .ZN(n8258) );
  INV_X1 U6149 ( .A(n6690), .ZN(n5028) );
  AND2_X1 U6150 ( .A1(n10065), .A2(n10133), .ZN(n4551) );
  INV_X1 U6151 ( .A(n5102), .ZN(n5756) );
  NOR2_X1 U6152 ( .A1(n4563), .A2(n9812), .ZN(n4552) );
  NAND2_X1 U6153 ( .A1(n8317), .A2(n4905), .ZN(n4907) );
  AND2_X1 U6154 ( .A1(n9259), .A2(n8938), .ZN(n4553) );
  OR2_X1 U6155 ( .A1(n7893), .A2(n7713), .ZN(n4554) );
  AND2_X1 U6156 ( .A1(n5046), .A2(n9039), .ZN(n4555) );
  OR2_X1 U6157 ( .A1(n7428), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4556) );
  NAND2_X1 U6158 ( .A1(n4539), .A2(n5290), .ZN(n4557) );
  INV_X1 U6159 ( .A(n5655), .ZN(n5656) );
  AND2_X1 U6160 ( .A1(n4941), .A2(n4540), .ZN(n4558) );
  AND2_X1 U6161 ( .A1(n4986), .A2(n4985), .ZN(n4559) );
  AND3_X1 U6162 ( .A1(n5784), .A2(n5783), .A3(n10518), .ZN(n9212) );
  NAND2_X1 U6163 ( .A1(n5534), .A2(n5533), .ZN(n9559) );
  INV_X1 U6164 ( .A(n9559), .ZN(n4940) );
  NAND2_X1 U6165 ( .A1(n5963), .A2(n5962), .ZN(n8332) );
  INV_X1 U6166 ( .A(n8332), .ZN(n4672) );
  NAND2_X1 U6167 ( .A1(n8036), .A2(n7945), .ZN(n7914) );
  INV_X1 U6168 ( .A(n8336), .ZN(n4845) );
  NAND2_X1 U6169 ( .A1(n7596), .A2(n4527), .ZN(n7415) );
  AND2_X1 U6170 ( .A1(n7148), .A2(n6519), .ZN(n4560) );
  NAND2_X1 U6171 ( .A1(n6013), .A2(n6012), .ZN(n10132) );
  INV_X1 U6172 ( .A(n10132), .ZN(n4909) );
  AOI21_X1 U6173 ( .B1(n7438), .B2(n6763), .A(n5060), .ZN(n7570) );
  NAND2_X1 U6174 ( .A1(n4970), .A2(n7315), .ZN(n7398) );
  NAND2_X1 U6175 ( .A1(n8036), .A2(n4778), .ZN(n4782) );
  AND2_X1 U6176 ( .A1(n4989), .A2(n7350), .ZN(n4561) );
  INV_X1 U6177 ( .A(n4805), .ZN(n4804) );
  OAI21_X1 U6178 ( .B1(n4806), .B2(n5737), .A(n5820), .ZN(n4805) );
  NAND2_X1 U6179 ( .A1(n5847), .A2(n5850), .ZN(n6458) );
  NAND4_X1 U6180 ( .A1(n6155), .A2(n6154), .A3(n6153), .A4(n6152), .ZN(n9831)
         );
  INV_X1 U6181 ( .A(n9831), .ZN(n4732) );
  NAND2_X1 U6182 ( .A1(n7371), .A2(n7372), .ZN(n7370) );
  AND2_X1 U6183 ( .A1(n6722), .A2(n6716), .ZN(n9802) );
  INV_X1 U6184 ( .A(n8877), .ZN(n7099) );
  INV_X1 U6185 ( .A(n7349), .ZN(n4992) );
  NAND2_X1 U6186 ( .A1(n7210), .A2(n7211), .ZN(n7209) );
  AND2_X1 U6187 ( .A1(n9316), .A2(n9297), .ZN(n4562) );
  INV_X1 U6188 ( .A(n5153), .ZN(n9565) );
  XNOR2_X1 U6189 ( .A(n5126), .B(n5125), .ZN(n8942) );
  NAND2_X1 U6190 ( .A1(n5103), .A2(n5104), .ZN(n9695) );
  NAND2_X1 U6191 ( .A1(n6470), .A2(n7095), .ZN(n7100) );
  INV_X1 U6192 ( .A(n9111), .ZN(n4706) );
  AOI21_X1 U6193 ( .B1(n9335), .B2(n10440), .A(n10165), .ZN(n4593) );
  NAND2_X1 U6194 ( .A1(n9337), .A2(n10440), .ZN(n4587) );
  INV_X1 U6195 ( .A(P2_U3966), .ZN(n9280) );
  OAI222_X1 U6196 ( .A1(n8906), .A2(n8479), .B1(P2_U3152), .B2(n8478), .C1(
        n8904), .C2(n8923), .ZN(P2_U3328) );
  INV_X2 U6197 ( .A(n9698), .ZN(n8906) );
  OAI21_X1 U6198 ( .B1(n4677), .B2(n9081), .A(n9119), .ZN(n4676) );
  OAI21_X1 U6199 ( .B1(n9015), .B2(n9119), .A(n4689), .ZN(n4688) );
  NOR2_X1 U6200 ( .A1(n9017), .A2(n9119), .ZN(n4687) );
  NOR2_X2 U6201 ( .A1(n7327), .A2(n10404), .ZN(n10327) );
  NAND2_X1 U6202 ( .A1(n8869), .A2(n10265), .ZN(n4675) );
  XNOR2_X1 U6203 ( .A(n4581), .B(n8862), .ZN(P1_U3552) );
  NAND2_X1 U6204 ( .A1(n4575), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4647) );
  AOI21_X2 U6205 ( .B1(n4497), .B2(n10438), .A(n8516), .ZN(n4581) );
  INV_X2 U6206 ( .A(n5175), .ZN(n5199) );
  MUX2_X1 U6207 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5175), .Z(n5198) );
  AND2_X2 U6208 ( .A1(n4646), .A2(n4645), .ZN(n5175) );
  AOI21_X2 U6209 ( .B1(n9960), .B2(n8504), .A(n8503), .ZN(n9942) );
  NAND3_X1 U6210 ( .A1(n4591), .A2(n4589), .A3(n4585), .ZN(P2_U3264) );
  INV_X1 U6211 ( .A(n9229), .ZN(n4612) );
  OAI21_X1 U6212 ( .B1(n9229), .B2(n5642), .A(n4509), .ZN(n4613) );
  NAND2_X1 U6213 ( .A1(n9149), .A2(n9152), .ZN(n4614) );
  INV_X1 U6214 ( .A(n4613), .ZN(n9151) );
  MUX2_X1 U6215 ( .A(n8884), .B(n8479), .S(n5199), .Z(n6237) );
  MUX2_X1 U6216 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n5199), .Z(n6252) );
  NAND2_X2 U6217 ( .A1(P1_U3084), .A2(n5199), .ZN(n8885) );
  NAND2_X2 U6218 ( .A1(P2_U3152), .A2(n5199), .ZN(n8904) );
  NAND2_X1 U6219 ( .A1(n7038), .A2(n4504), .ZN(n4619) );
  NAND2_X1 U6220 ( .A1(n4621), .A2(n4620), .ZN(n8435) );
  NAND3_X1 U6221 ( .A1(n4624), .A2(n4623), .A3(n9212), .ZN(n9251) );
  NAND2_X1 U6222 ( .A1(n7665), .A2(n4519), .ZN(n4627) );
  NAND2_X1 U6223 ( .A1(n4631), .A2(n6534), .ZN(n7348) );
  NAND2_X1 U6224 ( .A1(n4631), .A2(n4630), .ZN(n4634) );
  NAND2_X1 U6225 ( .A1(n4635), .A2(n4544), .ZN(n8324) );
  NAND3_X1 U6226 ( .A1(n9774), .A2(n6665), .A3(n6664), .ZN(n4644) );
  NAND3_X1 U6227 ( .A1(n5010), .A2(n4644), .A3(n4523), .ZN(n4639) );
  NAND2_X1 U6228 ( .A1(n4640), .A2(n4644), .ZN(n4643) );
  AND3_X2 U6229 ( .A1(n4774), .A2(n4773), .A3(n5833), .ZN(n5921) );
  INV_X2 U6230 ( .A(n6137), .ZN(n5833) );
  NAND2_X1 U6231 ( .A1(n5286), .A2(n5285), .ZN(n5289) );
  NAND2_X1 U6232 ( .A1(n5257), .A2(n5256), .ZN(n4648) );
  OAI22_X2 U6233 ( .A1(n8481), .A2(n8480), .B1(n9789), .B2(n9722), .ZN(n10044)
         );
  NAND2_X1 U6234 ( .A1(n4656), .A2(SI_1_), .ZN(n5174) );
  NAND2_X1 U6235 ( .A1(n5159), .A2(n6158), .ZN(n4656) );
  NAND2_X1 U6236 ( .A1(n8485), .A2(n4660), .ZN(n4657) );
  NAND2_X1 U6237 ( .A1(n4657), .A2(n4658), .ZN(n9953) );
  NAND2_X1 U6238 ( .A1(n5375), .A2(n4667), .ZN(n4666) );
  NAND2_X2 U6239 ( .A1(n5799), .A2(n9129), .ZN(n7723) );
  AND2_X1 U6240 ( .A1(n9038), .A2(n4543), .ZN(n4681) );
  OAI21_X1 U6241 ( .B1(n6339), .B2(n4719), .A(n4717), .ZN(n4716) );
  INV_X1 U6242 ( .A(n6339), .ZN(n6340) );
  NAND3_X1 U6243 ( .A1(n4731), .A2(n4545), .A3(n4729), .ZN(n4728) );
  NAND3_X1 U6244 ( .A1(n6308), .A2(n7403), .A3(n4730), .ZN(n4729) );
  NAND2_X1 U6245 ( .A1(n6161), .A2(n7213), .ZN(n4756) );
  XNOR2_X2 U6246 ( .A(n7222), .B(n4733), .ZN(n7215) );
  NAND2_X1 U6247 ( .A1(n6292), .A2(n9902), .ZN(n4735) );
  OAI211_X1 U6248 ( .C1(n7232), .C2(n6717), .A(n4739), .B(n7239), .ZN(n6306)
         );
  NAND2_X1 U6249 ( .A1(n4740), .A2(n6717), .ZN(n4739) );
  NAND4_X1 U6250 ( .A1(n4962), .A2(n4774), .A3(n4773), .A4(n4742), .ZN(n4744)
         );
  NAND2_X1 U6251 ( .A1(n5921), .A2(n4962), .ZN(n6463) );
  NAND3_X1 U6252 ( .A1(n4746), .A2(n6373), .A3(n6358), .ZN(n4745) );
  NAND2_X1 U6253 ( .A1(n4756), .A2(n7094), .ZN(n6178) );
  OAI21_X1 U6254 ( .B1(n4756), .B2(n6416), .A(n6415), .ZN(n6418) );
  XNOR2_X1 U6255 ( .A(n4756), .B(n7094), .ZN(n7098) );
  NAND2_X1 U6256 ( .A1(n7319), .A2(n7318), .ZN(n4758) );
  XNOR2_X1 U6257 ( .A(n4758), .B(n7320), .ZN(n7324) );
  NAND2_X1 U6258 ( .A1(n7758), .A2(n7757), .ZN(n10243) );
  NOR2_X1 U6259 ( .A1(n7926), .A2(n7925), .ZN(n8145) );
  INV_X1 U6260 ( .A(n4782), .ZN(n8271) );
  NAND2_X1 U6261 ( .A1(n5758), .A2(n4784), .ZN(n5148) );
  NAND2_X1 U6262 ( .A1(n5290), .A2(n4785), .ZN(n5497) );
  INV_X1 U6263 ( .A(n4786), .ZN(n9438) );
  AND2_X1 U6264 ( .A1(n9407), .A2(n4791), .ZN(n9347) );
  NAND2_X1 U6265 ( .A1(n9407), .A2(n4790), .ZN(n9346) );
  NAND2_X1 U6266 ( .A1(n9407), .A2(n4794), .ZN(n9369) );
  OAI21_X1 U6267 ( .B1(n5738), .B2(n4806), .A(n4804), .ZN(n6232) );
  INV_X1 U6268 ( .A(n4802), .ZN(n6231) );
  NAND2_X1 U6269 ( .A1(n5738), .A2(n5737), .ZN(n5816) );
  NAND2_X1 U6270 ( .A1(n5517), .A2(n4813), .ZN(n4812) );
  NAND2_X1 U6271 ( .A1(n4812), .A2(n4816), .ZN(n5566) );
  AOI21_X1 U6272 ( .B1(n5658), .B2(n5657), .A(n5656), .ZN(n5674) );
  NAND2_X1 U6273 ( .A1(n5711), .A2(n5710), .ZN(n5736) );
  NAND2_X1 U6274 ( .A1(n6235), .A2(n6234), .ZN(n6239) );
  NAND2_X1 U6275 ( .A1(n5289), .A2(n5288), .ZN(n5299) );
  NAND2_X1 U6276 ( .A1(n5634), .A2(n5633), .ZN(n5644) );
  NAND2_X1 U6277 ( .A1(n5736), .A2(n5735), .ZN(n5738) );
  NAND2_X1 U6278 ( .A1(n5709), .A2(n5708), .ZN(n5711) );
  AND2_X1 U6279 ( .A1(n5040), .A2(n5037), .ZN(n8934) );
  OAI21_X1 U6280 ( .B1(n9361), .B2(n5034), .A(n5033), .ZN(n5039) );
  INV_X1 U6281 ( .A(n6263), .ZN(n9906) );
  NAND2_X1 U6282 ( .A1(n5569), .A2(n5568), .ZN(n5591) );
  NAND2_X1 U6283 ( .A1(n5566), .A2(n5565), .ZN(n5569) );
  NAND2_X1 U6284 ( .A1(n4833), .A2(n5814), .ZN(P2_U3222) );
  OAI211_X1 U6285 ( .C1(n5790), .C2(n5782), .A(n4834), .B(n5791), .ZN(n4833)
         );
  NAND2_X1 U6286 ( .A1(n5790), .A2(n5789), .ZN(n4834) );
  NAND3_X1 U6287 ( .A1(n5176), .A2(n5031), .A3(n5086), .ZN(n5218) );
  INV_X1 U6288 ( .A(n8463), .ZN(n4842) );
  NAND3_X1 U6289 ( .A1(n4842), .A2(n4843), .A3(n4846), .ZN(n4839) );
  NAND2_X1 U6290 ( .A1(n4851), .A2(n4852), .ZN(n9141) );
  NAND2_X1 U6291 ( .A1(n9191), .A2(n4861), .ZN(n4859) );
  INV_X1 U6292 ( .A(n9188), .ZN(n4862) );
  NAND2_X1 U6293 ( .A1(n4539), .A2(n4864), .ZN(n5551) );
  OR2_X2 U6294 ( .A1(n8182), .A2(n8181), .ZN(n4871) );
  NOR2_X1 U6295 ( .A1(n5176), .A2(n9696), .ZN(n4879) );
  NAND3_X1 U6296 ( .A1(n4884), .A2(n4881), .A3(n4880), .ZN(P1_U3260) );
  AND2_X2 U6297 ( .A1(n8317), .A2(n4903), .ZN(n10046) );
  INV_X1 U6298 ( .A(n4907), .ZN(n10045) );
  AND2_X1 U6299 ( .A1(n5827), .A2(n5832), .ZN(n4908) );
  NAND2_X1 U6300 ( .A1(n4911), .A2(n10373), .ZN(n7291) );
  INV_X1 U6301 ( .A(n7289), .ZN(n4911) );
  NAND2_X1 U6302 ( .A1(n6826), .A2(n4510), .ZN(n6833) );
  NAND2_X1 U6303 ( .A1(n9424), .A2(n4926), .ZN(n4925) );
  NAND2_X1 U6304 ( .A1(n4936), .A2(n4932), .ZN(n4931) );
  INV_X1 U6305 ( .A(n4936), .ZN(n8259) );
  NAND2_X1 U6306 ( .A1(n8423), .A2(n4939), .ZN(n4938) );
  INV_X1 U6307 ( .A(n4941), .ZN(n8422) );
  NAND2_X1 U6308 ( .A1(n9494), .A2(n4948), .ZN(n4947) );
  INV_X1 U6309 ( .A(n4953), .ZN(n9493) );
  NAND2_X1 U6310 ( .A1(n7171), .A2(n7170), .ZN(n7238) );
  NAND2_X1 U6311 ( .A1(n7260), .A2(n7259), .ZN(n7262) );
  NAND2_X1 U6312 ( .A1(n7754), .A2(n4957), .ZN(n4954) );
  NAND2_X1 U6313 ( .A1(n4954), .A2(n4955), .ZN(n7918) );
  AND2_X1 U6314 ( .A1(n7815), .A2(n4958), .ZN(n4957) );
  NAND2_X1 U6315 ( .A1(n7754), .A2(n7753), .ZN(n10236) );
  NOR2_X1 U6316 ( .A1(n7756), .A2(n4961), .ZN(n4960) );
  INV_X1 U6317 ( .A(n7753), .ZN(n4961) );
  NOR2_X2 U6318 ( .A1(n4963), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n4962) );
  NAND2_X1 U6319 ( .A1(n7316), .A2(n4965), .ZN(n4964) );
  NAND2_X1 U6320 ( .A1(n4964), .A2(n4966), .ZN(n7751) );
  INV_X1 U6321 ( .A(n4986), .ZN(n8228) );
  NAND2_X1 U6322 ( .A1(n7348), .A2(n4990), .ZN(n4988) );
  NAND2_X1 U6323 ( .A1(n7543), .A2(n6562), .ZN(n4994) );
  OAI21_X1 U6324 ( .B1(n9765), .B2(n5005), .A(n5002), .ZN(n6657) );
  NAND2_X1 U6325 ( .A1(n9765), .A2(n5002), .ZN(n5001) );
  NAND3_X1 U6326 ( .A1(n9774), .A2(n5011), .A3(n6665), .ZN(n5010) );
  NAND2_X1 U6327 ( .A1(n5843), .A2(n5845), .ZN(n5850) );
  NAND2_X1 U6328 ( .A1(n5843), .A2(n5012), .ZN(n10153) );
  NAND3_X1 U6329 ( .A1(n6591), .A2(n5017), .A3(n6590), .ZN(n5015) );
  NAND2_X1 U6330 ( .A1(n6591), .A2(n6590), .ZN(n7982) );
  NOR2_X1 U6331 ( .A1(n7979), .A2(n7980), .ZN(n5016) );
  NAND2_X1 U6332 ( .A1(n7979), .A2(n7980), .ZN(n5017) );
  NAND2_X1 U6333 ( .A1(n9732), .A2(n5021), .ZN(n5018) );
  OAI211_X1 U6334 ( .C1(n9732), .C2(n5022), .A(n5019), .B(n5018), .ZN(P1_U3212) );
  NAND2_X1 U6335 ( .A1(n9740), .A2(n6620), .ZN(n6626) );
  INV_X1 U6336 ( .A(n9361), .ZN(n5032) );
  OAI21_X1 U6337 ( .B1(n5032), .B2(n5036), .A(n5035), .ZN(n8932) );
  AOI21_X1 U6338 ( .B1(n9361), .B2(n6818), .A(n9102), .ZN(n8922) );
  NAND2_X1 U6339 ( .A1(n8933), .A2(n9116), .ZN(n5040) );
  AOI21_X1 U6340 ( .B1(n5039), .B2(n5038), .A(n8969), .ZN(n5037) );
  NAND2_X1 U6341 ( .A1(n5041), .A2(n4546), .ZN(n6815) );
  NAND2_X1 U6342 ( .A1(n7910), .A2(n9041), .ZN(n5046) );
  AOI21_X1 U6343 ( .B1(n9516), .B2(n4541), .A(n5048), .ZN(n9460) );
  OAI21_X1 U6344 ( .B1(n8354), .B2(n5054), .A(n5053), .ZN(n9555) );
  INV_X1 U6345 ( .A(n5551), .ZN(n5118) );
  XNOR2_X1 U6346 ( .A(n5674), .B(n5672), .ZN(n7949) );
  AND2_X1 U6347 ( .A1(n10467), .A2(n5803), .ZN(n10475) );
  NAND2_X1 U6348 ( .A1(n9141), .A2(n5734), .ZN(n5790) );
  OAI21_X2 U6349 ( .B1(n8149), .B2(n8148), .A(n8147), .ZN(n8151) );
  NAND2_X1 U6350 ( .A1(n9435), .A2(n6781), .ZN(n9426) );
  NAND2_X1 U6351 ( .A1(n9437), .A2(n9436), .ZN(n9435) );
  OR2_X1 U6352 ( .A1(n7733), .A2(n9021), .ZN(n7895) );
  NAND2_X1 U6353 ( .A1(n9534), .A2(n5071), .ZN(n6776) );
  NAND2_X1 U6354 ( .A1(n7506), .A2(n6764), .ZN(n7733) );
  AND2_X1 U6355 ( .A1(n6695), .A2(n6697), .ZN(n10353) );
  INV_X1 U6356 ( .A(n9913), .ZN(n10262) );
  INV_X1 U6357 ( .A(n7068), .ZN(n6494) );
  NAND2_X1 U6358 ( .A1(n9529), .A2(n9078), .ZN(n9516) );
  INV_X1 U6359 ( .A(n7067), .ZN(n6493) );
  OAI22_X1 U6360 ( .A1(n7570), .A2(n8945), .B1(n7581), .B2(n9274), .ZN(n7507)
         );
  NAND2_X1 U6361 ( .A1(n7614), .A2(n6792), .ZN(n7509) );
  NAND2_X1 U6362 ( .A1(n6410), .A2(n6736), .ZN(n6488) );
  NOR2_X1 U6363 ( .A1(n6762), .A2(n6761), .ZN(n5060) );
  AND3_X1 U6364 ( .A1(n8296), .A2(n8297), .A3(n8299), .ZN(n5061) );
  OR2_X1 U6365 ( .A1(n4793), .A2(n9640), .ZN(n5063) );
  OR2_X1 U6366 ( .A1(n4793), .A2(n9692), .ZN(n5064) );
  INV_X1 U6367 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5215) );
  AND2_X1 U6368 ( .A1(n5374), .A2(n5354), .ZN(n5065) );
  NOR2_X1 U6369 ( .A1(n6038), .A2(n6037), .ZN(n5066) );
  AND2_X1 U6370 ( .A1(n5458), .A2(n5435), .ZN(n5067) );
  AND2_X1 U6371 ( .A1(n7284), .A2(n7166), .ZN(n5068) );
  AND2_X1 U6372 ( .A1(n9023), .A2(n10505), .ZN(n5069) );
  AND2_X1 U6373 ( .A1(n5211), .A2(n5210), .ZN(n5070) );
  OR2_X1 U6374 ( .A1(n9689), .A2(n9163), .ZN(n5071) );
  INV_X1 U6375 ( .A(n9689), .ZN(n9545) );
  AND2_X1 U6376 ( .A1(n5671), .A2(n5670), .ZN(n5072) );
  AND4_X1 U6377 ( .A1(n5562), .A2(n5561), .A3(n5560), .A4(n5559), .ZN(n9163)
         );
  NOR2_X1 U6378 ( .A1(n9798), .A2(n9799), .ZN(n5073) );
  AND2_X1 U6379 ( .A1(n7735), .A2(n9021), .ZN(n6794) );
  NOR2_X1 U6380 ( .A1(n6760), .A2(n6759), .ZN(n6761) );
  INV_X1 U6381 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5088) );
  NOR2_X1 U6382 ( .A1(n5093), .A2(n5092), .ZN(n5094) );
  INV_X1 U6383 ( .A(n6393), .ZN(n6398) );
  INV_X1 U6384 ( .A(n9945), .ZN(n8490) );
  INV_X1 U6385 ( .A(n7418), .ZN(n5207) );
  INV_X1 U6386 ( .A(n5509), .ZN(n5080) );
  INV_X1 U6387 ( .A(n5511), .ZN(n5081) );
  INV_X1 U6388 ( .A(n7467), .ZN(n8941) );
  INV_X1 U6389 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5087) );
  OR2_X1 U6390 ( .A1(n6083), .A2(n7030), .ZN(n6069) );
  AND2_X1 U6391 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6130) );
  INV_X1 U6392 ( .A(n7169), .ZN(n7170) );
  NAND2_X1 U6393 ( .A1(n6233), .A2(SI_29_), .ZN(n6234) );
  INV_X1 U6394 ( .A(n5592), .ZN(n5593) );
  INV_X1 U6395 ( .A(n5481), .ZN(n5482) );
  AND2_X1 U6396 ( .A1(n5347), .A2(n5346), .ZN(n5348) );
  INV_X1 U6397 ( .A(n5284), .ZN(n5285) );
  OR2_X1 U6398 ( .A1(n5617), .A2(n5084), .ZN(n5618) );
  INV_X1 U6399 ( .A(n8478), .ZN(n5110) );
  INV_X1 U6400 ( .A(n9425), .ZN(n9419) );
  NAND2_X1 U6401 ( .A1(n5085), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5665) );
  OR2_X1 U6402 ( .A1(n5407), .A2(n5406), .ZN(n5409) );
  INV_X1 U6403 ( .A(n10494), .ZN(n9214) );
  OR2_X1 U6404 ( .A1(n6016), .A2(n8697), .ZN(n6003) );
  NAND2_X1 U6405 ( .A1(n9773), .A2(n9776), .ZN(n6665) );
  NOR2_X1 U6406 ( .A1(n6069), .A2(n6051), .ZN(n6053) );
  AND2_X1 U6407 ( .A1(n10087), .A2(n10021), .ZN(n8486) );
  INV_X1 U6408 ( .A(n7239), .ZN(n7240) );
  OR3_X1 U6409 ( .A1(n5972), .A2(P1_IR_REG_15__SCAN_IN), .A3(
        P1_IR_REG_14__SCAN_IN), .ZN(n5960) );
  NAND2_X1 U6410 ( .A1(n5381), .A2(n5380), .ZN(n5430) );
  AND2_X1 U6411 ( .A1(n5734), .A2(n5732), .ZN(n9137) );
  OR2_X1 U6412 ( .A1(n5788), .A2(n5787), .ZN(n5789) );
  INV_X1 U6413 ( .A(n5670), .ZN(n5662) );
  OR2_X1 U6414 ( .A1(n5700), .A2(n9246), .ZN(n5721) );
  OR2_X1 U6415 ( .A1(n10450), .A2(n5801), .ZN(n7678) );
  NAND2_X1 U6416 ( .A1(n9689), .A2(n9163), .ZN(n6775) );
  OR2_X1 U6417 ( .A1(n7963), .A2(n8951), .ZN(n8023) );
  OR2_X1 U6418 ( .A1(n7007), .A2(n5800), .ZN(n9204) );
  INV_X1 U6419 ( .A(n10475), .ZN(n10518) );
  NOR2_X1 U6420 ( .A1(n6003), .A2(n5989), .ZN(n5991) );
  AND2_X1 U6421 ( .A1(n6685), .A2(n6684), .ZN(n6690) );
  NAND2_X1 U6422 ( .A1(n6494), .A2(n6493), .ZN(n7073) );
  OR2_X1 U6423 ( .A1(n5897), .A2(n8539), .ZN(n6198) );
  INV_X1 U6424 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9904) );
  OR2_X1 U6425 ( .A1(n10368), .A2(n7095), .ZN(n6996) );
  XNOR2_X1 U6426 ( .A(n5484), .B(SI_14_), .ZN(n5481) );
  NOR2_X1 U6427 ( .A1(n9367), .A2(n9230), .ZN(n5812) );
  INV_X1 U6428 ( .A(n9245), .ZN(n9390) );
  AND4_X1 U6429 ( .A1(n5604), .A2(n5603), .A3(n5602), .A4(n5601), .ZN(n9180)
         );
  INV_X1 U6430 ( .A(n10440), .ZN(n10442) );
  INV_X1 U6431 ( .A(n9552), .ZN(n10221) );
  AND2_X1 U6432 ( .A1(n10458), .A2(n5763), .ZN(n7377) );
  OR2_X1 U6433 ( .A1(n10528), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6832) );
  NOR2_X1 U6434 ( .A1(n6830), .A2(n6829), .ZN(n6836) );
  NAND2_X1 U6435 ( .A1(n7675), .A2(n10465), .ZN(n10450) );
  INV_X1 U6436 ( .A(n9732), .ZN(n9800) );
  AND4_X1 U6437 ( .A1(n5878), .A2(n5877), .A3(n5876), .A4(n5875), .ZN(n9945)
         );
  AND4_X1 U6438 ( .A1(n5920), .A2(n5919), .A3(n5918), .A4(n5917), .ZN(n9717)
         );
  AND4_X1 U6439 ( .A1(n5969), .A2(n5968), .A3(n5967), .A4(n5966), .ZN(n8316)
         );
  NAND2_X1 U6440 ( .A1(n9959), .A2(n8502), .ZN(n9971) );
  AND2_X1 U6441 ( .A1(n6355), .A2(n8497), .ZN(n10035) );
  OR2_X1 U6442 ( .A1(n6717), .A2(n7140), .ZN(n10368) );
  OR2_X1 U6443 ( .A1(n7978), .A2(n5777), .ZN(n7675) );
  AND2_X1 U6444 ( .A1(n5811), .A2(n5810), .ZN(n9230) );
  INV_X1 U6445 ( .A(n9212), .ZN(n9240) );
  AND2_X1 U6446 ( .A1(n5798), .A2(n5797), .ZN(n7185) );
  AND4_X1 U6447 ( .A1(n5451), .A2(n5450), .A3(n5449), .A4(n5448), .ZN(n9049)
         );
  NAND2_X1 U6448 ( .A1(n9540), .A2(n7391), .ZN(n9552) );
  AND2_X1 U6449 ( .A1(n8267), .A2(n8266), .ZN(n10230) );
  NAND2_X1 U6450 ( .A1(n10541), .A2(n10475), .ZN(n9640) );
  INV_X1 U6451 ( .A(n10541), .ZN(n10539) );
  INV_X1 U6452 ( .A(n9402), .ZN(n9660) );
  INV_X1 U6453 ( .A(n10528), .ZN(n10526) );
  INV_X1 U6454 ( .A(n10460), .ZN(n10462) );
  XNOR2_X1 U6455 ( .A(n5755), .B(n5754), .ZN(n7978) );
  INV_X1 U6456 ( .A(n10098), .ZN(n10032) );
  OR2_X1 U6457 ( .A1(n6472), .A2(n6471), .ZN(n6473) );
  AND4_X1 U6458 ( .A1(n5869), .A2(n5868), .A3(n5867), .A4(n5866), .ZN(n9927)
         );
  INV_X1 U6459 ( .A(n7155), .ZN(n9828) );
  AOI21_X1 U6460 ( .B1(n8513), .B2(n10343), .A(n8512), .ZN(n8872) );
  INV_X1 U6461 ( .A(n10424), .ZN(n10422) );
  INV_X1 U6462 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n8753) );
  CLKBUF_X2 U6463 ( .A(n8243), .Z(n10157) );
  NAND2_X1 U6464 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5245) );
  INV_X1 U6465 ( .A(n5245), .ZN(n5074) );
  NAND2_X1 U6466 ( .A1(n5074), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5276) );
  INV_X1 U6467 ( .A(n5276), .ZN(n5076) );
  AND2_X1 U6468 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_REG3_REG_6__SCAN_IN), 
        .ZN(n5075) );
  NAND2_X1 U6469 ( .A1(n5076), .A2(n5075), .ZN(n5312) );
  INV_X1 U6470 ( .A(n5312), .ZN(n5077) );
  NAND2_X1 U6471 ( .A1(n5077), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5336) );
  INV_X1 U6472 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5335) );
  INV_X1 U6473 ( .A(n5359), .ZN(n5078) );
  NAND2_X1 U6474 ( .A1(n5078), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5407) );
  INV_X1 U6475 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5406) );
  INV_X1 U6476 ( .A(n5409), .ZN(n5079) );
  NAND2_X1 U6477 ( .A1(n5079), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5445) );
  INV_X1 U6478 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5444) );
  INV_X1 U6479 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5468) );
  NAND2_X1 U6480 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_REG3_REG_18__SCAN_IN), 
        .ZN(n5082) );
  NAND2_X1 U6481 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(P2_REG3_REG_20__SCAN_IN), 
        .ZN(n5084) );
  XNOR2_X1 U6482 ( .A(n5665), .B(P2_REG3_REG_23__SCAN_IN), .ZN(n9453) );
  AND2_X2 U6483 ( .A1(n5261), .A2(n5087), .ZN(n5290) );
  INV_X1 U6484 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5089) );
  NAND4_X1 U6485 ( .A1(n5089), .A2(n5400), .A3(n5384), .A4(n5459), .ZN(n5093)
         );
  INV_X1 U6486 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5091) );
  INV_X1 U6487 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5090) );
  NAND4_X1 U6488 ( .A1(n5438), .A2(n5462), .A3(n5091), .A4(n5090), .ZN(n5092)
         );
  INV_X1 U6489 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5778) );
  INV_X1 U6490 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5127) );
  INV_X1 U6491 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5095) );
  AND3_X1 U6492 ( .A1(n5778), .A2(n5127), .A3(n5095), .ZN(n5099) );
  NOR2_X1 U6493 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5098) );
  NOR2_X1 U6494 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5097) );
  NOR2_X1 U6495 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n5096) );
  INV_X1 U6496 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5100) );
  INV_X1 U6497 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5146) );
  INV_X1 U6498 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5104) );
  XNOR2_X1 U6499 ( .A(n5108), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5106) );
  XNOR2_X2 U6500 ( .A(n5105), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5109) );
  INV_X1 U6501 ( .A(n5792), .ZN(n5705) );
  NAND2_X1 U6502 ( .A1(n9453), .A2(n5705), .ZN(n5115) );
  NAND2_X2 U6503 ( .A1(n5109), .A2(n8478), .ZN(n7014) );
  INV_X1 U6504 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9608) );
  NAND2_X1 U6505 ( .A1(n5189), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5112) );
  INV_X1 U6506 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8551) );
  OR2_X1 U6507 ( .A1(n5311), .A2(n8551), .ZN(n5111) );
  OAI211_X1 U6508 ( .C1(n7014), .C2(n9608), .A(n5112), .B(n5111), .ZN(n5113)
         );
  INV_X1 U6509 ( .A(n5113), .ZN(n5114) );
  NAND2_X1 U6510 ( .A1(n5115), .A2(n5114), .ZN(n9258) );
  INV_X1 U6511 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5116) );
  INV_X1 U6512 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5117) );
  NOR2_X1 U6513 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5120) );
  AND2_X1 U6514 ( .A1(n5120), .A2(n5095), .ZN(n5119) );
  INV_X1 U6515 ( .A(n9131), .ZN(n8902) );
  NAND2_X1 U6516 ( .A1(n5123), .A2(n5120), .ZN(n5121) );
  NAND2_X1 U6517 ( .A1(n5121), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5122) );
  XNOR2_X1 U6518 ( .A(n5122), .B(P2_IR_REG_21__SCAN_IN), .ZN(n5155) );
  NAND2_X1 U6519 ( .A1(n5128), .A2(n5127), .ZN(n5124) );
  NAND2_X1 U6520 ( .A1(n5124), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5126) );
  INV_X1 U6521 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5125) );
  XNOR2_X1 U6522 ( .A(n5128), .B(n5127), .ZN(n5153) );
  NAND2_X1 U6523 ( .A1(n9258), .A2(n8938), .ZN(n9152) );
  INV_X1 U6524 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n9470) );
  OR2_X1 U6525 ( .A1(n5311), .A2(n9470), .ZN(n5130) );
  INV_X1 U6526 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9674) );
  OR2_X1 U6527 ( .A1(n4498), .A2(n9674), .ZN(n5129) );
  AND2_X1 U6528 ( .A1(n5130), .A2(n5129), .ZN(n5134) );
  INV_X1 U6529 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9231) );
  NAND2_X1 U6530 ( .A1(n5618), .A2(n9231), .ZN(n5131) );
  NAND2_X1 U6531 ( .A1(n5665), .A2(n5131), .ZN(n9469) );
  OR2_X1 U6532 ( .A1(n9469), .A2(n5792), .ZN(n5133) );
  NAND2_X1 U6533 ( .A1(n6820), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5132) );
  INV_X1 U6534 ( .A(n9181), .ZN(n9259) );
  NAND2_X1 U6535 ( .A1(n7013), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5140) );
  INV_X1 U6536 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7662) );
  OR2_X1 U6537 ( .A1(n5792), .A2(n7662), .ZN(n5139) );
  INV_X1 U6538 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5135) );
  OR2_X1 U6539 ( .A1(n4498), .A2(n5135), .ZN(n5138) );
  INV_X1 U6540 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n5136) );
  INV_X1 U6541 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5142) );
  NAND2_X1 U6542 ( .A1(n5143), .A2(n5142), .ZN(n5145) );
  AND2_X1 U6543 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5144) );
  AND2_X1 U6544 ( .A1(n5145), .A2(n5159), .ZN(n9700) );
  NAND2_X1 U6545 ( .A1(n5148), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5149) );
  MUX2_X1 U6546 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5149), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5152) );
  INV_X1 U6547 ( .A(n5150), .ZN(n5151) );
  MUX2_X1 U6548 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9700), .S(n7723), .Z(n10466)
         );
  NAND2_X1 U6549 ( .A1(n9281), .A2(n10466), .ZN(n7452) );
  INV_X1 U6550 ( .A(n10467), .ZN(n5154) );
  NAND2_X1 U6551 ( .A1(n9131), .A2(n9565), .ZN(n8967) );
  NAND3_X1 U6552 ( .A1(n5154), .A2(n8931), .A3(n8967), .ZN(n5156) );
  NAND2_X1 U6553 ( .A1(n5155), .A2(n8942), .ZN(n7389) );
  INV_X1 U6554 ( .A(n10466), .ZN(n7655) );
  NAND2_X1 U6555 ( .A1(n5576), .A2(n7655), .ZN(n5157) );
  AND2_X1 U6556 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5158) );
  NAND2_X1 U6557 ( .A1(n5175), .A2(n5158), .ZN(n6158) );
  MUX2_X1 U6558 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5175), .Z(n5173) );
  XNOR2_X1 U6559 ( .A(n5172), .B(n5173), .ZN(n6148) );
  NAND2_X1 U6560 ( .A1(n4503), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5162) );
  NAND2_X1 U6561 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5160) );
  NAND2_X1 U6562 ( .A1(n7009), .A2(n7704), .ZN(n5161) );
  NAND2_X1 U6563 ( .A1(n7013), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5168) );
  INV_X1 U6564 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n8132) );
  OR2_X1 U6565 ( .A1(n5792), .A2(n8132), .ZN(n5167) );
  INV_X1 U6566 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5164) );
  OR2_X1 U6567 ( .A1(n4498), .A2(n5164), .ZN(n5166) );
  INV_X1 U6568 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7705) );
  AND2_X1 U6569 ( .A1(n9279), .A2(n8938), .ZN(n5169) );
  INV_X1 U6570 ( .A(n5169), .ZN(n5170) );
  NAND2_X1 U6571 ( .A1(n7584), .A2(n5170), .ZN(n5171) );
  NAND2_X1 U6572 ( .A1(n7370), .A2(n5171), .ZN(n5184) );
  XNOR2_X1 U6573 ( .A(n5197), .B(n5195), .ZN(n6169) );
  NAND2_X1 U6574 ( .A1(n4504), .A2(n6169), .ZN(n5179) );
  NAND2_X1 U6575 ( .A1(n5240), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5178) );
  NAND2_X1 U6576 ( .A1(n7009), .A2(n10164), .ZN(n5177) );
  XNOR2_X1 U6577 ( .A(n10482), .B(n5661), .ZN(n5187) );
  NAND2_X1 U6578 ( .A1(n7013), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5183) );
  NAND2_X1 U6579 ( .A1(n5189), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5182) );
  INV_X1 U6580 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7474) );
  OR2_X1 U6581 ( .A1(n5792), .A2(n7474), .ZN(n5181) );
  INV_X1 U6582 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7703) );
  OR2_X1 U6583 ( .A1(n7014), .A2(n7703), .ZN(n5180) );
  AND2_X1 U6584 ( .A1(n9278), .A2(n8938), .ZN(n5185) );
  XNOR2_X1 U6585 ( .A(n5187), .B(n5185), .ZN(n7586) );
  INV_X1 U6586 ( .A(n5185), .ZN(n5186) );
  NAND2_X1 U6587 ( .A1(n5187), .A2(n5186), .ZN(n5188) );
  NAND2_X1 U6588 ( .A1(n7013), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5194) );
  OR2_X1 U6589 ( .A1(n5792), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5193) );
  INV_X1 U6590 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5190) );
  INV_X1 U6591 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7702) );
  OR2_X1 U6592 ( .A1(n7014), .A2(n7702), .ZN(n5191) );
  NAND2_X1 U6593 ( .A1(n9277), .A2(n8938), .ZN(n5205) );
  INV_X1 U6594 ( .A(n5195), .ZN(n5196) );
  NAND2_X1 U6595 ( .A1(n5197), .A2(n5196), .ZN(n5213) );
  NAND2_X1 U6596 ( .A1(n5198), .A2(SI_2_), .ZN(n5209) );
  NAND2_X1 U6597 ( .A1(n5213), .A2(n5209), .ZN(n5200) );
  MUX2_X1 U6598 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n5199), .Z(n5208) );
  XNOR2_X1 U6599 ( .A(n5208), .B(SI_3_), .ZN(n5210) );
  XNOR2_X1 U6600 ( .A(n5200), .B(n5210), .ZN(n6100) );
  NAND2_X1 U6601 ( .A1(n4504), .A2(n6100), .ZN(n5204) );
  NAND2_X1 U6602 ( .A1(n5240), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5203) );
  NAND2_X1 U6603 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4529), .ZN(n5201) );
  XNOR2_X1 U6604 ( .A(n5201), .B(P2_IR_REG_3__SCAN_IN), .ZN(n7708) );
  NAND2_X1 U6605 ( .A1(n7009), .A2(n7708), .ZN(n5202) );
  XNOR2_X1 U6606 ( .A(n10489), .B(n5661), .ZN(n9222) );
  OR2_X1 U6607 ( .A1(n5205), .A2(n9222), .ZN(n5227) );
  NAND2_X1 U6608 ( .A1(n9222), .A2(n5205), .ZN(n5206) );
  NAND2_X1 U6609 ( .A1(n5227), .A2(n5206), .ZN(n7418) );
  NAND2_X1 U6610 ( .A1(n5208), .A2(SI_3_), .ZN(n5211) );
  AND2_X1 U6611 ( .A1(n5209), .A2(n5211), .ZN(n5212) );
  XNOR2_X1 U6612 ( .A(n5235), .B(n5233), .ZN(n6136) );
  NAND2_X1 U6613 ( .A1(n4504), .A2(n6136), .ZN(n5222) );
  NAND2_X1 U6614 ( .A1(n5240), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5221) );
  NAND2_X1 U6615 ( .A1(n5216), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5217) );
  MUX2_X1 U6616 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5217), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n5219) );
  AND2_X1 U6617 ( .A1(n5219), .A2(n5218), .ZN(n7709) );
  NAND2_X1 U6618 ( .A1(n7009), .A2(n7709), .ZN(n5220) );
  XNOR2_X1 U6619 ( .A(n10494), .B(n5661), .ZN(n5231) );
  NAND2_X1 U6620 ( .A1(n7013), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5226) );
  OAI21_X1 U6621 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n5245), .ZN(n7619) );
  OR2_X1 U6622 ( .A1(n5792), .A2(n7619), .ZN(n5225) );
  INV_X1 U6623 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5223) );
  AND2_X1 U6624 ( .A1(n9276), .A2(n8938), .ZN(n5229) );
  XNOR2_X1 U6625 ( .A(n5231), .B(n5229), .ZN(n9221) );
  AND2_X1 U6626 ( .A1(n9221), .A2(n5227), .ZN(n5228) );
  NAND2_X1 U6627 ( .A1(n7415), .A2(n5228), .ZN(n9211) );
  INV_X1 U6628 ( .A(n5229), .ZN(n5230) );
  NAND2_X1 U6629 ( .A1(n5231), .A2(n5230), .ZN(n5232) );
  INV_X1 U6630 ( .A(n5233), .ZN(n5234) );
  NAND2_X1 U6631 ( .A1(n5235), .A2(n5234), .ZN(n5238) );
  NAND2_X1 U6632 ( .A1(n5236), .A2(SI_4_), .ZN(n5237) );
  INV_X1 U6633 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n5239) );
  INV_X1 U6634 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6924) );
  MUX2_X1 U6635 ( .A(n5239), .B(n6924), .S(n6889), .Z(n5258) );
  XNOR2_X1 U6636 ( .A(n5257), .B(n5256), .ZN(n6925) );
  NAND2_X1 U6637 ( .A1(n5240), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5243) );
  NAND2_X1 U6638 ( .A1(n5218), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5241) );
  XNOR2_X1 U6639 ( .A(n5241), .B(P2_IR_REG_5__SCAN_IN), .ZN(n8216) );
  NAND2_X1 U6640 ( .A1(n7009), .A2(n8216), .ZN(n5242) );
  OAI211_X1 U6641 ( .C1(n4505), .C2(n6925), .A(n5243), .B(n5242), .ZN(n7524)
         );
  XNOR2_X1 U6642 ( .A(n7539), .B(n5661), .ZN(n5254) );
  NAND2_X1 U6643 ( .A1(n7013), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5251) );
  INV_X1 U6644 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5244) );
  OR2_X1 U6645 ( .A1(n7014), .A2(n5244), .ZN(n5250) );
  INV_X1 U6646 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8207) );
  NAND2_X1 U6647 ( .A1(n5245), .A2(n8207), .ZN(n5246) );
  NAND2_X1 U6648 ( .A1(n5276), .A2(n5246), .ZN(n7527) );
  OR2_X1 U6649 ( .A1(n5792), .A2(n7527), .ZN(n5249) );
  INV_X1 U6650 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5247) );
  OR2_X1 U6651 ( .A1(n4498), .A2(n5247), .ZN(n5248) );
  NAND2_X1 U6652 ( .A1(n9275), .A2(n8938), .ZN(n5253) );
  NAND2_X1 U6653 ( .A1(n5254), .A2(n5253), .ZN(n5252) );
  INV_X1 U6654 ( .A(n5253), .ZN(n5255) );
  INV_X1 U6655 ( .A(n5254), .ZN(n7522) );
  NAND2_X1 U6656 ( .A1(n5255), .A2(n7522), .ZN(n7529) );
  INV_X1 U6657 ( .A(n5258), .ZN(n5259) );
  NAND2_X1 U6658 ( .A1(n5259), .A2(SI_5_), .ZN(n5260) );
  MUX2_X1 U6659 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6889), .Z(n5287) );
  XNOR2_X1 U6660 ( .A(n5286), .B(n5284), .ZN(n6894) );
  NAND2_X1 U6661 ( .A1(n4504), .A2(n6894), .ZN(n5265) );
  NAND2_X1 U6662 ( .A1(n5240), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n5264) );
  OR2_X1 U6663 ( .A1(n5261), .A2(n9696), .ZN(n5262) );
  XNOR2_X1 U6664 ( .A(n5262), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7712) );
  NAND2_X1 U6665 ( .A1(n7009), .A2(n7712), .ZN(n5263) );
  XNOR2_X1 U6666 ( .A(n10501), .B(n5661), .ZN(n5273) );
  NAND2_X1 U6667 ( .A1(n7013), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5270) );
  INV_X1 U6668 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7713) );
  OR2_X1 U6669 ( .A1(n7014), .A2(n7713), .ZN(n5269) );
  INV_X1 U6670 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5275) );
  XNOR2_X1 U6671 ( .A(n5276), .B(n5275), .ZN(n7574) );
  OR2_X1 U6672 ( .A1(n5792), .A2(n7574), .ZN(n5268) );
  INV_X1 U6673 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5266) );
  OR2_X1 U6674 ( .A1(n4498), .A2(n5266), .ZN(n5267) );
  NAND4_X1 U6675 ( .A1(n5270), .A2(n5269), .A3(n5268), .A4(n5267), .ZN(n9274)
         );
  AND2_X1 U6676 ( .A1(n9274), .A2(n8938), .ZN(n5271) );
  XNOR2_X1 U6677 ( .A(n5273), .B(n5271), .ZN(n7559) );
  INV_X1 U6678 ( .A(n5271), .ZN(n5272) );
  NAND2_X1 U6679 ( .A1(n5273), .A2(n5272), .ZN(n5274) );
  NAND2_X1 U6680 ( .A1(n7013), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5283) );
  INV_X1 U6681 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7701) );
  OR2_X1 U6682 ( .A1(n7014), .A2(n7701), .ZN(n5282) );
  INV_X1 U6683 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7648) );
  OAI21_X1 U6684 ( .B1(n5276), .B2(n5275), .A(n7648), .ZN(n5277) );
  NAND2_X1 U6685 ( .A1(n5277), .A2(n5312), .ZN(n7654) );
  OR2_X1 U6686 ( .A1(n5792), .A2(n7654), .ZN(n5281) );
  INV_X1 U6687 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n5278) );
  OR2_X1 U6688 ( .A1(n4498), .A2(n5278), .ZN(n5280) );
  NAND2_X1 U6689 ( .A1(n9273), .A2(n8938), .ZN(n5295) );
  NAND2_X1 U6690 ( .A1(n5287), .A2(SI_6_), .ZN(n5288) );
  MUX2_X1 U6691 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6889), .Z(n5300) );
  XNOR2_X1 U6692 ( .A(n5299), .B(n5297), .ZN(n6907) );
  NAND2_X1 U6693 ( .A1(n4504), .A2(n6907), .ZN(n5294) );
  NAND2_X1 U6694 ( .A1(n5240), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n5293) );
  OR2_X1 U6695 ( .A1(n5290), .A2(n9696), .ZN(n5291) );
  XNOR2_X1 U6696 ( .A(n5291), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7700) );
  NAND2_X1 U6697 ( .A1(n7009), .A2(n7700), .ZN(n5292) );
  XNOR2_X1 U6698 ( .A(n7633), .B(n5661), .ZN(n7780) );
  OR2_X1 U6699 ( .A1(n5295), .A2(n7780), .ZN(n5324) );
  NAND2_X1 U6700 ( .A1(n7780), .A2(n5295), .ZN(n5296) );
  NAND2_X1 U6701 ( .A1(n5324), .A2(n5296), .ZN(n7645) );
  NAND2_X1 U6702 ( .A1(n5300), .A2(SI_7_), .ZN(n5301) );
  INV_X1 U6703 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6914) );
  MUX2_X1 U6704 ( .A(n6914), .B(n6921), .S(n6889), .Z(n5303) );
  INV_X1 U6705 ( .A(SI_8_), .ZN(n5302) );
  NAND2_X1 U6706 ( .A1(n5303), .A2(n5302), .ZN(n5347) );
  INV_X1 U6707 ( .A(n5303), .ZN(n5304) );
  NAND2_X1 U6708 ( .A1(n5304), .A2(SI_8_), .ZN(n5305) );
  XNOR2_X1 U6709 ( .A(n5325), .B(n5326), .ZN(n6913) );
  NAND2_X1 U6710 ( .A1(n6913), .A2(n4504), .ZN(n5310) );
  NAND2_X1 U6711 ( .A1(n5306), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5307) );
  MUX2_X1 U6712 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5307), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n5308) );
  AND2_X1 U6713 ( .A1(n5308), .A2(n5355), .ZN(n7715) );
  AOI22_X1 U6714 ( .A1(n5240), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7009), .B2(
        n7715), .ZN(n5309) );
  XNOR2_X1 U6715 ( .A(n5576), .B(n10505), .ZN(n5319) );
  NAND2_X1 U6716 ( .A1(n6820), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5318) );
  INV_X1 U6717 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7743) );
  OR2_X1 U6718 ( .A1(n5311), .A2(n7743), .ZN(n5317) );
  INV_X1 U6719 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8815) );
  NAND2_X1 U6720 ( .A1(n5312), .A2(n8815), .ZN(n5313) );
  NAND2_X1 U6721 ( .A1(n5336), .A2(n5313), .ZN(n7785) );
  OR2_X1 U6722 ( .A1(n5792), .A2(n7785), .ZN(n5316) );
  INV_X1 U6723 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5314) );
  OR2_X1 U6724 ( .A1(n4498), .A2(n5314), .ZN(n5315) );
  NAND2_X1 U6725 ( .A1(n9272), .A2(n8938), .ZN(n5320) );
  NAND2_X1 U6726 ( .A1(n5319), .A2(n5320), .ZN(n5322) );
  INV_X1 U6727 ( .A(n5319), .ZN(n8886) );
  INV_X1 U6728 ( .A(n5320), .ZN(n5321) );
  NAND2_X1 U6729 ( .A1(n8886), .A2(n5321), .ZN(n5343) );
  NAND2_X1 U6730 ( .A1(n5322), .A2(n5343), .ZN(n7777) );
  OR2_X1 U6731 ( .A1(n7645), .A2(n7777), .ZN(n5323) );
  OR2_X1 U6732 ( .A1(n7777), .A2(n5324), .ZN(n7781) );
  NAND2_X1 U6733 ( .A1(n5349), .A2(n5347), .ZN(n5331) );
  INV_X1 U6734 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6931) );
  MUX2_X1 U6735 ( .A(n6931), .B(n8753), .S(n6889), .Z(n5328) );
  INV_X1 U6736 ( .A(SI_9_), .ZN(n5327) );
  NAND2_X1 U6737 ( .A1(n5328), .A2(n5327), .ZN(n5346) );
  INV_X1 U6738 ( .A(n5328), .ZN(n5329) );
  AND2_X1 U6739 ( .A1(n5346), .A2(n5350), .ZN(n5330) );
  XNOR2_X1 U6740 ( .A(n5331), .B(n5330), .ZN(n6930) );
  NAND2_X1 U6741 ( .A1(n6930), .A2(n4504), .ZN(n5334) );
  NAND2_X1 U6742 ( .A1(n5355), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5332) );
  XNOR2_X1 U6743 ( .A(n5332), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7716) );
  AOI22_X1 U6744 ( .A1(n5240), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7009), .B2(
        n7716), .ZN(n5333) );
  NAND2_X1 U6745 ( .A1(n5334), .A2(n5333), .ZN(n8898) );
  XNOR2_X1 U6746 ( .A(n8898), .B(n5576), .ZN(n5372) );
  NAND2_X1 U6747 ( .A1(n6820), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5342) );
  INV_X1 U6748 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7901) );
  OR2_X1 U6749 ( .A1(n5311), .A2(n7901), .ZN(n5341) );
  NAND2_X1 U6750 ( .A1(n5336), .A2(n5335), .ZN(n5337) );
  NAND2_X1 U6751 ( .A1(n5359), .A2(n5337), .ZN(n8892) );
  OR2_X1 U6752 ( .A1(n5792), .A2(n8892), .ZN(n5340) );
  INV_X1 U6753 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5338) );
  OR2_X1 U6754 ( .A1(n4498), .A2(n5338), .ZN(n5339) );
  NOR2_X1 U6755 ( .A1(n7808), .A2(n7521), .ZN(n5370) );
  XNOR2_X1 U6756 ( .A(n5372), .B(n5370), .ZN(n8889) );
  AND2_X1 U6757 ( .A1(n8889), .A2(n5343), .ZN(n5344) );
  AND2_X1 U6758 ( .A1(n7781), .A2(n5344), .ZN(n5345) );
  INV_X1 U6759 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6978) );
  INV_X1 U6760 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6976) );
  MUX2_X1 U6761 ( .A(n6978), .B(n6976), .S(n6889), .Z(n5352) );
  INV_X1 U6762 ( .A(SI_10_), .ZN(n5351) );
  NAND2_X1 U6763 ( .A1(n5352), .A2(n5351), .ZN(n5374) );
  INV_X1 U6764 ( .A(n5352), .ZN(n5353) );
  NAND2_X1 U6765 ( .A1(n5353), .A2(SI_10_), .ZN(n5354) );
  NAND2_X1 U6766 ( .A1(n6975), .A2(n4504), .ZN(n5357) );
  NAND2_X1 U6767 ( .A1(n5386), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5401) );
  XNOR2_X1 U6768 ( .A(n5401), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7698) );
  AOI22_X1 U6769 ( .A1(n5240), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n7009), .B2(
        n7698), .ZN(n5356) );
  NAND2_X1 U6770 ( .A1(n5357), .A2(n5356), .ZN(n8040) );
  XNOR2_X1 U6771 ( .A(n8040), .B(n5661), .ZN(n5366) );
  NAND2_X1 U6772 ( .A1(n7013), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5365) );
  INV_X1 U6773 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7699) );
  OR2_X1 U6774 ( .A1(n7014), .A2(n7699), .ZN(n5364) );
  INV_X1 U6775 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5358) );
  NAND2_X1 U6776 ( .A1(n5359), .A2(n5358), .ZN(n5360) );
  NAND2_X1 U6777 ( .A1(n5407), .A2(n5360), .ZN(n8032) );
  OR2_X1 U6778 ( .A1(n5792), .A2(n8032), .ZN(n5363) );
  INV_X1 U6779 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5361) );
  OR2_X1 U6780 ( .A1(n4498), .A2(n5361), .ZN(n5362) );
  NOR2_X1 U6781 ( .A1(n8895), .A2(n7521), .ZN(n5367) );
  NAND2_X1 U6782 ( .A1(n5366), .A2(n5367), .ZN(n7935) );
  INV_X1 U6783 ( .A(n5366), .ZN(n7934) );
  INV_X1 U6784 ( .A(n5367), .ZN(n5368) );
  NAND2_X1 U6785 ( .A1(n7934), .A2(n5368), .ZN(n5369) );
  AND2_X1 U6786 ( .A1(n7935), .A2(n5369), .ZN(n7807) );
  INV_X1 U6787 ( .A(n5370), .ZN(n5371) );
  NAND2_X1 U6788 ( .A1(n5372), .A2(n5371), .ZN(n7804) );
  AND2_X1 U6789 ( .A1(n7807), .A2(n7804), .ZN(n7805) );
  NAND2_X1 U6790 ( .A1(n5373), .A2(n5065), .ZN(n5375) );
  INV_X1 U6791 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6995) );
  INV_X1 U6792 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6993) );
  MUX2_X1 U6793 ( .A(n6995), .B(n6993), .S(n6889), .Z(n5376) );
  INV_X1 U6794 ( .A(n5376), .ZN(n5377) );
  INV_X1 U6795 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7041) );
  INV_X1 U6796 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7039) );
  MUX2_X1 U6797 ( .A(n7041), .B(n7039), .S(n6889), .Z(n5381) );
  INV_X1 U6798 ( .A(SI_12_), .ZN(n5380) );
  INV_X1 U6799 ( .A(n5381), .ZN(n5382) );
  NAND2_X1 U6800 ( .A1(n5382), .A2(SI_12_), .ZN(n5383) );
  XNOR2_X1 U6801 ( .A(n5432), .B(n5431), .ZN(n7038) );
  NAND2_X1 U6802 ( .A1(n5400), .A2(n5384), .ZN(n5385) );
  NOR2_X1 U6803 ( .A1(n5386), .A2(n5385), .ZN(n5439) );
  OR2_X1 U6804 ( .A1(n5439), .A2(n9696), .ZN(n5387) );
  XNOR2_X1 U6805 ( .A(n5387), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8203) );
  AOI22_X1 U6806 ( .A1(n5240), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7009), .B2(
        n8203), .ZN(n5388) );
  NAND2_X1 U6807 ( .A1(n5189), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5393) );
  INV_X1 U6808 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7971) );
  OR2_X1 U6809 ( .A1(n5311), .A2(n7971), .ZN(n5392) );
  INV_X1 U6810 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8000) );
  NAND2_X1 U6811 ( .A1(n5409), .A2(n8000), .ZN(n5389) );
  NAND2_X1 U6812 ( .A1(n5445), .A2(n5389), .ZN(n8003) );
  OR2_X1 U6813 ( .A1(n5792), .A2(n8003), .ZN(n5391) );
  INV_X1 U6814 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7719) );
  OR2_X1 U6815 ( .A1(n7014), .A2(n7719), .ZN(n5390) );
  NOR2_X1 U6816 ( .A1(n8051), .A2(n7521), .ZN(n5395) );
  NAND2_X1 U6817 ( .A1(n5394), .A2(n5395), .ZN(n5415) );
  INV_X1 U6818 ( .A(n5395), .ZN(n5396) );
  NAND2_X1 U6819 ( .A1(n8047), .A2(n5396), .ZN(n5397) );
  XNOR2_X1 U6820 ( .A(n5399), .B(n5398), .ZN(n6992) );
  NAND2_X1 U6821 ( .A1(n6992), .A2(n4504), .ZN(n5405) );
  NAND2_X1 U6822 ( .A1(n5401), .A2(n5400), .ZN(n5402) );
  NAND2_X1 U6823 ( .A1(n5402), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5403) );
  XNOR2_X1 U6824 ( .A(n5403), .B(P2_IR_REG_11__SCAN_IN), .ZN(n9287) );
  AOI22_X1 U6825 ( .A1(n5240), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n7009), .B2(
        n9287), .ZN(n5404) );
  NAND2_X1 U6826 ( .A1(n5405), .A2(n5404), .ZN(n7957) );
  XNOR2_X1 U6827 ( .A(n7957), .B(n5661), .ZN(n5416) );
  NAND2_X1 U6828 ( .A1(n7013), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5414) );
  INV_X1 U6829 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7697) );
  OR2_X1 U6830 ( .A1(n7014), .A2(n7697), .ZN(n5413) );
  NAND2_X1 U6831 ( .A1(n5407), .A2(n5406), .ZN(n5408) );
  NAND2_X1 U6832 ( .A1(n5409), .A2(n5408), .ZN(n7952) );
  OR2_X1 U6833 ( .A1(n5792), .A2(n7952), .ZN(n5412) );
  INV_X1 U6834 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n5410) );
  OR2_X1 U6835 ( .A1(n4498), .A2(n5410), .ZN(n5411) );
  NOR2_X1 U6836 ( .A1(n7992), .A2(n7521), .ZN(n5417) );
  NAND2_X1 U6837 ( .A1(n5416), .A2(n5417), .ZN(n5420) );
  INV_X1 U6838 ( .A(n5416), .ZN(n7993) );
  INV_X1 U6839 ( .A(n5417), .ZN(n5418) );
  NAND2_X1 U6840 ( .A1(n7993), .A2(n5418), .ZN(n5419) );
  AND2_X1 U6841 ( .A1(n5420), .A2(n5419), .ZN(n7937) );
  AND2_X1 U6842 ( .A1(n7937), .A2(n5421), .ZN(n7994) );
  AND2_X1 U6843 ( .A1(n7805), .A2(n5424), .ZN(n5423) );
  NAND2_X1 U6844 ( .A1(n8901), .A2(n5423), .ZN(n5429) );
  INV_X1 U6845 ( .A(n5424), .ZN(n5427) );
  AND2_X1 U6846 ( .A1(n7935), .A2(n5425), .ZN(n5426) );
  OR2_X1 U6847 ( .A1(n5427), .A2(n5426), .ZN(n5428) );
  NAND2_X1 U6848 ( .A1(n5429), .A2(n5428), .ZN(n5456) );
  INV_X1 U6849 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7088) );
  INV_X1 U6850 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n7086) );
  MUX2_X1 U6851 ( .A(n7088), .B(n7086), .S(n6889), .Z(n5433) );
  INV_X1 U6852 ( .A(SI_13_), .ZN(n8796) );
  NAND2_X1 U6853 ( .A1(n5433), .A2(n8796), .ZN(n5458) );
  INV_X1 U6854 ( .A(n5433), .ZN(n5434) );
  NAND2_X1 U6855 ( .A1(n5434), .A2(SI_13_), .ZN(n5435) );
  XNOR2_X1 U6856 ( .A(n5457), .B(n5067), .ZN(n7085) );
  NAND2_X1 U6857 ( .A1(n7085), .A2(n4504), .ZN(n5442) );
  NAND2_X1 U6858 ( .A1(n5439), .A2(n5438), .ZN(n5440) );
  NAND2_X1 U6859 ( .A1(n5440), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5460) );
  XNOR2_X1 U6860 ( .A(n5460), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7835) );
  AOI22_X1 U6861 ( .A1(n5240), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n7009), .B2(
        n7835), .ZN(n5441) );
  XNOR2_X1 U6862 ( .A(n10220), .B(n5661), .ZN(n5452) );
  NAND2_X1 U6863 ( .A1(n7013), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5451) );
  INV_X1 U6864 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5443) );
  OR2_X1 U6865 ( .A1(n7014), .A2(n5443), .ZN(n5450) );
  NAND2_X1 U6866 ( .A1(n5445), .A2(n5444), .ZN(n5446) );
  NAND2_X1 U6867 ( .A1(n5469), .A2(n5446), .ZN(n10217) );
  OR2_X1 U6868 ( .A1(n5792), .A2(n10217), .ZN(n5449) );
  INV_X1 U6869 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n5447) );
  OR2_X1 U6870 ( .A1(n4498), .A2(n5447), .ZN(n5448) );
  NOR2_X1 U6871 ( .A1(n9049), .A2(n7521), .ZN(n5453) );
  NAND2_X1 U6872 ( .A1(n5452), .A2(n5453), .ZN(n5475) );
  INV_X1 U6873 ( .A(n5452), .ZN(n8907) );
  INV_X1 U6874 ( .A(n5453), .ZN(n5454) );
  NAND2_X1 U6875 ( .A1(n8907), .A2(n5454), .ZN(n5455) );
  AND2_X1 U6876 ( .A1(n5475), .A2(n5455), .ZN(n8044) );
  NAND2_X1 U6877 ( .A1(n5456), .A2(n8044), .ZN(n8048) );
  INV_X1 U6878 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n8520) );
  INV_X1 U6879 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7110) );
  MUX2_X1 U6880 ( .A(n8520), .B(n7110), .S(n6889), .Z(n5484) );
  XNOR2_X1 U6881 ( .A(n5483), .B(n5481), .ZN(n7109) );
  NAND2_X1 U6882 ( .A1(n7109), .A2(n4504), .ZN(n5466) );
  NAND2_X1 U6883 ( .A1(n5460), .A2(n5459), .ZN(n5461) );
  NAND2_X1 U6884 ( .A1(n5461), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5463) );
  NAND2_X1 U6885 ( .A1(n5463), .A2(n5462), .ZN(n5518) );
  OR2_X1 U6886 ( .A1(n5463), .A2(n5462), .ZN(n5464) );
  AND2_X1 U6887 ( .A1(n5518), .A2(n5464), .ZN(n8079) );
  AOI22_X1 U6888 ( .A1(n5240), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n7009), .B2(
        n8079), .ZN(n5465) );
  XNOR2_X1 U6889 ( .A(n8917), .B(n5576), .ZN(n5479) );
  NAND2_X1 U6890 ( .A1(n5189), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5474) );
  INV_X1 U6891 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n5467) );
  OR2_X1 U6892 ( .A1(n7014), .A2(n5467), .ZN(n5473) );
  INV_X1 U6893 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8171) );
  OR2_X1 U6894 ( .A1(n5311), .A2(n8171), .ZN(n5472) );
  NAND2_X1 U6895 ( .A1(n5469), .A2(n5468), .ZN(n5470) );
  NAND2_X1 U6896 ( .A1(n5509), .A2(n5470), .ZN(n8912) );
  OR2_X1 U6897 ( .A1(n5792), .A2(n8912), .ZN(n5471) );
  NOR2_X1 U6898 ( .A1(n8249), .A2(n7521), .ZN(n5477) );
  XNOR2_X1 U6899 ( .A(n5479), .B(n5477), .ZN(n8908) );
  AND2_X1 U6900 ( .A1(n8908), .A2(n5475), .ZN(n5476) );
  INV_X1 U6901 ( .A(n5477), .ZN(n5478) );
  NAND2_X1 U6902 ( .A1(n5479), .A2(n5478), .ZN(n5480) );
  INV_X1 U6903 ( .A(n5484), .ZN(n5485) );
  NAND2_X1 U6904 ( .A1(n5485), .A2(SI_14_), .ZN(n5486) );
  INV_X1 U6905 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n8653) );
  INV_X1 U6906 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n8662) );
  MUX2_X1 U6907 ( .A(n8653), .B(n8662), .S(n6889), .Z(n5489) );
  INV_X1 U6908 ( .A(SI_15_), .ZN(n5488) );
  INV_X1 U6909 ( .A(n5489), .ZN(n5490) );
  NAND2_X1 U6910 ( .A1(n5490), .A2(SI_15_), .ZN(n5491) );
  INV_X1 U6911 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5493) );
  INV_X1 U6912 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7202) );
  MUX2_X1 U6913 ( .A(n5493), .B(n7202), .S(n6889), .Z(n5494) );
  INV_X1 U6914 ( .A(SI_16_), .ZN(n8684) );
  NAND2_X1 U6915 ( .A1(n5494), .A2(n8684), .ZN(n5529) );
  INV_X1 U6916 ( .A(n5494), .ZN(n5495) );
  NAND2_X1 U6917 ( .A1(n5495), .A2(SI_16_), .ZN(n5496) );
  NAND2_X1 U6918 ( .A1(n7162), .A2(n4504), .ZN(n5500) );
  NAND2_X1 U6919 ( .A1(n5497), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5498) );
  XNOR2_X1 U6920 ( .A(n5498), .B(P2_IR_REG_16__SCAN_IN), .ZN(n9304) );
  AOI22_X1 U6921 ( .A1(n5240), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n7009), .B2(
        n9304), .ZN(n5499) );
  XNOR2_X1 U6922 ( .A(n9066), .B(n5661), .ZN(n8300) );
  NAND2_X1 U6923 ( .A1(n7013), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5506) );
  INV_X1 U6924 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8383) );
  OR2_X1 U6925 ( .A1(n7014), .A2(n8383), .ZN(n5505) );
  INV_X1 U6926 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8387) );
  NAND2_X1 U6927 ( .A1(n5511), .A2(n8387), .ZN(n5501) );
  NAND2_X1 U6928 ( .A1(n5557), .A2(n5501), .ZN(n8425) );
  OR2_X1 U6929 ( .A1(n5792), .A2(n8425), .ZN(n5504) );
  INV_X1 U6930 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n5502) );
  OR2_X1 U6931 ( .A1(n4498), .A2(n5502), .ZN(n5503) );
  NAND4_X1 U6932 ( .A1(n5506), .A2(n5505), .A3(n5504), .A4(n5503), .ZN(n9265)
         );
  AND2_X1 U6933 ( .A1(n9265), .A2(n8938), .ZN(n5524) );
  NAND2_X1 U6934 ( .A1(n5189), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5515) );
  INV_X1 U6935 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n5507) );
  OR2_X1 U6936 ( .A1(n7014), .A2(n5507), .ZN(n5514) );
  INV_X1 U6937 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n5508) );
  OR2_X1 U6938 ( .A1(n5311), .A2(n5508), .ZN(n5513) );
  INV_X1 U6939 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8252) );
  NAND2_X1 U6940 ( .A1(n5509), .A2(n8252), .ZN(n5510) );
  NAND2_X1 U6941 ( .A1(n5511), .A2(n5510), .ZN(n8248) );
  OR2_X1 U6942 ( .A1(n5792), .A2(n8248), .ZN(n5512) );
  NOR2_X1 U6943 ( .A1(n8303), .A2(n7521), .ZN(n5523) );
  XNOR2_X1 U6944 ( .A(n5517), .B(n5516), .ZN(n7160) );
  NAND2_X1 U6945 ( .A1(n7160), .A2(n4504), .ZN(n5521) );
  NAND2_X1 U6946 ( .A1(n5518), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5519) );
  XNOR2_X1 U6947 ( .A(n5519), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8380) );
  AOI22_X1 U6948 ( .A1(n5240), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n8380), .B2(
        n7009), .ZN(n5520) );
  XNOR2_X1 U6949 ( .A(n8361), .B(n5661), .ZN(n8245) );
  AOI22_X1 U6950 ( .A1(n8300), .A2(n5524), .B1(n5523), .B2(n8245), .ZN(n5522)
         );
  INV_X1 U6951 ( .A(n8300), .ZN(n5526) );
  OAI21_X1 U6952 ( .B1(n8245), .B2(n5523), .A(n5524), .ZN(n5525) );
  INV_X1 U6953 ( .A(n8245), .ZN(n8296) );
  INV_X1 U6954 ( .A(n5523), .ZN(n8297) );
  INV_X1 U6955 ( .A(n5524), .ZN(n8299) );
  AOI21_X1 U6956 ( .B1(n5526), .B2(n5525), .A(n5061), .ZN(n5527) );
  MUX2_X1 U6957 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n6889), .Z(n5548) );
  INV_X1 U6958 ( .A(SI_17_), .ZN(n5530) );
  XNOR2_X1 U6959 ( .A(n5548), .B(n5530), .ZN(n5547) );
  XNOR2_X1 U6960 ( .A(n5550), .B(n5547), .ZN(n7228) );
  NAND2_X1 U6961 ( .A1(n7228), .A2(n4504), .ZN(n5534) );
  NAND2_X1 U6962 ( .A1(n4557), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5531) );
  MUX2_X1 U6963 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5531), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n5532) );
  NAND2_X1 U6964 ( .A1(n5532), .A2(n5551), .ZN(n9311) );
  INV_X1 U6965 ( .A(n9311), .ZN(n9313) );
  AOI22_X1 U6966 ( .A1(n5240), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n7009), .B2(
        n9313), .ZN(n5533) );
  XNOR2_X1 U6967 ( .A(n9559), .B(n5661), .ZN(n5541) );
  NAND2_X1 U6968 ( .A1(n6820), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5540) );
  INV_X1 U6969 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n5535) );
  OR2_X1 U6970 ( .A1(n5311), .A2(n5535), .ZN(n5539) );
  INV_X1 U6971 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5556) );
  XNOR2_X1 U6972 ( .A(n5557), .B(n5556), .ZN(n9549) );
  OR2_X1 U6973 ( .A1(n5792), .A2(n9549), .ZN(n5538) );
  INV_X1 U6974 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n5536) );
  OR2_X1 U6975 ( .A1(n4498), .A2(n5536), .ZN(n5537) );
  NOR2_X1 U6976 ( .A1(n8341), .A2(n7521), .ZN(n5542) );
  NAND2_X1 U6977 ( .A1(n5541), .A2(n5542), .ZN(n5546) );
  INV_X1 U6978 ( .A(n5541), .ZN(n8337) );
  INV_X1 U6979 ( .A(n5542), .ZN(n5543) );
  NAND2_X1 U6980 ( .A1(n8337), .A2(n5543), .ZN(n5544) );
  NAND2_X1 U6981 ( .A1(n5546), .A2(n5544), .ZN(n8437) );
  INV_X1 U6982 ( .A(n8437), .ZN(n5545) );
  NAND2_X1 U6983 ( .A1(n8435), .A2(n5546), .ZN(n5563) );
  NAND2_X1 U6984 ( .A1(n5548), .A2(SI_17_), .ZN(n5549) );
  MUX2_X1 U6985 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6889), .Z(n5567) );
  XNOR2_X1 U6986 ( .A(n5567), .B(SI_18_), .ZN(n5564) );
  XNOR2_X1 U6987 ( .A(n5566), .B(n5564), .ZN(n7361) );
  NAND2_X1 U6988 ( .A1(n7361), .A2(n4504), .ZN(n5554) );
  NAND2_X1 U6989 ( .A1(n5551), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5552) );
  XNOR2_X1 U6990 ( .A(n5552), .B(P2_IR_REG_18__SCAN_IN), .ZN(n9320) );
  AOI22_X1 U6991 ( .A1(n5240), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n7009), .B2(
        n9320), .ZN(n5553) );
  XNOR2_X1 U6992 ( .A(n9689), .B(n5661), .ZN(n5583) );
  NAND2_X1 U6993 ( .A1(n5189), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5562) );
  INV_X1 U6994 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9634) );
  OR2_X1 U6995 ( .A1(n7014), .A2(n9634), .ZN(n5561) );
  INV_X1 U6996 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9539) );
  OR2_X1 U6997 ( .A1(n5311), .A2(n9539), .ZN(n5560) );
  INV_X1 U6998 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5555) );
  OAI21_X1 U6999 ( .B1(n5557), .B2(n5556), .A(n5555), .ZN(n5558) );
  NAND2_X1 U7000 ( .A1(n5558), .A2(n5577), .ZN(n9538) );
  OR2_X1 U7001 ( .A1(n5792), .A2(n9538), .ZN(n5559) );
  NOR2_X1 U7002 ( .A1(n9163), .A2(n7521), .ZN(n5584) );
  XNOR2_X1 U7003 ( .A(n5583), .B(n5584), .ZN(n8336) );
  INV_X1 U7004 ( .A(n5564), .ZN(n5565) );
  NAND2_X1 U7005 ( .A1(n5567), .A2(SI_18_), .ZN(n5568) );
  INV_X1 U7006 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n8781) );
  INV_X1 U7007 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7366) );
  MUX2_X1 U7008 ( .A(n8781), .B(n7366), .S(n6889), .Z(n5571) );
  INV_X1 U7009 ( .A(SI_19_), .ZN(n5570) );
  NAND2_X1 U7010 ( .A1(n5571), .A2(n5570), .ZN(n5609) );
  INV_X1 U7011 ( .A(n5571), .ZN(n5572) );
  NAND2_X1 U7012 ( .A1(n5572), .A2(SI_19_), .ZN(n5573) );
  NAND2_X1 U7013 ( .A1(n5609), .A2(n5573), .ZN(n5592) );
  XNOR2_X1 U7014 ( .A(n5591), .B(n5592), .ZN(n7365) );
  NAND2_X1 U7015 ( .A1(n7365), .A2(n4504), .ZN(n5575) );
  AOI22_X1 U7016 ( .A1(n5240), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7009), .B2(
        n9565), .ZN(n5574) );
  XNOR2_X1 U7017 ( .A(n6777), .B(n5576), .ZN(n9168) );
  NAND2_X1 U7018 ( .A1(n5189), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5582) );
  INV_X1 U7019 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n9514) );
  OR2_X1 U7020 ( .A1(n5311), .A2(n9514), .ZN(n5581) );
  INV_X1 U7021 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8681) );
  NAND2_X1 U7022 ( .A1(n5577), .A2(n8681), .ZN(n5578) );
  NAND2_X1 U7023 ( .A1(n5617), .A2(n5578), .ZN(n9513) );
  OR2_X1 U7024 ( .A1(n5792), .A2(n9513), .ZN(n5580) );
  INV_X1 U7025 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9334) );
  OR2_X1 U7026 ( .A1(n7014), .A2(n9334), .ZN(n5579) );
  NOR2_X1 U7027 ( .A1(n8464), .A2(n7521), .ZN(n5588) );
  AND2_X1 U7028 ( .A1(n9168), .A2(n5588), .ZN(n9167) );
  INV_X1 U7029 ( .A(n9167), .ZN(n5586) );
  INV_X1 U7030 ( .A(n5583), .ZN(n5585) );
  NAND2_X1 U7031 ( .A1(n5585), .A2(n5584), .ZN(n9171) );
  AND2_X1 U7032 ( .A1(n5586), .A2(n9171), .ZN(n5587) );
  INV_X1 U7033 ( .A(n9168), .ZN(n5590) );
  INV_X1 U7034 ( .A(n5588), .ZN(n5589) );
  NAND2_X1 U7035 ( .A1(n5590), .A2(n5589), .ZN(n9170) );
  NAND2_X1 U7036 ( .A1(n5612), .A2(n5609), .ZN(n5598) );
  INV_X1 U7037 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7538) );
  INV_X1 U7038 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7555) );
  MUX2_X1 U7039 ( .A(n7538), .B(n7555), .S(n6889), .Z(n5595) );
  INV_X1 U7040 ( .A(SI_20_), .ZN(n5594) );
  NAND2_X1 U7041 ( .A1(n5595), .A2(n5594), .ZN(n5608) );
  INV_X1 U7042 ( .A(n5595), .ZN(n5596) );
  NAND2_X1 U7043 ( .A1(n5596), .A2(SI_20_), .ZN(n5610) );
  AND2_X1 U7044 ( .A1(n5608), .A2(n5610), .ZN(n5597) );
  NAND2_X1 U7045 ( .A1(n7537), .A2(n4504), .ZN(n5600) );
  NAND2_X1 U7046 ( .A1(n5240), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5599) );
  XNOR2_X1 U7047 ( .A(n9503), .B(n5661), .ZN(n5606) );
  NAND2_X1 U7048 ( .A1(n7013), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5604) );
  INV_X1 U7049 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9682) );
  OR2_X1 U7050 ( .A1(n4498), .A2(n9682), .ZN(n5603) );
  INV_X1 U7051 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8467) );
  XNOR2_X1 U7052 ( .A(n5617), .B(n8467), .ZN(n9505) );
  OR2_X1 U7053 ( .A1(n5792), .A2(n9505), .ZN(n5602) );
  INV_X1 U7054 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9623) );
  OR2_X1 U7055 ( .A1(n7014), .A2(n9623), .ZN(n5601) );
  NOR2_X1 U7056 ( .A1(n9180), .A2(n7521), .ZN(n5605) );
  XNOR2_X1 U7057 ( .A(n5606), .B(n5605), .ZN(n8463) );
  NAND2_X1 U7058 ( .A1(n5606), .A2(n5605), .ZN(n5607) );
  MUX2_X1 U7059 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n6889), .Z(n5632) );
  INV_X1 U7060 ( .A(SI_21_), .ZN(n5613) );
  XNOR2_X1 U7061 ( .A(n5632), .B(n5613), .ZN(n5630) );
  XNOR2_X1 U7062 ( .A(n5629), .B(n5630), .ZN(n7568) );
  NAND2_X1 U7063 ( .A1(n7568), .A2(n4504), .ZN(n5615) );
  NAND2_X1 U7064 ( .A1(n5240), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5614) );
  XNOR2_X1 U7065 ( .A(n9486), .B(n5661), .ZN(n5627) );
  INV_X1 U7066 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5616) );
  OAI21_X1 U7067 ( .B1(n5617), .B2(n8467), .A(n5616), .ZN(n5619) );
  AND2_X1 U7068 ( .A1(n5619), .A2(n5618), .ZN(n9487) );
  NAND2_X1 U7069 ( .A1(n5705), .A2(n9487), .ZN(n5624) );
  NAND2_X1 U7070 ( .A1(n6820), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5623) );
  INV_X1 U7071 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n5620) );
  OR2_X1 U7072 ( .A1(n5311), .A2(n5620), .ZN(n5622) );
  INV_X1 U7073 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9678) );
  OR2_X1 U7074 ( .A1(n4498), .A2(n9678), .ZN(n5621) );
  NAND4_X1 U7075 ( .A1(n5624), .A2(n5623), .A3(n5622), .A4(n5621), .ZN(n9260)
         );
  NAND2_X1 U7076 ( .A1(n9260), .A2(n8938), .ZN(n5625) );
  XNOR2_X1 U7077 ( .A(n5627), .B(n5625), .ZN(n9178) );
  INV_X1 U7078 ( .A(n5625), .ZN(n5626) );
  AND2_X1 U7079 ( .A1(n5627), .A2(n5626), .ZN(n5628) );
  NAND2_X1 U7080 ( .A1(n5631), .A2(n5630), .ZN(n5634) );
  NAND2_X1 U7081 ( .A1(n5632), .A2(SI_21_), .ZN(n5633) );
  INV_X1 U7082 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8905) );
  INV_X1 U7083 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7802) );
  MUX2_X1 U7084 ( .A(n8905), .B(n7802), .S(n6889), .Z(n5635) );
  INV_X1 U7085 ( .A(SI_22_), .ZN(n8847) );
  NAND2_X1 U7086 ( .A1(n5635), .A2(n8847), .ZN(n5654) );
  INV_X1 U7087 ( .A(n5635), .ZN(n5636) );
  NAND2_X1 U7088 ( .A1(n5636), .A2(SI_22_), .ZN(n5637) );
  NAND2_X1 U7089 ( .A1(n5654), .A2(n5637), .ZN(n5643) );
  XNOR2_X1 U7090 ( .A(n5644), .B(n5643), .ZN(n7801) );
  NAND2_X1 U7091 ( .A1(n7801), .A2(n4504), .ZN(n5639) );
  NAND2_X1 U7092 ( .A1(n5240), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5638) );
  XNOR2_X1 U7093 ( .A(n9676), .B(n5661), .ZN(n5640) );
  XNOR2_X1 U7094 ( .A(n5641), .B(n5640), .ZN(n9236) );
  AND2_X1 U7095 ( .A1(n5641), .A2(n5640), .ZN(n5642) );
  NAND2_X1 U7096 ( .A1(n5658), .A2(n5654), .ZN(n5650) );
  INV_X1 U7097 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8698) );
  INV_X1 U7098 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5645) );
  MUX2_X1 U7099 ( .A(n8698), .B(n5645), .S(n6889), .Z(n5647) );
  INV_X1 U7100 ( .A(SI_23_), .ZN(n5646) );
  NAND2_X1 U7101 ( .A1(n5647), .A2(n5646), .ZN(n5653) );
  INV_X1 U7102 ( .A(n5647), .ZN(n5648) );
  NAND2_X1 U7103 ( .A1(n5648), .A2(SI_23_), .ZN(n5655) );
  AND2_X1 U7104 ( .A1(n5653), .A2(n5655), .ZN(n5649) );
  NAND2_X1 U7105 ( .A1(n7844), .A2(n4504), .ZN(n5652) );
  NAND2_X1 U7106 ( .A1(n5240), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5651) );
  AND2_X1 U7107 ( .A1(n5654), .A2(n5653), .ZN(n5657) );
  INV_X1 U7108 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8553) );
  INV_X1 U7109 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7950) );
  MUX2_X1 U7110 ( .A(n8553), .B(n7950), .S(n6889), .Z(n5675) );
  XNOR2_X1 U7111 ( .A(n5675), .B(SI_24_), .ZN(n5672) );
  NAND2_X1 U7112 ( .A1(n7949), .A2(n4504), .ZN(n5660) );
  NAND2_X1 U7113 ( .A1(n5240), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5659) );
  XNOR2_X1 U7114 ( .A(n9439), .B(n5661), .ZN(n5670) );
  XNOR2_X1 U7115 ( .A(n5671), .B(n5662), .ZN(n9200) );
  INV_X1 U7116 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n5663) );
  INV_X1 U7117 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9207) );
  OAI21_X1 U7118 ( .B1(n5665), .B2(n5663), .A(n9207), .ZN(n5666) );
  NAND2_X1 U7119 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(P2_REG3_REG_24__SCAN_IN), 
        .ZN(n5664) );
  NAND2_X1 U7120 ( .A1(n5666), .A2(n5685), .ZN(n9203) );
  OR2_X1 U7121 ( .A1(n9203), .A2(n5792), .ZN(n5669) );
  AOI22_X1 U7122 ( .A1(n6820), .A2(P2_REG1_REG_24__SCAN_IN), .B1(n7013), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n5668) );
  INV_X1 U7123 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9666) );
  OR2_X1 U7124 ( .A1(n4498), .A2(n9666), .ZN(n5667) );
  NOR2_X1 U7125 ( .A1(n9155), .A2(n7521), .ZN(n9199) );
  INV_X1 U7126 ( .A(n5672), .ZN(n5673) );
  INV_X1 U7127 ( .A(n5675), .ZN(n5676) );
  NAND2_X1 U7128 ( .A1(n5676), .A2(SI_24_), .ZN(n5677) );
  INV_X1 U7129 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8091) );
  INV_X1 U7130 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8241) );
  MUX2_X1 U7131 ( .A(n8091), .B(n8241), .S(n6889), .Z(n5679) );
  INV_X1 U7132 ( .A(SI_25_), .ZN(n5678) );
  NAND2_X1 U7133 ( .A1(n5679), .A2(n5678), .ZN(n5691) );
  INV_X1 U7134 ( .A(n5679), .ZN(n5680) );
  NAND2_X1 U7135 ( .A1(n5680), .A2(SI_25_), .ZN(n5681) );
  NAND2_X1 U7136 ( .A1(n5691), .A2(n5681), .ZN(n5692) );
  NAND2_X1 U7137 ( .A1(n8090), .A2(n4504), .ZN(n5683) );
  NAND2_X1 U7138 ( .A1(n5240), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5682) );
  XNOR2_X1 U7139 ( .A(n9664), .B(n5661), .ZN(n5690) );
  INV_X1 U7140 ( .A(n5685), .ZN(n5684) );
  NAND2_X1 U7141 ( .A1(n5684), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5700) );
  INV_X1 U7142 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9194) );
  NAND2_X1 U7143 ( .A1(n5685), .A2(n9194), .ZN(n5686) );
  NAND2_X1 U7144 ( .A1(n5700), .A2(n5686), .ZN(n9415) );
  OR2_X1 U7145 ( .A1(n9415), .A2(n5792), .ZN(n5689) );
  AOI22_X1 U7146 ( .A1(n6820), .A2(P2_REG1_REG_25__SCAN_IN), .B1(n7013), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n5688) );
  NAND2_X1 U7147 ( .A1(n5189), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5687) );
  NOR2_X1 U7148 ( .A1(n9244), .A2(n7521), .ZN(n9188) );
  INV_X1 U7149 ( .A(n5690), .ZN(n9189) );
  INV_X1 U7150 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8219) );
  INV_X1 U7151 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8178) );
  MUX2_X1 U7152 ( .A(n8219), .B(n8178), .S(n6889), .Z(n5695) );
  INV_X1 U7153 ( .A(SI_26_), .ZN(n5694) );
  NAND2_X1 U7154 ( .A1(n5695), .A2(n5694), .ZN(n5710) );
  INV_X1 U7155 ( .A(n5695), .ZN(n5696) );
  NAND2_X1 U7156 ( .A1(n5696), .A2(SI_26_), .ZN(n5697) );
  AND2_X1 U7157 ( .A1(n5710), .A2(n5697), .ZN(n5708) );
  NAND2_X1 U7158 ( .A1(n8177), .A2(n4504), .ZN(n5699) );
  NAND2_X1 U7159 ( .A1(n5240), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5698) );
  XNOR2_X1 U7160 ( .A(n9402), .B(n5661), .ZN(n9138) );
  INV_X1 U7161 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9246) );
  NAND2_X1 U7162 ( .A1(n5700), .A2(n9246), .ZN(n5701) );
  INV_X1 U7163 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9592) );
  NAND2_X1 U7164 ( .A1(n5189), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5703) );
  NAND2_X1 U7165 ( .A1(n7013), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5702) );
  OAI211_X1 U7166 ( .C1(n7014), .C2(n9592), .A(n5703), .B(n5702), .ZN(n5704)
         );
  AOI21_X1 U7167 ( .B1(n9408), .B2(n5705), .A(n5704), .ZN(n9391) );
  NOR2_X1 U7168 ( .A1(n9391), .A2(n7521), .ZN(n5706) );
  NAND2_X1 U7169 ( .A1(n9138), .A2(n5706), .ZN(n5707) );
  OAI21_X1 U7170 ( .B1(n9138), .B2(n5706), .A(n5707), .ZN(n9242) );
  INV_X1 U7171 ( .A(n5707), .ZN(n5733) );
  INV_X1 U7172 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8293) );
  INV_X1 U7173 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5712) );
  MUX2_X1 U7174 ( .A(n8293), .B(n5712), .S(n6889), .Z(n5714) );
  INV_X1 U7175 ( .A(SI_27_), .ZN(n5713) );
  NAND2_X1 U7176 ( .A1(n5714), .A2(n5713), .ZN(n5737) );
  INV_X1 U7177 ( .A(n5714), .ZN(n5715) );
  NAND2_X1 U7178 ( .A1(n5715), .A2(SI_27_), .ZN(n5716) );
  AND2_X1 U7179 ( .A1(n5737), .A2(n5716), .ZN(n5735) );
  NAND2_X1 U7180 ( .A1(n8256), .A2(n4504), .ZN(n5718) );
  NAND2_X1 U7181 ( .A1(n5240), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5717) );
  XNOR2_X1 U7182 ( .A(n9393), .B(n5661), .ZN(n5728) );
  INV_X1 U7183 ( .A(n5721), .ZN(n5719) );
  NAND2_X1 U7184 ( .A1(n5719), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5742) );
  INV_X1 U7185 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5720) );
  NAND2_X1 U7186 ( .A1(n5721), .A2(n5720), .ZN(n5722) );
  NAND2_X1 U7187 ( .A1(n5742), .A2(n5722), .ZN(n9143) );
  OR2_X1 U7188 ( .A1(n9143), .A2(n5792), .ZN(n5727) );
  INV_X1 U7189 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9654) );
  NAND2_X1 U7190 ( .A1(n6820), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5724) );
  NAND2_X1 U7191 ( .A1(n7013), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5723) );
  OAI211_X1 U7192 ( .C1(n9654), .C2(n4498), .A(n5724), .B(n5723), .ZN(n5725)
         );
  INV_X1 U7193 ( .A(n5725), .ZN(n5726) );
  NOR2_X1 U7194 ( .A1(n9243), .A2(n7521), .ZN(n5729) );
  NAND2_X1 U7195 ( .A1(n5728), .A2(n5729), .ZN(n5734) );
  INV_X1 U7196 ( .A(n5728), .ZN(n5731) );
  INV_X1 U7197 ( .A(n5729), .ZN(n5730) );
  NAND2_X1 U7198 ( .A1(n5731), .A2(n5730), .ZN(n5732) );
  MUX2_X1 U7199 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n6889), .Z(n5817) );
  INV_X1 U7200 ( .A(SI_28_), .ZN(n5818) );
  XNOR2_X1 U7201 ( .A(n5817), .B(n5818), .ZN(n5815) );
  NAND2_X1 U7202 ( .A1(n8347), .A2(n4504), .ZN(n5740) );
  NAND2_X1 U7203 ( .A1(n5240), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5739) );
  INV_X1 U7204 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5741) );
  NAND2_X1 U7205 ( .A1(n5742), .A2(n5741), .ZN(n5743) );
  NAND2_X1 U7206 ( .A1(n9353), .A2(n5743), .ZN(n9367) );
  OR2_X1 U7207 ( .A1(n9367), .A2(n5792), .ZN(n5748) );
  INV_X1 U7208 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9650) );
  NAND2_X1 U7209 ( .A1(n6820), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5745) );
  NAND2_X1 U7210 ( .A1(n7013), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5744) );
  OAI211_X1 U7211 ( .C1(n9650), .C2(n4498), .A(n5745), .B(n5744), .ZN(n5746)
         );
  INV_X1 U7212 ( .A(n5746), .ZN(n5747) );
  NOR2_X1 U7213 ( .A1(n9145), .A2(n7521), .ZN(n5749) );
  XNOR2_X1 U7214 ( .A(n5749), .B(n5661), .ZN(n5785) );
  INV_X1 U7215 ( .A(n5785), .ZN(n5786) );
  INV_X1 U7216 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5750) );
  NAND2_X1 U7217 ( .A1(n5751), .A2(n5750), .ZN(n5752) );
  NAND2_X1 U7218 ( .A1(n5752), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5779) );
  NAND2_X1 U7219 ( .A1(n5779), .A2(n5778), .ZN(n5753) );
  NAND2_X1 U7220 ( .A1(n5753), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5755) );
  INV_X1 U7221 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5754) );
  NAND2_X1 U7222 ( .A1(n5756), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5757) );
  XNOR2_X1 U7223 ( .A(n5757), .B(P2_IR_REG_26__SCAN_IN), .ZN(n5776) );
  INV_X1 U7224 ( .A(n5776), .ZN(n8220) );
  NAND2_X1 U7225 ( .A1(n7978), .A2(n8220), .ZN(n10458) );
  OR2_X1 U7226 ( .A1(n5758), .A2(n9696), .ZN(n5759) );
  XNOR2_X1 U7227 ( .A(n5759), .B(P2_IR_REG_25__SCAN_IN), .ZN(n5775) );
  INV_X1 U7228 ( .A(n5775), .ZN(n8092) );
  XNOR2_X1 U7229 ( .A(n7978), .B(P2_B_REG_SCAN_IN), .ZN(n5760) );
  NAND2_X1 U7230 ( .A1(n8092), .A2(n5760), .ZN(n5761) );
  INV_X1 U7231 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n5762) );
  NAND2_X1 U7232 ( .A1(n10451), .A2(n5762), .ZN(n5763) );
  INV_X1 U7233 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10463) );
  NOR2_X1 U7234 ( .A1(n5775), .A2(n5776), .ZN(n10464) );
  AOI21_X1 U7235 ( .B1(n10451), .B2(n10463), .A(n10464), .ZN(n6829) );
  NOR4_X1 U7236 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n5767) );
  NOR4_X1 U7237 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n5766) );
  NOR4_X1 U7238 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5765) );
  NOR4_X1 U7239 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n5764) );
  NAND4_X1 U7240 ( .A1(n5767), .A2(n5766), .A3(n5765), .A4(n5764), .ZN(n5773)
         );
  NOR2_X1 U7241 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .ZN(
        n5771) );
  NOR4_X1 U7242 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n5770) );
  NOR4_X1 U7243 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n5769) );
  NOR4_X1 U7244 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n5768) );
  NAND4_X1 U7245 ( .A1(n5771), .A2(n5770), .A3(n5769), .A4(n5768), .ZN(n5772)
         );
  OAI21_X1 U7246 ( .B1(n5773), .B2(n5772), .A(n10451), .ZN(n6828) );
  NAND2_X1 U7247 ( .A1(n6829), .A2(n6828), .ZN(n7376) );
  INV_X1 U7248 ( .A(n7376), .ZN(n5774) );
  NAND2_X1 U7249 ( .A1(n7377), .A2(n5774), .ZN(n5808) );
  NAND2_X1 U7250 ( .A1(n5776), .A2(n5775), .ZN(n5777) );
  XNOR2_X1 U7251 ( .A(n5779), .B(n5778), .ZN(n7008) );
  INV_X1 U7252 ( .A(n8942), .ZN(n9124) );
  AND2_X1 U7253 ( .A1(n10467), .A2(n9124), .ZN(n7391) );
  INV_X1 U7254 ( .A(n7391), .ZN(n5780) );
  OR2_X1 U7255 ( .A1(n10450), .A2(n5780), .ZN(n5807) );
  NAND2_X1 U7256 ( .A1(n9541), .A2(n9565), .ZN(n6827) );
  NOR3_X1 U7257 ( .A1(n9652), .A2(n10593), .A3(n5786), .ZN(n5781) );
  AOI21_X1 U7258 ( .B1(n9652), .B2(n5786), .A(n5781), .ZN(n5782) );
  AND2_X1 U7259 ( .A1(n9131), .A2(n5155), .ZN(n5801) );
  INV_X1 U7260 ( .A(n7678), .ZN(n5784) );
  INV_X1 U7261 ( .A(n5808), .ZN(n5783) );
  NAND2_X1 U7262 ( .A1(n8942), .A2(n9522), .ZN(n5803) );
  OAI21_X1 U7263 ( .B1(n9652), .B2(n9252), .A(n9240), .ZN(n5791) );
  NOR3_X1 U7264 ( .A1(n9652), .A2(n5785), .A3(n10593), .ZN(n5788) );
  NOR2_X1 U7265 ( .A1(n9372), .A2(n5786), .ZN(n5787) );
  OR2_X1 U7266 ( .A1(n9353), .A2(n5792), .ZN(n5798) );
  INV_X1 U7267 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n5795) );
  NAND2_X1 U7268 ( .A1(n6820), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5794) );
  NAND2_X1 U7269 ( .A1(n7013), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5793) );
  OAI211_X1 U7270 ( .C1(n5795), .C2(n4498), .A(n5794), .B(n5793), .ZN(n5796)
         );
  INV_X1 U7271 ( .A(n5796), .ZN(n5797) );
  INV_X1 U7272 ( .A(n5801), .ZN(n7007) );
  INV_X1 U7273 ( .A(n5799), .ZN(n5800) );
  OAI22_X1 U7274 ( .A1(n7185), .A2(n9204), .B1(n9243), .B2(n9390), .ZN(n9362)
         );
  NOR2_X2 U7275 ( .A1(n5808), .A2(n9130), .ZN(n9182) );
  AOI22_X1 U7276 ( .A1(n9362), .A2(n9182), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n5802) );
  INV_X1 U7277 ( .A(n5802), .ZN(n5813) );
  INV_X1 U7278 ( .A(n5803), .ZN(n5804) );
  OAI211_X1 U7279 ( .C1(n5804), .C2(n7007), .A(n7675), .B(n7008), .ZN(n5805)
         );
  AOI21_X1 U7280 ( .B1(n5808), .B2(n10518), .A(n5805), .ZN(n5806) );
  OR2_X1 U7281 ( .A1(n5806), .A2(P2_U3152), .ZN(n5811) );
  INV_X1 U7282 ( .A(n5807), .ZN(n5809) );
  NAND2_X1 U7283 ( .A1(n5809), .A2(n5808), .ZN(n5810) );
  NOR2_X1 U7284 ( .A1(n5813), .A2(n5812), .ZN(n5814) );
  INV_X1 U7285 ( .A(n5817), .ZN(n5819) );
  NAND2_X1 U7286 ( .A1(n5819), .A2(n5818), .ZN(n5820) );
  MUX2_X1 U7287 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n6889), .Z(n6230) );
  INV_X1 U7288 ( .A(SI_29_), .ZN(n6229) );
  XNOR2_X1 U7289 ( .A(n6230), .B(n6229), .ZN(n5821) );
  INV_X1 U7290 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5933) );
  INV_X1 U7291 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5824) );
  INV_X1 U7292 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5823) );
  INV_X1 U7293 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5822) );
  NOR2_X1 U7294 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5826) );
  AND2_X1 U7295 ( .A1(n5826), .A2(n5825), .ZN(n5828) );
  NOR2_X1 U7296 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5827) );
  NAND2_X1 U7297 ( .A1(n6101), .A2(n5831), .ZN(n6137) );
  INV_X1 U7298 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5834) );
  INV_X1 U7299 ( .A(n5840), .ZN(n5836) );
  NAND2_X1 U7300 ( .A1(n5836), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5837) );
  INV_X1 U7301 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5839) );
  NAND2_X1 U7302 ( .A1(n5840), .A2(n5839), .ZN(n5841) );
  INV_X1 U7303 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5845) );
  NAND2_X1 U7304 ( .A1(n5844), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5846) );
  MUX2_X1 U7305 ( .A(n5846), .B(P1_IR_REG_31__SCAN_IN), .S(n5845), .Z(n5847)
         );
  INV_X2 U7306 ( .A(n6177), .ZN(n6117) );
  NAND2_X1 U7307 ( .A1(n8472), .A2(n6117), .ZN(n5849) );
  NAND2_X1 U7308 ( .A1(n6244), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n5848) );
  INV_X1 U7309 ( .A(n5854), .ZN(n8883) );
  INV_X1 U7310 ( .A(n6164), .ZN(n5853) );
  NAND2_X1 U7311 ( .A1(n6106), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5869) );
  NAND2_X1 U7312 ( .A1(n6095), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5868) );
  INV_X1 U7313 ( .A(n6143), .ZN(n5894) );
  NAND2_X1 U7314 ( .A1(n6130), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6120) );
  NAND2_X1 U7315 ( .A1(n6108), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6083) );
  INV_X1 U7316 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7030) );
  INV_X1 U7317 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6051) );
  AND2_X1 U7318 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_12__SCAN_IN), 
        .ZN(n5855) );
  NAND2_X1 U7319 ( .A1(n6038), .A2(n5855), .ZN(n6016) );
  INV_X1 U7320 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n8697) );
  INV_X1 U7321 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5989) );
  NAND2_X1 U7322 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(n5991), .ZN(n5977) );
  NAND2_X1 U7323 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(n5965), .ZN(n5964) );
  INV_X1 U7324 ( .A(n5964), .ZN(n5856) );
  NAND2_X1 U7325 ( .A1(n5856), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5950) );
  INV_X1 U7326 ( .A(n5950), .ZN(n5857) );
  NAND2_X1 U7327 ( .A1(n5857), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5940) );
  INV_X1 U7328 ( .A(n5940), .ZN(n5859) );
  AND2_X1 U7329 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n5858) );
  NAND2_X1 U7330 ( .A1(n5859), .A2(n5858), .ZN(n5916) );
  INV_X1 U7331 ( .A(n5916), .ZN(n5860) );
  NAND2_X1 U7332 ( .A1(n5860), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5906) );
  INV_X1 U7333 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5895) );
  INV_X1 U7334 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8539) );
  INV_X1 U7335 ( .A(n6198), .ZN(n5862) );
  AND2_X1 U7336 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(P1_REG3_REG_25__SCAN_IN), 
        .ZN(n5861) );
  NAND2_X1 U7337 ( .A1(n5862), .A2(n5861), .ZN(n6214) );
  INV_X1 U7338 ( .A(n6214), .ZN(n5863) );
  NAND2_X1 U7339 ( .A1(n5863), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6216) );
  NAND2_X1 U7340 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5864) );
  OR2_X1 U7341 ( .A1(n6216), .A2(n5864), .ZN(n5873) );
  INV_X1 U7342 ( .A(n5873), .ZN(n8865) );
  NAND2_X1 U7343 ( .A1(n6004), .A2(n8865), .ZN(n5867) );
  INV_X1 U7344 ( .A(n5865), .ZN(n8474) );
  NAND2_X1 U7345 ( .A1(n6131), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5866) );
  NAND2_X1 U7346 ( .A1(n8347), .A2(n6117), .ZN(n5871) );
  NAND2_X1 U7347 ( .A1(n6244), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5870) );
  NAND2_X1 U7348 ( .A1(n6095), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5878) );
  NAND2_X1 U7349 ( .A1(n6106), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5877) );
  INV_X1 U7350 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6725) );
  INV_X1 U7351 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5872) );
  OAI21_X1 U7352 ( .B1(n6216), .B2(n6725), .A(n5872), .ZN(n5874) );
  NAND2_X1 U7353 ( .A1(n6004), .A2(n9929), .ZN(n5876) );
  NAND2_X1 U7354 ( .A1(n6131), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5875) );
  AND2_X1 U7355 ( .A1(n6390), .A2(n6380), .ZN(n6441) );
  NAND2_X1 U7356 ( .A1(n7949), .A2(n6117), .ZN(n5880) );
  NAND2_X1 U7357 ( .A1(n6244), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5879) );
  NAND2_X1 U7358 ( .A1(n6095), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5884) );
  NAND2_X1 U7359 ( .A1(n6131), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5883) );
  XNOR2_X1 U7360 ( .A(n6198), .B(P1_REG3_REG_24__SCAN_IN), .ZN(n9993) );
  NAND2_X1 U7361 ( .A1(n6004), .A2(n9993), .ZN(n5882) );
  NAND2_X1 U7362 ( .A1(n6106), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5881) );
  INV_X1 U7363 ( .A(n9973), .ZN(n10007) );
  NAND2_X1 U7364 ( .A1(n9996), .A2(n10007), .ZN(n6193) );
  NAND2_X1 U7365 ( .A1(n7844), .A2(n6117), .ZN(n5886) );
  NAND2_X1 U7366 ( .A1(n6244), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5885) );
  NAND2_X2 U7367 ( .A1(n5886), .A2(n5885), .ZN(n10087) );
  NAND2_X1 U7368 ( .A1(n6106), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5891) );
  NAND2_X1 U7369 ( .A1(n6095), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5890) );
  NAND2_X1 U7370 ( .A1(n5897), .A2(n8539), .ZN(n5887) );
  AND2_X1 U7371 ( .A1(n6198), .A2(n5887), .ZN(n10001) );
  NAND2_X1 U7372 ( .A1(n6004), .A2(n10001), .ZN(n5889) );
  NAND2_X1 U7373 ( .A1(n6131), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5888) );
  NAND4_X1 U7374 ( .A1(n5891), .A2(n5890), .A3(n5889), .A4(n5888), .ZN(n10021)
         );
  INV_X1 U7375 ( .A(n10021), .ZN(n9989) );
  OR2_X1 U7376 ( .A1(n10087), .A2(n9989), .ZN(n8500) );
  NAND2_X1 U7377 ( .A1(n6193), .A2(n8500), .ZN(n6365) );
  NAND2_X1 U7378 ( .A1(n7801), .A2(n6117), .ZN(n5893) );
  NAND2_X1 U7379 ( .A1(n6244), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5892) );
  NAND2_X1 U7380 ( .A1(n6106), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5901) );
  NAND2_X1 U7381 ( .A1(n6095), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5900) );
  NAND2_X1 U7382 ( .A1(n5906), .A2(n5895), .ZN(n5896) );
  AND2_X1 U7383 ( .A1(n5897), .A2(n5896), .ZN(n10016) );
  NAND2_X1 U7384 ( .A1(n6004), .A2(n10016), .ZN(n5899) );
  NAND2_X1 U7385 ( .A1(n6131), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5898) );
  NAND4_X1 U7386 ( .A1(n5901), .A2(n5900), .A3(n5899), .A4(n5898), .ZN(n10037)
         );
  INV_X1 U7387 ( .A(n10037), .ZN(n9728) );
  AND2_X1 U7388 ( .A1(n10092), .A2(n9728), .ZN(n8499) );
  NAND2_X1 U7389 ( .A1(n7568), .A2(n6117), .ZN(n5903) );
  NAND2_X1 U7390 ( .A1(n6244), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5902) );
  NAND2_X1 U7391 ( .A1(n6095), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5910) );
  NAND2_X1 U7392 ( .A1(n6106), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5909) );
  INV_X1 U7393 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5904) );
  NAND2_X1 U7394 ( .A1(n5916), .A2(n5904), .ZN(n5905) );
  AND2_X1 U7395 ( .A1(n5906), .A2(n5905), .ZN(n10030) );
  NAND2_X1 U7396 ( .A1(n6004), .A2(n10030), .ZN(n5908) );
  NAND2_X1 U7397 ( .A1(n6131), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5907) );
  NAND4_X1 U7398 ( .A1(n5910), .A2(n5909), .A3(n5908), .A4(n5907), .ZN(n10057)
         );
  INV_X1 U7399 ( .A(n10057), .ZN(n8482) );
  NAND2_X1 U7400 ( .A1(n10098), .A2(n8482), .ZN(n8497) );
  NOR2_X1 U7401 ( .A1(n8499), .A2(n4755), .ZN(n6353) );
  INV_X1 U7402 ( .A(n6353), .ZN(n6190) );
  OR2_X1 U7403 ( .A1(n10098), .A2(n8482), .ZN(n6355) );
  NAND2_X1 U7404 ( .A1(n7537), .A2(n6117), .ZN(n5912) );
  NAND2_X1 U7405 ( .A1(n6244), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5911) );
  NAND2_X1 U7406 ( .A1(n6095), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5920) );
  NAND2_X1 U7407 ( .A1(n6131), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5919) );
  INV_X1 U7408 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5914) );
  INV_X1 U7409 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5913) );
  OAI21_X1 U7410 ( .B1(n5940), .B2(n5914), .A(n5913), .ZN(n5915) );
  AND2_X1 U7411 ( .A1(n5916), .A2(n5915), .ZN(n10047) );
  NAND2_X1 U7412 ( .A1(n6004), .A2(n10047), .ZN(n5918) );
  NAND2_X1 U7413 ( .A1(n6106), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5917) );
  OR2_X1 U7414 ( .A1(n10102), .A2(n9717), .ZN(n6270) );
  NAND2_X1 U7415 ( .A1(n7365), .A2(n6117), .ZN(n5926) );
  INV_X1 U7416 ( .A(n5921), .ZN(n5922) );
  NAND2_X1 U7417 ( .A1(n5922), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5923) );
  OAI22_X1 U7418 ( .A1(n4502), .A2(n7366), .B1(n7367), .B2(n6844), .ZN(n5924)
         );
  INV_X1 U7419 ( .A(n5924), .ZN(n5925) );
  NAND2_X1 U7420 ( .A1(n6106), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5930) );
  NAND2_X1 U7421 ( .A1(n6095), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5929) );
  XNOR2_X1 U7422 ( .A(n5940), .B(P1_REG3_REG_19__SCAN_IN), .ZN(n9719) );
  NAND2_X1 U7423 ( .A1(n6004), .A2(n9719), .ZN(n5928) );
  NAND2_X1 U7424 ( .A1(n6131), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5927) );
  NAND2_X1 U7425 ( .A1(n10108), .A2(n9789), .ZN(n8494) );
  NAND2_X1 U7426 ( .A1(n7361), .A2(n6117), .ZN(n5937) );
  NOR2_X1 U7427 ( .A1(n5931), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n6114) );
  NAND2_X1 U7428 ( .A1(n6114), .A2(n6115), .ZN(n6061) );
  NOR2_X1 U7429 ( .A1(n6043), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n6045) );
  INV_X1 U7430 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5932) );
  NAND2_X1 U7431 ( .A1(n6045), .A2(n5932), .ZN(n6022) );
  NOR2_X1 U7432 ( .A1(n6010), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5996) );
  NAND2_X1 U7433 ( .A1(n5996), .A2(n5997), .ZN(n5972) );
  OAI21_X1 U7434 ( .B1(n5960), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5945) );
  NAND2_X1 U7435 ( .A1(n5945), .A2(n5933), .ZN(n5934) );
  NAND2_X1 U7436 ( .A1(n5934), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5935) );
  XNOR2_X1 U7437 ( .A(n5935), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9892) );
  AOI22_X1 U7438 ( .A1(n9892), .A2(n6173), .B1(n6244), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n5936) );
  NAND2_X1 U7439 ( .A1(n6106), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5944) );
  NAND2_X1 U7440 ( .A1(n6095), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5943) );
  INV_X1 U7441 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5938) );
  NAND2_X1 U7442 ( .A1(n5950), .A2(n5938), .ZN(n5939) );
  AND2_X1 U7443 ( .A1(n5940), .A2(n5939), .ZN(n9791) );
  NAND2_X1 U7444 ( .A1(n6143), .A2(n9791), .ZN(n5942) );
  NAND2_X1 U7445 ( .A1(n6131), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5941) );
  NAND2_X1 U7446 ( .A1(n10112), .A2(n9745), .ZN(n8454) );
  OR2_X1 U7447 ( .A1(n10112), .A2(n9745), .ZN(n6341) );
  NAND2_X1 U7448 ( .A1(n7228), .A2(n6117), .ZN(n5947) );
  XNOR2_X1 U7449 ( .A(n5945), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9877) );
  AOI22_X1 U7450 ( .A1(n9877), .A2(n6173), .B1(n6244), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n5946) );
  NAND2_X1 U7451 ( .A1(n6095), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5954) );
  NAND2_X1 U7452 ( .A1(n6131), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5953) );
  INV_X1 U7453 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5948) );
  NAND2_X1 U7454 ( .A1(n5964), .A2(n5948), .ZN(n5949) );
  AND2_X1 U7455 ( .A1(n5950), .A2(n5949), .ZN(n9747) );
  NAND2_X1 U7456 ( .A1(n6143), .A2(n9747), .ZN(n5952) );
  NAND2_X1 U7457 ( .A1(n6106), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5951) );
  NAND4_X1 U7458 ( .A1(n5954), .A2(n5953), .A3(n5952), .A4(n5951), .ZN(n9816)
         );
  INV_X1 U7459 ( .A(n9816), .ZN(n8329) );
  OR2_X1 U7460 ( .A1(n10119), .A2(n8329), .ZN(n6271) );
  NAND2_X1 U7461 ( .A1(n6341), .A2(n6271), .ZN(n8455) );
  NAND3_X1 U7462 ( .A1(n8494), .A2(n8454), .A3(n8455), .ZN(n5955) );
  NAND3_X1 U7463 ( .A1(n6270), .A2(n6346), .A3(n5955), .ZN(n5956) );
  NAND2_X1 U7464 ( .A1(n10102), .A2(n9717), .ZN(n8496) );
  NAND2_X1 U7465 ( .A1(n5956), .A2(n8496), .ZN(n5957) );
  AND2_X1 U7466 ( .A1(n6355), .A2(n5957), .ZN(n5958) );
  OAI21_X1 U7467 ( .B1(n6190), .B2(n5958), .A(n8498), .ZN(n5959) );
  NOR2_X1 U7468 ( .A1(n6365), .A2(n5959), .ZN(n6436) );
  AND2_X1 U7469 ( .A1(n10119), .A2(n8329), .ZN(n8407) );
  NAND2_X1 U7470 ( .A1(n7162), .A2(n6117), .ZN(n5963) );
  NAND2_X1 U7471 ( .A1(n5960), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5961) );
  XNOR2_X1 U7472 ( .A(n5961), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9858) );
  AOI22_X1 U7473 ( .A1(n9858), .A2(n6173), .B1(n6244), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n5962) );
  NAND2_X1 U7474 ( .A1(n6095), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5969) );
  NAND2_X1 U7475 ( .A1(n6131), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5968) );
  OAI21_X1 U7476 ( .B1(P1_REG3_REG_16__SCAN_IN), .B2(n5965), .A(n5964), .ZN(
        n8231) );
  INV_X1 U7477 ( .A(n8231), .ZN(n8331) );
  NAND2_X1 U7478 ( .A1(n6143), .A2(n8331), .ZN(n5967) );
  NAND2_X1 U7479 ( .A1(n6106), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5966) );
  INV_X1 U7480 ( .A(n8311), .ZN(n5970) );
  NOR2_X1 U7481 ( .A1(n8407), .A2(n5970), .ZN(n5971) );
  NAND2_X1 U7482 ( .A1(n5971), .A2(n8454), .ZN(n6094) );
  NAND2_X1 U7483 ( .A1(n7160), .A2(n6117), .ZN(n5976) );
  NAND2_X1 U7484 ( .A1(n5972), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5984) );
  NAND2_X1 U7485 ( .A1(n5984), .A2(n5983), .ZN(n5986) );
  NAND2_X1 U7486 ( .A1(n5986), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5973) );
  XNOR2_X1 U7487 ( .A(n5973), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9839) );
  NOR2_X1 U7488 ( .A1(n4502), .A2(n8662), .ZN(n5974) );
  AOI21_X1 U7489 ( .B1(n9839), .B2(n6173), .A(n5974), .ZN(n5975) );
  NAND2_X1 U7490 ( .A1(n6106), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5982) );
  NAND2_X1 U7491 ( .A1(n6095), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5981) );
  OR2_X1 U7492 ( .A1(n5991), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5978) );
  AND2_X1 U7493 ( .A1(n5978), .A2(n5977), .ZN(n8158) );
  NAND2_X1 U7494 ( .A1(n6004), .A2(n8158), .ZN(n5980) );
  NAND2_X1 U7495 ( .A1(n6131), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5979) );
  NAND2_X1 U7496 ( .A1(n6336), .A2(n8223), .ZN(n8312) );
  NAND2_X1 U7497 ( .A1(n7109), .A2(n6117), .ZN(n5988) );
  OR2_X1 U7498 ( .A1(n5984), .A2(n5983), .ZN(n5985) );
  AND2_X1 U7499 ( .A1(n5986), .A2(n5985), .ZN(n8010) );
  AOI22_X1 U7500 ( .A1(n6244), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n8010), .B2(
        n6173), .ZN(n5987) );
  NAND2_X1 U7501 ( .A1(n6106), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5995) );
  NAND2_X1 U7502 ( .A1(n6095), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5994) );
  AND2_X1 U7503 ( .A1(n6003), .A2(n5989), .ZN(n5990) );
  NOR2_X1 U7504 ( .A1(n5991), .A2(n5990), .ZN(n7987) );
  NAND2_X1 U7505 ( .A1(n6004), .A2(n7987), .ZN(n5993) );
  NAND2_X1 U7506 ( .A1(n6131), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5992) );
  NAND4_X1 U7507 ( .A1(n5995), .A2(n5994), .A3(n5993), .A4(n5992), .ZN(n9819)
         );
  INV_X1 U7508 ( .A(n9819), .ZN(n8146) );
  NOR2_X1 U7509 ( .A1(n10129), .A2(n8146), .ZN(n8143) );
  NAND2_X1 U7510 ( .A1(n7085), .A2(n6117), .ZN(n6001) );
  INV_X1 U7511 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6113) );
  OR2_X1 U7512 ( .A1(n5996), .A2(n6113), .ZN(n5998) );
  XNOR2_X1 U7513 ( .A(n5998), .B(n5997), .ZN(n8009) );
  OAI22_X1 U7514 ( .A1(n4502), .A2(n7086), .B1(n8009), .B2(n6844), .ZN(n5999)
         );
  INV_X1 U7515 ( .A(n5999), .ZN(n6000) );
  NAND2_X1 U7516 ( .A1(n6095), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6008) );
  NAND2_X1 U7517 ( .A1(n6131), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6007) );
  NAND2_X1 U7518 ( .A1(n6016), .A2(n8697), .ZN(n6002) );
  AND2_X1 U7519 ( .A1(n6003), .A2(n6002), .ZN(n7851) );
  NAND2_X1 U7520 ( .A1(n6004), .A2(n7851), .ZN(n6006) );
  NAND2_X1 U7521 ( .A1(n6106), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6005) );
  OR2_X1 U7522 ( .A1(n10270), .A2(n7928), .ZN(n6279) );
  INV_X1 U7523 ( .A(n6279), .ZN(n6009) );
  OR2_X1 U7524 ( .A1(n8143), .A2(n6009), .ZN(n6323) );
  NAND2_X1 U7525 ( .A1(n7038), .A2(n6117), .ZN(n6013) );
  NAND2_X1 U7526 ( .A1(n6010), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6011) );
  XNOR2_X1 U7527 ( .A(n6011), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7606) );
  AOI22_X1 U7528 ( .A1(n6244), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6173), .B2(
        n7606), .ZN(n6012) );
  NAND2_X1 U7529 ( .A1(n6095), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6021) );
  NAND2_X1 U7530 ( .A1(n6131), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6020) );
  NAND2_X1 U7531 ( .A1(n6038), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6015) );
  INV_X1 U7532 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6014) );
  NAND2_X1 U7533 ( .A1(n6015), .A2(n6014), .ZN(n6017) );
  AND2_X1 U7534 ( .A1(n6017), .A2(n6016), .ZN(n7822) );
  NAND2_X1 U7535 ( .A1(n6004), .A2(n7822), .ZN(n6019) );
  NAND2_X1 U7536 ( .A1(n6106), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6018) );
  NAND2_X1 U7537 ( .A1(n10132), .A2(n10248), .ZN(n7761) );
  NAND2_X1 U7538 ( .A1(n6992), .A2(n6117), .ZN(n6027) );
  NAND2_X1 U7539 ( .A1(n6022), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6024) );
  XNOR2_X1 U7540 ( .A(n6024), .B(n6023), .ZN(n7422) );
  OAI22_X1 U7541 ( .A1(n4502), .A2(n6993), .B1(n6844), .B2(n7422), .ZN(n6025)
         );
  INV_X1 U7542 ( .A(n6025), .ZN(n6026) );
  INV_X2 U7543 ( .A(n5853), .ZN(n6106) );
  NAND2_X1 U7544 ( .A1(n6106), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6032) );
  NAND2_X1 U7545 ( .A1(n6095), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6031) );
  INV_X1 U7546 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6028) );
  XNOR2_X1 U7547 ( .A(n6038), .B(n6028), .ZN(n10254) );
  NAND2_X1 U7548 ( .A1(n6004), .A2(n10254), .ZN(n6030) );
  NAND2_X1 U7549 ( .A1(n6131), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6029) );
  NAND4_X1 U7550 ( .A1(n6032), .A2(n6031), .A3(n6030), .A4(n6029), .ZN(n9822)
         );
  INV_X1 U7551 ( .A(n9822), .ZN(n7814) );
  NAND2_X1 U7552 ( .A1(n10237), .A2(n7814), .ZN(n6315) );
  NAND2_X1 U7553 ( .A1(n6975), .A2(n6117), .ZN(n6036) );
  OR2_X1 U7554 ( .A1(n6045), .A2(n6113), .ZN(n6033) );
  XNOR2_X1 U7555 ( .A(n6033), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7305) );
  INV_X1 U7556 ( .A(n7305), .ZN(n7299) );
  OAI22_X1 U7557 ( .A1(n4502), .A2(n6976), .B1(n6844), .B2(n7299), .ZN(n6034)
         );
  INV_X1 U7558 ( .A(n6034), .ZN(n6035) );
  NAND2_X1 U7559 ( .A1(n6036), .A2(n6035), .ZN(n7752) );
  NAND2_X1 U7560 ( .A1(n6095), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6042) );
  NAND2_X1 U7561 ( .A1(n6131), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6041) );
  NOR2_X1 U7562 ( .A1(n6053), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6037) );
  NAND2_X1 U7563 ( .A1(n6004), .A2(n5066), .ZN(n6040) );
  NAND2_X1 U7564 ( .A1(n6106), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6039) );
  NAND2_X1 U7565 ( .A1(n7752), .A2(n10339), .ZN(n10242) );
  OR2_X1 U7566 ( .A1(n7752), .A2(n10339), .ZN(n6312) );
  NAND2_X1 U7567 ( .A1(n6930), .A2(n6117), .ZN(n6050) );
  NAND2_X1 U7568 ( .A1(n6043), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6044) );
  MUX2_X1 U7569 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6044), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n6047) );
  INV_X1 U7570 ( .A(n6045), .ZN(n6046) );
  NAND2_X1 U7571 ( .A1(n6047), .A2(n6046), .ZN(n7192) );
  OAI22_X1 U7572 ( .A1(n4502), .A2(n8753), .B1(n6844), .B2(n7192), .ZN(n6048)
         );
  INV_X1 U7573 ( .A(n6048), .ZN(n6049) );
  NAND2_X1 U7574 ( .A1(n6050), .A2(n6049), .ZN(n7547) );
  AND2_X1 U7575 ( .A1(n6069), .A2(n6051), .ZN(n6052) );
  NOR2_X1 U7576 ( .A1(n6053), .A2(n6052), .ZN(n10346) );
  NAND2_X1 U7577 ( .A1(n6004), .A2(n10346), .ZN(n6057) );
  NAND2_X1 U7578 ( .A1(n6095), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6056) );
  NAND2_X1 U7579 ( .A1(n6131), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6055) );
  NAND2_X1 U7580 ( .A1(n6106), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6054) );
  NAND4_X1 U7581 ( .A1(n6057), .A2(n6056), .A3(n6055), .A4(n6054), .ZN(n9824)
         );
  INV_X1 U7582 ( .A(n9824), .ZN(n7321) );
  NAND2_X1 U7583 ( .A1(n7547), .A2(n7321), .ZN(n7403) );
  INV_X1 U7584 ( .A(n7403), .ZN(n6058) );
  NAND2_X1 U7585 ( .A1(n6312), .A2(n6058), .ZN(n6059) );
  AND4_X1 U7586 ( .A1(n7761), .A2(n6315), .A3(n10242), .A4(n6059), .ZN(n6060)
         );
  AND2_X1 U7587 ( .A1(n7924), .A2(n6060), .ZN(n6092) );
  INV_X1 U7588 ( .A(n6092), .ZN(n6077) );
  OR2_X1 U7589 ( .A1(n7547), .A2(n7321), .ZN(n6310) );
  NAND2_X1 U7590 ( .A1(n6913), .A2(n6117), .ZN(n6067) );
  NAND2_X1 U7591 ( .A1(n6061), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6088) );
  INV_X1 U7592 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n6062) );
  NAND2_X1 U7593 ( .A1(n6088), .A2(n6062), .ZN(n6063) );
  NAND2_X1 U7594 ( .A1(n6063), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6064) );
  XNOR2_X1 U7595 ( .A(n6064), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7031) );
  INV_X1 U7596 ( .A(n7031), .ZN(n6923) );
  OAI22_X1 U7597 ( .A1(n4502), .A2(n6921), .B1(n6844), .B2(n6923), .ZN(n6065)
         );
  INV_X1 U7598 ( .A(n6065), .ZN(n6066) );
  NAND2_X1 U7599 ( .A1(n6067), .A2(n6066), .ZN(n10404) );
  NAND2_X1 U7600 ( .A1(n6106), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6073) );
  NAND2_X1 U7601 ( .A1(n6095), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6072) );
  NAND2_X1 U7602 ( .A1(n6083), .A2(n7030), .ZN(n6068) );
  AND2_X1 U7603 ( .A1(n6069), .A2(n6068), .ZN(n7490) );
  NAND2_X1 U7604 ( .A1(n6143), .A2(n7490), .ZN(n6071) );
  NAND2_X1 U7605 ( .A1(n6131), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6070) );
  OR2_X1 U7606 ( .A1(n10404), .A2(n10341), .ZN(n10334) );
  AND2_X1 U7607 ( .A1(n6310), .A2(n10334), .ZN(n7402) );
  AND2_X1 U7608 ( .A1(n6312), .A2(n7402), .ZN(n6076) );
  OR2_X1 U7609 ( .A1(n10132), .A2(n10248), .ZN(n6319) );
  OR2_X1 U7610 ( .A1(n10237), .A2(n7814), .ZN(n7812) );
  NAND2_X1 U7611 ( .A1(n6319), .A2(n7812), .ZN(n6074) );
  NAND2_X1 U7612 ( .A1(n6074), .A2(n7761), .ZN(n7763) );
  INV_X1 U7613 ( .A(n7763), .ZN(n6321) );
  NAND2_X1 U7614 ( .A1(n6321), .A2(n7924), .ZN(n6075) );
  OAI21_X1 U7615 ( .B1(n6077), .B2(n6076), .A(n6075), .ZN(n6078) );
  NAND2_X1 U7616 ( .A1(n10122), .A2(n8226), .ZN(n6332) );
  NAND2_X1 U7617 ( .A1(n10129), .A2(n8146), .ZN(n6324) );
  OAI211_X1 U7618 ( .C1(n6323), .C2(n6078), .A(n6332), .B(n6324), .ZN(n6079)
         );
  INV_X1 U7619 ( .A(n6079), .ZN(n6080) );
  NOR2_X1 U7620 ( .A1(n8312), .A2(n6080), .ZN(n6081) );
  NOR2_X1 U7621 ( .A1(n6094), .A2(n6081), .ZN(n6428) );
  INV_X1 U7622 ( .A(n6332), .ZN(n8221) );
  NAND2_X1 U7623 ( .A1(n10404), .A2(n10341), .ZN(n7400) );
  NAND2_X1 U7624 ( .A1(n6095), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6087) );
  NAND2_X1 U7625 ( .A1(n6131), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6086) );
  OR2_X1 U7626 ( .A1(n6108), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6082) );
  AND2_X1 U7627 ( .A1(n6083), .A2(n6082), .ZN(n7357) );
  NAND2_X1 U7628 ( .A1(n6004), .A2(n7357), .ZN(n6085) );
  NAND2_X1 U7629 ( .A1(n6106), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6084) );
  NAND4_X1 U7630 ( .A1(n6087), .A2(n6086), .A3(n6085), .A4(n6084), .ZN(n9826)
         );
  INV_X1 U7631 ( .A(n9826), .ZN(n7322) );
  NAND2_X1 U7632 ( .A1(n6907), .A2(n6117), .ZN(n6091) );
  INV_X1 U7633 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6927) );
  XNOR2_X1 U7634 ( .A(n6088), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6864) );
  INV_X1 U7635 ( .A(n6864), .ZN(n6982) );
  OAI22_X1 U7636 ( .A1(n4502), .A2(n6927), .B1(n6844), .B2(n6982), .ZN(n6089)
         );
  INV_X1 U7637 ( .A(n6089), .ZN(n6090) );
  INV_X1 U7638 ( .A(n7312), .ZN(n7347) );
  NAND2_X1 U7639 ( .A1(n7322), .A2(n7347), .ZN(n7318) );
  NAND4_X1 U7640 ( .A1(n6324), .A2(n6092), .A3(n7400), .A4(n7318), .ZN(n6093)
         );
  OR3_X1 U7641 ( .A1(n6094), .A2(n8221), .A3(n6093), .ZN(n6431) );
  NAND2_X1 U7642 ( .A1(n6131), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6099) );
  NAND2_X1 U7643 ( .A1(n6095), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6098) );
  NAND2_X1 U7644 ( .A1(n6164), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6097) );
  INV_X1 U7645 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7292) );
  NAND2_X1 U7646 ( .A1(n6143), .A2(n7292), .ZN(n6096) );
  INV_X1 U7647 ( .A(n6100), .ZN(n6916) );
  NAND2_X1 U7648 ( .A1(n6244), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n6105) );
  INV_X1 U7649 ( .A(n6170), .ZN(n6103) );
  INV_X1 U7650 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6102) );
  NAND2_X1 U7651 ( .A1(n6103), .A2(n6102), .ZN(n6171) );
  NAND2_X1 U7652 ( .A1(n6173), .A2(n6915), .ZN(n6104) );
  OAI211_X1 U7653 ( .C1(n6916), .C2(n6177), .A(n6105), .B(n6104), .ZN(n6180)
         );
  NAND2_X1 U7654 ( .A1(n7099), .A2(n10373), .ZN(n6272) );
  NAND2_X1 U7655 ( .A1(n6095), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6112) );
  NAND2_X1 U7656 ( .A1(n6106), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6111) );
  AND2_X1 U7657 ( .A1(n6120), .A2(n8817), .ZN(n6107) );
  NOR2_X1 U7658 ( .A1(n6108), .A2(n6107), .ZN(n7243) );
  NAND2_X1 U7659 ( .A1(n6143), .A2(n7243), .ZN(n6110) );
  NAND2_X1 U7660 ( .A1(n6131), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6109) );
  OR2_X1 U7661 ( .A1(n6114), .A2(n6113), .ZN(n6116) );
  XNOR2_X1 U7662 ( .A(n6116), .B(n6115), .ZN(n6969) );
  NAND2_X1 U7663 ( .A1(n6894), .A2(n6117), .ZN(n6119) );
  NAND2_X1 U7664 ( .A1(n6244), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n6118) );
  OAI211_X1 U7665 ( .C1(n6844), .C2(n6969), .A(n6119), .B(n6118), .ZN(n7244)
         );
  NAND2_X1 U7666 ( .A1(n7258), .A2(n7244), .ZN(n6305) );
  NAND2_X1 U7667 ( .A1(n6106), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6124) );
  NAND2_X1 U7668 ( .A1(n6095), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6123) );
  OAI21_X1 U7669 ( .B1(n6130), .B2(P1_REG3_REG_5__SCAN_IN), .A(n6120), .ZN(
        n7175) );
  INV_X1 U7670 ( .A(n7175), .ZN(n7339) );
  NAND2_X1 U7671 ( .A1(n6143), .A2(n7339), .ZN(n6122) );
  NAND2_X1 U7672 ( .A1(n6131), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6121) );
  NAND2_X1 U7673 ( .A1(n6244), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n6127) );
  NAND2_X1 U7674 ( .A1(n5931), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6125) );
  XNOR2_X1 U7675 ( .A(n6125), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10311) );
  NAND2_X1 U7676 ( .A1(n6173), .A2(n10311), .ZN(n6126) );
  OAI211_X1 U7677 ( .C1(n6925), .C2(n6177), .A(n6127), .B(n6126), .ZN(n7236)
         );
  INV_X1 U7678 ( .A(n7236), .ZN(n7337) );
  NAND2_X1 U7679 ( .A1(n9828), .A2(n7337), .ZN(n6301) );
  INV_X1 U7680 ( .A(n6301), .ZN(n6182) );
  NAND2_X1 U7681 ( .A1(n6305), .A2(n6182), .ZN(n6128) );
  INV_X1 U7682 ( .A(n7258), .ZN(n9827) );
  NAND2_X1 U7683 ( .A1(n9827), .A2(n10391), .ZN(n6302) );
  NAND2_X1 U7684 ( .A1(n6128), .A2(n6302), .ZN(n6421) );
  NAND2_X1 U7685 ( .A1(n6106), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6135) );
  NAND2_X1 U7686 ( .A1(n6095), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6134) );
  NOR2_X1 U7687 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6129) );
  NOR2_X1 U7688 ( .A1(n6130), .A2(n6129), .ZN(n7151) );
  NAND2_X1 U7689 ( .A1(n6004), .A2(n7151), .ZN(n6133) );
  NAND2_X1 U7690 ( .A1(n6131), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6132) );
  INV_X1 U7691 ( .A(n6136), .ZN(n6919) );
  NAND2_X1 U7692 ( .A1(n6244), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n6141) );
  NAND2_X1 U7693 ( .A1(n6137), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6138) );
  MUX2_X1 U7694 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6138), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n6139) );
  AND2_X1 U7695 ( .A1(n5931), .A2(n6139), .ZN(n10293) );
  NAND2_X1 U7696 ( .A1(n6173), .A2(n10293), .ZN(n6140) );
  OAI211_X1 U7697 ( .C1(n6919), .C2(n6177), .A(n6141), .B(n6140), .ZN(n6179)
         );
  INV_X1 U7698 ( .A(n6179), .ZN(n7166) );
  INV_X1 U7699 ( .A(n7126), .ZN(n6142) );
  NOR2_X1 U7700 ( .A1(n6421), .A2(n6142), .ZN(n7250) );
  AND2_X1 U7701 ( .A1(n6272), .A2(n7250), .ZN(n6420) );
  NAND2_X1 U7702 ( .A1(n6162), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U7703 ( .A1(n6163), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6146) );
  NAND2_X1 U7704 ( .A1(n6143), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6145) );
  NAND2_X1 U7705 ( .A1(n6164), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6144) );
  INV_X1 U7706 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6892) );
  INV_X1 U7707 ( .A(n6148), .ZN(n6891) );
  NAND2_X1 U7708 ( .A1(n6173), .A2(n6890), .ZN(n6149) );
  NAND2_X1 U7709 ( .A1(n6143), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6155) );
  NAND2_X1 U7710 ( .A1(n6162), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6154) );
  NAND2_X1 U7711 ( .A1(n6163), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6153) );
  NAND2_X1 U7712 ( .A1(n6164), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6152) );
  INV_X1 U7713 ( .A(SI_0_), .ZN(n6157) );
  INV_X1 U7714 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6156) );
  AND2_X1 U7715 ( .A1(n6159), .A2(n6158), .ZN(n10159) );
  MUX2_X1 U7716 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10159), .S(n6160), .Z(n7205)
         );
  INV_X1 U7717 ( .A(n7222), .ZN(n7225) );
  NAND2_X1 U7718 ( .A1(n4733), .A2(n7225), .ZN(n6161) );
  NAND2_X1 U7719 ( .A1(n6143), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6168) );
  NAND2_X1 U7720 ( .A1(n6162), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6167) );
  NAND2_X1 U7721 ( .A1(n6163), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6166) );
  NAND2_X1 U7722 ( .A1(n6164), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6165) );
  INV_X1 U7723 ( .A(n6169), .ZN(n6910) );
  NAND2_X1 U7724 ( .A1(n6170), .A2(P1_IR_REG_2__SCAN_IN), .ZN(n6172) );
  NAND2_X1 U7725 ( .A1(n6173), .A2(n7052), .ZN(n6176) );
  INV_X1 U7726 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6893) );
  NAND2_X1 U7727 ( .A1(n7285), .A2(n8879), .ZN(n6414) );
  INV_X1 U7728 ( .A(n7285), .ZN(n7076) );
  NAND2_X1 U7729 ( .A1(n7076), .A2(n7272), .ZN(n6415) );
  NAND2_X1 U7730 ( .A1(n6414), .A2(n6415), .ZN(n7090) );
  INV_X1 U7731 ( .A(n7090), .ZN(n7094) );
  NAND2_X1 U7732 ( .A1(n6178), .A2(n6414), .ZN(n7280) );
  NAND2_X1 U7733 ( .A1(n6420), .A2(n7280), .ZN(n6187) );
  NAND2_X1 U7734 ( .A1(n7284), .A2(n6179), .ZN(n7127) );
  NAND2_X1 U7735 ( .A1(n7127), .A2(n6417), .ZN(n6181) );
  NAND2_X1 U7736 ( .A1(n6181), .A2(n7126), .ZN(n6183) );
  NAND2_X1 U7737 ( .A1(n7155), .A2(n7236), .ZN(n6300) );
  AOI21_X1 U7738 ( .B1(n6183), .B2(n6300), .A(n6182), .ZN(n6185) );
  INV_X1 U7739 ( .A(n6305), .ZN(n6184) );
  OAI21_X1 U7740 ( .B1(n6185), .B2(n6184), .A(n6302), .ZN(n6186) );
  NAND2_X1 U7741 ( .A1(n7312), .A2(n9826), .ZN(n6274) );
  INV_X1 U7742 ( .A(n6274), .ZN(n6426) );
  AOI21_X1 U7743 ( .B1(n6187), .B2(n6186), .A(n6426), .ZN(n6188) );
  NOR2_X1 U7744 ( .A1(n6431), .A2(n6188), .ZN(n6191) );
  NAND2_X1 U7745 ( .A1(n8496), .A2(n8494), .ZN(n6189) );
  NOR2_X1 U7746 ( .A1(n6190), .A2(n6189), .ZN(n6433) );
  OAI21_X1 U7747 ( .B1(n6428), .B2(n6191), .A(n6433), .ZN(n6205) );
  AND2_X1 U7748 ( .A1(n10084), .A2(n9973), .ZN(n8501) );
  NAND2_X1 U7749 ( .A1(n10087), .A2(n9989), .ZN(n6269) );
  INV_X1 U7750 ( .A(n6269), .ZN(n6192) );
  OR2_X1 U7751 ( .A1(n8501), .A2(n6192), .ZN(n6360) );
  NAND2_X1 U7752 ( .A1(n6360), .A2(n6193), .ZN(n6204) );
  NAND2_X1 U7753 ( .A1(n8090), .A2(n6117), .ZN(n6195) );
  NAND2_X1 U7754 ( .A1(n6244), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6194) );
  NAND2_X1 U7755 ( .A1(n6095), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6203) );
  NAND2_X1 U7756 ( .A1(n6131), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6202) );
  INV_X1 U7757 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6197) );
  INV_X1 U7758 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6196) );
  OAI21_X1 U7759 ( .B1(n6198), .B2(n6197), .A(n6196), .ZN(n6199) );
  AND2_X1 U7760 ( .A1(n6214), .A2(n6199), .ZN(n9977) );
  NAND2_X1 U7761 ( .A1(n6143), .A2(n9977), .ZN(n6201) );
  NAND2_X1 U7762 ( .A1(n6106), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6200) );
  NAND2_X1 U7763 ( .A1(n10079), .A2(n9990), .ZN(n8502) );
  NAND2_X1 U7764 ( .A1(n6204), .A2(n8502), .ZN(n6434) );
  AOI21_X1 U7765 ( .B1(n6436), .B2(n6205), .A(n6434), .ZN(n6222) );
  NAND2_X1 U7766 ( .A1(n6244), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6206) );
  NAND2_X1 U7767 ( .A1(n6095), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6211) );
  NAND2_X1 U7768 ( .A1(n6131), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6210) );
  XNOR2_X1 U7769 ( .A(n6216), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9940) );
  NAND2_X1 U7770 ( .A1(n6143), .A2(n9940), .ZN(n6209) );
  NAND2_X1 U7771 ( .A1(n6106), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6208) );
  NAND2_X1 U7772 ( .A1(n6244), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6212) );
  NAND2_X1 U7773 ( .A1(n6106), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6220) );
  NAND2_X1 U7774 ( .A1(n6095), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6219) );
  INV_X1 U7775 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9805) );
  NAND2_X1 U7776 ( .A1(n6214), .A2(n9805), .ZN(n6215) );
  AND2_X1 U7777 ( .A1(n6216), .A2(n6215), .ZN(n9956) );
  NAND2_X1 U7778 ( .A1(n6004), .A2(n9956), .ZN(n6218) );
  NAND2_X1 U7779 ( .A1(n6131), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6217) );
  AND2_X1 U7780 ( .A1(n6268), .A2(n9959), .ZN(n8504) );
  NAND2_X1 U7781 ( .A1(n9923), .A2(n8504), .ZN(n6438) );
  NAND2_X1 U7782 ( .A1(n10067), .A2(n9926), .ZN(n6295) );
  NAND2_X1 U7783 ( .A1(n10072), .A2(n9974), .ZN(n6267) );
  INV_X1 U7784 ( .A(n6267), .ZN(n8503) );
  NAND2_X1 U7785 ( .A1(n9923), .A2(n8503), .ZN(n6221) );
  AND3_X1 U7786 ( .A1(n8506), .A2(n6295), .A3(n6221), .ZN(n6408) );
  OAI21_X1 U7787 ( .B1(n6222), .B2(n6438), .A(n6408), .ZN(n6248) );
  NAND2_X1 U7788 ( .A1(n8515), .A2(n9927), .ZN(n6443) );
  INV_X1 U7789 ( .A(n6443), .ZN(n6247) );
  INV_X1 U7790 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n6225) );
  NAND2_X1 U7791 ( .A1(n6095), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6224) );
  NAND2_X1 U7792 ( .A1(n6131), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6223) );
  OAI211_X1 U7793 ( .C1(n5853), .C2(n6225), .A(n6224), .B(n6223), .ZN(n9813)
         );
  NAND2_X1 U7794 ( .A1(n6131), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6228) );
  NAND2_X1 U7795 ( .A1(n6095), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6227) );
  NAND2_X1 U7796 ( .A1(n6106), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6226) );
  NAND3_X1 U7797 ( .A1(n6228), .A2(n6227), .A3(n6226), .ZN(n9909) );
  NAND2_X1 U7798 ( .A1(n6231), .A2(n6230), .ZN(n6235) );
  INV_X1 U7799 ( .A(n6232), .ZN(n6233) );
  INV_X1 U7800 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8884) );
  INV_X1 U7801 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8479) );
  INV_X1 U7802 ( .A(SI_30_), .ZN(n6236) );
  NAND2_X1 U7803 ( .A1(n6237), .A2(n6236), .ZN(n6238) );
  NAND2_X1 U7804 ( .A1(n6239), .A2(n6238), .ZN(n6251) );
  NOR2_X1 U7805 ( .A1(n6237), .A2(n6236), .ZN(n6249) );
  INV_X1 U7806 ( .A(n6238), .ZN(n6241) );
  INV_X1 U7807 ( .A(n6239), .ZN(n6240) );
  NAND2_X1 U7808 ( .A1(n6244), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n6245) );
  AOI211_X1 U7809 ( .C1(n6441), .C2(n6248), .A(n6247), .B(n6397), .ZN(n6265)
         );
  INV_X1 U7810 ( .A(n6249), .ZN(n6250) );
  NAND2_X1 U7811 ( .A1(n6251), .A2(n6250), .ZN(n6254) );
  XNOR2_X1 U7812 ( .A(n6252), .B(SI_31_), .ZN(n6253) );
  MUX2_X1 U7813 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n9694), .S(n6889), .Z(n6255) );
  INV_X1 U7814 ( .A(n9813), .ZN(n6266) );
  NAND2_X1 U7815 ( .A1(n6290), .A2(n9909), .ZN(n6256) );
  NAND2_X1 U7816 ( .A1(n6263), .A2(n6256), .ZN(n6400) );
  INV_X1 U7817 ( .A(n6400), .ZN(n6264) );
  NAND2_X1 U7818 ( .A1(n6257), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6403) );
  INV_X1 U7819 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6258) );
  NAND2_X1 U7820 ( .A1(n6403), .A2(n6258), .ZN(n6259) );
  NAND2_X1 U7821 ( .A1(n6259), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6261) );
  INV_X1 U7822 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6260) );
  OR2_X1 U7823 ( .A1(n6261), .A2(n6260), .ZN(n6262) );
  NAND2_X1 U7824 ( .A1(n6261), .A2(n6260), .ZN(n6294) );
  AND2_X2 U7825 ( .A1(n6262), .A2(n6294), .ZN(n7095) );
  NAND2_X1 U7826 ( .A1(n9906), .A2(n9909), .ZN(n6404) );
  OAI211_X1 U7827 ( .C1(n6265), .C2(n6264), .A(n7095), .B(n6404), .ZN(n6293)
         );
  INV_X1 U7828 ( .A(n6404), .ZN(n6447) );
  AND2_X1 U7829 ( .A1(n9913), .A2(n6266), .ZN(n6442) );
  INV_X1 U7830 ( .A(n9943), .ZN(n8505) );
  INV_X1 U7831 ( .A(n9961), .ZN(n6288) );
  XNOR2_X1 U7832 ( .A(n10084), .B(n9973), .ZN(n9986) );
  NAND2_X1 U7833 ( .A1(n6270), .A2(n8496), .ZN(n10043) );
  NAND2_X1 U7834 ( .A1(n6341), .A2(n8454), .ZN(n8450) );
  INV_X1 U7835 ( .A(n8450), .ZN(n8410) );
  INV_X1 U7836 ( .A(n6271), .ZN(n8409) );
  OR2_X1 U7837 ( .A1(n8409), .A2(n8407), .ZN(n8314) );
  NAND2_X1 U7838 ( .A1(n6319), .A2(n7761), .ZN(n7815) );
  INV_X1 U7839 ( .A(n7815), .ZN(n6278) );
  NAND2_X1 U7840 ( .A1(n7812), .A2(n6315), .ZN(n10244) );
  INV_X1 U7841 ( .A(n10244), .ZN(n6314) );
  NAND2_X1 U7842 ( .A1(n6312), .A2(n10242), .ZN(n7750) );
  INV_X1 U7843 ( .A(n7750), .ZN(n7757) );
  NAND2_X1 U7844 ( .A1(n6417), .A2(n6272), .ZN(n7282) );
  INV_X1 U7845 ( .A(n7282), .ZN(n6297) );
  AND2_X1 U7846 ( .A1(n9831), .A2(n7221), .ZN(n6409) );
  NOR2_X1 U7847 ( .A1(n7214), .A2(n6409), .ZN(n7002) );
  NAND4_X1 U7848 ( .A1(n6297), .A2(n7002), .A3(n7094), .A4(n7215), .ZN(n6273)
         );
  INV_X1 U7849 ( .A(n6300), .ZN(n6422) );
  NAND2_X1 U7850 ( .A1(n6305), .A2(n7127), .ZN(n6423) );
  NOR3_X1 U7851 ( .A1(n6273), .A2(n6422), .A3(n6423), .ZN(n6275) );
  NAND2_X1 U7852 ( .A1(n6274), .A2(n7318), .ZN(n7261) );
  INV_X1 U7853 ( .A(n7261), .ZN(n7252) );
  NAND4_X1 U7854 ( .A1(n6275), .A2(n7320), .A3(n7252), .A4(n7250), .ZN(n6276)
         );
  NAND2_X1 U7855 ( .A1(n6310), .A2(n7403), .ZN(n10336) );
  NOR2_X1 U7856 ( .A1(n6276), .A2(n10336), .ZN(n6277) );
  NAND4_X1 U7857 ( .A1(n6278), .A2(n6314), .A3(n7757), .A4(n6277), .ZN(n6280)
         );
  NOR2_X1 U7858 ( .A1(n6280), .A2(n7917), .ZN(n6281) );
  XNOR2_X1 U7859 ( .A(n10129), .B(n9819), .ZN(n8144) );
  NAND4_X1 U7860 ( .A1(n8229), .A2(n8150), .A3(n6281), .A4(n8144), .ZN(n6282)
         );
  NOR2_X1 U7861 ( .A1(n8314), .A2(n6282), .ZN(n6283) );
  NAND3_X1 U7862 ( .A1(n8480), .A2(n8410), .A3(n6283), .ZN(n6284) );
  NOR2_X1 U7863 ( .A1(n10043), .A2(n6284), .ZN(n6285) );
  XNOR2_X1 U7864 ( .A(n10092), .B(n10037), .ZN(n10019) );
  NAND4_X1 U7865 ( .A1(n10005), .A2(n10035), .A3(n6285), .A4(n10019), .ZN(
        n6286) );
  NOR3_X1 U7866 ( .A1(n9971), .A2(n9986), .A3(n6286), .ZN(n6287) );
  NAND4_X1 U7867 ( .A1(n9922), .A2(n8505), .A3(n6288), .A4(n6287), .ZN(n6289)
         );
  NOR4_X1 U7868 ( .A1(n6447), .A2(n6442), .A3(n8507), .A4(n6289), .ZN(n6291)
         );
  OR2_X1 U7869 ( .A1(n9906), .A2(n9909), .ZN(n6394) );
  AND2_X1 U7870 ( .A1(n6394), .A2(n6290), .ZN(n6449) );
  AOI21_X1 U7871 ( .B1(n6291), .B2(n6449), .A(n7095), .ZN(n6401) );
  INV_X1 U7872 ( .A(n6401), .ZN(n6292) );
  NAND2_X1 U7873 ( .A1(n6293), .A2(n6292), .ZN(n6402) );
  MUX2_X1 U7874 ( .A(n9923), .B(n6295), .S(n6717), .Z(n6296) );
  NAND2_X1 U7875 ( .A1(n6296), .A2(n9922), .ZN(n6385) );
  INV_X1 U7876 ( .A(n6385), .ZN(n6389) );
  INV_X1 U7877 ( .A(n6717), .ZN(n6373) );
  OR2_X1 U7878 ( .A1(n9717), .A2(n6373), .ZN(n6352) );
  NAND2_X1 U7879 ( .A1(n7280), .A2(n6297), .ZN(n6298) );
  NAND2_X1 U7880 ( .A1(n6298), .A2(n6417), .ZN(n7251) );
  NAND2_X1 U7881 ( .A1(n7251), .A2(n7126), .ZN(n6299) );
  NAND2_X1 U7882 ( .A1(n6299), .A2(n7127), .ZN(n7164) );
  AND2_X1 U7883 ( .A1(n6300), .A2(n6301), .ZN(n7169) );
  AOI21_X1 U7884 ( .B1(n7164), .B2(n7169), .A(n6422), .ZN(n7232) );
  AND2_X1 U7885 ( .A1(n6305), .A2(n6302), .ZN(n7239) );
  NAND3_X1 U7886 ( .A1(n6306), .A2(n7252), .A3(n6302), .ZN(n6303) );
  NAND3_X1 U7887 ( .A1(n6303), .A2(n7320), .A3(n7318), .ZN(n6304) );
  NAND2_X1 U7888 ( .A1(n6304), .A2(n7402), .ZN(n6309) );
  OAI21_X1 U7889 ( .B1(n6307), .B2(n4757), .A(n7320), .ZN(n6308) );
  MUX2_X1 U7890 ( .A(n7403), .B(n6310), .S(n6717), .Z(n6311) );
  MUX2_X1 U7891 ( .A(n10242), .B(n6312), .S(n6373), .Z(n6313) );
  NAND2_X1 U7892 ( .A1(n7761), .A2(n6315), .ZN(n6316) );
  NAND2_X1 U7893 ( .A1(n6316), .A2(n6373), .ZN(n6317) );
  NAND2_X1 U7894 ( .A1(n6318), .A2(n6317), .ZN(n6320) );
  NAND2_X1 U7895 ( .A1(n6320), .A2(n6319), .ZN(n6331) );
  OAI21_X1 U7896 ( .B1(n6323), .B2(n6321), .A(n6717), .ZN(n6322) );
  AND3_X1 U7897 ( .A1(n6322), .A2(n7924), .A3(n6324), .ZN(n6330) );
  NAND2_X1 U7898 ( .A1(n6323), .A2(n6324), .ZN(n6327) );
  OAI21_X1 U7899 ( .B1(n8143), .B2(n7924), .A(n6324), .ZN(n6325) );
  INV_X1 U7900 ( .A(n6325), .ZN(n6326) );
  MUX2_X1 U7901 ( .A(n6327), .B(n6326), .S(n6717), .Z(n6328) );
  NAND2_X1 U7902 ( .A1(n6328), .A2(n8150), .ZN(n6329) );
  AOI21_X1 U7903 ( .B1(n6331), .B2(n6330), .A(n6329), .ZN(n6335) );
  NAND2_X1 U7904 ( .A1(n8311), .A2(n6332), .ZN(n6333) );
  MUX2_X1 U7905 ( .A(n6333), .B(n8312), .S(n6717), .Z(n6334) );
  OR2_X1 U7906 ( .A1(n6335), .A2(n6334), .ZN(n6338) );
  MUX2_X1 U7907 ( .A(n6336), .B(n8311), .S(n6717), .Z(n6337) );
  NAND2_X1 U7908 ( .A1(n6338), .A2(n6337), .ZN(n6339) );
  INV_X1 U7909 ( .A(n10119), .ZN(n9750) );
  NAND2_X1 U7910 ( .A1(n6340), .A2(n4550), .ZN(n6345) );
  NAND2_X1 U7911 ( .A1(n6346), .A2(n6341), .ZN(n6343) );
  NAND2_X1 U7912 ( .A1(n8494), .A2(n8454), .ZN(n6342) );
  MUX2_X1 U7913 ( .A(n6343), .B(n6342), .S(n6717), .Z(n6344) );
  INV_X1 U7914 ( .A(n8494), .ZN(n6348) );
  INV_X1 U7915 ( .A(n6346), .ZN(n6347) );
  MUX2_X1 U7916 ( .A(n6348), .B(n6347), .S(n6717), .Z(n6349) );
  INV_X1 U7917 ( .A(n10043), .ZN(n10053) );
  OAI21_X1 U7918 ( .B1(n6350), .B2(n6349), .A(n10053), .ZN(n6351) );
  OAI211_X1 U7919 ( .C1(n10102), .C2(n6352), .A(n6351), .B(n10035), .ZN(n6357)
         );
  NAND2_X1 U7920 ( .A1(n6357), .A2(n6353), .ZN(n6354) );
  NAND2_X1 U7921 ( .A1(n6354), .A2(n8498), .ZN(n6359) );
  INV_X1 U7922 ( .A(n8496), .ZN(n6356) );
  INV_X1 U7923 ( .A(n8499), .ZN(n6358) );
  NOR2_X1 U7924 ( .A1(n6360), .A2(n6365), .ZN(n6361) );
  NAND2_X1 U7925 ( .A1(n10072), .A2(n9959), .ZN(n6363) );
  INV_X1 U7926 ( .A(n9974), .ZN(n9814) );
  NAND2_X1 U7927 ( .A1(n8502), .A2(n9814), .ZN(n6362) );
  MUX2_X1 U7928 ( .A(n6363), .B(n6362), .S(n6717), .Z(n6383) );
  OR2_X1 U7929 ( .A1(n6434), .A2(n6717), .ZN(n6368) );
  INV_X1 U7930 ( .A(n8501), .ZN(n6364) );
  NAND2_X1 U7931 ( .A1(n6365), .A2(n6364), .ZN(n6366) );
  NAND3_X1 U7932 ( .A1(n6366), .A2(n9959), .A3(n6717), .ZN(n6367) );
  NAND2_X1 U7933 ( .A1(n6368), .A2(n6367), .ZN(n6384) );
  MUX2_X1 U7934 ( .A(n9814), .B(n10072), .S(n6373), .Z(n6369) );
  INV_X1 U7935 ( .A(n6369), .ZN(n6370) );
  NAND3_X1 U7936 ( .A1(n6379), .A2(n6384), .A3(n6370), .ZN(n6377) );
  NOR2_X1 U7937 ( .A1(n8502), .A2(n9814), .ZN(n6371) );
  NOR2_X1 U7938 ( .A1(n6371), .A2(n10072), .ZN(n6375) );
  INV_X1 U7939 ( .A(n10072), .ZN(n9958) );
  INV_X1 U7940 ( .A(n9959), .ZN(n6372) );
  AOI21_X1 U7941 ( .B1(n9958), .B2(n6372), .A(n9814), .ZN(n6374) );
  MUX2_X1 U7942 ( .A(n6375), .B(n6374), .S(n6373), .Z(n6376) );
  NAND2_X1 U7943 ( .A1(n6377), .A2(n6376), .ZN(n6378) );
  OAI211_X1 U7944 ( .C1(n6379), .C2(n6383), .A(n6378), .B(n8505), .ZN(n6388)
         );
  INV_X1 U7945 ( .A(n8506), .ZN(n6382) );
  INV_X1 U7946 ( .A(n6380), .ZN(n6381) );
  MUX2_X1 U7947 ( .A(n6382), .B(n6381), .S(n6717), .Z(n6387) );
  NOR3_X1 U7948 ( .A1(n6385), .A2(n6384), .A3(n6383), .ZN(n6386) );
  AOI211_X1 U7949 ( .C1(n6389), .C2(n6388), .A(n6387), .B(n6386), .ZN(n6392)
         );
  MUX2_X1 U7950 ( .A(n6443), .B(n6390), .S(n6717), .Z(n6391) );
  OAI211_X1 U7951 ( .C1(n6392), .C2(n8507), .A(n6391), .B(n6400), .ZN(n6393)
         );
  NAND2_X1 U7952 ( .A1(n6394), .A2(n6717), .ZN(n6395) );
  NAND2_X1 U7953 ( .A1(n6395), .A2(n6397), .ZN(n6396) );
  INV_X1 U7954 ( .A(n7100), .ZN(n7000) );
  XNOR2_X1 U7955 ( .A(n6403), .B(P1_IR_REG_20__SCAN_IN), .ZN(n7140) );
  NAND4_X1 U7956 ( .A1(n6405), .A2(n7095), .A3(n6404), .A4(n7803), .ZN(n6406)
         );
  NAND3_X1 U7957 ( .A1(n6407), .A2(n7140), .A3(n6406), .ZN(n6456) );
  INV_X1 U7958 ( .A(n6408), .ZN(n6440) );
  INV_X1 U7959 ( .A(n6409), .ZN(n6412) );
  NAND2_X1 U7960 ( .A1(n6410), .A2(n7222), .ZN(n6411) );
  NAND3_X1 U7961 ( .A1(n6412), .A2(n7095), .A3(n6411), .ZN(n6413) );
  NAND2_X1 U7962 ( .A1(n6414), .A2(n6413), .ZN(n6416) );
  NAND2_X1 U7963 ( .A1(n6418), .A2(n6417), .ZN(n6419) );
  NAND2_X1 U7964 ( .A1(n6420), .A2(n6419), .ZN(n6427) );
  INV_X1 U7965 ( .A(n6421), .ZN(n6425) );
  OR2_X1 U7966 ( .A1(n6423), .A2(n6422), .ZN(n6424) );
  NAND2_X1 U7967 ( .A1(n6425), .A2(n6424), .ZN(n7254) );
  AOI21_X1 U7968 ( .B1(n6427), .B2(n7254), .A(n6426), .ZN(n6430) );
  INV_X1 U7969 ( .A(n6428), .ZN(n6429) );
  OAI21_X1 U7970 ( .B1(n6431), .B2(n6430), .A(n6429), .ZN(n6432) );
  NAND2_X1 U7971 ( .A1(n6433), .A2(n6432), .ZN(n6435) );
  AOI21_X1 U7972 ( .B1(n6436), .B2(n6435), .A(n6434), .ZN(n6437) );
  NOR2_X1 U7973 ( .A1(n6438), .A2(n6437), .ZN(n6439) );
  NOR2_X1 U7974 ( .A1(n6440), .A2(n6439), .ZN(n6446) );
  INV_X1 U7975 ( .A(n6441), .ZN(n6445) );
  INV_X1 U7976 ( .A(n6442), .ZN(n6444) );
  OAI211_X1 U7977 ( .C1(n6446), .C2(n6445), .A(n6444), .B(n6443), .ZN(n6448)
         );
  AOI21_X1 U7978 ( .B1(n6449), .B2(n6448), .A(n6447), .ZN(n6451) );
  INV_X1 U7979 ( .A(n6451), .ZN(n6450) );
  NAND3_X1 U7980 ( .A1(n6450), .A2(n9902), .A3(n7557), .ZN(n6455) );
  AND2_X1 U7981 ( .A1(n7557), .A2(n7367), .ZN(n6719) );
  NAND2_X1 U7982 ( .A1(n6451), .A2(n6719), .ZN(n6454) );
  NAND2_X1 U7983 ( .A1(n6463), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6453) );
  INV_X1 U7984 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6452) );
  XNOR2_X1 U7985 ( .A(n6453), .B(n6452), .ZN(n6842) );
  OR2_X1 U7986 ( .A1(n6842), .A2(P1_U3084), .ZN(n6469) );
  INV_X1 U7987 ( .A(n6469), .ZN(n7827) );
  NAND4_X1 U7988 ( .A1(n6456), .A2(n6455), .A3(n6454), .A4(n7827), .ZN(n6474)
         );
  NOR2_X1 U7989 ( .A1(n6457), .A2(P1_U3084), .ZN(n9896) );
  NAND2_X1 U7990 ( .A1(n9896), .A2(n4500), .ZN(n6852) );
  INV_X1 U7991 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6462) );
  NAND2_X1 U7992 ( .A1(n6459), .A2(n6462), .ZN(n6461) );
  NAND2_X1 U7993 ( .A1(n6461), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6460) );
  OAI21_X1 U7994 ( .B1(n6459), .B2(n6462), .A(n6461), .ZN(n8244) );
  INV_X1 U7995 ( .A(n6463), .ZN(n6464) );
  NAND2_X1 U7996 ( .A1(n6465), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6467) );
  INV_X1 U7997 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6466) );
  NOR2_X1 U7998 ( .A1(n8244), .A2(n7951), .ZN(n6468) );
  INV_X1 U7999 ( .A(n6478), .ZN(n6481) );
  INV_X1 U8000 ( .A(n6842), .ZN(n6871) );
  NOR4_X1 U8001 ( .A1(n6852), .A2(n6481), .A3(n6871), .A4(n7172), .ZN(n6472)
         );
  OAI21_X1 U8002 ( .B1(n6470), .B2(n6469), .A(P1_B_REG_SCAN_IN), .ZN(n6471) );
  NAND2_X1 U8003 ( .A1(n6474), .A2(n6473), .ZN(P1_U3240) );
  NAND2_X1 U8004 ( .A1(n7095), .A2(n7557), .ZN(n7131) );
  AND2_X1 U8005 ( .A1(n7803), .A2(n6719), .ZN(n6475) );
  OR2_X4 U8006 ( .A1(n6487), .A2(n6475), .ZN(n6678) );
  NAND2_X1 U8007 ( .A1(n9831), .A2(n6476), .ZN(n6480) );
  INV_X1 U8008 ( .A(n7131), .ZN(n6477) );
  AND2_X4 U8009 ( .A1(n6478), .A2(n6477), .ZN(n6736) );
  AOI22_X1 U8010 ( .A1(n7205), .A2(n6736), .B1(n6481), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n6479) );
  NAND2_X1 U8011 ( .A1(n9831), .A2(n6736), .ZN(n6483) );
  AOI22_X1 U8012 ( .A1(n7205), .A2(n6731), .B1(n6481), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n6482) );
  NAND2_X1 U8013 ( .A1(n6483), .A2(n6482), .ZN(n7044) );
  NAND2_X1 U8014 ( .A1(n7045), .A2(n7044), .ZN(n7043) );
  INV_X1 U8015 ( .A(n7044), .ZN(n6485) );
  INV_X1 U8016 ( .A(n7095), .ZN(n7627) );
  OAI22_X1 U8017 ( .A1(n7803), .A2(n9902), .B1(n7627), .B2(n6715), .ZN(n6484)
         );
  NAND2_X2 U8018 ( .A1(n7172), .A2(n6484), .ZN(n7093) );
  NAND2_X4 U8019 ( .A1(n7093), .A2(n7131), .ZN(n7173) );
  NAND2_X1 U8020 ( .A1(n6485), .A2(n7173), .ZN(n6486) );
  OAI21_X1 U8021 ( .B1(n7222), .B2(n6487), .A(n6488), .ZN(n6489) );
  NAND2_X1 U8022 ( .A1(n7068), .A2(n7067), .ZN(n6492) );
  NAND2_X1 U8023 ( .A1(n6410), .A2(n6476), .ZN(n6491) );
  INV_X2 U8024 ( .A(n6736), .ZN(n6732) );
  OR2_X1 U8025 ( .A1(n7222), .A2(n6732), .ZN(n6490) );
  NAND2_X1 U8026 ( .A1(n6491), .A2(n6490), .ZN(n7070) );
  NAND2_X1 U8027 ( .A1(n6492), .A2(n7070), .ZN(n7069) );
  OAI22_X1 U8028 ( .A1(n7285), .A2(n6732), .B1(n7272), .B2(n6487), .ZN(n6495)
         );
  XNOR2_X1 U8029 ( .A(n6495), .B(n6660), .ZN(n6498) );
  OR2_X1 U8030 ( .A1(n7285), .A2(n6678), .ZN(n6497) );
  NAND2_X1 U8031 ( .A1(n8879), .A2(n6736), .ZN(n6496) );
  AND2_X1 U8032 ( .A1(n6497), .A2(n6496), .ZN(n6499) );
  NAND2_X1 U8033 ( .A1(n6498), .A2(n6499), .ZN(n7112) );
  INV_X1 U8034 ( .A(n6498), .ZN(n6501) );
  INV_X1 U8035 ( .A(n6499), .ZN(n6500) );
  NAND2_X1 U8036 ( .A1(n6501), .A2(n6500), .ZN(n6502) );
  AND2_X1 U8037 ( .A1(n7112), .A2(n6502), .ZN(n8874) );
  NAND2_X1 U8038 ( .A1(n8875), .A2(n8874), .ZN(n8873) );
  NAND2_X1 U8039 ( .A1(n8873), .A2(n7112), .ZN(n6511) );
  OAI22_X1 U8040 ( .A1(n8877), .A2(n6732), .B1(n10373), .B2(n6487), .ZN(n6503)
         );
  XNOR2_X1 U8041 ( .A(n6503), .B(n6676), .ZN(n6506) );
  OR2_X1 U8042 ( .A1(n8877), .A2(n6678), .ZN(n6505) );
  NAND2_X1 U8043 ( .A1(n6180), .A2(n6736), .ZN(n6504) );
  AND2_X1 U8044 ( .A1(n6505), .A2(n6504), .ZN(n6507) );
  NAND2_X1 U8045 ( .A1(n6506), .A2(n6507), .ZN(n6512) );
  INV_X1 U8046 ( .A(n6506), .ZN(n6509) );
  INV_X1 U8047 ( .A(n6507), .ZN(n6508) );
  NAND2_X1 U8048 ( .A1(n6509), .A2(n6508), .ZN(n6510) );
  AND2_X1 U8049 ( .A1(n6512), .A2(n6510), .ZN(n7114) );
  NAND2_X1 U8050 ( .A1(n6511), .A2(n7114), .ZN(n7115) );
  NAND2_X1 U8051 ( .A1(n7115), .A2(n6512), .ZN(n7149) );
  OAI22_X1 U8052 ( .A1(n7284), .A2(n6732), .B1(n7166), .B2(n6487), .ZN(n6513)
         );
  XNOR2_X1 U8053 ( .A(n6513), .B(n6676), .ZN(n6518) );
  OR2_X1 U8054 ( .A1(n7284), .A2(n6678), .ZN(n6515) );
  NAND2_X1 U8055 ( .A1(n6179), .A2(n6736), .ZN(n6514) );
  NAND2_X1 U8056 ( .A1(n6515), .A2(n6514), .ZN(n6516) );
  XNOR2_X1 U8057 ( .A(n6518), .B(n6516), .ZN(n7150) );
  NAND2_X1 U8058 ( .A1(n7149), .A2(n7150), .ZN(n7148) );
  INV_X1 U8059 ( .A(n6516), .ZN(n6517) );
  NAND2_X1 U8060 ( .A1(n6518), .A2(n6517), .ZN(n6519) );
  OAI22_X1 U8061 ( .A1(n7155), .A2(n6732), .B1(n7337), .B2(n6487), .ZN(n6520)
         );
  XNOR2_X1 U8062 ( .A(n6520), .B(n6676), .ZN(n6531) );
  OR2_X1 U8063 ( .A1(n7155), .A2(n6678), .ZN(n6522) );
  NAND2_X1 U8064 ( .A1(n7236), .A2(n6736), .ZN(n6521) );
  AND2_X1 U8065 ( .A1(n6522), .A2(n6521), .ZN(n7335) );
  AND2_X1 U8066 ( .A1(n6531), .A2(n7335), .ZN(n6535) );
  OAI22_X1 U8067 ( .A1(n7258), .A2(n6732), .B1(n10391), .B2(n6487), .ZN(n6523)
         );
  XNOR2_X1 U8068 ( .A(n6523), .B(n6676), .ZN(n6526) );
  OR2_X1 U8069 ( .A1(n7258), .A2(n6678), .ZN(n6525) );
  NAND2_X1 U8070 ( .A1(n7244), .A2(n6736), .ZN(n6524) );
  AND2_X1 U8071 ( .A1(n6525), .A2(n6524), .ZN(n6527) );
  NAND2_X1 U8072 ( .A1(n6526), .A2(n6527), .ZN(n7349) );
  INV_X1 U8073 ( .A(n6526), .ZN(n6529) );
  INV_X1 U8074 ( .A(n6527), .ZN(n6528) );
  NAND2_X1 U8075 ( .A1(n6529), .A2(n6528), .ZN(n6530) );
  NAND2_X1 U8076 ( .A1(n7349), .A2(n6530), .ZN(n6880) );
  INV_X1 U8077 ( .A(n6531), .ZN(n6877) );
  INV_X1 U8078 ( .A(n7335), .ZN(n6532) );
  AND2_X1 U8079 ( .A1(n6877), .A2(n6532), .ZN(n6533) );
  NOR2_X1 U8080 ( .A1(n6880), .A2(n6533), .ZN(n6534) );
  NAND2_X1 U8081 ( .A1(n9826), .A2(n6736), .ZN(n6536) );
  OAI21_X1 U8082 ( .B1(n7312), .B2(n6487), .A(n6536), .ZN(n6537) );
  XNOR2_X1 U8083 ( .A(n6537), .B(n6676), .ZN(n6540) );
  OR2_X1 U8084 ( .A1(n7312), .A2(n6732), .ZN(n6539) );
  NAND2_X1 U8085 ( .A1(n9826), .A2(n6476), .ZN(n6538) );
  AND2_X1 U8086 ( .A1(n6539), .A2(n6538), .ZN(n6541) );
  NAND2_X1 U8087 ( .A1(n6540), .A2(n6541), .ZN(n6545) );
  INV_X1 U8088 ( .A(n6540), .ZN(n6543) );
  INV_X1 U8089 ( .A(n6541), .ZN(n6542) );
  NAND2_X1 U8090 ( .A1(n6543), .A2(n6542), .ZN(n6544) );
  AND2_X1 U8091 ( .A1(n6545), .A2(n6544), .ZN(n7350) );
  NAND2_X1 U8092 ( .A1(n10404), .A2(n6736), .ZN(n6547) );
  OR2_X1 U8093 ( .A1(n10341), .A2(n6678), .ZN(n6546) );
  NAND2_X1 U8094 ( .A1(n10404), .A2(n6731), .ZN(n6549) );
  OR2_X1 U8095 ( .A1(n10341), .A2(n6732), .ZN(n6548) );
  NAND2_X1 U8096 ( .A1(n6549), .A2(n6548), .ZN(n6550) );
  XNOR2_X1 U8097 ( .A(n6550), .B(n7173), .ZN(n7487) );
  NAND2_X1 U8098 ( .A1(n7486), .A2(n7487), .ZN(n6551) );
  NAND2_X1 U8099 ( .A1(n6551), .A2(n4508), .ZN(n7543) );
  NAND2_X1 U8100 ( .A1(n7547), .A2(n6731), .ZN(n6553) );
  NAND2_X1 U8101 ( .A1(n9824), .A2(n6736), .ZN(n6552) );
  NAND2_X1 U8102 ( .A1(n6553), .A2(n6552), .ZN(n6554) );
  XNOR2_X1 U8103 ( .A(n6554), .B(n6676), .ZN(n6556) );
  AND2_X1 U8104 ( .A1(n9824), .A2(n6476), .ZN(n6555) );
  AOI21_X1 U8105 ( .B1(n7547), .B2(n6736), .A(n6555), .ZN(n6557) );
  NAND2_X1 U8106 ( .A1(n6556), .A2(n6557), .ZN(n6562) );
  INV_X1 U8107 ( .A(n6556), .ZN(n6559) );
  INV_X1 U8108 ( .A(n6557), .ZN(n6558) );
  NAND2_X1 U8109 ( .A1(n6559), .A2(n6558), .ZN(n6560) );
  NAND2_X1 U8110 ( .A1(n6562), .A2(n6560), .ZN(n7544) );
  INV_X1 U8111 ( .A(n7544), .ZN(n6561) );
  NAND2_X1 U8112 ( .A1(n7752), .A2(n6731), .ZN(n6564) );
  OR2_X1 U8113 ( .A1(n10339), .A2(n6732), .ZN(n6563) );
  NAND2_X1 U8114 ( .A1(n6564), .A2(n6563), .ZN(n6565) );
  XNOR2_X1 U8115 ( .A(n6565), .B(n7173), .ZN(n6571) );
  NOR2_X1 U8116 ( .A1(n10339), .A2(n6678), .ZN(n6566) );
  AOI21_X1 U8117 ( .B1(n7752), .B2(n6736), .A(n6566), .ZN(n6572) );
  XNOR2_X1 U8118 ( .A(n6571), .B(n6572), .ZN(n7638) );
  NAND2_X1 U8119 ( .A1(n10237), .A2(n6731), .ZN(n6568) );
  NAND2_X1 U8120 ( .A1(n9822), .A2(n6736), .ZN(n6567) );
  NAND2_X1 U8121 ( .A1(n6568), .A2(n6567), .ZN(n6569) );
  XNOR2_X1 U8122 ( .A(n6569), .B(n7173), .ZN(n6577) );
  AND2_X1 U8123 ( .A1(n9822), .A2(n6476), .ZN(n6570) );
  AOI21_X1 U8124 ( .B1(n10237), .B2(n6736), .A(n6570), .ZN(n6575) );
  XNOR2_X1 U8125 ( .A(n6577), .B(n6575), .ZN(n7667) );
  INV_X1 U8126 ( .A(n6571), .ZN(n6573) );
  NAND2_X1 U8127 ( .A1(n6573), .A2(n6572), .ZN(n7664) );
  AND2_X1 U8128 ( .A1(n7667), .A2(n7664), .ZN(n6574) );
  INV_X1 U8129 ( .A(n6575), .ZN(n6576) );
  NAND2_X1 U8130 ( .A1(n6577), .A2(n6576), .ZN(n6578) );
  NAND2_X1 U8131 ( .A1(n10132), .A2(n6731), .ZN(n6580) );
  OR2_X1 U8132 ( .A1(n10248), .A2(n6732), .ZN(n6579) );
  NAND2_X1 U8133 ( .A1(n6580), .A2(n6579), .ZN(n6581) );
  XNOR2_X1 U8134 ( .A(n6581), .B(n6676), .ZN(n6584) );
  NOR2_X1 U8135 ( .A1(n10248), .A2(n6678), .ZN(n6582) );
  AOI21_X1 U8136 ( .B1(n10132), .B2(n6736), .A(n6582), .ZN(n6583) );
  NAND2_X1 U8137 ( .A1(n6584), .A2(n6583), .ZN(n7791) );
  OR2_X1 U8138 ( .A1(n6584), .A2(n6583), .ZN(n7792) );
  NAND2_X1 U8139 ( .A1(n10270), .A2(n6731), .ZN(n6586) );
  OR2_X1 U8140 ( .A1(n7928), .A2(n6732), .ZN(n6585) );
  NAND2_X1 U8141 ( .A1(n6586), .A2(n6585), .ZN(n6587) );
  XNOR2_X1 U8142 ( .A(n6587), .B(n7173), .ZN(n7847) );
  NAND2_X1 U8143 ( .A1(n10270), .A2(n6736), .ZN(n6589) );
  OR2_X1 U8144 ( .A1(n7928), .A2(n6678), .ZN(n6588) );
  NAND2_X1 U8145 ( .A1(n6589), .A2(n6588), .ZN(n7848) );
  OAI21_X1 U8146 ( .B1(n7846), .B2(n7847), .A(n7848), .ZN(n6591) );
  NAND2_X1 U8147 ( .A1(n7846), .A2(n7847), .ZN(n6590) );
  NAND2_X1 U8148 ( .A1(n10129), .A2(n6736), .ZN(n6593) );
  NAND2_X1 U8149 ( .A1(n9819), .A2(n6476), .ZN(n6592) );
  NAND2_X1 U8150 ( .A1(n6593), .A2(n6592), .ZN(n7980) );
  NAND2_X1 U8151 ( .A1(n10129), .A2(n6731), .ZN(n6595) );
  NAND2_X1 U8152 ( .A1(n9819), .A2(n6736), .ZN(n6594) );
  NAND2_X1 U8153 ( .A1(n6595), .A2(n6594), .ZN(n6596) );
  XNOR2_X1 U8154 ( .A(n6596), .B(n7173), .ZN(n7979) );
  NAND2_X1 U8155 ( .A1(n10122), .A2(n6731), .ZN(n6598) );
  OR2_X1 U8156 ( .A1(n8226), .A2(n6732), .ZN(n6597) );
  NAND2_X1 U8157 ( .A1(n6598), .A2(n6597), .ZN(n6599) );
  XNOR2_X1 U8158 ( .A(n6599), .B(n6676), .ZN(n8070) );
  NOR2_X1 U8159 ( .A1(n8226), .A2(n6678), .ZN(n6600) );
  AOI21_X1 U8160 ( .B1(n10122), .B2(n6736), .A(n6600), .ZN(n6601) );
  INV_X1 U8161 ( .A(n8070), .ZN(n6602) );
  INV_X1 U8162 ( .A(n6601), .ZN(n8069) );
  NAND2_X1 U8163 ( .A1(n6602), .A2(n8069), .ZN(n6603) );
  NAND2_X1 U8164 ( .A1(n8332), .A2(n6731), .ZN(n6605) );
  OR2_X1 U8165 ( .A1(n8316), .A2(n6732), .ZN(n6604) );
  NAND2_X1 U8166 ( .A1(n6605), .A2(n6604), .ZN(n6606) );
  XNOR2_X1 U8167 ( .A(n6606), .B(n6676), .ZN(n6609) );
  NOR2_X1 U8168 ( .A1(n8316), .A2(n6678), .ZN(n6607) );
  AOI21_X1 U8169 ( .B1(n8332), .B2(n6736), .A(n6607), .ZN(n6608) );
  NAND2_X1 U8170 ( .A1(n6609), .A2(n6608), .ZN(n6612) );
  OR2_X1 U8171 ( .A1(n6609), .A2(n6608), .ZN(n6610) );
  NAND2_X1 U8172 ( .A1(n6612), .A2(n6610), .ZN(n8326) );
  INV_X1 U8173 ( .A(n8326), .ZN(n6611) );
  NAND2_X1 U8174 ( .A1(n8324), .A2(n6612), .ZN(n9741) );
  NAND2_X1 U8175 ( .A1(n10119), .A2(n6731), .ZN(n6614) );
  NAND2_X1 U8176 ( .A1(n9816), .A2(n6736), .ZN(n6613) );
  NAND2_X1 U8177 ( .A1(n6614), .A2(n6613), .ZN(n6615) );
  XNOR2_X1 U8178 ( .A(n6615), .B(n7173), .ZN(n6617) );
  AND2_X1 U8179 ( .A1(n9816), .A2(n6476), .ZN(n6616) );
  AOI21_X1 U8180 ( .B1(n10119), .B2(n6736), .A(n6616), .ZN(n6618) );
  XNOR2_X1 U8181 ( .A(n6617), .B(n6618), .ZN(n9742) );
  INV_X1 U8182 ( .A(n6617), .ZN(n6619) );
  NAND2_X1 U8183 ( .A1(n6619), .A2(n6618), .ZN(n6620) );
  NOR2_X1 U8184 ( .A1(n9745), .A2(n6732), .ZN(n6621) );
  AOI21_X1 U8185 ( .B1(n10112), .B2(n6731), .A(n6621), .ZN(n6622) );
  XNOR2_X1 U8186 ( .A(n6622), .B(n7173), .ZN(n6625) );
  INV_X1 U8187 ( .A(n6625), .ZN(n6623) );
  NOR2_X1 U8188 ( .A1(n9745), .A2(n6678), .ZN(n6624) );
  AOI21_X1 U8189 ( .B1(n10112), .B2(n6736), .A(n6624), .ZN(n9784) );
  NAND2_X1 U8190 ( .A1(n9783), .A2(n9784), .ZN(n9710) );
  NAND2_X1 U8191 ( .A1(n6626), .A2(n6625), .ZN(n9782) );
  NAND2_X1 U8192 ( .A1(n9710), .A2(n9782), .ZN(n6634) );
  NAND2_X1 U8193 ( .A1(n10108), .A2(n6731), .ZN(n6628) );
  OR2_X1 U8194 ( .A1(n9789), .A2(n6732), .ZN(n6627) );
  NAND2_X1 U8195 ( .A1(n6628), .A2(n6627), .ZN(n6629) );
  XNOR2_X1 U8196 ( .A(n6629), .B(n6676), .ZN(n6632) );
  NOR2_X1 U8197 ( .A1(n9789), .A2(n6678), .ZN(n6630) );
  AOI21_X1 U8198 ( .B1(n10108), .B2(n6736), .A(n6630), .ZN(n6631) );
  NAND2_X1 U8199 ( .A1(n6632), .A2(n6631), .ZN(n9761) );
  OR2_X1 U8200 ( .A1(n6632), .A2(n6631), .ZN(n6633) );
  AND2_X1 U8201 ( .A1(n9761), .A2(n6633), .ZN(n9711) );
  NAND2_X1 U8202 ( .A1(n6634), .A2(n9711), .ZN(n9714) );
  NAND2_X1 U8203 ( .A1(n9714), .A2(n9761), .ZN(n6642) );
  NAND2_X1 U8204 ( .A1(n10102), .A2(n6731), .ZN(n6636) );
  OR2_X1 U8205 ( .A1(n9717), .A2(n6732), .ZN(n6635) );
  NAND2_X1 U8206 ( .A1(n6636), .A2(n6635), .ZN(n6637) );
  XNOR2_X1 U8207 ( .A(n6637), .B(n6676), .ZN(n6640) );
  NOR2_X1 U8208 ( .A1(n9717), .A2(n6678), .ZN(n6638) );
  AOI21_X1 U8209 ( .B1(n10102), .B2(n6736), .A(n6638), .ZN(n6639) );
  NAND2_X1 U8210 ( .A1(n6640), .A2(n6639), .ZN(n6643) );
  OR2_X1 U8211 ( .A1(n6640), .A2(n6639), .ZN(n6641) );
  AND2_X1 U8212 ( .A1(n6643), .A2(n6641), .ZN(n9762) );
  NAND2_X1 U8213 ( .A1(n6642), .A2(n9762), .ZN(n9765) );
  NAND2_X1 U8214 ( .A1(n10098), .A2(n6731), .ZN(n6645) );
  NAND2_X1 U8215 ( .A1(n10057), .A2(n6736), .ZN(n6644) );
  NAND2_X1 U8216 ( .A1(n6645), .A2(n6644), .ZN(n6646) );
  XNOR2_X1 U8217 ( .A(n6646), .B(n7173), .ZN(n6648) );
  AND2_X1 U8218 ( .A1(n10057), .A2(n6476), .ZN(n6647) );
  AOI21_X1 U8219 ( .B1(n10098), .B2(n6736), .A(n6647), .ZN(n6649) );
  XNOR2_X1 U8220 ( .A(n6648), .B(n6649), .ZN(n9725) );
  INV_X1 U8221 ( .A(n6648), .ZN(n6650) );
  NAND2_X1 U8222 ( .A1(n6650), .A2(n6649), .ZN(n6651) );
  AND2_X1 U8223 ( .A1(n10037), .A2(n6476), .ZN(n6652) );
  AOI21_X1 U8224 ( .B1(n10092), .B2(n6736), .A(n6652), .ZN(n6656) );
  NAND2_X1 U8225 ( .A1(n10092), .A2(n6731), .ZN(n6654) );
  NAND2_X1 U8226 ( .A1(n10037), .A2(n6736), .ZN(n6653) );
  NAND2_X1 U8227 ( .A1(n6654), .A2(n6653), .ZN(n6655) );
  XNOR2_X1 U8228 ( .A(n6655), .B(n7173), .ZN(n9776) );
  NAND2_X1 U8229 ( .A1(n10087), .A2(n6731), .ZN(n6659) );
  NAND2_X1 U8230 ( .A1(n10021), .A2(n6736), .ZN(n6658) );
  NAND2_X1 U8231 ( .A1(n6659), .A2(n6658), .ZN(n6661) );
  XNOR2_X1 U8232 ( .A(n6661), .B(n6660), .ZN(n6664) );
  NAND2_X1 U8233 ( .A1(n10087), .A2(n6736), .ZN(n6663) );
  NAND2_X1 U8234 ( .A1(n10021), .A2(n6476), .ZN(n6662) );
  NAND2_X1 U8235 ( .A1(n6663), .A2(n6662), .ZN(n9701) );
  OAI22_X1 U8236 ( .A1(n9996), .A2(n6487), .B1(n9973), .B2(n6732), .ZN(n6666)
         );
  XNOR2_X1 U8237 ( .A(n6666), .B(n7173), .ZN(n6668) );
  OAI22_X1 U8238 ( .A1(n9996), .A2(n6732), .B1(n9973), .B2(n6678), .ZN(n6667)
         );
  NAND2_X1 U8239 ( .A1(n6668), .A2(n6667), .ZN(n6669) );
  NAND2_X1 U8240 ( .A1(n10079), .A2(n6731), .ZN(n6672) );
  OR2_X1 U8241 ( .A1(n9990), .A2(n6732), .ZN(n6671) );
  NAND2_X1 U8242 ( .A1(n6672), .A2(n6671), .ZN(n6673) );
  XNOR2_X1 U8243 ( .A(n6673), .B(n7173), .ZN(n6681) );
  OAI22_X1 U8244 ( .A1(n9980), .A2(n6732), .B1(n9990), .B2(n6678), .ZN(n6680)
         );
  XNOR2_X1 U8245 ( .A(n6681), .B(n6680), .ZN(n9733) );
  NAND2_X1 U8246 ( .A1(n10072), .A2(n6731), .ZN(n6675) );
  OR2_X1 U8247 ( .A1(n9974), .A2(n6732), .ZN(n6674) );
  NAND2_X1 U8248 ( .A1(n6675), .A2(n6674), .ZN(n6677) );
  XNOR2_X1 U8249 ( .A(n6677), .B(n6676), .ZN(n6682) );
  NOR2_X1 U8250 ( .A1(n9974), .A2(n6678), .ZN(n6679) );
  AOI21_X1 U8251 ( .B1(n10072), .B2(n6736), .A(n6679), .ZN(n6683) );
  XNOR2_X1 U8252 ( .A(n6682), .B(n6683), .ZN(n9798) );
  NOR2_X1 U8253 ( .A1(n6681), .A2(n6680), .ZN(n9799) );
  INV_X1 U8254 ( .A(n6682), .ZN(n6685) );
  INV_X1 U8255 ( .A(n6683), .ZN(n6684) );
  AOI22_X1 U8256 ( .A1(n10067), .A2(n6731), .B1(n6736), .B2(n9964), .ZN(n6686)
         );
  XNOR2_X1 U8257 ( .A(n6686), .B(n7173), .ZN(n6688) );
  AOI22_X1 U8258 ( .A1(n10067), .A2(n6736), .B1(n6476), .B2(n9964), .ZN(n6687)
         );
  NAND2_X1 U8259 ( .A1(n6688), .A2(n6687), .ZN(n6744) );
  OAI21_X1 U8260 ( .B1(n6688), .B2(n6687), .A(n6744), .ZN(n6689) );
  NAND3_X1 U8261 ( .A1(n8244), .A2(P1_B_REG_SCAN_IN), .A3(n7951), .ZN(n6694)
         );
  INV_X1 U8262 ( .A(n7951), .ZN(n6692) );
  INV_X1 U8263 ( .A(P1_B_REG_SCAN_IN), .ZN(n6691) );
  NAND2_X1 U8264 ( .A1(n6692), .A2(n6691), .ZN(n6693) );
  AND2_X1 U8265 ( .A1(n6694), .A2(n6693), .ZN(n6695) );
  INV_X1 U8266 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6696) );
  NAND2_X1 U8267 ( .A1(n10353), .A2(n6696), .ZN(n6699) );
  INV_X1 U8268 ( .A(n6697), .ZN(n8179) );
  NAND2_X1 U8269 ( .A1(n8179), .A2(n7951), .ZN(n6698) );
  AND2_X1 U8270 ( .A1(n6699), .A2(n6698), .ZN(n7019) );
  AND2_X1 U8271 ( .A1(n6842), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6840) );
  AND2_X1 U8272 ( .A1(n6478), .A2(n6840), .ZN(n10354) );
  AND2_X1 U8273 ( .A1(n7019), .A2(n10354), .ZN(n6896) );
  NOR4_X1 U8274 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6708) );
  NOR4_X1 U8275 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n6707) );
  INV_X1 U8276 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n10359) );
  INV_X1 U8277 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10364) );
  INV_X1 U8278 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10363) );
  INV_X1 U8279 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10360) );
  NAND4_X1 U8280 ( .A1(n10359), .A2(n10364), .A3(n10363), .A4(n10360), .ZN(
        n6705) );
  NOR4_X1 U8281 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6703) );
  NOR4_X1 U8282 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n6702) );
  NOR4_X1 U8283 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6701) );
  NOR4_X1 U8284 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n6700) );
  NAND4_X1 U8285 ( .A1(n6703), .A2(n6702), .A3(n6701), .A4(n6700), .ZN(n6704)
         );
  NOR4_X1 U8286 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n6705), .A4(n6704), .ZN(n6706) );
  NAND3_X1 U8287 ( .A1(n6708), .A2(n6707), .A3(n6706), .ZN(n6709) );
  NAND2_X1 U8288 ( .A1(n10353), .A2(n6709), .ZN(n6999) );
  INV_X1 U8289 ( .A(n6999), .ZN(n6713) );
  INV_X1 U8290 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6710) );
  NAND2_X1 U8291 ( .A1(n10353), .A2(n6710), .ZN(n6712) );
  NAND2_X1 U8292 ( .A1(n8179), .A2(n8244), .ZN(n6711) );
  NAND2_X1 U8293 ( .A1(n6712), .A2(n6711), .ZN(n6997) );
  NOR2_X1 U8294 ( .A1(n6713), .A2(n6997), .ZN(n6714) );
  AND2_X1 U8295 ( .A1(n6896), .A2(n6714), .ZN(n6722) );
  AND2_X1 U8296 ( .A1(n7803), .A2(n7627), .ZN(n7141) );
  NOR2_X1 U8297 ( .A1(n10133), .A2(n7000), .ZN(n6716) );
  INV_X1 U8298 ( .A(n6997), .ZN(n7128) );
  NAND3_X1 U8299 ( .A1(n7128), .A2(n7019), .A3(n6999), .ZN(n6718) );
  NAND2_X1 U8300 ( .A1(n6718), .A2(n6996), .ZN(n6721) );
  OR2_X1 U8301 ( .A1(n7100), .A2(n6719), .ZN(n6998) );
  AND3_X1 U8302 ( .A1(n6478), .A2(n6842), .A3(n6998), .ZN(n6720) );
  NAND2_X1 U8303 ( .A1(n6721), .A2(n6720), .ZN(n7066) );
  AND2_X2 U8304 ( .A1(n7066), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9809) );
  INV_X1 U8305 ( .A(n6722), .ZN(n6729) );
  INV_X1 U8306 ( .A(n7172), .ZN(n7001) );
  NAND2_X1 U8307 ( .A1(n7001), .A2(n4501), .ZN(n6723) );
  OR2_X1 U8308 ( .A1(n6729), .A2(n6723), .ZN(n9806) );
  NOR2_X1 U8309 ( .A1(n9806), .A2(n9945), .ZN(n6727) );
  NAND2_X1 U8310 ( .A1(n4500), .A2(n7001), .ZN(n6724) );
  OR2_X1 U8311 ( .A1(n6729), .A2(n6724), .ZN(n9804) );
  OAI22_X1 U8312 ( .A1(n9804), .A2(n9974), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6725), .ZN(n6726) );
  AOI211_X1 U8313 ( .C1(n9809), .C2(n9940), .A(n6727), .B(n6726), .ZN(n6730)
         );
  INV_X1 U8314 ( .A(n6996), .ZN(n6728) );
  NAND2_X1 U8315 ( .A1(n10354), .A2(n6728), .ZN(n8230) );
  NAND2_X1 U8316 ( .A1(n6729), .A2(n8230), .ZN(n7338) );
  NAND2_X1 U8317 ( .A1(n7338), .A2(n10133), .ZN(n9812) );
  INV_X1 U8318 ( .A(n6741), .ZN(n6739) );
  NAND2_X1 U8319 ( .A1(n10065), .A2(n6731), .ZN(n6734) );
  OR2_X1 U8320 ( .A1(n9945), .A2(n6732), .ZN(n6733) );
  NAND2_X1 U8321 ( .A1(n6734), .A2(n6733), .ZN(n6735) );
  XNOR2_X1 U8322 ( .A(n6735), .B(n7173), .ZN(n6738) );
  AOI22_X1 U8323 ( .A1(n10065), .A2(n6736), .B1(n6476), .B2(n8490), .ZN(n6737)
         );
  XNOR2_X1 U8324 ( .A(n6738), .B(n6737), .ZN(n6740) );
  INV_X1 U8325 ( .A(n6740), .ZN(n6745) );
  NAND2_X1 U8326 ( .A1(n6739), .A2(n4549), .ZN(n6750) );
  NAND3_X1 U8327 ( .A1(n6741), .A2(n6740), .A3(n9802), .ZN(n6749) );
  INV_X1 U8328 ( .A(n9812), .ZN(n9792) );
  INV_X1 U8329 ( .A(n9804), .ZN(n9786) );
  AOI22_X1 U8330 ( .A1(n9786), .A2(n9964), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n6743) );
  NAND2_X1 U8331 ( .A1(n9809), .A2(n9929), .ZN(n6742) );
  OAI211_X1 U8332 ( .C1(n9927), .C2(n9806), .A(n6743), .B(n6742), .ZN(n6747)
         );
  INV_X1 U8333 ( .A(n9802), .ZN(n9795) );
  NOR3_X1 U8334 ( .A1(n6745), .A2(n9795), .A3(n6744), .ZN(n6746) );
  AOI211_X1 U8335 ( .C1(n9792), .C2(n10065), .A(n6747), .B(n6746), .ZN(n6748)
         );
  NAND3_X1 U8336 ( .A1(n6750), .A2(n6749), .A3(n6748), .ZN(P1_U3218) );
  INV_X1 U8337 ( .A(n8464), .ZN(n9262) );
  INV_X1 U8338 ( .A(n8341), .ZN(n9264) );
  INV_X1 U8339 ( .A(n8303), .ZN(n9266) );
  NAND2_X1 U8340 ( .A1(n9279), .A2(n7457), .ZN(n9007) );
  NAND2_X2 U8341 ( .A1(n9008), .A2(n9007), .ZN(n8939) );
  NAND2_X1 U8342 ( .A1(n8939), .A2(n7452), .ZN(n6753) );
  INV_X1 U8343 ( .A(n9279), .ZN(n6751) );
  NAND2_X1 U8344 ( .A1(n6751), .A2(n7457), .ZN(n6752) );
  NAND2_X1 U8345 ( .A1(n6753), .A2(n6752), .ZN(n7464) );
  OR2_X2 U8346 ( .A1(n9278), .A2(n10482), .ZN(n9009) );
  NAND2_X1 U8347 ( .A1(n9278), .A2(n10482), .ZN(n9011) );
  NAND2_X1 U8348 ( .A1(n7464), .A2(n8941), .ZN(n6755) );
  INV_X1 U8349 ( .A(n10482), .ZN(n7588) );
  OR2_X1 U8350 ( .A1(n9278), .A2(n7588), .ZN(n6754) );
  NAND2_X1 U8351 ( .A1(n6755), .A2(n6754), .ZN(n7380) );
  OR2_X1 U8352 ( .A1(n9277), .A2(n10489), .ZN(n8996) );
  NAND2_X1 U8353 ( .A1(n9277), .A2(n10489), .ZN(n8988) );
  NAND2_X1 U8354 ( .A1(n7380), .A2(n8943), .ZN(n6757) );
  INV_X1 U8355 ( .A(n9277), .ZN(n7592) );
  NAND2_X1 U8356 ( .A1(n7592), .A2(n10489), .ZN(n6756) );
  NAND2_X1 U8357 ( .A1(n6757), .A2(n6756), .ZN(n7438) );
  NAND2_X1 U8358 ( .A1(n9275), .A2(n7524), .ZN(n6758) );
  AND2_X1 U8359 ( .A1(n8940), .A2(n6758), .ZN(n6763) );
  INV_X1 U8360 ( .A(n6758), .ZN(n6762) );
  NOR2_X1 U8361 ( .A1(n9275), .A2(n7524), .ZN(n6760) );
  OR2_X1 U8362 ( .A1(n9276), .A2(n9214), .ZN(n7439) );
  INV_X1 U8363 ( .A(n7439), .ZN(n6759) );
  NAND2_X1 U8364 ( .A1(n9274), .A2(n10501), .ZN(n9014) );
  NAND2_X1 U8365 ( .A1(n9273), .A2(n7633), .ZN(n9019) );
  NAND2_X1 U8366 ( .A1(n9018), .A2(n9019), .ZN(n9016) );
  NAND2_X1 U8367 ( .A1(n7507), .A2(n9016), .ZN(n7506) );
  INV_X1 U8368 ( .A(n7633), .ZN(n7651) );
  OR2_X1 U8369 ( .A1(n9273), .A2(n7651), .ZN(n6764) );
  XNOR2_X2 U8370 ( .A(n9272), .B(n10505), .ZN(n9021) );
  NOR2_X1 U8371 ( .A1(n7733), .A2(n9021), .ZN(n6768) );
  OR2_X1 U8372 ( .A1(n8898), .A2(n7808), .ZN(n9033) );
  NAND2_X1 U8373 ( .A1(n8898), .A2(n7808), .ZN(n9028) );
  INV_X1 U8374 ( .A(n8895), .ZN(n9270) );
  AND2_X1 U8375 ( .A1(n8040), .A2(n9270), .ZN(n6769) );
  OR2_X1 U8376 ( .A1(n8951), .A2(n6769), .ZN(n7906) );
  INV_X1 U8377 ( .A(n7992), .ZN(n9269) );
  AND2_X1 U8378 ( .A1(n7957), .A2(n9269), .ZN(n6770) );
  OR2_X1 U8379 ( .A1(n7906), .A2(n6770), .ZN(n7962) );
  NAND2_X1 U8380 ( .A1(n6765), .A2(n8051), .ZN(n9045) );
  NOR2_X1 U8381 ( .A1(n7962), .A2(n8956), .ZN(n6766) );
  NAND2_X1 U8382 ( .A1(n9272), .A2(n10505), .ZN(n7894) );
  NAND2_X1 U8383 ( .A1(n6766), .A2(n7894), .ZN(n6767) );
  NOR2_X1 U8384 ( .A1(n6768), .A2(n6767), .ZN(n6774) );
  NAND2_X1 U8385 ( .A1(n8040), .A2(n8895), .ZN(n9031) );
  NAND2_X1 U8386 ( .A1(n9032), .A2(n9031), .ZN(n8025) );
  INV_X1 U8387 ( .A(n7808), .ZN(n9271) );
  OR2_X1 U8388 ( .A1(n8898), .A2(n9271), .ZN(n8021) );
  INV_X1 U8389 ( .A(n8051), .ZN(n9268) );
  OR2_X1 U8390 ( .A1(n6765), .A2(n9268), .ZN(n6771) );
  NAND2_X1 U8391 ( .A1(n6772), .A2(n6771), .ZN(n6773) );
  XNOR2_X1 U8392 ( .A(n10220), .B(n9049), .ZN(n9055) );
  NAND2_X1 U8393 ( .A1(n8917), .A2(n8249), .ZN(n9057) );
  INV_X1 U8394 ( .A(n8249), .ZN(n9267) );
  NAND2_X1 U8395 ( .A1(n8361), .A2(n8303), .ZN(n9060) );
  NAND2_X1 U8396 ( .A1(n9061), .A2(n9060), .ZN(n8351) );
  NAND2_X1 U8397 ( .A1(n8352), .A2(n8351), .ZN(n8350) );
  OAI21_X1 U8398 ( .B1(n9266), .B2(n8361), .A(n8350), .ZN(n8423) );
  XNOR2_X1 U8399 ( .A(n9066), .B(n9265), .ZN(n9063) );
  NAND2_X1 U8400 ( .A1(n9559), .A2(n8341), .ZN(n9071) );
  NAND2_X1 U8401 ( .A1(n9527), .A2(n9071), .ZN(n9554) );
  INV_X1 U8402 ( .A(n9163), .ZN(n9263) );
  OAI21_X1 U8403 ( .B1(n6777), .B2(n8464), .A(n9512), .ZN(n6778) );
  NAND2_X1 U8404 ( .A1(n9503), .A2(n9180), .ZN(n9085) );
  INV_X1 U8405 ( .A(n9180), .ZN(n9261) );
  NOR2_X1 U8406 ( .A1(n9486), .A2(n9260), .ZN(n6779) );
  INV_X1 U8407 ( .A(n9486), .ZN(n9680) );
  INV_X1 U8408 ( .A(n9260), .ZN(n6809) );
  NAND2_X1 U8409 ( .A1(n9468), .A2(n9181), .ZN(n8983) );
  NOR2_X1 U8410 ( .A1(n9451), .A2(n9452), .ZN(n9450) );
  INV_X1 U8411 ( .A(n9258), .ZN(n9091) );
  NOR2_X1 U8412 ( .A1(n9672), .A2(n9091), .ZN(n6780) );
  NAND2_X1 U8413 ( .A1(n9439), .A2(n9155), .ZN(n9096) );
  INV_X1 U8414 ( .A(n9155), .ZN(n9257) );
  NAND2_X1 U8415 ( .A1(n9427), .A2(n9244), .ZN(n8975) );
  NAND2_X1 U8416 ( .A1(n9426), .A2(n9425), .ZN(n9424) );
  NAND2_X1 U8417 ( .A1(n9664), .A2(n9244), .ZN(n6782) );
  NAND2_X1 U8418 ( .A1(n9402), .A2(n9391), .ZN(n9380) );
  NAND2_X1 U8419 ( .A1(n9660), .A2(n9391), .ZN(n6783) );
  NAND2_X1 U8420 ( .A1(n9656), .A2(n9243), .ZN(n6784) );
  NAND2_X1 U8421 ( .A1(n9372), .A2(n9145), .ZN(n6785) );
  NAND2_X1 U8422 ( .A1(n9366), .A2(n9365), .ZN(n9364) );
  NAND2_X1 U8423 ( .A1(n9652), .A2(n9145), .ZN(n6786) );
  NAND2_X1 U8424 ( .A1(n9364), .A2(n6786), .ZN(n6789) );
  NAND2_X1 U8425 ( .A1(n8472), .A2(n4504), .ZN(n6788) );
  NAND2_X1 U8426 ( .A1(n5240), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6787) );
  NAND2_X1 U8427 ( .A1(n6834), .A2(n7185), .ZN(n9113) );
  XNOR2_X1 U8428 ( .A(n6789), .B(n8921), .ZN(n9351) );
  XNOR2_X1 U8429 ( .A(n9131), .B(n7389), .ZN(n9562) );
  NAND2_X1 U8430 ( .A1(n9562), .A2(n9522), .ZN(n8260) );
  AND2_X1 U8431 ( .A1(n8942), .A2(n9565), .ZN(n6790) );
  NAND2_X1 U8432 ( .A1(n8902), .A2(n6790), .ZN(n8272) );
  NAND2_X1 U8433 ( .A1(n8260), .A2(n8272), .ZN(n10524) );
  NAND2_X1 U8434 ( .A1(n9351), .A2(n10524), .ZN(n6826) );
  NAND2_X1 U8435 ( .A1(n9008), .A2(n7498), .ZN(n8993) );
  AND2_X1 U8436 ( .A1(n8993), .A2(n9007), .ZN(n7466) );
  NAND2_X1 U8437 ( .A1(n7465), .A2(n9009), .ZN(n6791) );
  INV_X1 U8438 ( .A(n8943), .ZN(n8999) );
  NAND2_X1 U8439 ( .A1(n6791), .A2(n8999), .ZN(n7383) );
  OR2_X1 U8440 ( .A1(n9275), .A2(n7539), .ZN(n9001) );
  AND2_X1 U8441 ( .A1(n8997), .A2(n9001), .ZN(n6792) );
  INV_X1 U8442 ( .A(n9001), .ZN(n6793) );
  OR2_X1 U8443 ( .A1(n6793), .A2(n8989), .ZN(n7508) );
  AND2_X1 U8444 ( .A1(n8945), .A2(n9019), .ZN(n7735) );
  NAND2_X1 U8445 ( .A1(n7509), .A2(n6795), .ZN(n6801) );
  INV_X1 U8446 ( .A(n9272), .ZN(n9023) );
  INV_X1 U8447 ( .A(n9021), .ZN(n6798) );
  INV_X1 U8448 ( .A(n9019), .ZN(n6797) );
  AND2_X1 U8449 ( .A1(n9017), .A2(n9018), .ZN(n6796) );
  OR2_X1 U8450 ( .A1(n6797), .A2(n6796), .ZN(n7737) );
  NOR2_X1 U8451 ( .A1(n5069), .A2(n6799), .ZN(n6800) );
  NAND2_X1 U8452 ( .A1(n6801), .A2(n6800), .ZN(n7897) );
  NAND2_X1 U8453 ( .A1(n7897), .A2(n9033), .ZN(n6802) );
  NAND2_X1 U8454 ( .A1(n6802), .A2(n9028), .ZN(n8028) );
  INV_X1 U8455 ( .A(n8025), .ZN(n8950) );
  NAND2_X1 U8456 ( .A1(n8028), .A2(n8950), .ZN(n8027) );
  NAND2_X1 U8457 ( .A1(n8027), .A2(n9031), .ZN(n7910) );
  INV_X1 U8458 ( .A(n8956), .ZN(n6803) );
  NAND2_X1 U8459 ( .A1(n7967), .A2(n9043), .ZN(n8261) );
  NAND2_X1 U8460 ( .A1(n10220), .A2(n9049), .ZN(n6804) );
  NAND2_X1 U8461 ( .A1(n8165), .A2(n9056), .ZN(n8354) );
  INV_X1 U8462 ( .A(n8351), .ZN(n9059) );
  INV_X1 U8463 ( .A(n9063), .ZN(n8958) );
  INV_X1 U8464 ( .A(n9265), .ZN(n9065) );
  INV_X1 U8465 ( .A(n9555), .ZN(n6806) );
  INV_X1 U8466 ( .A(n9554), .ZN(n6805) );
  OR2_X1 U8467 ( .A1(n9545), .A2(n9163), .ZN(n9075) );
  NAND2_X1 U8468 ( .A1(n9545), .A2(n9163), .ZN(n9078) );
  NAND2_X1 U8469 ( .A1(n9075), .A2(n9078), .ZN(n9535) );
  INV_X1 U8470 ( .A(n9527), .ZN(n6807) );
  NOR2_X1 U8471 ( .A1(n9535), .A2(n6807), .ZN(n6808) );
  OR2_X1 U8472 ( .A1(n9626), .A2(n8464), .ZN(n9076) );
  NAND2_X1 U8473 ( .A1(n9626), .A2(n8464), .ZN(n9080) );
  INV_X1 U8474 ( .A(n9495), .ZN(n9497) );
  OR2_X1 U8475 ( .A1(n9486), .A2(n6809), .ZN(n8979) );
  NAND2_X1 U8476 ( .A1(n9486), .A2(n6809), .ZN(n8981) );
  NAND2_X1 U8477 ( .A1(n8979), .A2(n8981), .ZN(n9479) );
  INV_X1 U8478 ( .A(n9478), .ZN(n9077) );
  NOR2_X1 U8479 ( .A1(n9479), .A2(n9077), .ZN(n6810) );
  NAND2_X1 U8480 ( .A1(n9460), .A2(n9463), .ZN(n9459) );
  AND2_X1 U8481 ( .A1(n9432), .A2(n8975), .ZN(n6811) );
  INV_X1 U8482 ( .A(n8975), .ZN(n6813) );
  AND2_X1 U8483 ( .A1(n9417), .A2(n8976), .ZN(n6812) );
  INV_X1 U8484 ( .A(n9382), .ZN(n9099) );
  AND2_X1 U8485 ( .A1(n9380), .A2(n9099), .ZN(n6816) );
  NAND2_X1 U8486 ( .A1(n9379), .A2(n6816), .ZN(n9378) );
  OR2_X1 U8487 ( .A1(n9393), .A2(n9243), .ZN(n9105) );
  OR2_X1 U8488 ( .A1(n9382), .A2(n9381), .ZN(n9377) );
  AND2_X1 U8489 ( .A1(n9105), .A2(n9377), .ZN(n6817) );
  NAND2_X1 U8490 ( .A1(n9378), .A2(n6817), .ZN(n9361) );
  INV_X1 U8491 ( .A(n9365), .ZN(n6818) );
  INV_X1 U8492 ( .A(n9106), .ZN(n9102) );
  XNOR2_X1 U8493 ( .A(n8922), .B(n8921), .ZN(n6824) );
  NAND2_X1 U8494 ( .A1(n5155), .A2(n9124), .ZN(n8937) );
  AND2_X1 U8495 ( .A1(n8967), .A2(n8937), .ZN(n9553) );
  INV_X1 U8496 ( .A(n9145), .ZN(n9387) );
  INV_X1 U8497 ( .A(P2_B_REG_SCAN_IN), .ZN(n8756) );
  NOR2_X1 U8498 ( .A1(n9129), .A2(n8756), .ZN(n6819) );
  NOR2_X1 U8499 ( .A1(n9204), .A2(n6819), .ZN(n9342) );
  INV_X1 U8500 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8691) );
  NAND2_X1 U8501 ( .A1(n7013), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6822) );
  NAND2_X1 U8502 ( .A1(n6820), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6821) );
  OAI211_X1 U8503 ( .C1(n4498), .C2(n8691), .A(n6822), .B(n6821), .ZN(n9253)
         );
  AOI22_X1 U8504 ( .A1(n9387), .A2(n9245), .B1(n9342), .B2(n9253), .ZN(n6823)
         );
  NAND2_X1 U8505 ( .A1(n7472), .A2(n10489), .ZN(n7618) );
  INV_X1 U8506 ( .A(n8040), .ZN(n10512) );
  INV_X1 U8507 ( .A(n7957), .ZN(n7945) );
  INV_X1 U8508 ( .A(n8917), .ZN(n8375) );
  INV_X1 U8509 ( .A(n8361), .ZN(n8449) );
  NAND2_X1 U8510 ( .A1(n8357), .A2(n8449), .ZN(n8358) );
  NAND2_X1 U8511 ( .A1(n9542), .A2(n9689), .ZN(n9519) );
  AND2_X2 U8512 ( .A1(n9660), .A2(n9414), .ZN(n9407) );
  AOI211_X1 U8513 ( .C1(n6834), .C2(n9369), .A(n10520), .B(n9347), .ZN(n9352)
         );
  NOR2_X1 U8514 ( .A1(n9358), .A2(n9352), .ZN(n6825) );
  NAND2_X1 U8515 ( .A1(n7678), .A2(n9130), .ZN(n7379) );
  NAND3_X1 U8516 ( .A1(n6828), .A2(n6827), .A3(n7379), .ZN(n6830) );
  INV_X1 U8517 ( .A(n7377), .ZN(n6831) );
  AND2_X2 U8518 ( .A1(n6836), .A2(n6831), .ZN(n10528) );
  NAND2_X1 U8519 ( .A1(n6833), .A2(n6832), .ZN(n6835) );
  NAND2_X1 U8520 ( .A1(n6835), .A2(n5064), .ZN(P2_U3517) );
  AND2_X2 U8521 ( .A1(n6836), .A2(n7377), .ZN(n10541) );
  OR2_X1 U8522 ( .A1(n10541), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6837) );
  NAND2_X1 U8523 ( .A1(n6838), .A2(n6837), .ZN(n6839) );
  NAND2_X1 U8524 ( .A1(n6839), .A2(n5063), .ZN(P2_U3549) );
  INV_X1 U8525 ( .A(n6840), .ZN(n6841) );
  OR2_X1 U8526 ( .A1(n6478), .A2(n6841), .ZN(n9830) );
  INV_X2 U8527 ( .A(n9830), .ZN(P1_U4006) );
  NAND2_X1 U8528 ( .A1(n6478), .A2(n7100), .ZN(n6843) );
  NAND2_X1 U8529 ( .A1(n6843), .A2(n6842), .ZN(n9897) );
  NAND2_X1 U8530 ( .A1(n9897), .A2(n6844), .ZN(n6845) );
  NAND2_X1 U8531 ( .A1(n6845), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U8532 ( .A(n10465), .ZN(n10459) );
  NOR2_X2 U8533 ( .A1(n7675), .A2(n10459), .ZN(P2_U3966) );
  AND2_X1 U8534 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7548) );
  INV_X1 U8535 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n8694) );
  AOI22_X1 U8536 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n7031), .B1(n6923), .B2(
        n8694), .ZN(n7029) );
  NOR2_X1 U8537 ( .A1(n6864), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6846) );
  AOI21_X1 U8538 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n6864), .A(n6846), .ZN(
        n6980) );
  INV_X1 U8539 ( .A(n6969), .ZN(n6850) );
  XOR2_X1 U8540 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n6969), .Z(n6962) );
  NAND2_X1 U8541 ( .A1(n10311), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6847) );
  OAI21_X1 U8542 ( .B1(n10311), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6847), .ZN(
        n10316) );
  INV_X1 U8543 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6848) );
  MUX2_X1 U8544 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6848), .S(n7052), .Z(n6849)
         );
  NAND2_X1 U8545 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n7042) );
  NOR2_X1 U8546 ( .A1(n7042), .A2(n6934), .ZN(n6933) );
  AOI21_X1 U8547 ( .B1(n6890), .B2(P1_REG2_REG_1__SCAN_IN), .A(n6933), .ZN(
        n7058) );
  INV_X1 U8548 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7144) );
  XNOR2_X1 U8549 ( .A(n10293), .B(n7144), .ZN(n10292) );
  OAI21_X1 U8550 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n10293), .A(n10291), .ZN(
        n10315) );
  OAI21_X1 U8551 ( .B1(n6864), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6979), .ZN(
        n7028) );
  NAND2_X1 U8552 ( .A1(n7029), .A2(n7028), .ZN(n7027) );
  OR2_X1 U8553 ( .A1(n7031), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6851) );
  XNOR2_X1 U8554 ( .A(n7192), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n6854) );
  INV_X1 U8555 ( .A(n6852), .ZN(n6853) );
  AND2_X1 U8556 ( .A1(n6853), .A2(n9897), .ZN(n10294) );
  OAI21_X1 U8557 ( .B1(n6855), .B2(n6854), .A(n10294), .ZN(n6856) );
  NOR2_X1 U8558 ( .A1(n6856), .A2(n7193), .ZN(n6876) );
  NOR2_X1 U8559 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(n7031), .ZN(n6866) );
  NOR2_X1 U8560 ( .A1(n6864), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6865) );
  INV_X1 U8561 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10430) );
  MUX2_X1 U8562 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n10430), .S(n6969), .Z(n6965)
         );
  INV_X1 U8563 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10428) );
  INV_X1 U8564 ( .A(n10311), .ZN(n6926) );
  MUX2_X1 U8565 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10428), .S(n10311), .Z(
        n10320) );
  INV_X1 U8566 ( .A(n10293), .ZN(n6918) );
  INV_X1 U8567 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6863) );
  NAND2_X1 U8568 ( .A1(n6890), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6858) );
  INV_X1 U8569 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6857) );
  MUX2_X1 U8570 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n6857), .S(n6890), .Z(n6937)
         );
  NAND3_X1 U8571 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .A3(n6937), .ZN(n6936) );
  NAND2_X1 U8572 ( .A1(n6858), .A2(n6936), .ZN(n7051) );
  INV_X1 U8573 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6859) );
  MUX2_X1 U8574 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n6859), .S(n7052), .Z(n6860)
         );
  AND2_X1 U8575 ( .A1(n7051), .A2(n6860), .ZN(n7053) );
  AND2_X1 U8576 ( .A1(n7052), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6951) );
  INV_X1 U8577 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6861) );
  MUX2_X1 U8578 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6861), .S(n6915), .Z(n6950)
         );
  OAI21_X1 U8579 ( .B1(n7053), .B2(n6951), .A(n6950), .ZN(n6949) );
  NAND2_X1 U8580 ( .A1(n6915), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6862) );
  NAND2_X1 U8581 ( .A1(n6949), .A2(n6862), .ZN(n10297) );
  MUX2_X1 U8582 ( .A(n6863), .B(P1_REG1_REG_4__SCAN_IN), .S(n10293), .Z(n10296) );
  NOR2_X1 U8583 ( .A1(n10297), .A2(n10296), .ZN(n10298) );
  AOI21_X1 U8584 ( .B1(n6918), .B2(n6863), .A(n10298), .ZN(n10321) );
  NAND2_X1 U8585 ( .A1(n10320), .A2(n10321), .ZN(n10318) );
  OAI21_X1 U8586 ( .B1(n10428), .B2(n6926), .A(n10318), .ZN(n6966) );
  NOR2_X1 U8587 ( .A1(n6965), .A2(n6966), .ZN(n6964) );
  AOI21_X1 U8588 ( .B1(n10430), .B2(n6969), .A(n6964), .ZN(n6985) );
  INV_X1 U8589 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10432) );
  AOI22_X1 U8590 ( .A1(n6864), .A2(n10432), .B1(P1_REG1_REG_7__SCAN_IN), .B2(
        n6982), .ZN(n6984) );
  NOR2_X1 U8591 ( .A1(n6985), .A2(n6984), .ZN(n6983) );
  NOR2_X1 U8592 ( .A1(n6865), .A2(n6983), .ZN(n7026) );
  INV_X1 U8593 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10434) );
  AOI22_X1 U8594 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(n6923), .B1(n7031), .B2(
        n10434), .ZN(n7025) );
  NOR2_X1 U8595 ( .A1(n7026), .A2(n7025), .ZN(n7024) );
  NOR2_X1 U8596 ( .A1(n6866), .A2(n7024), .ZN(n6869) );
  INV_X1 U8597 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6867) );
  MUX2_X1 U8598 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n6867), .S(n7192), .Z(n6868)
         );
  OR2_X1 U8599 ( .A1(n6869), .A2(n6868), .ZN(n7187) );
  NAND2_X1 U8600 ( .A1(n6869), .A2(n6868), .ZN(n6870) );
  NOR2_X1 U8601 ( .A1(n4501), .A2(P1_U3084), .ZN(n8348) );
  AND3_X1 U8602 ( .A1(n6457), .A2(n8348), .A3(n9897), .ZN(n10319) );
  INV_X1 U8603 ( .A(n10319), .ZN(n9895) );
  AOI21_X1 U8604 ( .B1(n7187), .B2(n6870), .A(n9895), .ZN(n6875) );
  NOR2_X1 U8605 ( .A1(n6478), .A2(n6871), .ZN(n6872) );
  OR2_X1 U8606 ( .A1(P1_U3083), .A2(n6872), .ZN(n10305) );
  INV_X1 U8607 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10580) );
  AND2_X1 U8608 ( .A1(n4501), .A2(n9896), .ZN(n6873) );
  NAND2_X1 U8609 ( .A1(n9897), .A2(n6873), .ZN(n9899) );
  OAI22_X1 U8610 ( .A1(n10305), .A2(n10580), .B1(n7192), .B2(n9899), .ZN(n6874) );
  OR4_X1 U8611 ( .A1(n7548), .A2(n6876), .A3(n6875), .A4(n6874), .ZN(P1_U3250)
         );
  NOR2_X1 U8612 ( .A1(n4560), .A2(n6877), .ZN(n6878) );
  AOI21_X1 U8613 ( .B1(n4560), .B2(n6877), .A(n6878), .ZN(n7334) );
  NAND2_X1 U8614 ( .A1(n7334), .A2(n7335), .ZN(n7333) );
  INV_X1 U8615 ( .A(n6878), .ZN(n6879) );
  NAND3_X1 U8616 ( .A1(n7333), .A2(n6880), .A3(n6879), .ZN(n6881) );
  AOI21_X1 U8617 ( .B1(n6881), .B2(n7348), .A(n9795), .ZN(n6886) );
  NOR2_X1 U8618 ( .A1(n9812), .A2(n10391), .ZN(n6885) );
  AND2_X1 U8619 ( .A1(n9809), .A2(n7243), .ZN(n6884) );
  NAND2_X1 U8620 ( .A1(n9786), .A2(n9828), .ZN(n6882) );
  OR2_X1 U8621 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8817), .ZN(n6968) );
  OAI211_X1 U8622 ( .C1(n7322), .C2(n9806), .A(n6882), .B(n6968), .ZN(n6883)
         );
  OR4_X1 U8623 ( .A1(n6886), .A2(n6885), .A3(n6884), .A4(n6883), .ZN(P1_U3237)
         );
  INV_X1 U8624 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6887) );
  INV_X1 U8625 ( .A(n7704), .ZN(n8140) );
  OAI222_X1 U8626 ( .A1(n8906), .A2(n6887), .B1(n8904), .B2(n6891), .C1(
        P2_U3152), .C2(n8140), .ZN(P2_U3357) );
  NAND2_X1 U8627 ( .A1(n7128), .A2(n10354), .ZN(n6888) );
  OAI21_X1 U8628 ( .B1(n10354), .B2(n6710), .A(n6888), .ZN(P1_U3441) );
  NAND2_X1 U8629 ( .A1(n6889), .A2(P1_U3084), .ZN(n8243) );
  INV_X1 U8630 ( .A(n6890), .ZN(n6940) );
  OAI222_X1 U8631 ( .A1(n8885), .A2(n6892), .B1(n10157), .B2(n6891), .C1(n6940), .C2(P1_U3084), .ZN(P1_U3352) );
  INV_X1 U8632 ( .A(n7052), .ZN(n7060) );
  OAI222_X1 U8633 ( .A1(n8885), .A2(n6893), .B1(n10157), .B2(n6910), .C1(n7060), .C2(P1_U3084), .ZN(P1_U3351) );
  INV_X1 U8634 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6895) );
  INV_X1 U8635 ( .A(n6894), .ZN(n6908) );
  OAI222_X1 U8636 ( .A1(n8885), .A2(n6895), .B1(n10157), .B2(n6908), .C1(n6969), .C2(P1_U3084), .ZN(P1_U3347) );
  INV_X1 U8637 ( .A(n6896), .ZN(n6897) );
  OAI21_X1 U8638 ( .B1(n10354), .B2(n6696), .A(n6897), .ZN(P1_U3440) );
  INV_X1 U8639 ( .A(n8904), .ZN(n7843) );
  AOI22_X1 U8640 ( .A1(n8216), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n9698), .ZN(n6898) );
  OAI21_X1 U8641 ( .B1(n6925), .B2(n8904), .A(n6898), .ZN(P2_U3353) );
  INV_X1 U8642 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6906) );
  INV_X1 U8643 ( .A(n6457), .ZN(n8509) );
  INV_X1 U8644 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6899) );
  AOI21_X1 U8645 ( .B1(n8509), .B2(n6899), .A(n4501), .ZN(n7050) );
  XNOR2_X1 U8646 ( .A(n7050), .B(P1_IR_REG_0__SCAN_IN), .ZN(n6902) );
  INV_X1 U8647 ( .A(n9897), .ZN(n6901) );
  INV_X1 U8648 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n7023) );
  AOI21_X1 U8649 ( .B1(n8348), .B2(P1_REG1_REG_0__SCAN_IN), .A(n9896), .ZN(
        n6900) );
  NOR3_X1 U8650 ( .A1(n6902), .A2(n6901), .A3(n6900), .ZN(n6903) );
  AOI21_X1 U8651 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(P1_U3084), .A(n6903), .ZN(
        n6905) );
  NAND3_X1 U8652 ( .A1(n10319), .A2(P1_IR_REG_0__SCAN_IN), .A3(n7023), .ZN(
        n6904) );
  OAI211_X1 U8653 ( .C1(n6906), .C2(n10305), .A(n6905), .B(n6904), .ZN(
        P1_U3241) );
  INV_X1 U8654 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n8839) );
  INV_X1 U8655 ( .A(n6907), .ZN(n6928) );
  INV_X1 U8656 ( .A(n7700), .ZN(n8126) );
  OAI222_X1 U8657 ( .A1(n8906), .A2(n8839), .B1(n8904), .B2(n6928), .C1(
        P2_U3152), .C2(n8126), .ZN(P2_U3351) );
  INV_X1 U8658 ( .A(n7709), .ZN(n8191) );
  OAI222_X1 U8659 ( .A1(n8906), .A2(n5215), .B1(n8904), .B2(n6919), .C1(
        P2_U3152), .C2(n8191), .ZN(P2_U3354) );
  INV_X1 U8660 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6909) );
  INV_X1 U8661 ( .A(n7712), .ZN(n7893) );
  OAI222_X1 U8662 ( .A1(n8906), .A2(n6909), .B1(n8904), .B2(n6908), .C1(
        P2_U3152), .C2(n7893), .ZN(P2_U3352) );
  INV_X1 U8663 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6911) );
  INV_X1 U8664 ( .A(n10164), .ZN(n7706) );
  OAI222_X1 U8665 ( .A1(n8906), .A2(n6911), .B1(n8904), .B2(n6910), .C1(
        P2_U3152), .C2(n7706), .ZN(P2_U3356) );
  INV_X1 U8666 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6912) );
  INV_X1 U8667 ( .A(n7708), .ZN(n8102) );
  OAI222_X1 U8668 ( .A1(n8906), .A2(n6912), .B1(n8904), .B2(n6916), .C1(
        P2_U3152), .C2(n8102), .ZN(P2_U3355) );
  INV_X1 U8669 ( .A(n6913), .ZN(n6922) );
  INV_X1 U8670 ( .A(n7715), .ZN(n7880) );
  OAI222_X1 U8671 ( .A1(n8906), .A2(n6914), .B1(n8904), .B2(n6922), .C1(
        P2_U3152), .C2(n7880), .ZN(P2_U3350) );
  INV_X1 U8672 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6917) );
  INV_X1 U8673 ( .A(n6915), .ZN(n6955) );
  OAI222_X1 U8674 ( .A1(n8885), .A2(n6917), .B1(n10157), .B2(n6916), .C1(n6955), .C2(P1_U3084), .ZN(P1_U3350) );
  INV_X1 U8675 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6920) );
  OAI222_X1 U8676 ( .A1(n8885), .A2(n6920), .B1(n10157), .B2(n6919), .C1(n6918), .C2(P1_U3084), .ZN(P1_U3349) );
  OAI222_X1 U8677 ( .A1(n6923), .A2(P1_U3084), .B1(n10157), .B2(n6922), .C1(
        n6921), .C2(n8885), .ZN(P1_U3345) );
  OAI222_X1 U8678 ( .A1(n6926), .A2(P1_U3084), .B1(n10157), .B2(n6925), .C1(
        n6924), .C2(n8885), .ZN(P1_U3348) );
  OAI222_X1 U8679 ( .A1(n6982), .A2(P1_U3084), .B1(n10157), .B2(n6928), .C1(
        n6927), .C2(n8885), .ZN(P1_U3346) );
  INV_X1 U8680 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8748) );
  NAND2_X1 U8681 ( .A1(n9909), .A2(P1_U4006), .ZN(n6929) );
  OAI21_X1 U8682 ( .B1(P1_U4006), .B2(n8748), .A(n6929), .ZN(P1_U3586) );
  INV_X1 U8683 ( .A(n6930), .ZN(n6932) );
  INV_X1 U8684 ( .A(n7716), .ZN(n7869) );
  OAI222_X1 U8685 ( .A1(n8906), .A2(n6931), .B1(n8904), .B2(n6932), .C1(n7869), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  OAI222_X1 U8686 ( .A1(P1_U3084), .A2(n7192), .B1(n10157), .B2(n6932), .C1(
        n8753), .C2(n8885), .ZN(P1_U3344) );
  INV_X1 U8687 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6945) );
  INV_X1 U8688 ( .A(n10294), .ZN(n10313) );
  AOI211_X1 U8689 ( .C1(n7042), .C2(n6934), .A(n6933), .B(n10313), .ZN(n6943)
         );
  INV_X1 U8690 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6935) );
  NOR2_X1 U8691 ( .A1(n6935), .A2(n7023), .ZN(n6938) );
  OAI211_X1 U8692 ( .C1(n6938), .C2(n6937), .A(n10319), .B(n6936), .ZN(n6939)
         );
  INV_X1 U8693 ( .A(n6939), .ZN(n6942) );
  INV_X1 U8694 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7223) );
  OAI22_X1 U8695 ( .A1(n9899), .A2(n6940), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7223), .ZN(n6941) );
  NOR3_X1 U8696 ( .A1(n6943), .A2(n6942), .A3(n6941), .ZN(n6944) );
  OAI21_X1 U8697 ( .B1(n10305), .B2(n6945), .A(n6944), .ZN(P1_U3242) );
  INV_X1 U8698 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6960) );
  AOI211_X1 U8699 ( .C1(n6948), .C2(n6947), .A(n6946), .B(n10313), .ZN(n6958)
         );
  INV_X1 U8700 ( .A(n6949), .ZN(n6953) );
  NOR3_X1 U8701 ( .A1(n7053), .A2(n6951), .A3(n6950), .ZN(n6952) );
  NOR3_X1 U8702 ( .A1(n9895), .A2(n6953), .A3(n6952), .ZN(n6957) );
  NOR2_X1 U8703 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7292), .ZN(n7119) );
  INV_X1 U8704 ( .A(n7119), .ZN(n6954) );
  OAI21_X1 U8705 ( .B1(n9899), .B2(n6955), .A(n6954), .ZN(n6956) );
  NOR3_X1 U8706 ( .A1(n6958), .A2(n6957), .A3(n6956), .ZN(n6959) );
  OAI21_X1 U8707 ( .B1(n10305), .B2(n6960), .A(n6959), .ZN(P1_U3244) );
  INV_X1 U8708 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6974) );
  AOI211_X1 U8709 ( .C1(n6963), .C2(n6962), .A(n6961), .B(n10313), .ZN(n6972)
         );
  AOI21_X1 U8710 ( .B1(n6966), .B2(n6965), .A(n6964), .ZN(n6967) );
  NOR2_X1 U8711 ( .A1(n9895), .A2(n6967), .ZN(n6971) );
  OAI21_X1 U8712 ( .B1(n9899), .B2(n6969), .A(n6968), .ZN(n6970) );
  NOR3_X1 U8713 ( .A1(n6972), .A2(n6971), .A3(n6970), .ZN(n6973) );
  OAI21_X1 U8714 ( .B1(n10305), .B2(n6974), .A(n6973), .ZN(P1_U3247) );
  INV_X1 U8715 ( .A(n6975), .ZN(n6977) );
  OAI222_X1 U8716 ( .A1(P1_U3084), .A2(n7299), .B1(n10157), .B2(n6977), .C1(
        n6976), .C2(n8885), .ZN(P1_U3343) );
  INV_X1 U8717 ( .A(n7698), .ZN(n8114) );
  OAI222_X1 U8718 ( .A1(n8906), .A2(n6978), .B1(n8904), .B2(n6977), .C1(n8114), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U8719 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6991) );
  OAI21_X1 U8720 ( .B1(n6981), .B2(n6980), .A(n6979), .ZN(n6989) );
  NAND2_X1 U8721 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7353) );
  OAI21_X1 U8722 ( .B1(n9899), .B2(n6982), .A(n7353), .ZN(n6988) );
  AOI21_X1 U8723 ( .B1(n6985), .B2(n6984), .A(n6983), .ZN(n6986) );
  NOR2_X1 U8724 ( .A1(n9895), .A2(n6986), .ZN(n6987) );
  AOI211_X1 U8725 ( .C1(n10294), .C2(n6989), .A(n6988), .B(n6987), .ZN(n6990)
         );
  OAI21_X1 U8726 ( .B1(n6991), .B2(n10305), .A(n6990), .ZN(P1_U3248) );
  INV_X1 U8727 ( .A(n6992), .ZN(n6994) );
  OAI222_X1 U8728 ( .A1(n8885), .A2(n6993), .B1(n10157), .B2(n6994), .C1(
        P1_U3084), .C2(n7422), .ZN(P1_U3342) );
  INV_X1 U8729 ( .A(n9287), .ZN(n7718) );
  OAI222_X1 U8730 ( .A1(n8906), .A2(n6995), .B1(n8904), .B2(n6994), .C1(n7718), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  AND2_X1 U8731 ( .A1(n6997), .A2(n6996), .ZN(n7020) );
  INV_X1 U8732 ( .A(n7019), .ZN(n7130) );
  AND3_X1 U8733 ( .A1(n6999), .A2(n10354), .A3(n6998), .ZN(n7129) );
  AND3_X2 U8734 ( .A1(n7020), .A2(n7130), .A3(n7129), .ZN(n10424) );
  INV_X1 U8735 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7006) );
  INV_X1 U8736 ( .A(n7141), .ZN(n7004) );
  NAND2_X1 U8737 ( .A1(n4501), .A2(n7000), .ZN(n10338) );
  INV_X1 U8738 ( .A(n10338), .ZN(n10056) );
  NOR3_X1 U8739 ( .A1(n7002), .A2(n7001), .A3(n7141), .ZN(n7003) );
  AOI21_X1 U8740 ( .B1(n10056), .B2(n6410), .A(n7003), .ZN(n7203) );
  OAI21_X1 U8741 ( .B1(n7221), .B2(n7004), .A(n7203), .ZN(n7021) );
  NAND2_X1 U8742 ( .A1(n7021), .A2(n10424), .ZN(n7005) );
  OAI21_X1 U8743 ( .B1(n10424), .B2(n7006), .A(n7005), .ZN(P1_U3454) );
  OR2_X1 U8744 ( .A1(n10450), .A2(n7007), .ZN(n7012) );
  OR2_X1 U8745 ( .A1(n7008), .A2(P2_U3152), .ZN(n9134) );
  NAND2_X1 U8746 ( .A1(n10450), .A2(n9134), .ZN(n7010) );
  NAND2_X1 U8747 ( .A1(n7010), .A2(n7009), .ZN(n7011) );
  AND2_X1 U8748 ( .A1(n7012), .A2(n7011), .ZN(n9339) );
  NOR2_X1 U8749 ( .A1(n10441), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8750 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n7018) );
  INV_X1 U8751 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n9642) );
  NAND2_X1 U8752 ( .A1(n7013), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n7016) );
  INV_X1 U8753 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9571) );
  OR2_X1 U8754 ( .A1(n7014), .A2(n9571), .ZN(n7015) );
  OAI211_X1 U8755 ( .C1(n4498), .C2(n9642), .A(n7016), .B(n7015), .ZN(n9343)
         );
  NAND2_X1 U8756 ( .A1(n9343), .A2(P2_U3966), .ZN(n7017) );
  OAI21_X1 U8757 ( .B1(P2_U3966), .B2(n7018), .A(n7017), .ZN(P2_U3583) );
  NAND3_X1 U8758 ( .A1(n7020), .A2(n7129), .A3(n7019), .ZN(n10436) );
  NAND2_X1 U8759 ( .A1(n7021), .A2(n10438), .ZN(n7022) );
  OAI21_X1 U8760 ( .B1(n10438), .B2(n7023), .A(n7022), .ZN(P1_U3523) );
  AOI21_X1 U8761 ( .B1(n7026), .B2(n7025), .A(n7024), .ZN(n7037) );
  OAI21_X1 U8762 ( .B1(n7029), .B2(n7028), .A(n7027), .ZN(n7035) );
  INV_X1 U8763 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10583) );
  NOR2_X1 U8764 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7030), .ZN(n7489) );
  INV_X1 U8765 ( .A(n7489), .ZN(n7033) );
  INV_X1 U8766 ( .A(n9899), .ZN(n10310) );
  NAND2_X1 U8767 ( .A1(n10310), .A2(n7031), .ZN(n7032) );
  OAI211_X1 U8768 ( .C1(n10305), .C2(n10583), .A(n7033), .B(n7032), .ZN(n7034)
         );
  AOI21_X1 U8769 ( .B1(n7035), .B2(n10294), .A(n7034), .ZN(n7036) );
  OAI21_X1 U8770 ( .B1(n7037), .B2(n9895), .A(n7036), .ZN(P1_U3249) );
  INV_X1 U8771 ( .A(n7606), .ZN(n7598) );
  INV_X1 U8772 ( .A(n7038), .ZN(n7040) );
  OAI222_X1 U8773 ( .A1(n7598), .A2(P1_U3084), .B1(n8243), .B2(n7040), .C1(
        n7039), .C2(n8885), .ZN(P1_U3341) );
  INV_X1 U8774 ( .A(n8203), .ZN(n7720) );
  OAI222_X1 U8775 ( .A1(n8906), .A2(n7041), .B1(n8904), .B2(n7040), .C1(
        P2_U3152), .C2(n7720), .ZN(P2_U3346) );
  INV_X1 U8776 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7065) );
  INV_X1 U8777 ( .A(n7042), .ZN(n7047) );
  OAI21_X1 U8778 ( .B1(n7045), .B2(n7044), .A(n7043), .ZN(n7081) );
  INV_X1 U8779 ( .A(n7081), .ZN(n7046) );
  MUX2_X1 U8780 ( .A(n7047), .B(n7046), .S(n6457), .Z(n7048) );
  NAND2_X1 U8781 ( .A1(n7048), .A2(n4500), .ZN(n7049) );
  OAI211_X1 U8782 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n7050), .A(n7049), .B(
        P1_U4006), .ZN(n10307) );
  INV_X1 U8783 ( .A(n7051), .ZN(n7055) );
  MUX2_X1 U8784 ( .A(n6859), .B(P1_REG1_REG_2__SCAN_IN), .S(n7052), .Z(n7054)
         );
  AOI211_X1 U8785 ( .C1(n7055), .C2(n7054), .A(n7053), .B(n9895), .ZN(n7063)
         );
  AOI211_X1 U8786 ( .C1(n7058), .C2(n7057), .A(n7056), .B(n10313), .ZN(n7062)
         );
  INV_X1 U8787 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7059) );
  OAI22_X1 U8788 ( .A1(n9899), .A2(n7060), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7059), .ZN(n7061) );
  NOR3_X1 U8789 ( .A1(n7063), .A2(n7062), .A3(n7061), .ZN(n7064) );
  OAI211_X1 U8790 ( .C1(n7065), .C2(n10305), .A(n10307), .B(n7064), .ZN(
        P1_U3243) );
  NOR2_X1 U8791 ( .A1(n7066), .A2(P1_U3084), .ZN(n8882) );
  INV_X1 U8792 ( .A(n7070), .ZN(n7074) );
  XOR2_X1 U8793 ( .A(n7068), .B(n7067), .Z(n7071) );
  OAI21_X1 U8794 ( .B1(n7071), .B2(n7070), .A(n7069), .ZN(n7072) );
  OAI21_X1 U8795 ( .B1(n7074), .B2(n7073), .A(n7072), .ZN(n7075) );
  NAND2_X1 U8796 ( .A1(n7075), .A2(n9802), .ZN(n7079) );
  INV_X1 U8797 ( .A(n9806), .ZN(n9768) );
  INV_X1 U8798 ( .A(n7338), .ZN(n7360) );
  INV_X1 U8799 ( .A(n10133), .ZN(n10414) );
  OR2_X1 U8800 ( .A1(n7222), .A2(n10414), .ZN(n10367) );
  OAI22_X1 U8801 ( .A1(n7360), .A2(n10367), .B1(n9804), .B2(n4732), .ZN(n7077)
         );
  AOI21_X1 U8802 ( .B1(n9768), .B2(n7076), .A(n7077), .ZN(n7078) );
  OAI211_X1 U8803 ( .C1(n8882), .C2(n7223), .A(n7079), .B(n7078), .ZN(P1_U3220) );
  NAND2_X1 U8804 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(n9280), .ZN(n7080) );
  OAI21_X1 U8805 ( .B1(n9049), .B2(n9280), .A(n7080), .ZN(P2_U3565) );
  INV_X1 U8806 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7084) );
  NAND2_X1 U8807 ( .A1(n7081), .A2(n9802), .ZN(n7083) );
  AOI22_X1 U8808 ( .A1(n9792), .A2(n7205), .B1(n9768), .B2(n6410), .ZN(n7082)
         );
  OAI211_X1 U8809 ( .C1(n8882), .C2(n7084), .A(n7083), .B(n7082), .ZN(P1_U3230) );
  INV_X1 U8810 ( .A(n7085), .ZN(n7087) );
  OAI222_X1 U8811 ( .A1(n8885), .A2(n7086), .B1(n10157), .B2(n7087), .C1(
        P1_U3084), .C2(n8009), .ZN(P1_U3340) );
  INV_X1 U8812 ( .A(n7835), .ZN(n7831) );
  OAI222_X1 U8813 ( .A1(n8906), .A2(n7088), .B1(n8904), .B2(n7087), .C1(n7831), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U8814 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n7106) );
  INV_X1 U8815 ( .A(n10368), .ZN(n10410) );
  NAND2_X1 U8816 ( .A1(n9831), .A2(n7205), .ZN(n7210) );
  NAND2_X1 U8817 ( .A1(n4733), .A2(n7222), .ZN(n7089) );
  NAND2_X1 U8818 ( .A1(n7209), .A2(n7089), .ZN(n7091) );
  NAND2_X1 U8819 ( .A1(n7091), .A2(n7090), .ZN(n7124) );
  OR2_X1 U8820 ( .A1(n7091), .A2(n7090), .ZN(n7092) );
  NAND2_X1 U8821 ( .A1(n7124), .A2(n7092), .ZN(n7277) );
  AND2_X1 U8822 ( .A1(n7141), .A2(n7557), .ZN(n10265) );
  OAI211_X1 U8823 ( .C1(n7219), .C2(n7272), .A(n10265), .B(n7289), .ZN(n7275)
         );
  OAI21_X1 U8824 ( .B1(n7272), .B2(n10414), .A(n7275), .ZN(n7104) );
  INV_X1 U8825 ( .A(n7093), .ZN(n10253) );
  NAND2_X1 U8826 ( .A1(n7277), .A2(n10253), .ZN(n7103) );
  OR2_X1 U8827 ( .A1(n7803), .A2(n7367), .ZN(n7097) );
  NAND2_X1 U8828 ( .A1(n7095), .A2(n7140), .ZN(n7096) );
  NAND2_X1 U8829 ( .A1(n7097), .A2(n7096), .ZN(n10343) );
  NAND2_X1 U8830 ( .A1(n7098), .A2(n10343), .ZN(n7102) );
  NOR2_X2 U8831 ( .A1(n4501), .A2(n7100), .ZN(n10054) );
  AOI22_X1 U8832 ( .A1(n7099), .A2(n10056), .B1(n10054), .B2(n6410), .ZN(n7101) );
  NAND3_X1 U8833 ( .A1(n7103), .A2(n7102), .A3(n7101), .ZN(n7270) );
  AOI211_X1 U8834 ( .C1(n10410), .C2(n7277), .A(n7104), .B(n7270), .ZN(n7107)
         );
  OR2_X1 U8835 ( .A1(n7107), .A2(n10422), .ZN(n7105) );
  OAI21_X1 U8836 ( .B1(n10424), .B2(n7106), .A(n7105), .ZN(P1_U3460) );
  OR2_X1 U8837 ( .A1(n7107), .A2(n10436), .ZN(n7108) );
  OAI21_X1 U8838 ( .B1(n10438), .B2(n6859), .A(n7108), .ZN(P1_U3525) );
  INV_X1 U8839 ( .A(n7109), .ZN(n7111) );
  INV_X1 U8840 ( .A(n8079), .ZN(n8086) );
  OAI222_X1 U8841 ( .A1(n8906), .A2(n8520), .B1(n8904), .B2(n7111), .C1(n8086), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U8842 ( .A(n8010), .ZN(n8284) );
  OAI222_X1 U8843 ( .A1(P1_U3084), .A2(n8284), .B1(n10157), .B2(n7111), .C1(
        n7110), .C2(n8885), .ZN(P1_U3339) );
  INV_X1 U8844 ( .A(n7112), .ZN(n7113) );
  NOR2_X1 U8845 ( .A1(n7114), .A2(n7113), .ZN(n7117) );
  INV_X1 U8846 ( .A(n7115), .ZN(n7116) );
  AOI21_X1 U8847 ( .B1(n7117), .B2(n8873), .A(n7116), .ZN(n7122) );
  NOR2_X1 U8848 ( .A1(n9804), .A2(n7285), .ZN(n7118) );
  AOI211_X1 U8849 ( .C1(n9768), .C2(n9829), .A(n7119), .B(n7118), .ZN(n7121)
         );
  AOI22_X1 U8850 ( .A1(n9792), .A2(n6180), .B1(n9809), .B2(n7292), .ZN(n7120)
         );
  OAI211_X1 U8851 ( .C1(n7122), .C2(n9795), .A(n7121), .B(n7120), .ZN(P1_U3216) );
  NAND2_X1 U8852 ( .A1(n7285), .A2(n7272), .ZN(n7123) );
  NAND2_X1 U8853 ( .A1(n7124), .A2(n7123), .ZN(n7283) );
  NAND2_X1 U8854 ( .A1(n7283), .A2(n7282), .ZN(n7281) );
  NAND2_X1 U8855 ( .A1(n8877), .A2(n10373), .ZN(n7125) );
  NAND2_X1 U8856 ( .A1(n7281), .A2(n7125), .ZN(n7168) );
  NAND2_X1 U8857 ( .A1(n7127), .A2(n7126), .ZN(n7167) );
  XOR2_X1 U8858 ( .A(n7168), .B(n7167), .Z(n10379) );
  NAND3_X1 U8859 ( .A1(n7130), .A2(n7129), .A3(n7128), .ZN(n7139) );
  NAND2_X1 U8860 ( .A1(n7139), .A2(n8230), .ZN(n10349) );
  NOR2_X1 U8861 ( .A1(n7131), .A2(n7367), .ZN(n7132) );
  NAND2_X1 U8862 ( .A1(n10349), .A2(n7132), .ZN(n8161) );
  XOR2_X1 U8863 ( .A(n7167), .B(n7251), .Z(n7134) );
  INV_X1 U8864 ( .A(n10054), .ZN(n10340) );
  OAI22_X1 U8865 ( .A1(n8877), .A2(n10340), .B1(n7155), .B2(n10338), .ZN(n7133) );
  AOI21_X1 U8866 ( .B1(n7134), .B2(n10343), .A(n7133), .ZN(n7135) );
  OAI21_X1 U8867 ( .B1(n10379), .B2(n7093), .A(n7135), .ZN(n10380) );
  NAND2_X1 U8868 ( .A1(n10380), .A2(n10349), .ZN(n7147) );
  XNOR2_X1 U8869 ( .A(n7291), .B(n7166), .ZN(n7136) );
  NAND2_X1 U8870 ( .A1(n7136), .A2(n10265), .ZN(n7138) );
  NAND2_X1 U8871 ( .A1(n6179), .A2(n10133), .ZN(n7137) );
  NAND2_X1 U8872 ( .A1(n7138), .A2(n7137), .ZN(n10381) );
  OR2_X1 U8873 ( .A1(n7139), .A2(n9902), .ZN(n8235) );
  INV_X1 U8874 ( .A(n10265), .ZN(n10416) );
  NOR2_X2 U8875 ( .A1(n8235), .A2(n10416), .ZN(n10331) );
  INV_X1 U8876 ( .A(n10331), .ZN(n7774) );
  AND2_X1 U8877 ( .A1(n7141), .A2(n7140), .ZN(n7142) );
  NAND2_X1 U8878 ( .A1(n10349), .A2(n7142), .ZN(n10256) );
  NAND2_X1 U8879 ( .A1(n7774), .A2(n10256), .ZN(n7206) );
  INV_X1 U8880 ( .A(n7151), .ZN(n7143) );
  OAI22_X1 U8881 ( .A1(n10349), .A2(n7144), .B1(n7143), .B2(n8230), .ZN(n7145)
         );
  AOI21_X1 U8882 ( .B1(n10381), .B2(n7206), .A(n7145), .ZN(n7146) );
  OAI211_X1 U8883 ( .C1(n10379), .C2(n8161), .A(n7147), .B(n7146), .ZN(
        P1_U3287) );
  OAI21_X1 U8884 ( .B1(n7150), .B2(n7149), .A(n7148), .ZN(n7157) );
  AOI22_X1 U8885 ( .A1(n9792), .A2(n6179), .B1(n7151), .B2(n9809), .ZN(n7154)
         );
  INV_X1 U8886 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n7152) );
  NOR2_X1 U8887 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7152), .ZN(n10301) );
  AOI21_X1 U8888 ( .B1(n9786), .B2(n7099), .A(n10301), .ZN(n7153) );
  OAI211_X1 U8889 ( .C1(n7155), .C2(n9806), .A(n7154), .B(n7153), .ZN(n7156)
         );
  AOI21_X1 U8890 ( .B1(n7157), .B2(n9802), .A(n7156), .ZN(n7158) );
  INV_X1 U8891 ( .A(n7158), .ZN(P1_U3228) );
  NAND2_X1 U8892 ( .A1(n9830), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7159) );
  OAI21_X1 U8893 ( .B1(n9927), .B2(n9830), .A(n7159), .ZN(P1_U3584) );
  INV_X1 U8894 ( .A(n9839), .ZN(n9832) );
  INV_X1 U8895 ( .A(n7160), .ZN(n7161) );
  OAI222_X1 U8896 ( .A1(n9832), .A2(P1_U3084), .B1(n10157), .B2(n7161), .C1(
        n8662), .C2(n8885), .ZN(P1_U3338) );
  INV_X1 U8897 ( .A(n8380), .ZN(n8391) );
  OAI222_X1 U8898 ( .A1(n8906), .A2(n8653), .B1(n8904), .B2(n7161), .C1(
        P2_U3152), .C2(n8391), .ZN(P2_U3343) );
  INV_X1 U8899 ( .A(n7162), .ZN(n7201) );
  AOI22_X1 U8900 ( .A1(n9304), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n9698), .ZN(n7163) );
  OAI21_X1 U8901 ( .B1(n7201), .B2(n8904), .A(n7163), .ZN(P2_U3342) );
  XOR2_X1 U8902 ( .A(n7169), .B(n7164), .Z(n7165) );
  INV_X1 U8903 ( .A(n10343), .ZN(n9988) );
  OAI222_X1 U8904 ( .A1(n10340), .A2(n7284), .B1(n10338), .B2(n7258), .C1(
        n7165), .C2(n9988), .ZN(n10388) );
  AOI21_X1 U8905 ( .B1(n7168), .B2(n7167), .A(n5068), .ZN(n7171) );
  OAI21_X1 U8906 ( .B1(n7171), .B2(n7170), .A(n7238), .ZN(n10384) );
  AND2_X1 U8907 ( .A1(n7173), .A2(n7172), .ZN(n7174) );
  AND2_X1 U8908 ( .A1(n10349), .A2(n7174), .ZN(n8864) );
  INV_X1 U8909 ( .A(n8864), .ZN(n10062) );
  INV_X1 U8910 ( .A(n10256), .ZN(n8238) );
  INV_X1 U8911 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7176) );
  OAI22_X1 U8912 ( .A1(n10349), .A2(n7176), .B1(n7175), .B2(n8230), .ZN(n7177)
         );
  AOI21_X1 U8913 ( .B1(n8238), .B2(n7236), .A(n7177), .ZN(n7181) );
  OAI21_X1 U8914 ( .B1(n7178), .B2(n7337), .A(n10265), .ZN(n7179) );
  NOR2_X1 U8915 ( .A1(n7179), .A2(n7242), .ZN(n10385) );
  INV_X1 U8916 ( .A(n8235), .ZN(n10041) );
  NAND2_X1 U8917 ( .A1(n10385), .A2(n10041), .ZN(n7180) );
  OAI211_X1 U8918 ( .C1(n10384), .C2(n10062), .A(n7181), .B(n7180), .ZN(n7182)
         );
  AOI21_X1 U8919 ( .B1(n10388), .B2(n10349), .A(n7182), .ZN(n7183) );
  INV_X1 U8920 ( .A(n7183), .ZN(P1_U3286) );
  NAND2_X1 U8921 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n9280), .ZN(n7184) );
  OAI21_X1 U8922 ( .B1(n7185), .B2(n9280), .A(n7184), .ZN(P2_U3581) );
  NAND2_X1 U8923 ( .A1(n7192), .A2(n6867), .ZN(n7186) );
  AND2_X1 U8924 ( .A1(n7187), .A2(n7186), .ZN(n7189) );
  INV_X1 U8925 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10179) );
  AOI22_X1 U8926 ( .A1(n7305), .A2(n10179), .B1(P1_REG1_REG_10__SCAN_IN), .B2(
        n7299), .ZN(n7188) );
  NOR2_X1 U8927 ( .A1(n7189), .A2(n7188), .ZN(n7298) );
  AOI21_X1 U8928 ( .B1(n7189), .B2(n7188), .A(n7298), .ZN(n7200) );
  INV_X1 U8929 ( .A(n10305), .ZN(n10312) );
  INV_X1 U8930 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7190) );
  NOR2_X1 U8931 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7190), .ZN(n7640) );
  INV_X1 U8932 ( .A(n7640), .ZN(n7191) );
  OAI21_X1 U8933 ( .B1(n9899), .B2(n7299), .A(n7191), .ZN(n7198) );
  NAND2_X1 U8934 ( .A1(n7305), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7194) );
  OAI21_X1 U8935 ( .B1(n7305), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7194), .ZN(
        n7195) );
  AOI211_X1 U8936 ( .C1(n7196), .C2(n7195), .A(n10313), .B(n7304), .ZN(n7197)
         );
  AOI211_X1 U8937 ( .C1(n10312), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n7198), .B(
        n7197), .ZN(n7199) );
  OAI21_X1 U8938 ( .B1(n7200), .B2(n9895), .A(n7199), .ZN(P1_U3251) );
  INV_X1 U8939 ( .A(n9858), .ZN(n9853) );
  OAI222_X1 U8940 ( .A1(n8885), .A2(n7202), .B1(n10157), .B2(n7201), .C1(
        P1_U3084), .C2(n9853), .ZN(P1_U3337) );
  INV_X1 U8941 ( .A(n8230), .ZN(n10345) );
  INV_X1 U8942 ( .A(n7203), .ZN(n7204) );
  AOI21_X1 U8943 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n10345), .A(n7204), .ZN(
        n7208) );
  AOI22_X1 U8944 ( .A1(n7206), .A2(n7205), .B1(P1_REG2_REG_0__SCAN_IN), .B2(
        n10048), .ZN(n7207) );
  OAI21_X1 U8945 ( .B1(n7208), .B2(n10048), .A(n7207), .ZN(P1_U3291) );
  OAI21_X1 U8946 ( .B1(n7211), .B2(n7210), .A(n7209), .ZN(n7212) );
  INV_X1 U8947 ( .A(n7212), .ZN(n10369) );
  OAI21_X1 U8948 ( .B1(n7215), .B2(n7214), .A(n7213), .ZN(n7217) );
  OAI22_X1 U8949 ( .A1(n4732), .A2(n10340), .B1(n7285), .B2(n10338), .ZN(n7216) );
  AOI21_X1 U8950 ( .B1(n7217), .B2(n10343), .A(n7216), .ZN(n7218) );
  OAI21_X1 U8951 ( .B1(n10369), .B2(n7093), .A(n7218), .ZN(n10371) );
  INV_X1 U8952 ( .A(n7219), .ZN(n7220) );
  OAI211_X1 U8953 ( .C1(n7222), .C2(n7221), .A(n7220), .B(n10265), .ZN(n10366)
         );
  OAI22_X1 U8954 ( .A1(n10366), .A2(n9902), .B1(n8230), .B2(n7223), .ZN(n7224)
         );
  OAI21_X1 U8955 ( .B1(n10371), .B2(n7224), .A(n10349), .ZN(n7227) );
  AOI22_X1 U8956 ( .A1(n8238), .A2(n7225), .B1(n10048), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n7226) );
  OAI211_X1 U8957 ( .C1(n10369), .C2(n8161), .A(n7227), .B(n7226), .ZN(
        P1_U3290) );
  INV_X1 U8958 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7229) );
  INV_X1 U8959 ( .A(n7228), .ZN(n7231) );
  OAI222_X1 U8960 ( .A1(n8906), .A2(n7229), .B1(n8904), .B2(n7231), .C1(n9311), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  INV_X1 U8961 ( .A(n9877), .ZN(n9871) );
  INV_X1 U8962 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7230) );
  OAI222_X1 U8963 ( .A1(P1_U3084), .A2(n9871), .B1(n10157), .B2(n7231), .C1(
        n7230), .C2(n8885), .ZN(P1_U3336) );
  XNOR2_X1 U8964 ( .A(n7232), .B(n7240), .ZN(n7233) );
  NAND2_X1 U8965 ( .A1(n7233), .A2(n10343), .ZN(n7235) );
  AOI22_X1 U8966 ( .A1(n9828), .A2(n10054), .B1(n10056), .B2(n9826), .ZN(n7234) );
  NAND2_X1 U8967 ( .A1(n7235), .A2(n7234), .ZN(n10392) );
  INV_X1 U8968 ( .A(n10392), .ZN(n7249) );
  NAND2_X1 U8969 ( .A1(n9828), .A2(n7236), .ZN(n7237) );
  OAI21_X1 U8970 ( .B1(n7241), .B2(n7240), .A(n7260), .ZN(n10394) );
  NAND2_X1 U8971 ( .A1(n7242), .A2(n10391), .ZN(n7263) );
  OAI211_X1 U8972 ( .C1(n7242), .C2(n10391), .A(n10265), .B(n7263), .ZN(n10390) );
  AOI22_X1 U8973 ( .A1(n10048), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7243), .B2(
        n10345), .ZN(n7246) );
  NAND2_X1 U8974 ( .A1(n8238), .A2(n7244), .ZN(n7245) );
  OAI211_X1 U8975 ( .C1(n10390), .C2(n8235), .A(n7246), .B(n7245), .ZN(n7247)
         );
  AOI21_X1 U8976 ( .B1(n10394), .B2(n8864), .A(n7247), .ZN(n7248) );
  OAI21_X1 U8977 ( .B1(n10048), .B2(n7249), .A(n7248), .ZN(P1_U3285) );
  NAND2_X1 U8978 ( .A1(n7251), .A2(n7250), .ZN(n7255) );
  NAND2_X1 U8979 ( .A1(n7255), .A2(n7254), .ZN(n7253) );
  NAND2_X1 U8980 ( .A1(n7253), .A2(n7252), .ZN(n7319) );
  NAND3_X1 U8981 ( .A1(n7255), .A2(n7261), .A3(n7254), .ZN(n7256) );
  NAND2_X1 U8982 ( .A1(n7319), .A2(n7256), .ZN(n7257) );
  INV_X1 U8983 ( .A(n10341), .ZN(n9825) );
  AOI222_X1 U8984 ( .A1(n10343), .A2(n7257), .B1(n9825), .B2(n10056), .C1(
        n9827), .C2(n10054), .ZN(n10397) );
  NAND2_X1 U8985 ( .A1(n7258), .A2(n10391), .ZN(n7259) );
  NAND2_X1 U8986 ( .A1(n7262), .A2(n7261), .ZN(n7314) );
  OAI21_X1 U8987 ( .B1(n7262), .B2(n7261), .A(n7314), .ZN(n10400) );
  NAND2_X1 U8988 ( .A1(n10400), .A2(n8864), .ZN(n7269) );
  INV_X1 U8989 ( .A(n7263), .ZN(n7264) );
  OR2_X2 U8990 ( .A1(n7263), .A2(n7347), .ZN(n7327) );
  OAI21_X1 U8991 ( .B1(n7264), .B2(n7312), .A(n7327), .ZN(n10398) );
  INV_X1 U8992 ( .A(n10398), .ZN(n7267) );
  AOI22_X1 U8993 ( .A1(n10048), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7357), .B2(
        n10345), .ZN(n7265) );
  OAI21_X1 U8994 ( .B1(n7312), .B2(n10256), .A(n7265), .ZN(n7266) );
  AOI21_X1 U8995 ( .B1(n7267), .B2(n10331), .A(n7266), .ZN(n7268) );
  OAI211_X1 U8996 ( .C1(n10397), .C2(n10048), .A(n7269), .B(n7268), .ZN(
        P1_U3284) );
  MUX2_X1 U8997 ( .A(n7270), .B(P1_REG2_REG_2__SCAN_IN), .S(n10048), .Z(n7271)
         );
  INV_X1 U8998 ( .A(n7271), .ZN(n7279) );
  INV_X1 U8999 ( .A(n8161), .ZN(n10332) );
  OAI22_X1 U9000 ( .A1(n10256), .A2(n7272), .B1(n8230), .B2(n7059), .ZN(n7273)
         );
  INV_X1 U9001 ( .A(n7273), .ZN(n7274) );
  OAI21_X1 U9002 ( .B1(n7275), .B2(n8235), .A(n7274), .ZN(n7276) );
  AOI21_X1 U9003 ( .B1(n7277), .B2(n10332), .A(n7276), .ZN(n7278) );
  NAND2_X1 U9004 ( .A1(n7279), .A2(n7278), .ZN(P1_U3289) );
  XNOR2_X1 U9005 ( .A(n7282), .B(n7280), .ZN(n7288) );
  OAI21_X1 U9006 ( .B1(n7283), .B2(n7282), .A(n7281), .ZN(n10377) );
  OAI22_X1 U9007 ( .A1(n7285), .A2(n10340), .B1(n7284), .B2(n10338), .ZN(n7286) );
  AOI21_X1 U9008 ( .B1(n10377), .B2(n10253), .A(n7286), .ZN(n7287) );
  OAI21_X1 U9009 ( .B1(n9988), .B2(n7288), .A(n7287), .ZN(n10375) );
  INV_X1 U9010 ( .A(n10375), .ZN(n7297) );
  NAND2_X1 U9011 ( .A1(n7289), .A2(n6180), .ZN(n7290) );
  NAND2_X1 U9012 ( .A1(n7291), .A2(n7290), .ZN(n10374) );
  AOI22_X1 U9013 ( .A1(n10048), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n10345), .B2(
        n7292), .ZN(n7294) );
  NAND2_X1 U9014 ( .A1(n8238), .A2(n6180), .ZN(n7293) );
  OAI211_X1 U9015 ( .C1(n7774), .C2(n10374), .A(n7294), .B(n7293), .ZN(n7295)
         );
  AOI21_X1 U9016 ( .B1(n10377), .B2(n10332), .A(n7295), .ZN(n7296) );
  OAI21_X1 U9017 ( .B1(n7297), .B2(n10048), .A(n7296), .ZN(P1_U3288) );
  AOI21_X1 U9018 ( .B1(n7299), .B2(n10179), .A(n7298), .ZN(n7302) );
  INV_X1 U9019 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7300) );
  MUX2_X1 U9020 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n7300), .S(n7422), .Z(n7301)
         );
  NOR2_X1 U9021 ( .A1(n7302), .A2(n7301), .ZN(n7425) );
  AOI21_X1 U9022 ( .B1(n7302), .B2(n7301), .A(n7425), .ZN(n7311) );
  INV_X1 U9023 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7303) );
  XNOR2_X1 U9024 ( .A(n7422), .B(n7303), .ZN(n7430) );
  XNOR2_X1 U9025 ( .A(n7430), .B(n7429), .ZN(n7309) );
  NAND2_X1 U9026 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7669) );
  OAI21_X1 U9027 ( .B1(n9899), .B2(n7422), .A(n7669), .ZN(n7308) );
  INV_X1 U9028 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7306) );
  NOR2_X1 U9029 ( .A1(n10305), .A2(n7306), .ZN(n7307) );
  AOI211_X1 U9030 ( .C1(n10294), .C2(n7309), .A(n7308), .B(n7307), .ZN(n7310)
         );
  OAI21_X1 U9031 ( .B1(n7311), .B2(n9895), .A(n7310), .ZN(P1_U3252) );
  NAND2_X1 U9032 ( .A1(n7312), .A2(n7322), .ZN(n7313) );
  NAND2_X1 U9033 ( .A1(n7314), .A2(n7313), .ZN(n7316) );
  NAND2_X1 U9034 ( .A1(n7316), .A2(n7320), .ZN(n7317) );
  NAND2_X1 U9035 ( .A1(n7398), .A2(n7317), .ZN(n10403) );
  OAI22_X1 U9036 ( .A1(n7322), .A2(n10340), .B1(n7321), .B2(n10338), .ZN(n7323) );
  AOI21_X1 U9037 ( .B1(n7324), .B2(n10343), .A(n7323), .ZN(n7325) );
  OAI21_X1 U9038 ( .B1(n10403), .B2(n7093), .A(n7325), .ZN(n10407) );
  NAND2_X1 U9039 ( .A1(n10407), .A2(n10349), .ZN(n7332) );
  INV_X1 U9040 ( .A(n7490), .ZN(n7326) );
  OAI22_X1 U9041 ( .A1(n10349), .A2(n8694), .B1(n7326), .B2(n8230), .ZN(n7330)
         );
  AND2_X1 U9042 ( .A1(n7327), .A2(n10404), .ZN(n7328) );
  OR2_X1 U9043 ( .A1(n7328), .A2(n10327), .ZN(n10406) );
  NOR2_X1 U9044 ( .A1(n10406), .A2(n7774), .ZN(n7329) );
  AOI211_X1 U9045 ( .C1(n8238), .C2(n10404), .A(n7330), .B(n7329), .ZN(n7331)
         );
  OAI211_X1 U9046 ( .C1(n10403), .C2(n8161), .A(n7332), .B(n7331), .ZN(
        P1_U3283) );
  OAI21_X1 U9047 ( .B1(n7335), .B2(n7334), .A(n7333), .ZN(n7345) );
  NAND2_X1 U9048 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10324) );
  INV_X1 U9049 ( .A(n10324), .ZN(n7336) );
  AOI21_X1 U9050 ( .B1(n9786), .B2(n9829), .A(n7336), .ZN(n7343) );
  NOR2_X1 U9051 ( .A1(n7337), .A2(n10414), .ZN(n10386) );
  NAND2_X1 U9052 ( .A1(n10386), .A2(n7338), .ZN(n7342) );
  NAND2_X1 U9053 ( .A1(n9809), .A2(n7339), .ZN(n7341) );
  NAND2_X1 U9054 ( .A1(n9768), .A2(n9827), .ZN(n7340) );
  NAND4_X1 U9055 ( .A1(n7343), .A2(n7342), .A3(n7341), .A4(n7340), .ZN(n7344)
         );
  AOI21_X1 U9056 ( .B1(n7345), .B2(n9802), .A(n7344), .ZN(n7346) );
  INV_X1 U9057 ( .A(n7346), .ZN(P1_U3225) );
  NAND2_X1 U9058 ( .A1(n7347), .A2(n10133), .ZN(n10396) );
  INV_X1 U9059 ( .A(n7348), .ZN(n7351) );
  NOR3_X1 U9060 ( .A1(n7351), .A2(n4992), .A3(n7350), .ZN(n7352) );
  OAI21_X1 U9061 ( .B1(n7352), .B2(n4561), .A(n9802), .ZN(n7359) );
  INV_X1 U9062 ( .A(n7353), .ZN(n7354) );
  AOI21_X1 U9063 ( .B1(n9786), .B2(n9827), .A(n7354), .ZN(n7355) );
  OAI21_X1 U9064 ( .B1(n10341), .B2(n9806), .A(n7355), .ZN(n7356) );
  AOI21_X1 U9065 ( .B1(n7357), .B2(n9809), .A(n7356), .ZN(n7358) );
  OAI211_X1 U9066 ( .C1(n7360), .C2(n10396), .A(n7359), .B(n7358), .ZN(
        P1_U3211) );
  INV_X1 U9067 ( .A(n9892), .ZN(n9887) );
  INV_X1 U9068 ( .A(n7361), .ZN(n7363) );
  INV_X1 U9069 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7362) );
  OAI222_X1 U9070 ( .A1(n9887), .A2(P1_U3084), .B1(n10157), .B2(n7363), .C1(
        n7362), .C2(n8885), .ZN(P1_U3335) );
  INV_X1 U9071 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7364) );
  INV_X1 U9072 ( .A(n9320), .ZN(n9332) );
  OAI222_X1 U9073 ( .A1(n8906), .A2(n7364), .B1(n8904), .B2(n7363), .C1(
        P2_U3152), .C2(n9332), .ZN(P2_U3340) );
  INV_X1 U9074 ( .A(n7365), .ZN(n7368) );
  OAI222_X1 U9075 ( .A1(P1_U3084), .A2(n7367), .B1(n10157), .B2(n7368), .C1(
        n7366), .C2(n8885), .ZN(P1_U3334) );
  OAI222_X1 U9076 ( .A1(n8906), .A2(n8781), .B1(n8904), .B2(n7368), .C1(n9522), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  NAND2_X1 U9077 ( .A1(n9230), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7589) );
  INV_X1 U9078 ( .A(n7589), .ZN(n7663) );
  INV_X1 U9079 ( .A(n9278), .ZN(n7369) );
  INV_X1 U9080 ( .A(n9281), .ZN(n7656) );
  OAI22_X1 U9081 ( .A1(n7369), .A2(n9204), .B1(n7656), .B2(n9390), .ZN(n7460)
         );
  AOI22_X1 U9082 ( .A1(n9182), .A2(n7460), .B1(n10593), .B2(n10474), .ZN(n7375) );
  OAI21_X1 U9083 ( .B1(n7372), .B2(n7371), .A(n7370), .ZN(n7373) );
  NAND2_X1 U9084 ( .A1(n7373), .A2(n9212), .ZN(n7374) );
  OAI211_X1 U9085 ( .C1(n7663), .C2(n8132), .A(n7375), .B(n7374), .ZN(P2_U3224) );
  NOR2_X1 U9086 ( .A1(n7377), .A2(n7376), .ZN(n7378) );
  NAND2_X1 U9087 ( .A1(n7379), .A2(n7378), .ZN(n7455) );
  NAND2_X2 U9088 ( .A1(n7455), .A2(n9537), .ZN(n9540) );
  XNOR2_X1 U9089 ( .A(n7380), .B(n8943), .ZN(n10491) );
  INV_X1 U9090 ( .A(n8260), .ZN(n7381) );
  NAND2_X1 U9091 ( .A1(n10491), .A2(n7381), .ZN(n7388) );
  NAND3_X1 U9092 ( .A1(n7465), .A2(n8943), .A3(n9009), .ZN(n7382) );
  NAND2_X1 U9093 ( .A1(n7383), .A2(n7382), .ZN(n7386) );
  INV_X2 U9094 ( .A(n9553), .ZN(n9532) );
  INV_X1 U9095 ( .A(n9204), .ZN(n9386) );
  NAND2_X1 U9096 ( .A1(n9276), .A2(n9386), .ZN(n7385) );
  NAND2_X1 U9097 ( .A1(n9278), .A2(n9245), .ZN(n7384) );
  NAND2_X1 U9098 ( .A1(n7385), .A2(n7384), .ZN(n7413) );
  AOI21_X1 U9099 ( .B1(n7386), .B2(n9532), .A(n7413), .ZN(n7387) );
  AND2_X1 U9100 ( .A1(n7388), .A2(n7387), .ZN(n10493) );
  OR2_X1 U9101 ( .A1(n7389), .A2(n9522), .ZN(n7453) );
  INV_X1 U9102 ( .A(n7453), .ZN(n7390) );
  NAND2_X1 U9103 ( .A1(n9540), .A2(n7390), .ZN(n8043) );
  INV_X1 U9104 ( .A(n8043), .ZN(n10227) );
  NOR2_X2 U9105 ( .A1(n7455), .A2(n9565), .ZN(n9504) );
  OAI211_X1 U9106 ( .C1(n7472), .C2(n10489), .A(n7618), .B(n9541), .ZN(n10488)
         );
  INV_X1 U9107 ( .A(n10488), .ZN(n7392) );
  INV_X1 U9108 ( .A(n9537), .ZN(n10218) );
  INV_X1 U9109 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n8522) );
  AOI22_X1 U9110 ( .A1(n9504), .A2(n7392), .B1(n10218), .B2(n8522), .ZN(n7394)
         );
  NAND2_X1 U9111 ( .A1(n4499), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7393) );
  OAI211_X1 U9112 ( .C1(n9552), .C2(n10489), .A(n7394), .B(n7393), .ZN(n7395)
         );
  AOI21_X1 U9113 ( .B1(n10227), .B2(n10491), .A(n7395), .ZN(n7396) );
  OAI21_X1 U9114 ( .B1(n4499), .B2(n10493), .A(n7396), .ZN(P2_U3293) );
  NAND2_X1 U9115 ( .A1(n10404), .A2(n9825), .ZN(n7397) );
  AND2_X1 U9116 ( .A1(n7547), .A2(n9824), .ZN(n7399) );
  XNOR2_X1 U9117 ( .A(n7751), .B(n7750), .ZN(n10175) );
  INV_X1 U9118 ( .A(n7400), .ZN(n7401) );
  NAND2_X1 U9119 ( .A1(n10335), .A2(n7402), .ZN(n7404) );
  XNOR2_X1 U9120 ( .A(n7758), .B(n7750), .ZN(n7406) );
  AOI22_X1 U9121 ( .A1(n10054), .A2(n9824), .B1(n9822), .B2(n10056), .ZN(n7405) );
  OAI21_X1 U9122 ( .B1(n7406), .B2(n9988), .A(n7405), .ZN(n7407) );
  AOI21_X1 U9123 ( .B1(n10175), .B2(n10253), .A(n7407), .ZN(n10177) );
  INV_X1 U9124 ( .A(n7547), .ZN(n10415) );
  INV_X1 U9125 ( .A(n7752), .ZN(n10172) );
  NAND2_X1 U9126 ( .A1(n10329), .A2(n10172), .ZN(n10238) );
  OR2_X1 U9127 ( .A1(n10329), .A2(n10172), .ZN(n7408) );
  NAND2_X1 U9128 ( .A1(n10238), .A2(n7408), .ZN(n10173) );
  AOI22_X1 U9129 ( .A1(n10048), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n5066), .B2(
        n10345), .ZN(n7410) );
  NAND2_X1 U9130 ( .A1(n7752), .A2(n8238), .ZN(n7409) );
  OAI211_X1 U9131 ( .C1(n10173), .C2(n7774), .A(n7410), .B(n7409), .ZN(n7411)
         );
  AOI21_X1 U9132 ( .B1(n10175), .B2(n10332), .A(n7411), .ZN(n7412) );
  OAI21_X1 U9133 ( .B1(n10177), .B2(n10048), .A(n7412), .ZN(P1_U3281) );
  INV_X1 U9134 ( .A(n9230), .ZN(n9249) );
  AOI22_X1 U9135 ( .A1(n9182), .A2(n7413), .B1(P2_U3152), .B2(
        P2_REG3_REG_3__SCAN_IN), .ZN(n7414) );
  OAI21_X1 U9136 ( .B1(n9252), .B2(n10489), .A(n7414), .ZN(n7420) );
  INV_X1 U9137 ( .A(n7415), .ZN(n7416) );
  AOI211_X1 U9138 ( .C1(n7418), .C2(n7417), .A(n9240), .B(n7416), .ZN(n7419)
         );
  AOI211_X1 U9139 ( .C1(n8522), .C2(n9249), .A(n7420), .B(n7419), .ZN(n7421)
         );
  INV_X1 U9140 ( .A(n7421), .ZN(P2_U3220) );
  INV_X1 U9141 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7437) );
  INV_X1 U9142 ( .A(n7422), .ZN(n7428) );
  NOR2_X1 U9143 ( .A1(n7428), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7423) );
  INV_X1 U9144 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7597) );
  MUX2_X1 U9145 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n7597), .S(n7606), .Z(n7424)
         );
  OAI21_X1 U9146 ( .B1(n7425), .B2(n7423), .A(n7424), .ZN(n7602) );
  INV_X1 U9147 ( .A(n7602), .ZN(n7427) );
  NOR3_X1 U9148 ( .A1(n7425), .A2(n7424), .A3(n7423), .ZN(n7426) );
  OAI21_X1 U9149 ( .B1(n7427), .B2(n7426), .A(n10319), .ZN(n7436) );
  NOR2_X1 U9150 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6014), .ZN(n7795) );
  NAND2_X1 U9151 ( .A1(n7606), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7431) );
  OAI21_X1 U9152 ( .B1(n7606), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7431), .ZN(
        n7432) );
  AOI211_X1 U9153 ( .C1(n7433), .C2(n7432), .A(n7605), .B(n10313), .ZN(n7434)
         );
  AOI211_X1 U9154 ( .C1(n10310), .C2(n7606), .A(n7795), .B(n7434), .ZN(n7435)
         );
  OAI211_X1 U9155 ( .C1(n7437), .C2(n10305), .A(n7436), .B(n7435), .ZN(
        P1_U3253) );
  INV_X1 U9156 ( .A(n10524), .ZN(n10478) );
  NAND2_X1 U9157 ( .A1(n7438), .A2(n8940), .ZN(n7440) );
  NAND2_X1 U9158 ( .A1(n7440), .A2(n7439), .ZN(n7442) );
  XNOR2_X1 U9159 ( .A(n9275), .B(n7539), .ZN(n8948) );
  INV_X1 U9160 ( .A(n8948), .ZN(n7441) );
  XNOR2_X1 U9161 ( .A(n7442), .B(n7441), .ZN(n7485) );
  NAND2_X1 U9162 ( .A1(n7614), .A2(n8997), .ZN(n7444) );
  NAND2_X1 U9163 ( .A1(n7444), .A2(n7443), .ZN(n7445) );
  XNOR2_X1 U9164 ( .A(n7445), .B(n8948), .ZN(n7448) );
  NAND2_X1 U9165 ( .A1(n9276), .A2(n9245), .ZN(n7447) );
  NAND2_X1 U9166 ( .A1(n9274), .A2(n9386), .ZN(n7446) );
  NAND2_X1 U9167 ( .A1(n7447), .A2(n7446), .ZN(n7523) );
  AOI21_X1 U9168 ( .B1(n7448), .B2(n9532), .A(n7523), .ZN(n7478) );
  OAI21_X1 U9169 ( .B1(n7618), .B2(n9214), .A(n7524), .ZN(n7449) );
  NAND3_X1 U9170 ( .A1(n7449), .A2(n9541), .A3(n7571), .ZN(n7479) );
  OAI211_X1 U9171 ( .C1(n10478), .C2(n7485), .A(n7478), .B(n7479), .ZN(n7541)
         );
  OAI22_X1 U9172 ( .A1(n9640), .A2(n7539), .B1(n10541), .B2(n5244), .ZN(n7450)
         );
  AOI21_X1 U9173 ( .B1(n7541), .B2(n10541), .A(n7450), .ZN(n7451) );
  INV_X1 U9174 ( .A(n7451), .ZN(P2_U3525) );
  XOR2_X1 U9175 ( .A(n7452), .B(n8939), .Z(n10479) );
  NAND2_X1 U9176 ( .A1(n8260), .A2(n7453), .ZN(n7454) );
  NAND2_X1 U9177 ( .A1(n9540), .A2(n7454), .ZN(n9536) );
  INV_X1 U9178 ( .A(n7455), .ZN(n7456) );
  NAND2_X1 U9179 ( .A1(n7456), .A2(n7521), .ZN(n8037) );
  NOR2_X1 U9180 ( .A1(n7457), .A2(n7655), .ZN(n10472) );
  OR2_X1 U9181 ( .A1(n10472), .A2(n10471), .ZN(n7458) );
  OAI22_X1 U9182 ( .A1(n8037), .A2(n7458), .B1(n8132), .B2(n9537), .ZN(n7459)
         );
  AOI21_X1 U9183 ( .B1(n10221), .B2(n10474), .A(n7459), .ZN(n7463) );
  XNOR2_X1 U9184 ( .A(n8939), .B(n7498), .ZN(n7461) );
  AOI21_X1 U9185 ( .B1(n9532), .B2(n7461), .A(n7460), .ZN(n10477) );
  INV_X1 U9186 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7682) );
  MUX2_X1 U9187 ( .A(n10477), .B(n7682), .S(n4499), .Z(n7462) );
  OAI211_X1 U9188 ( .C1(n10479), .C2(n9536), .A(n7463), .B(n7462), .ZN(
        P2_U3295) );
  XNOR2_X1 U9189 ( .A(n7464), .B(n7467), .ZN(n10481) );
  OAI21_X1 U9190 ( .B1(n7467), .B2(n7466), .A(n7465), .ZN(n7468) );
  NAND2_X1 U9191 ( .A1(n7468), .A2(n9532), .ZN(n7470) );
  AOI22_X1 U9192 ( .A1(n9245), .A2(n9279), .B1(n9277), .B2(n9386), .ZN(n7469)
         );
  NAND2_X1 U9193 ( .A1(n7470), .A2(n7469), .ZN(n10484) );
  MUX2_X1 U9194 ( .A(n10484), .B(P2_REG2_REG_2__SCAN_IN), .S(n4499), .Z(n7471)
         );
  INV_X1 U9195 ( .A(n7471), .ZN(n7477) );
  INV_X1 U9196 ( .A(n7472), .ZN(n7473) );
  OAI21_X1 U9197 ( .B1(n10482), .B2(n10471), .A(n7473), .ZN(n10483) );
  OAI22_X1 U9198 ( .A1(n8037), .A2(n10483), .B1(n7474), .B2(n9537), .ZN(n7475)
         );
  AOI21_X1 U9199 ( .B1(n10221), .B2(n7588), .A(n7475), .ZN(n7476) );
  OAI211_X1 U9200 ( .C1(n10481), .C2(n9536), .A(n7477), .B(n7476), .ZN(
        P2_U3294) );
  OAI21_X1 U9201 ( .B1(n9565), .B2(n7479), .A(n7478), .ZN(n7480) );
  NAND2_X1 U9202 ( .A1(n7480), .A2(n9540), .ZN(n7484) );
  INV_X1 U9203 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7481) );
  OAI22_X1 U9204 ( .A1(n9540), .A2(n7481), .B1(n7527), .B2(n9537), .ZN(n7482)
         );
  AOI21_X1 U9205 ( .B1(n10221), .B2(n7524), .A(n7482), .ZN(n7483) );
  OAI211_X1 U9206 ( .C1(n7485), .C2(n9536), .A(n7484), .B(n7483), .ZN(P2_U3291) );
  NAND2_X1 U9207 ( .A1(n4508), .A2(n7486), .ZN(n7488) );
  XNOR2_X1 U9208 ( .A(n7488), .B(n7487), .ZN(n7496) );
  NAND2_X1 U9209 ( .A1(n9792), .A2(n10404), .ZN(n7494) );
  AOI21_X1 U9210 ( .B1(n9786), .B2(n9826), .A(n7489), .ZN(n7493) );
  NAND2_X1 U9211 ( .A1(n9809), .A2(n7490), .ZN(n7492) );
  NAND2_X1 U9212 ( .A1(n9768), .A2(n9824), .ZN(n7491) );
  NAND4_X1 U9213 ( .A1(n7494), .A2(n7493), .A3(n7492), .A4(n7491), .ZN(n7495)
         );
  AOI21_X1 U9214 ( .B1(n7496), .B2(n9802), .A(n7495), .ZN(n7497) );
  INV_X1 U9215 ( .A(n7497), .ZN(P1_U3219) );
  NAND2_X1 U9216 ( .A1(n9281), .A2(n7655), .ZN(n9006) );
  NAND2_X1 U9217 ( .A1(n7498), .A2(n9006), .ZN(n10468) );
  AND2_X1 U9218 ( .A1(n9279), .A2(n9386), .ZN(n7499) );
  AOI21_X1 U9219 ( .B1(n10468), .B2(n9532), .A(n7499), .ZN(n10470) );
  OAI22_X1 U9220 ( .A1(n4499), .A2(n10470), .B1(n7662), .B2(n9537), .ZN(n7502)
         );
  INV_X1 U9221 ( .A(n10468), .ZN(n7500) );
  NOR2_X1 U9222 ( .A1(n9536), .A2(n7500), .ZN(n7501) );
  AOI211_X1 U9223 ( .C1(n4499), .C2(P2_REG2_REG_0__SCAN_IN), .A(n7502), .B(
        n7501), .ZN(n7505) );
  INV_X1 U9224 ( .A(n8037), .ZN(n7503) );
  OAI21_X1 U9225 ( .B1(n10221), .B2(n7503), .A(n10466), .ZN(n7504) );
  NAND2_X1 U9226 ( .A1(n7505), .A2(n7504), .ZN(P2_U3296) );
  OAI21_X1 U9227 ( .B1(n7507), .B2(n9016), .A(n7506), .ZN(n7630) );
  INV_X1 U9228 ( .A(n7630), .ZN(n7520) );
  AND2_X1 U9229 ( .A1(n7509), .A2(n7508), .ZN(n7736) );
  NAND2_X1 U9230 ( .A1(n7736), .A2(n8945), .ZN(n7510) );
  NAND2_X1 U9231 ( .A1(n7510), .A2(n9017), .ZN(n7511) );
  XNOR2_X1 U9232 ( .A(n7511), .B(n9016), .ZN(n7512) );
  AOI22_X1 U9233 ( .A1(n9386), .A2(n9272), .B1(n9274), .B2(n9245), .ZN(n7649)
         );
  OAI21_X1 U9234 ( .B1(n7512), .B2(n9553), .A(n7649), .ZN(n7628) );
  NAND2_X1 U9235 ( .A1(n7628), .A2(n9540), .ZN(n7519) );
  INV_X1 U9236 ( .A(n7513), .ZN(n7573) );
  INV_X1 U9237 ( .A(n7744), .ZN(n7514) );
  AOI211_X1 U9238 ( .C1(n7651), .C2(n7573), .A(n10520), .B(n7514), .ZN(n7629)
         );
  NOR2_X1 U9239 ( .A1(n9552), .A2(n7633), .ZN(n7517) );
  INV_X1 U9240 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7515) );
  OAI22_X1 U9241 ( .A1(n9540), .A2(n7515), .B1(n7654), .B2(n9537), .ZN(n7516)
         );
  AOI211_X1 U9242 ( .C1(n7629), .C2(n9504), .A(n7517), .B(n7516), .ZN(n7518)
         );
  OAI211_X1 U9243 ( .C1(n7520), .C2(n9536), .A(n7519), .B(n7518), .ZN(P2_U3289) );
  INV_X1 U9244 ( .A(n7560), .ZN(n7536) );
  AOI22_X1 U9245 ( .A1(n9235), .A2(n9275), .B1(n9212), .B2(n7522), .ZN(n7535)
         );
  AOI22_X1 U9246 ( .A1(n9182), .A2(n7523), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        P2_U3152), .ZN(n7526) );
  NAND2_X1 U9247 ( .A1(n10593), .A2(n7524), .ZN(n7525) );
  OAI211_X1 U9248 ( .C1(n9230), .C2(n7527), .A(n7526), .B(n7525), .ZN(n7528)
         );
  INV_X1 U9249 ( .A(n7528), .ZN(n7534) );
  INV_X1 U9250 ( .A(n7529), .ZN(n7531) );
  OAI211_X1 U9251 ( .C1(n7532), .C2(n7531), .A(n7530), .B(n9212), .ZN(n7533)
         );
  OAI211_X1 U9252 ( .C1(n7536), .C2(n7535), .A(n7534), .B(n7533), .ZN(P2_U3229) );
  INV_X1 U9253 ( .A(n7537), .ZN(n7556) );
  OAI222_X1 U9254 ( .A1(n8904), .A2(n7556), .B1(P2_U3152), .B2(n8942), .C1(
        n7538), .C2(n8906), .ZN(P2_U3338) );
  OAI22_X1 U9255 ( .A1(n9692), .A2(n7539), .B1(n10528), .B2(n5247), .ZN(n7540)
         );
  AOI21_X1 U9256 ( .B1(n7541), .B2(n10528), .A(n7540), .ZN(n7542) );
  INV_X1 U9257 ( .A(n7542), .ZN(P2_U3466) );
  NAND2_X1 U9258 ( .A1(n7543), .A2(n7544), .ZN(n7545) );
  AOI21_X1 U9259 ( .B1(n7546), .B2(n7545), .A(n9795), .ZN(n7554) );
  NAND2_X1 U9260 ( .A1(n7547), .A2(n9792), .ZN(n7552) );
  AOI21_X1 U9261 ( .B1(n9786), .B2(n9825), .A(n7548), .ZN(n7551) );
  NAND2_X1 U9262 ( .A1(n9809), .A2(n10346), .ZN(n7550) );
  INV_X1 U9263 ( .A(n10339), .ZN(n9823) );
  NAND2_X1 U9264 ( .A1(n9768), .A2(n9823), .ZN(n7549) );
  NAND4_X1 U9265 ( .A1(n7552), .A2(n7551), .A3(n7550), .A4(n7549), .ZN(n7553)
         );
  OR2_X1 U9266 ( .A1(n7554), .A2(n7553), .ZN(P1_U3229) );
  OAI222_X1 U9267 ( .A1(n7557), .A2(P1_U3084), .B1(n10157), .B2(n7556), .C1(
        n7555), .C2(n8885), .ZN(P1_U3333) );
  OAI21_X1 U9268 ( .B1(n7560), .B2(n7559), .A(n7558), .ZN(n7566) );
  NAND2_X1 U9269 ( .A1(n9273), .A2(n9386), .ZN(n7562) );
  NAND2_X1 U9270 ( .A1(n9275), .A2(n9245), .ZN(n7561) );
  NAND2_X1 U9271 ( .A1(n7562), .A2(n7561), .ZN(n7577) );
  AND2_X1 U9272 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n7885) );
  AOI21_X1 U9273 ( .B1(n9182), .B2(n7577), .A(n7885), .ZN(n7564) );
  NAND2_X1 U9274 ( .A1(n10593), .A2(n7581), .ZN(n7563) );
  OAI211_X1 U9275 ( .C1(n9230), .C2(n7574), .A(n7564), .B(n7563), .ZN(n7565)
         );
  AOI21_X1 U9276 ( .B1(n7566), .B2(n9212), .A(n7565), .ZN(n7567) );
  INV_X1 U9277 ( .A(n7567), .ZN(P2_U3241) );
  INV_X1 U9278 ( .A(n7568), .ZN(n7626) );
  INV_X1 U9279 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7569) );
  OAI222_X1 U9280 ( .A1(n8904), .A2(n7626), .B1(P2_U3152), .B2(n8931), .C1(
        n7569), .C2(n8906), .ZN(P2_U3337) );
  XNOR2_X1 U9281 ( .A(n7570), .B(n8945), .ZN(n10503) );
  INV_X1 U9282 ( .A(n10503), .ZN(n7583) );
  AOI21_X1 U9283 ( .B1(n7571), .B2(n7581), .A(n10520), .ZN(n7572) );
  NAND2_X1 U9284 ( .A1(n7573), .A2(n7572), .ZN(n10499) );
  INV_X1 U9285 ( .A(n9504), .ZN(n10224) );
  NOR2_X1 U9286 ( .A1(n9537), .A2(n7574), .ZN(n7575) );
  AOI21_X1 U9287 ( .B1(n4499), .B2(P2_REG2_REG_6__SCAN_IN), .A(n7575), .ZN(
        n7576) );
  OAI21_X1 U9288 ( .B1(n10499), .B2(n10224), .A(n7576), .ZN(n7580) );
  XNOR2_X1 U9289 ( .A(n7736), .B(n8945), .ZN(n7578) );
  AOI21_X1 U9290 ( .B1(n7578), .B2(n9532), .A(n7577), .ZN(n10500) );
  NOR2_X1 U9291 ( .A1(n10500), .A2(n4499), .ZN(n7579) );
  AOI211_X1 U9292 ( .C1(n10221), .C2(n7581), .A(n7580), .B(n7579), .ZN(n7582)
         );
  OAI21_X1 U9293 ( .B1(n9536), .B2(n7583), .A(n7582), .ZN(P2_U3290) );
  INV_X1 U9294 ( .A(n7584), .ZN(n7585) );
  AOI22_X1 U9295 ( .A1(n9235), .A2(n9279), .B1(n9212), .B2(n7585), .ZN(n7587)
         );
  NOR2_X1 U9296 ( .A1(n7587), .A2(n7586), .ZN(n7594) );
  NAND2_X1 U9297 ( .A1(n9182), .A2(n9386), .ZN(n9218) );
  AND2_X1 U9298 ( .A1(n9182), .A2(n9245), .ZN(n9224) );
  AOI22_X1 U9299 ( .A1(n9224), .A2(n9279), .B1(n7588), .B2(n10593), .ZN(n7591)
         );
  NAND2_X1 U9300 ( .A1(n7589), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n7590) );
  OAI211_X1 U9301 ( .C1(n7592), .C2(n9218), .A(n7591), .B(n7590), .ZN(n7593)
         );
  AOI21_X1 U9302 ( .B1(n7594), .B2(n7370), .A(n7593), .ZN(n7595) );
  OAI21_X1 U9303 ( .B1(n7596), .B2(n9240), .A(n7595), .ZN(P2_U3239) );
  NAND2_X1 U9304 ( .A1(n7598), .A2(n7597), .ZN(n7600) );
  INV_X1 U9305 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7599) );
  MUX2_X1 U9306 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n7599), .S(n8009), .Z(n7601)
         );
  AOI21_X1 U9307 ( .B1(n7602), .B2(n7600), .A(n7601), .ZN(n8008) );
  INV_X1 U9308 ( .A(n8008), .ZN(n7604) );
  NAND3_X1 U9309 ( .A1(n7602), .A2(n7601), .A3(n7600), .ZN(n7603) );
  AOI21_X1 U9310 ( .B1(n7604), .B2(n7603), .A(n9895), .ZN(n7613) );
  XOR2_X1 U9311 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n8009), .Z(n7607) );
  AOI211_X1 U9312 ( .C1(n7608), .C2(n7607), .A(n10313), .B(n8014), .ZN(n7612)
         );
  INV_X1 U9313 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7610) );
  INV_X1 U9314 ( .A(n8009), .ZN(n8015) );
  NOR2_X1 U9315 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8697), .ZN(n7850) );
  AOI21_X1 U9316 ( .B1(n10310), .B2(n8015), .A(n7850), .ZN(n7609) );
  OAI21_X1 U9317 ( .B1(n10305), .B2(n7610), .A(n7609), .ZN(n7611) );
  OR3_X1 U9318 ( .A1(n7613), .A2(n7612), .A3(n7611), .ZN(P1_U3254) );
  XNOR2_X1 U9319 ( .A(n7614), .B(n8940), .ZN(n7615) );
  NAND2_X1 U9320 ( .A1(n7615), .A2(n9532), .ZN(n7617) );
  AOI22_X1 U9321 ( .A1(n9245), .A2(n9277), .B1(n9275), .B2(n9386), .ZN(n7616)
         );
  NAND2_X1 U9322 ( .A1(n7617), .A2(n7616), .ZN(n10496) );
  INV_X1 U9323 ( .A(n10496), .ZN(n7624) );
  INV_X1 U9324 ( .A(n9536), .ZN(n9465) );
  XNOR2_X1 U9325 ( .A(n7438), .B(n8940), .ZN(n10498) );
  XNOR2_X1 U9326 ( .A(n7618), .B(n9214), .ZN(n10495) );
  NAND2_X1 U9327 ( .A1(n10221), .A2(n9214), .ZN(n7621) );
  INV_X1 U9328 ( .A(n7619), .ZN(n9220) );
  AOI22_X1 U9329 ( .A1(n4499), .A2(P2_REG2_REG_4__SCAN_IN), .B1(n9220), .B2(
        n10218), .ZN(n7620) );
  OAI211_X1 U9330 ( .C1(n8037), .C2(n10495), .A(n7621), .B(n7620), .ZN(n7622)
         );
  AOI21_X1 U9331 ( .B1(n9465), .B2(n10498), .A(n7622), .ZN(n7623) );
  OAI21_X1 U9332 ( .B1(n7624), .B2(n4499), .A(n7623), .ZN(P2_U3292) );
  INV_X1 U9333 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7625) );
  OAI222_X1 U9334 ( .A1(n7627), .A2(P1_U3084), .B1(n10157), .B2(n7626), .C1(
        n7625), .C2(n8885), .ZN(P1_U3332) );
  AOI211_X1 U9335 ( .C1(n10524), .C2(n7630), .A(n7629), .B(n7628), .ZN(n7636)
         );
  OAI22_X1 U9336 ( .A1(n9640), .A2(n7633), .B1(n10541), .B2(n7701), .ZN(n7631)
         );
  INV_X1 U9337 ( .A(n7631), .ZN(n7632) );
  OAI21_X1 U9338 ( .B1(n7636), .B2(n10539), .A(n7632), .ZN(P2_U3527) );
  OAI22_X1 U9339 ( .A1(n9692), .A2(n7633), .B1(n10528), .B2(n5278), .ZN(n7634)
         );
  INV_X1 U9340 ( .A(n7634), .ZN(n7635) );
  OAI21_X1 U9341 ( .B1(n7636), .B2(n10526), .A(n7635), .ZN(P2_U3472) );
  OAI21_X1 U9342 ( .B1(n7638), .B2(n7637), .A(n7665), .ZN(n7639) );
  NAND2_X1 U9343 ( .A1(n7639), .A2(n9802), .ZN(n7644) );
  AOI21_X1 U9344 ( .B1(n9786), .B2(n9824), .A(n7640), .ZN(n7641) );
  OAI21_X1 U9345 ( .B1(n7814), .B2(n9806), .A(n7641), .ZN(n7642) );
  AOI21_X1 U9346 ( .B1(n5066), .B2(n9809), .A(n7642), .ZN(n7643) );
  OAI211_X1 U9347 ( .C1(n10172), .C2(n9812), .A(n7644), .B(n7643), .ZN(
        P1_U3215) );
  AOI21_X1 U9348 ( .B1(n7646), .B2(n7645), .A(n9240), .ZN(n7647) );
  OR2_X1 U9349 ( .A1(n7646), .A2(n7645), .ZN(n7778) );
  NAND2_X1 U9350 ( .A1(n7647), .A2(n7778), .ZN(n7653) );
  INV_X1 U9351 ( .A(n9182), .ZN(n9247) );
  OAI22_X1 U9352 ( .A1(n9247), .A2(n7649), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7648), .ZN(n7650) );
  AOI21_X1 U9353 ( .B1(n7651), .B2(n10593), .A(n7650), .ZN(n7652) );
  OAI211_X1 U9354 ( .C1(n9230), .C2(n7654), .A(n7653), .B(n7652), .ZN(P2_U3215) );
  INV_X1 U9355 ( .A(n9235), .ZN(n9223) );
  OAI22_X1 U9356 ( .A1(n9223), .A2(n7656), .B1(n7655), .B2(n9240), .ZN(n7658)
         );
  NAND2_X1 U9357 ( .A1(n7658), .A2(n7657), .ZN(n7661) );
  INV_X1 U9358 ( .A(n9218), .ZN(n7659) );
  AOI22_X1 U9359 ( .A1(n7659), .A2(n9279), .B1(n10466), .B2(n10593), .ZN(n7660) );
  OAI211_X1 U9360 ( .C1(n7663), .C2(n7662), .A(n7661), .B(n7660), .ZN(P2_U3234) );
  INV_X1 U9361 ( .A(n10237), .ZN(n10277) );
  AND2_X1 U9362 ( .A1(n7665), .A2(n7664), .ZN(n7668) );
  OAI211_X1 U9363 ( .C1(n7668), .C2(n7667), .A(n9802), .B(n7666), .ZN(n7674)
         );
  INV_X1 U9364 ( .A(n7669), .ZN(n7670) );
  AOI21_X1 U9365 ( .B1(n9786), .B2(n9823), .A(n7670), .ZN(n7671) );
  OAI21_X1 U9366 ( .B1(n10248), .B2(n9806), .A(n7671), .ZN(n7672) );
  AOI21_X1 U9367 ( .B1(n10254), .B2(n9809), .A(n7672), .ZN(n7673) );
  OAI211_X1 U9368 ( .C1(n10277), .C2(n9812), .A(n7674), .B(n7673), .ZN(
        P1_U3234) );
  OR2_X1 U9369 ( .A1(n5799), .A2(P2_U3152), .ZN(n8377) );
  OAI21_X1 U9370 ( .B1(n7675), .B2(n8377), .A(n9134), .ZN(n7676) );
  INV_X1 U9371 ( .A(n7676), .ZN(n7677) );
  NAND2_X1 U9372 ( .A1(n7678), .A2(n7677), .ZN(n7725) );
  NAND2_X1 U9373 ( .A1(n7725), .A2(n7723), .ZN(n7679) );
  NAND2_X1 U9374 ( .A1(n7679), .A2(n9280), .ZN(n7726) );
  INV_X1 U9375 ( .A(n7726), .ZN(n7680) );
  NOR3_X2 U9376 ( .A1(n7680), .A2(n9129), .A3(n5799), .ZN(n10440) );
  NAND2_X1 U9377 ( .A1(n8203), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7681) );
  OAI21_X1 U9378 ( .B1(n8203), .B2(P2_REG2_REG_12__SCAN_IN), .A(n7681), .ZN(
        n8199) );
  XNOR2_X1 U9379 ( .A(n7709), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n8181) );
  MUX2_X1 U9380 ( .A(n7682), .B(P2_REG2_REG_1__SCAN_IN), .S(n7704), .Z(n8130)
         );
  NAND2_X1 U9381 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n8131) );
  NOR2_X1 U9382 ( .A1(n8130), .A2(n8131), .ZN(n8129) );
  AOI21_X1 U9383 ( .B1(n7704), .B2(P2_REG2_REG_1__SCAN_IN), .A(n8129), .ZN(
        n10162) );
  INV_X1 U9384 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7683) );
  MUX2_X1 U9385 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n7683), .S(n10164), .Z(n7684)
         );
  INV_X1 U9386 ( .A(n7684), .ZN(n10161) );
  NOR2_X1 U9387 ( .A1(n10162), .A2(n10161), .ZN(n10160) );
  AOI21_X1 U9388 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n10164), .A(n10160), .ZN(
        n8095) );
  NAND2_X1 U9389 ( .A1(n7708), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7685) );
  OAI21_X1 U9390 ( .B1(n7708), .B2(P2_REG2_REG_3__SCAN_IN), .A(n7685), .ZN(
        n8094) );
  NOR2_X1 U9391 ( .A1(n8095), .A2(n8094), .ZN(n8093) );
  NAND2_X1 U9392 ( .A1(n8216), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7686) );
  OAI21_X1 U9393 ( .B1(n8216), .B2(P2_REG2_REG_5__SCAN_IN), .A(n7686), .ZN(
        n8212) );
  AOI21_X1 U9394 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n8216), .A(n8211), .ZN(
        n7887) );
  XNOR2_X1 U9395 ( .A(n7712), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n7886) );
  OR2_X1 U9396 ( .A1(n7700), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7688) );
  NAND2_X1 U9397 ( .A1(n7700), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7687) );
  NAND2_X1 U9398 ( .A1(n7688), .A2(n7687), .ZN(n8118) );
  AOI21_X1 U9399 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n7700), .A(n8117), .ZN(
        n7689) );
  INV_X1 U9400 ( .A(n7689), .ZN(n7876) );
  MUX2_X1 U9401 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n7743), .S(n7715), .Z(n7877)
         );
  NAND2_X1 U9402 ( .A1(n7876), .A2(n7877), .ZN(n7875) );
  OAI21_X1 U9403 ( .B1(n7743), .B2(n7880), .A(n7875), .ZN(n7865) );
  NAND2_X1 U9404 ( .A1(n7716), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7690) );
  OAI21_X1 U9405 ( .B1(n7716), .B2(P2_REG2_REG_9__SCAN_IN), .A(n7690), .ZN(
        n7691) );
  INV_X1 U9406 ( .A(n7691), .ZN(n7866) );
  NAND2_X1 U9407 ( .A1(n7865), .A2(n7866), .ZN(n7864) );
  NAND2_X1 U9408 ( .A1(n7698), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7692) );
  OAI21_X1 U9409 ( .B1(n7698), .B2(P2_REG2_REG_10__SCAN_IN), .A(n7692), .ZN(
        n8106) );
  NOR2_X1 U9410 ( .A1(n9287), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7693) );
  AOI21_X1 U9411 ( .B1(n9287), .B2(P2_REG2_REG_11__SCAN_IN), .A(n7693), .ZN(
        n9284) );
  NAND2_X1 U9412 ( .A1(n9283), .A2(n9284), .ZN(n9282) );
  OAI21_X1 U9413 ( .B1(n9287), .B2(P2_REG2_REG_11__SCAN_IN), .A(n9282), .ZN(
        n8200) );
  NOR2_X1 U9414 ( .A1(n8199), .A2(n8200), .ZN(n8198) );
  NOR2_X1 U9415 ( .A1(n7835), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7694) );
  AOI21_X1 U9416 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n7835), .A(n7694), .ZN(
        n7695) );
  OAI21_X1 U9417 ( .B1(n7696), .B2(n7695), .A(n7834), .ZN(n7731) );
  MUX2_X1 U9418 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n7697), .S(n9287), .Z(n9289)
         );
  MUX2_X1 U9419 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n7699), .S(n7698), .Z(n8109)
         );
  INV_X1 U9420 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n8062) );
  NAND2_X1 U9421 ( .A1(n7700), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7714) );
  MUX2_X1 U9422 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n7701), .S(n7700), .Z(n8123)
         );
  NAND2_X1 U9423 ( .A1(n8216), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7711) );
  INV_X1 U9424 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10533) );
  MUX2_X1 U9425 ( .A(n10533), .B(P2_REG1_REG_4__SCAN_IN), .S(n7709), .Z(n8185)
         );
  MUX2_X1 U9426 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n7702), .S(n7708), .Z(n8098)
         );
  MUX2_X1 U9427 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n7703), .S(n10164), .Z(n10167) );
  MUX2_X1 U9428 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n7705), .S(n7704), .Z(n8136)
         );
  AND2_X1 U9429 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(
        n8137) );
  NAND2_X1 U9430 ( .A1(n8136), .A2(n8137), .ZN(n8135) );
  OAI21_X1 U9431 ( .B1(n8140), .B2(n7705), .A(n8135), .ZN(n10168) );
  NAND2_X1 U9432 ( .A1(n10167), .A2(n10168), .ZN(n10166) );
  OAI21_X1 U9433 ( .B1(n7703), .B2(n7706), .A(n10166), .ZN(n8099) );
  NAND2_X1 U9434 ( .A1(n8098), .A2(n8099), .ZN(n8097) );
  INV_X1 U9435 ( .A(n8097), .ZN(n7707) );
  MUX2_X1 U9436 ( .A(n5244), .B(P2_REG1_REG_5__SCAN_IN), .S(n8216), .Z(n8205)
         );
  AND2_X1 U9437 ( .A1(n7711), .A2(n7710), .ZN(n7883) );
  MUX2_X1 U9438 ( .A(n7713), .B(P2_REG1_REG_6__SCAN_IN), .S(n7712), .Z(n7882)
         );
  AND2_X1 U9439 ( .A1(n7714), .A2(n8121), .ZN(n7872) );
  INV_X1 U9440 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10536) );
  MUX2_X1 U9441 ( .A(n10536), .B(P2_REG1_REG_8__SCAN_IN), .S(n7715), .Z(n7871)
         );
  NAND2_X1 U9442 ( .A1(n7715), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7858) );
  MUX2_X1 U9443 ( .A(n8062), .B(P2_REG1_REG_9__SCAN_IN), .S(n7716), .Z(n7857)
         );
  OAI21_X1 U9444 ( .B1(n8062), .B2(n7869), .A(n7717), .ZN(n8110) );
  NAND2_X1 U9445 ( .A1(n8109), .A2(n8110), .ZN(n8108) );
  OAI21_X1 U9446 ( .B1(n8114), .B2(n7699), .A(n8108), .ZN(n9290) );
  NAND2_X1 U9447 ( .A1(n9289), .A2(n9290), .ZN(n9288) );
  OAI21_X1 U9448 ( .B1(n7718), .B2(n7697), .A(n9288), .ZN(n8193) );
  MUX2_X1 U9449 ( .A(n7719), .B(P2_REG1_REG_12__SCAN_IN), .S(n8203), .Z(n8194)
         );
  NOR2_X1 U9450 ( .A1(n8193), .A2(n8194), .ZN(n8192) );
  AOI21_X1 U9451 ( .B1(n7720), .B2(n7719), .A(n8192), .ZN(n7722) );
  AOI22_X1 U9452 ( .A1(n7835), .A2(n5443), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n7831), .ZN(n7721) );
  AOI21_X1 U9453 ( .B1(n7722), .B2(n7721), .A(n7830), .ZN(n7729) );
  AND2_X1 U9454 ( .A1(n7723), .A2(n9129), .ZN(n7724) );
  NAND2_X1 U9455 ( .A1(n7725), .A2(n7724), .ZN(n10444) );
  AND2_X1 U9456 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8055) );
  AOI21_X1 U9457 ( .B1(n10441), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n8055), .ZN(
        n7728) );
  NAND2_X1 U9458 ( .A1(n7726), .A2(n5799), .ZN(n10443) );
  INV_X1 U9459 ( .A(n10443), .ZN(n10165) );
  NAND2_X1 U9460 ( .A1(n10165), .A2(n7835), .ZN(n7727) );
  OAI211_X1 U9461 ( .C1(n7729), .C2(n10444), .A(n7728), .B(n7727), .ZN(n7730)
         );
  AOI21_X1 U9462 ( .B1(n10440), .B2(n7731), .A(n7730), .ZN(n7732) );
  INV_X1 U9463 ( .A(n7732), .ZN(P2_U3258) );
  NAND2_X1 U9464 ( .A1(n7733), .A2(n9021), .ZN(n7734) );
  NAND2_X1 U9465 ( .A1(n7895), .A2(n7734), .ZN(n10504) );
  AOI22_X1 U9466 ( .A1(n9271), .A2(n9386), .B1(n9245), .B2(n9273), .ZN(n7742)
         );
  NAND2_X1 U9467 ( .A1(n7736), .A2(n7735), .ZN(n7738) );
  NAND2_X1 U9468 ( .A1(n7738), .A2(n7737), .ZN(n7739) );
  XNOR2_X1 U9469 ( .A(n7739), .B(n9021), .ZN(n7740) );
  NAND2_X1 U9470 ( .A1(n7740), .A2(n9532), .ZN(n7741) );
  OAI211_X1 U9471 ( .C1(n10504), .C2(n8260), .A(n7742), .B(n7741), .ZN(n10508)
         );
  NAND2_X1 U9472 ( .A1(n10508), .A2(n9540), .ZN(n7749) );
  OAI22_X1 U9473 ( .A1(n9540), .A2(n7743), .B1(n7785), .B2(n9537), .ZN(n7747)
         );
  NAND2_X1 U9474 ( .A1(n7744), .A2(n10505), .ZN(n7745) );
  NAND2_X1 U9475 ( .A1(n4514), .A2(n7745), .ZN(n10507) );
  NOR2_X1 U9476 ( .A1(n10507), .A2(n8037), .ZN(n7746) );
  AOI211_X1 U9477 ( .C1(n10221), .C2(n10505), .A(n7747), .B(n7746), .ZN(n7748)
         );
  OAI211_X1 U9478 ( .C1(n10504), .C2(n8043), .A(n7749), .B(n7748), .ZN(
        P2_U3288) );
  NAND2_X1 U9479 ( .A1(n7751), .A2(n7750), .ZN(n7754) );
  OR2_X1 U9480 ( .A1(n7752), .A2(n9823), .ZN(n7753) );
  NOR2_X1 U9481 ( .A1(n10237), .A2(n9822), .ZN(n7756) );
  NAND2_X1 U9482 ( .A1(n10237), .A2(n9822), .ZN(n7755) );
  INV_X1 U9483 ( .A(n10248), .ZN(n9821) );
  XNOR2_X1 U9484 ( .A(n7918), .B(n4763), .ZN(n10274) );
  INV_X1 U9485 ( .A(n10242), .ZN(n7759) );
  NOR2_X1 U9486 ( .A1(n10244), .A2(n7759), .ZN(n7760) );
  INV_X1 U9487 ( .A(n7761), .ZN(n7762) );
  NAND2_X1 U9488 ( .A1(n7764), .A2(n7763), .ZN(n7765) );
  AND2_X1 U9489 ( .A1(n7765), .A2(n7917), .ZN(n7766) );
  OAI21_X1 U9490 ( .B1(n7926), .B2(n7766), .A(n10343), .ZN(n7768) );
  AOI22_X1 U9491 ( .A1(n9821), .A2(n10054), .B1(n10056), .B2(n9819), .ZN(n7767) );
  NAND2_X1 U9492 ( .A1(n7768), .A2(n7767), .ZN(n7769) );
  AOI21_X1 U9493 ( .B1(n10274), .B2(n10253), .A(n7769), .ZN(n10276) );
  INV_X1 U9494 ( .A(n7921), .ZN(n7771) );
  NAND2_X1 U9495 ( .A1(n7820), .A2(n10270), .ZN(n7770) );
  NAND2_X1 U9496 ( .A1(n7771), .A2(n7770), .ZN(n10272) );
  AOI22_X1 U9497 ( .A1(n10048), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7851), .B2(
        n10345), .ZN(n7773) );
  NAND2_X1 U9498 ( .A1(n10270), .A2(n8238), .ZN(n7772) );
  OAI211_X1 U9499 ( .C1(n10272), .C2(n7774), .A(n7773), .B(n7772), .ZN(n7775)
         );
  AOI21_X1 U9500 ( .B1(n10274), .B2(n10332), .A(n7775), .ZN(n7776) );
  OAI21_X1 U9501 ( .B1(n10276), .B2(n10048), .A(n7776), .ZN(P1_U3278) );
  AOI21_X1 U9502 ( .B1(n7778), .B2(n7777), .A(n9240), .ZN(n7784) );
  INV_X1 U9503 ( .A(n9273), .ZN(n7779) );
  NOR3_X1 U9504 ( .A1(n9223), .A2(n7780), .A3(n7779), .ZN(n7783) );
  AND2_X1 U9505 ( .A1(n7782), .A2(n7781), .ZN(n8888) );
  OAI21_X1 U9506 ( .B1(n7784), .B2(n7783), .A(n8888), .ZN(n7790) );
  AOI22_X1 U9507 ( .A1(n9224), .A2(n9273), .B1(P2_REG3_REG_8__SCAN_IN), .B2(
        P2_U3152), .ZN(n7787) );
  OR2_X1 U9508 ( .A1(n9230), .A2(n7785), .ZN(n7786) );
  OAI211_X1 U9509 ( .C1(n7808), .C2(n9218), .A(n7787), .B(n7786), .ZN(n7788)
         );
  AOI21_X1 U9510 ( .B1(n10505), .B2(n10593), .A(n7788), .ZN(n7789) );
  NAND2_X1 U9511 ( .A1(n7790), .A2(n7789), .ZN(P2_U3223) );
  NAND2_X1 U9512 ( .A1(n7792), .A2(n7791), .ZN(n7794) );
  XOR2_X1 U9513 ( .A(n7794), .B(n7793), .Z(n7800) );
  INV_X1 U9514 ( .A(n7928), .ZN(n9820) );
  AOI21_X1 U9515 ( .B1(n9768), .B2(n9820), .A(n7795), .ZN(n7797) );
  NAND2_X1 U9516 ( .A1(n9809), .A2(n7822), .ZN(n7796) );
  OAI211_X1 U9517 ( .C1(n7814), .C2(n9804), .A(n7797), .B(n7796), .ZN(n7798)
         );
  AOI21_X1 U9518 ( .B1(n10132), .B2(n9792), .A(n7798), .ZN(n7799) );
  OAI21_X1 U9519 ( .B1(n7800), .B2(n9795), .A(n7799), .ZN(P1_U3222) );
  INV_X1 U9520 ( .A(n7801), .ZN(n8903) );
  OAI222_X1 U9521 ( .A1(P1_U3084), .A2(n7803), .B1(n8243), .B2(n8903), .C1(
        n7802), .C2(n8885), .ZN(P1_U3331) );
  AND2_X1 U9522 ( .A1(n8901), .A2(n7804), .ZN(n7806) );
  NAND2_X1 U9523 ( .A1(n8901), .A2(n7805), .ZN(n7936) );
  OAI211_X1 U9524 ( .C1(n7807), .C2(n7806), .A(n7936), .B(n9212), .ZN(n7811)
         );
  OAI22_X1 U9525 ( .A1(n7808), .A2(n9390), .B1(n7992), .B2(n9204), .ZN(n8029)
         );
  AND2_X1 U9526 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n8111) );
  NOR2_X1 U9527 ( .A1(n9230), .A2(n8032), .ZN(n7809) );
  AOI211_X1 U9528 ( .C1(n9182), .C2(n8029), .A(n8111), .B(n7809), .ZN(n7810)
         );
  OAI211_X1 U9529 ( .C1(n10512), .C2(n9252), .A(n7811), .B(n7810), .ZN(
        P2_U3219) );
  NAND2_X1 U9530 ( .A1(n10246), .A2(n7812), .ZN(n7813) );
  XNOR2_X1 U9531 ( .A(n7813), .B(n7815), .ZN(n7819) );
  OAI22_X1 U9532 ( .A1(n7814), .A2(n10340), .B1(n7928), .B2(n10338), .ZN(n7818) );
  XNOR2_X1 U9533 ( .A(n7816), .B(n7815), .ZN(n10137) );
  NOR2_X1 U9534 ( .A1(n10137), .A2(n7093), .ZN(n7817) );
  AOI211_X1 U9535 ( .C1(n10343), .C2(n7819), .A(n7818), .B(n7817), .ZN(n10136)
         );
  INV_X1 U9536 ( .A(n7820), .ZN(n7821) );
  AOI21_X1 U9537 ( .B1(n10132), .B2(n10240), .A(n7821), .ZN(n10134) );
  AOI22_X1 U9538 ( .A1(n10048), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7822), .B2(
        n10345), .ZN(n7823) );
  OAI21_X1 U9539 ( .B1(n4909), .B2(n10256), .A(n7823), .ZN(n7825) );
  NOR2_X1 U9540 ( .A1(n10137), .A2(n8161), .ZN(n7824) );
  AOI211_X1 U9541 ( .C1(n10134), .C2(n10331), .A(n7825), .B(n7824), .ZN(n7826)
         );
  OAI21_X1 U9542 ( .B1(n10136), .B2(n10048), .A(n7826), .ZN(P1_U3279) );
  INV_X1 U9543 ( .A(n7844), .ZN(n7829) );
  INV_X1 U9544 ( .A(n8885), .ZN(n10155) );
  AOI21_X1 U9545 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n10155), .A(n7827), .ZN(
        n7828) );
  OAI21_X1 U9546 ( .B1(n7829), .B2(n10157), .A(n7828), .ZN(P1_U3330) );
  AOI22_X1 U9547 ( .A1(n8079), .A2(n5467), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n8086), .ZN(n7832) );
  AOI21_X1 U9548 ( .B1(n7833), .B2(n7832), .A(n8085), .ZN(n7842) );
  AOI22_X1 U9549 ( .A1(n8079), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8171), .B2(
        n8086), .ZN(n7837) );
  OAI21_X1 U9550 ( .B1(n7837), .B2(n7836), .A(n8078), .ZN(n7840) );
  NAND2_X1 U9551 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8913) );
  NAND2_X1 U9552 ( .A1(n10441), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n7838) );
  OAI211_X1 U9553 ( .C1(n10443), .C2(n8086), .A(n8913), .B(n7838), .ZN(n7839)
         );
  AOI21_X1 U9554 ( .B1(n7840), .B2(n10440), .A(n7839), .ZN(n7841) );
  OAI21_X1 U9555 ( .B1(n7842), .B2(n10444), .A(n7841), .ZN(P2_U3259) );
  NAND2_X1 U9556 ( .A1(n7844), .A2(n7843), .ZN(n7845) );
  OAI211_X1 U9557 ( .C1(n8698), .C2(n8906), .A(n7845), .B(n9134), .ZN(P2_U3335) );
  XOR2_X1 U9558 ( .A(n7848), .B(n7847), .Z(n7849) );
  XNOR2_X1 U9559 ( .A(n7846), .B(n7849), .ZN(n7856) );
  AOI21_X1 U9560 ( .B1(n9768), .B2(n9819), .A(n7850), .ZN(n7853) );
  NAND2_X1 U9561 ( .A1(n9809), .A2(n7851), .ZN(n7852) );
  OAI211_X1 U9562 ( .C1(n10248), .C2(n9804), .A(n7853), .B(n7852), .ZN(n7854)
         );
  AOI21_X1 U9563 ( .B1(n10270), .B2(n9792), .A(n7854), .ZN(n7855) );
  OAI21_X1 U9564 ( .B1(n7856), .B2(n9795), .A(n7855), .ZN(P1_U3232) );
  NAND2_X1 U9565 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n8893) );
  INV_X1 U9566 ( .A(n8893), .ZN(n7863) );
  AND3_X1 U9567 ( .A1(n7859), .A2(n7858), .A3(n7857), .ZN(n7860) );
  NOR3_X1 U9568 ( .A1(n7861), .A2(n7860), .A3(n10444), .ZN(n7862) );
  AOI211_X1 U9569 ( .C1(P2_ADDR_REG_9__SCAN_IN), .C2(n10441), .A(n7863), .B(
        n7862), .ZN(n7868) );
  OAI211_X1 U9570 ( .C1(n7866), .C2(n7865), .A(n10440), .B(n7864), .ZN(n7867)
         );
  OAI211_X1 U9571 ( .C1(n10443), .C2(n7869), .A(n7868), .B(n7867), .ZN(
        P2_U3254) );
  NOR2_X1 U9572 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8815), .ZN(n7874) );
  AOI211_X1 U9573 ( .C1(n7872), .C2(n7871), .A(n7870), .B(n10444), .ZN(n7873)
         );
  AOI211_X1 U9574 ( .C1(P2_ADDR_REG_8__SCAN_IN), .C2(n10441), .A(n7874), .B(
        n7873), .ZN(n7879) );
  OAI211_X1 U9575 ( .C1(n7877), .C2(n7876), .A(n10440), .B(n7875), .ZN(n7878)
         );
  OAI211_X1 U9576 ( .C1(n10443), .C2(n7880), .A(n7879), .B(n7878), .ZN(
        P2_U3253) );
  AOI211_X1 U9577 ( .C1(n7883), .C2(n7882), .A(n7881), .B(n10444), .ZN(n7884)
         );
  AOI211_X1 U9578 ( .C1(P2_ADDR_REG_6__SCAN_IN), .C2(n10441), .A(n7885), .B(
        n7884), .ZN(n7892) );
  INV_X1 U9579 ( .A(n7886), .ZN(n7890) );
  INV_X1 U9580 ( .A(n7887), .ZN(n7889) );
  OAI211_X1 U9581 ( .C1(n7890), .C2(n7889), .A(n10440), .B(n7888), .ZN(n7891)
         );
  OAI211_X1 U9582 ( .C1(n10443), .C2(n7893), .A(n7892), .B(n7891), .ZN(
        P2_U3251) );
  NAND2_X1 U9583 ( .A1(n7895), .A2(n7894), .ZN(n7963) );
  INV_X1 U9584 ( .A(n8023), .ZN(n7896) );
  AOI21_X1 U9585 ( .B1(n8951), .B2(n7963), .A(n7896), .ZN(n8058) );
  XNOR2_X1 U9586 ( .A(n7897), .B(n8951), .ZN(n7899) );
  OAI22_X1 U9587 ( .A1(n9023), .A2(n9390), .B1(n8895), .B2(n9204), .ZN(n7898)
         );
  AOI21_X1 U9588 ( .B1(n7899), .B2(n9532), .A(n7898), .ZN(n7900) );
  OAI21_X1 U9589 ( .B1(n8058), .B2(n8260), .A(n7900), .ZN(n8059) );
  NAND2_X1 U9590 ( .A1(n8059), .A2(n9540), .ZN(n7905) );
  AOI211_X1 U9591 ( .C1(n8898), .C2(n4514), .A(n10520), .B(n8034), .ZN(n8060)
         );
  INV_X1 U9592 ( .A(n8898), .ZN(n8065) );
  NOR2_X1 U9593 ( .A1(n9552), .A2(n8065), .ZN(n7903) );
  OAI22_X1 U9594 ( .A1(n9540), .A2(n7901), .B1(n8892), .B2(n9537), .ZN(n7902)
         );
  AOI211_X1 U9595 ( .C1(n8060), .C2(n9504), .A(n7903), .B(n7902), .ZN(n7904)
         );
  OAI211_X1 U9596 ( .C1(n8058), .C2(n8043), .A(n7905), .B(n7904), .ZN(P2_U3287) );
  OR2_X1 U9597 ( .A1(n7963), .A2(n7906), .ZN(n7908) );
  AND2_X1 U9598 ( .A1(n7908), .A2(n7907), .ZN(n7909) );
  XNOR2_X1 U9599 ( .A(n7909), .B(n8953), .ZN(n7958) );
  XOR2_X1 U9600 ( .A(n7910), .B(n8953), .Z(n7913) );
  OR2_X1 U9601 ( .A1(n8051), .A2(n9204), .ZN(n7912) );
  OR2_X1 U9602 ( .A1(n8895), .A2(n9390), .ZN(n7911) );
  NAND2_X1 U9603 ( .A1(n7912), .A2(n7911), .ZN(n7940) );
  AOI21_X1 U9604 ( .B1(n7913), .B2(n9532), .A(n7940), .ZN(n7961) );
  OAI211_X1 U9605 ( .C1(n8036), .C2(n7945), .A(n9541), .B(n7914), .ZN(n7954)
         );
  OAI211_X1 U9606 ( .C1(n7958), .C2(n10478), .A(n7961), .B(n7954), .ZN(n7947)
         );
  OAI22_X1 U9607 ( .A1(n9640), .A2(n7945), .B1(n10541), .B2(n7697), .ZN(n7915)
         );
  AOI21_X1 U9608 ( .B1(n7947), .B2(n10541), .A(n7915), .ZN(n7916) );
  INV_X1 U9609 ( .A(n7916), .ZN(P2_U3531) );
  NAND2_X1 U9610 ( .A1(n7918), .A2(n7917), .ZN(n7920) );
  NAND2_X1 U9611 ( .A1(n10270), .A2(n9820), .ZN(n7919) );
  XOR2_X1 U9612 ( .A(n8144), .B(n8149), .Z(n10131) );
  INV_X1 U9613 ( .A(n10129), .ZN(n7984) );
  OR2_X1 U9614 ( .A1(n7921), .A2(n7984), .ZN(n7922) );
  AND3_X1 U9615 ( .A1(n7922), .A2(n8156), .A3(n10265), .ZN(n10128) );
  INV_X1 U9616 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7923) );
  OAI22_X1 U9617 ( .A1(n7984), .A2(n10256), .B1(n7923), .B2(n10349), .ZN(n7931) );
  XNOR2_X1 U9618 ( .A(n8145), .B(n8144), .ZN(n7927) );
  OAI222_X1 U9619 ( .A1(n10338), .A2(n8226), .B1(n10340), .B2(n7928), .C1(
        n9988), .C2(n7927), .ZN(n10127) );
  AOI21_X1 U9620 ( .B1(n7987), .B2(n10345), .A(n10127), .ZN(n7929) );
  NOR2_X1 U9621 ( .A1(n7929), .A2(n10048), .ZN(n7930) );
  AOI211_X1 U9622 ( .C1(n10128), .C2(n10041), .A(n7931), .B(n7930), .ZN(n7932)
         );
  OAI21_X1 U9623 ( .B1(n10131), .B2(n10062), .A(n7932), .ZN(P1_U3277) );
  INV_X1 U9624 ( .A(n7937), .ZN(n7933) );
  AOI21_X1 U9625 ( .B1(n7936), .B2(n7933), .A(n9240), .ZN(n7939) );
  NOR3_X1 U9626 ( .A1(n9223), .A2(n7934), .A3(n8895), .ZN(n7938) );
  NAND2_X1 U9627 ( .A1(n7936), .A2(n7935), .ZN(n7995) );
  NAND2_X1 U9628 ( .A1(n7995), .A2(n7937), .ZN(n7991) );
  OAI21_X1 U9629 ( .B1(n7939), .B2(n7938), .A(n7991), .ZN(n7944) );
  AOI22_X1 U9630 ( .A1(n9182), .A2(n7940), .B1(P2_REG3_REG_11__SCAN_IN), .B2(
        P2_U3152), .ZN(n7941) );
  OAI21_X1 U9631 ( .B1(n9230), .B2(n7952), .A(n7941), .ZN(n7942) );
  INV_X1 U9632 ( .A(n7942), .ZN(n7943) );
  OAI211_X1 U9633 ( .C1(n7945), .C2(n9252), .A(n7944), .B(n7943), .ZN(P2_U3238) );
  OAI22_X1 U9634 ( .A1(n9692), .A2(n7945), .B1(n10528), .B2(n5410), .ZN(n7946)
         );
  AOI21_X1 U9635 ( .B1(n7947), .B2(n10528), .A(n7946), .ZN(n7948) );
  INV_X1 U9636 ( .A(n7948), .ZN(P2_U3484) );
  INV_X1 U9637 ( .A(n7949), .ZN(n7977) );
  OAI222_X1 U9638 ( .A1(n7951), .A2(P1_U3084), .B1(n8243), .B2(n7977), .C1(
        n7950), .C2(n8885), .ZN(P1_U3329) );
  INV_X1 U9639 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7953) );
  OAI22_X1 U9640 ( .A1(n9540), .A2(n7953), .B1(n7952), .B2(n9537), .ZN(n7956)
         );
  NOR2_X1 U9641 ( .A1(n7954), .A2(n10224), .ZN(n7955) );
  AOI211_X1 U9642 ( .C1(n10221), .C2(n7957), .A(n7956), .B(n7955), .ZN(n7960)
         );
  OR2_X1 U9643 ( .A1(n7958), .A2(n9536), .ZN(n7959) );
  OAI211_X1 U9644 ( .C1(n7961), .C2(n4499), .A(n7960), .B(n7959), .ZN(P2_U3285) );
  OR2_X1 U9645 ( .A1(n7963), .A2(n7962), .ZN(n7965) );
  AND2_X1 U9646 ( .A1(n7965), .A2(n7964), .ZN(n7966) );
  XNOR2_X1 U9647 ( .A(n7966), .B(n8956), .ZN(n10525) );
  INV_X1 U9648 ( .A(n10525), .ZN(n7976) );
  OAI211_X1 U9649 ( .C1(n4555), .C2(n8956), .A(n7967), .B(n9532), .ZN(n7969)
         );
  NAND2_X1 U9650 ( .A1(n9269), .A2(n9245), .ZN(n7968) );
  OAI211_X1 U9651 ( .C1(n9049), .C2(n9204), .A(n7969), .B(n7968), .ZN(n10522)
         );
  INV_X1 U9652 ( .A(n7914), .ZN(n7970) );
  INV_X1 U9653 ( .A(n6765), .ZN(n10519) );
  OAI21_X1 U9654 ( .B1(n7970), .B2(n10519), .A(n8268), .ZN(n10521) );
  OAI22_X1 U9655 ( .A1(n9540), .A2(n7971), .B1(n8003), .B2(n9537), .ZN(n7972)
         );
  AOI21_X1 U9656 ( .B1(n10221), .B2(n6765), .A(n7972), .ZN(n7973) );
  OAI21_X1 U9657 ( .B1(n10521), .B2(n8037), .A(n7973), .ZN(n7974) );
  AOI21_X1 U9658 ( .B1(n10522), .B2(n9540), .A(n7974), .ZN(n7975) );
  OAI21_X1 U9659 ( .B1(n7976), .B2(n9536), .A(n7975), .ZN(P2_U3284) );
  OAI222_X1 U9660 ( .A1(n7978), .A2(P2_U3152), .B1(n8906), .B2(n8553), .C1(
        n8904), .C2(n7977), .ZN(P2_U3334) );
  XOR2_X1 U9661 ( .A(n7980), .B(n7979), .Z(n7981) );
  XNOR2_X1 U9662 ( .A(n7982), .B(n7981), .ZN(n7989) );
  NAND2_X1 U9663 ( .A1(n9786), .A2(n9820), .ZN(n7983) );
  NAND2_X1 U9664 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3084), .ZN(n8013) );
  OAI211_X1 U9665 ( .C1(n8226), .C2(n9806), .A(n7983), .B(n8013), .ZN(n7986)
         );
  NOR2_X1 U9666 ( .A1(n7984), .A2(n9812), .ZN(n7985) );
  AOI211_X1 U9667 ( .C1(n9809), .C2(n7987), .A(n7986), .B(n7985), .ZN(n7988)
         );
  OAI21_X1 U9668 ( .B1(n7989), .B2(n9795), .A(n7988), .ZN(P1_U3213) );
  AOI21_X1 U9669 ( .B1(n7991), .B2(n7990), .A(n9240), .ZN(n7999) );
  NOR3_X1 U9670 ( .A1(n7993), .A2(n9223), .A3(n7992), .ZN(n7998) );
  NAND2_X1 U9671 ( .A1(n7995), .A2(n7994), .ZN(n7997) );
  AND2_X1 U9672 ( .A1(n7997), .A2(n7996), .ZN(n8046) );
  OAI21_X1 U9673 ( .B1(n7999), .B2(n7998), .A(n8046), .ZN(n8007) );
  NAND2_X1 U9674 ( .A1(n9224), .A2(n9269), .ZN(n8002) );
  NOR2_X1 U9675 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8000), .ZN(n8195) );
  INV_X1 U9676 ( .A(n8195), .ZN(n8001) );
  OAI211_X1 U9677 ( .C1(n9049), .C2(n9218), .A(n8002), .B(n8001), .ZN(n8005)
         );
  NOR2_X1 U9678 ( .A1(n9230), .A2(n8003), .ZN(n8004) );
  NOR2_X1 U9679 ( .A1(n8005), .A2(n8004), .ZN(n8006) );
  OAI211_X1 U9680 ( .C1(n10519), .C2(n9252), .A(n8007), .B(n8006), .ZN(
        P2_U3226) );
  AOI21_X1 U9681 ( .B1(n7599), .B2(n8009), .A(n8008), .ZN(n8012) );
  INV_X1 U9682 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n8285) );
  AOI22_X1 U9683 ( .A1(P1_REG1_REG_14__SCAN_IN), .A2(n8284), .B1(n8010), .B2(
        n8285), .ZN(n8011) );
  NOR2_X1 U9684 ( .A1(n8012), .A2(n8011), .ZN(n8283) );
  AOI21_X1 U9685 ( .B1(n8012), .B2(n8011), .A(n8283), .ZN(n8020) );
  OAI21_X1 U9686 ( .B1(n8284), .B2(n9899), .A(n8013), .ZN(n8018) );
  AOI211_X1 U9687 ( .C1(n8016), .C2(n7923), .A(n8279), .B(n10313), .ZN(n8017)
         );
  AOI211_X1 U9688 ( .C1(n10312), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n8018), .B(
        n8017), .ZN(n8019) );
  OAI21_X1 U9689 ( .B1(n8020), .B2(n9895), .A(n8019), .ZN(P1_U3255) );
  AND2_X1 U9690 ( .A1(n8023), .A2(n8021), .ZN(n8026) );
  NAND2_X1 U9691 ( .A1(n8023), .A2(n8022), .ZN(n8024) );
  OAI21_X1 U9692 ( .B1(n8026), .B2(n8025), .A(n8024), .ZN(n10511) );
  OAI21_X1 U9693 ( .B1(n8950), .B2(n8028), .A(n8027), .ZN(n8030) );
  AOI21_X1 U9694 ( .B1(n8030), .B2(n9532), .A(n8029), .ZN(n8031) );
  OAI21_X1 U9695 ( .B1(n10511), .B2(n8260), .A(n8031), .ZN(n10514) );
  NAND2_X1 U9696 ( .A1(n10514), .A2(n9540), .ZN(n8042) );
  INV_X1 U9697 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8033) );
  OAI22_X1 U9698 ( .A1(n9540), .A2(n8033), .B1(n8032), .B2(n9537), .ZN(n8039)
         );
  NOR2_X1 U9699 ( .A1(n8034), .A2(n10512), .ZN(n8035) );
  OR2_X1 U9700 ( .A1(n8036), .A2(n8035), .ZN(n10513) );
  NOR2_X1 U9701 ( .A1(n10513), .A2(n8037), .ZN(n8038) );
  AOI211_X1 U9702 ( .C1(n10221), .C2(n8040), .A(n8039), .B(n8038), .ZN(n8041)
         );
  OAI211_X1 U9703 ( .C1(n10511), .C2(n8043), .A(n8042), .B(n8041), .ZN(
        P2_U3286) );
  INV_X1 U9704 ( .A(n8044), .ZN(n8045) );
  AOI21_X1 U9705 ( .B1(n8046), .B2(n8045), .A(n9240), .ZN(n8050) );
  NOR3_X1 U9706 ( .A1(n8047), .A2(n8051), .A3(n9223), .ZN(n8049) );
  OAI21_X1 U9707 ( .B1(n8050), .B2(n8049), .A(n8048), .ZN(n8057) );
  OR2_X1 U9708 ( .A1(n8249), .A2(n9204), .ZN(n8053) );
  OR2_X1 U9709 ( .A1(n8051), .A2(n9390), .ZN(n8052) );
  NAND2_X1 U9710 ( .A1(n8053), .A2(n8052), .ZN(n8264) );
  NOR2_X1 U9711 ( .A1(n9230), .A2(n10217), .ZN(n8054) );
  AOI211_X1 U9712 ( .C1(n9182), .C2(n8264), .A(n8055), .B(n8054), .ZN(n8056)
         );
  OAI211_X1 U9713 ( .C1(n4780), .C2(n9252), .A(n8057), .B(n8056), .ZN(P2_U3236) );
  INV_X1 U9714 ( .A(n8272), .ZN(n10517) );
  INV_X1 U9715 ( .A(n8058), .ZN(n8061) );
  AOI211_X1 U9716 ( .C1(n10517), .C2(n8061), .A(n8060), .B(n8059), .ZN(n8068)
         );
  OAI22_X1 U9717 ( .A1(n9640), .A2(n8065), .B1(n10541), .B2(n8062), .ZN(n8063)
         );
  INV_X1 U9718 ( .A(n8063), .ZN(n8064) );
  OAI21_X1 U9719 ( .B1(n8068), .B2(n10539), .A(n8064), .ZN(P2_U3529) );
  OAI22_X1 U9720 ( .A1(n9692), .A2(n8065), .B1(n10528), .B2(n5338), .ZN(n8066)
         );
  INV_X1 U9721 ( .A(n8066), .ZN(n8067) );
  OAI21_X1 U9722 ( .B1(n8068), .B2(n10526), .A(n8067), .ZN(P2_U3478) );
  XNOR2_X1 U9723 ( .A(n8070), .B(n8069), .ZN(n8071) );
  XNOR2_X1 U9724 ( .A(n8072), .B(n8071), .ZN(n8077) );
  INV_X1 U9725 ( .A(n8316), .ZN(n9817) );
  INV_X1 U9726 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n8693) );
  NOR2_X1 U9727 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8693), .ZN(n8287) );
  AOI21_X1 U9728 ( .B1(n9768), .B2(n9817), .A(n8287), .ZN(n8074) );
  NAND2_X1 U9729 ( .A1(n9809), .A2(n8158), .ZN(n8073) );
  OAI211_X1 U9730 ( .C1(n8146), .C2(n9804), .A(n8074), .B(n8073), .ZN(n8075)
         );
  AOI21_X1 U9731 ( .B1(n10122), .B2(n9792), .A(n8075), .ZN(n8076) );
  OAI21_X1 U9732 ( .B1(n8077), .B2(n9795), .A(n8076), .ZN(P1_U3239) );
  OAI21_X1 U9733 ( .B1(n8079), .B2(P2_REG2_REG_14__SCAN_IN), .A(n8078), .ZN(
        n8390) );
  XNOR2_X1 U9734 ( .A(n8390), .B(n8380), .ZN(n8080) );
  NAND2_X1 U9735 ( .A1(n8080), .A2(n5508), .ZN(n8392) );
  OAI21_X1 U9736 ( .B1(n8080), .B2(n5508), .A(n8392), .ZN(n8084) );
  AND2_X1 U9737 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8081) );
  AOI21_X1 U9738 ( .B1(n10441), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n8081), .ZN(
        n8082) );
  OAI21_X1 U9739 ( .B1(n10443), .B2(n8391), .A(n8082), .ZN(n8083) );
  AOI21_X1 U9740 ( .B1(n8084), .B2(n10440), .A(n8083), .ZN(n8089) );
  XNOR2_X1 U9741 ( .A(n8379), .B(n8391), .ZN(n8087) );
  INV_X1 U9742 ( .A(n10444), .ZN(n10439) );
  NAND2_X1 U9743 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n8087), .ZN(n8381) );
  OAI211_X1 U9744 ( .C1(n8087), .C2(P2_REG1_REG_15__SCAN_IN), .A(n10439), .B(
        n8381), .ZN(n8088) );
  NAND2_X1 U9745 ( .A1(n8089), .A2(n8088), .ZN(P2_U3260) );
  INV_X1 U9746 ( .A(n8090), .ZN(n8242) );
  OAI222_X1 U9747 ( .A1(P2_U3152), .A2(n8092), .B1(n8904), .B2(n8242), .C1(
        n8091), .C2(n8906), .ZN(P2_U3333) );
  AOI211_X1 U9748 ( .C1(n8095), .C2(n8094), .A(n8093), .B(n10442), .ZN(n8104)
         );
  NOR2_X1 U9749 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8522), .ZN(n8096) );
  AOI21_X1 U9750 ( .B1(n10441), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n8096), .ZN(
        n8101) );
  OAI211_X1 U9751 ( .C1(n8099), .C2(n8098), .A(n10439), .B(n8097), .ZN(n8100)
         );
  OAI211_X1 U9752 ( .C1(n10443), .C2(n8102), .A(n8101), .B(n8100), .ZN(n8103)
         );
  OR2_X1 U9753 ( .A1(n8104), .A2(n8103), .ZN(P2_U3248) );
  AOI211_X1 U9754 ( .C1(n8107), .C2(n8106), .A(n8105), .B(n10442), .ZN(n8116)
         );
  OAI211_X1 U9755 ( .C1(n8110), .C2(n8109), .A(n8108), .B(n10439), .ZN(n8113)
         );
  AOI21_X1 U9756 ( .B1(n10441), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n8111), .ZN(
        n8112) );
  OAI211_X1 U9757 ( .C1(n10443), .C2(n8114), .A(n8113), .B(n8112), .ZN(n8115)
         );
  OR2_X1 U9758 ( .A1(n8116), .A2(n8115), .ZN(P2_U3255) );
  AOI211_X1 U9759 ( .C1(n8119), .C2(n8118), .A(n8117), .B(n10442), .ZN(n8128)
         );
  AND2_X1 U9760 ( .A1(P2_U3152), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8120) );
  AOI21_X1 U9761 ( .B1(n10441), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n8120), .ZN(
        n8125) );
  OAI211_X1 U9762 ( .C1(n8123), .C2(n8122), .A(n10439), .B(n8121), .ZN(n8124)
         );
  OAI211_X1 U9763 ( .C1(n10443), .C2(n8126), .A(n8125), .B(n8124), .ZN(n8127)
         );
  OR2_X1 U9764 ( .A1(n8128), .A2(n8127), .ZN(P2_U3252) );
  AOI211_X1 U9765 ( .C1(n8131), .C2(n8130), .A(n8129), .B(n10442), .ZN(n8142)
         );
  INV_X1 U9766 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n8133) );
  OAI22_X1 U9767 ( .A1(n9339), .A2(n8133), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8132), .ZN(n8134) );
  INV_X1 U9768 ( .A(n8134), .ZN(n8139) );
  OAI211_X1 U9769 ( .C1(n8137), .C2(n8136), .A(n10439), .B(n8135), .ZN(n8138)
         );
  OAI211_X1 U9770 ( .C1(n10443), .C2(n8140), .A(n8139), .B(n8138), .ZN(n8141)
         );
  OR2_X1 U9771 ( .A1(n8142), .A2(n8141), .ZN(P2_U3246) );
  XNOR2_X1 U9772 ( .A(n8222), .B(n8150), .ZN(n8155) );
  OAI22_X1 U9773 ( .A1(n8146), .A2(n10340), .B1(n8316), .B2(n10338), .ZN(n8154) );
  AND2_X1 U9774 ( .A1(n10129), .A2(n9819), .ZN(n8148) );
  OR2_X1 U9775 ( .A1(n10129), .A2(n9819), .ZN(n8147) );
  AND2_X1 U9776 ( .A1(n8151), .A2(n8150), .ZN(n8152) );
  OR2_X1 U9777 ( .A1(n8228), .A2(n8152), .ZN(n10126) );
  NOR2_X1 U9778 ( .A1(n10126), .A2(n7093), .ZN(n8153) );
  AOI211_X1 U9779 ( .C1(n10343), .C2(n8155), .A(n8154), .B(n8153), .ZN(n10125)
         );
  NAND2_X1 U9780 ( .A1(n8156), .A2(n10122), .ZN(n8157) );
  AND2_X1 U9781 ( .A1(n8233), .A2(n8157), .ZN(n10123) );
  INV_X1 U9782 ( .A(n10122), .ZN(n8160) );
  AOI22_X1 U9783 ( .A1(n10048), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n8158), .B2(
        n10345), .ZN(n8159) );
  OAI21_X1 U9784 ( .B1(n8160), .B2(n10256), .A(n8159), .ZN(n8163) );
  NOR2_X1 U9785 ( .A1(n10126), .A2(n8161), .ZN(n8162) );
  AOI211_X1 U9786 ( .C1(n10123), .C2(n10331), .A(n8163), .B(n8162), .ZN(n8164)
         );
  OAI21_X1 U9787 ( .B1(n10125), .B2(n10048), .A(n8164), .ZN(P1_U3276) );
  OAI211_X1 U9788 ( .C1(n8166), .C2(n9054), .A(n8165), .B(n9532), .ZN(n8169)
         );
  OR2_X1 U9789 ( .A1(n8303), .A2(n9204), .ZN(n8168) );
  OR2_X1 U9790 ( .A1(n9049), .A2(n9390), .ZN(n8167) );
  AND2_X1 U9791 ( .A1(n8168), .A2(n8167), .ZN(n8914) );
  NAND2_X1 U9792 ( .A1(n8169), .A2(n8914), .ZN(n8368) );
  INV_X1 U9793 ( .A(n8368), .ZN(n8176) );
  XNOR2_X1 U9794 ( .A(n8170), .B(n9054), .ZN(n8370) );
  NAND2_X1 U9795 ( .A1(n8370), .A2(n9465), .ZN(n8175) );
  AOI211_X1 U9796 ( .C1(n8917), .C2(n4782), .A(n10520), .B(n8357), .ZN(n8369)
         );
  NOR2_X1 U9797 ( .A1(n8375), .A2(n9552), .ZN(n8173) );
  OAI22_X1 U9798 ( .A1(n9540), .A2(n8171), .B1(n8912), .B2(n9537), .ZN(n8172)
         );
  AOI211_X1 U9799 ( .C1(n8369), .C2(n9504), .A(n8173), .B(n8172), .ZN(n8174)
         );
  OAI211_X1 U9800 ( .C1(n4499), .C2(n8176), .A(n8175), .B(n8174), .ZN(P2_U3282) );
  INV_X1 U9801 ( .A(n8177), .ZN(n8218) );
  OAI222_X1 U9802 ( .A1(n8179), .A2(P1_U3084), .B1(n10157), .B2(n8218), .C1(
        n8178), .C2(n8885), .ZN(P1_U3327) );
  AOI211_X1 U9803 ( .C1(n8182), .C2(n8181), .A(n8180), .B(n10442), .ZN(n8183)
         );
  INV_X1 U9804 ( .A(n8183), .ZN(n8190) );
  NAND2_X1 U9805 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n9216) );
  INV_X1 U9806 ( .A(n9216), .ZN(n8188) );
  AOI211_X1 U9807 ( .C1(n8186), .C2(n8185), .A(n8184), .B(n10444), .ZN(n8187)
         );
  AOI211_X1 U9808 ( .C1(P2_ADDR_REG_4__SCAN_IN), .C2(n10441), .A(n8188), .B(
        n8187), .ZN(n8189) );
  OAI211_X1 U9809 ( .C1(n10443), .C2(n8191), .A(n8190), .B(n8189), .ZN(
        P2_U3249) );
  AOI21_X1 U9810 ( .B1(n8194), .B2(n8193), .A(n8192), .ZN(n8197) );
  AOI21_X1 U9811 ( .B1(n10441), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n8195), .ZN(
        n8196) );
  OAI21_X1 U9812 ( .B1(n8197), .B2(n10444), .A(n8196), .ZN(n8202) );
  AOI211_X1 U9813 ( .C1(n8200), .C2(n8199), .A(n8198), .B(n10442), .ZN(n8201)
         );
  AOI211_X1 U9814 ( .C1(n10165), .C2(n8203), .A(n8202), .B(n8201), .ZN(n8204)
         );
  INV_X1 U9815 ( .A(n8204), .ZN(P2_U3257) );
  XNOR2_X1 U9816 ( .A(n8206), .B(n8205), .ZN(n8210) );
  NOR2_X1 U9817 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8207), .ZN(n8208) );
  AOI21_X1 U9818 ( .B1(n10441), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n8208), .ZN(
        n8209) );
  OAI21_X1 U9819 ( .B1(n10444), .B2(n8210), .A(n8209), .ZN(n8215) );
  AOI211_X1 U9820 ( .C1(n8213), .C2(n8212), .A(n8211), .B(n10442), .ZN(n8214)
         );
  AOI211_X1 U9821 ( .C1(n10165), .C2(n8216), .A(n8215), .B(n8214), .ZN(n8217)
         );
  INV_X1 U9822 ( .A(n8217), .ZN(P2_U3250) );
  OAI222_X1 U9823 ( .A1(n8220), .A2(P2_U3152), .B1(n8906), .B2(n8219), .C1(
        n8904), .C2(n8218), .ZN(P2_U3332) );
  INV_X1 U9824 ( .A(n8223), .ZN(n8224) );
  NOR2_X1 U9825 ( .A1(n8313), .A2(n8224), .ZN(n8225) );
  XNOR2_X1 U9826 ( .A(n8225), .B(n8229), .ZN(n8227) );
  INV_X1 U9827 ( .A(n8226), .ZN(n9818) );
  AOI222_X1 U9828 ( .A1(n10343), .A2(n8227), .B1(n9816), .B2(n10056), .C1(
        n9818), .C2(n10054), .ZN(n10267) );
  AOI21_X1 U9829 ( .B1(n4559), .B2(n8229), .A(n8310), .ZN(n10269) );
  NAND2_X1 U9830 ( .A1(n10269), .A2(n8864), .ZN(n8240) );
  INV_X1 U9831 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n8232) );
  OAI22_X1 U9832 ( .A1(n10349), .A2(n8232), .B1(n8231), .B2(n8230), .ZN(n8237)
         );
  INV_X1 U9833 ( .A(n8233), .ZN(n8234) );
  INV_X1 U9834 ( .A(n8317), .ZN(n8319) );
  OAI211_X1 U9835 ( .C1(n4672), .C2(n8234), .A(n8319), .B(n10265), .ZN(n10266)
         );
  NOR2_X1 U9836 ( .A1(n10266), .A2(n8235), .ZN(n8236) );
  AOI211_X1 U9837 ( .C1(n8238), .C2(n8332), .A(n8237), .B(n8236), .ZN(n8239)
         );
  OAI211_X1 U9838 ( .C1(n10048), .C2(n10267), .A(n8240), .B(n8239), .ZN(
        P1_U3275) );
  OAI222_X1 U9839 ( .A1(P1_U3084), .A2(n8244), .B1(n8243), .B2(n8242), .C1(
        n8241), .C2(n8885), .ZN(P1_U3328) );
  NAND2_X1 U9840 ( .A1(n9235), .A2(n9266), .ZN(n8247) );
  NAND2_X1 U9841 ( .A1(n9212), .A2(n8297), .ZN(n8246) );
  XNOR2_X1 U9842 ( .A(n8295), .B(n8245), .ZN(n8298) );
  MUX2_X1 U9843 ( .A(n8247), .B(n8246), .S(n8298), .Z(n8255) );
  INV_X1 U9844 ( .A(n8248), .ZN(n8362) );
  OR2_X1 U9845 ( .A1(n8249), .A2(n9390), .ZN(n8251) );
  NAND2_X1 U9846 ( .A1(n9265), .A2(n9386), .ZN(n8250) );
  AND2_X1 U9847 ( .A1(n8251), .A2(n8250), .ZN(n8355) );
  OAI22_X1 U9848 ( .A1(n9247), .A2(n8355), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8252), .ZN(n8253) );
  AOI21_X1 U9849 ( .B1(n8362), .B2(n9249), .A(n8253), .ZN(n8254) );
  OAI211_X1 U9850 ( .C1(n8449), .C2(n9252), .A(n8255), .B(n8254), .ZN(P2_U3243) );
  INV_X1 U9851 ( .A(n8256), .ZN(n8294) );
  AOI21_X1 U9852 ( .B1(P2_DATAO_REG_27__SCAN_IN), .B2(n10155), .A(n9896), .ZN(
        n8257) );
  OAI21_X1 U9853 ( .B1(n8294), .B2(n10157), .A(n8257), .ZN(P1_U3326) );
  OAI21_X1 U9854 ( .B1(n8259), .B2(n9055), .A(n8258), .ZN(n10216) );
  OR2_X1 U9855 ( .A1(n10216), .A2(n8260), .ZN(n8267) );
  NAND2_X1 U9856 ( .A1(n8261), .A2(n9055), .ZN(n8262) );
  NAND2_X1 U9857 ( .A1(n8263), .A2(n8262), .ZN(n8265) );
  AOI21_X1 U9858 ( .B1(n8265), .B2(n9532), .A(n8264), .ZN(n8266) );
  NAND2_X1 U9859 ( .A1(n8268), .A2(n10220), .ZN(n8269) );
  NAND2_X1 U9860 ( .A1(n8269), .A2(n9541), .ZN(n8270) );
  OR2_X1 U9861 ( .A1(n8271), .A2(n8270), .ZN(n10225) );
  OAI21_X1 U9862 ( .B1(n10216), .B2(n8272), .A(n10225), .ZN(n8273) );
  INV_X1 U9863 ( .A(n8273), .ZN(n8274) );
  AND2_X1 U9864 ( .A1(n10230), .A2(n8274), .ZN(n8276) );
  MUX2_X1 U9865 ( .A(n8276), .B(n5447), .S(n10526), .Z(n8275) );
  OAI21_X1 U9866 ( .B1(n4780), .B2(n9692), .A(n8275), .ZN(P2_U3490) );
  MUX2_X1 U9867 ( .A(n5443), .B(n8276), .S(n10541), .Z(n8277) );
  OAI21_X1 U9868 ( .B1(n4780), .B2(n9640), .A(n8277), .ZN(P2_U3533) );
  NOR2_X1 U9869 ( .A1(n8278), .A2(n8284), .ZN(n8280) );
  INV_X1 U9870 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n8281) );
  NOR2_X1 U9871 ( .A1(n8281), .A2(n8282), .ZN(n9834) );
  AOI211_X1 U9872 ( .C1(n8282), .C2(n8281), .A(n9834), .B(n10313), .ZN(n8292)
         );
  INV_X1 U9873 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n8290) );
  AOI21_X1 U9874 ( .B1(n8285), .B2(n8284), .A(n8283), .ZN(n9838) );
  XNOR2_X1 U9875 ( .A(n9832), .B(n9838), .ZN(n8286) );
  NAND2_X1 U9876 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n8286), .ZN(n9840) );
  OAI211_X1 U9877 ( .C1(n8286), .C2(P1_REG1_REG_15__SCAN_IN), .A(n10319), .B(
        n9840), .ZN(n8289) );
  AOI21_X1 U9878 ( .B1(n9839), .B2(n10310), .A(n8287), .ZN(n8288) );
  OAI211_X1 U9879 ( .C1(n8290), .C2(n10305), .A(n8289), .B(n8288), .ZN(n8291)
         );
  OR2_X1 U9880 ( .A1(n8292), .A2(n8291), .ZN(P1_U3256) );
  OAI222_X1 U9881 ( .A1(n8904), .A2(n8294), .B1(P2_U3152), .B2(n9129), .C1(
        n8293), .C2(n8906), .ZN(P2_U3331) );
  AOI22_X1 U9882 ( .A1(n8298), .A2(n8297), .B1(n8296), .B2(n8295), .ZN(n8302)
         );
  XNOR2_X1 U9883 ( .A(n8300), .B(n8299), .ZN(n8301) );
  XNOR2_X1 U9884 ( .A(n8302), .B(n8301), .ZN(n8309) );
  NOR2_X1 U9885 ( .A1(n9230), .A2(n8425), .ZN(n8307) );
  OR2_X1 U9886 ( .A1(n8303), .A2(n9390), .ZN(n8305) );
  OR2_X1 U9887 ( .A1(n8341), .A2(n9204), .ZN(n8304) );
  AND2_X1 U9888 ( .A1(n8305), .A2(n8304), .ZN(n8420) );
  OAI22_X1 U9889 ( .A1(n9247), .A2(n8420), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8387), .ZN(n8306) );
  AOI211_X1 U9890 ( .C1(n9066), .C2(n10593), .A(n8307), .B(n8306), .ZN(n8308)
         );
  OAI21_X1 U9891 ( .B1(n8309), .B2(n9240), .A(n8308), .ZN(P2_U3228) );
  XOR2_X1 U9892 ( .A(n8314), .B(n8402), .Z(n10121) );
  XNOR2_X1 U9893 ( .A(n8408), .B(n8314), .ZN(n8315) );
  OAI222_X1 U9894 ( .A1(n10338), .A2(n9745), .B1(n10340), .B2(n8316), .C1(
        n8315), .C2(n9988), .ZN(n10117) );
  INV_X1 U9895 ( .A(n8404), .ZN(n8318) );
  AOI211_X1 U9896 ( .C1(n10119), .C2(n8319), .A(n10416), .B(n8318), .ZN(n10118) );
  NAND2_X1 U9897 ( .A1(n10118), .A2(n10041), .ZN(n8321) );
  AOI22_X1 U9898 ( .A1(n10048), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9747), .B2(
        n10345), .ZN(n8320) );
  OAI211_X1 U9899 ( .C1(n9750), .C2(n10256), .A(n8321), .B(n8320), .ZN(n8322)
         );
  AOI21_X1 U9900 ( .B1(n10117), .B2(n10349), .A(n8322), .ZN(n8323) );
  OAI21_X1 U9901 ( .B1(n10121), .B2(n10062), .A(n8323), .ZN(P1_U3274) );
  INV_X1 U9902 ( .A(n8324), .ZN(n8325) );
  AOI21_X1 U9903 ( .B1(n8327), .B2(n8326), .A(n8325), .ZN(n8335) );
  NAND2_X1 U9904 ( .A1(n9786), .A2(n9818), .ZN(n8328) );
  NAND2_X1 U9905 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9845) );
  OAI211_X1 U9906 ( .C1(n8329), .C2(n9806), .A(n8328), .B(n9845), .ZN(n8330)
         );
  AOI21_X1 U9907 ( .B1(n8331), .B2(n9809), .A(n8330), .ZN(n8334) );
  NAND2_X1 U9908 ( .A1(n8332), .A2(n9792), .ZN(n8333) );
  OAI211_X1 U9909 ( .C1(n8335), .C2(n9795), .A(n8334), .B(n8333), .ZN(P1_U3224) );
  AOI21_X1 U9910 ( .B1(n8435), .B2(n4845), .A(n9240), .ZN(n8340) );
  NOR3_X1 U9911 ( .A1(n8337), .A2(n8341), .A3(n9223), .ZN(n8339) );
  OAI21_X1 U9912 ( .B1(n8340), .B2(n8339), .A(n8338), .ZN(n8346) );
  OR2_X1 U9913 ( .A1(n8464), .A2(n9204), .ZN(n8343) );
  OR2_X1 U9914 ( .A1(n8341), .A2(n9390), .ZN(n8342) );
  NAND2_X1 U9915 ( .A1(n8343), .A2(n8342), .ZN(n9531) );
  AND2_X1 U9916 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n9321) );
  NOR2_X1 U9917 ( .A1(n9230), .A2(n9538), .ZN(n8344) );
  AOI211_X1 U9918 ( .C1(n9182), .C2(n9531), .A(n9321), .B(n8344), .ZN(n8345)
         );
  OAI211_X1 U9919 ( .C1(n9689), .C2(n9252), .A(n8346), .B(n8345), .ZN(P2_U3240) );
  INV_X1 U9920 ( .A(n8347), .ZN(n8378) );
  AOI21_X1 U9921 ( .B1(n10155), .B2(P2_DATAO_REG_28__SCAN_IN), .A(n8348), .ZN(
        n8349) );
  OAI21_X1 U9922 ( .B1(n8378), .B2(n10157), .A(n8349), .ZN(P1_U3325) );
  OAI21_X1 U9923 ( .B1(n8352), .B2(n8351), .A(n8350), .ZN(n8444) );
  INV_X1 U9924 ( .A(n8444), .ZN(n8367) );
  OAI211_X1 U9925 ( .C1(n8354), .C2(n9059), .A(n8353), .B(n9532), .ZN(n8356)
         );
  NAND2_X1 U9926 ( .A1(n8356), .A2(n8355), .ZN(n8442) );
  INV_X1 U9927 ( .A(n8357), .ZN(n8360) );
  INV_X1 U9928 ( .A(n8358), .ZN(n8359) );
  AOI211_X1 U9929 ( .C1(n8361), .C2(n8360), .A(n10520), .B(n8359), .ZN(n8443)
         );
  NAND2_X1 U9930 ( .A1(n8443), .A2(n9504), .ZN(n8364) );
  AOI22_X1 U9931 ( .A1(n4499), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8362), .B2(
        n10218), .ZN(n8363) );
  OAI211_X1 U9932 ( .C1(n8449), .C2(n9552), .A(n8364), .B(n8363), .ZN(n8365)
         );
  AOI21_X1 U9933 ( .B1(n8442), .B2(n9540), .A(n8365), .ZN(n8366) );
  OAI21_X1 U9934 ( .B1(n8367), .B2(n9536), .A(n8366), .ZN(P2_U3281) );
  AOI211_X1 U9935 ( .C1(n8370), .C2(n10524), .A(n8369), .B(n8368), .ZN(n8372)
         );
  MUX2_X1 U9936 ( .A(n5467), .B(n8372), .S(n10541), .Z(n8371) );
  OAI21_X1 U9937 ( .B1(n8375), .B2(n9640), .A(n8371), .ZN(P2_U3534) );
  INV_X1 U9938 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8373) );
  MUX2_X1 U9939 ( .A(n8373), .B(n8372), .S(n10528), .Z(n8374) );
  OAI21_X1 U9940 ( .B1(n8375), .B2(n9692), .A(n8374), .ZN(P2_U3493) );
  NAND2_X1 U9941 ( .A1(n9698), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8376) );
  OAI211_X1 U9942 ( .C1(n8378), .C2(n8904), .A(n8377), .B(n8376), .ZN(P2_U3330) );
  NAND2_X1 U9943 ( .A1(n8380), .A2(n8379), .ZN(n8382) );
  NAND2_X1 U9944 ( .A1(n8382), .A2(n8381), .ZN(n8386) );
  NOR2_X1 U9945 ( .A1(n9304), .A2(n8383), .ZN(n8384) );
  AOI21_X1 U9946 ( .B1(n8383), .B2(n9304), .A(n8384), .ZN(n8385) );
  AOI21_X1 U9947 ( .B1(n8386), .B2(n8385), .A(n9295), .ZN(n8400) );
  NOR2_X1 U9948 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8387), .ZN(n8388) );
  AOI21_X1 U9949 ( .B1(n10441), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8388), .ZN(
        n8389) );
  INV_X1 U9950 ( .A(n8389), .ZN(n8398) );
  NAND2_X1 U9951 ( .A1(n8391), .A2(n8390), .ZN(n8393) );
  NAND2_X1 U9952 ( .A1(n8393), .A2(n8392), .ZN(n8396) );
  NAND2_X1 U9953 ( .A1(n9304), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8394) );
  OAI21_X1 U9954 ( .B1(n9304), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8394), .ZN(
        n8395) );
  NOR2_X1 U9955 ( .A1(n8395), .A2(n8396), .ZN(n9303) );
  AOI211_X1 U9956 ( .C1(n8396), .C2(n8395), .A(n9303), .B(n10442), .ZN(n8397)
         );
  AOI211_X1 U9957 ( .C1(n10165), .C2(n9304), .A(n8398), .B(n8397), .ZN(n8399)
         );
  OAI21_X1 U9958 ( .B1(n8400), .B2(n10444), .A(n8399), .ZN(P2_U3261) );
  NOR2_X1 U9959 ( .A1(n10119), .A2(n9816), .ZN(n8401) );
  XNOR2_X1 U9960 ( .A(n8451), .B(n8450), .ZN(n10116) );
  INV_X1 U9961 ( .A(n8452), .ZN(n8403) );
  AOI21_X1 U9962 ( .B1(n10112), .B2(n8404), .A(n8403), .ZN(n10113) );
  INV_X1 U9963 ( .A(n10112), .ZN(n8406) );
  AOI22_X1 U9964 ( .A1(n10048), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9791), .B2(
        n10345), .ZN(n8405) );
  OAI21_X1 U9965 ( .B1(n8406), .B2(n10256), .A(n8405), .ZN(n8414) );
  NOR2_X1 U9966 ( .A1(n8456), .A2(n8409), .ZN(n8411) );
  XNOR2_X1 U9967 ( .A(n8411), .B(n8410), .ZN(n8412) );
  INV_X1 U9968 ( .A(n9789), .ZN(n10055) );
  AOI222_X1 U9969 ( .A1(n10343), .A2(n8412), .B1(n10055), .B2(n10056), .C1(
        n9816), .C2(n10054), .ZN(n10115) );
  NOR2_X1 U9970 ( .A1(n10115), .A2(n10048), .ZN(n8413) );
  AOI211_X1 U9971 ( .C1(n10113), .C2(n10331), .A(n8414), .B(n8413), .ZN(n8415)
         );
  OAI21_X1 U9972 ( .B1(n10116), .B2(n10062), .A(n8415), .ZN(P1_U3273) );
  NAND2_X1 U9973 ( .A1(n8416), .A2(n8958), .ZN(n8417) );
  NAND2_X1 U9974 ( .A1(n8418), .A2(n8417), .ZN(n8419) );
  NAND2_X1 U9975 ( .A1(n8419), .A2(n9532), .ZN(n8421) );
  NAND2_X1 U9976 ( .A1(n8421), .A2(n8420), .ZN(n9636) );
  INV_X1 U9977 ( .A(n9636), .ZN(n8431) );
  AOI21_X1 U9978 ( .B1(n9063), .B2(n8423), .A(n8422), .ZN(n9638) );
  NAND2_X1 U9979 ( .A1(n9638), .A2(n9465), .ZN(n8430) );
  INV_X1 U9980 ( .A(n9560), .ZN(n8424) );
  AOI211_X1 U9981 ( .C1(n9066), .C2(n8358), .A(n10520), .B(n8424), .ZN(n9637)
         );
  INV_X1 U9982 ( .A(n9066), .ZN(n9693) );
  NOR2_X1 U9983 ( .A1(n9693), .A2(n9552), .ZN(n8428) );
  INV_X1 U9984 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8426) );
  OAI22_X1 U9985 ( .A1(n9540), .A2(n8426), .B1(n8425), .B2(n9537), .ZN(n8427)
         );
  AOI211_X1 U9986 ( .C1(n9637), .C2(n9504), .A(n8428), .B(n8427), .ZN(n8429)
         );
  OAI211_X1 U9987 ( .C1(n4499), .C2(n8431), .A(n8430), .B(n8429), .ZN(P2_U3280) );
  OR2_X1 U9988 ( .A1(n9163), .A2(n9204), .ZN(n8433) );
  NAND2_X1 U9989 ( .A1(n9265), .A2(n9245), .ZN(n8432) );
  NAND2_X1 U9990 ( .A1(n8433), .A2(n8432), .ZN(n9556) );
  AOI22_X1 U9991 ( .A1(n9182), .A2(n9556), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3152), .ZN(n8434) );
  OAI21_X1 U9992 ( .B1(n9230), .B2(n9549), .A(n8434), .ZN(n8440) );
  INV_X1 U9993 ( .A(n8435), .ZN(n8436) );
  AOI211_X1 U9994 ( .C1(n8438), .C2(n8437), .A(n9240), .B(n8436), .ZN(n8439)
         );
  AOI211_X1 U9995 ( .C1(n9559), .C2(n10593), .A(n8440), .B(n8439), .ZN(n8441)
         );
  INV_X1 U9996 ( .A(n8441), .ZN(P2_U3230) );
  AOI211_X1 U9997 ( .C1(n8444), .C2(n10524), .A(n8443), .B(n8442), .ZN(n8446)
         );
  MUX2_X1 U9998 ( .A(n5507), .B(n8446), .S(n10541), .Z(n8445) );
  OAI21_X1 U9999 ( .B1(n8449), .B2(n9640), .A(n8445), .ZN(P2_U3535) );
  INV_X1 U10000 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8447) );
  MUX2_X1 U10001 ( .A(n8447), .B(n8446), .S(n10528), .Z(n8448) );
  OAI21_X1 U10002 ( .B1(n8449), .B2(n9692), .A(n8448), .ZN(P2_U3496) );
  INV_X1 U10003 ( .A(n9745), .ZN(n9815) );
  XNOR2_X1 U10004 ( .A(n8481), .B(n8480), .ZN(n10111) );
  AOI211_X1 U10005 ( .C1(n10108), .C2(n8452), .A(n10416), .B(n10045), .ZN(
        n10107) );
  INV_X1 U10006 ( .A(n10108), .ZN(n9722) );
  AOI22_X1 U10007 ( .A1(n10048), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9719), 
        .B2(n10345), .ZN(n8453) );
  OAI21_X1 U10008 ( .B1(n9722), .B2(n10256), .A(n8453), .ZN(n8460) );
  NAND2_X1 U10009 ( .A1(n8457), .A2(n8480), .ZN(n8495) );
  OAI21_X1 U10010 ( .B1(n8480), .B2(n8457), .A(n8495), .ZN(n8458) );
  INV_X1 U10011 ( .A(n9717), .ZN(n10036) );
  AOI222_X1 U10012 ( .A1(n10343), .A2(n8458), .B1(n10036), .B2(n10056), .C1(
        n9815), .C2(n10054), .ZN(n10110) );
  NOR2_X1 U10013 ( .A1(n10110), .A2(n10048), .ZN(n8459) );
  AOI211_X1 U10014 ( .C1(n10107), .C2(n10041), .A(n8460), .B(n8459), .ZN(n8461) );
  OAI21_X1 U10015 ( .B1(n10111), .B2(n10062), .A(n8461), .ZN(P1_U3272) );
  XNOR2_X1 U10016 ( .A(n8462), .B(n8463), .ZN(n8471) );
  NOR2_X1 U10017 ( .A1(n9230), .A2(n9505), .ZN(n8469) );
  OR2_X1 U10018 ( .A1(n8464), .A2(n9390), .ZN(n8466) );
  NAND2_X1 U10019 ( .A1(n9260), .A2(n9386), .ZN(n8465) );
  AND2_X1 U10020 ( .A1(n8466), .A2(n8465), .ZN(n9499) );
  OAI22_X1 U10021 ( .A1(n9247), .A2(n9499), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8467), .ZN(n8468) );
  AOI211_X1 U10022 ( .C1(n9503), .C2(n10593), .A(n8469), .B(n8468), .ZN(n8470)
         );
  OAI21_X1 U10023 ( .B1(n8471), .B2(n9240), .A(n8470), .ZN(P2_U3235) );
  INV_X1 U10024 ( .A(n8472), .ZN(n8475) );
  INV_X1 U10025 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8473) );
  OAI222_X1 U10026 ( .A1(P1_U3084), .A2(n8474), .B1(n10157), .B2(n8475), .C1(
        n8473), .C2(n8885), .ZN(P1_U3324) );
  INV_X1 U10027 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8477) );
  OAI222_X1 U10028 ( .A1(n8906), .A2(n8477), .B1(P2_U3152), .B2(n8476), .C1(
        n8904), .C2(n8475), .ZN(P2_U3329) );
  INV_X1 U10029 ( .A(n10087), .ZN(n10003) );
  AOI22_X1 U10030 ( .A1(n10044), .A2(n10043), .B1(n10036), .B2(n10102), .ZN(
        n10026) );
  NAND2_X1 U10031 ( .A1(n10098), .A2(n10057), .ZN(n8483) );
  NAND2_X1 U10032 ( .A1(n10013), .A2(n8484), .ZN(n8485) );
  INV_X1 U10033 ( .A(n10092), .ZN(n10018) );
  NAND2_X1 U10034 ( .A1(n9996), .A2(n9973), .ZN(n8487) );
  NAND2_X1 U10035 ( .A1(n9953), .A2(n9961), .ZN(n9952) );
  NAND2_X1 U10036 ( .A1(n9952), .A2(n8488), .ZN(n9936) );
  NAND2_X1 U10037 ( .A1(n9936), .A2(n9943), .ZN(n9935) );
  NAND2_X1 U10038 ( .A1(n9935), .A2(n8489), .ZN(n9917) );
  OR2_X2 U10039 ( .A1(n9917), .A2(n9922), .ZN(n9918) );
  INV_X1 U10040 ( .A(n10065), .ZN(n9932) );
  NAND2_X1 U10041 ( .A1(n7093), .A2(n10368), .ZN(n10401) );
  NAND2_X1 U10042 ( .A1(n10004), .A2(n8500), .ZN(n9985) );
  NAND2_X1 U10043 ( .A1(n9942), .A2(n8505), .ZN(n9947) );
  NAND3_X1 U10044 ( .A1(n9947), .A2(n9922), .A3(n9923), .ZN(n9921) );
  NAND2_X1 U10045 ( .A1(n9921), .A2(n8506), .ZN(n8508) );
  AND2_X1 U10046 ( .A1(n8509), .A2(P1_B_REG_SCAN_IN), .ZN(n8510) );
  NOR2_X1 U10047 ( .A1(n10338), .A2(n8510), .ZN(n9908) );
  INV_X1 U10048 ( .A(n8511), .ZN(n8512) );
  INV_X1 U10049 ( .A(n10102), .ZN(n10050) );
  NAND2_X1 U10050 ( .A1(n10046), .A2(n10032), .ZN(n10027) );
  INV_X1 U10051 ( .A(n9928), .ZN(n8514) );
  INV_X1 U10052 ( .A(n8515), .ZN(n8867) );
  NOR2_X1 U10053 ( .A1(n10438), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n8516) );
  INV_X1 U10054 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10395) );
  AOI22_X1 U10055 ( .A1(n10395), .A2(keyinput191), .B1(keyinput175), .B2(n5125), .ZN(n8517) );
  OAI221_X1 U10056 ( .B1(n10395), .B2(keyinput191), .C1(n5125), .C2(
        keyinput175), .A(n8517), .ZN(n8526) );
  INV_X1 U10057 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n10456) );
  AOI22_X1 U10058 ( .A1(n7300), .A2(keyinput200), .B1(keyinput138), .B2(n10456), .ZN(n8518) );
  OAI221_X1 U10059 ( .B1(n7300), .B2(keyinput200), .C1(n10456), .C2(
        keyinput138), .A(n8518), .ZN(n8525) );
  INV_X1 U10060 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n10452) );
  AOI22_X1 U10061 ( .A1(n8520), .A2(keyinput211), .B1(keyinput254), .B2(n10452), .ZN(n8519) );
  OAI221_X1 U10062 ( .B1(n8520), .B2(keyinput211), .C1(n10452), .C2(
        keyinput254), .A(n8519), .ZN(n8524) );
  AOI22_X1 U10063 ( .A1(n9674), .A2(keyinput169), .B1(n8522), .B2(keyinput237), 
        .ZN(n8521) );
  OAI221_X1 U10064 ( .B1(n9674), .B2(keyinput169), .C1(n8522), .C2(keyinput237), .A(n8521), .ZN(n8523) );
  NOR4_X1 U10065 ( .A1(n8526), .A2(n8525), .A3(n8524), .A4(n8523), .ZN(n8573)
         );
  AOI22_X1 U10066 ( .A1(n8756), .A2(keyinput228), .B1(keyinput186), .B2(n10533), .ZN(n8527) );
  OAI221_X1 U10067 ( .B1(n8756), .B2(keyinput228), .C1(n10533), .C2(
        keyinput186), .A(n8527), .ZN(n8535) );
  INV_X1 U10068 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n10358) );
  AOI22_X1 U10069 ( .A1(n10358), .A2(keyinput131), .B1(n8847), .B2(keyinput189), .ZN(n8528) );
  OAI221_X1 U10070 ( .B1(n10358), .B2(keyinput131), .C1(n8847), .C2(
        keyinput189), .A(n8528), .ZN(n8534) );
  XNOR2_X1 U10071 ( .A(P1_REG2_REG_29__SCAN_IN), .B(keyinput158), .ZN(n8532)
         );
  XNOR2_X1 U10072 ( .A(P2_IR_REG_10__SCAN_IN), .B(keyinput209), .ZN(n8531) );
  XNOR2_X1 U10073 ( .A(P2_IR_REG_16__SCAN_IN), .B(keyinput235), .ZN(n8530) );
  XNOR2_X1 U10074 ( .A(SI_0_), .B(keyinput213), .ZN(n8529) );
  NAND4_X1 U10075 ( .A1(n8532), .A2(n8531), .A3(n8530), .A4(n8529), .ZN(n8533)
         );
  NOR3_X1 U10076 ( .A1(n8535), .A2(n8534), .A3(n8533), .ZN(n8572) );
  AOI22_X1 U10077 ( .A1(n7923), .A2(keyinput222), .B1(keyinput171), .B2(n5754), 
        .ZN(n8536) );
  OAI221_X1 U10078 ( .B1(n7923), .B2(keyinput222), .C1(n5754), .C2(keyinput171), .A(n8536), .ZN(n8547) );
  INV_X1 U10079 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n10453) );
  AOI22_X1 U10080 ( .A1(n9608), .A2(keyinput144), .B1(n10453), .B2(keyinput218), .ZN(n8537) );
  OAI221_X1 U10081 ( .B1(n9608), .B2(keyinput144), .C1(n10453), .C2(
        keyinput218), .A(n8537), .ZN(n8546) );
  AOI22_X1 U10082 ( .A1(n10583), .A2(keyinput206), .B1(n8539), .B2(keyinput201), .ZN(n8538) );
  OAI221_X1 U10083 ( .B1(n10583), .B2(keyinput206), .C1(n8539), .C2(
        keyinput201), .A(n8538), .ZN(n8545) );
  XOR2_X1 U10084 ( .A(n5467), .B(keyinput221), .Z(n8543) );
  XNOR2_X1 U10085 ( .A(P2_IR_REG_11__SCAN_IN), .B(keyinput163), .ZN(n8542) );
  XNOR2_X1 U10086 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput252), .ZN(n8541) );
  XNOR2_X1 U10087 ( .A(P2_IR_REG_25__SCAN_IN), .B(keyinput134), .ZN(n8540) );
  NAND4_X1 U10088 ( .A1(n8543), .A2(n8542), .A3(n8541), .A4(n8540), .ZN(n8544)
         );
  NOR4_X1 U10089 ( .A1(n8547), .A2(n8546), .A3(n8545), .A4(n8544), .ZN(n8571)
         );
  INV_X1 U10090 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8549) );
  AOI22_X1 U10091 ( .A1(n8549), .A2(keyinput149), .B1(n10359), .B2(keyinput247), .ZN(n8548) );
  OAI221_X1 U10092 ( .B1(n8549), .B2(keyinput149), .C1(n10359), .C2(
        keyinput247), .A(n8548), .ZN(n8556) );
  AOI22_X1 U10093 ( .A1(n8697), .A2(keyinput190), .B1(keyinput137), .B2(n8551), 
        .ZN(n8550) );
  OAI221_X1 U10094 ( .B1(n8697), .B2(keyinput190), .C1(n8551), .C2(keyinput137), .A(n8550), .ZN(n8555) );
  AOI22_X1 U10095 ( .A1(n9805), .A2(keyinput181), .B1(n8553), .B2(keyinput176), 
        .ZN(n8552) );
  OAI221_X1 U10096 ( .B1(n9805), .B2(keyinput181), .C1(n8553), .C2(keyinput176), .A(n8552), .ZN(n8554) );
  NOR3_X1 U10097 ( .A1(n8556), .A2(n8555), .A3(n8554), .ZN(n8569) );
  INV_X1 U10098 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n8557) );
  XNOR2_X1 U10099 ( .A(keyinput198), .B(n8557), .ZN(n8559) );
  INV_X1 U10100 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10178) );
  XNOR2_X1 U10101 ( .A(keyinput227), .B(n10178), .ZN(n8558) );
  NOR2_X1 U10102 ( .A1(n8559), .A2(n8558), .ZN(n8568) );
  AOI22_X1 U10103 ( .A1(P1_D_REG_0__SCAN_IN), .A2(keyinput174), .B1(n8817), 
        .B2(keyinput244), .ZN(n8560) );
  OAI221_X1 U10104 ( .B1(P1_D_REG_0__SCAN_IN), .B2(keyinput174), .C1(n8817), 
        .C2(keyinput244), .A(n8560), .ZN(n8563) );
  AOI22_X1 U10105 ( .A1(P2_REG0_REG_31__SCAN_IN), .A2(keyinput150), .B1(
        P2_IR_REG_23__SCAN_IN), .B2(keyinput128), .ZN(n8561) );
  OAI221_X1 U10106 ( .B1(P2_REG0_REG_31__SCAN_IN), .B2(keyinput150), .C1(
        P2_IR_REG_23__SCAN_IN), .C2(keyinput128), .A(n8561), .ZN(n8562) );
  NOR2_X1 U10107 ( .A1(n8563), .A2(n8562), .ZN(n8567) );
  AOI22_X1 U10108 ( .A1(n9231), .A2(keyinput133), .B1(n9194), .B2(keyinput185), 
        .ZN(n8564) );
  OAI221_X1 U10109 ( .B1(n9231), .B2(keyinput133), .C1(n9194), .C2(keyinput185), .A(n8564), .ZN(n8565) );
  INV_X1 U10110 ( .A(n8565), .ZN(n8566) );
  AND4_X1 U10111 ( .A1(n8569), .A2(n8568), .A3(n8567), .A4(n8566), .ZN(n8570)
         );
  NAND4_X1 U10112 ( .A1(n8573), .A2(n8572), .A3(n8571), .A4(n8570), .ZN(n8648)
         );
  AOI22_X1 U10113 ( .A1(P2_D_REG_15__SCAN_IN), .A2(keyinput183), .B1(
        P2_D_REG_13__SCAN_IN), .B2(keyinput147), .ZN(n8574) );
  OAI221_X1 U10114 ( .B1(P2_D_REG_15__SCAN_IN), .B2(keyinput183), .C1(
        P2_D_REG_13__SCAN_IN), .C2(keyinput147), .A(n8574), .ZN(n8581) );
  AOI22_X1 U10115 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(keyinput156), .B1(SI_1_), 
        .B2(keyinput199), .ZN(n8575) );
  OAI221_X1 U10116 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(keyinput156), .C1(SI_1_), 
        .C2(keyinput199), .A(n8575), .ZN(n8580) );
  AOI22_X1 U10117 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(keyinput159), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(keyinput167), .ZN(n8576) );
  OAI221_X1 U10118 ( .B1(P1_REG3_REG_12__SCAN_IN), .B2(keyinput159), .C1(
        P1_DATAO_REG_9__SCAN_IN), .C2(keyinput167), .A(n8576), .ZN(n8579) );
  AOI22_X1 U10119 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(keyinput210), .B1(
        P1_REG2_REG_20__SCAN_IN), .B2(keyinput196), .ZN(n8577) );
  OAI221_X1 U10120 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(keyinput210), .C1(
        P1_REG2_REG_20__SCAN_IN), .C2(keyinput196), .A(n8577), .ZN(n8578) );
  NOR4_X1 U10121 ( .A1(n8581), .A2(n8580), .A3(n8579), .A4(n8578), .ZN(n8609)
         );
  AOI22_X1 U10122 ( .A1(P1_D_REG_28__SCAN_IN), .A2(keyinput177), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(keyinput219), .ZN(n8582) );
  OAI221_X1 U10123 ( .B1(P1_D_REG_28__SCAN_IN), .B2(keyinput177), .C1(
        P1_DATAO_REG_13__SCAN_IN), .C2(keyinput219), .A(n8582), .ZN(n8589) );
  AOI22_X1 U10124 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(keyinput207), .B1(
        P1_REG1_REG_21__SCAN_IN), .B2(keyinput231), .ZN(n8583) );
  OAI221_X1 U10125 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(keyinput207), .C1(
        P1_REG1_REG_21__SCAN_IN), .C2(keyinput231), .A(n8583), .ZN(n8588) );
  AOI22_X1 U10126 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(keyinput205), .B1(
        P1_REG3_REG_18__SCAN_IN), .B2(keyinput187), .ZN(n8584) );
  OAI221_X1 U10127 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(keyinput205), .C1(
        P1_REG3_REG_18__SCAN_IN), .C2(keyinput187), .A(n8584), .ZN(n8587) );
  AOI22_X1 U10128 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(keyinput182), .B1(
        P1_REG2_REG_24__SCAN_IN), .B2(keyinput245), .ZN(n8585) );
  OAI221_X1 U10129 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(keyinput182), .C1(
        P1_REG2_REG_24__SCAN_IN), .C2(keyinput245), .A(n8585), .ZN(n8586) );
  NOR4_X1 U10130 ( .A1(n8589), .A2(n8588), .A3(n8587), .A4(n8586), .ZN(n8608)
         );
  AOI22_X1 U10131 ( .A1(P1_REG0_REG_5__SCAN_IN), .A2(keyinput239), .B1(
        P1_REG1_REG_19__SCAN_IN), .B2(keyinput145), .ZN(n8590) );
  OAI221_X1 U10132 ( .B1(P1_REG0_REG_5__SCAN_IN), .B2(keyinput239), .C1(
        P1_REG1_REG_19__SCAN_IN), .C2(keyinput145), .A(n8590), .ZN(n8597) );
  AOI22_X1 U10133 ( .A1(P1_REG1_REG_6__SCAN_IN), .A2(keyinput195), .B1(
        P1_REG0_REG_26__SCAN_IN), .B2(keyinput143), .ZN(n8591) );
  OAI221_X1 U10134 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(keyinput195), .C1(
        P1_REG0_REG_26__SCAN_IN), .C2(keyinput143), .A(n8591), .ZN(n8596) );
  AOI22_X1 U10135 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(keyinput160), .B1(
        P1_REG1_REG_5__SCAN_IN), .B2(keyinput161), .ZN(n8592) );
  OAI221_X1 U10136 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(keyinput160), .C1(
        P1_REG1_REG_5__SCAN_IN), .C2(keyinput161), .A(n8592), .ZN(n8595) );
  AOI22_X1 U10137 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(keyinput220), .B1(
        P1_REG3_REG_4__SCAN_IN), .B2(keyinput142), .ZN(n8593) );
  OAI221_X1 U10138 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput220), .C1(
        P1_REG3_REG_4__SCAN_IN), .C2(keyinput142), .A(n8593), .ZN(n8594) );
  NOR4_X1 U10139 ( .A1(n8597), .A2(n8596), .A3(n8595), .A4(n8594), .ZN(n8607)
         );
  AOI22_X1 U10140 ( .A1(P1_REG2_REG_31__SCAN_IN), .A2(keyinput243), .B1(
        P2_REG1_REG_26__SCAN_IN), .B2(keyinput172), .ZN(n8598) );
  OAI221_X1 U10141 ( .B1(P1_REG2_REG_31__SCAN_IN), .B2(keyinput243), .C1(
        P2_REG1_REG_26__SCAN_IN), .C2(keyinput172), .A(n8598), .ZN(n8605) );
  AOI22_X1 U10142 ( .A1(P2_REG1_REG_20__SCAN_IN), .A2(keyinput240), .B1(
        P1_D_REG_3__SCAN_IN), .B2(keyinput250), .ZN(n8599) );
  OAI221_X1 U10143 ( .B1(P2_REG1_REG_20__SCAN_IN), .B2(keyinput240), .C1(
        P1_D_REG_3__SCAN_IN), .C2(keyinput250), .A(n8599), .ZN(n8604) );
  AOI22_X1 U10144 ( .A1(P2_D_REG_21__SCAN_IN), .A2(keyinput165), .B1(
        P2_D_REG_1__SCAN_IN), .B2(keyinput251), .ZN(n8600) );
  OAI221_X1 U10145 ( .B1(P2_D_REG_21__SCAN_IN), .B2(keyinput165), .C1(
        P2_D_REG_1__SCAN_IN), .C2(keyinput251), .A(n8600), .ZN(n8603) );
  AOI22_X1 U10146 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(keyinput146), .B1(SI_17_), .B2(keyinput255), .ZN(n8601) );
  OAI221_X1 U10147 ( .B1(P1_DATAO_REG_7__SCAN_IN), .B2(keyinput146), .C1(
        SI_17_), .C2(keyinput255), .A(n8601), .ZN(n8602) );
  NOR4_X1 U10148 ( .A1(n8605), .A2(n8604), .A3(n8603), .A4(n8602), .ZN(n8606)
         );
  NAND4_X1 U10149 ( .A1(n8609), .A2(n8608), .A3(n8607), .A4(n8606), .ZN(n8647)
         );
  AOI22_X1 U10150 ( .A1(P2_REG2_REG_24__SCAN_IN), .A2(keyinput130), .B1(SI_28_), .B2(keyinput212), .ZN(n8610) );
  OAI221_X1 U10151 ( .B1(P2_REG2_REG_24__SCAN_IN), .B2(keyinput130), .C1(
        SI_28_), .C2(keyinput212), .A(n8610), .ZN(n8617) );
  AOI22_X1 U10152 ( .A1(P1_D_REG_2__SCAN_IN), .A2(keyinput238), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(keyinput132), .ZN(n8611) );
  OAI221_X1 U10153 ( .B1(P1_D_REG_2__SCAN_IN), .B2(keyinput238), .C1(
        P1_DATAO_REG_19__SCAN_IN), .C2(keyinput132), .A(n8611), .ZN(n8616) );
  AOI22_X1 U10154 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(keyinput170), .B1(SI_13_), 
        .B2(keyinput151), .ZN(n8612) );
  OAI221_X1 U10155 ( .B1(P2_IR_REG_12__SCAN_IN), .B2(keyinput170), .C1(SI_13_), 
        .C2(keyinput151), .A(n8612), .ZN(n8615) );
  AOI22_X1 U10156 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(keyinput233), .B1(
        P1_IR_REG_28__SCAN_IN), .B2(keyinput208), .ZN(n8613) );
  OAI221_X1 U10157 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput233), .C1(
        P1_IR_REG_28__SCAN_IN), .C2(keyinput208), .A(n8613), .ZN(n8614) );
  NOR4_X1 U10158 ( .A1(n8617), .A2(n8616), .A3(n8615), .A4(n8614), .ZN(n8645)
         );
  AOI22_X1 U10159 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(keyinput236), .B1(SI_21_), .B2(keyinput193), .ZN(n8618) );
  OAI221_X1 U10160 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(keyinput236), .C1(
        SI_21_), .C2(keyinput193), .A(n8618), .ZN(n8625) );
  AOI22_X1 U10161 ( .A1(P2_D_REG_3__SCAN_IN), .A2(keyinput232), .B1(
        P1_REG0_REG_20__SCAN_IN), .B2(keyinput226), .ZN(n8619) );
  OAI221_X1 U10162 ( .B1(P2_D_REG_3__SCAN_IN), .B2(keyinput232), .C1(
        P1_REG0_REG_20__SCAN_IN), .C2(keyinput226), .A(n8619), .ZN(n8624) );
  AOI22_X1 U10163 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(keyinput178), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(keyinput216), .ZN(n8620) );
  OAI221_X1 U10164 ( .B1(P1_DATAO_REG_8__SCAN_IN), .B2(keyinput178), .C1(
        P1_DATAO_REG_23__SCAN_IN), .C2(keyinput216), .A(n8620), .ZN(n8623) );
  AOI22_X1 U10165 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(keyinput162), .B1(SI_27_), .B2(keyinput154), .ZN(n8621) );
  OAI221_X1 U10166 ( .B1(P2_DATAO_REG_9__SCAN_IN), .B2(keyinput162), .C1(
        SI_27_), .C2(keyinput154), .A(n8621), .ZN(n8622) );
  NOR4_X1 U10167 ( .A1(n8625), .A2(n8624), .A3(n8623), .A4(n8622), .ZN(n8644)
         );
  AOI22_X1 U10168 ( .A1(P1_REG2_REG_26__SCAN_IN), .A2(keyinput215), .B1(
        P1_D_REG_20__SCAN_IN), .B2(keyinput242), .ZN(n8626) );
  OAI221_X1 U10169 ( .B1(P1_REG2_REG_26__SCAN_IN), .B2(keyinput215), .C1(
        P1_D_REG_20__SCAN_IN), .C2(keyinput242), .A(n8626), .ZN(n8633) );
  AOI22_X1 U10170 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(keyinput197), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(keyinput234), .ZN(n8627) );
  OAI221_X1 U10171 ( .B1(P2_DATAO_REG_16__SCAN_IN), .B2(keyinput197), .C1(
        P1_DATAO_REG_17__SCAN_IN), .C2(keyinput234), .A(n8627), .ZN(n8632) );
  AOI22_X1 U10172 ( .A1(P1_REG1_REG_9__SCAN_IN), .A2(keyinput166), .B1(
        P1_REG1_REG_10__SCAN_IN), .B2(keyinput249), .ZN(n8628) );
  OAI221_X1 U10173 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(keyinput166), .C1(
        P1_REG1_REG_10__SCAN_IN), .C2(keyinput249), .A(n8628), .ZN(n8631) );
  AOI22_X1 U10174 ( .A1(P2_REG0_REG_24__SCAN_IN), .A2(keyinput225), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(keyinput241), .ZN(n8629) );
  OAI221_X1 U10175 ( .B1(P2_REG0_REG_24__SCAN_IN), .B2(keyinput225), .C1(
        P1_DATAO_REG_22__SCAN_IN), .C2(keyinput241), .A(n8629), .ZN(n8630) );
  NOR4_X1 U10176 ( .A1(n8633), .A2(n8632), .A3(n8631), .A4(n8630), .ZN(n8643)
         );
  AOI22_X1 U10177 ( .A1(P1_REG0_REG_4__SCAN_IN), .A2(keyinput168), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(keyinput248), .ZN(n8634) );
  OAI221_X1 U10178 ( .B1(P1_REG0_REG_4__SCAN_IN), .B2(keyinput168), .C1(
        P2_DATAO_REG_7__SCAN_IN), .C2(keyinput248), .A(n8634), .ZN(n8641) );
  AOI22_X1 U10179 ( .A1(P1_D_REG_5__SCAN_IN), .A2(keyinput192), .B1(SI_25_), 
        .B2(keyinput202), .ZN(n8635) );
  OAI221_X1 U10180 ( .B1(P1_D_REG_5__SCAN_IN), .B2(keyinput192), .C1(SI_25_), 
        .C2(keyinput202), .A(n8635), .ZN(n8640) );
  AOI22_X1 U10181 ( .A1(P2_REG2_REG_22__SCAN_IN), .A2(keyinput188), .B1(
        P1_D_REG_11__SCAN_IN), .B2(keyinput184), .ZN(n8636) );
  OAI221_X1 U10182 ( .B1(P2_REG2_REG_22__SCAN_IN), .B2(keyinput188), .C1(
        P1_D_REG_11__SCAN_IN), .C2(keyinput184), .A(n8636), .ZN(n8639) );
  AOI22_X1 U10183 ( .A1(P2_REG2_REG_1__SCAN_IN), .A2(keyinput140), .B1(
        P2_REG1_REG_16__SCAN_IN), .B2(keyinput179), .ZN(n8637) );
  OAI221_X1 U10184 ( .B1(P2_REG2_REG_1__SCAN_IN), .B2(keyinput140), .C1(
        P2_REG1_REG_16__SCAN_IN), .C2(keyinput179), .A(n8637), .ZN(n8638) );
  NOR4_X1 U10185 ( .A1(n8641), .A2(n8640), .A3(n8639), .A4(n8638), .ZN(n8642)
         );
  NAND4_X1 U10186 ( .A1(n8645), .A2(n8644), .A3(n8643), .A4(n8642), .ZN(n8646)
         );
  NOR3_X1 U10187 ( .A1(n8648), .A2(n8647), .A3(n8646), .ZN(n8679) );
  INV_X1 U10188 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10423) );
  AOI22_X1 U10189 ( .A1(n10423), .A2(keyinput204), .B1(keyinput139), .B2(n7719), .ZN(n8649) );
  OAI221_X1 U10190 ( .B1(n10423), .B2(keyinput204), .C1(n7719), .C2(
        keyinput139), .A(n8649), .ZN(n8658) );
  INV_X1 U10191 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10357) );
  INV_X1 U10192 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n8651) );
  AOI22_X1 U10193 ( .A1(n10357), .A2(keyinput224), .B1(keyinput246), .B2(n8651), .ZN(n8650) );
  OAI221_X1 U10194 ( .B1(n10357), .B2(keyinput224), .C1(n8651), .C2(
        keyinput246), .A(n8650), .ZN(n8657) );
  AOI22_X1 U10195 ( .A1(n10536), .A2(keyinput180), .B1(n8653), .B2(keyinput203), .ZN(n8652) );
  OAI221_X1 U10196 ( .B1(n10536), .B2(keyinput180), .C1(n8653), .C2(
        keyinput203), .A(n8652), .ZN(n8656) );
  INV_X1 U10197 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10289) );
  AOI22_X1 U10198 ( .A1(n8693), .A2(keyinput129), .B1(keyinput217), .B2(n10289), .ZN(n8654) );
  OAI221_X1 U10199 ( .B1(n8693), .B2(keyinput129), .C1(n10289), .C2(
        keyinput217), .A(n8654), .ZN(n8655) );
  NOR4_X1 U10200 ( .A1(n8658), .A2(n8657), .A3(n8656), .A4(n8655), .ZN(n8678)
         );
  AOI22_X1 U10201 ( .A1(n5164), .A2(keyinput230), .B1(n5895), .B2(keyinput135), 
        .ZN(n8659) );
  OAI221_X1 U10202 ( .B1(n5164), .B2(keyinput230), .C1(n5895), .C2(keyinput135), .A(n8659), .ZN(n8667) );
  AOI22_X1 U10203 ( .A1(n7702), .A2(keyinput148), .B1(n8684), .B2(keyinput157), 
        .ZN(n8660) );
  OAI221_X1 U10204 ( .B1(n7702), .B2(keyinput148), .C1(n8684), .C2(keyinput157), .A(n8660), .ZN(n8666) );
  INV_X1 U10205 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n10457) );
  AOI22_X1 U10206 ( .A1(n8662), .A2(keyinput152), .B1(keyinput253), .B2(n10457), .ZN(n8661) );
  OAI221_X1 U10207 ( .B1(n8662), .B2(keyinput152), .C1(n10457), .C2(
        keyinput253), .A(n8661), .ZN(n8665) );
  INV_X1 U10208 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10576) );
  AOI22_X1 U10209 ( .A1(n10576), .A2(keyinput173), .B1(n8748), .B2(keyinput194), .ZN(n8663) );
  OAI221_X1 U10210 ( .B1(n10576), .B2(keyinput173), .C1(n8748), .C2(
        keyinput194), .A(n8663), .ZN(n8664) );
  NOR4_X1 U10211 ( .A1(n8667), .A2(n8666), .A3(n8665), .A4(n8664), .ZN(n8677)
         );
  AOI22_X1 U10212 ( .A1(P2_REG0_REG_5__SCAN_IN), .A2(keyinput214), .B1(
        P2_REG3_REG_8__SCAN_IN), .B2(keyinput136), .ZN(n8668) );
  OAI221_X1 U10213 ( .B1(P2_REG0_REG_5__SCAN_IN), .B2(keyinput214), .C1(
        P2_REG3_REG_8__SCAN_IN), .C2(keyinput136), .A(n8668), .ZN(n8675) );
  AOI22_X1 U10214 ( .A1(P1_REG1_REG_13__SCAN_IN), .A2(keyinput155), .B1(
        P1_REG2_REG_27__SCAN_IN), .B2(keyinput223), .ZN(n8669) );
  OAI221_X1 U10215 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(keyinput155), .C1(
        P1_REG2_REG_27__SCAN_IN), .C2(keyinput223), .A(n8669), .ZN(n8674) );
  AOI22_X1 U10216 ( .A1(P2_REG0_REG_30__SCAN_IN), .A2(keyinput164), .B1(
        P1_REG0_REG_24__SCAN_IN), .B2(keyinput141), .ZN(n8670) );
  OAI221_X1 U10217 ( .B1(P2_REG0_REG_30__SCAN_IN), .B2(keyinput164), .C1(
        P1_REG0_REG_24__SCAN_IN), .C2(keyinput141), .A(n8670), .ZN(n8673) );
  AOI22_X1 U10218 ( .A1(P1_REG0_REG_12__SCAN_IN), .A2(keyinput229), .B1(
        P1_REG2_REG_28__SCAN_IN), .B2(keyinput153), .ZN(n8671) );
  OAI221_X1 U10219 ( .B1(P1_REG0_REG_12__SCAN_IN), .B2(keyinput229), .C1(
        P1_REG2_REG_28__SCAN_IN), .C2(keyinput153), .A(n8671), .ZN(n8672) );
  NOR4_X1 U10220 ( .A1(n8675), .A2(n8674), .A3(n8673), .A4(n8672), .ZN(n8676)
         );
  NAND4_X1 U10221 ( .A1(n8679), .A2(n8678), .A3(n8677), .A4(n8676), .ZN(n8714)
         );
  INV_X1 U10222 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10356) );
  AOI22_X1 U10223 ( .A1(n10356), .A2(keyinput49), .B1(keyinput105), .B2(n8681), 
        .ZN(n8680) );
  OAI221_X1 U10224 ( .B1(n10356), .B2(keyinput49), .C1(n8681), .C2(keyinput105), .A(n8680), .ZN(n8689) );
  AOI22_X1 U10225 ( .A1(n9470), .A2(keyinput60), .B1(n5443), .B2(keyinput108), 
        .ZN(n8682) );
  OAI221_X1 U10226 ( .B1(n9470), .B2(keyinput60), .C1(n5443), .C2(keyinput108), 
        .A(n8682), .ZN(n8688) );
  AOI22_X1 U10227 ( .A1(n8684), .A2(keyinput29), .B1(keyinput63), .B2(n10395), 
        .ZN(n8683) );
  OAI221_X1 U10228 ( .B1(n8684), .B2(keyinput29), .C1(n10395), .C2(keyinput63), 
        .A(n8683), .ZN(n8687) );
  AOI22_X1 U10229 ( .A1(n10178), .A2(keyinput99), .B1(keyinput10), .B2(n10456), 
        .ZN(n8685) );
  OAI221_X1 U10230 ( .B1(n10178), .B2(keyinput99), .C1(n10456), .C2(keyinput10), .A(n8685), .ZN(n8686) );
  NOR4_X1 U10231 ( .A1(n8689), .A2(n8688), .A3(n8687), .A4(n8686), .ZN(n8713)
         );
  AOI22_X1 U10232 ( .A1(n7923), .A2(keyinput94), .B1(keyinput36), .B2(n8691), 
        .ZN(n8690) );
  OAI221_X1 U10233 ( .B1(n7923), .B2(keyinput94), .C1(n8691), .C2(keyinput36), 
        .A(n8690), .ZN(n8702) );
  AOI22_X1 U10234 ( .A1(n8694), .A2(keyinput28), .B1(n8693), .B2(keyinput1), 
        .ZN(n8692) );
  OAI221_X1 U10235 ( .B1(n8694), .B2(keyinput28), .C1(n8693), .C2(keyinput1), 
        .A(n8692), .ZN(n8701) );
  INV_X1 U10236 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10383) );
  AOI22_X1 U10237 ( .A1(n10383), .A2(keyinput40), .B1(n6696), .B2(keyinput46), 
        .ZN(n8695) );
  OAI221_X1 U10238 ( .B1(n10383), .B2(keyinput40), .C1(n6696), .C2(keyinput46), 
        .A(n8695), .ZN(n8700) );
  AOI22_X1 U10239 ( .A1(n8698), .A2(keyinput88), .B1(keyinput62), .B2(n8697), 
        .ZN(n8696) );
  OAI221_X1 U10240 ( .B1(n8698), .B2(keyinput88), .C1(n8697), .C2(keyinput62), 
        .A(n8696), .ZN(n8699) );
  NOR4_X1 U10241 ( .A1(n8702), .A2(n8701), .A3(n8700), .A4(n8699), .ZN(n8712)
         );
  AOI22_X1 U10242 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(keyinput93), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(keyinput83), .ZN(n8703) );
  OAI221_X1 U10243 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(keyinput93), .C1(
        P1_DATAO_REG_14__SCAN_IN), .C2(keyinput83), .A(n8703), .ZN(n8710) );
  AOI22_X1 U10244 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(keyinput50), .B1(SI_21_), 
        .B2(keyinput65), .ZN(n8704) );
  OAI221_X1 U10245 ( .B1(P1_DATAO_REG_8__SCAN_IN), .B2(keyinput50), .C1(SI_21_), .C2(keyinput65), .A(n8704), .ZN(n8709) );
  AOI22_X1 U10246 ( .A1(P1_D_REG_14__SCAN_IN), .A2(keyinput119), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(keyinput120), .ZN(n8705) );
  OAI221_X1 U10247 ( .B1(P1_D_REG_14__SCAN_IN), .B2(keyinput119), .C1(
        P2_DATAO_REG_7__SCAN_IN), .C2(keyinput120), .A(n8705), .ZN(n8708) );
  AOI22_X1 U10248 ( .A1(P2_REG0_REG_24__SCAN_IN), .A2(keyinput97), .B1(
        P1_REG3_REG_22__SCAN_IN), .B2(keyinput7), .ZN(n8706) );
  OAI221_X1 U10249 ( .B1(P2_REG0_REG_24__SCAN_IN), .B2(keyinput97), .C1(
        P1_REG3_REG_22__SCAN_IN), .C2(keyinput7), .A(n8706), .ZN(n8707) );
  NOR4_X1 U10250 ( .A1(n8710), .A2(n8709), .A3(n8708), .A4(n8707), .ZN(n8711)
         );
  NAND4_X1 U10251 ( .A1(n8714), .A2(n8713), .A3(n8712), .A4(n8711), .ZN(n8861)
         );
  OAI22_X1 U10252 ( .A1(P1_D_REG_3__SCAN_IN), .A2(keyinput122), .B1(keyinput51), .B2(P2_REG1_REG_16__SCAN_IN), .ZN(n8715) );
  AOI221_X1 U10253 ( .B1(P1_D_REG_3__SCAN_IN), .B2(keyinput122), .C1(
        P2_REG1_REG_16__SCAN_IN), .C2(keyinput51), .A(n8715), .ZN(n8722) );
  OAI22_X1 U10254 ( .A1(SI_27_), .A2(keyinput26), .B1(keyinput82), .B2(
        P2_ADDR_REG_3__SCAN_IN), .ZN(n8716) );
  AOI221_X1 U10255 ( .B1(SI_27_), .B2(keyinput26), .C1(P2_ADDR_REG_3__SCAN_IN), 
        .C2(keyinput82), .A(n8716), .ZN(n8721) );
  OAI22_X1 U10256 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(keyinput124), .B1(
        P2_REG1_REG_12__SCAN_IN), .B2(keyinput11), .ZN(n8717) );
  AOI221_X1 U10257 ( .B1(P1_IR_REG_26__SCAN_IN), .B2(keyinput124), .C1(
        keyinput11), .C2(P2_REG1_REG_12__SCAN_IN), .A(n8717), .ZN(n8720) );
  OAI22_X1 U10258 ( .A1(P1_D_REG_11__SCAN_IN), .A2(keyinput56), .B1(
        P2_REG2_REG_24__SCAN_IN), .B2(keyinput2), .ZN(n8718) );
  AOI221_X1 U10259 ( .B1(P1_D_REG_11__SCAN_IN), .B2(keyinput56), .C1(keyinput2), .C2(P2_REG2_REG_24__SCAN_IN), .A(n8718), .ZN(n8719) );
  NAND4_X1 U10260 ( .A1(n8722), .A2(n8721), .A3(n8720), .A4(n8719), .ZN(n8775)
         );
  OAI22_X1 U10261 ( .A1(SI_28_), .A2(keyinput84), .B1(keyinput19), .B2(
        P2_D_REG_13__SCAN_IN), .ZN(n8723) );
  AOI221_X1 U10262 ( .B1(SI_28_), .B2(keyinput84), .C1(P2_D_REG_13__SCAN_IN), 
        .C2(keyinput19), .A(n8723), .ZN(n8730) );
  OAI22_X1 U10263 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(keyinput42), .B1(keyinput9), .B2(P2_REG2_REG_23__SCAN_IN), .ZN(n8724) );
  AOI221_X1 U10264 ( .B1(P2_IR_REG_12__SCAN_IN), .B2(keyinput42), .C1(
        P2_REG2_REG_23__SCAN_IN), .C2(keyinput9), .A(n8724), .ZN(n8729) );
  OAI22_X1 U10265 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(keyinput24), .B1(
        P1_REG0_REG_5__SCAN_IN), .B2(keyinput111), .ZN(n8725) );
  AOI221_X1 U10266 ( .B1(P2_DATAO_REG_15__SCAN_IN), .B2(keyinput24), .C1(
        keyinput111), .C2(P1_REG0_REG_5__SCAN_IN), .A(n8725), .ZN(n8728) );
  OAI22_X1 U10267 ( .A1(SI_17_), .A2(keyinput127), .B1(P1_DATAO_REG_9__SCAN_IN), .B2(keyinput39), .ZN(n8726) );
  AOI221_X1 U10268 ( .B1(SI_17_), .B2(keyinput127), .C1(keyinput39), .C2(
        P1_DATAO_REG_9__SCAN_IN), .A(n8726), .ZN(n8727) );
  NAND4_X1 U10269 ( .A1(n8730), .A2(n8729), .A3(n8728), .A4(n8727), .ZN(n8774)
         );
  AOI22_X1 U10270 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(keyinput54), .B1(
        P1_REG3_REG_26__SCAN_IN), .B2(keyinput53), .ZN(n8731) );
  OAI221_X1 U10271 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(keyinput54), .C1(
        P1_REG3_REG_26__SCAN_IN), .C2(keyinput53), .A(n8731), .ZN(n8738) );
  AOI22_X1 U10272 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(keyinput91), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(keyinput48), .ZN(n8732) );
  OAI221_X1 U10273 ( .B1(P1_DATAO_REG_13__SCAN_IN), .B2(keyinput91), .C1(
        P1_DATAO_REG_24__SCAN_IN), .C2(keyinput48), .A(n8732), .ZN(n8737) );
  AOI22_X1 U10274 ( .A1(P1_REG2_REG_25__SCAN_IN), .A2(keyinput70), .B1(
        P1_REG3_REG_16__SCAN_IN), .B2(keyinput21), .ZN(n8733) );
  OAI221_X1 U10275 ( .B1(P1_REG2_REG_25__SCAN_IN), .B2(keyinput70), .C1(
        P1_REG3_REG_16__SCAN_IN), .C2(keyinput21), .A(n8733), .ZN(n8736) );
  AOI22_X1 U10276 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(keyinput45), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(keyinput75), .ZN(n8734) );
  OAI221_X1 U10277 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(keyinput45), .C1(
        P1_DATAO_REG_15__SCAN_IN), .C2(keyinput75), .A(n8734), .ZN(n8735) );
  NOR4_X1 U10278 ( .A1(n8738), .A2(n8737), .A3(n8736), .A4(n8735), .ZN(n8772)
         );
  AOI22_X1 U10279 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(keyinput118), .B1(
        P1_D_REG_22__SCAN_IN), .B2(keyinput3), .ZN(n8739) );
  OAI221_X1 U10280 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(keyinput118), .C1(
        P1_D_REG_22__SCAN_IN), .C2(keyinput3), .A(n8739), .ZN(n8746) );
  AOI22_X1 U10281 ( .A1(P2_D_REG_1__SCAN_IN), .A2(keyinput123), .B1(
        P1_D_REG_20__SCAN_IN), .B2(keyinput114), .ZN(n8740) );
  OAI221_X1 U10282 ( .B1(P2_D_REG_1__SCAN_IN), .B2(keyinput123), .C1(
        P1_D_REG_20__SCAN_IN), .C2(keyinput114), .A(n8740), .ZN(n8745) );
  AOI22_X1 U10283 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(keyinput78), .B1(
        P1_REG2_REG_20__SCAN_IN), .B2(keyinput68), .ZN(n8741) );
  OAI221_X1 U10284 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(keyinput78), .C1(
        P1_REG2_REG_20__SCAN_IN), .C2(keyinput68), .A(n8741), .ZN(n8744) );
  AOI22_X1 U10285 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput109), .B1(
        P1_REG3_REG_18__SCAN_IN), .B2(keyinput59), .ZN(n8742) );
  OAI221_X1 U10286 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput109), .C1(
        P1_REG3_REG_18__SCAN_IN), .C2(keyinput59), .A(n8742), .ZN(n8743) );
  NOR4_X1 U10287 ( .A1(n8746), .A2(n8745), .A3(n8744), .A4(n8743), .ZN(n8771)
         );
  AOI22_X1 U10288 ( .A1(n7599), .A2(keyinput27), .B1(keyinput66), .B2(n8748), 
        .ZN(n8747) );
  OAI221_X1 U10289 ( .B1(n7599), .B2(keyinput27), .C1(n8748), .C2(keyinput66), 
        .A(n8747), .ZN(n8760) );
  INV_X1 U10290 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n8750) );
  AOI22_X1 U10291 ( .A1(n5778), .A2(keyinput0), .B1(n8750), .B2(keyinput103), 
        .ZN(n8749) );
  OAI221_X1 U10292 ( .B1(n5778), .B2(keyinput0), .C1(n8750), .C2(keyinput103), 
        .A(n8749), .ZN(n8759) );
  INV_X1 U10293 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n8752) );
  AOI22_X1 U10294 ( .A1(n8753), .A2(keyinput34), .B1(keyinput115), .B2(n8752), 
        .ZN(n8751) );
  OAI221_X1 U10295 ( .B1(n8753), .B2(keyinput34), .C1(n8752), .C2(keyinput115), 
        .A(n8751), .ZN(n8758) );
  INV_X1 U10296 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n8755) );
  AOI22_X1 U10297 ( .A1(n8756), .A2(keyinput100), .B1(n8755), .B2(keyinput101), 
        .ZN(n8754) );
  OAI221_X1 U10298 ( .B1(n8756), .B2(keyinput100), .C1(n8755), .C2(keyinput101), .A(n8754), .ZN(n8757) );
  NOR4_X1 U10299 ( .A1(n8760), .A2(n8759), .A3(n8758), .A4(n8757), .ZN(n8770)
         );
  AOI22_X1 U10300 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(keyinput43), .B1(SI_1_), 
        .B2(keyinput71), .ZN(n8761) );
  OAI221_X1 U10301 ( .B1(P2_IR_REG_24__SCAN_IN), .B2(keyinput43), .C1(SI_1_), 
        .C2(keyinput71), .A(n8761), .ZN(n8768) );
  AOI22_X1 U10302 ( .A1(P2_D_REG_3__SCAN_IN), .A2(keyinput104), .B1(
        P2_IR_REG_25__SCAN_IN), .B2(keyinput6), .ZN(n8762) );
  OAI221_X1 U10303 ( .B1(P2_D_REG_3__SCAN_IN), .B2(keyinput104), .C1(
        P2_IR_REG_25__SCAN_IN), .C2(keyinput6), .A(n8762), .ZN(n8767) );
  AOI22_X1 U10304 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(keyinput69), .B1(n9608), 
        .B2(keyinput16), .ZN(n8763) );
  OAI221_X1 U10305 ( .B1(P2_DATAO_REG_16__SCAN_IN), .B2(keyinput69), .C1(n9608), .C2(keyinput16), .A(n8763), .ZN(n8766) );
  AOI22_X1 U10306 ( .A1(P1_REG0_REG_24__SCAN_IN), .A2(keyinput13), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(keyinput106), .ZN(n8764) );
  OAI221_X1 U10307 ( .B1(P1_REG0_REG_24__SCAN_IN), .B2(keyinput13), .C1(
        P1_DATAO_REG_17__SCAN_IN), .C2(keyinput106), .A(n8764), .ZN(n8765) );
  NOR4_X1 U10308 ( .A1(n8768), .A2(n8767), .A3(n8766), .A4(n8765), .ZN(n8769)
         );
  NAND4_X1 U10309 ( .A1(n8772), .A2(n8771), .A3(n8770), .A4(n8769), .ZN(n8773)
         );
  NOR3_X1 U10310 ( .A1(n8775), .A2(n8774), .A3(n8773), .ZN(n8859) );
  INV_X1 U10311 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n10455) );
  AOI22_X1 U10312 ( .A1(n10533), .A2(keyinput58), .B1(n10455), .B2(keyinput55), 
        .ZN(n8776) );
  OAI221_X1 U10313 ( .B1(n10533), .B2(keyinput58), .C1(n10455), .C2(keyinput55), .A(n8776), .ZN(n8786) );
  INV_X1 U10314 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n8778) );
  AOI22_X1 U10315 ( .A1(n8778), .A2(keyinput87), .B1(n8905), .B2(keyinput113), 
        .ZN(n8777) );
  OAI221_X1 U10316 ( .B1(n8778), .B2(keyinput87), .C1(n8905), .C2(keyinput113), 
        .A(n8777), .ZN(n8785) );
  AOI22_X1 U10317 ( .A1(n10457), .A2(keyinput125), .B1(keyinput126), .B2(
        n10452), .ZN(n8779) );
  OAI221_X1 U10318 ( .B1(n10457), .B2(keyinput125), .C1(n10452), .C2(
        keyinput126), .A(n8779), .ZN(n8784) );
  INV_X1 U10319 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n8782) );
  AOI22_X1 U10320 ( .A1(n8782), .A2(keyinput15), .B1(n8781), .B2(keyinput4), 
        .ZN(n8780) );
  OAI221_X1 U10321 ( .B1(n8782), .B2(keyinput15), .C1(n8781), .C2(keyinput4), 
        .A(n8780), .ZN(n8783) );
  NOR4_X1 U10322 ( .A1(n8786), .A2(n8785), .A3(n8784), .A4(n8783), .ZN(n8836)
         );
  AOI22_X1 U10323 ( .A1(P2_REG1_REG_26__SCAN_IN), .A2(keyinput44), .B1(
        P2_D_REG_23__SCAN_IN), .B2(keyinput90), .ZN(n8787) );
  OAI221_X1 U10324 ( .B1(P2_REG1_REG_26__SCAN_IN), .B2(keyinput44), .C1(
        P2_D_REG_23__SCAN_IN), .C2(keyinput90), .A(n8787), .ZN(n8794) );
  AOI22_X1 U10325 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(keyinput77), .B1(
        P1_REG3_REG_23__SCAN_IN), .B2(keyinput73), .ZN(n8788) );
  OAI221_X1 U10326 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(keyinput77), .C1(
        P1_REG3_REG_23__SCAN_IN), .C2(keyinput73), .A(n8788), .ZN(n8793) );
  AOI22_X1 U10327 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(keyinput52), .B1(
        P1_IR_REG_28__SCAN_IN), .B2(keyinput80), .ZN(n8789) );
  OAI221_X1 U10328 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(keyinput52), .C1(
        P1_IR_REG_28__SCAN_IN), .C2(keyinput80), .A(n8789), .ZN(n8792) );
  AOI22_X1 U10329 ( .A1(P2_REG0_REG_22__SCAN_IN), .A2(keyinput41), .B1(
        P1_D_REG_2__SCAN_IN), .B2(keyinput110), .ZN(n8790) );
  OAI221_X1 U10330 ( .B1(P2_REG0_REG_22__SCAN_IN), .B2(keyinput41), .C1(
        P1_D_REG_2__SCAN_IN), .C2(keyinput110), .A(n8790), .ZN(n8791) );
  NOR4_X1 U10331 ( .A1(n8794), .A2(n8793), .A3(n8792), .A4(n8791), .ZN(n8835)
         );
  INV_X1 U10332 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n10454) );
  AOI22_X1 U10333 ( .A1(n10454), .A2(keyinput37), .B1(n8796), .B2(keyinput23), 
        .ZN(n8795) );
  OAI221_X1 U10334 ( .B1(n10454), .B2(keyinput37), .C1(n8796), .C2(keyinput23), 
        .A(n8795), .ZN(n8801) );
  INV_X1 U10335 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n8799) );
  INV_X1 U10336 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n8798) );
  AOI22_X1 U10337 ( .A1(n8799), .A2(keyinput30), .B1(n8798), .B2(keyinput95), 
        .ZN(n8797) );
  OAI221_X1 U10338 ( .B1(n8799), .B2(keyinput30), .C1(n8798), .C2(keyinput95), 
        .A(n8797), .ZN(n8800) );
  NOR2_X1 U10339 ( .A1(n8801), .A2(n8800), .ZN(n8813) );
  XNOR2_X1 U10340 ( .A(P1_REG3_REG_4__SCAN_IN), .B(keyinput14), .ZN(n8805) );
  XNOR2_X1 U10341 ( .A(P2_IR_REG_10__SCAN_IN), .B(keyinput81), .ZN(n8804) );
  XNOR2_X1 U10342 ( .A(SI_0_), .B(keyinput85), .ZN(n8803) );
  XNOR2_X1 U10343 ( .A(SI_25_), .B(keyinput74), .ZN(n8802) );
  NAND4_X1 U10344 ( .A1(n8805), .A2(n8804), .A3(n8803), .A4(n8802), .ZN(n8811)
         );
  XNOR2_X1 U10345 ( .A(P1_REG0_REG_20__SCAN_IN), .B(keyinput98), .ZN(n8809) );
  XNOR2_X1 U10346 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput92), .ZN(n8808) );
  XNOR2_X1 U10347 ( .A(P2_IR_REG_11__SCAN_IN), .B(keyinput35), .ZN(n8807) );
  XNOR2_X1 U10348 ( .A(P2_IR_REG_16__SCAN_IN), .B(keyinput107), .ZN(n8806) );
  NAND4_X1 U10349 ( .A1(n8809), .A2(n8808), .A3(n8807), .A4(n8806), .ZN(n8810)
         );
  NOR2_X1 U10350 ( .A1(n8811), .A2(n8810), .ZN(n8812) );
  AND2_X1 U10351 ( .A1(n8813), .A2(n8812), .ZN(n8833) );
  AOI22_X1 U10352 ( .A1(n10430), .A2(keyinput67), .B1(keyinput8), .B2(n8815), 
        .ZN(n8814) );
  OAI221_X1 U10353 ( .B1(n10430), .B2(keyinput67), .C1(n8815), .C2(keyinput8), 
        .A(n8814), .ZN(n8819) );
  AOI22_X1 U10354 ( .A1(n10357), .A2(keyinput96), .B1(keyinput116), .B2(n8817), 
        .ZN(n8816) );
  OAI221_X1 U10355 ( .B1(n10357), .B2(keyinput96), .C1(n8817), .C2(keyinput116), .A(n8816), .ZN(n8818) );
  NOR2_X1 U10356 ( .A1(n8819), .A2(n8818), .ZN(n8832) );
  INV_X1 U10357 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n8821) );
  AOI22_X1 U10358 ( .A1(n8821), .A2(keyinput25), .B1(keyinput76), .B2(n10423), 
        .ZN(n8820) );
  OAI221_X1 U10359 ( .B1(n8821), .B2(keyinput25), .C1(n10423), .C2(keyinput76), 
        .A(n8820), .ZN(n8824) );
  AOI22_X1 U10360 ( .A1(n10428), .A2(keyinput33), .B1(n10179), .B2(keyinput121), .ZN(n8822) );
  OAI221_X1 U10361 ( .B1(n10428), .B2(keyinput33), .C1(n10179), .C2(
        keyinput121), .A(n8822), .ZN(n8823) );
  NOR2_X1 U10362 ( .A1(n8824), .A2(n8823), .ZN(n8831) );
  AOI22_X1 U10363 ( .A1(n9194), .A2(keyinput57), .B1(n6867), .B2(keyinput38), 
        .ZN(n8825) );
  OAI221_X1 U10364 ( .B1(n9194), .B2(keyinput57), .C1(n6867), .C2(keyinput38), 
        .A(n8825), .ZN(n8829) );
  INV_X1 U10365 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n8827) );
  AOI22_X1 U10366 ( .A1(n8827), .A2(keyinput117), .B1(n6014), .B2(keyinput31), 
        .ZN(n8826) );
  OAI221_X1 U10367 ( .B1(n8827), .B2(keyinput117), .C1(n6014), .C2(keyinput31), 
        .A(n8826), .ZN(n8828) );
  NOR2_X1 U10368 ( .A1(n8829), .A2(n8828), .ZN(n8830) );
  AND4_X1 U10369 ( .A1(n8833), .A2(n8832), .A3(n8831), .A4(n8830), .ZN(n8834)
         );
  AND3_X1 U10370 ( .A1(n8836), .A2(n8835), .A3(n8834), .ZN(n8858) );
  AOI22_X1 U10371 ( .A1(n9231), .A2(keyinput5), .B1(keyinput112), .B2(n9623), 
        .ZN(n8837) );
  OAI221_X1 U10372 ( .B1(n9231), .B2(keyinput5), .C1(n9623), .C2(keyinput112), 
        .A(n8837), .ZN(n8845) );
  AOI22_X1 U10373 ( .A1(n8839), .A2(keyinput18), .B1(keyinput22), .B2(n9642), 
        .ZN(n8838) );
  OAI221_X1 U10374 ( .B1(n8839), .B2(keyinput18), .C1(n9642), .C2(keyinput22), 
        .A(n8838), .ZN(n8844) );
  INV_X1 U10375 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9889) );
  AOI22_X1 U10376 ( .A1(n5247), .A2(keyinput86), .B1(n9889), .B2(keyinput17), 
        .ZN(n8840) );
  OAI221_X1 U10377 ( .B1(n5247), .B2(keyinput86), .C1(n9889), .C2(keyinput17), 
        .A(n8840), .ZN(n8843) );
  AOI22_X1 U10378 ( .A1(n7682), .A2(keyinput12), .B1(n10289), .B2(keyinput89), 
        .ZN(n8841) );
  OAI221_X1 U10379 ( .B1(n7682), .B2(keyinput12), .C1(n10289), .C2(keyinput89), 
        .A(n8841), .ZN(n8842) );
  NOR4_X1 U10380 ( .A1(n8845), .A2(n8844), .A3(n8843), .A4(n8842), .ZN(n8857)
         );
  AOI22_X1 U10381 ( .A1(n8847), .A2(keyinput61), .B1(keyinput72), .B2(n7300), 
        .ZN(n8846) );
  OAI221_X1 U10382 ( .B1(n8847), .B2(keyinput61), .C1(n7300), .C2(keyinput72), 
        .A(n8846), .ZN(n8855) );
  AOI22_X1 U10383 ( .A1(n7743), .A2(keyinput32), .B1(keyinput102), .B2(n5164), 
        .ZN(n8848) );
  OAI221_X1 U10384 ( .B1(n7743), .B2(keyinput32), .C1(n5164), .C2(keyinput102), 
        .A(n8848), .ZN(n8854) );
  AOI22_X1 U10385 ( .A1(n5125), .A2(keyinput47), .B1(keyinput20), .B2(n7702), 
        .ZN(n8849) );
  OAI221_X1 U10386 ( .B1(n5125), .B2(keyinput47), .C1(n7702), .C2(keyinput20), 
        .A(n8849), .ZN(n8853) );
  INV_X1 U10387 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10361) );
  INV_X1 U10388 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n8851) );
  AOI22_X1 U10389 ( .A1(n10361), .A2(keyinput64), .B1(keyinput79), .B2(n8851), 
        .ZN(n8850) );
  OAI221_X1 U10390 ( .B1(n10361), .B2(keyinput64), .C1(n8851), .C2(keyinput79), 
        .A(n8850), .ZN(n8852) );
  NOR4_X1 U10391 ( .A1(n8855), .A2(n8854), .A3(n8853), .A4(n8852), .ZN(n8856)
         );
  NAND4_X1 U10392 ( .A1(n8859), .A2(n8858), .A3(n8857), .A4(n8856), .ZN(n8860)
         );
  OR2_X1 U10393 ( .A1(n8861), .A2(n8860), .ZN(n8862) );
  NAND2_X1 U10394 ( .A1(n8863), .A2(n8864), .ZN(n8871) );
  AOI22_X1 U10395 ( .A1(n10048), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n8865), 
        .B2(n10345), .ZN(n8866) );
  OAI21_X1 U10396 ( .B1(n8867), .B2(n10256), .A(n8866), .ZN(n8868) );
  AOI21_X1 U10397 ( .B1(n8869), .B2(n10331), .A(n8868), .ZN(n8870) );
  OAI211_X1 U10398 ( .C1(n8872), .C2(n10048), .A(n8871), .B(n8870), .ZN(
        P1_U3355) );
  OAI21_X1 U10399 ( .B1(n8875), .B2(n8874), .A(n8873), .ZN(n8876) );
  NAND2_X1 U10400 ( .A1(n8876), .A2(n9802), .ZN(n8881) );
  OAI22_X1 U10401 ( .A1(n8877), .A2(n9806), .B1(n9804), .B2(n4733), .ZN(n8878)
         );
  AOI21_X1 U10402 ( .B1(n9792), .B2(n8879), .A(n8878), .ZN(n8880) );
  OAI211_X1 U10403 ( .C1(n8882), .C2(n7059), .A(n8881), .B(n8880), .ZN(
        P1_U3235) );
  OAI222_X1 U10404 ( .A1(n8885), .A2(n8884), .B1(n8883), .B2(P1_U3084), .C1(
        n10157), .C2(n8923), .ZN(P1_U3323) );
  NAND3_X1 U10405 ( .A1(n9235), .A2(n8886), .A3(n9272), .ZN(n8887) );
  OAI21_X1 U10406 ( .B1(n8888), .B2(n9240), .A(n8887), .ZN(n8891) );
  INV_X1 U10407 ( .A(n8889), .ZN(n8890) );
  NAND2_X1 U10408 ( .A1(n8891), .A2(n8890), .ZN(n8900) );
  NOR2_X1 U10409 ( .A1(n9230), .A2(n8892), .ZN(n8897) );
  NAND2_X1 U10410 ( .A1(n9224), .A2(n9272), .ZN(n8894) );
  OAI211_X1 U10411 ( .C1(n8895), .C2(n9218), .A(n8894), .B(n8893), .ZN(n8896)
         );
  AOI211_X1 U10412 ( .C1(n8898), .C2(n10593), .A(n8897), .B(n8896), .ZN(n8899)
         );
  OAI211_X1 U10413 ( .C1(n9240), .C2(n8901), .A(n8900), .B(n8899), .ZN(
        P2_U3233) );
  OAI222_X1 U10414 ( .A1(n8906), .A2(n8905), .B1(n8904), .B2(n8903), .C1(n8902), .C2(P2_U3152), .ZN(P2_U3336) );
  NOR2_X1 U10415 ( .A1(n8048), .A2(n9240), .ZN(n8911) );
  NOR3_X1 U10416 ( .A1(n8907), .A2(n9049), .A3(n9223), .ZN(n8910) );
  INV_X1 U10417 ( .A(n8908), .ZN(n8909) );
  OAI21_X1 U10418 ( .B1(n8911), .B2(n8910), .A(n8909), .ZN(n8919) );
  NOR2_X1 U10419 ( .A1(n9230), .A2(n8912), .ZN(n8916) );
  OAI21_X1 U10420 ( .B1(n9247), .B2(n8914), .A(n8913), .ZN(n8915) );
  AOI211_X1 U10421 ( .C1(n8917), .C2(n10593), .A(n8916), .B(n8915), .ZN(n8918)
         );
  OAI211_X1 U10422 ( .C1(n9240), .C2(n8920), .A(n8919), .B(n8918), .ZN(
        P2_U3217) );
  INV_X1 U10423 ( .A(n8921), .ZN(n9108) );
  INV_X1 U10424 ( .A(n8932), .ZN(n8933) );
  NAND2_X1 U10425 ( .A1(n5240), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8924) );
  INV_X1 U10426 ( .A(n9253), .ZN(n8929) );
  NAND2_X1 U10427 ( .A1(n9694), .A2(n4504), .ZN(n8927) );
  NAND2_X1 U10428 ( .A1(n5240), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8926) );
  INV_X1 U10429 ( .A(n9343), .ZN(n8928) );
  OR2_X1 U10430 ( .A1(n9340), .A2(n8928), .ZN(n9118) );
  NAND2_X1 U10431 ( .A1(n8930), .A2(n8929), .ZN(n9115) );
  NAND2_X1 U10432 ( .A1(n9118), .A2(n9115), .ZN(n8969) );
  NOR2_X1 U10433 ( .A1(n8934), .A2(n9121), .ZN(n8935) );
  XNOR2_X1 U10434 ( .A(n8935), .B(n9565), .ZN(n8936) );
  AOI21_X1 U10435 ( .B1(n8938), .B2(n8937), .A(n8936), .ZN(n9128) );
  NOR2_X1 U10436 ( .A1(n8940), .A2(n8939), .ZN(n8947) );
  NOR2_X1 U10437 ( .A1(n8941), .A2(n10468), .ZN(n8946) );
  NOR2_X1 U10438 ( .A1(n8943), .A2(n8942), .ZN(n8944) );
  NAND4_X1 U10439 ( .A1(n8947), .A2(n8946), .A3(n8945), .A4(n8944), .ZN(n8949)
         );
  NOR3_X1 U10440 ( .A1(n8949), .A2(n8948), .A3(n9016), .ZN(n8952) );
  NAND4_X1 U10441 ( .A1(n8952), .A2(n8951), .A3(n8950), .A4(n9021), .ZN(n8954)
         );
  NOR2_X1 U10442 ( .A1(n8954), .A2(n8953), .ZN(n8955) );
  AND4_X1 U10443 ( .A1(n9054), .A2(n8956), .A3(n8955), .A4(n4935), .ZN(n8957)
         );
  NAND2_X1 U10444 ( .A1(n9059), .A2(n8957), .ZN(n8959) );
  OR3_X1 U10445 ( .A1(n9554), .A2(n8959), .A3(n8958), .ZN(n8960) );
  NOR2_X1 U10446 ( .A1(n9535), .A2(n8960), .ZN(n8961) );
  NAND3_X1 U10447 ( .A1(n9495), .A2(n9515), .A3(n8961), .ZN(n8962) );
  NOR2_X1 U10448 ( .A1(n9479), .A2(n8962), .ZN(n8963) );
  NAND4_X1 U10449 ( .A1(n9432), .A2(n9463), .A3(n8963), .A4(n9452), .ZN(n8964)
         );
  NOR4_X1 U10450 ( .A1(n9365), .A2(n9403), .A3(n9425), .A4(n8964), .ZN(n8965)
         );
  OAI22_X1 U10451 ( .A1(n8966), .A2(n5155), .B1(n9124), .B2(n8967), .ZN(n9126)
         );
  INV_X1 U10452 ( .A(n8967), .ZN(n8968) );
  NOR2_X1 U10453 ( .A1(n8968), .A2(n10467), .ZN(n9125) );
  INV_X1 U10454 ( .A(n8969), .ZN(n8973) );
  NOR2_X1 U10455 ( .A1(n9121), .A2(n8970), .ZN(n8972) );
  NAND2_X1 U10456 ( .A1(n5155), .A2(n9565), .ZN(n8971) );
  OR2_X1 U10457 ( .A1(n9131), .A2(n8971), .ZN(n9119) );
  MUX2_X1 U10458 ( .A(n8973), .B(n8972), .S(n9119), .Z(n9123) );
  AND2_X1 U10459 ( .A1(n9393), .A2(n9243), .ZN(n8974) );
  OAI21_X1 U10460 ( .B1(n9365), .B2(n8974), .A(n9119), .ZN(n9104) );
  OR2_X1 U10461 ( .A1(n9403), .A2(n6813), .ZN(n8978) );
  NAND2_X1 U10462 ( .A1(n9381), .A2(n8976), .ZN(n8977) );
  INV_X1 U10463 ( .A(n9119), .ZN(n9111) );
  MUX2_X1 U10464 ( .A(n8978), .B(n8977), .S(n9111), .Z(n9101) );
  AND2_X1 U10465 ( .A1(n8980), .A2(n8979), .ZN(n9086) );
  INV_X1 U10466 ( .A(n9086), .ZN(n8982) );
  OR2_X1 U10467 ( .A1(n8982), .A2(n8981), .ZN(n8984) );
  AND2_X1 U10468 ( .A1(n8984), .A2(n8983), .ZN(n9089) );
  NAND2_X1 U10469 ( .A1(n8997), .A2(n9001), .ZN(n8986) );
  MUX2_X1 U10470 ( .A(n8986), .B(n8985), .S(n9119), .Z(n9004) );
  NAND2_X1 U10471 ( .A1(n9004), .A2(n8987), .ZN(n8992) );
  NAND2_X1 U10472 ( .A1(n8989), .A2(n8988), .ZN(n8991) );
  INV_X1 U10473 ( .A(n9014), .ZN(n8990) );
  AOI21_X1 U10474 ( .B1(n8992), .B2(n8991), .A(n8990), .ZN(n9015) );
  AND2_X1 U10475 ( .A1(n9006), .A2(n5155), .ZN(n8994) );
  OAI211_X1 U10476 ( .C1(n8994), .C2(n8993), .A(n9011), .B(n9007), .ZN(n8995)
         );
  NAND3_X1 U10477 ( .A1(n8995), .A2(n9009), .A3(n9119), .ZN(n9000) );
  AOI21_X1 U10478 ( .B1(n8997), .B2(n8996), .A(n9111), .ZN(n8998) );
  AOI21_X1 U10479 ( .B1(n9000), .B2(n8999), .A(n8998), .ZN(n9005) );
  NAND2_X1 U10480 ( .A1(n9017), .A2(n9001), .ZN(n9002) );
  NAND2_X1 U10481 ( .A1(n9002), .A2(n9119), .ZN(n9003) );
  NAND2_X1 U10482 ( .A1(n9007), .A2(n9006), .ZN(n9010) );
  NAND3_X1 U10483 ( .A1(n9010), .A2(n9009), .A3(n9008), .ZN(n9012) );
  NAND3_X1 U10484 ( .A1(n9012), .A2(n9111), .A3(n9011), .ZN(n9013) );
  MUX2_X1 U10485 ( .A(n9019), .B(n9018), .S(n9119), .Z(n9020) );
  NAND3_X1 U10486 ( .A1(n9022), .A2(n9021), .A3(n9020), .ZN(n9027) );
  NAND2_X1 U10487 ( .A1(n9272), .A2(n9119), .ZN(n9025) );
  NAND2_X1 U10488 ( .A1(n9023), .A2(n9111), .ZN(n9024) );
  MUX2_X1 U10489 ( .A(n9025), .B(n9024), .S(n10505), .Z(n9026) );
  AOI21_X1 U10490 ( .B1(n9031), .B2(n9028), .A(n9111), .ZN(n9030) );
  NAND2_X1 U10491 ( .A1(n9032), .A2(n9033), .ZN(n9029) );
  NAND2_X1 U10492 ( .A1(n9039), .A2(n9031), .ZN(n9036) );
  INV_X1 U10493 ( .A(n9031), .ZN(n9034) );
  OAI211_X1 U10494 ( .C1(n9034), .C2(n9033), .A(n9041), .B(n9032), .ZN(n9035)
         );
  MUX2_X1 U10495 ( .A(n9036), .B(n9035), .S(n9119), .Z(n9037) );
  INV_X1 U10496 ( .A(n9037), .ZN(n9038) );
  NAND2_X1 U10497 ( .A1(n9040), .A2(n9043), .ZN(n9048) );
  NAND2_X1 U10498 ( .A1(n9042), .A2(n9041), .ZN(n9046) );
  INV_X1 U10499 ( .A(n9043), .ZN(n9044) );
  AOI21_X1 U10500 ( .B1(n9046), .B2(n9045), .A(n9044), .ZN(n9047) );
  NOR2_X1 U10501 ( .A1(n10220), .A2(n9119), .ZN(n9051) );
  AND2_X1 U10502 ( .A1(n10220), .A2(n9119), .ZN(n9050) );
  MUX2_X1 U10503 ( .A(n9051), .B(n9050), .S(n9049), .Z(n9052) );
  INV_X1 U10504 ( .A(n9052), .ZN(n9053) );
  MUX2_X1 U10505 ( .A(n9057), .B(n9056), .S(n9119), .Z(n9058) );
  MUX2_X1 U10506 ( .A(n9061), .B(n9060), .S(n9119), .Z(n9062) );
  NAND2_X1 U10507 ( .A1(n9064), .A2(n9063), .ZN(n9070) );
  NOR2_X1 U10508 ( .A1(n9066), .A2(n9065), .ZN(n9067) );
  MUX2_X1 U10509 ( .A(n9067), .B(n4537), .S(n9119), .Z(n9068) );
  NOR2_X1 U10510 ( .A1(n9554), .A2(n9068), .ZN(n9069) );
  NAND2_X1 U10511 ( .A1(n9070), .A2(n9069), .ZN(n9074) );
  AND2_X1 U10512 ( .A1(n9078), .A2(n9071), .ZN(n9072) );
  MUX2_X1 U10513 ( .A(n9527), .B(n9072), .S(n9111), .Z(n9073) );
  NAND2_X1 U10514 ( .A1(n9074), .A2(n9073), .ZN(n9079) );
  AND2_X1 U10515 ( .A1(n9076), .A2(n9075), .ZN(n9082) );
  NAND2_X1 U10516 ( .A1(n9085), .A2(n9080), .ZN(n9081) );
  NAND3_X1 U10517 ( .A1(n9083), .A2(n9086), .A3(n9478), .ZN(n9084) );
  INV_X1 U10518 ( .A(n9085), .ZN(n9087) );
  OAI21_X1 U10519 ( .B1(n9088), .B2(n9087), .A(n9086), .ZN(n9090) );
  NAND3_X1 U10520 ( .A1(n9159), .A2(n9091), .A3(n9119), .ZN(n9093) );
  OR3_X1 U10521 ( .A1(n9159), .A2(n9091), .A3(n9119), .ZN(n9092) );
  NAND2_X1 U10522 ( .A1(n9093), .A2(n9092), .ZN(n9094) );
  NOR2_X1 U10523 ( .A1(n9436), .A2(n9094), .ZN(n9095) );
  MUX2_X1 U10524 ( .A(n9096), .B(n9417), .S(n9119), .Z(n9097) );
  MUX2_X1 U10525 ( .A(n9380), .B(n9381), .S(n9119), .Z(n9098) );
  OAI211_X1 U10526 ( .C1(n9101), .C2(n9100), .A(n9099), .B(n9098), .ZN(n9103)
         );
  AOI21_X1 U10527 ( .B1(n9104), .B2(n9103), .A(n9102), .ZN(n9110) );
  AOI21_X1 U10528 ( .B1(n9106), .B2(n9105), .A(n9119), .ZN(n9109) );
  NAND3_X1 U10529 ( .A1(n9372), .A2(n9145), .A3(n9111), .ZN(n9107) );
  OAI211_X1 U10530 ( .C1(n9110), .C2(n9109), .A(n9108), .B(n9107), .ZN(n9117)
         );
  MUX2_X1 U10531 ( .A(n9113), .B(n9112), .S(n9111), .Z(n9114) );
  INV_X1 U10532 ( .A(n9118), .ZN(n9120) );
  MUX2_X1 U10533 ( .A(n9121), .B(n9120), .S(n4706), .Z(n9122) );
  NOR3_X1 U10534 ( .A1(n9130), .A2(n9129), .A3(n9390), .ZN(n9133) );
  OAI21_X1 U10535 ( .B1(n9134), .B2(n9131), .A(P2_B_REG_SCAN_IN), .ZN(n9132)
         );
  OAI22_X1 U10536 ( .A1(n9135), .A2(n9134), .B1(n9133), .B2(n9132), .ZN(
        P2_U3244) );
  NAND2_X1 U10537 ( .A1(n10422), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n9136) );
  OAI21_X1 U10538 ( .B1(n4497), .B2(n10422), .A(n9136), .ZN(P1_U3520) );
  NOR2_X1 U10539 ( .A1(n9239), .A2(n9137), .ZN(n9140) );
  INV_X1 U10540 ( .A(n9391), .ZN(n9255) );
  NAND3_X1 U10541 ( .A1(n9138), .A2(n9235), .A3(n9255), .ZN(n9139) );
  OAI21_X1 U10542 ( .B1(n9140), .B2(n9240), .A(n9139), .ZN(n9142) );
  NAND2_X1 U10543 ( .A1(n9142), .A2(n9141), .ZN(n9148) );
  INV_X1 U10544 ( .A(n9143), .ZN(n9394) );
  AOI22_X1 U10545 ( .A1(n9255), .A2(n9224), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3152), .ZN(n9144) );
  OAI21_X1 U10546 ( .B1(n9145), .B2(n9218), .A(n9144), .ZN(n9146) );
  AOI21_X1 U10547 ( .B1(n9394), .B2(n9249), .A(n9146), .ZN(n9147) );
  OAI211_X1 U10548 ( .C1(n9656), .C2(n9252), .A(n9148), .B(n9147), .ZN(
        P2_U3216) );
  INV_X1 U10549 ( .A(n9149), .ZN(n9150) );
  NOR2_X1 U10550 ( .A1(n9151), .A2(n9150), .ZN(n9153) );
  NAND3_X1 U10551 ( .A1(n9153), .A2(n9212), .A3(n9152), .ZN(n9162) );
  INV_X1 U10552 ( .A(n9153), .ZN(n9154) );
  NAND3_X1 U10553 ( .A1(n9154), .A2(n9235), .A3(n9258), .ZN(n9161) );
  INV_X1 U10554 ( .A(n9453), .ZN(n9157) );
  OAI22_X1 U10555 ( .A1(n9155), .A2(n9204), .B1(n9181), .B2(n9390), .ZN(n9448)
         );
  AOI22_X1 U10556 ( .A1(n9448), .A2(n9182), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n9156) );
  OAI21_X1 U10557 ( .B1(n9230), .B2(n9157), .A(n9156), .ZN(n9158) );
  AOI21_X1 U10558 ( .B1(n9159), .B2(n10593), .A(n9158), .ZN(n9160) );
  NAND3_X1 U10559 ( .A1(n9162), .A2(n9161), .A3(n9160), .ZN(P2_U3218) );
  OR2_X1 U10560 ( .A1(n9180), .A2(n9204), .ZN(n9165) );
  OR2_X1 U10561 ( .A1(n9163), .A2(n9390), .ZN(n9164) );
  NAND2_X1 U10562 ( .A1(n9165), .A2(n9164), .ZN(n9517) );
  AOI22_X1 U10563 ( .A1(n9182), .A2(n9517), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3152), .ZN(n9166) );
  OAI21_X1 U10564 ( .B1(n9230), .B2(n9513), .A(n9166), .ZN(n9176) );
  NOR3_X1 U10565 ( .A1(n4844), .A2(n9167), .A3(n9240), .ZN(n9174) );
  NAND3_X1 U10566 ( .A1(n9168), .A2(n9235), .A3(n9262), .ZN(n9169) );
  OAI21_X1 U10567 ( .B1(n9170), .B2(n9240), .A(n9169), .ZN(n9173) );
  NAND2_X1 U10568 ( .A1(n8338), .A2(n9171), .ZN(n9172) );
  MUX2_X1 U10569 ( .A(n9174), .B(n9173), .S(n9172), .Z(n9175) );
  AOI211_X1 U10570 ( .C1(n9626), .C2(n10593), .A(n9176), .B(n9175), .ZN(n9177)
         );
  INV_X1 U10571 ( .A(n9177), .ZN(P2_U3221) );
  XNOR2_X1 U10572 ( .A(n9179), .B(n9178), .ZN(n9187) );
  INV_X1 U10573 ( .A(n9487), .ZN(n9184) );
  OAI22_X1 U10574 ( .A1(n9181), .A2(n9204), .B1(n9180), .B2(n9390), .ZN(n9482)
         );
  AOI22_X1 U10575 ( .A1(n9482), .A2(n9182), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3152), .ZN(n9183) );
  OAI21_X1 U10576 ( .B1(n9230), .B2(n9184), .A(n9183), .ZN(n9185) );
  AOI21_X1 U10577 ( .B1(n9486), .B2(n10593), .A(n9185), .ZN(n9186) );
  OAI21_X1 U10578 ( .B1(n9187), .B2(n9240), .A(n9186), .ZN(P2_U3225) );
  XNOR2_X1 U10579 ( .A(n9189), .B(n9188), .ZN(n9190) );
  XNOR2_X1 U10580 ( .A(n9191), .B(n9190), .ZN(n9198) );
  NOR2_X1 U10581 ( .A1(n9230), .A2(n9415), .ZN(n9196) );
  OR2_X1 U10582 ( .A1(n9391), .A2(n9204), .ZN(n9193) );
  NAND2_X1 U10583 ( .A1(n9257), .A2(n9245), .ZN(n9192) );
  AND2_X1 U10584 ( .A1(n9193), .A2(n9192), .ZN(n9421) );
  OAI22_X1 U10585 ( .A1(n9421), .A2(n9247), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9194), .ZN(n9195) );
  AOI211_X1 U10586 ( .C1(n9427), .C2(n10593), .A(n9196), .B(n9195), .ZN(n9197)
         );
  OAI21_X1 U10587 ( .B1(n9198), .B2(n9240), .A(n9197), .ZN(P2_U3227) );
  INV_X1 U10588 ( .A(n9439), .ZN(n9668) );
  NAND2_X1 U10589 ( .A1(n9235), .A2(n9257), .ZN(n9202) );
  OR2_X1 U10590 ( .A1(n9240), .A2(n9199), .ZN(n9201) );
  MUX2_X1 U10591 ( .A(n9202), .B(n9201), .S(n9200), .Z(n9210) );
  INV_X1 U10592 ( .A(n9203), .ZN(n9440) );
  OR2_X1 U10593 ( .A1(n9244), .A2(n9204), .ZN(n9206) );
  NAND2_X1 U10594 ( .A1(n9258), .A2(n9245), .ZN(n9205) );
  AND2_X1 U10595 ( .A1(n9206), .A2(n9205), .ZN(n9433) );
  OAI22_X1 U10596 ( .A1(n9433), .A2(n9247), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9207), .ZN(n9208) );
  AOI21_X1 U10597 ( .B1(n9440), .B2(n9249), .A(n9208), .ZN(n9209) );
  OAI211_X1 U10598 ( .C1(n9668), .C2(n9252), .A(n9210), .B(n9209), .ZN(
        P2_U3231) );
  OAI21_X1 U10599 ( .B1(n9221), .B2(n7415), .A(n9211), .ZN(n9213) );
  NAND2_X1 U10600 ( .A1(n9213), .A2(n9212), .ZN(n9228) );
  INV_X1 U10601 ( .A(n9275), .ZN(n9217) );
  NAND2_X1 U10602 ( .A1(n10593), .A2(n9214), .ZN(n9215) );
  OAI211_X1 U10603 ( .C1(n9218), .C2(n9217), .A(n9216), .B(n9215), .ZN(n9219)
         );
  AOI21_X1 U10604 ( .B1(n9220), .B2(n9249), .A(n9219), .ZN(n9227) );
  NOR3_X1 U10605 ( .A1(n9223), .A2(n9222), .A3(n9221), .ZN(n9225) );
  OAI21_X1 U10606 ( .B1(n9225), .B2(n9224), .A(n9277), .ZN(n9226) );
  NAND3_X1 U10607 ( .A1(n9228), .A2(n9227), .A3(n9226), .ZN(P2_U3232) );
  NOR2_X1 U10608 ( .A1(n9230), .A2(n9469), .ZN(n9233) );
  AOI22_X1 U10609 ( .A1(n9258), .A2(n9386), .B1(n9245), .B2(n9260), .ZN(n9461)
         );
  OAI22_X1 U10610 ( .A1(n9247), .A2(n9461), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9231), .ZN(n9232) );
  AOI211_X1 U10611 ( .C1(n9468), .C2(n10593), .A(n9233), .B(n9232), .ZN(n9238)
         );
  NAND3_X1 U10612 ( .A1(n9236), .A2(n9235), .A3(n9259), .ZN(n9237) );
  OAI211_X1 U10613 ( .C1(n4612), .C2(n9240), .A(n9238), .B(n9237), .ZN(
        P2_U3237) );
  INV_X1 U10614 ( .A(n9243), .ZN(n9254) );
  INV_X1 U10615 ( .A(n9244), .ZN(n9256) );
  AOI22_X1 U10616 ( .A1(n9254), .A2(n9386), .B1(n9245), .B2(n9256), .ZN(n9404)
         );
  OAI22_X1 U10617 ( .A1(n9404), .A2(n9247), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9246), .ZN(n9248) );
  AOI21_X1 U10618 ( .B1(n9408), .B2(n9249), .A(n9248), .ZN(n9250) );
  OAI211_X1 U10619 ( .C1(n9660), .C2(n9252), .A(n9251), .B(n9250), .ZN(
        P2_U3242) );
  MUX2_X1 U10620 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n9253), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U10621 ( .A(n9387), .B(P2_DATAO_REG_28__SCAN_IN), .S(n9280), .Z(
        P2_U3580) );
  MUX2_X1 U10622 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n9254), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U10623 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n9255), .S(P2_U3966), .Z(
        P2_U3578) );
  MUX2_X1 U10624 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n9256), .S(P2_U3966), .Z(
        P2_U3577) );
  MUX2_X1 U10625 ( .A(n9257), .B(P2_DATAO_REG_24__SCAN_IN), .S(n9280), .Z(
        P2_U3576) );
  MUX2_X1 U10626 ( .A(n9258), .B(P2_DATAO_REG_23__SCAN_IN), .S(n9280), .Z(
        P2_U3575) );
  MUX2_X1 U10627 ( .A(n9259), .B(P2_DATAO_REG_22__SCAN_IN), .S(n9280), .Z(
        P2_U3574) );
  MUX2_X1 U10628 ( .A(n9260), .B(P2_DATAO_REG_21__SCAN_IN), .S(n9280), .Z(
        P2_U3573) );
  MUX2_X1 U10629 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n9261), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U10630 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n9262), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U10631 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n9263), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U10632 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n9264), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U10633 ( .A(n9265), .B(P2_DATAO_REG_16__SCAN_IN), .S(n9280), .Z(
        P2_U3568) );
  MUX2_X1 U10634 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n9266), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U10635 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n9267), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U10636 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n9268), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U10637 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n9269), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U10638 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n9270), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U10639 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n9271), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U10640 ( .A(n9272), .B(P2_DATAO_REG_8__SCAN_IN), .S(n9280), .Z(
        P2_U3560) );
  MUX2_X1 U10641 ( .A(n9273), .B(P2_DATAO_REG_7__SCAN_IN), .S(n9280), .Z(
        P2_U3559) );
  MUX2_X1 U10642 ( .A(n9274), .B(P2_DATAO_REG_6__SCAN_IN), .S(n9280), .Z(
        P2_U3558) );
  MUX2_X1 U10643 ( .A(n9275), .B(P2_DATAO_REG_5__SCAN_IN), .S(n9280), .Z(
        P2_U3557) );
  MUX2_X1 U10644 ( .A(n9276), .B(P2_DATAO_REG_4__SCAN_IN), .S(n9280), .Z(
        P2_U3556) );
  MUX2_X1 U10645 ( .A(n9277), .B(P2_DATAO_REG_3__SCAN_IN), .S(n9280), .Z(
        P2_U3555) );
  MUX2_X1 U10646 ( .A(n9278), .B(P2_DATAO_REG_2__SCAN_IN), .S(n9280), .Z(
        P2_U3554) );
  MUX2_X1 U10647 ( .A(n9279), .B(P2_DATAO_REG_1__SCAN_IN), .S(n9280), .Z(
        P2_U3553) );
  MUX2_X1 U10648 ( .A(n9281), .B(P2_DATAO_REG_0__SCAN_IN), .S(n9280), .Z(
        P2_U3552) );
  OAI21_X1 U10649 ( .B1(n9284), .B2(n9283), .A(n9282), .ZN(n9285) );
  NAND2_X1 U10650 ( .A1(n10440), .A2(n9285), .ZN(n9294) );
  AND2_X1 U10651 ( .A1(P2_U3152), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n9286) );
  AOI21_X1 U10652 ( .B1(n10441), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n9286), .ZN(
        n9293) );
  NAND2_X1 U10653 ( .A1(n10165), .A2(n9287), .ZN(n9292) );
  OAI211_X1 U10654 ( .C1(n9290), .C2(n9289), .A(n10439), .B(n9288), .ZN(n9291)
         );
  NAND4_X1 U10655 ( .A1(n9294), .A2(n9293), .A3(n9292), .A4(n9291), .ZN(
        P2_U3256) );
  AND2_X1 U10656 ( .A1(P2_U3152), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9302) );
  NAND2_X1 U10657 ( .A1(n9313), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n9316) );
  INV_X1 U10658 ( .A(n9304), .ZN(n9296) );
  INV_X1 U10659 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n10234) );
  NAND2_X1 U10660 ( .A1(n9311), .A2(n10234), .ZN(n9297) );
  NOR2_X1 U10661 ( .A1(n9311), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n9298) );
  AOI211_X1 U10662 ( .C1(n9311), .C2(P2_REG1_REG_17__SCAN_IN), .A(n9299), .B(
        n9298), .ZN(n9300) );
  NOR3_X1 U10663 ( .A1(n10444), .A2(n9315), .A3(n9300), .ZN(n9301) );
  AOI211_X1 U10664 ( .C1(P2_ADDR_REG_17__SCAN_IN), .C2(n10441), .A(n9302), .B(
        n9301), .ZN(n9310) );
  XNOR2_X1 U10665 ( .A(n9313), .B(P2_REG2_REG_17__SCAN_IN), .ZN(n9306) );
  INV_X1 U10666 ( .A(n9306), .ZN(n9308) );
  AOI21_X1 U10667 ( .B1(n9304), .B2(P2_REG2_REG_16__SCAN_IN), .A(n9303), .ZN(
        n9305) );
  INV_X1 U10668 ( .A(n9305), .ZN(n9307) );
  OAI211_X1 U10669 ( .C1(n9308), .C2(n9307), .A(n10440), .B(n9312), .ZN(n9309)
         );
  OAI211_X1 U10670 ( .C1(n10443), .C2(n9311), .A(n9310), .B(n9309), .ZN(
        P2_U3262) );
  NOR2_X1 U10671 ( .A1(n9539), .A2(n9314), .ZN(n9328) );
  AOI211_X1 U10672 ( .C1(n9314), .C2(n9539), .A(n9328), .B(n10442), .ZN(n9326)
         );
  NAND2_X1 U10673 ( .A1(n9317), .A2(n9316), .ZN(n9319) );
  AOI22_X1 U10674 ( .A1(n9320), .A2(n9634), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n9332), .ZN(n9318) );
  NOR2_X1 U10675 ( .A1(n9319), .A2(n9318), .ZN(n9331) );
  AOI21_X1 U10676 ( .B1(n9319), .B2(n9318), .A(n9331), .ZN(n9324) );
  NAND2_X1 U10677 ( .A1(n10165), .A2(n9320), .ZN(n9323) );
  AOI21_X1 U10678 ( .B1(n10441), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n9321), .ZN(
        n9322) );
  OAI211_X1 U10679 ( .C1(n9324), .C2(n10444), .A(n9323), .B(n9322), .ZN(n9325)
         );
  OR2_X1 U10680 ( .A1(n9326), .A2(n9325), .ZN(P2_U3263) );
  NOR2_X1 U10681 ( .A1(n9327), .A2(n9332), .ZN(n9329) );
  NOR2_X1 U10682 ( .A1(n9329), .A2(n9328), .ZN(n9330) );
  XNOR2_X1 U10683 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n9330), .ZN(n9337) );
  INV_X1 U10684 ( .A(n9337), .ZN(n9335) );
  AOI21_X1 U10685 ( .B1(n9332), .B2(n9634), .A(n9331), .ZN(n9333) );
  XNOR2_X1 U10686 ( .A(n9334), .B(n9333), .ZN(n9336) );
  NAND2_X1 U10687 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3152), .ZN(n9338) );
  XNOR2_X1 U10688 ( .A(n9346), .B(n9340), .ZN(n9341) );
  NAND2_X1 U10689 ( .A1(n9570), .A2(n9504), .ZN(n9345) );
  AND2_X1 U10690 ( .A1(n9343), .A2(n9342), .ZN(n9569) );
  INV_X1 U10691 ( .A(n9569), .ZN(n9573) );
  NOR2_X1 U10692 ( .A1(n4499), .A2(n9573), .ZN(n9349) );
  AOI21_X1 U10693 ( .B1(n4499), .B2(P2_REG2_REG_31__SCAN_IN), .A(n9349), .ZN(
        n9344) );
  OAI211_X1 U10694 ( .C1(n9644), .C2(n9552), .A(n9345), .B(n9344), .ZN(
        P2_U3265) );
  OAI211_X1 U10695 ( .C1(n9648), .C2(n9347), .A(n9541), .B(n9346), .ZN(n9574)
         );
  NOR2_X1 U10696 ( .A1(n9648), .A2(n9552), .ZN(n9348) );
  AOI211_X1 U10697 ( .C1(n4499), .C2(P2_REG2_REG_30__SCAN_IN), .A(n9349), .B(
        n9348), .ZN(n9350) );
  OAI21_X1 U10698 ( .B1(n10224), .B2(n9574), .A(n9350), .ZN(P2_U3266) );
  INV_X1 U10699 ( .A(n9351), .ZN(n9360) );
  NAND2_X1 U10700 ( .A1(n9352), .A2(n9504), .ZN(n9356) );
  INV_X1 U10701 ( .A(n9353), .ZN(n9354) );
  AOI22_X1 U10702 ( .A1(P2_REG2_REG_29__SCAN_IN), .A2(n4499), .B1(n9354), .B2(
        n10218), .ZN(n9355) );
  OAI211_X1 U10703 ( .C1(n4793), .C2(n9552), .A(n9356), .B(n9355), .ZN(n9357)
         );
  AOI21_X1 U10704 ( .B1(n9358), .B2(n9540), .A(n9357), .ZN(n9359) );
  OAI21_X1 U10705 ( .B1(n9360), .B2(n9536), .A(n9359), .ZN(P2_U3267) );
  XNOR2_X1 U10706 ( .A(n9361), .B(n9365), .ZN(n9363) );
  OAI21_X1 U10707 ( .B1(n9366), .B2(n9365), .A(n9364), .ZN(n9580) );
  NAND2_X1 U10708 ( .A1(n9580), .A2(n9465), .ZN(n9374) );
  INV_X1 U10709 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n9368) );
  OAI22_X1 U10710 ( .A1(n9540), .A2(n9368), .B1(n9537), .B2(n9367), .ZN(n9371)
         );
  OAI211_X1 U10711 ( .C1(n9652), .C2(n4516), .A(n9541), .B(n9369), .ZN(n9577)
         );
  NOR2_X1 U10712 ( .A1(n9577), .A2(n10224), .ZN(n9370) );
  AOI211_X1 U10713 ( .C1(n10221), .C2(n9372), .A(n9371), .B(n9370), .ZN(n9373)
         );
  OAI211_X1 U10714 ( .C1(n9578), .C2(n4499), .A(n9374), .B(n9373), .ZN(
        P2_U3268) );
  OAI21_X1 U10715 ( .B1(n9376), .B2(n9382), .A(n9375), .ZN(n9585) );
  INV_X1 U10716 ( .A(n9585), .ZN(n9399) );
  AND2_X1 U10717 ( .A1(n9378), .A2(n9377), .ZN(n9385) );
  NAND2_X1 U10718 ( .A1(n9379), .A2(n9380), .ZN(n9383) );
  NAND3_X1 U10719 ( .A1(n9383), .A2(n9382), .A3(n9381), .ZN(n9384) );
  NAND3_X1 U10720 ( .A1(n9385), .A2(n9532), .A3(n9384), .ZN(n9389) );
  NAND2_X1 U10721 ( .A1(n9387), .A2(n9386), .ZN(n9388) );
  OAI211_X1 U10722 ( .C1(n9391), .C2(n9390), .A(n9389), .B(n9388), .ZN(n9583)
         );
  INV_X1 U10723 ( .A(n9407), .ZN(n9392) );
  AOI211_X1 U10724 ( .C1(n9393), .C2(n9392), .A(n10520), .B(n4516), .ZN(n9584)
         );
  NAND2_X1 U10725 ( .A1(n9584), .A2(n9504), .ZN(n9396) );
  AOI22_X1 U10726 ( .A1(P2_REG2_REG_27__SCAN_IN), .A2(n4499), .B1(n9394), .B2(
        n10218), .ZN(n9395) );
  OAI211_X1 U10727 ( .C1(n9656), .C2(n9552), .A(n9396), .B(n9395), .ZN(n9397)
         );
  AOI21_X1 U10728 ( .B1(n9583), .B2(n9540), .A(n9397), .ZN(n9398) );
  OAI21_X1 U10729 ( .B1(n9399), .B2(n9536), .A(n9398), .ZN(P2_U3269) );
  OAI21_X1 U10730 ( .B1(n9401), .B2(n9403), .A(n9400), .ZN(n9591) );
  INV_X1 U10731 ( .A(n9591), .ZN(n9413) );
  AOI22_X1 U10732 ( .A1(n9402), .A2(n10221), .B1(n4499), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n9412) );
  XOR2_X1 U10733 ( .A(n9403), .B(n9379), .Z(n9405) );
  NOR2_X1 U10734 ( .A1(n9660), .A2(n9414), .ZN(n9406) );
  INV_X1 U10735 ( .A(n9408), .ZN(n9409) );
  OAI22_X1 U10736 ( .A1(n9588), .A2(n9565), .B1(n9537), .B2(n9409), .ZN(n9410)
         );
  OAI21_X1 U10737 ( .B1(n9589), .B2(n9410), .A(n9540), .ZN(n9411) );
  OAI211_X1 U10738 ( .C1(n9413), .C2(n9536), .A(n9412), .B(n9411), .ZN(
        P2_U3270) );
  AOI211_X1 U10739 ( .C1(n9427), .C2(n9438), .A(n10520), .B(n9414), .ZN(n9595)
         );
  NOR2_X1 U10740 ( .A1(n9537), .A2(n9415), .ZN(n9423) );
  NAND2_X1 U10741 ( .A1(n9416), .A2(n9432), .ZN(n9431) );
  NAND2_X1 U10742 ( .A1(n9431), .A2(n9417), .ZN(n9420) );
  NAND2_X1 U10743 ( .A1(n9420), .A2(n9419), .ZN(n9418) );
  OAI211_X1 U10744 ( .C1(n9420), .C2(n9419), .A(n9418), .B(n9532), .ZN(n9422)
         );
  NAND2_X1 U10745 ( .A1(n9422), .A2(n9421), .ZN(n9594) );
  AOI211_X1 U10746 ( .C1(n9595), .C2(n9522), .A(n9423), .B(n9594), .ZN(n9430)
         );
  OAI21_X1 U10747 ( .B1(n9426), .B2(n9425), .A(n9424), .ZN(n9596) );
  NAND2_X1 U10748 ( .A1(n9596), .A2(n9465), .ZN(n9429) );
  AOI22_X1 U10749 ( .A1(n9427), .A2(n10221), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n4499), .ZN(n9428) );
  OAI211_X1 U10750 ( .C1(n4499), .C2(n9430), .A(n9429), .B(n9428), .ZN(
        P2_U3271) );
  OAI211_X1 U10751 ( .C1(n9416), .C2(n9432), .A(n9431), .B(n9532), .ZN(n9434)
         );
  NAND2_X1 U10752 ( .A1(n9434), .A2(n9433), .ZN(n9599) );
  INV_X1 U10753 ( .A(n9599), .ZN(n9445) );
  OAI21_X1 U10754 ( .B1(n9437), .B2(n9436), .A(n9435), .ZN(n9601) );
  NAND2_X1 U10755 ( .A1(n9601), .A2(n9465), .ZN(n9444) );
  AOI211_X1 U10756 ( .C1(n9439), .C2(n4512), .A(n10520), .B(n4786), .ZN(n9600)
         );
  AOI22_X1 U10757 ( .A1(n4499), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n9440), .B2(
        n10218), .ZN(n9441) );
  OAI21_X1 U10758 ( .B1(n9668), .B2(n9552), .A(n9441), .ZN(n9442) );
  AOI21_X1 U10759 ( .B1(n9600), .B2(n9504), .A(n9442), .ZN(n9443) );
  OAI211_X1 U10760 ( .C1(n4499), .C2(n9445), .A(n9444), .B(n9443), .ZN(
        P2_U3272) );
  XNOR2_X1 U10761 ( .A(n9447), .B(n9446), .ZN(n9449) );
  AOI21_X1 U10762 ( .B1(n9449), .B2(n9532), .A(n9448), .ZN(n9605) );
  AOI21_X1 U10763 ( .B1(n9452), .B2(n9451), .A(n9450), .ZN(n9607) );
  NAND2_X1 U10764 ( .A1(n9607), .A2(n9465), .ZN(n9458) );
  OAI211_X1 U10765 ( .C1(n9466), .C2(n9672), .A(n9541), .B(n4512), .ZN(n9604)
         );
  INV_X1 U10766 ( .A(n9604), .ZN(n9456) );
  AOI22_X1 U10767 ( .A1(n4499), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n9453), .B2(
        n10218), .ZN(n9454) );
  OAI21_X1 U10768 ( .B1(n9672), .B2(n9552), .A(n9454), .ZN(n9455) );
  AOI21_X1 U10769 ( .B1(n9456), .B2(n9504), .A(n9455), .ZN(n9457) );
  OAI211_X1 U10770 ( .C1(n4499), .C2(n9605), .A(n9458), .B(n9457), .ZN(
        P2_U3273) );
  OAI211_X1 U10771 ( .C1(n9460), .C2(n9463), .A(n9459), .B(n9532), .ZN(n9462)
         );
  NAND2_X1 U10772 ( .A1(n9462), .A2(n9461), .ZN(n9610) );
  INV_X1 U10773 ( .A(n9610), .ZN(n9475) );
  XNOR2_X1 U10774 ( .A(n9464), .B(n9463), .ZN(n9612) );
  NAND2_X1 U10775 ( .A1(n9612), .A2(n9465), .ZN(n9474) );
  INV_X1 U10776 ( .A(n9485), .ZN(n9467) );
  AOI211_X1 U10777 ( .C1(n9468), .C2(n9467), .A(n10520), .B(n9466), .ZN(n9611)
         );
  NOR2_X1 U10778 ( .A1(n9676), .A2(n9552), .ZN(n9472) );
  OAI22_X1 U10779 ( .A1(n9540), .A2(n9470), .B1(n9469), .B2(n9537), .ZN(n9471)
         );
  AOI211_X1 U10780 ( .C1(n9611), .C2(n9504), .A(n9472), .B(n9471), .ZN(n9473)
         );
  OAI211_X1 U10781 ( .C1(n4499), .C2(n9475), .A(n9474), .B(n9473), .ZN(
        P2_U3274) );
  XNOR2_X1 U10782 ( .A(n9476), .B(n9479), .ZN(n9617) );
  INV_X1 U10783 ( .A(n9617), .ZN(n9492) );
  NAND2_X1 U10784 ( .A1(n9477), .A2(n9478), .ZN(n9480) );
  XNOR2_X1 U10785 ( .A(n9480), .B(n9479), .ZN(n9481) );
  NAND2_X1 U10786 ( .A1(n9481), .A2(n9532), .ZN(n9484) );
  INV_X1 U10787 ( .A(n9482), .ZN(n9483) );
  NAND2_X1 U10788 ( .A1(n9484), .A2(n9483), .ZN(n9615) );
  AOI211_X1 U10789 ( .C1(n9486), .C2(n9501), .A(n10520), .B(n9485), .ZN(n9616)
         );
  NAND2_X1 U10790 ( .A1(n9616), .A2(n9504), .ZN(n9489) );
  AOI22_X1 U10791 ( .A1(n4499), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n9487), .B2(
        n10218), .ZN(n9488) );
  OAI211_X1 U10792 ( .C1(n9680), .C2(n9552), .A(n9489), .B(n9488), .ZN(n9490)
         );
  AOI21_X1 U10793 ( .B1(n9615), .B2(n9540), .A(n9490), .ZN(n9491) );
  OAI21_X1 U10794 ( .B1(n9492), .B2(n9536), .A(n9491), .ZN(P2_U3275) );
  AOI21_X1 U10795 ( .B1(n9495), .B2(n9494), .A(n9493), .ZN(n9622) );
  INV_X1 U10796 ( .A(n9622), .ZN(n9511) );
  NAND2_X1 U10797 ( .A1(n9496), .A2(n9497), .ZN(n9498) );
  NAND3_X1 U10798 ( .A1(n9477), .A2(n9532), .A3(n9498), .ZN(n9500) );
  NAND2_X1 U10799 ( .A1(n9500), .A2(n9499), .ZN(n9620) );
  INV_X1 U10800 ( .A(n9503), .ZN(n9684) );
  INV_X1 U10801 ( .A(n9501), .ZN(n9502) );
  AOI211_X1 U10802 ( .C1(n9503), .C2(n9520), .A(n10520), .B(n9502), .ZN(n9621)
         );
  NAND2_X1 U10803 ( .A1(n9621), .A2(n9504), .ZN(n9508) );
  INV_X1 U10804 ( .A(n9505), .ZN(n9506) );
  AOI22_X1 U10805 ( .A1(n4499), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9506), .B2(
        n10218), .ZN(n9507) );
  OAI211_X1 U10806 ( .C1(n9684), .C2(n9552), .A(n9508), .B(n9507), .ZN(n9509)
         );
  AOI21_X1 U10807 ( .B1(n9620), .B2(n9540), .A(n9509), .ZN(n9510) );
  OAI21_X1 U10808 ( .B1(n9511), .B2(n9536), .A(n9510), .ZN(P2_U3276) );
  XNOR2_X1 U10809 ( .A(n9512), .B(n9515), .ZN(n9629) );
  OAI22_X1 U10810 ( .A1(n9540), .A2(n9514), .B1(n9513), .B2(n9537), .ZN(n9525)
         );
  XNOR2_X1 U10811 ( .A(n9516), .B(n9515), .ZN(n9518) );
  AOI21_X1 U10812 ( .B1(n9518), .B2(n9532), .A(n9517), .ZN(n9628) );
  INV_X1 U10813 ( .A(n9520), .ZN(n9521) );
  AOI211_X1 U10814 ( .C1(n9626), .C2(n9519), .A(n10520), .B(n9521), .ZN(n9625)
         );
  NAND2_X1 U10815 ( .A1(n9625), .A2(n9522), .ZN(n9523) );
  AOI21_X1 U10816 ( .B1(n9628), .B2(n9523), .A(n4499), .ZN(n9524) );
  AOI211_X1 U10817 ( .C1(n10221), .C2(n9626), .A(n9525), .B(n9524), .ZN(n9526)
         );
  OAI21_X1 U10818 ( .B1(n9629), .B2(n9536), .A(n9526), .ZN(P2_U3277) );
  NAND2_X1 U10819 ( .A1(n9557), .A2(n9527), .ZN(n9528) );
  NAND2_X1 U10820 ( .A1(n9528), .A2(n9535), .ZN(n9530) );
  NAND2_X1 U10821 ( .A1(n9530), .A2(n9529), .ZN(n9533) );
  AOI21_X1 U10822 ( .B1(n9533), .B2(n9532), .A(n9531), .ZN(n9631) );
  XOR2_X1 U10823 ( .A(n9535), .B(n9534), .Z(n9632) );
  OR2_X1 U10824 ( .A1(n9632), .A2(n9536), .ZN(n9547) );
  OAI22_X1 U10825 ( .A1(n9540), .A2(n9539), .B1(n9538), .B2(n9537), .ZN(n9544)
         );
  OAI211_X1 U10826 ( .C1(n9542), .C2(n9689), .A(n9519), .B(n9541), .ZN(n9630)
         );
  NOR2_X1 U10827 ( .A1(n9630), .A2(n10224), .ZN(n9543) );
  AOI211_X1 U10828 ( .C1(n10221), .C2(n9545), .A(n9544), .B(n9543), .ZN(n9546)
         );
  OAI211_X1 U10829 ( .C1(n4499), .C2(n9631), .A(n9547), .B(n9546), .ZN(
        P2_U3278) );
  OAI21_X1 U10830 ( .B1(n4558), .B2(n9554), .A(n9548), .ZN(n10233) );
  INV_X1 U10831 ( .A(n9549), .ZN(n9550) );
  AOI22_X1 U10832 ( .A1(n4499), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n9550), .B2(
        n10218), .ZN(n9551) );
  OAI21_X1 U10833 ( .B1(n4940), .B2(n9552), .A(n9551), .ZN(n9567) );
  AOI21_X1 U10834 ( .B1(n9555), .B2(n9554), .A(n9553), .ZN(n9558) );
  AOI21_X1 U10835 ( .B1(n9558), .B2(n9557), .A(n9556), .ZN(n9564) );
  XNOR2_X1 U10836 ( .A(n9560), .B(n9559), .ZN(n9561) );
  OAI21_X1 U10837 ( .B1(n10520), .B2(n9561), .A(n9564), .ZN(n10231) );
  AOI21_X1 U10838 ( .B1(n10233), .B2(n9562), .A(n10231), .ZN(n9563) );
  AOI211_X1 U10839 ( .C1(n9565), .C2(n9564), .A(n4499), .B(n9563), .ZN(n9566)
         );
  AOI211_X1 U10840 ( .C1(n10227), .C2(n10233), .A(n9567), .B(n9566), .ZN(n9568) );
  INV_X1 U10841 ( .A(n9568), .ZN(P2_U3279) );
  NOR2_X1 U10842 ( .A1(n9570), .A2(n9569), .ZN(n9641) );
  MUX2_X1 U10843 ( .A(n9571), .B(n9641), .S(n10541), .Z(n9572) );
  OAI21_X1 U10844 ( .B1(n9644), .B2(n9640), .A(n9572), .ZN(P2_U3551) );
  NAND2_X1 U10845 ( .A1(n9574), .A2(n9573), .ZN(n9645) );
  MUX2_X1 U10846 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9645), .S(n10541), .Z(
        n9575) );
  INV_X1 U10847 ( .A(n9575), .ZN(n9576) );
  OAI21_X1 U10848 ( .B1(n9648), .B2(n9640), .A(n9576), .ZN(P2_U3550) );
  INV_X1 U10849 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9581) );
  NAND2_X1 U10850 ( .A1(n9578), .A2(n9577), .ZN(n9579) );
  AOI21_X1 U10851 ( .B1(n9580), .B2(n10524), .A(n9579), .ZN(n9649) );
  MUX2_X1 U10852 ( .A(n9581), .B(n9649), .S(n10541), .Z(n9582) );
  OAI21_X1 U10853 ( .B1(n9652), .B2(n9640), .A(n9582), .ZN(P2_U3548) );
  INV_X1 U10854 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9586) );
  AOI211_X1 U10855 ( .C1(n9585), .C2(n10524), .A(n9584), .B(n9583), .ZN(n9653)
         );
  MUX2_X1 U10856 ( .A(n9586), .B(n9653), .S(n10541), .Z(n9587) );
  OAI21_X1 U10857 ( .B1(n9656), .B2(n9640), .A(n9587), .ZN(P2_U3547) );
  INV_X1 U10858 ( .A(n9588), .ZN(n9590) );
  MUX2_X1 U10859 ( .A(n9592), .B(n9657), .S(n10541), .Z(n9593) );
  OAI21_X1 U10860 ( .B1(n9660), .B2(n9640), .A(n9593), .ZN(P2_U3546) );
  INV_X1 U10861 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9597) );
  AOI211_X1 U10862 ( .C1(n9596), .C2(n10524), .A(n9595), .B(n9594), .ZN(n9661)
         );
  MUX2_X1 U10863 ( .A(n9597), .B(n9661), .S(n10541), .Z(n9598) );
  OAI21_X1 U10864 ( .B1(n9664), .B2(n9640), .A(n9598), .ZN(P2_U3545) );
  INV_X1 U10865 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9602) );
  AOI211_X1 U10866 ( .C1(n9601), .C2(n10524), .A(n9600), .B(n9599), .ZN(n9665)
         );
  MUX2_X1 U10867 ( .A(n9602), .B(n9665), .S(n10541), .Z(n9603) );
  OAI21_X1 U10868 ( .B1(n9668), .B2(n9640), .A(n9603), .ZN(P2_U3544) );
  NAND2_X1 U10869 ( .A1(n9605), .A2(n9604), .ZN(n9606) );
  AOI21_X1 U10870 ( .B1(n9607), .B2(n10524), .A(n9606), .ZN(n9669) );
  MUX2_X1 U10871 ( .A(n9608), .B(n9669), .S(n10541), .Z(n9609) );
  OAI21_X1 U10872 ( .B1(n9672), .B2(n9640), .A(n9609), .ZN(P2_U3543) );
  INV_X1 U10873 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9613) );
  AOI211_X1 U10874 ( .C1(n9612), .C2(n10524), .A(n9611), .B(n9610), .ZN(n9673)
         );
  MUX2_X1 U10875 ( .A(n9613), .B(n9673), .S(n10541), .Z(n9614) );
  OAI21_X1 U10876 ( .B1(n9676), .B2(n9640), .A(n9614), .ZN(P2_U3542) );
  INV_X1 U10877 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9618) );
  AOI211_X1 U10878 ( .C1(n9617), .C2(n10524), .A(n9616), .B(n9615), .ZN(n9677)
         );
  MUX2_X1 U10879 ( .A(n9618), .B(n9677), .S(n10541), .Z(n9619) );
  OAI21_X1 U10880 ( .B1(n9680), .B2(n9640), .A(n9619), .ZN(P2_U3541) );
  AOI211_X1 U10881 ( .C1(n9622), .C2(n10524), .A(n9621), .B(n9620), .ZN(n9681)
         );
  MUX2_X1 U10882 ( .A(n9623), .B(n9681), .S(n10541), .Z(n9624) );
  OAI21_X1 U10883 ( .B1(n9684), .B2(n9640), .A(n9624), .ZN(P2_U3540) );
  AOI21_X1 U10884 ( .B1(n10475), .B2(n9626), .A(n9625), .ZN(n9627) );
  OAI211_X1 U10885 ( .C1(n9629), .C2(n10478), .A(n9628), .B(n9627), .ZN(n9685)
         );
  MUX2_X1 U10886 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9685), .S(n10541), .Z(
        P2_U3539) );
  OAI211_X1 U10887 ( .C1(n9632), .C2(n10478), .A(n9631), .B(n9630), .ZN(n9633)
         );
  INV_X1 U10888 ( .A(n9633), .ZN(n9686) );
  MUX2_X1 U10889 ( .A(n9634), .B(n9686), .S(n10541), .Z(n9635) );
  OAI21_X1 U10890 ( .B1(n9689), .B2(n9640), .A(n9635), .ZN(P2_U3538) );
  AOI211_X1 U10891 ( .C1(n9638), .C2(n10524), .A(n9637), .B(n9636), .ZN(n9690)
         );
  MUX2_X1 U10892 ( .A(n8383), .B(n9690), .S(n10541), .Z(n9639) );
  OAI21_X1 U10893 ( .B1(n9693), .B2(n9640), .A(n9639), .ZN(P2_U3536) );
  MUX2_X1 U10894 ( .A(n9642), .B(n9641), .S(n10528), .Z(n9643) );
  OAI21_X1 U10895 ( .B1(n9644), .B2(n9692), .A(n9643), .ZN(P2_U3519) );
  MUX2_X1 U10896 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n9645), .S(n10528), .Z(
        n9646) );
  INV_X1 U10897 ( .A(n9646), .ZN(n9647) );
  OAI21_X1 U10898 ( .B1(n9648), .B2(n9692), .A(n9647), .ZN(P2_U3518) );
  MUX2_X1 U10899 ( .A(n9650), .B(n9649), .S(n10528), .Z(n9651) );
  OAI21_X1 U10900 ( .B1(n9652), .B2(n9692), .A(n9651), .ZN(P2_U3516) );
  MUX2_X1 U10901 ( .A(n9654), .B(n9653), .S(n10528), .Z(n9655) );
  OAI21_X1 U10902 ( .B1(n9656), .B2(n9692), .A(n9655), .ZN(P2_U3515) );
  INV_X1 U10903 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9658) );
  MUX2_X1 U10904 ( .A(n9658), .B(n9657), .S(n10528), .Z(n9659) );
  OAI21_X1 U10905 ( .B1(n9660), .B2(n9692), .A(n9659), .ZN(P2_U3514) );
  INV_X1 U10906 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9662) );
  MUX2_X1 U10907 ( .A(n9662), .B(n9661), .S(n10528), .Z(n9663) );
  OAI21_X1 U10908 ( .B1(n9664), .B2(n9692), .A(n9663), .ZN(P2_U3513) );
  MUX2_X1 U10909 ( .A(n9666), .B(n9665), .S(n10528), .Z(n9667) );
  OAI21_X1 U10910 ( .B1(n9668), .B2(n9692), .A(n9667), .ZN(P2_U3512) );
  INV_X1 U10911 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9670) );
  MUX2_X1 U10912 ( .A(n9670), .B(n9669), .S(n10528), .Z(n9671) );
  OAI21_X1 U10913 ( .B1(n9672), .B2(n9692), .A(n9671), .ZN(P2_U3511) );
  MUX2_X1 U10914 ( .A(n9674), .B(n9673), .S(n10528), .Z(n9675) );
  OAI21_X1 U10915 ( .B1(n9676), .B2(n9692), .A(n9675), .ZN(P2_U3510) );
  MUX2_X1 U10916 ( .A(n9678), .B(n9677), .S(n10528), .Z(n9679) );
  OAI21_X1 U10917 ( .B1(n9680), .B2(n9692), .A(n9679), .ZN(P2_U3509) );
  MUX2_X1 U10918 ( .A(n9682), .B(n9681), .S(n10528), .Z(n9683) );
  OAI21_X1 U10919 ( .B1(n9684), .B2(n9692), .A(n9683), .ZN(P2_U3508) );
  MUX2_X1 U10920 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9685), .S(n10528), .Z(
        P2_U3507) );
  INV_X1 U10921 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9687) );
  MUX2_X1 U10922 ( .A(n9687), .B(n9686), .S(n10528), .Z(n9688) );
  OAI21_X1 U10923 ( .B1(n9689), .B2(n9692), .A(n9688), .ZN(P2_U3505) );
  MUX2_X1 U10924 ( .A(n5502), .B(n9690), .S(n10528), .Z(n9691) );
  OAI21_X1 U10925 ( .B1(n9693), .B2(n9692), .A(n9691), .ZN(P2_U3499) );
  INV_X1 U10926 ( .A(n9694), .ZN(n10158) );
  NOR4_X1 U10927 ( .A1(n9695), .A2(P2_IR_REG_30__SCAN_IN), .A3(n9696), .A4(
        P2_U3152), .ZN(n9697) );
  AOI21_X1 U10928 ( .B1(n9698), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9697), .ZN(
        n9699) );
  OAI21_X1 U10929 ( .B1(n10158), .B2(n8904), .A(n9699), .ZN(P2_U3327) );
  MUX2_X1 U10930 ( .A(n9700), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  INV_X1 U10931 ( .A(n9754), .ZN(n9704) );
  OAI21_X1 U10932 ( .B1(n9702), .B2(n9753), .A(n9701), .ZN(n9703) );
  OAI21_X1 U10933 ( .B1(n9704), .B2(n9753), .A(n9703), .ZN(n9705) );
  NAND2_X1 U10934 ( .A1(n9705), .A2(n9802), .ZN(n9709) );
  AOI22_X1 U10935 ( .A1(n9768), .A2(n10007), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9706) );
  OAI21_X1 U10936 ( .B1(n9728), .B2(n9804), .A(n9706), .ZN(n9707) );
  AOI21_X1 U10937 ( .B1(n10001), .B2(n9809), .A(n9707), .ZN(n9708) );
  OAI211_X1 U10938 ( .C1(n10003), .C2(n9812), .A(n9709), .B(n9708), .ZN(
        P1_U3214) );
  INV_X1 U10939 ( .A(n9710), .ZN(n9713) );
  INV_X1 U10940 ( .A(n9782), .ZN(n9712) );
  NOR3_X1 U10941 ( .A1(n9713), .A2(n9712), .A3(n9711), .ZN(n9715) );
  INV_X1 U10942 ( .A(n9714), .ZN(n9764) );
  OAI21_X1 U10943 ( .B1(n9715), .B2(n9764), .A(n9802), .ZN(n9721) );
  NAND2_X1 U10944 ( .A1(n9786), .A2(n9815), .ZN(n9716) );
  NAND2_X1 U10945 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9903) );
  OAI211_X1 U10946 ( .C1(n9717), .C2(n9806), .A(n9716), .B(n9903), .ZN(n9718)
         );
  AOI21_X1 U10947 ( .B1(n9719), .B2(n9809), .A(n9718), .ZN(n9720) );
  OAI211_X1 U10948 ( .C1(n9722), .C2(n9812), .A(n9721), .B(n9720), .ZN(
        P1_U3217) );
  OAI21_X1 U10949 ( .B1(n9725), .B2(n9724), .A(n9723), .ZN(n9726) );
  NAND2_X1 U10950 ( .A1(n9726), .A2(n9802), .ZN(n9731) );
  AOI22_X1 U10951 ( .A1(n9786), .A2(n10036), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9727) );
  OAI21_X1 U10952 ( .B1(n9728), .B2(n9806), .A(n9727), .ZN(n9729) );
  AOI21_X1 U10953 ( .B1(n10030), .B2(n9809), .A(n9729), .ZN(n9730) );
  OAI211_X1 U10954 ( .C1(n10032), .C2(n9812), .A(n9731), .B(n9730), .ZN(
        P1_U3221) );
  AOI21_X1 U10955 ( .B1(n9734), .B2(n9733), .A(n9800), .ZN(n9739) );
  AOI22_X1 U10956 ( .A1(n9768), .A2(n9814), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n9736) );
  NAND2_X1 U10957 ( .A1(n9809), .A2(n9977), .ZN(n9735) );
  OAI211_X1 U10958 ( .C1(n9973), .C2(n9804), .A(n9736), .B(n9735), .ZN(n9737)
         );
  AOI21_X1 U10959 ( .B1(n10079), .B2(n9792), .A(n9737), .ZN(n9738) );
  OAI21_X1 U10960 ( .B1(n9739), .B2(n9795), .A(n9738), .ZN(P1_U3223) );
  OAI21_X1 U10961 ( .B1(n9742), .B2(n9741), .A(n9740), .ZN(n9743) );
  NAND2_X1 U10962 ( .A1(n9743), .A2(n9802), .ZN(n9749) );
  NAND2_X1 U10963 ( .A1(n9786), .A2(n9817), .ZN(n9744) );
  NAND2_X1 U10964 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9855) );
  OAI211_X1 U10965 ( .C1(n9745), .C2(n9806), .A(n9744), .B(n9855), .ZN(n9746)
         );
  AOI21_X1 U10966 ( .B1(n9747), .B2(n9809), .A(n9746), .ZN(n9748) );
  OAI211_X1 U10967 ( .C1(n9750), .C2(n9812), .A(n9749), .B(n9748), .ZN(
        P1_U3226) );
  INV_X1 U10968 ( .A(n9751), .ZN(n9756) );
  NOR3_X1 U10969 ( .A1(n9754), .A2(n9753), .A3(n9752), .ZN(n9755) );
  OAI21_X1 U10970 ( .B1(n9756), .B2(n9755), .A(n9802), .ZN(n9760) );
  INV_X1 U10971 ( .A(n9990), .ZN(n9963) );
  AOI22_X1 U10972 ( .A1(n9768), .A2(n9963), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n9757) );
  OAI21_X1 U10973 ( .B1(n9989), .B2(n9804), .A(n9757), .ZN(n9758) );
  AOI21_X1 U10974 ( .B1(n9993), .B2(n9809), .A(n9758), .ZN(n9759) );
  OAI211_X1 U10975 ( .C1(n9996), .C2(n9812), .A(n9760), .B(n9759), .ZN(
        P1_U3227) );
  INV_X1 U10976 ( .A(n9761), .ZN(n9763) );
  NOR3_X1 U10977 ( .A1(n9764), .A2(n9763), .A3(n9762), .ZN(n9767) );
  INV_X1 U10978 ( .A(n9765), .ZN(n9766) );
  OAI21_X1 U10979 ( .B1(n9767), .B2(n9766), .A(n9802), .ZN(n9772) );
  AOI22_X1 U10980 ( .A1(n9768), .A2(n10057), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9769) );
  OAI21_X1 U10981 ( .B1(n9789), .B2(n9804), .A(n9769), .ZN(n9770) );
  AOI21_X1 U10982 ( .B1(n10047), .B2(n9809), .A(n9770), .ZN(n9771) );
  OAI211_X1 U10983 ( .C1(n10050), .C2(n9812), .A(n9772), .B(n9771), .ZN(
        P1_U3231) );
  NAND2_X1 U10984 ( .A1(n9774), .A2(n9773), .ZN(n9775) );
  XOR2_X1 U10985 ( .A(n9776), .B(n9775), .Z(n9781) );
  AOI22_X1 U10986 ( .A1(n9786), .A2(n10057), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9778) );
  NAND2_X1 U10987 ( .A1(n9809), .A2(n10016), .ZN(n9777) );
  OAI211_X1 U10988 ( .C1(n9989), .C2(n9806), .A(n9778), .B(n9777), .ZN(n9779)
         );
  AOI21_X1 U10989 ( .B1(n10092), .B2(n9792), .A(n9779), .ZN(n9780) );
  OAI21_X1 U10990 ( .B1(n9781), .B2(n9795), .A(n9780), .ZN(P1_U3233) );
  NAND2_X1 U10991 ( .A1(n9783), .A2(n9782), .ZN(n9785) );
  XNOR2_X1 U10992 ( .A(n9785), .B(n9784), .ZN(n9796) );
  NAND2_X1 U10993 ( .A1(n9786), .A2(n9816), .ZN(n9788) );
  NAND2_X1 U10994 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9874) );
  OAI211_X1 U10995 ( .C1(n9789), .C2(n9806), .A(n9788), .B(n9874), .ZN(n9790)
         );
  AOI21_X1 U10996 ( .B1(n9791), .B2(n9809), .A(n9790), .ZN(n9794) );
  NAND2_X1 U10997 ( .A1(n10112), .A2(n9792), .ZN(n9793) );
  OAI211_X1 U10998 ( .C1(n9796), .C2(n9795), .A(n9794), .B(n9793), .ZN(
        P1_U3236) );
  INV_X1 U10999 ( .A(n9797), .ZN(n9803) );
  OAI21_X1 U11000 ( .B1(n9800), .B2(n9799), .A(n9798), .ZN(n9801) );
  NAND3_X1 U11001 ( .A1(n9803), .A2(n9802), .A3(n9801), .ZN(n9811) );
  NOR2_X1 U11002 ( .A1(n9804), .A2(n9990), .ZN(n9808) );
  OAI22_X1 U11003 ( .A1(n9806), .A2(n9926), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9805), .ZN(n9807) );
  AOI211_X1 U11004 ( .C1(n9809), .C2(n9956), .A(n9808), .B(n9807), .ZN(n9810)
         );
  OAI211_X1 U11005 ( .C1(n9958), .C2(n9812), .A(n9811), .B(n9810), .ZN(
        P1_U3238) );
  MUX2_X1 U11006 ( .A(n9813), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9830), .Z(
        P1_U3585) );
  MUX2_X1 U11007 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n8490), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U11008 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9964), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U11009 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9814), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U11010 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9963), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U11011 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n10007), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U11012 ( .A(n10021), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9830), .Z(
        P1_U3578) );
  MUX2_X1 U11013 ( .A(n10037), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9830), .Z(
        P1_U3577) );
  MUX2_X1 U11014 ( .A(n10057), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9830), .Z(
        P1_U3576) );
  MUX2_X1 U11015 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n10036), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U11016 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n10055), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U11017 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9815), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U11018 ( .A(n9816), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9830), .Z(
        P1_U3572) );
  MUX2_X1 U11019 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9817), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U11020 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9818), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U11021 ( .A(n9819), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9830), .Z(
        P1_U3569) );
  MUX2_X1 U11022 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9820), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U11023 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9821), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U11024 ( .A(n9822), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9830), .Z(
        P1_U3566) );
  MUX2_X1 U11025 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9823), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U11026 ( .A(n9824), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9830), .Z(
        P1_U3564) );
  MUX2_X1 U11027 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9825), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U11028 ( .A(n9826), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9830), .Z(
        P1_U3562) );
  MUX2_X1 U11029 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9827), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U11030 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9828), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U11031 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9829), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U11032 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n7099), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U11033 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n7076), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U11034 ( .A(n6410), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9830), .Z(
        P1_U3556) );
  MUX2_X1 U11035 ( .A(n9831), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9830), .Z(
        P1_U3555) );
  NOR2_X1 U11036 ( .A1(n9833), .A2(n9832), .ZN(n9835) );
  XNOR2_X1 U11037 ( .A(n9858), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n9836) );
  AOI211_X1 U11038 ( .C1(n9837), .C2(n9836), .A(n10313), .B(n9857), .ZN(n9851)
         );
  INV_X1 U11039 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9849) );
  NAND2_X1 U11040 ( .A1(n9839), .A2(n9838), .ZN(n9841) );
  NAND2_X1 U11041 ( .A1(n9841), .A2(n9840), .ZN(n9844) );
  INV_X1 U11042 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9842) );
  MUX2_X1 U11043 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9842), .S(n9858), .Z(n9843) );
  NAND2_X1 U11044 ( .A1(n9844), .A2(n9843), .ZN(n9852) );
  OAI211_X1 U11045 ( .C1(n9844), .C2(n9843), .A(n9852), .B(n10319), .ZN(n9848)
         );
  INV_X1 U11046 ( .A(n9845), .ZN(n9846) );
  AOI21_X1 U11047 ( .B1(n10310), .B2(n9858), .A(n9846), .ZN(n9847) );
  OAI211_X1 U11048 ( .C1(n9849), .C2(n10305), .A(n9848), .B(n9847), .ZN(n9850)
         );
  OR2_X1 U11049 ( .A1(n9851), .A2(n9850), .ZN(P1_U3257) );
  OAI21_X1 U11050 ( .B1(n9842), .B2(n9853), .A(n9852), .ZN(n9868) );
  XNOR2_X1 U11051 ( .A(n9877), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9866) );
  XNOR2_X1 U11052 ( .A(n9868), .B(n9866), .ZN(n9864) );
  INV_X1 U11053 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9856) );
  NAND2_X1 U11054 ( .A1(n9877), .A2(n10310), .ZN(n9854) );
  OAI211_X1 U11055 ( .C1(n10305), .C2(n9856), .A(n9855), .B(n9854), .ZN(n9863)
         );
  NAND2_X1 U11056 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9877), .ZN(n9859) );
  OAI21_X1 U11057 ( .B1(n9877), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9859), .ZN(
        n9860) );
  AOI211_X1 U11058 ( .C1(n9861), .C2(n9860), .A(n10313), .B(n9876), .ZN(n9862)
         );
  AOI211_X1 U11059 ( .C1(n10319), .C2(n9864), .A(n9863), .B(n9862), .ZN(n9865)
         );
  INV_X1 U11060 ( .A(n9865), .ZN(P1_U3258) );
  INV_X1 U11061 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9888) );
  AOI22_X1 U11062 ( .A1(n9892), .A2(n9888), .B1(P1_REG1_REG_18__SCAN_IN), .B2(
        n9887), .ZN(n9873) );
  INV_X1 U11063 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9870) );
  INV_X1 U11064 ( .A(n9866), .ZN(n9867) );
  NAND2_X1 U11065 ( .A1(n9868), .A2(n9867), .ZN(n9869) );
  OAI21_X1 U11066 ( .B1(n9871), .B2(n9870), .A(n9869), .ZN(n9872) );
  NOR2_X1 U11067 ( .A1(n9873), .A2(n9872), .ZN(n9886) );
  AOI21_X1 U11068 ( .B1(n9873), .B2(n9872), .A(n9886), .ZN(n9885) );
  NAND2_X1 U11069 ( .A1(n9892), .A2(n10310), .ZN(n9875) );
  NAND2_X1 U11070 ( .A1(n9875), .A2(n9874), .ZN(n9883) );
  AOI21_X1 U11071 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n9877), .A(n9876), .ZN(
        n9881) );
  INV_X1 U11072 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9878) );
  MUX2_X1 U11073 ( .A(P1_REG2_REG_18__SCAN_IN), .B(n9878), .S(n9892), .Z(n9879) );
  INV_X1 U11074 ( .A(n9879), .ZN(n9880) );
  NOR2_X1 U11075 ( .A1(n9881), .A2(n9880), .ZN(n9891) );
  AOI211_X1 U11076 ( .C1(n9881), .C2(n9880), .A(n9891), .B(n10313), .ZN(n9882)
         );
  AOI211_X1 U11077 ( .C1(n10312), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n9883), .B(
        n9882), .ZN(n9884) );
  OAI21_X1 U11078 ( .B1(n9885), .B2(n9895), .A(n9884), .ZN(P1_U3259) );
  AOI21_X1 U11079 ( .B1(n9888), .B2(n9887), .A(n9886), .ZN(n9890) );
  XOR2_X1 U11080 ( .A(n9890), .B(n9889), .Z(n9898) );
  AOI21_X1 U11081 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n9892), .A(n9891), .ZN(
        n9893) );
  XNOR2_X1 U11082 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9893), .ZN(n9901) );
  NAND2_X1 U11083 ( .A1(n9901), .A2(n10294), .ZN(n9894) );
  NAND2_X1 U11084 ( .A1(n9897), .A2(n9896), .ZN(n9900) );
  OAI21_X1 U11085 ( .B1(n10305), .B2(n9904), .A(n9903), .ZN(n9905) );
  NAND2_X1 U11086 ( .A1(n10262), .A2(n9912), .ZN(n9907) );
  XNOR2_X1 U11087 ( .A(n9906), .B(n9907), .ZN(n10212) );
  NAND2_X1 U11088 ( .A1(n10212), .A2(n10331), .ZN(n9911) );
  NAND2_X1 U11089 ( .A1(n9909), .A2(n9908), .ZN(n10261) );
  NOR2_X1 U11090 ( .A1(n10048), .A2(n10261), .ZN(n9914) );
  AOI21_X1 U11091 ( .B1(n10048), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9914), .ZN(
        n9910) );
  OAI211_X1 U11092 ( .C1(n10256), .C2(n9906), .A(n9911), .B(n9910), .ZN(
        P1_U3261) );
  XNOR2_X1 U11093 ( .A(n9913), .B(n9912), .ZN(n10264) );
  NAND2_X1 U11094 ( .A1(n10264), .A2(n10331), .ZN(n9916) );
  AOI21_X1 U11095 ( .B1(n10048), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9914), .ZN(
        n9915) );
  OAI211_X1 U11096 ( .C1(n10262), .C2(n10256), .A(n9916), .B(n9915), .ZN(
        P1_U3262) );
  INV_X1 U11097 ( .A(n9917), .ZN(n9920) );
  INV_X1 U11098 ( .A(n9922), .ZN(n9919) );
  INV_X1 U11099 ( .A(n9921), .ZN(n9925) );
  AOI21_X1 U11100 ( .B1(n9947), .B2(n9923), .A(n9922), .ZN(n9924) );
  AOI211_X1 U11101 ( .C1(n10065), .C2(n9938), .A(n10416), .B(n9928), .ZN(
        n10064) );
  NAND2_X1 U11102 ( .A1(n10064), .A2(n10041), .ZN(n9931) );
  AOI22_X1 U11103 ( .A1(n10048), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9929), 
        .B2(n10345), .ZN(n9930) );
  OAI211_X1 U11104 ( .C1(n9932), .C2(n10256), .A(n9931), .B(n9930), .ZN(n9933)
         );
  AOI21_X1 U11105 ( .B1(n10063), .B2(n10349), .A(n9933), .ZN(n9934) );
  OAI21_X1 U11106 ( .B1(n10066), .B2(n10062), .A(n9934), .ZN(P1_U3263) );
  OAI21_X1 U11107 ( .B1(n9936), .B2(n9943), .A(n9935), .ZN(n9937) );
  INV_X1 U11108 ( .A(n9937), .ZN(n10071) );
  INV_X1 U11109 ( .A(n9938), .ZN(n9939) );
  AOI21_X1 U11110 ( .B1(n10067), .B2(n9955), .A(n9939), .ZN(n10068) );
  AOI22_X1 U11111 ( .A1(n10048), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9940), 
        .B2(n10345), .ZN(n9941) );
  OAI21_X1 U11112 ( .B1(n4563), .B2(n10256), .A(n9941), .ZN(n9950) );
  INV_X1 U11113 ( .A(n9942), .ZN(n9944) );
  AOI21_X1 U11114 ( .B1(n9944), .B2(n9943), .A(n9988), .ZN(n9948) );
  OAI22_X1 U11115 ( .A1(n9974), .A2(n10340), .B1(n9945), .B2(n10338), .ZN(
        n9946) );
  AOI21_X1 U11116 ( .B1(n9948), .B2(n9947), .A(n9946), .ZN(n10070) );
  NOR2_X1 U11117 ( .A1(n10070), .A2(n10048), .ZN(n9949) );
  AOI211_X1 U11118 ( .C1(n10068), .C2(n10331), .A(n9950), .B(n9949), .ZN(n9951) );
  OAI21_X1 U11119 ( .B1(n10071), .B2(n10062), .A(n9951), .ZN(P1_U3264) );
  OAI21_X1 U11120 ( .B1(n9953), .B2(n9961), .A(n9952), .ZN(n9954) );
  INV_X1 U11121 ( .A(n9954), .ZN(n10076) );
  AOI21_X1 U11122 ( .B1(n10072), .B2(n9975), .A(n4564), .ZN(n10073) );
  AOI22_X1 U11123 ( .A1(n10048), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9956), 
        .B2(n10345), .ZN(n9957) );
  OAI21_X1 U11124 ( .B1(n9958), .B2(n10256), .A(n9957), .ZN(n9967) );
  NAND2_X1 U11125 ( .A1(n9960), .A2(n9959), .ZN(n9962) );
  XNOR2_X1 U11126 ( .A(n9962), .B(n9961), .ZN(n9965) );
  AOI222_X1 U11127 ( .A1(n10343), .A2(n9965), .B1(n9964), .B2(n10056), .C1(
        n9963), .C2(n10054), .ZN(n10075) );
  NOR2_X1 U11128 ( .A1(n10075), .A2(n10048), .ZN(n9966) );
  AOI211_X1 U11129 ( .C1(n10073), .C2(n10331), .A(n9967), .B(n9966), .ZN(n9968) );
  OAI21_X1 U11130 ( .B1(n10076), .B2(n10062), .A(n9968), .ZN(P1_U3265) );
  XOR2_X1 U11131 ( .A(n9971), .B(n9969), .Z(n10081) );
  XOR2_X1 U11132 ( .A(n9971), .B(n9970), .Z(n9972) );
  OAI222_X1 U11133 ( .A1(n10338), .A2(n9974), .B1(n10340), .B2(n9973), .C1(
        n9972), .C2(n9988), .ZN(n10077) );
  INV_X1 U11134 ( .A(n9991), .ZN(n9976) );
  AOI211_X1 U11135 ( .C1(n10079), .C2(n9976), .A(n10416), .B(n4912), .ZN(
        n10078) );
  NAND2_X1 U11136 ( .A1(n10078), .A2(n10041), .ZN(n9979) );
  AOI22_X1 U11137 ( .A1(n10048), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9977), 
        .B2(n10345), .ZN(n9978) );
  OAI211_X1 U11138 ( .C1(n9980), .C2(n10256), .A(n9979), .B(n9978), .ZN(n9981)
         );
  AOI21_X1 U11139 ( .B1(n10077), .B2(n10349), .A(n9981), .ZN(n9982) );
  OAI21_X1 U11140 ( .B1(n10081), .B2(n10062), .A(n9982), .ZN(P1_U3266) );
  XNOR2_X1 U11141 ( .A(n9983), .B(n9986), .ZN(n10086) );
  AOI21_X1 U11142 ( .B1(n9986), .B2(n9985), .A(n9984), .ZN(n9987) );
  OAI222_X1 U11143 ( .A1(n10338), .A2(n9990), .B1(n10340), .B2(n9989), .C1(
        n9988), .C2(n9987), .ZN(n10082) );
  INV_X1 U11144 ( .A(n10000), .ZN(n9992) );
  AOI211_X1 U11145 ( .C1(n10084), .C2(n9992), .A(n10416), .B(n9991), .ZN(
        n10083) );
  NAND2_X1 U11146 ( .A1(n10083), .A2(n10041), .ZN(n9995) );
  AOI22_X1 U11147 ( .A1(n10048), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9993), 
        .B2(n10345), .ZN(n9994) );
  OAI211_X1 U11148 ( .C1(n9996), .C2(n10256), .A(n9995), .B(n9994), .ZN(n9997)
         );
  AOI21_X1 U11149 ( .B1(n10082), .B2(n10349), .A(n9997), .ZN(n9998) );
  OAI21_X1 U11150 ( .B1(n10086), .B2(n10062), .A(n9998), .ZN(P1_U3267) );
  XOR2_X1 U11151 ( .A(n9999), .B(n10005), .Z(n10091) );
  AOI21_X1 U11152 ( .B1(n10087), .B2(n10014), .A(n10000), .ZN(n10088) );
  AOI22_X1 U11153 ( .A1(n10048), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n10001), 
        .B2(n10345), .ZN(n10002) );
  OAI21_X1 U11154 ( .B1(n10003), .B2(n10256), .A(n10002), .ZN(n10011) );
  OAI211_X1 U11155 ( .C1(n10006), .C2(n10005), .A(n10004), .B(n10343), .ZN(
        n10009) );
  AOI22_X1 U11156 ( .A1(n10007), .A2(n10056), .B1(n10054), .B2(n10037), .ZN(
        n10008) );
  AND2_X1 U11157 ( .A1(n10009), .A2(n10008), .ZN(n10090) );
  NOR2_X1 U11158 ( .A1(n10090), .A2(n10048), .ZN(n10010) );
  AOI211_X1 U11159 ( .C1(n10088), .C2(n10331), .A(n10011), .B(n10010), .ZN(
        n10012) );
  OAI21_X1 U11160 ( .B1(n10091), .B2(n10062), .A(n10012), .ZN(P1_U3268) );
  XOR2_X1 U11161 ( .A(n10013), .B(n10019), .Z(n10096) );
  INV_X1 U11162 ( .A(n10014), .ZN(n10015) );
  AOI21_X1 U11163 ( .B1(n10092), .B2(n10027), .A(n10015), .ZN(n10093) );
  AOI22_X1 U11164 ( .A1(n10048), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n10016), 
        .B2(n10345), .ZN(n10017) );
  OAI21_X1 U11165 ( .B1(n10018), .B2(n10256), .A(n10017), .ZN(n10024) );
  XNOR2_X1 U11166 ( .A(n10020), .B(n10019), .ZN(n10022) );
  AOI222_X1 U11167 ( .A1(n10343), .A2(n10022), .B1(n10021), .B2(n10056), .C1(
        n10057), .C2(n10054), .ZN(n10095) );
  NOR2_X1 U11168 ( .A1(n10095), .A2(n10048), .ZN(n10023) );
  AOI211_X1 U11169 ( .C1(n10093), .C2(n10331), .A(n10024), .B(n10023), .ZN(
        n10025) );
  OAI21_X1 U11170 ( .B1(n10096), .B2(n10062), .A(n10025), .ZN(P1_U3269) );
  XNOR2_X1 U11171 ( .A(n10026), .B(n10035), .ZN(n10101) );
  INV_X1 U11172 ( .A(n10046), .ZN(n10029) );
  INV_X1 U11173 ( .A(n10027), .ZN(n10028) );
  AOI211_X1 U11174 ( .C1(n10098), .C2(n10029), .A(n10416), .B(n10028), .ZN(
        n10097) );
  AOI22_X1 U11175 ( .A1(n10048), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n10030), 
        .B2(n10345), .ZN(n10031) );
  OAI21_X1 U11176 ( .B1(n10032), .B2(n10256), .A(n10031), .ZN(n10040) );
  OAI21_X1 U11177 ( .B1(n10035), .B2(n10034), .A(n10033), .ZN(n10038) );
  AOI222_X1 U11178 ( .A1(n10343), .A2(n10038), .B1(n10037), .B2(n10056), .C1(
        n10036), .C2(n10054), .ZN(n10100) );
  NOR2_X1 U11179 ( .A1(n10100), .A2(n10048), .ZN(n10039) );
  AOI211_X1 U11180 ( .C1(n10097), .C2(n10041), .A(n10040), .B(n10039), .ZN(
        n10042) );
  OAI21_X1 U11181 ( .B1(n10101), .B2(n10062), .A(n10042), .ZN(P1_U3270) );
  XNOR2_X1 U11182 ( .A(n10044), .B(n10043), .ZN(n10106) );
  AOI21_X1 U11183 ( .B1(n10102), .B2(n4907), .A(n10046), .ZN(n10103) );
  AOI22_X1 U11184 ( .A1(n10048), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n10047), 
        .B2(n10345), .ZN(n10049) );
  OAI21_X1 U11185 ( .B1(n10050), .B2(n10256), .A(n10049), .ZN(n10060) );
  OAI21_X1 U11186 ( .B1(n10053), .B2(n10052), .A(n10051), .ZN(n10058) );
  AOI222_X1 U11187 ( .A1(n10343), .A2(n10058), .B1(n10057), .B2(n10056), .C1(
        n10055), .C2(n10054), .ZN(n10105) );
  NOR2_X1 U11188 ( .A1(n10105), .A2(n10048), .ZN(n10059) );
  AOI211_X1 U11189 ( .C1(n10103), .C2(n10331), .A(n10060), .B(n10059), .ZN(
        n10061) );
  OAI21_X1 U11190 ( .B1(n10106), .B2(n10062), .A(n10061), .ZN(P1_U3271) );
  INV_X1 U11191 ( .A(n10401), .ZN(n10412) );
  MUX2_X1 U11192 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n10138), .S(n10438), .Z(
        P1_U3551) );
  AOI22_X1 U11193 ( .A1(n10068), .A2(n10265), .B1(n10133), .B2(n10067), .ZN(
        n10069) );
  OAI211_X1 U11194 ( .C1(n10071), .C2(n10412), .A(n10070), .B(n10069), .ZN(
        n10139) );
  MUX2_X1 U11195 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10139), .S(n10438), .Z(
        P1_U3550) );
  AOI22_X1 U11196 ( .A1(n10073), .A2(n10265), .B1(n10133), .B2(n10072), .ZN(
        n10074) );
  OAI211_X1 U11197 ( .C1(n10076), .C2(n10412), .A(n10075), .B(n10074), .ZN(
        n10140) );
  MUX2_X1 U11198 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10140), .S(n10438), .Z(
        P1_U3549) );
  AOI211_X1 U11199 ( .C1(n10133), .C2(n10079), .A(n10078), .B(n10077), .ZN(
        n10080) );
  OAI21_X1 U11200 ( .B1(n10081), .B2(n10412), .A(n10080), .ZN(n10141) );
  MUX2_X1 U11201 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10141), .S(n10438), .Z(
        P1_U3548) );
  AOI211_X1 U11202 ( .C1(n10133), .C2(n10084), .A(n10083), .B(n10082), .ZN(
        n10085) );
  OAI21_X1 U11203 ( .B1(n10086), .B2(n10412), .A(n10085), .ZN(n10142) );
  MUX2_X1 U11204 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10142), .S(n10438), .Z(
        P1_U3547) );
  AOI22_X1 U11205 ( .A1(n10088), .A2(n10265), .B1(n10133), .B2(n10087), .ZN(
        n10089) );
  OAI211_X1 U11206 ( .C1(n10091), .C2(n10412), .A(n10090), .B(n10089), .ZN(
        n10143) );
  MUX2_X1 U11207 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10143), .S(n10438), .Z(
        P1_U3546) );
  AOI22_X1 U11208 ( .A1(n10093), .A2(n10265), .B1(n10133), .B2(n10092), .ZN(
        n10094) );
  OAI211_X1 U11209 ( .C1(n10096), .C2(n10412), .A(n10095), .B(n10094), .ZN(
        n10144) );
  MUX2_X1 U11210 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10144), .S(n10438), .Z(
        P1_U3545) );
  AOI21_X1 U11211 ( .B1(n10133), .B2(n10098), .A(n10097), .ZN(n10099) );
  OAI211_X1 U11212 ( .C1(n10101), .C2(n10412), .A(n10100), .B(n10099), .ZN(
        n10145) );
  MUX2_X1 U11213 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10145), .S(n10438), .Z(
        P1_U3544) );
  AOI22_X1 U11214 ( .A1(n10103), .A2(n10265), .B1(n10133), .B2(n10102), .ZN(
        n10104) );
  OAI211_X1 U11215 ( .C1(n10106), .C2(n10412), .A(n10105), .B(n10104), .ZN(
        n10146) );
  MUX2_X1 U11216 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10146), .S(n10438), .Z(
        P1_U3543) );
  AOI21_X1 U11217 ( .B1(n10133), .B2(n10108), .A(n10107), .ZN(n10109) );
  OAI211_X1 U11218 ( .C1(n10111), .C2(n10412), .A(n10110), .B(n10109), .ZN(
        n10147) );
  MUX2_X1 U11219 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10147), .S(n10438), .Z(
        P1_U3542) );
  AOI22_X1 U11220 ( .A1(n10113), .A2(n10265), .B1(n10133), .B2(n10112), .ZN(
        n10114) );
  OAI211_X1 U11221 ( .C1(n10116), .C2(n10412), .A(n10115), .B(n10114), .ZN(
        n10148) );
  MUX2_X1 U11222 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10148), .S(n10438), .Z(
        P1_U3541) );
  AOI211_X1 U11223 ( .C1(n10133), .C2(n10119), .A(n10118), .B(n10117), .ZN(
        n10120) );
  OAI21_X1 U11224 ( .B1(n10121), .B2(n10412), .A(n10120), .ZN(n10149) );
  MUX2_X1 U11225 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10149), .S(n10438), .Z(
        P1_U3540) );
  AOI22_X1 U11226 ( .A1(n10123), .A2(n10265), .B1(n10133), .B2(n10122), .ZN(
        n10124) );
  OAI211_X1 U11227 ( .C1(n10368), .C2(n10126), .A(n10125), .B(n10124), .ZN(
        n10150) );
  MUX2_X1 U11228 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n10150), .S(n10438), .Z(
        P1_U3538) );
  AOI211_X1 U11229 ( .C1(n10133), .C2(n10129), .A(n10128), .B(n10127), .ZN(
        n10130) );
  OAI21_X1 U11230 ( .B1(n10131), .B2(n10412), .A(n10130), .ZN(n10151) );
  MUX2_X1 U11231 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10151), .S(n10438), .Z(
        P1_U3537) );
  AOI22_X1 U11232 ( .A1(n10134), .A2(n10265), .B1(n10133), .B2(n10132), .ZN(
        n10135) );
  OAI211_X1 U11233 ( .C1(n10368), .C2(n10137), .A(n10136), .B(n10135), .ZN(
        n10152) );
  MUX2_X1 U11234 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10152), .S(n10438), .Z(
        P1_U3535) );
  MUX2_X1 U11235 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n10138), .S(n10424), .Z(
        P1_U3519) );
  MUX2_X1 U11236 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10139), .S(n10424), .Z(
        P1_U3518) );
  MUX2_X1 U11237 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10140), .S(n10424), .Z(
        P1_U3517) );
  MUX2_X1 U11238 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10141), .S(n10424), .Z(
        P1_U3516) );
  MUX2_X1 U11239 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10142), .S(n10424), .Z(
        P1_U3515) );
  MUX2_X1 U11240 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10143), .S(n10424), .Z(
        P1_U3514) );
  MUX2_X1 U11241 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10144), .S(n10424), .Z(
        P1_U3513) );
  MUX2_X1 U11242 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10145), .S(n10424), .Z(
        P1_U3512) );
  MUX2_X1 U11243 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10146), .S(n10424), .Z(
        P1_U3511) );
  MUX2_X1 U11244 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10147), .S(n10424), .Z(
        P1_U3510) );
  MUX2_X1 U11245 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10148), .S(n10424), .Z(
        P1_U3508) );
  MUX2_X1 U11246 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10149), .S(n10424), .Z(
        P1_U3505) );
  MUX2_X1 U11247 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n10150), .S(n10424), .Z(
        P1_U3499) );
  MUX2_X1 U11248 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10151), .S(n10424), .Z(
        P1_U3496) );
  MUX2_X1 U11249 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n10152), .S(n10424), .Z(
        P1_U3490) );
  NOR4_X1 U11250 ( .A1(n10153), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), 
        .A4(n6113), .ZN(n10154) );
  AOI21_X1 U11251 ( .B1(n10155), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n10154), 
        .ZN(n10156) );
  OAI21_X1 U11252 ( .B1(n10158), .B2(n10157), .A(n10156), .ZN(P1_U3322) );
  MUX2_X1 U11253 ( .A(n10159), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  AOI22_X1 U11254 ( .A1(n10441), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n10171) );
  AOI211_X1 U11255 ( .C1(n10162), .C2(n10161), .A(n10160), .B(n10442), .ZN(
        n10163) );
  AOI21_X1 U11256 ( .B1(n10165), .B2(n10164), .A(n10163), .ZN(n10170) );
  OAI211_X1 U11257 ( .C1(n10168), .C2(n10167), .A(n10439), .B(n10166), .ZN(
        n10169) );
  NAND3_X1 U11258 ( .A1(n10171), .A2(n10170), .A3(n10169), .ZN(P2_U3247) );
  OAI22_X1 U11259 ( .A1(n10173), .A2(n10416), .B1(n10172), .B2(n10414), .ZN(
        n10174) );
  AOI21_X1 U11260 ( .B1(n10175), .B2(n10410), .A(n10174), .ZN(n10176) );
  AND2_X1 U11261 ( .A1(n10177), .A2(n10176), .ZN(n10180) );
  AOI22_X1 U11262 ( .A1(n10424), .A2(n10180), .B1(n10178), .B2(n10422), .ZN(
        P1_U3484) );
  AOI22_X1 U11263 ( .A1(n10438), .A2(n10180), .B1(n10179), .B2(n10436), .ZN(
        P1_U3533) );
  NOR2_X1 U11264 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10181) );
  AOI21_X1 U11265 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n10181), .ZN(n10548) );
  NOR2_X1 U11266 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10182) );
  AOI21_X1 U11267 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n10182), .ZN(n10551) );
  NOR2_X1 U11268 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10183) );
  AOI21_X1 U11269 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n10183), .ZN(n10554) );
  NOR2_X1 U11270 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(P2_ADDR_REG_14__SCAN_IN), 
        .ZN(n10184) );
  AOI21_X1 U11271 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10184), .ZN(n10557) );
  NOR2_X1 U11272 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(P2_ADDR_REG_13__SCAN_IN), 
        .ZN(n10185) );
  AOI21_X1 U11273 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10185), .ZN(n10560) );
  NOR2_X1 U11274 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10191) );
  XNOR2_X1 U11275 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10590) );
  NAND2_X1 U11276 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n10189) );
  XOR2_X1 U11277 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(P1_ADDR_REG_3__SCAN_IN), .Z(
        n10588) );
  NAND2_X1 U11278 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n10187) );
  XOR2_X1 U11279 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10586) );
  AOI21_X1 U11280 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10542) );
  NAND3_X1 U11281 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10544) );
  OAI21_X1 U11282 ( .B1(n10542), .B2(n8133), .A(n10544), .ZN(n10585) );
  NAND2_X1 U11283 ( .A1(n10586), .A2(n10585), .ZN(n10186) );
  NAND2_X1 U11284 ( .A1(n10187), .A2(n10186), .ZN(n10587) );
  NAND2_X1 U11285 ( .A1(n10588), .A2(n10587), .ZN(n10188) );
  NAND2_X1 U11286 ( .A1(n10189), .A2(n10188), .ZN(n10589) );
  NOR2_X1 U11287 ( .A1(n10590), .A2(n10589), .ZN(n10190) );
  NOR2_X1 U11288 ( .A1(n10191), .A2(n10190), .ZN(n10192) );
  NOR2_X1 U11289 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10192), .ZN(n10572) );
  AND2_X1 U11290 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10192), .ZN(n10571) );
  NOR2_X1 U11291 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10571), .ZN(n10193) );
  NOR2_X1 U11292 ( .A1(n10572), .A2(n10193), .ZN(n10194) );
  NAND2_X1 U11293 ( .A1(n10194), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n10196) );
  XOR2_X1 U11294 ( .A(n10194), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10570) );
  NAND2_X1 U11295 ( .A1(n10570), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n10195) );
  NAND2_X1 U11296 ( .A1(n10196), .A2(n10195), .ZN(n10197) );
  NAND2_X1 U11297 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n10197), .ZN(n10199) );
  XOR2_X1 U11298 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n10197), .Z(n10584) );
  NAND2_X1 U11299 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10584), .ZN(n10198) );
  NAND2_X1 U11300 ( .A1(n10199), .A2(n10198), .ZN(n10200) );
  AND2_X1 U11301 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10200), .ZN(n10201) );
  XNOR2_X1 U11302 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10200), .ZN(n10582) );
  NOR2_X1 U11303 ( .A1(n10583), .A2(n10582), .ZN(n10581) );
  NOR2_X1 U11304 ( .A1(n10201), .A2(n10581), .ZN(n10202) );
  INV_X1 U11305 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10203) );
  NOR2_X1 U11306 ( .A1(n10202), .A2(n10203), .ZN(n10204) );
  XNOR2_X1 U11307 ( .A(n10203), .B(n10202), .ZN(n10579) );
  NOR2_X1 U11308 ( .A1(n10580), .A2(n10579), .ZN(n10578) );
  NOR2_X1 U11309 ( .A1(n10204), .A2(n10578), .ZN(n10569) );
  NAND2_X1 U11310 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n10205) );
  OAI21_X1 U11311 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10205), .ZN(n10568) );
  NOR2_X1 U11312 ( .A1(n10569), .A2(n10568), .ZN(n10567) );
  AOI21_X1 U11313 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n10567), .ZN(n10566) );
  NAND2_X1 U11314 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n10206) );
  OAI21_X1 U11315 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n10206), .ZN(n10565) );
  NOR2_X1 U11316 ( .A1(n10566), .A2(n10565), .ZN(n10564) );
  AOI21_X1 U11317 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10564), .ZN(n10563) );
  NOR2_X1 U11318 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10207) );
  AOI21_X1 U11319 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n10207), .ZN(n10562) );
  NAND2_X1 U11320 ( .A1(n10563), .A2(n10562), .ZN(n10561) );
  OAI21_X1 U11321 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10561), .ZN(n10559) );
  NAND2_X1 U11322 ( .A1(n10560), .A2(n10559), .ZN(n10558) );
  OAI21_X1 U11323 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n10558), .ZN(n10556) );
  NAND2_X1 U11324 ( .A1(n10557), .A2(n10556), .ZN(n10555) );
  OAI21_X1 U11325 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n10555), .ZN(n10553) );
  NAND2_X1 U11326 ( .A1(n10554), .A2(n10553), .ZN(n10552) );
  OAI21_X1 U11327 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10552), .ZN(n10550) );
  NAND2_X1 U11328 ( .A1(n10551), .A2(n10550), .ZN(n10549) );
  OAI21_X1 U11329 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10549), .ZN(n10547) );
  NAND2_X1 U11330 ( .A1(n10548), .A2(n10547), .ZN(n10546) );
  OAI21_X1 U11331 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10546), .ZN(n10575) );
  NOR2_X1 U11332 ( .A1(n10576), .A2(n10575), .ZN(n10208) );
  NAND2_X1 U11333 ( .A1(n10576), .A2(n10575), .ZN(n10574) );
  OAI21_X1 U11334 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n10208), .A(n10574), 
        .ZN(n10210) );
  XOR2_X1 U11335 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .Z(n10209) );
  XNOR2_X1 U11336 ( .A(n10210), .B(n10209), .ZN(ADD_1071_U4) );
  OAI21_X1 U11337 ( .B1(n9906), .B2(n10414), .A(n10261), .ZN(n10211) );
  AOI21_X1 U11338 ( .B1(n10212), .B2(n10265), .A(n10211), .ZN(n10215) );
  INV_X1 U11339 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n10213) );
  AOI22_X1 U11340 ( .A1(n10438), .A2(n10215), .B1(n10213), .B2(n10436), .ZN(
        P1_U3554) );
  INV_X1 U11341 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n10214) );
  AOI22_X1 U11342 ( .A1(n10424), .A2(n10215), .B1(n10214), .B2(n10422), .ZN(
        P1_U3522) );
  INV_X1 U11343 ( .A(n10216), .ZN(n10228) );
  INV_X1 U11344 ( .A(n10217), .ZN(n10219) );
  AOI22_X1 U11345 ( .A1(n4499), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n10219), 
        .B2(n10218), .ZN(n10223) );
  NAND2_X1 U11346 ( .A1(n10221), .A2(n10220), .ZN(n10222) );
  OAI211_X1 U11347 ( .C1(n10225), .C2(n10224), .A(n10223), .B(n10222), .ZN(
        n10226) );
  AOI21_X1 U11348 ( .B1(n10228), .B2(n10227), .A(n10226), .ZN(n10229) );
  OAI21_X1 U11349 ( .B1(n4499), .B2(n10230), .A(n10229), .ZN(P2_U3283) );
  NOR2_X1 U11350 ( .A1(n4940), .A2(n10518), .ZN(n10232) );
  AOI211_X1 U11351 ( .C1(n10233), .C2(n10524), .A(n10232), .B(n10231), .ZN(
        n10235) );
  AOI22_X1 U11352 ( .A1(n10541), .A2(n10235), .B1(n10234), .B2(n10539), .ZN(
        P2_U3537) );
  AOI22_X1 U11353 ( .A1(n10528), .A2(n10235), .B1(n5536), .B2(n10526), .ZN(
        P2_U3502) );
  XNOR2_X1 U11354 ( .A(n10236), .B(n10244), .ZN(n10280) );
  NAND2_X1 U11355 ( .A1(n10238), .A2(n10237), .ZN(n10239) );
  NAND2_X1 U11356 ( .A1(n10240), .A2(n10239), .ZN(n10278) );
  INV_X1 U11357 ( .A(n10278), .ZN(n10241) );
  AOI22_X1 U11358 ( .A1(n10280), .A2(n10332), .B1(n10331), .B2(n10241), .ZN(
        n10260) );
  NAND2_X1 U11359 ( .A1(n10243), .A2(n10242), .ZN(n10245) );
  NAND2_X1 U11360 ( .A1(n10245), .A2(n10244), .ZN(n10247) );
  NAND3_X1 U11361 ( .A1(n10247), .A2(n10343), .A3(n10246), .ZN(n10251) );
  OAI22_X1 U11362 ( .A1(n10339), .A2(n10340), .B1(n10248), .B2(n10338), .ZN(
        n10249) );
  INV_X1 U11363 ( .A(n10249), .ZN(n10250) );
  NAND2_X1 U11364 ( .A1(n10251), .A2(n10250), .ZN(n10252) );
  AOI21_X1 U11365 ( .B1(n10280), .B2(n10253), .A(n10252), .ZN(n10282) );
  INV_X1 U11366 ( .A(n10282), .ZN(n10258) );
  AOI22_X1 U11367 ( .A1(n10048), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n10254), 
        .B2(n10345), .ZN(n10255) );
  OAI21_X1 U11368 ( .B1(n10277), .B2(n10256), .A(n10255), .ZN(n10257) );
  AOI21_X1 U11369 ( .B1(n10258), .B2(n10349), .A(n10257), .ZN(n10259) );
  NAND2_X1 U11370 ( .A1(n10260), .A2(n10259), .ZN(P1_U3280) );
  OAI21_X1 U11371 ( .B1(n10262), .B2(n10414), .A(n10261), .ZN(n10263) );
  AOI21_X1 U11372 ( .B1(n10265), .B2(n10264), .A(n10263), .ZN(n10284) );
  AOI22_X1 U11373 ( .A1(n10438), .A2(n10284), .B1(n6225), .B2(n10436), .ZN(
        P1_U3553) );
  OAI211_X1 U11374 ( .C1(n4672), .C2(n10414), .A(n10267), .B(n10266), .ZN(
        n10268) );
  AOI21_X1 U11375 ( .B1(n10269), .B2(n10401), .A(n10268), .ZN(n10286) );
  AOI22_X1 U11376 ( .A1(n10438), .A2(n10286), .B1(n9842), .B2(n10436), .ZN(
        P1_U3539) );
  INV_X1 U11377 ( .A(n10270), .ZN(n10271) );
  OAI22_X1 U11378 ( .A1(n10272), .A2(n10416), .B1(n10271), .B2(n10414), .ZN(
        n10273) );
  AOI21_X1 U11379 ( .B1(n10274), .B2(n10410), .A(n10273), .ZN(n10275) );
  AND2_X1 U11380 ( .A1(n10276), .A2(n10275), .ZN(n10288) );
  AOI22_X1 U11381 ( .A1(n10438), .A2(n10288), .B1(n7599), .B2(n10436), .ZN(
        P1_U3536) );
  OAI22_X1 U11382 ( .A1(n10278), .A2(n10416), .B1(n10277), .B2(n10414), .ZN(
        n10279) );
  AOI21_X1 U11383 ( .B1(n10280), .B2(n10410), .A(n10279), .ZN(n10281) );
  AND2_X1 U11384 ( .A1(n10282), .A2(n10281), .ZN(n10290) );
  AOI22_X1 U11385 ( .A1(n10438), .A2(n10290), .B1(n7300), .B2(n10436), .ZN(
        P1_U3534) );
  INV_X1 U11386 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10283) );
  AOI22_X1 U11387 ( .A1(n10424), .A2(n10284), .B1(n10283), .B2(n10422), .ZN(
        P1_U3521) );
  INV_X1 U11388 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n10285) );
  AOI22_X1 U11389 ( .A1(n10424), .A2(n10286), .B1(n10285), .B2(n10422), .ZN(
        P1_U3502) );
  INV_X1 U11390 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10287) );
  AOI22_X1 U11391 ( .A1(n10424), .A2(n10288), .B1(n10287), .B2(n10422), .ZN(
        P1_U3493) );
  AOI22_X1 U11392 ( .A1(n10424), .A2(n10290), .B1(n10289), .B2(n10422), .ZN(
        P1_U3487) );
  XNOR2_X1 U11393 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11394 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  OAI21_X1 U11395 ( .B1(n10292), .B2(n4520), .A(n10291), .ZN(n10295) );
  AOI22_X1 U11396 ( .A1(n10295), .A2(n10294), .B1(n10293), .B2(n10310), .ZN(
        n10309) );
  INV_X1 U11397 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10304) );
  NAND2_X1 U11398 ( .A1(n10297), .A2(n10296), .ZN(n10300) );
  INV_X1 U11399 ( .A(n10298), .ZN(n10299) );
  NAND2_X1 U11400 ( .A1(n10300), .A2(n10299), .ZN(n10302) );
  AOI21_X1 U11401 ( .B1(n10319), .B2(n10302), .A(n10301), .ZN(n10303) );
  OAI21_X1 U11402 ( .B1(n10305), .B2(n10304), .A(n10303), .ZN(n10306) );
  INV_X1 U11403 ( .A(n10306), .ZN(n10308) );
  NAND3_X1 U11404 ( .A1(n10309), .A2(n10308), .A3(n10307), .ZN(P1_U3245) );
  AOI22_X1 U11405 ( .A1(n10312), .A2(P1_ADDR_REG_5__SCAN_IN), .B1(n10311), 
        .B2(n10310), .ZN(n10325) );
  AOI211_X1 U11406 ( .C1(n10316), .C2(n10315), .A(n10314), .B(n10313), .ZN(
        n10317) );
  INV_X1 U11407 ( .A(n10317), .ZN(n10323) );
  OAI211_X1 U11408 ( .C1(n10321), .C2(n10320), .A(n10319), .B(n10318), .ZN(
        n10322) );
  NAND4_X1 U11409 ( .A1(n10325), .A2(n10324), .A3(n10323), .A4(n10322), .ZN(
        P1_U3246) );
  XNOR2_X1 U11410 ( .A(n10326), .B(n10336), .ZN(n10413) );
  INV_X1 U11411 ( .A(n10413), .ZN(n10333) );
  NOR2_X1 U11412 ( .A1(n10327), .A2(n10415), .ZN(n10328) );
  OR2_X1 U11413 ( .A1(n10329), .A2(n10328), .ZN(n10417) );
  INV_X1 U11414 ( .A(n10417), .ZN(n10330) );
  AOI22_X1 U11415 ( .A1(n10333), .A2(n10332), .B1(n10331), .B2(n10330), .ZN(
        n10352) );
  NAND2_X1 U11416 ( .A1(n10335), .A2(n10334), .ZN(n10337) );
  XNOR2_X1 U11417 ( .A(n10337), .B(n10336), .ZN(n10344) );
  OAI22_X1 U11418 ( .A1(n10341), .A2(n10340), .B1(n10339), .B2(n10338), .ZN(
        n10342) );
  AOI21_X1 U11419 ( .B1(n10344), .B2(n10343), .A(n10342), .ZN(n10420) );
  OAI21_X1 U11420 ( .B1(n10413), .B2(n7093), .A(n10420), .ZN(n10350) );
  AOI22_X1 U11421 ( .A1(n10048), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n10346), 
        .B2(n10345), .ZN(n10347) );
  OAI21_X1 U11422 ( .B1(n10415), .B2(n10256), .A(n10347), .ZN(n10348) );
  AOI21_X1 U11423 ( .B1(n10350), .B2(n10349), .A(n10348), .ZN(n10351) );
  NAND2_X1 U11424 ( .A1(n10352), .A2(n10351), .ZN(P1_U3282) );
  INV_X1 U11425 ( .A(n10353), .ZN(n10355) );
  AND2_X1 U11426 ( .A1(n10355), .A2(n10354), .ZN(n10365) );
  INV_X1 U11427 ( .A(n10365), .ZN(n10362) );
  AND2_X1 U11428 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10362), .ZN(P1_U3292) );
  AND2_X1 U11429 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10362), .ZN(P1_U3293) );
  AND2_X1 U11430 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10362), .ZN(P1_U3294) );
  NOR2_X1 U11431 ( .A1(n10365), .A2(n10356), .ZN(P1_U3295) );
  NOR2_X1 U11432 ( .A1(n10365), .A2(n10357), .ZN(P1_U3296) );
  AND2_X1 U11433 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10362), .ZN(P1_U3297) );
  AND2_X1 U11434 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10362), .ZN(P1_U3298) );
  AND2_X1 U11435 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10362), .ZN(P1_U3299) );
  AND2_X1 U11436 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10362), .ZN(P1_U3300) );
  NOR2_X1 U11437 ( .A1(n10365), .A2(n10358), .ZN(P1_U3301) );
  AND2_X1 U11438 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10362), .ZN(P1_U3302) );
  AND2_X1 U11439 ( .A1(n10362), .A2(P1_D_REG_20__SCAN_IN), .ZN(P1_U3303) );
  AND2_X1 U11440 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10362), .ZN(P1_U3304) );
  AND2_X1 U11441 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10362), .ZN(P1_U3305) );
  AND2_X1 U11442 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10362), .ZN(P1_U3306) );
  AND2_X1 U11443 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10362), .ZN(P1_U3307) );
  AND2_X1 U11444 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10362), .ZN(P1_U3308) );
  NOR2_X1 U11445 ( .A1(n10365), .A2(n10359), .ZN(P1_U3309) );
  AND2_X1 U11446 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10362), .ZN(P1_U3310) );
  AND2_X1 U11447 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10362), .ZN(P1_U3311) );
  NOR2_X1 U11448 ( .A1(n10365), .A2(n10360), .ZN(P1_U3312) );
  AND2_X1 U11449 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10362), .ZN(P1_U3313) );
  AND2_X1 U11450 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10362), .ZN(P1_U3314) );
  AND2_X1 U11451 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10362), .ZN(P1_U3315) );
  AND2_X1 U11452 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10362), .ZN(P1_U3316) );
  AND2_X1 U11453 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10362), .ZN(P1_U3317) );
  NOR2_X1 U11454 ( .A1(n10365), .A2(n10361), .ZN(P1_U3318) );
  AND2_X1 U11455 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10362), .ZN(P1_U3319) );
  NOR2_X1 U11456 ( .A1(n10365), .A2(n10363), .ZN(P1_U3320) );
  NOR2_X1 U11457 ( .A1(n10365), .A2(n10364), .ZN(P1_U3321) );
  OAI211_X1 U11458 ( .C1(n10369), .C2(n10368), .A(n10367), .B(n10366), .ZN(
        n10370) );
  NOR2_X1 U11459 ( .A1(n10371), .A2(n10370), .ZN(n10425) );
  INV_X1 U11460 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10372) );
  AOI22_X1 U11461 ( .A1(n10424), .A2(n10425), .B1(n10372), .B2(n10422), .ZN(
        P1_U3457) );
  OAI22_X1 U11462 ( .A1(n10374), .A2(n10416), .B1(n10373), .B2(n10414), .ZN(
        n10376) );
  AOI211_X1 U11463 ( .C1(n10410), .C2(n10377), .A(n10376), .B(n10375), .ZN(
        n10426) );
  INV_X1 U11464 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10378) );
  AOI22_X1 U11465 ( .A1(n10424), .A2(n10426), .B1(n10378), .B2(n10422), .ZN(
        P1_U3463) );
  INV_X1 U11466 ( .A(n10379), .ZN(n10382) );
  AOI211_X1 U11467 ( .C1(n10410), .C2(n10382), .A(n10381), .B(n10380), .ZN(
        n10427) );
  AOI22_X1 U11468 ( .A1(n10424), .A2(n10427), .B1(n10383), .B2(n10422), .ZN(
        P1_U3466) );
  NOR2_X1 U11469 ( .A1(n10384), .A2(n10412), .ZN(n10387) );
  NOR4_X1 U11470 ( .A1(n10388), .A2(n10387), .A3(n10386), .A4(n10385), .ZN(
        n10429) );
  INV_X1 U11471 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10389) );
  AOI22_X1 U11472 ( .A1(n10424), .A2(n10429), .B1(n10389), .B2(n10422), .ZN(
        P1_U3469) );
  OAI21_X1 U11473 ( .B1(n10391), .B2(n10414), .A(n10390), .ZN(n10393) );
  AOI211_X1 U11474 ( .C1(n10401), .C2(n10394), .A(n10393), .B(n10392), .ZN(
        n10431) );
  AOI22_X1 U11475 ( .A1(n10424), .A2(n10431), .B1(n10395), .B2(n10422), .ZN(
        P1_U3472) );
  OAI211_X1 U11476 ( .C1(n10416), .C2(n10398), .A(n10397), .B(n10396), .ZN(
        n10399) );
  AOI21_X1 U11477 ( .B1(n10401), .B2(n10400), .A(n10399), .ZN(n10433) );
  INV_X1 U11478 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10402) );
  AOI22_X1 U11479 ( .A1(n10424), .A2(n10433), .B1(n10402), .B2(n10422), .ZN(
        P1_U3475) );
  INV_X1 U11480 ( .A(n10403), .ZN(n10409) );
  INV_X1 U11481 ( .A(n10404), .ZN(n10405) );
  OAI22_X1 U11482 ( .A1(n10406), .A2(n10416), .B1(n10405), .B2(n10414), .ZN(
        n10408) );
  AOI211_X1 U11483 ( .C1(n10410), .C2(n10409), .A(n10408), .B(n10407), .ZN(
        n10435) );
  INV_X1 U11484 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10411) );
  AOI22_X1 U11485 ( .A1(n10424), .A2(n10435), .B1(n10411), .B2(n10422), .ZN(
        P1_U3478) );
  OR2_X1 U11486 ( .A1(n10413), .A2(n10412), .ZN(n10421) );
  OAI22_X1 U11487 ( .A1(n10417), .A2(n10416), .B1(n10415), .B2(n10414), .ZN(
        n10418) );
  INV_X1 U11488 ( .A(n10418), .ZN(n10419) );
  AND3_X1 U11489 ( .A1(n10421), .A2(n10420), .A3(n10419), .ZN(n10437) );
  AOI22_X1 U11490 ( .A1(n10424), .A2(n10437), .B1(n10423), .B2(n10422), .ZN(
        P1_U3481) );
  AOI22_X1 U11491 ( .A1(n10438), .A2(n10425), .B1(n6857), .B2(n10436), .ZN(
        P1_U3524) );
  AOI22_X1 U11492 ( .A1(n10438), .A2(n10426), .B1(n6861), .B2(n10436), .ZN(
        P1_U3526) );
  AOI22_X1 U11493 ( .A1(n10438), .A2(n10427), .B1(n6863), .B2(n10436), .ZN(
        P1_U3527) );
  AOI22_X1 U11494 ( .A1(n10438), .A2(n10429), .B1(n10428), .B2(n10436), .ZN(
        P1_U3528) );
  AOI22_X1 U11495 ( .A1(n10438), .A2(n10431), .B1(n10430), .B2(n10436), .ZN(
        P1_U3529) );
  AOI22_X1 U11496 ( .A1(n10438), .A2(n10433), .B1(n10432), .B2(n10436), .ZN(
        P1_U3530) );
  AOI22_X1 U11497 ( .A1(n10438), .A2(n10435), .B1(n10434), .B2(n10436), .ZN(
        P1_U3531) );
  AOI22_X1 U11498 ( .A1(n10438), .A2(n10437), .B1(n6867), .B2(n10436), .ZN(
        P1_U3532) );
  AOI22_X1 U11499 ( .A1(n10440), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10439), .ZN(n10449) );
  AOI22_X1 U11500 ( .A1(n10441), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10448) );
  NOR2_X1 U11501 ( .A1(n10442), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n10446) );
  OAI21_X1 U11502 ( .B1(P2_REG1_REG_0__SCAN_IN), .B2(n10444), .A(n10443), .ZN(
        n10445) );
  OAI21_X1 U11503 ( .B1(n10446), .B2(n10445), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n10447) );
  OAI211_X1 U11504 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n10449), .A(n10448), .B(
        n10447), .ZN(P2_U3245) );
  NOR2_X1 U11505 ( .A1(n10451), .A2(n10450), .ZN(n10460) );
  AND2_X1 U11506 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10462), .ZN(P2_U3297) );
  AND2_X1 U11507 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10462), .ZN(P2_U3298) );
  AND2_X1 U11508 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10462), .ZN(P2_U3299) );
  AND2_X1 U11509 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10462), .ZN(P2_U3300) );
  AND2_X1 U11510 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10462), .ZN(P2_U3301) );
  AND2_X1 U11511 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10462), .ZN(P2_U3302) );
  AND2_X1 U11512 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10462), .ZN(P2_U3303) );
  NOR2_X1 U11513 ( .A1(n10460), .A2(n10452), .ZN(P2_U3304) );
  NOR2_X1 U11514 ( .A1(n10460), .A2(n10453), .ZN(P2_U3305) );
  AND2_X1 U11515 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10462), .ZN(P2_U3306) );
  NOR2_X1 U11516 ( .A1(n10460), .A2(n10454), .ZN(P2_U3307) );
  AND2_X1 U11517 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10462), .ZN(P2_U3308) );
  AND2_X1 U11518 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10462), .ZN(P2_U3309) );
  AND2_X1 U11519 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10462), .ZN(P2_U3310) );
  AND2_X1 U11520 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10462), .ZN(P2_U3311) );
  AND2_X1 U11521 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10462), .ZN(P2_U3312) );
  NOR2_X1 U11522 ( .A1(n10460), .A2(n10455), .ZN(P2_U3313) );
  NOR2_X1 U11523 ( .A1(n10460), .A2(n10456), .ZN(P2_U3314) );
  AND2_X1 U11524 ( .A1(n10462), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3315) );
  AND2_X1 U11525 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10462), .ZN(P2_U3316) );
  NOR2_X1 U11526 ( .A1(n10460), .A2(n10457), .ZN(P2_U3317) );
  AND2_X1 U11527 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10462), .ZN(P2_U3318) );
  AND2_X1 U11528 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10462), .ZN(P2_U3319) );
  AND2_X1 U11529 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10462), .ZN(P2_U3320) );
  AND2_X1 U11530 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10462), .ZN(P2_U3321) );
  AND2_X1 U11531 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10462), .ZN(P2_U3322) );
  AND2_X1 U11532 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10462), .ZN(P2_U3323) );
  AND2_X1 U11533 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10462), .ZN(P2_U3324) );
  AND2_X1 U11534 ( .A1(n10462), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3325) );
  AND2_X1 U11535 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10462), .ZN(P2_U3326) );
  OAI22_X1 U11536 ( .A1(P2_D_REG_0__SCAN_IN), .A2(n10460), .B1(n10459), .B2(
        n10458), .ZN(n10461) );
  INV_X1 U11537 ( .A(n10461), .ZN(P2_U3437) );
  AOI22_X1 U11538 ( .A1(n10465), .A2(n10464), .B1(n10463), .B2(n10462), .ZN(
        P2_U3438) );
  AOI22_X1 U11539 ( .A1(n10468), .A2(n10524), .B1(n10467), .B2(n10466), .ZN(
        n10469) );
  AND2_X1 U11540 ( .A1(n10470), .A2(n10469), .ZN(n10529) );
  AOI22_X1 U11541 ( .A1(n10528), .A2(n10529), .B1(n5135), .B2(n10526), .ZN(
        P2_U3451) );
  NOR3_X1 U11542 ( .A1(n10472), .A2(n10471), .A3(n10520), .ZN(n10473) );
  AOI21_X1 U11543 ( .B1(n10475), .B2(n10474), .A(n10473), .ZN(n10476) );
  OAI211_X1 U11544 ( .C1(n10479), .C2(n10478), .A(n10477), .B(n10476), .ZN(
        n10480) );
  INV_X1 U11545 ( .A(n10480), .ZN(n10530) );
  AOI22_X1 U11546 ( .A1(n10528), .A2(n10530), .B1(n5164), .B2(n10526), .ZN(
        P2_U3454) );
  INV_X1 U11547 ( .A(n10481), .ZN(n10486) );
  OAI22_X1 U11548 ( .A1(n10483), .A2(n10520), .B1(n10482), .B2(n10518), .ZN(
        n10485) );
  AOI211_X1 U11549 ( .C1(n10524), .C2(n10486), .A(n10485), .B(n10484), .ZN(
        n10531) );
  INV_X1 U11550 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10487) );
  AOI22_X1 U11551 ( .A1(n10528), .A2(n10531), .B1(n10487), .B2(n10526), .ZN(
        P2_U3457) );
  OAI21_X1 U11552 ( .B1(n10489), .B2(n10518), .A(n10488), .ZN(n10490) );
  AOI21_X1 U11553 ( .B1(n10491), .B2(n10517), .A(n10490), .ZN(n10492) );
  AND2_X1 U11554 ( .A1(n10493), .A2(n10492), .ZN(n10532) );
  AOI22_X1 U11555 ( .A1(n10528), .A2(n10532), .B1(n5190), .B2(n10526), .ZN(
        P2_U3460) );
  OAI22_X1 U11556 ( .A1(n10495), .A2(n10520), .B1(n10494), .B2(n10518), .ZN(
        n10497) );
  AOI211_X1 U11557 ( .C1(n10524), .C2(n10498), .A(n10497), .B(n10496), .ZN(
        n10534) );
  AOI22_X1 U11558 ( .A1(n10528), .A2(n10534), .B1(n5223), .B2(n10526), .ZN(
        P2_U3463) );
  OAI211_X1 U11559 ( .C1(n10501), .C2(n10518), .A(n10500), .B(n10499), .ZN(
        n10502) );
  AOI21_X1 U11560 ( .B1(n10503), .B2(n10524), .A(n10502), .ZN(n10535) );
  AOI22_X1 U11561 ( .A1(n10528), .A2(n10535), .B1(n5266), .B2(n10526), .ZN(
        P2_U3469) );
  INV_X1 U11562 ( .A(n10504), .ZN(n10510) );
  INV_X1 U11563 ( .A(n10505), .ZN(n10506) );
  OAI22_X1 U11564 ( .A1(n10507), .A2(n10520), .B1(n10506), .B2(n10518), .ZN(
        n10509) );
  AOI211_X1 U11565 ( .C1(n10517), .C2(n10510), .A(n10509), .B(n10508), .ZN(
        n10537) );
  AOI22_X1 U11566 ( .A1(n10528), .A2(n10537), .B1(n5314), .B2(n10526), .ZN(
        P2_U3475) );
  INV_X1 U11567 ( .A(n10511), .ZN(n10516) );
  OAI22_X1 U11568 ( .A1(n10513), .A2(n10520), .B1(n10512), .B2(n10518), .ZN(
        n10515) );
  AOI211_X1 U11569 ( .C1(n10517), .C2(n10516), .A(n10515), .B(n10514), .ZN(
        n10538) );
  AOI22_X1 U11570 ( .A1(n10528), .A2(n10538), .B1(n5361), .B2(n10526), .ZN(
        P2_U3481) );
  OAI22_X1 U11571 ( .A1(n10521), .A2(n10520), .B1(n10519), .B2(n10518), .ZN(
        n10523) );
  AOI211_X1 U11572 ( .C1(n10525), .C2(n10524), .A(n10523), .B(n10522), .ZN(
        n10540) );
  INV_X1 U11573 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10527) );
  AOI22_X1 U11574 ( .A1(n10528), .A2(n10540), .B1(n10527), .B2(n10526), .ZN(
        P2_U3487) );
  AOI22_X1 U11575 ( .A1(n10541), .A2(n10529), .B1(n5136), .B2(n10539), .ZN(
        P2_U3520) );
  AOI22_X1 U11576 ( .A1(n10541), .A2(n10530), .B1(n7705), .B2(n10539), .ZN(
        P2_U3521) );
  AOI22_X1 U11577 ( .A1(n10541), .A2(n10531), .B1(n7703), .B2(n10539), .ZN(
        P2_U3522) );
  AOI22_X1 U11578 ( .A1(n10541), .A2(n10532), .B1(n7702), .B2(n10539), .ZN(
        P2_U3523) );
  AOI22_X1 U11579 ( .A1(n10541), .A2(n10534), .B1(n10533), .B2(n10539), .ZN(
        P2_U3524) );
  AOI22_X1 U11580 ( .A1(n10541), .A2(n10535), .B1(n7713), .B2(n10539), .ZN(
        P2_U3526) );
  AOI22_X1 U11581 ( .A1(n10541), .A2(n10537), .B1(n10536), .B2(n10539), .ZN(
        P2_U3528) );
  AOI22_X1 U11582 ( .A1(n10541), .A2(n10538), .B1(n7699), .B2(n10539), .ZN(
        P2_U3530) );
  AOI22_X1 U11583 ( .A1(n10541), .A2(n10540), .B1(n7719), .B2(n10539), .ZN(
        P2_U3532) );
  INV_X1 U11584 ( .A(n10542), .ZN(n10543) );
  NAND2_X1 U11585 ( .A1(n10544), .A2(n10543), .ZN(n10545) );
  XNOR2_X1 U11586 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10545), .ZN(ADD_1071_U5)
         );
  XOR2_X1 U11587 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11588 ( .B1(n10548), .B2(n10547), .A(n10546), .ZN(ADD_1071_U56) );
  OAI21_X1 U11589 ( .B1(n10551), .B2(n10550), .A(n10549), .ZN(ADD_1071_U57) );
  OAI21_X1 U11590 ( .B1(n10554), .B2(n10553), .A(n10552), .ZN(ADD_1071_U58) );
  OAI21_X1 U11591 ( .B1(n10557), .B2(n10556), .A(n10555), .ZN(ADD_1071_U59) );
  OAI21_X1 U11592 ( .B1(n10560), .B2(n10559), .A(n10558), .ZN(ADD_1071_U60) );
  OAI21_X1 U11593 ( .B1(n10563), .B2(n10562), .A(n10561), .ZN(ADD_1071_U61) );
  AOI21_X1 U11594 ( .B1(n10566), .B2(n10565), .A(n10564), .ZN(ADD_1071_U62) );
  AOI21_X1 U11595 ( .B1(n10569), .B2(n10568), .A(n10567), .ZN(ADD_1071_U63) );
  XOR2_X1 U11596 ( .A(n10570), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11597 ( .A1(n10572), .A2(n10571), .ZN(n10573) );
  XOR2_X1 U11598 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10573), .Z(ADD_1071_U51) );
  OAI21_X1 U11599 ( .B1(n10576), .B2(n10575), .A(n10574), .ZN(n10577) );
  XNOR2_X1 U11600 ( .A(n10577), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11601 ( .B1(n10580), .B2(n10579), .A(n10578), .ZN(ADD_1071_U47) );
  AOI21_X1 U11602 ( .B1(n10583), .B2(n10582), .A(n10581), .ZN(ADD_1071_U48) );
  XOR2_X1 U11603 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10584), .Z(ADD_1071_U49) );
  XOR2_X1 U11604 ( .A(n10586), .B(n10585), .Z(ADD_1071_U54) );
  XOR2_X1 U11605 ( .A(n10588), .B(n10587), .Z(ADD_1071_U53) );
  XNOR2_X1 U11606 ( .A(n10590), .B(n10589), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U5088 ( .A(n9234), .Z(n10593) );
  OAI21_X1 U11607 ( .B1(n5808), .B2(n5807), .A(n9537), .ZN(n9234) );
endmodule

