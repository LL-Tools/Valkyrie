

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, 
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, 
        keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, 
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, 
        keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, 
        keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, 
        keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, 
        keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, 
        keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, 
        keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, 
        keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, 
        keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941;

  AOI211_X1 U2364 ( .C1(n2998), .C2(n2530), .A(n4838), .B(n2997), .ZN(n2999)
         );
  NAND2_X1 U2365 ( .A1(n2281), .A2(n2280), .ZN(n4570) );
  CLKBUF_X1 U2366 ( .A(n3941), .Z(n2127) );
  NAND2_X1 U2367 ( .A1(n2580), .A2(n2579), .ZN(n3380) );
  INV_X1 U2368 ( .A(n3152), .ZN(n3218) );
  CLKBUF_X2 U2369 ( .A(n3026), .Z(n3611) );
  CLKBUF_X2 U2370 ( .A(n2469), .Z(n2789) );
  INV_X1 U2371 ( .A(n3611), .ZN(n3554) );
  OR2_X1 U2372 ( .A1(n2880), .A2(n2261), .ZN(n2260) );
  OAI21_X1 U2373 ( .B1(n2748), .B2(n2747), .A(IR_REG_31__SCAN_IN), .ZN(n2749)
         );
  BUF_X1 U2374 ( .A(n2496), .Z(n2941) );
  MUX2_X1 U2375 ( .A(n3946), .B(n3945), .S(n3944), .Z(n3947) );
  OR2_X1 U2376 ( .A1(n2780), .A2(n2923), .ZN(n2815) );
  XNOR2_X1 U2377 ( .A(n2751), .B(IR_REG_22__SCAN_IN), .ZN(n3950) );
  OR2_X1 U2378 ( .A1(n3053), .A2(n3048), .ZN(n3801) );
  NOR2_X1 U2379 ( .A1(n2527), .A2(n2526), .ZN(n4779) );
  AND4_X1 U2380 ( .A1(n2331), .A2(n2485), .A3(n2443), .A4(n2444), .ZN(n2122)
         );
  NOR2_X2 U2381 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2440)
         );
  XNOR2_X2 U2382 ( .A(n2841), .B(n2869), .ZN(n2990) );
  AND2_X2 U2383 ( .A1(n2246), .A2(n2150), .ZN(n2841) );
  NAND2_X2 U2384 ( .A1(n3150), .A2(n3149), .ZN(n3207) );
  NAND2_X2 U2385 ( .A1(n3089), .A2(n3038), .ZN(n3150) );
  OAI21_X2 U2386 ( .B1(n3732), .B2(n3735), .A(n3733), .ZN(n3634) );
  OAI21_X2 U2387 ( .B1(n2135), .B2(n3507), .A(n3506), .ZN(n3732) );
  NAND2_X2 U2388 ( .A1(n2304), .A2(IR_REG_31__SCAN_IN), .ZN(n2856) );
  XNOR2_X2 U2389 ( .A(n2890), .B(n4883), .ZN(n4825) );
  OR2_X1 U2390 ( .A1(n4127), .A2(n2709), .ZN(n2311) );
  NAND2_X1 U2391 ( .A1(n2893), .A2(n4881), .ZN(n2895) );
  XNOR2_X1 U2392 ( .A(n2887), .B(n4886), .ZN(n4803) );
  NAND4_X1 U2393 ( .A1(n2483), .A2(n2482), .A3(n2481), .A4(n2480), .ZN(n3226)
         );
  INV_X1 U2394 ( .A(n2126), .ZN(n2475) );
  NAND2_X1 U2395 ( .A1(n2311), .A2(n2330), .ZN(n4110) );
  AOI21_X1 U2396 ( .B1(n2895), .B2(REG2_REG_16__SCAN_IN), .A(n2253), .ZN(n2251) );
  AND2_X1 U2397 ( .A1(n2353), .A2(n2350), .ZN(n4479) );
  AOI21_X2 U2398 ( .B1(n4533), .B2(n4540), .A(n2667), .ZN(n4512) );
  NAND2_X1 U2399 ( .A1(n3918), .A2(n3903), .ZN(n4596) );
  NAND2_X1 U2400 ( .A1(n4803), .A2(REG2_REG_12__SCAN_IN), .ZN(n4802) );
  NAND2_X1 U2401 ( .A1(n2568), .A2(n2567), .ZN(n3346) );
  AND2_X1 U2402 ( .A1(n3810), .A2(n3869), .ZN(n4066) );
  OR2_X1 U2403 ( .A1(n4098), .A2(n4077), .ZN(n3810) );
  NAND3_X1 U2404 ( .A1(n2206), .A2(n2405), .A3(n2138), .ZN(n3362) );
  OAI21_X1 U2405 ( .B1(n3111), .B2(n4395), .A(n2215), .ZN(n3232) );
  OAI21_X1 U2406 ( .B1(n3135), .B2(n3134), .A(n3847), .ZN(n3122) );
  NAND2_X1 U2407 ( .A1(n2237), .A2(n2154), .ZN(n2236) );
  NAND2_X2 U2408 ( .A1(n3077), .A2(n4592), .ZN(n4585) );
  NAND2_X1 U2409 ( .A1(n3979), .A2(n3978), .ZN(n3977) );
  INV_X1 U2410 ( .A(n3963), .ZN(n3059) );
  AND4_X1 U2411 ( .A1(n2542), .A2(n2541), .A3(n2540), .A4(n2539), .ZN(n3330)
         );
  INV_X2 U2412 ( .A(n2478), .ZN(n3758) );
  INV_X2 U2413 ( .A(n3597), .ZN(n2123) );
  AND4_X2 U2414 ( .A1(n2471), .A2(n2473), .A3(n2472), .A4(n2474), .ZN(n2478)
         );
  CLKBUF_X3 U2415 ( .A(n2495), .Z(n3803) );
  INV_X1 U2416 ( .A(n3084), .ZN(n2959) );
  NAND2_X2 U2417 ( .A1(n3084), .A2(n3054), .ZN(n3612) );
  NAND2_X1 U2418 ( .A1(n2807), .A2(IR_REG_31__SCAN_IN), .ZN(n2379) );
  NAND2_X1 U2419 ( .A1(n2973), .A2(n2972), .ZN(n2971) );
  XNOR2_X1 U2420 ( .A(n2813), .B(IR_REG_25__SCAN_IN), .ZN(n4774) );
  NAND2_X1 U2421 ( .A1(n2743), .A2(IR_REG_31__SCAN_IN), .ZN(n2745) );
  OAI21_X1 U2422 ( .B1(n2811), .B2(n2810), .A(IR_REG_31__SCAN_IN), .ZN(n2813)
         );
  NOR2_X2 U2423 ( .A1(n2570), .A2(n2569), .ZN(n2586) );
  OAI21_X1 U2424 ( .B1(n2856), .B2(n2782), .A(n2466), .ZN(n2468) );
  NAND2_X1 U2425 ( .A1(n2924), .A2(IR_REG_31__SCAN_IN), .ZN(n2451) );
  NAND2_X1 U2426 ( .A1(n2856), .A2(n4160), .ZN(n2466) );
  INV_X1 U2427 ( .A(n2839), .ZN(n2373) );
  NOR2_X1 U2428 ( .A1(n2747), .A2(n2410), .ZN(n2411) );
  AND2_X1 U2429 ( .A1(n2431), .A2(n2781), .ZN(n2303) );
  AND4_X1 U2430 ( .A1(n2809), .A2(n2806), .A3(n2750), .A4(n2812), .ZN(n2431)
         );
  NAND2_X1 U2431 ( .A1(n4160), .A2(IR_REG_27__SCAN_IN), .ZN(n2467) );
  NOR2_X1 U2432 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2446)
         );
  INV_X1 U2433 ( .A(IR_REG_20__SCAN_IN), .ZN(n2744) );
  NOR2_X1 U2434 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_3__SCAN_IN), .ZN(n2331)
         );
  NOR2_X1 U2435 ( .A1(IR_REG_2__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2443)
         );
  NOR2_X1 U2436 ( .A1(IR_REG_4__SCAN_IN), .A2(IR_REG_13__SCAN_IN), .ZN(n2444)
         );
  NOR2_X1 U2437 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2442)
         );
  NOR2_X1 U2438 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2441)
         );
  AOI21_X2 U2439 ( .B1(n3224), .B2(n3225), .A(n3025), .ZN(n3755) );
  BUF_X4 U2440 ( .A(n2123), .Z(n2124) );
  BUF_X4 U2441 ( .A(n3807), .Z(n2125) );
  BUF_X4 U2442 ( .A(n3807), .Z(n2126) );
  NAND2_X2 U2443 ( .A1(n2468), .A2(n2467), .ZN(n3807) );
  NOR2_X2 U2444 ( .A1(n2606), .A2(n4217), .ZN(n2617) );
  XNOR2_X1 U2445 ( .A(n2749), .B(IR_REG_21__SCAN_IN), .ZN(n3941) );
  OAI211_X2 U2446 ( .C1(IR_REG_31__SCAN_IN), .C2(IR_REG_1__SCAN_IN), .A(n2332), 
        .B(n2238), .ZN(n3965) );
  CLKBUF_X3 U2447 ( .A(n2504), .Z(n3806) );
  AOI21_X1 U2448 ( .B1(n2134), .B2(n2295), .A(n2175), .ZN(n2292) );
  OAI22_X1 U2449 ( .A1(n3615), .A2(n2478), .B1(n3021), .B2(n3151), .ZN(n3023)
         );
  NAND2_X1 U2450 ( .A1(n2454), .A2(n4772), .ZN(n2504) );
  NOR2_X1 U2451 ( .A1(n3990), .A2(n4407), .ZN(n2374) );
  AND2_X1 U2452 ( .A1(n2324), .A2(n2165), .ZN(n2322) );
  NAND2_X1 U2453 ( .A1(n4578), .A2(n3895), .ZN(n2766) );
  INV_X1 U2454 ( .A(n3612), .ZN(n3589) );
  AND2_X1 U2456 ( .A1(n2395), .A2(n2402), .ZN(n2392) );
  OAI21_X1 U2457 ( .B1(n3572), .B2(n2415), .A(n2413), .ZN(n3585) );
  AOI21_X1 U2458 ( .B1(n3577), .B2(n2417), .A(n2414), .ZN(n2413) );
  AND2_X1 U2459 ( .A1(n3024), .A2(n3023), .ZN(n3025) );
  AND2_X1 U2460 ( .A1(n3950), .A2(n2127), .ZN(n3046) );
  INV_X1 U2461 ( .A(n2789), .ZN(n2716) );
  OAI21_X1 U2462 ( .B1(n4780), .B2(REG2_REG_2__SCAN_IN), .A(n2211), .ZN(n2975)
         );
  NAND2_X1 U2463 ( .A1(n4780), .A2(REG2_REG_2__SCAN_IN), .ZN(n2211) );
  NAND2_X1 U2464 ( .A1(n4847), .A2(n2356), .ZN(n2900) );
  NAND2_X1 U2465 ( .A1(n4880), .A2(n4205), .ZN(n2356) );
  OAI21_X1 U2466 ( .B1(n4836), .B2(n2248), .A(n2247), .ZN(n4003) );
  NAND2_X1 U2467 ( .A1(n4853), .A2(n2378), .ZN(n2247) );
  NAND2_X1 U2468 ( .A1(n2249), .A2(n2378), .ZN(n2248) );
  NAND2_X1 U2469 ( .A1(n4880), .A2(n4663), .ZN(n2378) );
  NAND2_X1 U2470 ( .A1(n4059), .A2(n2789), .ZN(n2740) );
  NAND2_X1 U2471 ( .A1(n2164), .A2(n2128), .ZN(n2288) );
  NOR2_X1 U2472 ( .A1(n2308), .A2(n2158), .ZN(n2306) );
  NAND2_X1 U2473 ( .A1(n2276), .A2(n2272), .ZN(n3199) );
  INV_X1 U2474 ( .A(n2273), .ZN(n2272) );
  NAND2_X1 U2475 ( .A1(n3133), .A2(n2277), .ZN(n2276) );
  OAI21_X1 U2476 ( .B1(n2278), .B2(n2274), .A(n2163), .ZN(n2273) );
  NAND2_X1 U2477 ( .A1(n2297), .A2(n2300), .ZN(n2294) );
  NAND2_X1 U2478 ( .A1(n2301), .A2(n2299), .ZN(n2298) );
  NAND2_X1 U2479 ( .A1(n4717), .A2(n4941), .ZN(n2212) );
  NOR2_X1 U2480 ( .A1(n2891), .A2(n2432), .ZN(n2225) );
  INV_X1 U2481 ( .A(n4812), .ZN(n2254) );
  INV_X1 U2482 ( .A(n2234), .ZN(n2231) );
  INV_X1 U2483 ( .A(n2227), .ZN(n2226) );
  INV_X1 U2484 ( .A(n2223), .ZN(n2222) );
  OAI21_X1 U2485 ( .B1(n3990), .B2(n4883), .A(n2228), .ZN(n2227) );
  INV_X1 U2486 ( .A(n2322), .ZN(n2321) );
  INV_X1 U2487 ( .A(n2330), .ZN(n2318) );
  INV_X1 U2488 ( .A(n2384), .ZN(n2383) );
  OAI21_X1 U2489 ( .B1(n2129), .B2(n2385), .A(n3655), .ZN(n2384) );
  NAND2_X1 U2490 ( .A1(n2373), .A2(REG1_REG_2__SCAN_IN), .ZN(n2372) );
  OAI21_X1 U2491 ( .B1(n2843), .B2(n2842), .A(n3977), .ZN(n2844) );
  INV_X1 U2492 ( .A(n3236), .ZN(n2267) );
  NAND2_X1 U2493 ( .A1(n3395), .A2(n2209), .ZN(n2887) );
  NAND2_X1 U2494 ( .A1(n2210), .A2(REG2_REG_11__SCAN_IN), .ZN(n2209) );
  INV_X1 U2495 ( .A(n4039), .ZN(n2338) );
  AOI21_X1 U2496 ( .B1(n2342), .B2(n2777), .A(n2341), .ZN(n2340) );
  INV_X1 U2497 ( .A(n3810), .ZN(n2341) );
  OAI21_X1 U2498 ( .B1(n4479), .B2(n4444), .A(n4443), .ZN(n4459) );
  NAND2_X1 U2499 ( .A1(n3376), .A2(n3817), .ZN(n3404) );
  AOI21_X1 U2500 ( .B1(n2322), .B2(n2320), .A(n2159), .ZN(n2319) );
  INV_X1 U2501 ( .A(n2327), .ZN(n2320) );
  NOR2_X1 U2502 ( .A1(n2321), .A2(n2318), .ZN(n2317) );
  NOR3_X1 U2503 ( .A1(n2321), .A2(n2318), .A3(n2314), .ZN(n2313) );
  INV_X1 U2504 ( .A(n2709), .ZN(n2314) );
  NAND2_X1 U2505 ( .A1(n4132), .A2(n3865), .ZN(n4116) );
  NOR2_X1 U2506 ( .A1(n3812), .A2(n2355), .ZN(n2354) );
  NAND2_X1 U2507 ( .A1(n4481), .A2(n3879), .ZN(n2300) );
  INV_X1 U2508 ( .A(n3332), .ZN(n3325) );
  INV_X1 U2509 ( .A(n4774), .ZN(n2817) );
  NOR2_X1 U2510 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2447)
         );
  INV_X1 U2511 ( .A(IR_REG_6__SCAN_IN), .ZN(n2439) );
  NOR2_X1 U2512 ( .A1(n2615), .A2(IR_REG_6__SCAN_IN), .ZN(n2565) );
  NAND2_X1 U2513 ( .A1(n2141), .A2(n2181), .ZN(n2407) );
  AND2_X1 U2514 ( .A1(n2181), .A2(n3208), .ZN(n2404) );
  INV_X1 U2515 ( .A(n2424), .ZN(n2423) );
  OAI21_X1 U2516 ( .B1(n3452), .B2(n2428), .A(n3451), .ZN(n2424) );
  NAND2_X1 U2517 ( .A1(n2427), .A2(n2426), .ZN(n2425) );
  INV_X1 U2518 ( .A(n2430), .ZN(n2427) );
  AND2_X1 U2519 ( .A1(n2423), .A2(n2135), .ZN(n2422) );
  INV_X1 U2520 ( .A(n3504), .ZN(n2421) );
  OR2_X1 U2521 ( .A1(n3061), .A2(n3949), .ZN(n3068) );
  OR2_X1 U2522 ( .A1(n3061), .A2(n3052), .ZN(n3053) );
  NAND2_X1 U2523 ( .A1(n2454), .A2(n2136), .ZN(n2474) );
  NAND2_X1 U2524 ( .A1(n2863), .A2(n2862), .ZN(n2977) );
  AND2_X1 U2525 ( .A1(n2243), .A2(REG1_REG_3__SCAN_IN), .ZN(n2240) );
  XNOR2_X1 U2526 ( .A(n2844), .B(n2874), .ZN(n2998) );
  AND2_X1 U2527 ( .A1(n2880), .A2(n4778), .ZN(n2268) );
  OAI211_X1 U2528 ( .C1(n2268), .C2(n3112), .A(n2267), .B(n2266), .ZN(n2269)
         );
  OR2_X1 U2529 ( .A1(n2268), .A2(REG2_REG_8__SCAN_IN), .ZN(n2266) );
  NAND2_X1 U2530 ( .A1(n3112), .A2(REG2_REG_8__SCAN_IN), .ZN(n2262) );
  OR2_X1 U2531 ( .A1(n2581), .A2(IR_REG_10__SCAN_IN), .ZN(n2582) );
  INV_X1 U2532 ( .A(IR_REG_11__SCAN_IN), .ZN(n2583) );
  NAND2_X1 U2533 ( .A1(n2217), .A2(n2216), .ZN(n2849) );
  NAND2_X1 U2534 ( .A1(n2210), .A2(REG1_REG_11__SCAN_IN), .ZN(n2216) );
  NAND2_X1 U2535 ( .A1(n3394), .A2(n2218), .ZN(n2217) );
  INV_X1 U2536 ( .A(n3393), .ZN(n2218) );
  NAND2_X1 U2537 ( .A1(n2192), .A2(n2155), .ZN(n2208) );
  NAND2_X1 U2538 ( .A1(n4490), .A2(n3880), .ZN(n2302) );
  NOR2_X1 U2539 ( .A1(n4560), .A2(n2666), .ZN(n2667) );
  CLKBUF_X1 U2540 ( .A(n2642), .Z(n2187) );
  AND2_X1 U2541 ( .A1(n2131), .A2(n3472), .ZN(n2370) );
  NAND2_X1 U2542 ( .A1(n2617), .A2(REG3_REG_14__SCAN_IN), .ZN(n2626) );
  NAND2_X1 U2543 ( .A1(n2586), .A2(REG3_REG_11__SCAN_IN), .ZN(n2598) );
  OAI21_X1 U2544 ( .B1(n3193), .B2(n2759), .A(n3839), .ZN(n3308) );
  AND2_X1 U2545 ( .A1(n3226), .A2(n3189), .ZN(n3174) );
  NAND2_X1 U2546 ( .A1(n2300), .A2(n2301), .ZN(n2295) );
  AND2_X1 U2547 ( .A1(n2674), .A2(n2673), .ZN(n4527) );
  AOI21_X1 U2548 ( .B1(n2133), .B2(n2285), .A(n2161), .ZN(n2280) );
  AOI21_X1 U2549 ( .B1(n2130), .B2(n2284), .A(n2162), .ZN(n2283) );
  INV_X1 U2550 ( .A(n2145), .ZN(n2284) );
  INV_X1 U2551 ( .A(n2130), .ZN(n2285) );
  NOR2_X1 U2552 ( .A1(n3263), .A2(n3332), .ZN(n2308) );
  NAND2_X1 U2553 ( .A1(n2544), .A2(n2309), .ZN(n2307) );
  NOR2_X1 U2554 ( .A1(n2310), .A2(n2556), .ZN(n2309) );
  INV_X1 U2555 ( .A(n2543), .ZN(n2310) );
  OAI22_X1 U2556 ( .A1(n3039), .A2(D_REG_0__SCAN_IN), .B1(n2818), .B2(n4773), 
        .ZN(n3075) );
  INV_X1 U2557 ( .A(IR_REG_27__SCAN_IN), .ZN(n2782) );
  INV_X1 U2558 ( .A(IR_REG_28__SCAN_IN), .ZN(n4160) );
  INV_X1 U2559 ( .A(IR_REG_12__SCAN_IN), .ZN(n2594) );
  INV_X1 U2560 ( .A(IR_REG_3__SCAN_IN), .ZN(n2509) );
  NAND2_X1 U2561 ( .A1(n2357), .A2(n2485), .ZN(n2332) );
  INV_X1 U2562 ( .A(IR_REG_1__SCAN_IN), .ZN(n2357) );
  NAND2_X1 U2563 ( .A1(n3165), .A2(n3166), .ZN(n3324) );
  NOR2_X1 U2564 ( .A1(n2390), .A2(n2402), .ZN(n2388) );
  NAND2_X1 U2565 ( .A1(n2392), .A2(n2390), .ZN(n2389) );
  INV_X1 U2566 ( .A(n2394), .ZN(n2393) );
  OAI21_X1 U2567 ( .B1(n2395), .B2(n2402), .A(n2401), .ZN(n2394) );
  INV_X1 U2568 ( .A(n2392), .ZN(n2391) );
  NAND2_X1 U2569 ( .A1(n3148), .A2(n3147), .ZN(n3149) );
  OR2_X1 U2570 ( .A1(n3068), .A2(n4783), .ZN(n3780) );
  INV_X1 U2571 ( .A(n4504), .ZN(n3879) );
  AND4_X1 U2572 ( .A1(n2603), .A2(n2602), .A3(n2601), .A4(n2600), .ZN(n3738)
         );
  OR2_X1 U2573 ( .A1(n3068), .A2(n3067), .ZN(n3769) );
  OAI21_X1 U2574 ( .B1(n3053), .B2(n4565), .A(n4592), .ZN(n3772) );
  NAND2_X1 U2575 ( .A1(n3066), .A2(STATE_REG_SCAN_IN), .ZN(n3778) );
  INV_X1 U2576 ( .A(n3330), .ZN(n3960) );
  NAND2_X1 U2577 ( .A1(n2845), .A2(n4778), .ZN(n2215) );
  XNOR2_X1 U2578 ( .A(n2846), .B(n2882), .ZN(n4799) );
  XNOR2_X1 U2579 ( .A(n2849), .B(n4886), .ZN(n4808) );
  NOR2_X1 U2580 ( .A1(n2900), .A2(n2899), .ZN(n4007) );
  NAND2_X1 U2581 ( .A1(n2900), .A2(n2899), .ZN(n2902) );
  XNOR2_X1 U2582 ( .A(n4003), .B(n2377), .ZN(n2857) );
  INV_X1 U2583 ( .A(n4002), .ZN(n2377) );
  AOI21_X1 U2584 ( .B1(ADDR_REG_18__SCAN_IN), .B2(n4851), .A(n2906), .ZN(n2361) );
  OR2_X1 U2585 ( .A1(n4791), .A2(n4784), .ZN(n4838) );
  AOI21_X1 U2586 ( .B1(n4003), .B2(n4002), .A(n2250), .ZN(n4006) );
  NOR2_X1 U2587 ( .A1(n2905), .A2(n4661), .ZN(n2250) );
  AOI21_X1 U2588 ( .B1(n4076), .B2(n4607), .A(n4075), .ZN(n4624) );
  OAI21_X1 U2589 ( .B1(n4110), .B2(n2717), .A(n2328), .ZN(n4086) );
  INV_X1 U2590 ( .A(n4708), .ZN(n4632) );
  INV_X1 U2591 ( .A(n4012), .ZN(n4004) );
  AND2_X1 U2592 ( .A1(n4539), .A2(n4924), .ZN(n4576) );
  OR2_X1 U2593 ( .A1(n4699), .A2(n4670), .ZN(n2196) );
  NAND2_X1 U2594 ( .A1(n2323), .A2(n2324), .ZN(n4067) );
  NAND2_X1 U2595 ( .A1(n4110), .A2(n2327), .ZN(n2323) );
  NAND2_X1 U2596 ( .A1(n2214), .A2(n2213), .ZN(n4717) );
  NOR2_X1 U2597 ( .A1(n4451), .A2(n4450), .ZN(n2213) );
  XNOR2_X1 U2598 ( .A(n2742), .B(n2741), .ZN(n4012) );
  NOR2_X1 U2599 ( .A1(n3236), .A2(n2265), .ZN(n2264) );
  NAND2_X1 U2600 ( .A1(n2374), .A2(n4883), .ZN(n2228) );
  OAI21_X1 U2601 ( .B1(n3990), .B2(n2182), .A(n2224), .ZN(n2223) );
  AOI21_X1 U2602 ( .B1(n2374), .B2(n2225), .A(n2184), .ZN(n2224) );
  AND2_X1 U2603 ( .A1(n4066), .A2(n4118), .ZN(n2186) );
  NAND2_X1 U2604 ( .A1(n2264), .A2(n4778), .ZN(n2261) );
  NAND2_X1 U2605 ( .A1(n2259), .A2(n2258), .ZN(n2257) );
  NAND2_X1 U2606 ( .A1(n2267), .A2(n4778), .ZN(n2258) );
  NAND2_X1 U2607 ( .A1(n2264), .A2(n3115), .ZN(n2259) );
  NOR2_X1 U2608 ( .A1(n2172), .A2(n2352), .ZN(n2351) );
  INV_X1 U2609 ( .A(n3925), .ZN(n2352) );
  INV_X1 U2610 ( .A(n3582), .ZN(n2414) );
  INV_X1 U2611 ( .A(n3577), .ZN(n2415) );
  OAI22_X1 U2612 ( .A1(n2123), .A2(n3292), .B1(n3615), .B2(n3246), .ZN(n3028)
         );
  NOR2_X1 U2613 ( .A1(n3529), .A2(n2435), .ZN(n3530) );
  NOR2_X1 U2614 ( .A1(n3681), .A2(n3680), .ZN(n3529) );
  OR3_X1 U2615 ( .A1(n2435), .A2(n3531), .A3(n3684), .ZN(n3542) );
  NAND2_X1 U2616 ( .A1(n2255), .A2(n2358), .ZN(n2890) );
  OR2_X1 U2617 ( .A1(n2889), .A2(REG2_REG_13__SCAN_IN), .ZN(n2358) );
  NAND2_X1 U2618 ( .A1(n4802), .A2(n2151), .ZN(n2255) );
  NAND2_X1 U2619 ( .A1(n2219), .A2(n2229), .ZN(n2852) );
  NOR2_X1 U2620 ( .A1(n2232), .A2(n2231), .ZN(n2230) );
  INV_X1 U2621 ( .A(n2853), .ZN(n2249) );
  NAND2_X1 U2622 ( .A1(n2528), .A2(n2275), .ZN(n2274) );
  INV_X1 U2623 ( .A(n2538), .ZN(n2275) );
  INV_X1 U2624 ( .A(n2529), .ZN(n2278) );
  NOR2_X1 U2625 ( .A1(n2278), .A2(n2538), .ZN(n2277) );
  NAND2_X1 U2626 ( .A1(n2188), .A2(n3825), .ZN(n3244) );
  NAND2_X1 U2627 ( .A1(n3246), .A2(n3760), .ZN(n3825) );
  INV_X1 U2628 ( .A(n3819), .ZN(n3822) );
  NAND2_X1 U2629 ( .A1(n3021), .A2(n3758), .ZN(n3820) );
  NAND2_X1 U2630 ( .A1(n2486), .A2(n2478), .ZN(n3824) );
  NOR2_X1 U2631 ( .A1(n4030), .A2(n4079), .ZN(n4017) );
  NAND2_X1 U2632 ( .A1(n4448), .A2(n4135), .ZN(n2330) );
  NOR2_X1 U2633 ( .A1(n4128), .A2(n2369), .ZN(n2368) );
  INV_X1 U2634 ( .A(n4462), .ZN(n4469) );
  INV_X1 U2635 ( .A(n2302), .ZN(n2299) );
  NAND2_X1 U2636 ( .A1(n2766), .A2(n3813), .ZN(n4517) );
  NOR2_X1 U2637 ( .A1(n4555), .A2(n4579), .ZN(n2366) );
  OR2_X1 U2638 ( .A1(n3052), .A2(n3063), .ZN(n3074) );
  INV_X1 U2639 ( .A(IR_REG_18__SCAN_IN), .ZN(n2664) );
  OR2_X1 U2640 ( .A1(n2652), .A2(IR_REG_17__SCAN_IN), .ZN(n2663) );
  OR2_X1 U2641 ( .A1(n2576), .A2(IR_REG_9__SCAN_IN), .ZN(n2581) );
  INV_X1 U2642 ( .A(n3609), .ZN(n2402) );
  INV_X1 U2643 ( .A(n2398), .ZN(n2390) );
  INV_X1 U2644 ( .A(n3765), .ZN(n2386) );
  NAND2_X1 U2645 ( .A1(n2396), .A2(n2160), .ZN(n2395) );
  NOR2_X1 U2646 ( .A1(n2132), .A2(n2399), .ZN(n2398) );
  INV_X1 U2647 ( .A(n2407), .ZN(n2406) );
  XNOR2_X1 U2648 ( .A(n3033), .B(n3589), .ZN(n3146) );
  NOR2_X1 U2649 ( .A1(n3017), .A2(n2964), .ZN(n3019) );
  AOI21_X1 U2650 ( .B1(n2383), .B2(n2385), .A(n2139), .ZN(n2381) );
  NAND2_X1 U2651 ( .A1(n2191), .A2(n2171), .ZN(n3572) );
  NAND2_X1 U2652 ( .A1(n3434), .A2(n3435), .ZN(n2428) );
  OR2_X1 U2653 ( .A1(n3424), .A2(n2430), .ZN(n2429) );
  INV_X1 U2654 ( .A(n3615), .ZN(n3602) );
  OR2_X1 U2655 ( .A1(n2971), .A2(n2245), .ZN(n2241) );
  NAND2_X1 U2656 ( .A1(n2971), .A2(n2242), .ZN(n2239) );
  NAND2_X1 U2657 ( .A1(n3983), .A2(n2873), .ZN(n2875) );
  NAND2_X1 U2658 ( .A1(n2376), .A2(n2375), .ZN(n2845) );
  NAND2_X1 U2659 ( .A1(n3004), .A2(REG1_REG_7__SCAN_IN), .ZN(n2375) );
  NAND2_X1 U2660 ( .A1(n2236), .A2(n2174), .ZN(n2376) );
  NAND2_X1 U2661 ( .A1(n4818), .A2(n2432), .ZN(n2221) );
  INV_X1 U2662 ( .A(n3993), .ZN(n2207) );
  XNOR2_X1 U2663 ( .A(n2852), .B(n2894), .ZN(n4837) );
  NOR2_X1 U2664 ( .A1(REG1_REG_16__SCAN_IN), .A2(n4837), .ZN(n4836) );
  AOI21_X1 U2665 ( .B1(n2343), .B2(n2340), .A(n2338), .ZN(n2337) );
  NAND2_X1 U2666 ( .A1(n2336), .A2(n2340), .ZN(n4040) );
  NAND2_X1 U2667 ( .A1(n4116), .A2(n2342), .ZN(n2336) );
  NAND2_X1 U2668 ( .A1(n2344), .A2(n2342), .ZN(n4071) );
  INV_X1 U2669 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3649) );
  NOR2_X2 U2670 ( .A1(n2642), .A2(n2437), .ZN(n2656) );
  INV_X1 U2671 ( .A(REG3_REG_15__SCAN_IN), .ZN(n3794) );
  NAND2_X1 U2672 ( .A1(n3381), .A2(n2370), .ZN(n3496) );
  INV_X1 U2673 ( .A(REG3_REG_13__SCAN_IN), .ZN(n4217) );
  INV_X1 U2674 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2597) );
  OR2_X2 U2675 ( .A1(n2598), .A2(n2597), .ZN(n2606) );
  NAND2_X1 U2676 ( .A1(n2760), .A2(n3844), .ZN(n3376) );
  INV_X1 U2677 ( .A(n2547), .ZN(n2202) );
  INV_X1 U2678 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2515) );
  INV_X1 U2679 ( .A(n3100), .ZN(n3105) );
  NAND2_X1 U2680 ( .A1(n3256), .A2(n3105), .ZN(n3143) );
  NOR2_X1 U2681 ( .A1(n3291), .A2(n3254), .ZN(n3256) );
  NAND2_X1 U2682 ( .A1(n2333), .A2(n3824), .ZN(n3279) );
  NAND2_X1 U2683 ( .A1(n2334), .A2(n3822), .ZN(n2333) );
  INV_X1 U2684 ( .A(n2753), .ZN(n2334) );
  AND2_X1 U2685 ( .A1(n3021), .A2(n3080), .ZN(n3293) );
  NOR2_X1 U2686 ( .A1(n4037), .A2(n4024), .ZN(n4023) );
  NAND2_X1 U2687 ( .A1(n2316), .A2(n2312), .ZN(n4032) );
  NOR2_X1 U2688 ( .A1(n2315), .A2(n2313), .ZN(n2312) );
  INV_X1 U2689 ( .A(n2319), .ZN(n2315) );
  NAND2_X1 U2690 ( .A1(n4087), .A2(n4077), .ZN(n4079) );
  AOI21_X1 U2691 ( .B1(n2325), .B2(n2328), .A(n2156), .ZN(n2324) );
  NOR2_X1 U2692 ( .A1(n2725), .A2(n2326), .ZN(n2325) );
  INV_X1 U2693 ( .A(n2717), .ZN(n2326) );
  NOR2_X1 U2694 ( .A1(n2725), .A2(n2329), .ZN(n2327) );
  AND2_X1 U2695 ( .A1(n4642), .A2(n2367), .ZN(n4087) );
  AND2_X1 U2696 ( .A1(n2142), .A2(n4099), .ZN(n2367) );
  NAND2_X1 U2697 ( .A1(n4642), .A2(n2142), .ZN(n4111) );
  NAND2_X1 U2698 ( .A1(n4642), .A2(n2368), .ZN(n4130) );
  NAND2_X1 U2699 ( .A1(n4642), .A2(n4449), .ZN(n4439) );
  AND2_X1 U2700 ( .A1(n4476), .A2(n4469), .ZN(n4642) );
  CLKBUF_X1 U2701 ( .A(n4436), .Z(n4457) );
  INV_X1 U2702 ( .A(n2172), .ZN(n2350) );
  AND2_X1 U2703 ( .A1(n2695), .A2(n2694), .ZN(n4483) );
  NOR2_X1 U2704 ( .A1(n2143), .A2(n4480), .ZN(n4476) );
  AND2_X1 U2705 ( .A1(n4571), .A2(n2364), .ZN(n4536) );
  NOR2_X1 U2706 ( .A1(n2365), .A2(n2666), .ZN(n2364) );
  INV_X1 U2707 ( .A(n2366), .ZN(n2365) );
  NAND2_X1 U2708 ( .A1(n4571), .A2(n2366), .ZN(n4553) );
  AND2_X1 U2709 ( .A1(n3884), .A2(n4518), .ZN(n4557) );
  NAND2_X1 U2710 ( .A1(n4571), .A2(n2825), .ZN(n4572) );
  NAND2_X1 U2711 ( .A1(n3381), .A2(n2131), .ZN(n3485) );
  AND2_X1 U2712 ( .A1(n3381), .A2(n3437), .ZN(n3410) );
  AND2_X1 U2713 ( .A1(n3067), .A2(n3046), .ZN(n4601) );
  NAND2_X1 U2714 ( .A1(n2348), .A2(n3838), .ZN(n3262) );
  NOR2_X1 U2715 ( .A1(n3200), .A2(n3201), .ZN(n3313) );
  NAND2_X1 U2716 ( .A1(n3256), .A2(n2146), .ZN(n3141) );
  NAND2_X1 U2717 ( .A1(n4502), .A2(n4894), .ZN(n4928) );
  NAND2_X1 U2718 ( .A1(n4773), .A2(n2816), .ZN(n3039) );
  NAND2_X1 U2719 ( .A1(n2960), .A2(n4877), .ZN(n3052) );
  NAND4_X1 U2720 ( .A1(n2448), .A2(n2445), .A3(n2303), .A4(n2122), .ZN(n2304)
         );
  NAND2_X1 U2721 ( .A1(n2750), .A2(n2806), .ZN(n2410) );
  INV_X1 U2722 ( .A(IR_REG_23__SCAN_IN), .ZN(n2820) );
  INV_X1 U2723 ( .A(IR_REG_19__SCAN_IN), .ZN(n2741) );
  OR2_X1 U2724 ( .A1(n2565), .A2(n2923), .ZN(n2553) );
  XNOR2_X1 U2725 ( .A(n2553), .B(IR_REG_7__SCAN_IN), .ZN(n3004) );
  NAND2_X1 U2726 ( .A1(n2525), .A2(n2524), .ZN(n2615) );
  AND2_X1 U2727 ( .A1(n2522), .A2(n2521), .ZN(n2525) );
  NOR2_X1 U2728 ( .A1(IR_REG_3__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2521)
         );
  NAND2_X1 U2729 ( .A1(n2408), .A2(n2407), .ZN(n3166) );
  AND4_X1 U2731 ( .A1(n2591), .A2(n2590), .A3(n2589), .A4(n2588), .ZN(n3457)
         );
  NAND2_X1 U2732 ( .A1(n2382), .A2(n3764), .ZN(n3654) );
  NAND2_X1 U2733 ( .A1(n3547), .A2(n2129), .ZN(n2382) );
  XNOR2_X1 U2734 ( .A(n3022), .B(n3024), .ZN(n3225) );
  OAI22_X1 U2735 ( .A1(n3019), .A2(n3018), .B1(n3612), .B2(n3017), .ZN(n3224)
         );
  NAND2_X1 U2736 ( .A1(n3721), .A2(n3725), .ZN(n3663) );
  INV_X1 U2737 ( .A(n3568), .ZN(n4480) );
  AND2_X1 U2738 ( .A1(n2687), .A2(n2686), .ZN(n4465) );
  INV_X1 U2739 ( .A(n3415), .ZN(n3443) );
  AOI21_X1 U2740 ( .B1(n2425), .B2(n2422), .A(n2421), .ZN(n2420) );
  NAND2_X1 U2741 ( .A1(n3572), .A2(n3571), .ZN(n3745) );
  NAND2_X1 U2742 ( .A1(n3547), .A2(n3546), .ZN(n3767) );
  NAND2_X1 U2743 ( .A1(n3208), .A2(n3207), .ZN(n2409) );
  INV_X1 U2744 ( .A(n3796), .ZN(n3759) );
  AOI21_X1 U2745 ( .B1(n3673), .B2(n3670), .A(n3671), .ZN(n3777) );
  INV_X1 U2746 ( .A(n3780), .ZN(n3798) );
  INV_X1 U2747 ( .A(n3778), .ZN(n3793) );
  INV_X1 U2748 ( .A(n3769), .ZN(n3791) );
  OR2_X1 U2749 ( .A1(n2124), .A2(n3056), .ZN(n3949) );
  NAND2_X1 U2750 ( .A1(n4080), .A2(n2789), .ZN(n2730) );
  INV_X1 U2751 ( .A(n4465), .ZN(n3957) );
  INV_X1 U2752 ( .A(n4483), .ZN(n3664) );
  NAND2_X1 U2753 ( .A1(n2680), .A2(n2679), .ZN(n4500) );
  INV_X1 U2754 ( .A(n4527), .ZN(n4481) );
  OAI211_X1 U2755 ( .C1(n4593), .C2(n2716), .A(n2629), .B(n2628), .ZN(n4580)
         );
  OAI211_X1 U2756 ( .C1(n3638), .C2(n2716), .A(n2621), .B(n2620), .ZN(n4602)
         );
  INV_X1 U2757 ( .A(n3457), .ZN(n3958) );
  OR2_X1 U2758 ( .A1(n2504), .A2(n2963), .ZN(n2483) );
  OAI21_X1 U2759 ( .B1(n3965), .B2(REG2_REG_1__SCAN_IN), .A(n2193), .ZN(n3973)
         );
  NAND2_X1 U2760 ( .A1(n3965), .A2(REG2_REG_1__SCAN_IN), .ZN(n2193) );
  NAND2_X1 U2761 ( .A1(n3970), .A2(n3969), .ZN(n3968) );
  NAND2_X1 U2762 ( .A1(n2989), .A2(n2194), .ZN(n3979) );
  INV_X1 U2763 ( .A(n2237), .ZN(n2997) );
  INV_X1 U2764 ( .A(n2236), .ZN(n3007) );
  XNOR2_X1 U2765 ( .A(n2845), .B(n4778), .ZN(n3111) );
  AND2_X1 U2766 ( .A1(n2263), .A2(n2262), .ZN(n3237) );
  INV_X1 U2767 ( .A(n2268), .ZN(n2263) );
  NAND2_X1 U2768 ( .A1(n4798), .A2(n2848), .ZN(n3394) );
  NAND2_X1 U2769 ( .A1(n2847), .A2(n2882), .ZN(n2848) );
  NAND2_X1 U2770 ( .A1(n4808), .A2(REG1_REG_12__SCAN_IN), .ZN(n4807) );
  NAND2_X1 U2771 ( .A1(n4802), .A2(n2888), .ZN(n4814) );
  NAND2_X1 U2772 ( .A1(n4830), .A2(REG1_REG_14__SCAN_IN), .ZN(n4829) );
  NAND2_X1 U2773 ( .A1(n4829), .A2(n2851), .ZN(n3989) );
  NAND2_X1 U2774 ( .A1(n2221), .A2(n2891), .ZN(n2851) );
  NAND2_X1 U2775 ( .A1(n4835), .A2(n4834), .ZN(n4833) );
  INV_X1 U2776 ( .A(n4848), .ZN(n2253) );
  NAND2_X1 U2777 ( .A1(n4833), .A2(n2895), .ZN(n4846) );
  NOR2_X1 U2778 ( .A1(n4854), .A2(n4853), .ZN(n4855) );
  INV_X1 U2779 ( .A(n4838), .ZN(n4852) );
  AND2_X1 U2780 ( .A1(n2719), .A2(n2734), .ZN(n4105) );
  NAND2_X1 U2781 ( .A1(n2296), .A2(n2301), .ZN(n4489) );
  NAND2_X1 U2782 ( .A1(n3381), .A2(n2137), .ZN(n4678) );
  NAND2_X1 U2783 ( .A1(n3409), .A2(n2145), .ZN(n2287) );
  AND2_X1 U2784 ( .A1(n2289), .A2(n2290), .ZN(n3484) );
  NAND2_X1 U2785 ( .A1(n3409), .A2(n2605), .ZN(n2289) );
  NAND2_X1 U2786 ( .A1(n2544), .A2(n2543), .ZN(n3312) );
  INV_X1 U2787 ( .A(n4588), .ZN(n4613) );
  NAND2_X1 U2788 ( .A1(n2279), .A2(n2529), .ZN(n3121) );
  OR2_X1 U2789 ( .A1(n3133), .A2(n2528), .ZN(n2279) );
  INV_X1 U2790 ( .A(n4592), .ZN(n4574) );
  XNOR2_X1 U2791 ( .A(n4023), .B(n4020), .ZN(n4693) );
  NAND2_X1 U2792 ( .A1(n2199), .A2(n2198), .ZN(n4708) );
  NOR2_X1 U2793 ( .A1(n4122), .A2(n4121), .ZN(n2198) );
  NAND2_X1 U2794 ( .A1(n4123), .A2(n4607), .ZN(n2199) );
  NAND2_X1 U2795 ( .A1(n2293), .A2(n2294), .ZN(n4475) );
  OR2_X1 U2796 ( .A1(n4512), .A2(n2295), .ZN(n2293) );
  NAND2_X1 U2797 ( .A1(n2282), .A2(n2283), .ZN(n4589) );
  OR2_X1 U2798 ( .A1(n3409), .A2(n2285), .ZN(n2282) );
  INV_X1 U2799 ( .A(n2307), .ZN(n2305) );
  NOR2_X1 U2800 ( .A1(n2449), .A2(IR_REG_29__SCAN_IN), .ZN(n2346) );
  NAND2_X1 U2801 ( .A1(n2452), .A2(IR_REG_31__SCAN_IN), .ZN(n2453) );
  INV_X1 U2802 ( .A(n2449), .ZN(n2345) );
  AND2_X1 U2803 ( .A1(n2854), .A2(STATE_REG_SCAN_IN), .ZN(n4877) );
  NOR2_X1 U2804 ( .A1(n2747), .A2(IR_REG_21__SCAN_IN), .ZN(n2412) );
  XNOR2_X1 U2805 ( .A(n2595), .B(n2594), .ZN(n4886) );
  XNOR2_X1 U2806 ( .A(n2566), .B(IR_REG_9__SCAN_IN), .ZN(n4777) );
  NAND2_X1 U2807 ( .A1(n2332), .A2(IR_REG_31__SCAN_IN), .ZN(n2270) );
  NAND2_X1 U2808 ( .A1(n2400), .A2(n3608), .ZN(U3211) );
  NAND2_X1 U2809 ( .A1(n2362), .A2(n2360), .ZN(U3258) );
  INV_X1 U2810 ( .A(n2904), .ZN(n2362) );
  AND2_X1 U2811 ( .A1(n2907), .A2(n2361), .ZN(n2360) );
  AOI21_X1 U2812 ( .B1(n4014), .B2(n2901), .A(n4013), .ZN(n4015) );
  AND2_X1 U2813 ( .A1(n4056), .A2(n4057), .ZN(n2271) );
  NAND2_X1 U2814 ( .A1(n2197), .A2(n2157), .ZN(U3547) );
  NAND2_X1 U2815 ( .A1(n4698), .A2(n4941), .ZN(n2197) );
  OR2_X1 U2816 ( .A1(n4061), .A2(n4675), .ZN(n2834) );
  OR2_X1 U2817 ( .A1(n4703), .A2(n4670), .ZN(n2185) );
  NAND2_X1 U2818 ( .A1(n2212), .A2(n2169), .ZN(n4640) );
  NAND2_X1 U2819 ( .A1(n4930), .A2(REG0_REG_29__SCAN_IN), .ZN(n2189) );
  OR2_X1 U2820 ( .A1(n4699), .A2(n4758), .ZN(n2200) );
  NAND2_X1 U2821 ( .A1(n4698), .A2(n4932), .ZN(n2190) );
  NAND2_X1 U2822 ( .A1(n2205), .A2(n4755), .ZN(n2204) );
  INV_X1 U2823 ( .A(n4707), .ZN(n2205) );
  OR2_X1 U2824 ( .A1(n3636), .A2(n3740), .ZN(n2128) );
  AND2_X1 U2825 ( .A1(n2386), .A2(n3546), .ZN(n2129) );
  AND2_X1 U2826 ( .A1(n2288), .A2(n2286), .ZN(n2130) );
  AND2_X1 U2827 ( .A1(n3454), .A2(n3437), .ZN(n2131) );
  INV_X1 U2828 ( .A(n3220), .ZN(n2363) );
  NOR2_X1 U2829 ( .A1(n3596), .A2(n3595), .ZN(n2132) );
  AND2_X1 U2830 ( .A1(n2283), .A2(n2149), .ZN(n2133) );
  AND2_X1 U2831 ( .A1(n2294), .A2(n2173), .ZN(n2134) );
  XOR2_X1 U2832 ( .A(n3453), .B(n3612), .Z(n2135) );
  AND2_X1 U2833 ( .A1(n4772), .A2(REG1_REG_1__SCAN_IN), .ZN(n2136) );
  AND2_X1 U2834 ( .A1(n2370), .A2(n2625), .ZN(n2137) );
  NAND2_X1 U2835 ( .A1(n3323), .A2(n3322), .ZN(n2138) );
  NOR2_X1 U2836 ( .A1(n3559), .A2(n3558), .ZN(n2139) );
  NAND2_X1 U2837 ( .A1(n2221), .A2(n4883), .ZN(n2140) );
  INV_X1 U2838 ( .A(n4448), .ZN(n3956) );
  AND2_X1 U2839 ( .A1(n2708), .A2(n2707), .ZN(n4448) );
  NAND2_X1 U2840 ( .A1(n3215), .A2(n2148), .ZN(n2141) );
  XNOR2_X1 U2841 ( .A(n2880), .B(n3115), .ZN(n3112) );
  AND2_X1 U2842 ( .A1(n2368), .A2(n4120), .ZN(n2142) );
  OR2_X1 U2843 ( .A1(n4503), .A2(n3879), .ZN(n2143) );
  INV_X1 U2844 ( .A(n2470), .ZN(n2613) );
  INV_X1 U2845 ( .A(IR_REG_25__SCAN_IN), .ZN(n2812) );
  AND2_X1 U2846 ( .A1(n3636), .A2(n3740), .ZN(n2144) );
  INV_X4 U2847 ( .A(n3151), .ZN(n3597) );
  INV_X1 U2848 ( .A(IR_REG_31__SCAN_IN), .ZN(n2923) );
  AND2_X1 U2849 ( .A1(n2128), .A2(n2605), .ZN(n2145) );
  AND2_X1 U2850 ( .A1(n2824), .A2(n3105), .ZN(n2146) );
  NAND2_X1 U2851 ( .A1(n2460), .A2(n2459), .ZN(n4547) );
  INV_X1 U2852 ( .A(n4547), .ZN(n4490) );
  AND3_X1 U2853 ( .A1(n2500), .A2(n2497), .A3(n2499), .ZN(n2147) );
  NAND2_X1 U2854 ( .A1(n3156), .A2(n3155), .ZN(n2148) );
  NAND2_X1 U2855 ( .A1(n2287), .A2(n2288), .ZN(n3490) );
  INV_X1 U2856 ( .A(IR_REG_5__SCAN_IN), .ZN(n2524) );
  OR2_X1 U2857 ( .A1(n4580), .A2(n4600), .ZN(n2149) );
  NAND2_X1 U2858 ( .A1(n2371), .A2(n2865), .ZN(n2150) );
  NOR2_X1 U2859 ( .A1(n2626), .A2(n3794), .ZN(n2201) );
  BUF_X1 U2860 ( .A(n2461), .Z(n2748) );
  AND2_X1 U2861 ( .A1(n2888), .A2(n2254), .ZN(n2151) );
  NAND2_X1 U2862 ( .A1(n3415), .A2(n3419), .ZN(n2152) );
  AND3_X1 U2863 ( .A1(n4160), .A2(n2782), .A3(n2781), .ZN(n2153) );
  NAND2_X1 U2864 ( .A1(n2844), .A2(n2874), .ZN(n2154) );
  OR2_X1 U2865 ( .A1(n4883), .A2(n2890), .ZN(n2155) );
  INV_X1 U2866 ( .A(n2417), .ZN(n2416) );
  NAND2_X1 U2867 ( .A1(n2418), .A2(n3571), .ZN(n2417) );
  AND2_X1 U2868 ( .A1(n4119), .A2(n4099), .ZN(n2156) );
  AND2_X1 U2869 ( .A1(n2196), .A2(n2195), .ZN(n2157) );
  INV_X1 U2870 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2840) );
  NOR2_X1 U2871 ( .A1(n3959), .A2(n3373), .ZN(n2158) );
  NOR2_X1 U2872 ( .A1(n2731), .A2(n4077), .ZN(n2159) );
  NAND2_X1 U2873 ( .A1(n2403), .A2(n3775), .ZN(n2160) );
  INV_X1 U2874 ( .A(n2329), .ZN(n2328) );
  NOR2_X1 U2875 ( .A1(n3781), .A2(n4120), .ZN(n2329) );
  NOR2_X1 U2876 ( .A1(n3692), .A2(n3795), .ZN(n2161) );
  INV_X1 U2877 ( .A(IR_REG_29__SCAN_IN), .ZN(n2450) );
  NOR2_X1 U2878 ( .A1(n4602), .A2(n3641), .ZN(n2162) );
  NAND2_X1 U2879 ( .A1(n3961), .A2(n3220), .ZN(n2163) );
  INV_X1 U2880 ( .A(n2343), .ZN(n2342) );
  NAND2_X1 U2881 ( .A1(n4066), .A2(n3871), .ZN(n2343) );
  OR2_X1 U2882 ( .A1(n2604), .A2(n2144), .ZN(n2164) );
  INV_X1 U2883 ( .A(IR_REG_21__SCAN_IN), .ZN(n2750) );
  NAND2_X1 U2884 ( .A1(n2675), .A2(n2298), .ZN(n2297) );
  OR2_X1 U2885 ( .A1(n4098), .A2(n3607), .ZN(n2165) );
  AND2_X1 U2886 ( .A1(REG3_REG_7__SCAN_IN), .A2(REG3_REG_8__SCAN_IN), .ZN(
        n2166) );
  AND2_X1 U2887 ( .A1(n2146), .A2(n2363), .ZN(n2167) );
  INV_X1 U2888 ( .A(IR_REG_26__SCAN_IN), .ZN(n2781) );
  AND2_X1 U2889 ( .A1(n2393), .A2(n2389), .ZN(n2168) );
  INV_X1 U2890 ( .A(n3813), .ZN(n2355) );
  OR2_X1 U2891 ( .A1(n4941), .A2(n4337), .ZN(n2169) );
  INV_X1 U2892 ( .A(n2132), .ZN(n2396) );
  INV_X1 U2893 ( .A(n3670), .ZN(n2399) );
  OAI21_X1 U2894 ( .B1(n4537), .B2(n2716), .A(n2662), .ZN(n4560) );
  AND2_X1 U2895 ( .A1(n4777), .A2(REG1_REG_9__SCAN_IN), .ZN(n2170) );
  AND2_X1 U2896 ( .A1(n4595), .A2(n3814), .ZN(n3903) );
  INV_X1 U2897 ( .A(n3903), .ZN(n2286) );
  OR2_X1 U2898 ( .A1(n3661), .A2(n3660), .ZN(n2171) );
  AND2_X1 U2899 ( .A1(n3923), .A2(n3922), .ZN(n2172) );
  OR2_X1 U2900 ( .A1(n4500), .A2(n4480), .ZN(n2173) );
  NAND2_X1 U2901 ( .A1(n3008), .A2(n3005), .ZN(n2174) );
  NAND2_X1 U2902 ( .A1(n4547), .A2(n4525), .ZN(n2301) );
  AND2_X1 U2903 ( .A1(n4500), .A2(n4480), .ZN(n2175) );
  INV_X1 U2904 ( .A(n3671), .ZN(n2403) );
  OR2_X1 U2905 ( .A1(n2305), .A2(n2308), .ZN(n2176) );
  OR2_X1 U2906 ( .A1(n4582), .A2(n4564), .ZN(n2177) );
  AND2_X1 U2907 ( .A1(n2429), .A2(n2428), .ZN(n2178) );
  AND2_X1 U2908 ( .A1(n2409), .A2(n2148), .ZN(n2179) );
  OR2_X1 U2909 ( .A1(n2881), .A2(n3272), .ZN(n2180) );
  INV_X1 U2910 ( .A(n3801), .ZN(n2401) );
  INV_X1 U2911 ( .A(n2891), .ZN(n4883) );
  INV_X1 U2912 ( .A(n4449), .ZN(n2369) );
  INV_X1 U2913 ( .A(n3452), .ZN(n2426) );
  INV_X1 U2914 ( .A(n3764), .ZN(n2385) );
  INV_X1 U2915 ( .A(n4113), .ZN(n4120) );
  NOR2_X1 U2916 ( .A1(n2748), .A2(n2449), .ZN(n2780) );
  NAND2_X1 U2917 ( .A1(n3163), .A2(n3162), .ZN(n2181) );
  OR2_X1 U2918 ( .A1(n2432), .A2(n4883), .ZN(n2182) );
  NAND2_X1 U2919 ( .A1(n3079), .A2(n3045), .ZN(n2183) );
  AND2_X1 U2920 ( .A1(n2653), .A2(n2663), .ZN(n2896) );
  INV_X1 U2921 ( .A(n2896), .ZN(n4880) );
  AND2_X1 U2922 ( .A1(n3997), .A2(REG1_REG_15__SCAN_IN), .ZN(n2184) );
  XNOR2_X1 U2923 ( .A(n2577), .B(IR_REG_10__SCAN_IN), .ZN(n2882) );
  INV_X1 U2924 ( .A(n2882), .ZN(n2359) );
  INV_X1 U2925 ( .A(REG2_REG_8__SCAN_IN), .ZN(n2265) );
  NAND2_X1 U2926 ( .A1(n2593), .A2(n2585), .ZN(n4776) );
  INV_X1 U2927 ( .A(n4776), .ZN(n2210) );
  NAND2_X1 U2928 ( .A1(n4939), .A2(REG1_REG_29__SCAN_IN), .ZN(n2195) );
  INV_X2 U2929 ( .A(n4939), .ZN(n4941) );
  NAND2_X1 U2930 ( .A1(n4627), .A2(n2185), .ZN(U3545) );
  NAND2_X1 U2931 ( .A1(n2344), .A2(n3871), .ZN(n4069) );
  NAND2_X1 U2932 ( .A1(n2531), .A2(REG3_REG_6__SCAN_IN), .ZN(n2547) );
  OR2_X4 U2933 ( .A1(n2688), .A2(n2681), .ZN(n2690) );
  NAND3_X1 U2934 ( .A1(n4029), .A2(n4095), .A3(n2186), .ZN(n3889) );
  AND2_X2 U2935 ( .A1(n4039), .A2(n4041), .ZN(n4029) );
  AND2_X2 U2936 ( .A1(n4054), .A2(n2735), .ZN(n4059) );
  NAND2_X1 U2937 ( .A1(n2202), .A2(n2166), .ZN(n2557) );
  NAND2_X1 U2938 ( .A1(n2658), .A2(REG3_REG_19__SCAN_IN), .ZN(n2668) );
  INV_X1 U2939 ( .A(n4074), .ZN(n4051) );
  OAI21_X1 U2940 ( .B1(n3362), .B2(n3361), .A(n3360), .ZN(n3364) );
  NAND2_X1 U2941 ( .A1(n2380), .A2(n2381), .ZN(n3722) );
  NOR2_X2 U2942 ( .A1(n3365), .A2(n3366), .ZN(n3424) );
  OAI22_X1 U2943 ( .A1(n3059), .A2(n2123), .B1(n3245), .B2(n3611), .ZN(n3032)
         );
  INV_X1 U2944 ( .A(n3663), .ZN(n2191) );
  NAND2_X1 U2945 ( .A1(n3647), .A2(n2434), .ZN(n3711) );
  NAND2_X1 U2946 ( .A1(n3279), .A2(n3282), .ZN(n2188) );
  NAND3_X1 U2947 ( .A1(n2190), .A2(n2200), .A3(n2189), .ZN(U3515) );
  INV_X1 U2948 ( .A(n4717), .ZN(n4639) );
  NAND2_X1 U2949 ( .A1(n4452), .A2(n4607), .ZN(n2214) );
  NAND2_X1 U2950 ( .A1(n3543), .A2(n2436), .ZN(n3547) );
  INV_X1 U2951 ( .A(n2208), .ZN(n3994) );
  INV_X1 U2952 ( .A(n4824), .ZN(n2192) );
  OAI21_X2 U2953 ( .B1(n4835), .B2(n2252), .A(n2251), .ZN(n4847) );
  NAND2_X1 U2954 ( .A1(n2977), .A2(n2864), .ZN(n2866) );
  NAND2_X1 U2955 ( .A1(n2208), .A2(n2207), .ZN(n3991) );
  NAND2_X2 U2956 ( .A1(n4819), .A2(n4820), .ZN(n4818) );
  OR2_X1 U2957 ( .A1(n2841), .A2(n2986), .ZN(n2194) );
  XNOR2_X2 U2958 ( .A(n2510), .B(IR_REG_3__SCAN_IN), .ZN(n2865) );
  NAND2_X1 U2959 ( .A1(n4792), .A2(n2884), .ZN(n3397) );
  NAND2_X1 U2960 ( .A1(n4793), .A2(REG2_REG_10__SCAN_IN), .ZN(n4792) );
  NAND2_X1 U2961 ( .A1(n2880), .A2(n2257), .ZN(n2256) );
  NAND2_X2 U2962 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n4177) );
  INV_X1 U2963 ( .A(n2201), .ZN(n2642) );
  INV_X1 U2964 ( .A(n2340), .ZN(n2339) );
  XNOR2_X2 U2965 ( .A(n2734), .B(REG3_REG_27__SCAN_IN), .ZN(n4080) );
  NAND2_X1 U2966 ( .A1(n3153), .A2(n2203), .ZN(n3154) );
  NAND2_X1 U2967 ( .A1(n3152), .A2(n3597), .ZN(n2203) );
  NAND2_X1 U2968 ( .A1(n4706), .A2(n2204), .ZN(U3512) );
  NAND3_X1 U2969 ( .A1(n2346), .A2(n2347), .A3(n2153), .ZN(n2924) );
  OAI22_X2 U2970 ( .A1(n3242), .A2(n2501), .B1(n3059), .B2(n3245), .ZN(n3098)
         );
  AOI21_X4 U2971 ( .B1(n3380), .B2(n3902), .A(n2592), .ZN(n3409) );
  INV_X1 U2972 ( .A(n2827), .ZN(n3079) );
  NAND2_X1 U2973 ( .A1(n2791), .A2(n2792), .ZN(n2827) );
  NAND2_X2 U2974 ( .A1(n3586), .A2(n3712), .ZN(n3673) );
  OAI21_X2 U2975 ( .B1(n3424), .B2(n2425), .A(n2423), .ZN(n3505) );
  NAND2_X1 U2976 ( .A1(n3644), .A2(n3577), .ZN(n3647) );
  NAND2_X1 U2977 ( .A1(n2397), .A2(n2395), .ZN(n3610) );
  OR2_X4 U2978 ( .A1(n4924), .A2(n3026), .ZN(n3615) );
  NAND3_X1 U2979 ( .A1(n3207), .A2(n3165), .A3(n2404), .ZN(n2206) );
  NAND2_X1 U2980 ( .A1(n2965), .A2(n3226), .ZN(n2968) );
  XNOR2_X1 U2981 ( .A(n2883), .B(n2359), .ZN(n4793) );
  NAND2_X1 U2982 ( .A1(n2349), .A2(n3836), .ZN(n3193) );
  NAND2_X1 U2983 ( .A1(n3308), .A2(n3840), .ZN(n2348) );
  NAND2_X1 U2984 ( .A1(n2122), .A2(n2445), .ZN(n2461) );
  INV_X1 U2985 ( .A(n2613), .ZN(n2496) );
  NAND2_X1 U2987 ( .A1(n3122), .A2(n3845), .ZN(n2349) );
  NAND2_X1 U2988 ( .A1(n4799), .A2(REG1_REG_10__SCAN_IN), .ZN(n4798) );
  AOI21_X2 U2989 ( .B1(n3232), .B2(n3231), .A(n2170), .ZN(n2846) );
  INV_X1 U2990 ( .A(n2220), .ZN(n2219) );
  OAI21_X2 U2991 ( .B1(n4818), .B2(n2226), .A(n2222), .ZN(n2220) );
  NAND2_X1 U2992 ( .A1(n4818), .A2(n2234), .ZN(n2233) );
  NAND2_X1 U2993 ( .A1(n4818), .A2(n2230), .ZN(n2229) );
  NAND2_X1 U2994 ( .A1(n2140), .A2(n2233), .ZN(n4830) );
  INV_X1 U2995 ( .A(n2374), .ZN(n2232) );
  NOR2_X1 U2996 ( .A1(n2235), .A2(n4883), .ZN(n2234) );
  INV_X1 U2997 ( .A(n2432), .ZN(n2235) );
  OR2_X2 U2998 ( .A1(n2998), .A2(n2530), .ZN(n2237) );
  MUX2_X1 U2999 ( .A(n2838), .B(REG1_REG_1__SCAN_IN), .S(n3965), .Z(n3970) );
  NAND3_X1 U3000 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .A3(
        IR_REG_0__SCAN_IN), .ZN(n2238) );
  NAND3_X1 U3001 ( .A1(n2241), .A2(n2243), .A3(n2239), .ZN(n2936) );
  NAND3_X1 U3002 ( .A1(n2241), .A2(n2240), .A3(n2239), .ZN(n2246) );
  NAND2_X1 U3003 ( .A1(n2971), .A2(n2372), .ZN(n2371) );
  NOR2_X1 U3004 ( .A1(n2244), .A2(n2865), .ZN(n2242) );
  NAND2_X1 U3005 ( .A1(n2244), .A2(n2865), .ZN(n2243) );
  INV_X1 U3006 ( .A(n2372), .ZN(n2244) );
  INV_X1 U3007 ( .A(n2865), .ZN(n2245) );
  INV_X1 U3008 ( .A(n2246), .ZN(n2935) );
  NOR2_X1 U3009 ( .A1(n4836), .A2(n2853), .ZN(n4854) );
  INV_X1 U3010 ( .A(n2895), .ZN(n2252) );
  XNOR2_X2 U3011 ( .A(n2893), .B(n2894), .ZN(n4835) );
  NAND3_X1 U3012 ( .A1(n2260), .A2(n2256), .A3(n2180), .ZN(n2883) );
  INV_X1 U3013 ( .A(n2269), .ZN(n3235) );
  XNOR2_X2 U3014 ( .A(n2270), .B(IR_REG_2__SCAN_IN), .ZN(n4780) );
  NAND2_X2 U3015 ( .A1(n3820), .A2(n3824), .ZN(n2753) );
  INV_X2 U3016 ( .A(n2486), .ZN(n3021) );
  NAND2_X2 U3017 ( .A1(n2477), .A2(n2476), .ZN(n2486) );
  OAI21_X1 U3018 ( .B1(n4699), .B2(n4588), .A(n2271), .ZN(U3354) );
  NAND2_X1 U3019 ( .A1(n3409), .A2(n2133), .ZN(n2281) );
  INV_X1 U3020 ( .A(n2604), .ZN(n2290) );
  NAND2_X1 U3021 ( .A1(n2291), .A2(n2292), .ZN(n4436) );
  NAND2_X1 U3022 ( .A1(n4512), .A2(n2134), .ZN(n2291) );
  NAND2_X1 U3023 ( .A1(n4512), .A2(n2302), .ZN(n2296) );
  NAND2_X1 U3024 ( .A1(n2448), .A2(n2431), .ZN(n2449) );
  NAND2_X1 U3025 ( .A1(n2307), .A2(n2306), .ZN(n2568) );
  NAND2_X1 U3026 ( .A1(n4127), .A2(n2317), .ZN(n2316) );
  NOR2_X1 U3027 ( .A1(n2332), .A2(IR_REG_2__SCAN_IN), .ZN(n2522) );
  OR2_X1 U3028 ( .A1(n4116), .A2(n2339), .ZN(n2335) );
  NAND2_X1 U3029 ( .A1(n2335), .A2(n2337), .ZN(n4042) );
  OR2_X1 U3030 ( .A1(n4116), .A2(n2777), .ZN(n2344) );
  NAND3_X1 U3031 ( .A1(n2347), .A2(n2153), .A3(n2345), .ZN(n2452) );
  INV_X2 U3032 ( .A(n2461), .ZN(n2347) );
  OAI21_X2 U3033 ( .B1(n3262), .B2(n3849), .A(n3841), .ZN(n3342) );
  OAI21_X2 U3034 ( .B1(n3404), .B2(n2761), .A(n3853), .ZN(n3918) );
  NAND2_X1 U3035 ( .A1(n2353), .A2(n2351), .ZN(n2776) );
  NAND2_X1 U3036 ( .A1(n2766), .A2(n2354), .ZN(n2353) );
  NAND2_X1 U3037 ( .A1(n2934), .A2(REG2_REG_3__SCAN_IN), .ZN(n2868) );
  XNOR2_X2 U3038 ( .A(n2866), .B(n2245), .ZN(n2934) );
  AND2_X2 U3039 ( .A1(n3991), .A2(n2892), .ZN(n2893) );
  NAND2_X1 U3040 ( .A1(n2167), .A2(n3256), .ZN(n3200) );
  NAND2_X2 U3041 ( .A1(n3084), .A2(n2960), .ZN(n3026) );
  NAND3_X2 U3042 ( .A1(n2818), .A2(n4774), .A3(n4773), .ZN(n2960) );
  XNOR2_X2 U3043 ( .A(n2379), .B(IR_REG_24__SCAN_IN), .ZN(n2818) );
  NAND2_X1 U3044 ( .A1(n3547), .A2(n2383), .ZN(n2380) );
  NAND2_X1 U3045 ( .A1(n3673), .A2(n2388), .ZN(n2387) );
  NAND2_X1 U3046 ( .A1(n3673), .A2(n2398), .ZN(n2397) );
  OAI211_X1 U3047 ( .C1(n3673), .C2(n2391), .A(n2168), .B(n2387), .ZN(n2400)
         );
  NAND2_X1 U3048 ( .A1(n3207), .A2(n2404), .ZN(n2408) );
  NAND2_X1 U3049 ( .A1(n2406), .A2(n3165), .ZN(n2405) );
  NAND2_X1 U3050 ( .A1(n2347), .A2(n2411), .ZN(n2811) );
  NAND2_X1 U3051 ( .A1(n2347), .A2(n2412), .ZN(n2805) );
  NAND2_X1 U3052 ( .A1(n3572), .A2(n2416), .ZN(n3644) );
  INV_X1 U3053 ( .A(n3746), .ZN(n2418) );
  NAND2_X1 U3054 ( .A1(n2419), .A2(n2420), .ZN(n3506) );
  NAND2_X1 U3055 ( .A1(n3424), .A2(n2422), .ZN(n2419) );
  INV_X1 U3056 ( .A(n2429), .ZN(n3433) );
  OR2_X1 U3057 ( .A1(n3423), .A2(n3426), .ZN(n2430) );
  NAND2_X2 U3058 ( .A1(n3010), .A2(n2879), .ZN(n2880) );
  NAND2_X1 U3059 ( .A1(n4807), .A2(n2850), .ZN(n4819) );
  NAND2_X1 U3060 ( .A1(n2902), .A2(n2901), .ZN(n2903) );
  NOR2_X2 U3061 ( .A1(n4678), .A2(n4600), .ZN(n4571) );
  NAND2_X1 U3062 ( .A1(n4536), .A2(n3880), .ZN(n4503) );
  NAND2_X1 U3063 ( .A1(n4017), .A2(n4049), .ZN(n4037) );
  INV_X1 U3064 ( .A(n4017), .ZN(n4035) );
  OAI21_X1 U3065 ( .B1(n4007), .B2(n2903), .A(n3768), .ZN(n2904) );
  NAND2_X1 U3066 ( .A1(n3807), .A2(DATAI_0_), .ZN(n2484) );
  AND2_X1 U3067 ( .A1(n2968), .A2(n2967), .ZN(n3018) );
  NAND2_X2 U3068 ( .A1(n2701), .A2(n2700), .ZN(n4127) );
  OAI22_X1 U3069 ( .A1(n2478), .A2(n3151), .B1(n3026), .B2(n3021), .ZN(n3020)
         );
  INV_X1 U3070 ( .A(n4780), .ZN(n2839) );
  INV_X1 U3071 ( .A(n4845), .ZN(n2901) );
  AND2_X2 U3072 ( .A1(n2823), .A2(n3075), .ZN(n4932) );
  OR2_X1 U3073 ( .A1(n4885), .A2(n4222), .ZN(n2432) );
  AND2_X1 U3074 ( .A1(n2633), .A2(n2639), .ZN(n3997) );
  INV_X1 U3075 ( .A(n4544), .ZN(n2666) );
  INV_X1 U3076 ( .A(n4582), .ZN(n3691) );
  NAND2_X1 U3077 ( .A1(n2811), .A2(IR_REG_31__SCAN_IN), .ZN(n2819) );
  OR2_X1 U3078 ( .A1(n4621), .A2(n4900), .ZN(n2433) );
  INV_X1 U3079 ( .A(n4564), .ZN(n4555) );
  AND2_X1 U3080 ( .A1(n3582), .A2(n3583), .ZN(n2434) );
  NAND2_X1 U3081 ( .A1(n3534), .A2(n3528), .ZN(n2435) );
  AND3_X1 U3082 ( .A1(n3542), .A2(n3541), .A3(n3540), .ZN(n2436) );
  NOR2_X2 U3083 ( .A1(IR_REG_15__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .ZN(n2462)
         );
  AND2_X1 U3084 ( .A1(n3885), .A2(n4093), .ZN(n3931) );
  INV_X1 U3085 ( .A(n4066), .ZN(n4068) );
  INV_X1 U3086 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2569) );
  INV_X1 U3087 ( .A(REG3_REG_9__SCAN_IN), .ZN(n3233) );
  OAI21_X1 U3088 ( .B1(n2698), .B2(n4437), .A(n2697), .ZN(n2699) );
  NAND2_X1 U3089 ( .A1(n2125), .A2(DATAI_1_), .ZN(n2476) );
  OR2_X1 U3090 ( .A1(n3026), .A2(n3080), .ZN(n2961) );
  INV_X1 U3091 ( .A(n3701), .ZN(n3544) );
  INV_X1 U3092 ( .A(n3715), .ZN(n4140) );
  OR2_X1 U3093 ( .A1(n4506), .A2(n2716), .ZN(n2674) );
  INV_X1 U3094 ( .A(n2699), .ZN(n2700) );
  INV_X1 U3095 ( .A(n3211), .ZN(n2824) );
  INV_X1 U3096 ( .A(n2755), .ZN(n3282) );
  AND2_X1 U3097 ( .A1(n3517), .A2(n3516), .ZN(n3680) );
  AND2_X1 U3098 ( .A1(n3537), .A2(n3536), .ZN(n3701) );
  AND2_X1 U3099 ( .A1(n3049), .A2(n3050), .ZN(n3038) );
  INV_X1 U3100 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3727) );
  NAND2_X1 U3101 ( .A1(n3545), .A2(n3544), .ZN(n3546) );
  AND2_X1 U3102 ( .A1(n2648), .A2(n2647), .ZN(n4582) );
  AND2_X1 U3103 ( .A1(n3886), .A2(n3885), .ZN(n4095) );
  INV_X1 U3104 ( .A(n4601), .ZN(n4545) );
  INV_X1 U3105 ( .A(n3760), .ZN(n3292) );
  INV_X1 U3106 ( .A(n4565), .ZN(n4599) );
  OR2_X1 U3107 ( .A1(n2827), .A2(n2828), .ZN(n4565) );
  NAND2_X1 U3108 ( .A1(n2433), .A2(n4623), .ZN(n4698) );
  INV_X1 U3109 ( .A(n4099), .ZN(n4088) );
  NAND2_X1 U3110 ( .A1(n4582), .A2(n4564), .ZN(n2654) );
  AND2_X1 U3111 ( .A1(n2779), .A2(n2778), .ZN(n4496) );
  NOR2_X1 U3112 ( .A1(n2748), .A2(IR_REG_14__SCAN_IN), .ZN(n2650) );
  INV_X1 U3113 ( .A(n2625), .ZN(n3641) );
  INV_X1 U3114 ( .A(n3772), .ZN(n3796) );
  INV_X1 U3115 ( .A(n4135), .ZN(n4128) );
  AND2_X1 U3116 ( .A1(n2125), .A2(DATAI_22_), .ZN(n4462) );
  OR2_X1 U3117 ( .A1(n2718), .A2(n2711), .ZN(n3674) );
  NAND2_X1 U3118 ( .A1(n2638), .A2(n2637), .ZN(n4561) );
  NOR2_X1 U3119 ( .A1(n4858), .A2(n2905), .ZN(n2906) );
  INV_X1 U3120 ( .A(n4604), .ZN(n4559) );
  AND2_X1 U3121 ( .A1(n4585), .A2(n4012), .ZN(n4539) );
  OR2_X1 U3122 ( .A1(n3052), .A2(n3060), .ZN(n4592) );
  INV_X1 U3123 ( .A(n4675), .ZN(n4667) );
  OR2_X1 U3124 ( .A1(n4932), .A2(n4312), .ZN(n2829) );
  OR2_X1 U3125 ( .A1(n3078), .A2(n3950), .ZN(n4894) );
  INV_X1 U3126 ( .A(n4496), .ZN(n4607) );
  INV_X1 U3127 ( .A(n4766), .ZN(n4755) );
  INV_X1 U3128 ( .A(n2818), .ZN(n2808) );
  AND2_X1 U3129 ( .A1(n2860), .A2(n2859), .ZN(n4851) );
  OR2_X1 U3130 ( .A1(n2960), .A2(n2908), .ZN(n3962) );
  OR2_X1 U3131 ( .A1(n4791), .A2(n3948), .ZN(n4845) );
  OR2_X1 U3132 ( .A1(n4791), .A2(n3067), .ZN(n4858) );
  INV_X1 U3133 ( .A(n4576), .ZN(n4594) );
  AND2_X1 U3134 ( .A1(n4511), .A2(n3132), .ZN(n4588) );
  AND2_X1 U3135 ( .A1(n2834), .A2(n2833), .ZN(n2835) );
  NAND2_X1 U3136 ( .A1(n4941), .A2(n4924), .ZN(n4675) );
  OR2_X1 U3137 ( .A1(n2832), .A2(n3075), .ZN(n4939) );
  AND2_X1 U3138 ( .A1(n2830), .A2(n2829), .ZN(n2831) );
  INV_X1 U3139 ( .A(n4932), .ZN(n4930) );
  INV_X1 U3140 ( .A(n4876), .ZN(n4875) );
  NAND2_X1 U3141 ( .A1(n3039), .A2(n2932), .ZN(n4876) );
  INV_X1 U3142 ( .A(n2894), .ZN(n4881) );
  INV_X2 U3143 ( .A(n3962), .ZN(U4043) );
  NOR2_X2 U3144 ( .A1(n4177), .A2(n2515), .ZN(n2531) );
  OR2_X2 U3145 ( .A1(n2557), .A2(n3233), .ZN(n2570) );
  NAND2_X1 U3146 ( .A1(REG3_REG_17__SCAN_IN), .A2(REG3_REG_16__SCAN_IN), .ZN(
        n2437) );
  AND2_X2 U3147 ( .A1(n2656), .A2(REG3_REG_18__SCAN_IN), .ZN(n2658) );
  OR2_X1 U31480 ( .A1(n2658), .A2(REG3_REG_19__SCAN_IN), .ZN(n2438) );
  AND2_X1 U31490 ( .A1(n2668), .A2(n2438), .ZN(n4515) );
  NAND4_X1 U3150 ( .A1(n2442), .A2(n2441), .A3(n2440), .A4(n2439), .ZN(n2614)
         );
  INV_X1 U3151 ( .A(n2614), .ZN(n2445) );
  NAND4_X1 U3152 ( .A1(n2462), .A2(n2447), .A3(n2446), .A4(n2744), .ZN(n2746)
         );
  INV_X1 U3153 ( .A(n2746), .ZN(n2448) );
  NOR2_X2 U3154 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2809)
         );
  XNOR2_X2 U3155 ( .A(n2451), .B(IR_REG_30__SCAN_IN), .ZN(n4771) );
  XNOR2_X2 U3156 ( .A(n2453), .B(IR_REG_29__SCAN_IN), .ZN(n4772) );
  AND2_X2 U3157 ( .A1(n4771), .A2(n4772), .ZN(n2469) );
  NAND2_X1 U3158 ( .A1(n4515), .A2(n2789), .ZN(n2460) );
  INV_X1 U3159 ( .A(n4771), .ZN(n2454) );
  INV_X1 U3160 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4656) );
  INV_X1 U3161 ( .A(n4772), .ZN(n2455) );
  AND2_X2 U3162 ( .A1(n4771), .A2(n2455), .ZN(n2470) );
  NAND2_X1 U3163 ( .A1(n2941), .A2(REG2_REG_19__SCAN_IN), .ZN(n2457) );
  NOR2_X1 U3164 ( .A1(n4771), .A2(n4772), .ZN(n2479) );
  NAND2_X1 U3165 ( .A1(n3803), .A2(REG0_REG_19__SCAN_IN), .ZN(n2456) );
  OAI211_X1 U3166 ( .C1(n3806), .C2(n4656), .A(n2457), .B(n2456), .ZN(n2458)
         );
  INV_X1 U3167 ( .A(n2458), .ZN(n2459) );
  INV_X1 U3168 ( .A(IR_REG_16__SCAN_IN), .ZN(n2464) );
  INV_X1 U3169 ( .A(IR_REG_17__SCAN_IN), .ZN(n2463) );
  NAND4_X1 U3170 ( .A1(n2462), .A2(n2464), .A3(n2664), .A4(n2463), .ZN(n2465)
         );
  OAI21_X2 U3171 ( .B1(n2461), .B2(n2465), .A(IR_REG_31__SCAN_IN), .ZN(n2742)
         );
  MUX2_X1 U3172 ( .A(n4004), .B(DATAI_19_), .S(n2126), .Z(n4525) );
  INV_X1 U3173 ( .A(n4525), .ZN(n3880) );
  INV_X1 U3174 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2838) );
  NAND2_X1 U3175 ( .A1(n2479), .A2(REG0_REG_1__SCAN_IN), .ZN(n2473) );
  NAND2_X1 U3176 ( .A1(n2469), .A2(REG3_REG_1__SCAN_IN), .ZN(n2472) );
  NAND2_X1 U3177 ( .A1(n2470), .A2(REG2_REG_1__SCAN_IN), .ZN(n2471) );
  INV_X1 U3178 ( .A(n3965), .ZN(n4781) );
  NAND2_X1 U3179 ( .A1(n2475), .A2(n4781), .ZN(n2477) );
  INV_X1 U3180 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2963) );
  NAND2_X1 U3181 ( .A1(n2469), .A2(REG3_REG_0__SCAN_IN), .ZN(n2482) );
  NAND2_X1 U3182 ( .A1(n2479), .A2(REG0_REG_0__SCAN_IN), .ZN(n2481) );
  NAND2_X1 U3183 ( .A1(n2470), .A2(REG2_REG_0__SCAN_IN), .ZN(n2480) );
  INV_X2 U3184 ( .A(IR_REG_0__SCAN_IN), .ZN(n2485) );
  OAI21_X2 U3185 ( .B1(n2126), .B2(n2485), .A(n2484), .ZN(n3189) );
  NAND2_X1 U3186 ( .A1(n2753), .A2(n3174), .ZN(n3176) );
  NAND2_X1 U3187 ( .A1(n3758), .A2(n2486), .ZN(n2487) );
  NAND2_X1 U3188 ( .A1(n3176), .A2(n2487), .ZN(n3281) );
  INV_X1 U3189 ( .A(n3281), .ZN(n2492) );
  MUX2_X1 U3190 ( .A(n4780), .B(DATAI_2_), .S(n2125), .Z(n3760) );
  OR2_X1 U3191 ( .A1(n2504), .A2(n2840), .ZN(n2491) );
  NAND2_X1 U3192 ( .A1(n2495), .A2(REG0_REG_2__SCAN_IN), .ZN(n2490) );
  NAND2_X1 U3193 ( .A1(n2470), .A2(REG2_REG_2__SCAN_IN), .ZN(n2489) );
  NAND2_X1 U3194 ( .A1(n2469), .A2(REG3_REG_2__SCAN_IN), .ZN(n2488) );
  AND4_X2 U3195 ( .A1(n2491), .A2(n2490), .A3(n2489), .A4(n2488), .ZN(n3246)
         );
  INV_X1 U3196 ( .A(n3246), .ZN(n3964) );
  NAND2_X1 U3197 ( .A1(n3292), .A2(n3964), .ZN(n3828) );
  NAND2_X1 U3198 ( .A1(n3828), .A2(n3825), .ZN(n2755) );
  NAND2_X1 U3199 ( .A1(n2492), .A2(n2755), .ZN(n3280) );
  NAND2_X1 U3200 ( .A1(n3246), .A2(n3292), .ZN(n2493) );
  NAND2_X1 U3201 ( .A1(n3280), .A2(n2493), .ZN(n3242) );
  INV_X1 U3202 ( .A(REG1_REG_3__SCAN_IN), .ZN(n2494) );
  OR2_X1 U3203 ( .A1(n2504), .A2(n2494), .ZN(n2500) );
  NAND2_X1 U3204 ( .A1(n2495), .A2(REG0_REG_3__SCAN_IN), .ZN(n2499) );
  NAND2_X1 U3205 ( .A1(n2496), .A2(REG2_REG_3__SCAN_IN), .ZN(n2498) );
  NAND2_X1 U3206 ( .A1(n2469), .A2(n4237), .ZN(n2497) );
  OR2_X1 U3207 ( .A1(n2522), .A2(n2923), .ZN(n2510) );
  MUX2_X1 U3208 ( .A(n2865), .B(DATAI_3_), .S(n2125), .Z(n3254) );
  NOR2_X1 U3209 ( .A1(n3963), .A2(n3254), .ZN(n2501) );
  INV_X1 U32100 ( .A(n3254), .ZN(n3245) );
  NAND2_X1 U32110 ( .A1(n3803), .A2(REG0_REG_4__SCAN_IN), .ZN(n2508) );
  NAND2_X1 U32120 ( .A1(n2496), .A2(REG2_REG_4__SCAN_IN), .ZN(n2507) );
  OAI21_X1 U32130 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        n4177), .ZN(n3106) );
  INV_X1 U32140 ( .A(n3106), .ZN(n2502) );
  NAND2_X1 U32150 ( .A1(n2789), .A2(n2502), .ZN(n2506) );
  INV_X1 U32160 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2503) );
  OR2_X1 U32170 ( .A1(n3806), .A2(n2503), .ZN(n2505) );
  AND4_X2 U32180 ( .A1(n2508), .A2(n2507), .A3(n2506), .A4(n2505), .ZN(n3247)
         );
  NAND2_X1 U32190 ( .A1(n2510), .A2(n2509), .ZN(n2511) );
  NAND2_X1 U32200 ( .A1(n2511), .A2(IR_REG_31__SCAN_IN), .ZN(n2512) );
  XNOR2_X1 U32210 ( .A(n2512), .B(IR_REG_4__SCAN_IN), .ZN(n2869) );
  MUX2_X1 U32220 ( .A(n2869), .B(DATAI_4_), .S(n2126), .Z(n3100) );
  NAND2_X1 U32230 ( .A1(n3247), .A2(n3100), .ZN(n3831) );
  INV_X1 U32240 ( .A(n3247), .ZN(n3136) );
  NAND2_X1 U32250 ( .A1(n3136), .A2(n3105), .ZN(n3834) );
  NAND2_X1 U32260 ( .A1(n3831), .A2(n3834), .ZN(n3900) );
  NAND2_X1 U32270 ( .A1(n3098), .A2(n3900), .ZN(n2514) );
  NAND2_X1 U32280 ( .A1(n3136), .A2(n3100), .ZN(n2513) );
  NAND2_X1 U32290 ( .A1(n2514), .A2(n2513), .ZN(n3133) );
  INV_X1 U32300 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2842) );
  OR2_X1 U32310 ( .A1(n3806), .A2(n2842), .ZN(n2520) );
  NAND2_X1 U32320 ( .A1(n3803), .A2(REG0_REG_5__SCAN_IN), .ZN(n2519) );
  AND2_X1 U32330 ( .A1(n4177), .A2(n2515), .ZN(n2516) );
  NOR2_X1 U32340 ( .A1(n2531), .A2(n2516), .ZN(n3209) );
  NAND2_X1 U32350 ( .A1(n2789), .A2(n3209), .ZN(n2518) );
  NAND2_X1 U32360 ( .A1(n2496), .A2(REG2_REG_5__SCAN_IN), .ZN(n2517) );
  NAND4_X1 U32370 ( .A1(n2520), .A2(n2519), .A3(n2518), .A4(n2517), .ZN(n3152)
         );
  NOR2_X1 U32380 ( .A1(n2525), .A2(n2923), .ZN(n2523) );
  MUX2_X1 U32390 ( .A(n2923), .B(n2523), .S(IR_REG_5__SCAN_IN), .Z(n2527) );
  INV_X1 U32400 ( .A(n2615), .ZN(n2526) );
  MUX2_X1 U32410 ( .A(n4779), .B(DATAI_5_), .S(n2125), .Z(n3211) );
  AND2_X1 U32420 ( .A1(n3152), .A2(n3211), .ZN(n2528) );
  NAND2_X1 U32430 ( .A1(n3218), .A2(n2824), .ZN(n2529) );
  INV_X1 U32440 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2530) );
  OR2_X1 U32450 ( .A1(n3806), .A2(n2530), .ZN(n2536) );
  NAND2_X1 U32460 ( .A1(n3803), .A2(REG0_REG_6__SCAN_IN), .ZN(n2535) );
  NAND2_X1 U32470 ( .A1(n2496), .A2(REG2_REG_6__SCAN_IN), .ZN(n2534) );
  OR2_X1 U32480 ( .A1(n2531), .A2(REG3_REG_6__SCAN_IN), .ZN(n2532) );
  AND2_X1 U32490 ( .A1(n2547), .A2(n2532), .ZN(n3301) );
  NAND2_X1 U32500 ( .A1(n2789), .A2(n3301), .ZN(n2533) );
  NAND4_X1 U32510 ( .A1(n2536), .A2(n2535), .A3(n2534), .A4(n2533), .ZN(n3961)
         );
  NAND2_X1 U32520 ( .A1(n2615), .A2(IR_REG_31__SCAN_IN), .ZN(n2537) );
  XNOR2_X1 U32530 ( .A(n2537), .B(IR_REG_6__SCAN_IN), .ZN(n2874) );
  MUX2_X1 U32540 ( .A(n2874), .B(DATAI_6_), .S(n2126), .Z(n3220) );
  NOR2_X1 U32550 ( .A1(n3961), .A2(n3220), .ZN(n2538) );
  NAND2_X1 U32560 ( .A1(n3803), .A2(REG0_REG_7__SCAN_IN), .ZN(n2542) );
  NAND2_X1 U32570 ( .A1(n2496), .A2(REG2_REG_7__SCAN_IN), .ZN(n2541) );
  XNOR2_X1 U32580 ( .A(n2547), .B(REG3_REG_7__SCAN_IN), .ZN(n3169) );
  NAND2_X1 U32590 ( .A1(n2789), .A2(n3169), .ZN(n2540) );
  INV_X1 U32600 ( .A(REG1_REG_7__SCAN_IN), .ZN(n3005) );
  OR2_X1 U32610 ( .A1(n3806), .A2(n3005), .ZN(n2539) );
  MUX2_X1 U32620 ( .A(n3004), .B(DATAI_7_), .S(n2125), .Z(n3201) );
  NAND2_X1 U32630 ( .A1(n3330), .A2(n3201), .ZN(n2758) );
  INV_X1 U32640 ( .A(n3201), .ZN(n3194) );
  NAND2_X1 U32650 ( .A1(n3960), .A2(n3194), .ZN(n3839) );
  NAND2_X1 U32660 ( .A1(n2758), .A2(n3839), .ZN(n3899) );
  NAND2_X1 U32670 ( .A1(n3199), .A2(n3899), .ZN(n2544) );
  NAND2_X1 U32680 ( .A1(n3960), .A2(n3201), .ZN(n2543) );
  INV_X1 U32690 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4395) );
  OR2_X1 U32700 ( .A1(n3806), .A2(n4395), .ZN(n2552) );
  NAND2_X1 U32710 ( .A1(n3803), .A2(REG0_REG_8__SCAN_IN), .ZN(n2551) );
  INV_X1 U32720 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2546) );
  INV_X1 U32730 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2545) );
  OAI21_X1 U32740 ( .B1(n2547), .B2(n2546), .A(n2545), .ZN(n2548) );
  AND2_X1 U32750 ( .A1(n2548), .A2(n2557), .ZN(n3328) );
  NAND2_X1 U32760 ( .A1(n2789), .A2(n3328), .ZN(n2550) );
  NAND2_X1 U32770 ( .A1(n2941), .A2(REG2_REG_8__SCAN_IN), .ZN(n2549) );
  NAND4_X1 U32780 ( .A1(n2552), .A2(n2551), .A3(n2550), .A4(n2549), .ZN(n3263)
         );
  INV_X1 U32790 ( .A(IR_REG_7__SCAN_IN), .ZN(n4161) );
  NAND2_X1 U32800 ( .A1(n2553), .A2(n4161), .ZN(n2554) );
  NAND2_X1 U32810 ( .A1(n2554), .A2(IR_REG_31__SCAN_IN), .ZN(n2555) );
  XNOR2_X1 U32820 ( .A(n2555), .B(IR_REG_8__SCAN_IN), .ZN(n4778) );
  MUX2_X1 U32830 ( .A(n4778), .B(DATAI_8_), .S(n2126), .Z(n3332) );
  AND2_X1 U32840 ( .A1(n3263), .A2(n3332), .ZN(n2556) );
  INV_X1 U32850 ( .A(REG1_REG_9__SCAN_IN), .ZN(n4219) );
  OR2_X1 U32860 ( .A1(n3806), .A2(n4219), .ZN(n2563) );
  NAND2_X1 U32870 ( .A1(n3803), .A2(REG0_REG_9__SCAN_IN), .ZN(n2562) );
  NAND2_X1 U32880 ( .A1(n2941), .A2(REG2_REG_9__SCAN_IN), .ZN(n2561) );
  NAND2_X1 U32890 ( .A1(n2557), .A2(n3233), .ZN(n2558) );
  NAND2_X1 U32900 ( .A1(n2570), .A2(n2558), .ZN(n3370) );
  INV_X1 U32910 ( .A(n3370), .ZN(n2559) );
  NAND2_X1 U32920 ( .A1(n2789), .A2(n2559), .ZN(n2560) );
  NAND4_X1 U32930 ( .A1(n2563), .A2(n2562), .A3(n2561), .A4(n2560), .ZN(n3959)
         );
  NOR2_X1 U32940 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2564)
         );
  NAND2_X1 U32950 ( .A1(n2565), .A2(n2564), .ZN(n2576) );
  NAND2_X1 U32960 ( .A1(n2576), .A2(IR_REG_31__SCAN_IN), .ZN(n2566) );
  MUX2_X1 U32970 ( .A(n4777), .B(DATAI_9_), .S(n2126), .Z(n3373) );
  NAND2_X1 U32980 ( .A1(n3959), .A2(n3373), .ZN(n2567) );
  INV_X1 U32990 ( .A(n3346), .ZN(n2578) );
  INV_X1 U33000 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4378) );
  OR2_X1 U33010 ( .A1(n3806), .A2(n4378), .ZN(n2575) );
  NAND2_X1 U33020 ( .A1(n3803), .A2(REG0_REG_10__SCAN_IN), .ZN(n2574) );
  AND2_X1 U33030 ( .A1(n2570), .A2(n2569), .ZN(n2571) );
  NOR2_X1 U33040 ( .A1(n2586), .A2(n2571), .ZN(n3349) );
  NAND2_X1 U33050 ( .A1(n2789), .A2(n3349), .ZN(n2573) );
  NAND2_X1 U33060 ( .A1(n2941), .A2(REG2_REG_10__SCAN_IN), .ZN(n2572) );
  NAND4_X1 U33070 ( .A1(n2575), .A2(n2574), .A3(n2573), .A4(n2572), .ZN(n3415)
         );
  NAND2_X1 U33080 ( .A1(n2581), .A2(IR_REG_31__SCAN_IN), .ZN(n2577) );
  MUX2_X1 U33090 ( .A(n2882), .B(DATAI_10_), .S(n2126), .Z(n3419) );
  NAND2_X1 U33100 ( .A1(n2578), .A2(n2152), .ZN(n2580) );
  INV_X1 U33110 ( .A(n3419), .ZN(n3429) );
  NAND2_X1 U33120 ( .A1(n3443), .A2(n3429), .ZN(n2579) );
  NAND2_X1 U33130 ( .A1(n2582), .A2(IR_REG_31__SCAN_IN), .ZN(n2584) );
  NAND2_X1 U33140 ( .A1(n2584), .A2(n2583), .ZN(n2593) );
  OR2_X1 U33150 ( .A1(n2584), .A2(n2583), .ZN(n2585) );
  INV_X1 U33160 ( .A(DATAI_11_), .ZN(n4380) );
  MUX2_X1 U33170 ( .A(n4776), .B(n4380), .S(n2126), .Z(n3437) );
  INV_X1 U33180 ( .A(n3437), .ZN(n3448) );
  NAND2_X1 U33190 ( .A1(n3803), .A2(REG0_REG_11__SCAN_IN), .ZN(n2591) );
  OR2_X1 U33200 ( .A1(n2586), .A2(REG3_REG_11__SCAN_IN), .ZN(n2587) );
  AND2_X1 U33210 ( .A1(n2587), .A2(n2598), .ZN(n3444) );
  NAND2_X1 U33220 ( .A1(n2789), .A2(n3444), .ZN(n2590) );
  NAND2_X1 U33230 ( .A1(n2941), .A2(REG2_REG_11__SCAN_IN), .ZN(n2589) );
  INV_X1 U33240 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4221) );
  OR2_X1 U33250 ( .A1(n3806), .A2(n4221), .ZN(n2588) );
  NAND2_X1 U33260 ( .A1(n3448), .A2(n3457), .ZN(n3403) );
  NAND2_X1 U33270 ( .A1(n3437), .A2(n3958), .ZN(n3817) );
  NAND2_X1 U33280 ( .A1(n3403), .A2(n3817), .ZN(n3902) );
  NOR2_X1 U33290 ( .A1(n3448), .A2(n3958), .ZN(n2592) );
  INV_X1 U33300 ( .A(DATAI_12_), .ZN(n2596) );
  NAND2_X1 U33310 ( .A1(n2593), .A2(IR_REG_31__SCAN_IN), .ZN(n2595) );
  MUX2_X1 U33320 ( .A(n2596), .B(n4886), .S(n2475), .Z(n3454) );
  NAND2_X1 U33330 ( .A1(n3803), .A2(REG0_REG_12__SCAN_IN), .ZN(n2603) );
  NAND2_X1 U33340 ( .A1(n2941), .A2(REG2_REG_12__SCAN_IN), .ZN(n2602) );
  NAND2_X1 U33350 ( .A1(n2598), .A2(n2597), .ZN(n2599) );
  AND2_X1 U33360 ( .A1(n2606), .A2(n2599), .ZN(n3456) );
  NAND2_X1 U33370 ( .A1(n2789), .A2(n3456), .ZN(n2601) );
  INV_X1 U33380 ( .A(REG1_REG_12__SCAN_IN), .ZN(n3466) );
  OR2_X1 U33390 ( .A1(n3806), .A2(n3466), .ZN(n2600) );
  NAND2_X1 U33400 ( .A1(n3454), .A2(n3738), .ZN(n2605) );
  NOR2_X1 U33410 ( .A1(n3454), .A2(n3738), .ZN(n2604) );
  INV_X1 U33420 ( .A(REG2_REG_13__SCAN_IN), .ZN(n2612) );
  AND2_X1 U33430 ( .A1(n2606), .A2(n4217), .ZN(n2607) );
  NOR2_X1 U33440 ( .A1(n2617), .A2(n2607), .ZN(n3737) );
  NAND2_X1 U33450 ( .A1(n3737), .A2(n2789), .ZN(n2611) );
  NAND2_X1 U33460 ( .A1(n3803), .A2(REG0_REG_13__SCAN_IN), .ZN(n2609) );
  INV_X1 U33470 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4222) );
  OR2_X1 U33480 ( .A1(n3806), .A2(n4222), .ZN(n2608) );
  AND2_X1 U33490 ( .A1(n2609), .A2(n2608), .ZN(n2610) );
  OAI211_X1 U33500 ( .C1(n2613), .C2(n2612), .A(n2611), .B(n2610), .ZN(n3636)
         );
  OAI21_X1 U33510 ( .B1(n2615), .B2(n2614), .A(IR_REG_31__SCAN_IN), .ZN(n2616)
         );
  XNOR2_X1 U33520 ( .A(n2616), .B(IR_REG_13__SCAN_IN), .ZN(n2889) );
  MUX2_X1 U3353 ( .A(n2889), .B(DATAI_13_), .S(n2125), .Z(n3740) );
  OR2_X1 U33540 ( .A1(n2617), .A2(REG3_REG_14__SCAN_IN), .ZN(n2618) );
  NAND2_X1 U3355 ( .A1(n2626), .A2(n2618), .ZN(n3638) );
  INV_X1 U3356 ( .A(n3806), .ZN(n2619) );
  AOI22_X1 U3357 ( .A1(n2619), .A2(REG1_REG_14__SCAN_IN), .B1(n3803), .B2(
        REG0_REG_14__SCAN_IN), .ZN(n2621) );
  NAND2_X1 U3358 ( .A1(n2941), .A2(REG2_REG_14__SCAN_IN), .ZN(n2620) );
  NAND2_X1 U3359 ( .A1(n2748), .A2(IR_REG_31__SCAN_IN), .ZN(n2622) );
  MUX2_X1 U3360 ( .A(IR_REG_31__SCAN_IN), .B(n2622), .S(IR_REG_14__SCAN_IN), 
        .Z(n2623) );
  INV_X1 U3361 ( .A(n2623), .ZN(n2624) );
  NOR2_X1 U3362 ( .A1(n2624), .A2(n2650), .ZN(n2891) );
  INV_X1 U3363 ( .A(DATAI_14_), .ZN(n4882) );
  MUX2_X1 U3364 ( .A(n4883), .B(n4882), .S(n2126), .Z(n2625) );
  OR2_X1 U3365 ( .A1(n4602), .A2(n2625), .ZN(n4595) );
  NAND2_X1 U3366 ( .A1(n4602), .A2(n2625), .ZN(n3814) );
  NAND2_X1 U3367 ( .A1(n2626), .A2(n3794), .ZN(n2627) );
  NAND2_X1 U3368 ( .A1(n2187), .A2(n2627), .ZN(n4593) );
  AOI22_X1 U3369 ( .A1(n3803), .A2(REG0_REG_15__SCAN_IN), .B1(n2941), .B2(
        REG2_REG_15__SCAN_IN), .ZN(n2629) );
  INV_X1 U3370 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4672) );
  OR2_X1 U3371 ( .A1(n3806), .A2(n4672), .ZN(n2628) );
  OR2_X1 U3372 ( .A1(n2650), .A2(n2923), .ZN(n2632) );
  INV_X1 U3373 ( .A(n2632), .ZN(n2630) );
  NAND2_X1 U3374 ( .A1(n2630), .A2(IR_REG_15__SCAN_IN), .ZN(n2633) );
  INV_X1 U3375 ( .A(IR_REG_15__SCAN_IN), .ZN(n2631) );
  NAND2_X1 U3376 ( .A1(n2632), .A2(n2631), .ZN(n2639) );
  MUX2_X1 U3377 ( .A(n3997), .B(DATAI_15_), .S(n2125), .Z(n4600) );
  INV_X1 U3378 ( .A(n4580), .ZN(n3692) );
  INV_X1 U3379 ( .A(n4600), .ZN(n3795) );
  XNOR2_X1 U3380 ( .A(n2187), .B(REG3_REG_16__SCAN_IN), .ZN(n4575) );
  NAND2_X1 U3381 ( .A1(n4575), .A2(n2789), .ZN(n2638) );
  INV_X1 U3382 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4666) );
  NAND2_X1 U3383 ( .A1(n3803), .A2(REG0_REG_16__SCAN_IN), .ZN(n2635) );
  NAND2_X1 U3384 ( .A1(n2941), .A2(REG2_REG_16__SCAN_IN), .ZN(n2634) );
  OAI211_X1 U3385 ( .C1(n4666), .C2(n3806), .A(n2635), .B(n2634), .ZN(n2636)
         );
  INV_X1 U3386 ( .A(n2636), .ZN(n2637) );
  NAND2_X1 U3387 ( .A1(n2639), .A2(IR_REG_31__SCAN_IN), .ZN(n2640) );
  XNOR2_X1 U3388 ( .A(n2640), .B(IR_REG_16__SCAN_IN), .ZN(n2894) );
  INV_X1 U3389 ( .A(DATAI_16_), .ZN(n2641) );
  MUX2_X1 U3390 ( .A(n4881), .B(n2641), .S(n2125), .Z(n2825) );
  OR2_X1 U3391 ( .A1(n4561), .A2(n2825), .ZN(n3920) );
  NAND2_X1 U3392 ( .A1(n4561), .A2(n2825), .ZN(n3813) );
  NAND2_X1 U3393 ( .A1(n3920), .A2(n3813), .ZN(n4577) );
  INV_X1 U3394 ( .A(n2825), .ZN(n4579) );
  AOI22_X1 U3395 ( .A1(n4570), .A2(n4577), .B1(n4579), .B2(n4561), .ZN(n4552)
         );
  AOI21_X1 U3396 ( .B1(n2201), .B2(REG3_REG_16__SCAN_IN), .A(
        REG3_REG_17__SCAN_IN), .ZN(n2643) );
  OR2_X1 U3397 ( .A1(n2643), .A2(n2656), .ZN(n3706) );
  INV_X1 U3398 ( .A(n3706), .ZN(n4556) );
  NAND2_X1 U3399 ( .A1(n4556), .A2(n2789), .ZN(n2648) );
  INV_X1 U3400 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4663) );
  NAND2_X1 U3401 ( .A1(n2941), .A2(REG2_REG_17__SCAN_IN), .ZN(n2645) );
  NAND2_X1 U3402 ( .A1(n3803), .A2(REG0_REG_17__SCAN_IN), .ZN(n2644) );
  OAI211_X1 U3403 ( .C1(n3806), .C2(n4663), .A(n2645), .B(n2644), .ZN(n2646)
         );
  INV_X1 U3404 ( .A(n2646), .ZN(n2647) );
  NOR2_X1 U3405 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2649)
         );
  NAND2_X1 U3406 ( .A1(n2650), .A2(n2649), .ZN(n2652) );
  NAND2_X1 U3407 ( .A1(n2652), .A2(IR_REG_31__SCAN_IN), .ZN(n2651) );
  MUX2_X1 U3408 ( .A(IR_REG_31__SCAN_IN), .B(n2651), .S(IR_REG_17__SCAN_IN), 
        .Z(n2653) );
  INV_X1 U3409 ( .A(DATAI_17_), .ZN(n4879) );
  MUX2_X1 U3410 ( .A(n4880), .B(n4879), .S(n2125), .Z(n4564) );
  NAND2_X1 U3411 ( .A1(n4552), .A2(n2177), .ZN(n2655) );
  NAND2_X1 U3412 ( .A1(n2655), .A2(n2654), .ZN(n4533) );
  NOR2_X1 U3413 ( .A1(n2656), .A2(REG3_REG_18__SCAN_IN), .ZN(n2657) );
  OR2_X1 U3414 ( .A1(n2658), .A2(n2657), .ZN(n4537) );
  INV_X1 U3415 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4661) );
  NAND2_X1 U3416 ( .A1(n2941), .A2(REG2_REG_18__SCAN_IN), .ZN(n2660) );
  NAND2_X1 U3417 ( .A1(n3803), .A2(REG0_REG_18__SCAN_IN), .ZN(n2659) );
  OAI211_X1 U3418 ( .C1(n3806), .C2(n4661), .A(n2660), .B(n2659), .ZN(n2661)
         );
  INV_X1 U3419 ( .A(n2661), .ZN(n2662) );
  NAND2_X1 U3420 ( .A1(n2663), .A2(IR_REG_31__SCAN_IN), .ZN(n2665) );
  XNOR2_X1 U3421 ( .A(n2665), .B(n2664), .ZN(n2905) );
  INV_X1 U3422 ( .A(DATAI_18_), .ZN(n4327) );
  MUX2_X1 U3423 ( .A(n2905), .B(n4327), .S(n2125), .Z(n4544) );
  OR2_X1 U3424 ( .A1(n4560), .A2(n4544), .ZN(n4520) );
  NAND2_X1 U3425 ( .A1(n4560), .A2(n4544), .ZN(n4521) );
  NAND2_X1 U3426 ( .A1(n4520), .A2(n4521), .ZN(n4540) );
  INV_X1 U3427 ( .A(n4560), .ZN(n3705) );
  OR2_X2 U3428 ( .A1(n2668), .A2(n3727), .ZN(n2688) );
  NAND2_X1 U3429 ( .A1(n2668), .A2(n3727), .ZN(n2669) );
  NAND2_X1 U3430 ( .A1(n2688), .A2(n2669), .ZN(n4506) );
  INV_X1 U3431 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4654) );
  NAND2_X1 U3432 ( .A1(n3803), .A2(REG0_REG_20__SCAN_IN), .ZN(n2671) );
  NAND2_X1 U3433 ( .A1(n2941), .A2(REG2_REG_20__SCAN_IN), .ZN(n2670) );
  OAI211_X1 U3434 ( .C1(n4654), .C2(n3806), .A(n2671), .B(n2670), .ZN(n2672)
         );
  INV_X1 U3435 ( .A(n2672), .ZN(n2673) );
  NAND2_X1 U3436 ( .A1(n2126), .A2(DATAI_20_), .ZN(n4504) );
  NAND2_X1 U3437 ( .A1(n4527), .A2(n4504), .ZN(n2675) );
  XNOR2_X1 U3438 ( .A(n2688), .B(REG3_REG_21__SCAN_IN), .ZN(n4477) );
  NAND2_X1 U3439 ( .A1(n4477), .A2(n2789), .ZN(n2680) );
  INV_X1 U3440 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4648) );
  NAND2_X1 U3441 ( .A1(n3803), .A2(REG0_REG_21__SCAN_IN), .ZN(n2677) );
  NAND2_X1 U3442 ( .A1(n2941), .A2(REG2_REG_21__SCAN_IN), .ZN(n2676) );
  OAI211_X1 U3443 ( .C1(n4648), .C2(n3806), .A(n2677), .B(n2676), .ZN(n2678)
         );
  INV_X1 U3444 ( .A(n2678), .ZN(n2679) );
  NAND2_X1 U3445 ( .A1(n2126), .A2(DATAI_21_), .ZN(n3568) );
  NAND2_X1 U3446 ( .A1(REG3_REG_21__SCAN_IN), .A2(REG3_REG_22__SCAN_IN), .ZN(
        n2681) );
  NOR2_X4 U3447 ( .A1(n2690), .A2(n3649), .ZN(n2702) );
  AND2_X1 U3448 ( .A1(n2690), .A2(n3649), .ZN(n2682) );
  NOR2_X1 U3449 ( .A1(n2702), .A2(n2682), .ZN(n4442) );
  NAND2_X1 U3450 ( .A1(n4442), .A2(n2789), .ZN(n2687) );
  INV_X1 U3451 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4337) );
  NAND2_X1 U3452 ( .A1(n2941), .A2(REG2_REG_23__SCAN_IN), .ZN(n2684) );
  NAND2_X1 U3453 ( .A1(n3803), .A2(REG0_REG_23__SCAN_IN), .ZN(n2683) );
  OAI211_X1 U3454 ( .C1(n3806), .C2(n4337), .A(n2684), .B(n2683), .ZN(n2685)
         );
  INV_X1 U3455 ( .A(n2685), .ZN(n2686) );
  NAND2_X1 U3456 ( .A1(n2125), .A2(DATAI_23_), .ZN(n4449) );
  NAND2_X1 U3457 ( .A1(n4465), .A2(n4449), .ZN(n2696) );
  INV_X1 U34580 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3665) );
  INV_X1 U34590 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3747) );
  OAI21_X1 U3460 ( .B1(n2688), .B2(n3665), .A(n3747), .ZN(n2689) );
  AND2_X1 U3461 ( .A1(n2690), .A2(n2689), .ZN(n4470) );
  NAND2_X1 U3462 ( .A1(n4470), .A2(n2789), .ZN(n2695) );
  INV_X1 U3463 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4646) );
  NAND2_X1 U3464 ( .A1(n2941), .A2(REG2_REG_22__SCAN_IN), .ZN(n2692) );
  NAND2_X1 U3465 ( .A1(n3803), .A2(REG0_REG_22__SCAN_IN), .ZN(n2691) );
  OAI211_X1 U3466 ( .C1(n3806), .C2(n4646), .A(n2692), .B(n2691), .ZN(n2693)
         );
  INV_X1 U34670 ( .A(n2693), .ZN(n2694) );
  NAND2_X1 U3468 ( .A1(n4483), .A2(n4462), .ZN(n4445) );
  NAND2_X1 U34690 ( .A1(n3664), .A2(n4469), .ZN(n2774) );
  NAND2_X1 U3470 ( .A1(n4445), .A2(n2774), .ZN(n4456) );
  NAND3_X1 U34710 ( .A1(n4436), .A2(n2696), .A3(n4456), .ZN(n2701) );
  INV_X1 U3472 ( .A(n2696), .ZN(n2698) );
  NAND2_X1 U34730 ( .A1(n3664), .A2(n4462), .ZN(n4437) );
  NAND2_X1 U3474 ( .A1(n3957), .A2(n2369), .ZN(n2697) );
  AND2_X2 U34750 ( .A1(n2702), .A2(REG3_REG_24__SCAN_IN), .ZN(n2710) );
  NOR2_X1 U3476 ( .A1(n2702), .A2(REG3_REG_24__SCAN_IN), .ZN(n2703) );
  OR2_X1 U34770 ( .A1(n2710), .A2(n2703), .ZN(n3715) );
  NAND2_X1 U3478 ( .A1(n4140), .A2(n2789), .ZN(n2708) );
  INV_X1 U34790 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4637) );
  NAND2_X1 U3480 ( .A1(n2941), .A2(REG2_REG_24__SCAN_IN), .ZN(n2705) );
  NAND2_X1 U34810 ( .A1(n3803), .A2(REG0_REG_24__SCAN_IN), .ZN(n2704) );
  OAI211_X1 U3482 ( .C1(n3806), .C2(n4637), .A(n2705), .B(n2704), .ZN(n2706)
         );
  INV_X1 U34830 ( .A(n2706), .ZN(n2707) );
  NAND2_X1 U3484 ( .A1(n2126), .A2(DATAI_24_), .ZN(n4135) );
  NOR2_X1 U34850 ( .A1(n4448), .A2(n4135), .ZN(n2709) );
  AND2_X2 U3486 ( .A1(n2710), .A2(REG3_REG_25__SCAN_IN), .ZN(n2718) );
  NOR2_X1 U34870 ( .A1(n2710), .A2(REG3_REG_25__SCAN_IN), .ZN(n2711) );
  INV_X1 U3488 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4322) );
  NAND2_X1 U34890 ( .A1(n3803), .A2(REG0_REG_25__SCAN_IN), .ZN(n2713) );
  NAND2_X1 U3490 ( .A1(n2941), .A2(REG2_REG_25__SCAN_IN), .ZN(n2712) );
  OAI211_X1 U34910 ( .C1(n4322), .C2(n3806), .A(n2713), .B(n2712), .ZN(n2714)
         );
  INV_X1 U3492 ( .A(n2714), .ZN(n2715) );
  OAI21_X2 U34930 ( .B1(n3674), .B2(n2716), .A(n2715), .ZN(n4137) );
  AND2_X1 U3494 ( .A1(n2125), .A2(DATAI_25_), .ZN(n4113) );
  NOR2_X1 U34950 ( .A1(n4137), .A2(n4113), .ZN(n2717) );
  INV_X1 U3496 ( .A(n4137), .ZN(n3781) );
  OR2_X1 U34970 ( .A1(n2718), .A2(REG3_REG_26__SCAN_IN), .ZN(n2719) );
  NAND2_X2 U3498 ( .A1(n2718), .A2(REG3_REG_26__SCAN_IN), .ZN(n2734) );
  NAND2_X1 U34990 ( .A1(n4105), .A2(n2789), .ZN(n2724) );
  INV_X1 U3500 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4630) );
  NAND2_X1 U35010 ( .A1(n2941), .A2(REG2_REG_26__SCAN_IN), .ZN(n2721) );
  NAND2_X1 U3502 ( .A1(n3803), .A2(REG0_REG_26__SCAN_IN), .ZN(n2720) );
  OAI211_X1 U35030 ( .C1(n3806), .C2(n4630), .A(n2721), .B(n2720), .ZN(n2722)
         );
  INV_X1 U3504 ( .A(n2722), .ZN(n2723) );
  AND2_X2 U35050 ( .A1(n2724), .A2(n2723), .ZN(n4119) );
  NAND2_X1 U35060 ( .A1(n2126), .A2(DATAI_26_), .ZN(n4099) );
  NOR2_X1 U35070 ( .A1(n4119), .A2(n4099), .ZN(n2725) );
  INV_X1 U35080 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4306) );
  NAND2_X1 U35090 ( .A1(n2941), .A2(REG2_REG_27__SCAN_IN), .ZN(n2727) );
  NAND2_X1 U35100 ( .A1(n3803), .A2(REG0_REG_27__SCAN_IN), .ZN(n2726) );
  OAI211_X1 U35110 ( .C1(n3806), .C2(n4306), .A(n2727), .B(n2726), .ZN(n2728)
         );
  INV_X1 U35120 ( .A(n2728), .ZN(n2729) );
  NAND2_X2 U35130 ( .A1(n2730), .A2(n2729), .ZN(n4098) );
  NAND2_X1 U35140 ( .A1(n2125), .A2(DATAI_27_), .ZN(n4077) );
  INV_X1 U35150 ( .A(n4077), .ZN(n3607) );
  INV_X1 U35160 ( .A(n4098), .ZN(n2731) );
  INV_X1 U35170 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3603) );
  INV_X1 U35180 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2732) );
  OAI21_X1 U35190 ( .B1(n2734), .B2(n3603), .A(n2732), .ZN(n2735) );
  NAND2_X1 U35200 ( .A1(REG3_REG_27__SCAN_IN), .A2(REG3_REG_28__SCAN_IN), .ZN(
        n2733) );
  OR2_X2 U35210 ( .A1(n2734), .A2(n2733), .ZN(n4054) );
  INV_X1 U35220 ( .A(REG1_REG_28__SCAN_IN), .ZN(n4313) );
  NAND2_X1 U35230 ( .A1(n3803), .A2(REG0_REG_28__SCAN_IN), .ZN(n2737) );
  NAND2_X1 U35240 ( .A1(n2941), .A2(REG2_REG_28__SCAN_IN), .ZN(n2736) );
  OAI211_X1 U35250 ( .C1(n4313), .C2(n3806), .A(n2737), .B(n2736), .ZN(n2738)
         );
  INV_X1 U35260 ( .A(n2738), .ZN(n2739) );
  AND2_X2 U35270 ( .A1(n2740), .A2(n2739), .ZN(n4074) );
  AND2_X1 U35280 ( .A1(n2125), .A2(DATAI_28_), .ZN(n4030) );
  NAND2_X1 U35290 ( .A1(n4074), .A2(n4030), .ZN(n4041) );
  INV_X1 U35300 ( .A(n4030), .ZN(n3614) );
  NAND2_X1 U35310 ( .A1(n4051), .A2(n3614), .ZN(n4039) );
  XNOR2_X1 U35320 ( .A(n4032), .B(n4029), .ZN(n4058) );
  NAND2_X1 U35330 ( .A1(n2742), .A2(n2741), .ZN(n2743) );
  XNOR2_X2 U35340 ( .A(n2745), .B(n2744), .ZN(n2828) );
  BUF_X1 U35350 ( .A(n2746), .Z(n2747) );
  NAND2_X2 U35360 ( .A1(n2828), .A2(n3941), .ZN(n3084) );
  NAND2_X1 U35370 ( .A1(n2805), .A2(IR_REG_31__SCAN_IN), .ZN(n2751) );
  XNOR2_X1 U35380 ( .A(n3084), .B(n3950), .ZN(n2752) );
  NAND2_X1 U35390 ( .A1(n2752), .A2(n4012), .ZN(n4502) );
  NAND2_X1 U35400 ( .A1(n2828), .A2(n4004), .ZN(n3078) );
  INV_X1 U35410 ( .A(n3226), .ZN(n2754) );
  NAND2_X1 U35420 ( .A1(n2754), .A2(n3189), .ZN(n3819) );
  NAND2_X1 U35430 ( .A1(n3059), .A2(n3254), .ZN(n3830) );
  NAND2_X1 U35440 ( .A1(n3963), .A2(n3245), .ZN(n3827) );
  AND2_X1 U35450 ( .A1(n3830), .A2(n3827), .ZN(n3243) );
  INV_X1 U35460 ( .A(n3830), .ZN(n2756) );
  AOI21_X1 U35470 ( .B1(n3244), .B2(n3243), .A(n2756), .ZN(n3099) );
  NAND2_X1 U35480 ( .A1(n3099), .A2(n3831), .ZN(n2757) );
  NAND2_X1 U35490 ( .A1(n2757), .A2(n3834), .ZN(n3135) );
  AND2_X1 U35500 ( .A1(n3152), .A2(n2824), .ZN(n3134) );
  NAND2_X1 U35510 ( .A1(n3218), .A2(n3211), .ZN(n3847) );
  NAND2_X1 U35520 ( .A1(n3961), .A2(n2363), .ZN(n3845) );
  INV_X1 U35530 ( .A(n3961), .ZN(n3195) );
  NAND2_X1 U35540 ( .A1(n3195), .A2(n3220), .ZN(n3836) );
  INV_X1 U35550 ( .A(n2758), .ZN(n2759) );
  INV_X1 U35560 ( .A(n3263), .ZN(n3369) );
  NAND2_X1 U35570 ( .A1(n3369), .A2(n3332), .ZN(n3840) );
  NAND2_X1 U35580 ( .A1(n3263), .A2(n3325), .ZN(n3838) );
  INV_X1 U35590 ( .A(n3373), .ZN(n3358) );
  AND2_X1 U35600 ( .A1(n3959), .A2(n3358), .ZN(n3849) );
  INV_X1 U35610 ( .A(n3959), .ZN(n3359) );
  NAND2_X1 U35620 ( .A1(n3359), .A2(n3373), .ZN(n3841) );
  NAND2_X1 U35630 ( .A1(n3429), .A2(n3415), .ZN(n3816) );
  NAND2_X1 U35640 ( .A1(n3342), .A2(n3816), .ZN(n2760) );
  NAND2_X1 U35650 ( .A1(n3443), .A2(n3419), .ZN(n3844) );
  INV_X1 U35660 ( .A(n3738), .ZN(n2954) );
  NAND2_X1 U35670 ( .A1(n3454), .A2(n2954), .ZN(n3477) );
  INV_X1 U35680 ( .A(n3740), .ZN(n3472) );
  NAND2_X1 U35690 ( .A1(n3636), .A2(n3472), .ZN(n3473) );
  NAND2_X1 U35700 ( .A1(n3477), .A2(n3473), .ZN(n2761) );
  INV_X1 U35710 ( .A(n3454), .ZN(n3459) );
  NAND2_X1 U35720 ( .A1(n3459), .A2(n3738), .ZN(n3476) );
  NAND2_X1 U35730 ( .A1(n3476), .A2(n3403), .ZN(n2762) );
  INV_X1 U35740 ( .A(n2761), .ZN(n3818) );
  NOR2_X1 U35750 ( .A1(n3636), .A2(n3472), .ZN(n3474) );
  AOI21_X1 U35760 ( .B1(n2762), .B2(n3818), .A(n3474), .ZN(n3853) );
  OR2_X1 U35770 ( .A1(n4580), .A2(n3795), .ZN(n3852) );
  NAND2_X1 U35780 ( .A1(n4580), .A2(n3795), .ZN(n3815) );
  NAND2_X1 U35790 ( .A1(n3852), .A2(n3815), .ZN(n4597) );
  INV_X1 U35800 ( .A(n4595), .ZN(n2763) );
  NOR2_X1 U35810 ( .A1(n4597), .A2(n2763), .ZN(n2764) );
  NAND2_X1 U3582 ( .A1(n4596), .A2(n2764), .ZN(n2765) );
  NAND2_X1 U3583 ( .A1(n2765), .A2(n3815), .ZN(n4578) );
  INV_X1 U3584 ( .A(n4577), .ZN(n3895) );
  NAND2_X1 U3585 ( .A1(n4547), .A2(n3880), .ZN(n2767) );
  NAND2_X1 U3586 ( .A1(n2767), .A2(n4521), .ZN(n2768) );
  AND2_X1 U3587 ( .A1(n3691), .A2(n4564), .ZN(n4516) );
  NOR2_X1 U3588 ( .A1(n2768), .A2(n4516), .ZN(n4492) );
  NAND2_X1 U3589 ( .A1(n4481), .A2(n4504), .ZN(n3922) );
  NAND2_X1 U3590 ( .A1(n4492), .A2(n3922), .ZN(n3812) );
  INV_X1 U3591 ( .A(n2768), .ZN(n2770) );
  OR2_X1 U3592 ( .A1(n3691), .A2(n4564), .ZN(n4518) );
  NAND2_X1 U3593 ( .A1(n4520), .A2(n4518), .ZN(n2769) );
  NAND2_X1 U3594 ( .A1(n2770), .A2(n2769), .ZN(n2772) );
  NAND2_X1 U3595 ( .A1(n4490), .A2(n4525), .ZN(n2771) );
  NAND2_X1 U3596 ( .A1(n2772), .A2(n2771), .ZN(n4491) );
  NOR2_X1 U3597 ( .A1(n4481), .A2(n4504), .ZN(n2773) );
  OR2_X1 U3598 ( .A1(n4491), .A2(n2773), .ZN(n3923) );
  OR2_X1 U3599 ( .A1(n4500), .A2(n3568), .ZN(n4443) );
  AND2_X1 U3600 ( .A1(n4445), .A2(n4443), .ZN(n3925) );
  NAND2_X1 U3601 ( .A1(n3957), .A2(n4449), .ZN(n3883) );
  NAND2_X1 U3602 ( .A1(n3883), .A2(n2774), .ZN(n3867) );
  AND2_X1 U3603 ( .A1(n4500), .A2(n3568), .ZN(n4444) );
  AND2_X1 U3604 ( .A1(n4445), .A2(n4444), .ZN(n2775) );
  NOR2_X1 U3605 ( .A1(n3867), .A2(n2775), .ZN(n3928) );
  NAND2_X1 U3606 ( .A1(n2776), .A2(n3928), .ZN(n4132) );
  OR2_X1 U3607 ( .A1(n3956), .A2(n4135), .ZN(n3878) );
  OR2_X1 U3608 ( .A1(n3957), .A2(n4449), .ZN(n4131) );
  NAND2_X1 U3609 ( .A1(n3878), .A2(n4131), .ZN(n3927) );
  INV_X1 U3610 ( .A(n3927), .ZN(n3865) );
  NAND2_X1 U3611 ( .A1(n4119), .A2(n4088), .ZN(n3885) );
  OR2_X1 U3612 ( .A1(n4137), .A2(n4120), .ZN(n4093) );
  INV_X1 U3613 ( .A(n3931), .ZN(n2777) );
  NAND2_X1 U3614 ( .A1(n4137), .A2(n4120), .ZN(n3887) );
  NAND2_X1 U3615 ( .A1(n3956), .A2(n4135), .ZN(n4115) );
  NAND2_X1 U3616 ( .A1(n3887), .A2(n4115), .ZN(n4091) );
  INV_X1 U3617 ( .A(n4119), .ZN(n3955) );
  AND2_X1 U3618 ( .A1(n3955), .A2(n4099), .ZN(n3915) );
  AOI21_X1 U3619 ( .B1(n3931), .B2(n4091), .A(n3915), .ZN(n3871) );
  NAND2_X1 U3620 ( .A1(n4098), .A2(n4077), .ZN(n3869) );
  XOR2_X1 U3621 ( .A(n4029), .B(n4040), .Z(n2795) );
  NAND2_X1 U3622 ( .A1(n3950), .A2(n4004), .ZN(n2779) );
  INV_X1 U3623 ( .A(n2828), .ZN(n3944) );
  NAND2_X1 U3624 ( .A1(n3944), .A2(n2127), .ZN(n2778) );
  NAND3_X1 U3625 ( .A1(n2780), .A2(n2782), .A3(n2781), .ZN(n2783) );
  NAND2_X1 U3626 ( .A1(n2783), .A2(IR_REG_31__SCAN_IN), .ZN(n2784) );
  XNOR2_X1 U3627 ( .A(n2784), .B(n4160), .ZN(n4783) );
  INV_X1 U3628 ( .A(n4783), .ZN(n3067) );
  INV_X1 U3629 ( .A(n4054), .ZN(n2790) );
  INV_X1 U3630 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2787) );
  NAND2_X1 U3631 ( .A1(n3803), .A2(REG0_REG_29__SCAN_IN), .ZN(n2786) );
  NAND2_X1 U3632 ( .A1(n2941), .A2(REG2_REG_29__SCAN_IN), .ZN(n2785) );
  OAI211_X1 U3633 ( .C1(n3806), .C2(n2787), .A(n2786), .B(n2785), .ZN(n2788)
         );
  AOI21_X1 U3634 ( .B1(n2790), .B2(n2789), .A(n2788), .ZN(n3877) );
  NAND2_X1 U3635 ( .A1(n3046), .A2(n4783), .ZN(n4604) );
  INV_X1 U3636 ( .A(n3950), .ZN(n2792) );
  INV_X1 U3637 ( .A(n3941), .ZN(n2791) );
  OAI22_X1 U3638 ( .A1(n3877), .A2(n4604), .B1(n3614), .B2(n4565), .ZN(n2793)
         );
  AOI21_X1 U3639 ( .B1(n4601), .B2(n4098), .A(n2793), .ZN(n2794) );
  OAI21_X1 U3640 ( .B1(n2795), .B2(n4496), .A(n2794), .ZN(n4063) );
  AOI21_X1 U3641 ( .B1(n4058), .B2(n4928), .A(n4063), .ZN(n2837) );
  NOR4_X1 U3642 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_12__SCAN_IN), .A3(
        D_REG_13__SCAN_IN), .A4(D_REG_19__SCAN_IN), .ZN(n2799) );
  NOR4_X1 U3643 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_4__SCAN_IN), .A3(
        D_REG_2__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n2798) );
  INV_X1 U3644 ( .A(D_REG_15__SCAN_IN), .ZN(n4869) );
  INV_X1 U3645 ( .A(D_REG_21__SCAN_IN), .ZN(n4866) );
  INV_X1 U3646 ( .A(D_REG_22__SCAN_IN), .ZN(n4865) );
  INV_X1 U3647 ( .A(D_REG_18__SCAN_IN), .ZN(n4867) );
  NAND4_X1 U3648 ( .A1(n4869), .A2(n4866), .A3(n4865), .A4(n4867), .ZN(n2796)
         );
  NOR2_X1 U3649 ( .A1(D_REG_31__SCAN_IN), .A2(n2796), .ZN(n4187) );
  NOR4_X1 U3650 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_20__SCAN_IN), .A3(
        D_REG_14__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n2797) );
  NAND4_X1 U3651 ( .A1(n2799), .A2(n2798), .A3(n4187), .A4(n2797), .ZN(n2804)
         );
  NOR4_X1 U3652 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(
        D_REG_10__SCAN_IN), .A4(D_REG_6__SCAN_IN), .ZN(n2802) );
  NOR4_X1 U3653 ( .A1(D_REG_25__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_16__SCAN_IN), .A4(D_REG_9__SCAN_IN), .ZN(n2801) );
  NOR4_X1 U3654 ( .A1(D_REG_30__SCAN_IN), .A2(D_REG_24__SCAN_IN), .A3(
        D_REG_5__SCAN_IN), .A4(D_REG_3__SCAN_IN), .ZN(n2800) );
  INV_X1 U3655 ( .A(D_REG_23__SCAN_IN), .ZN(n4864) );
  NAND4_X1 U3656 ( .A1(n2802), .A2(n2801), .A3(n2800), .A4(n4864), .ZN(n2803)
         );
  NOR2_X1 U3657 ( .A1(n2804), .A2(n2803), .ZN(n3040) );
  INV_X1 U3658 ( .A(IR_REG_22__SCAN_IN), .ZN(n2806) );
  NAND2_X1 U3659 ( .A1(n2819), .A2(n2820), .ZN(n2807) );
  INV_X1 U3660 ( .A(n2809), .ZN(n2810) );
  NAND2_X1 U3661 ( .A1(n2808), .A2(n2817), .ZN(n2814) );
  MUX2_X1 U3662 ( .A(n2808), .B(n2814), .S(B_REG_SCAN_IN), .Z(n2816) );
  XNOR2_X2 U3663 ( .A(n2815), .B(IR_REG_26__SCAN_IN), .ZN(n4773) );
  XNOR2_X1 U3664 ( .A(n2819), .B(n2820), .ZN(n2854) );
  NAND2_X1 U3665 ( .A1(n2828), .A2(n4012), .ZN(n3045) );
  AND2_X1 U3666 ( .A1(n3046), .A2(n3045), .ZN(n3063) );
  NOR2_X1 U3667 ( .A1(n4894), .A2(n2127), .ZN(n3051) );
  NOR2_X1 U3668 ( .A1(n3074), .A2(n3051), .ZN(n2822) );
  INV_X1 U3669 ( .A(n4773), .ZN(n3501) );
  NAND2_X1 U3670 ( .A1(n2817), .A2(n3501), .ZN(n2933) );
  OAI21_X1 U3671 ( .B1(n3039), .B2(D_REG_1__SCAN_IN), .A(n2933), .ZN(n2821) );
  OAI211_X1 U3672 ( .C1(n3040), .C2(n3039), .A(n2822), .B(n2821), .ZN(n2832)
         );
  INV_X1 U3673 ( .A(n2832), .ZN(n2823) );
  INV_X1 U3674 ( .A(n3189), .ZN(n3080) );
  NAND2_X1 U3675 ( .A1(n3293), .A2(n3292), .ZN(n3291) );
  NAND2_X1 U3676 ( .A1(n3313), .A2(n3325), .ZN(n3314) );
  OR2_X2 U3677 ( .A1(n3314), .A2(n3373), .ZN(n3347) );
  NOR2_X4 U3678 ( .A1(n3347), .A2(n3419), .ZN(n3381) );
  INV_X1 U3679 ( .A(n4079), .ZN(n2826) );
  OAI21_X1 U3680 ( .B1(n2826), .B2(n3614), .A(n4035), .ZN(n4061) );
  AND2_X2 U3681 ( .A1(n3079), .A2(n2828), .ZN(n4924) );
  NAND2_X1 U3682 ( .A1(n4932), .A2(n4924), .ZN(n4766) );
  OR2_X1 U3683 ( .A1(n4061), .A2(n4766), .ZN(n2830) );
  INV_X1 U3684 ( .A(REG0_REG_28__SCAN_IN), .ZN(n4312) );
  OAI21_X1 U3685 ( .B1(n2837), .B2(n4930), .A(n2831), .ZN(U3514) );
  INV_X1 U3686 ( .A(n4941), .ZN(n2836) );
  NAND2_X1 U3687 ( .A1(n2836), .A2(REG1_REG_28__SCAN_IN), .ZN(n2833) );
  OAI21_X1 U3688 ( .B1(n2837), .B2(n2836), .A(n2835), .ZN(U3546) );
  INV_X2 U3689 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  XNOR2_X1 U3690 ( .A(n2905), .B(REG1_REG_18__SCAN_IN), .ZN(n4002) );
  INV_X1 U3691 ( .A(n4779), .ZN(n2843) );
  MUX2_X1 U3692 ( .A(REG1_REG_2__SCAN_IN), .B(n2840), .S(n2373), .Z(n2973) );
  NAND2_X1 U3693 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n4164) );
  INV_X1 U3694 ( .A(n4164), .ZN(n3969) );
  OAI21_X1 U3695 ( .B1(n3965), .B2(n2838), .A(n3968), .ZN(n2972) );
  INV_X1 U3696 ( .A(n2869), .ZN(n2986) );
  NAND2_X1 U3697 ( .A1(n2990), .A2(REG1_REG_4__SCAN_IN), .ZN(n2989) );
  MUX2_X1 U3698 ( .A(REG1_REG_5__SCAN_IN), .B(n2842), .S(n4779), .Z(n3978) );
  INV_X1 U3699 ( .A(n3004), .ZN(n3008) );
  INV_X1 U3700 ( .A(n4778), .ZN(n3115) );
  XOR2_X1 U3701 ( .A(REG1_REG_9__SCAN_IN), .B(n4777), .Z(n3231) );
  INV_X1 U3702 ( .A(n2846), .ZN(n2847) );
  XOR2_X1 U3703 ( .A(REG1_REG_11__SCAN_IN), .B(n4776), .Z(n3393) );
  INV_X1 U3704 ( .A(n4886), .ZN(n2886) );
  NAND2_X1 U3705 ( .A1(n2849), .A2(n2886), .ZN(n2850) );
  INV_X1 U3706 ( .A(n2889), .ZN(n4885) );
  AOI22_X1 U3707 ( .A1(n2889), .A2(REG1_REG_13__SCAN_IN), .B1(n4222), .B2(
        n4885), .ZN(n4820) );
  XNOR2_X1 U3708 ( .A(n3997), .B(REG1_REG_15__SCAN_IN), .ZN(n3990) );
  INV_X1 U3709 ( .A(n3997), .ZN(n2930) );
  NOR2_X1 U3710 ( .A1(n2894), .A2(n2852), .ZN(n2853) );
  AOI22_X1 U3711 ( .A1(REG1_REG_17__SCAN_IN), .A2(n4880), .B1(n2896), .B2(
        n4663), .ZN(n4853) );
  INV_X1 U3712 ( .A(n2854), .ZN(n3062) );
  NAND2_X1 U3713 ( .A1(n3062), .A2(STATE_REG_SCAN_IN), .ZN(n3953) );
  NAND2_X1 U3714 ( .A1(n3052), .A2(n3953), .ZN(n2860) );
  NAND2_X1 U3715 ( .A1(n3046), .A2(n2854), .ZN(n2855) );
  AND2_X1 U3716 ( .A1(n2855), .A2(n2125), .ZN(n2858) );
  NAND2_X1 U3717 ( .A1(n2860), .A2(n2858), .ZN(n4791) );
  XNOR2_X1 U3718 ( .A(n2856), .B(IR_REG_27__SCAN_IN), .ZN(n4784) );
  NAND2_X1 U3719 ( .A1(n2857), .A2(n4852), .ZN(n2907) );
  INV_X1 U3720 ( .A(n2858), .ZN(n2859) );
  INV_X1 U3721 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4205) );
  AOI22_X1 U3722 ( .A1(REG2_REG_17__SCAN_IN), .A2(n2896), .B1(n4880), .B2(
        n4205), .ZN(n4848) );
  NOR2_X1 U3723 ( .A1(n4885), .A2(n2612), .ZN(n4812) );
  INV_X1 U3724 ( .A(REG2_REG_11__SCAN_IN), .ZN(n2885) );
  INV_X1 U3725 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3272) );
  INV_X1 U3726 ( .A(n4777), .ZN(n2881) );
  AND2_X1 U3727 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n2861)
         );
  NAND2_X1 U3728 ( .A1(n3973), .A2(n2861), .ZN(n3972) );
  NAND2_X1 U3729 ( .A1(n4781), .A2(REG2_REG_1__SCAN_IN), .ZN(n2974) );
  NAND2_X1 U3730 ( .A1(n3972), .A2(n2974), .ZN(n2863) );
  INV_X1 U3731 ( .A(n2975), .ZN(n2862) );
  NAND2_X1 U3732 ( .A1(n4780), .A2(REG2_REG_2__SCAN_IN), .ZN(n2864) );
  NAND2_X1 U3733 ( .A1(n2866), .A2(n2865), .ZN(n2867) );
  NAND2_X1 U3734 ( .A1(n2868), .A2(n2867), .ZN(n2870) );
  XNOR2_X1 U3735 ( .A(n2870), .B(n2986), .ZN(n2984) );
  NAND2_X1 U3736 ( .A1(n2984), .A2(REG2_REG_4__SCAN_IN), .ZN(n2872) );
  NAND2_X1 U3737 ( .A1(n2870), .A2(n2869), .ZN(n2871) );
  NAND2_X1 U3738 ( .A1(n2872), .A2(n2871), .ZN(n3984) );
  INV_X1 U3739 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3140) );
  MUX2_X1 U3740 ( .A(REG2_REG_5__SCAN_IN), .B(n3140), .S(n4779), .Z(n3985) );
  NAND2_X1 U3741 ( .A1(n3984), .A2(n3985), .ZN(n3983) );
  NAND2_X1 U3742 ( .A1(n4779), .A2(REG2_REG_5__SCAN_IN), .ZN(n2873) );
  INV_X1 U3743 ( .A(n2874), .ZN(n2996) );
  XNOR2_X1 U3744 ( .A(n2875), .B(n2996), .ZN(n2994) );
  NAND2_X1 U3745 ( .A1(n2994), .A2(REG2_REG_6__SCAN_IN), .ZN(n2877) );
  NAND2_X1 U3746 ( .A1(n2875), .A2(n2874), .ZN(n2876) );
  NAND2_X1 U3747 ( .A1(n2877), .A2(n2876), .ZN(n3012) );
  INV_X1 U3748 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2878) );
  MUX2_X1 U3749 ( .A(REG2_REG_7__SCAN_IN), .B(n2878), .S(n3004), .Z(n3011) );
  NAND2_X1 U3750 ( .A1(n3012), .A2(n3011), .ZN(n3010) );
  NAND2_X1 U3751 ( .A1(n3004), .A2(REG2_REG_7__SCAN_IN), .ZN(n2879) );
  MUX2_X1 U3752 ( .A(n3272), .B(REG2_REG_9__SCAN_IN), .S(n4777), .Z(n3236) );
  NAND2_X1 U3753 ( .A1(n2882), .A2(n2883), .ZN(n2884) );
  MUX2_X1 U3754 ( .A(n2885), .B(REG2_REG_11__SCAN_IN), .S(n4776), .Z(n3396) );
  NAND2_X1 U3755 ( .A1(n3397), .A2(n3396), .ZN(n3395) );
  NAND2_X1 U3756 ( .A1(n2887), .A2(n2886), .ZN(n2888) );
  INV_X1 U3757 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4826) );
  NOR2_X2 U3758 ( .A1(n4825), .A2(n4826), .ZN(n4824) );
  NAND2_X1 U3759 ( .A1(n3997), .A2(REG2_REG_15__SCAN_IN), .ZN(n2892) );
  OAI21_X1 U3760 ( .B1(n3997), .B2(REG2_REG_15__SCAN_IN), .A(n2892), .ZN(n3993) );
  INV_X1 U3761 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4834) );
  INV_X1 U3762 ( .A(n2905), .ZN(n4775) );
  INV_X1 U3763 ( .A(REG2_REG_18__SCAN_IN), .ZN(n2898) );
  NOR2_X1 U3764 ( .A1(n4775), .A2(n2898), .ZN(n2897) );
  AOI21_X1 U3765 ( .B1(n4775), .B2(n2898), .A(n2897), .ZN(n2899) );
  NAND2_X1 U3766 ( .A1(n3067), .A2(n4784), .ZN(n3948) );
  NAND2_X1 U3767 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n3768) );
  INV_X1 U3768 ( .A(n4877), .ZN(n2908) );
  INV_X1 U3769 ( .A(DATAI_3_), .ZN(n2909) );
  MUX2_X1 U3770 ( .A(n2245), .B(n2909), .S(U3149), .Z(n2910) );
  INV_X1 U3771 ( .A(n2910), .ZN(U3349) );
  INV_X1 U3772 ( .A(DATAI_4_), .ZN(n2911) );
  MUX2_X1 U3773 ( .A(n2986), .B(n2911), .S(U3149), .Z(n2912) );
  INV_X1 U3774 ( .A(n2912), .ZN(U3348) );
  INV_X1 U3775 ( .A(DATAI_19_), .ZN(n2913) );
  MUX2_X1 U3776 ( .A(n4012), .B(n2913), .S(U3149), .Z(n2914) );
  INV_X1 U3777 ( .A(n2914), .ZN(U3333) );
  INV_X1 U3778 ( .A(DATAI_21_), .ZN(n2916) );
  NAND2_X1 U3779 ( .A1(n2127), .A2(STATE_REG_SCAN_IN), .ZN(n2915) );
  OAI21_X1 U3780 ( .B1(STATE_REG_SCAN_IN), .B2(n2916), .A(n2915), .ZN(U3331)
         );
  INV_X1 U3781 ( .A(DATAI_6_), .ZN(n2917) );
  MUX2_X1 U3782 ( .A(n2917), .B(n2996), .S(STATE_REG_SCAN_IN), .Z(n2918) );
  INV_X1 U3783 ( .A(n2918), .ZN(U3346) );
  INV_X1 U3784 ( .A(DATAI_22_), .ZN(n4246) );
  NAND2_X1 U3785 ( .A1(n3950), .A2(STATE_REG_SCAN_IN), .ZN(n2919) );
  OAI21_X1 U3786 ( .B1(STATE_REG_SCAN_IN), .B2(n4246), .A(n2919), .ZN(U3330)
         );
  INV_X1 U3787 ( .A(DATAI_20_), .ZN(n2921) );
  NAND2_X1 U3788 ( .A1(n3944), .A2(STATE_REG_SCAN_IN), .ZN(n2920) );
  OAI21_X1 U3789 ( .B1(STATE_REG_SCAN_IN), .B2(n2921), .A(n2920), .ZN(U3332)
         );
  INV_X1 U3790 ( .A(DATAI_27_), .ZN(n4230) );
  NAND2_X1 U3791 ( .A1(n4784), .A2(STATE_REG_SCAN_IN), .ZN(n2922) );
  OAI21_X1 U3792 ( .B1(STATE_REG_SCAN_IN), .B2(n4230), .A(n2922), .ZN(U3325)
         );
  INV_X1 U3793 ( .A(DATAI_31_), .ZN(n2926) );
  OR4_X1 U3794 ( .A1(n2924), .A2(IR_REG_30__SCAN_IN), .A3(n2923), .A4(U3149), 
        .ZN(n2925) );
  OAI21_X1 U3795 ( .B1(STATE_REG_SCAN_IN), .B2(n2926), .A(n2925), .ZN(U3321)
         );
  INV_X1 U3796 ( .A(DATAI_7_), .ZN(n2927) );
  MUX2_X1 U3797 ( .A(n2927), .B(n3008), .S(STATE_REG_SCAN_IN), .Z(n2928) );
  INV_X1 U3798 ( .A(n2928), .ZN(U3345) );
  INV_X1 U3799 ( .A(DATAI_15_), .ZN(n2929) );
  MUX2_X1 U3800 ( .A(n2930), .B(n2929), .S(U3149), .Z(n2931) );
  INV_X1 U3801 ( .A(n2931), .ZN(U3337) );
  INV_X1 U3802 ( .A(n3052), .ZN(n2932) );
  INV_X1 U3803 ( .A(D_REG_1__SCAN_IN), .ZN(n4252) );
  INV_X1 U3804 ( .A(n2933), .ZN(n3041) );
  AOI22_X1 U3805 ( .A1(n4876), .A2(n4252), .B1(n3041), .B2(n4877), .ZN(U3459)
         );
  NOR2_X1 U3806 ( .A1(n4851), .A2(U4043), .ZN(U3148) );
  XOR2_X1 U3807 ( .A(n2934), .B(REG2_REG_3__SCAN_IN), .Z(n2938) );
  AOI211_X1 U3808 ( .C1(n2494), .C2(n2936), .A(n2935), .B(n4838), .ZN(n2937)
         );
  AOI21_X1 U3809 ( .B1(n2901), .B2(n2938), .A(n2937), .ZN(n2940) );
  INV_X1 U3810 ( .A(REG3_REG_3__SCAN_IN), .ZN(n4237) );
  NOR2_X1 U3811 ( .A1(STATE_REG_SCAN_IN), .A2(n4237), .ZN(n3092) );
  AOI21_X1 U3812 ( .B1(n4851), .B2(ADDR_REG_3__SCAN_IN), .A(n3092), .ZN(n2939)
         );
  OAI211_X1 U3813 ( .C1(n2245), .C2(n4858), .A(n2940), .B(n2939), .ZN(U3243)
         );
  INV_X1 U3814 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n4320) );
  INV_X1 U3815 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4615) );
  NAND2_X1 U3816 ( .A1(n2941), .A2(REG2_REG_31__SCAN_IN), .ZN(n2943) );
  NAND2_X1 U3817 ( .A1(n3803), .A2(REG0_REG_31__SCAN_IN), .ZN(n2942) );
  OAI211_X1 U3818 ( .C1(n3806), .C2(n4615), .A(n2943), .B(n2942), .ZN(n4019)
         );
  NAND2_X1 U3819 ( .A1(U4043), .A2(n4019), .ZN(n2944) );
  OAI21_X1 U3820 ( .B1(U4043), .B2(n4320), .A(n2944), .ZN(U3581) );
  NAND2_X1 U3821 ( .A1(U4043), .A2(n3226), .ZN(n2945) );
  OAI21_X1 U3822 ( .B1(U4043), .B2(n4172), .A(n2945), .ZN(U3550) );
  INV_X1 U3823 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n4328) );
  NAND2_X1 U3824 ( .A1(U4043), .A2(n3152), .ZN(n2946) );
  OAI21_X1 U3825 ( .B1(U4043), .B2(n4328), .A(n2946), .ZN(U3555) );
  INV_X1 U3826 ( .A(DATAO_REG_10__SCAN_IN), .ZN(n4408) );
  NAND2_X1 U3827 ( .A1(U4043), .A2(n3415), .ZN(n2947) );
  OAI21_X1 U3828 ( .B1(U4043), .B2(n4408), .A(n2947), .ZN(U3560) );
  INV_X1 U3829 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n4256) );
  NAND2_X1 U3830 ( .A1(U4043), .A2(n3263), .ZN(n2948) );
  OAI21_X1 U3831 ( .B1(U4043), .B2(n4256), .A(n2948), .ZN(U3558) );
  INV_X1 U3832 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n4335) );
  NAND2_X1 U3833 ( .A1(n3758), .A2(U4043), .ZN(n2949) );
  OAI21_X1 U3834 ( .B1(n4335), .B2(U4043), .A(n2949), .ZN(U3551) );
  INV_X1 U3835 ( .A(DATAO_REG_4__SCAN_IN), .ZN(n4323) );
  NAND2_X1 U3836 ( .A1(n3136), .A2(U4043), .ZN(n2950) );
  OAI21_X1 U3837 ( .B1(U4043), .B2(n4323), .A(n2950), .ZN(U3554) );
  INV_X1 U3838 ( .A(DATAO_REG_16__SCAN_IN), .ZN(n4402) );
  NAND2_X1 U3839 ( .A1(n4561), .A2(U4043), .ZN(n2951) );
  OAI21_X1 U3840 ( .B1(U4043), .B2(n4402), .A(n2951), .ZN(U3566) );
  INV_X1 U3841 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n4331) );
  NAND2_X1 U3842 ( .A1(n4560), .A2(U4043), .ZN(n2952) );
  OAI21_X1 U3843 ( .B1(U4043), .B2(n4331), .A(n2952), .ZN(U3568) );
  INV_X1 U3844 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n4258) );
  NAND2_X1 U3845 ( .A1(n3691), .A2(U4043), .ZN(n2953) );
  OAI21_X1 U3846 ( .B1(U4043), .B2(n4258), .A(n2953), .ZN(U3567) );
  INV_X1 U3847 ( .A(DATAO_REG_12__SCAN_IN), .ZN(n4264) );
  NAND2_X1 U3848 ( .A1(n2954), .A2(U4043), .ZN(n2955) );
  OAI21_X1 U3849 ( .B1(U4043), .B2(n4264), .A(n2955), .ZN(U3562) );
  INV_X1 U3850 ( .A(DATAO_REG_15__SCAN_IN), .ZN(n4416) );
  NAND2_X1 U3851 ( .A1(n4580), .A2(U4043), .ZN(n2956) );
  OAI21_X1 U3852 ( .B1(U4043), .B2(n4416), .A(n2956), .ZN(U3565) );
  INV_X1 U3853 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n4403) );
  NAND2_X1 U3854 ( .A1(n3636), .A2(U4043), .ZN(n2957) );
  OAI21_X1 U3855 ( .B1(U4043), .B2(n4403), .A(n2957), .ZN(U3563) );
  INV_X1 U3856 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n4389) );
  NAND2_X1 U3857 ( .A1(n4547), .A2(U4043), .ZN(n2958) );
  OAI21_X1 U3858 ( .B1(U4043), .B2(n4389), .A(n2958), .ZN(U3569) );
  NAND2_X2 U3859 ( .A1(n2959), .A2(n2960), .ZN(n3151) );
  NAND2_X1 U3860 ( .A1(n3597), .A2(n3226), .ZN(n2962) );
  NAND2_X1 U3861 ( .A1(n2962), .A2(n2961), .ZN(n3017) );
  NOR2_X1 U3862 ( .A1(n2960), .A2(n2963), .ZN(n2964) );
  INV_X1 U3863 ( .A(n3615), .ZN(n2965) );
  INV_X1 U3864 ( .A(n2960), .ZN(n2966) );
  AOI22_X1 U3865 ( .A1(n3597), .A2(n3189), .B1(n2966), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n2967) );
  XNOR2_X1 U3866 ( .A(n3019), .B(n3018), .ZN(n3192) );
  NOR2_X1 U3867 ( .A1(n4784), .A2(n4783), .ZN(n2970) );
  INV_X1 U3868 ( .A(REG2_REG_0__SCAN_IN), .ZN(n3088) );
  AOI21_X1 U3869 ( .B1(n4784), .B2(n3088), .A(n4783), .ZN(n4785) );
  NAND2_X1 U3870 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3971) );
  OAI22_X1 U3871 ( .A1(n4785), .A2(IR_REG_0__SCAN_IN), .B1(n3948), .B2(n3971), 
        .ZN(n2969) );
  AOI211_X1 U3872 ( .C1(n3192), .C2(n2970), .A(n3962), .B(n2969), .ZN(n2988)
         );
  OAI211_X1 U3873 ( .C1(n2973), .C2(n2972), .A(n4852), .B(n2971), .ZN(n2981)
         );
  NAND3_X1 U3874 ( .A1(n3972), .A2(n2975), .A3(n2974), .ZN(n2976) );
  NAND3_X1 U3875 ( .A1(n2901), .A2(n2977), .A3(n2976), .ZN(n2980) );
  INV_X1 U3876 ( .A(n4858), .ZN(n3998) );
  NAND2_X1 U3877 ( .A1(n3998), .A2(n2373), .ZN(n2979) );
  AOI22_X1 U3878 ( .A1(n4851), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n2978) );
  NAND4_X1 U3879 ( .A1(n2981), .A2(n2980), .A3(n2979), .A4(n2978), .ZN(n2982)
         );
  OR2_X1 U3880 ( .A1(n2988), .A2(n2982), .ZN(U3242) );
  INV_X1 U3881 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n4421) );
  NAND2_X1 U3882 ( .A1(n4500), .A2(U4043), .ZN(n2983) );
  OAI21_X1 U3883 ( .B1(U4043), .B2(n4421), .A(n2983), .ZN(U3571) );
  XNOR2_X1 U3884 ( .A(n2984), .B(REG2_REG_4__SCAN_IN), .ZN(n2993) );
  INV_X1 U3885 ( .A(REG3_REG_4__SCAN_IN), .ZN(n4391) );
  NOR2_X1 U3886 ( .A1(STATE_REG_SCAN_IN), .A2(n4391), .ZN(n3057) );
  AOI21_X1 U3887 ( .B1(n4851), .B2(ADDR_REG_4__SCAN_IN), .A(n3057), .ZN(n2985)
         );
  OAI21_X1 U3888 ( .B1(n4858), .B2(n2986), .A(n2985), .ZN(n2987) );
  NOR2_X1 U3889 ( .A1(n2988), .A2(n2987), .ZN(n2992) );
  OAI211_X1 U3890 ( .C1(n2990), .C2(REG1_REG_4__SCAN_IN), .A(n2989), .B(n4852), 
        .ZN(n2991) );
  OAI211_X1 U3891 ( .C1(n2993), .C2(n4845), .A(n2992), .B(n2991), .ZN(U3244)
         );
  XOR2_X1 U3892 ( .A(n2994), .B(REG2_REG_6__SCAN_IN), .Z(n3001) );
  NAND2_X1 U3893 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3217) );
  NAND2_X1 U3894 ( .A1(n4851), .A2(ADDR_REG_6__SCAN_IN), .ZN(n2995) );
  OAI211_X1 U3895 ( .C1(n4858), .C2(n2996), .A(n3217), .B(n2995), .ZN(n3000)
         );
  AOI211_X1 U3896 ( .C1(n2901), .C2(n3001), .A(n3000), .B(n2999), .ZN(n3002)
         );
  INV_X1 U3897 ( .A(n3002), .ZN(U3246) );
  INV_X1 U3898 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n4295) );
  NAND2_X1 U3899 ( .A1(n4481), .A2(U4043), .ZN(n3003) );
  OAI21_X1 U3900 ( .B1(U4043), .B2(n4295), .A(n3003), .ZN(U3570) );
  MUX2_X1 U3901 ( .A(n3005), .B(REG1_REG_7__SCAN_IN), .S(n3004), .Z(n3006) );
  XNOR2_X1 U3902 ( .A(n3007), .B(n3006), .ZN(n3015) );
  AND2_X1 U3903 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3167) );
  NOR2_X1 U3904 ( .A1(n4858), .A2(n3008), .ZN(n3009) );
  AOI211_X1 U3905 ( .C1(n4851), .C2(ADDR_REG_7__SCAN_IN), .A(n3167), .B(n3009), 
        .ZN(n3014) );
  OAI211_X1 U3906 ( .C1(n3012), .C2(n3011), .A(n3010), .B(n2901), .ZN(n3013)
         );
  OAI211_X1 U3907 ( .C1(n3015), .C2(n4838), .A(n3014), .B(n3013), .ZN(U3247)
         );
  INV_X1 U3908 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n4269) );
  NAND2_X1 U3909 ( .A1(n3664), .A2(U4043), .ZN(n3016) );
  OAI21_X1 U3910 ( .B1(U4043), .B2(n4269), .A(n3016), .ZN(U3572) );
  NAND2_X1 U3911 ( .A1(n3950), .A2(n4012), .ZN(n3054) );
  XNOR2_X1 U3912 ( .A(n3020), .B(n3612), .ZN(n3024) );
  INV_X1 U3913 ( .A(n3023), .ZN(n3022) );
  OAI22_X1 U3914 ( .A1(n3246), .A2(n3151), .B1(n3292), .B2(n3026), .ZN(n3027)
         );
  XNOR2_X1 U3915 ( .A(n3027), .B(n3612), .ZN(n3029) );
  NOR2_X1 U3916 ( .A1(n3029), .A2(n3028), .ZN(n3030) );
  AOI21_X1 U3917 ( .B1(n3029), .B2(n3028), .A(n3030), .ZN(n3754) );
  NAND2_X1 U3918 ( .A1(n3755), .A2(n3754), .ZN(n3753) );
  INV_X1 U3919 ( .A(n3030), .ZN(n3031) );
  NAND2_X1 U3920 ( .A1(n3753), .A2(n3031), .ZN(n3090) );
  OAI22_X1 U3921 ( .A1(n3059), .A2(n3615), .B1(n3245), .B2(n2123), .ZN(n3035)
         );
  XNOR2_X1 U3922 ( .A(n3032), .B(n3612), .ZN(n3034) );
  XOR2_X1 U3923 ( .A(n3035), .B(n3034), .Z(n3091) );
  NAND2_X1 U3924 ( .A1(n3090), .A2(n3091), .ZN(n3089) );
  OAI22_X1 U3925 ( .A1(n3247), .A2(n2123), .B1(n3105), .B2(n3611), .ZN(n3033)
         );
  OAI22_X1 U3926 ( .A1(n3247), .A2(n3615), .B1(n3105), .B2(n2124), .ZN(n3147)
         );
  XNOR2_X1 U3927 ( .A(n3146), .B(n3147), .ZN(n3049) );
  INV_X1 U3928 ( .A(n3034), .ZN(n3037) );
  INV_X1 U3929 ( .A(n3035), .ZN(n3036) );
  NAND2_X1 U3930 ( .A1(n3037), .A2(n3036), .ZN(n3050) );
  INV_X1 U3931 ( .A(n3075), .ZN(n3044) );
  INV_X1 U3932 ( .A(n3039), .ZN(n3043) );
  NAND2_X1 U3933 ( .A1(n3040), .A2(D_REG_1__SCAN_IN), .ZN(n3042) );
  AOI21_X1 U3934 ( .B1(n3043), .B2(n3042), .A(n3041), .ZN(n3076) );
  NAND2_X1 U3935 ( .A1(n3044), .A2(n3076), .ZN(n3061) );
  INV_X1 U3936 ( .A(n3046), .ZN(n3047) );
  NAND2_X1 U3937 ( .A1(n2183), .A2(n3047), .ZN(n3048) );
  NAND2_X1 U3938 ( .A1(n3150), .A2(n2401), .ZN(n3073) );
  AOI21_X1 U3939 ( .B1(n3089), .B2(n3050), .A(n3049), .ZN(n3072) );
  INV_X1 U3940 ( .A(n3051), .ZN(n3060) );
  INV_X1 U3941 ( .A(n3054), .ZN(n3055) );
  NAND2_X1 U3942 ( .A1(n4877), .A2(n3055), .ZN(n3056) );
  INV_X1 U3943 ( .A(n3057), .ZN(n3058) );
  OAI21_X1 U3944 ( .B1(n3780), .B2(n3059), .A(n3058), .ZN(n3070) );
  NAND2_X1 U3945 ( .A1(n3061), .A2(n3060), .ZN(n3188) );
  NOR2_X1 U3946 ( .A1(n3063), .A2(n3062), .ZN(n3064) );
  AND2_X1 U3947 ( .A1(n2960), .A2(n3064), .ZN(n3065) );
  NAND2_X1 U3948 ( .A1(n3188), .A2(n3065), .ZN(n3066) );
  OAI22_X1 U3949 ( .A1(n3778), .A2(n3106), .B1(n3769), .B2(n3218), .ZN(n3069)
         );
  AOI211_X1 U3950 ( .C1(n3100), .C2(n3772), .A(n3070), .B(n3069), .ZN(n3071)
         );
  OAI21_X1 U3951 ( .B1(n3073), .B2(n3072), .A(n3071), .ZN(U3227) );
  INV_X1 U3952 ( .A(n3074), .ZN(n3187) );
  NAND3_X1 U3953 ( .A1(n3076), .A2(n3187), .A3(n3075), .ZN(n3077) );
  INV_X1 U3954 ( .A(n3078), .ZN(n3082) );
  NAND2_X1 U3955 ( .A1(n3189), .A2(n3079), .ZN(n4888) );
  NAND2_X1 U3956 ( .A1(n3080), .A2(n3226), .ZN(n3821) );
  NAND2_X1 U3957 ( .A1(n3819), .A2(n3821), .ZN(n4892) );
  NAND2_X1 U3958 ( .A1(n4502), .A2(n4496), .ZN(n3081) );
  AOI22_X1 U3959 ( .A1(n4892), .A2(n3081), .B1(n4559), .B2(n3758), .ZN(n4889)
         );
  OAI21_X1 U3960 ( .B1(n3082), .B2(n4888), .A(n4889), .ZN(n3083) );
  AOI22_X1 U3961 ( .A1(n3083), .A2(n4585), .B1(REG3_REG_0__SCAN_IN), .B2(n4574), .ZN(n3087) );
  NOR2_X1 U3962 ( .A1(n3084), .A2(n4012), .ZN(n3085) );
  NAND2_X1 U3963 ( .A1(n4585), .A2(n3085), .ZN(n4511) );
  INV_X1 U3964 ( .A(n4511), .ZN(n3499) );
  NAND2_X1 U3965 ( .A1(n3499), .A2(n4892), .ZN(n3086) );
  OAI211_X1 U3966 ( .C1(n4585), .C2(n3088), .A(n3087), .B(n3086), .ZN(U3290)
         );
  OAI21_X1 U3967 ( .B1(n3091), .B2(n3090), .A(n3089), .ZN(n3096) );
  OAI22_X1 U3968 ( .A1(n3778), .A2(REG3_REG_3__SCAN_IN), .B1(n3769), .B2(n3247), .ZN(n3095) );
  AOI21_X1 U3969 ( .B1(n3798), .B2(n3964), .A(n3092), .ZN(n3093) );
  OAI21_X1 U3970 ( .B1(n3796), .B2(n3245), .A(n3093), .ZN(n3094) );
  AOI211_X1 U3971 ( .C1(n3096), .C2(n2401), .A(n3095), .B(n3094), .ZN(n3097)
         );
  INV_X1 U3972 ( .A(n3097), .ZN(U3215) );
  XNOR2_X1 U3973 ( .A(n3098), .B(n3900), .ZN(n3108) );
  XNOR2_X1 U3974 ( .A(n3099), .B(n3900), .ZN(n3103) );
  AOI22_X1 U3975 ( .A1(n3963), .A2(n4601), .B1(n3100), .B2(n4599), .ZN(n3101)
         );
  OAI21_X1 U3976 ( .B1(n3218), .B2(n4604), .A(n3101), .ZN(n3102) );
  AOI21_X1 U3977 ( .B1(n3103), .B2(n4607), .A(n3102), .ZN(n3104) );
  OAI21_X1 U3978 ( .B1(n3108), .B2(n4502), .A(n3104), .ZN(n4913) );
  OAI211_X1 U3979 ( .C1(n3256), .C2(n3105), .A(n3143), .B(n4924), .ZN(n4912)
         );
  OAI22_X1 U3980 ( .A1(n4912), .A2(n4004), .B1(n4592), .B2(n3106), .ZN(n3107)
         );
  OAI21_X1 U3981 ( .B1(n4913), .B2(n3107), .A(n4585), .ZN(n3110) );
  INV_X1 U3982 ( .A(n3108), .ZN(n4916) );
  INV_X2 U3983 ( .A(n4585), .ZN(n4609) );
  AOI22_X1 U3984 ( .A1(n4916), .A2(n3499), .B1(REG2_REG_4__SCAN_IN), .B2(n4609), .ZN(n3109) );
  NAND2_X1 U3985 ( .A1(n3110), .A2(n3109), .ZN(U3286) );
  XOR2_X1 U3986 ( .A(n3111), .B(REG1_REG_8__SCAN_IN), .Z(n3119) );
  XOR2_X1 U3987 ( .A(REG2_REG_8__SCAN_IN), .B(n3112), .Z(n3113) );
  NAND2_X1 U3988 ( .A1(n2901), .A2(n3113), .ZN(n3114) );
  NAND2_X1 U3989 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3329) );
  NAND2_X1 U3990 ( .A1(n3114), .A2(n3329), .ZN(n3117) );
  NOR2_X1 U3991 ( .A1(n4858), .A2(n3115), .ZN(n3116) );
  AOI211_X1 U3992 ( .C1(n4851), .C2(ADDR_REG_8__SCAN_IN), .A(n3117), .B(n3116), 
        .ZN(n3118) );
  OAI21_X1 U3993 ( .B1(n3119), .B2(n4838), .A(n3118), .ZN(U3248) );
  NAND2_X1 U3994 ( .A1(n3962), .A2(DATAO_REG_29__SCAN_IN), .ZN(n3120) );
  OAI21_X1 U3995 ( .B1(n3877), .B2(n3962), .A(n3120), .ZN(U3579) );
  NAND2_X1 U3996 ( .A1(n3836), .A2(n3845), .ZN(n3904) );
  XNOR2_X1 U3997 ( .A(n3121), .B(n3904), .ZN(n3305) );
  XNOR2_X1 U3998 ( .A(n3122), .B(n3904), .ZN(n3125) );
  OAI22_X1 U3999 ( .A1(n3218), .A2(n4545), .B1(n2363), .B2(n4565), .ZN(n3123)
         );
  AOI21_X1 U4000 ( .B1(n4559), .B2(n3960), .A(n3123), .ZN(n3124) );
  OAI21_X1 U4001 ( .B1(n3125), .B2(n4496), .A(n3124), .ZN(n3299) );
  AOI21_X1 U4002 ( .B1(n4928), .B2(n3305), .A(n3299), .ZN(n3131) );
  INV_X1 U4003 ( .A(n3200), .ZN(n3126) );
  AOI21_X1 U4004 ( .B1(n3220), .B2(n3141), .A(n3126), .ZN(n3300) );
  INV_X1 U4005 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3127) );
  NOR2_X1 U4006 ( .A1(n4932), .A2(n3127), .ZN(n3128) );
  AOI21_X1 U4007 ( .B1(n3300), .B2(n4755), .A(n3128), .ZN(n3129) );
  OAI21_X1 U4008 ( .B1(n3131), .B2(n4930), .A(n3129), .ZN(U3479) );
  AOI22_X1 U4009 ( .A1(n3300), .A2(n4667), .B1(n4939), .B2(REG1_REG_6__SCAN_IN), .ZN(n3130) );
  OAI21_X1 U4010 ( .B1(n3131), .B2(n4939), .A(n3130), .ZN(U3524) );
  INV_X1 U4011 ( .A(n4502), .ZN(n3495) );
  NAND2_X1 U4012 ( .A1(n4585), .A2(n3495), .ZN(n3132) );
  INV_X1 U4013 ( .A(n3134), .ZN(n3833) );
  NAND2_X1 U4014 ( .A1(n3833), .A2(n3847), .ZN(n3897) );
  XNOR2_X1 U4015 ( .A(n3133), .B(n3897), .ZN(n4919) );
  XNOR2_X1 U4016 ( .A(n3135), .B(n3897), .ZN(n3139) );
  AOI22_X1 U4017 ( .A1(n3136), .A2(n4601), .B1(n3211), .B2(n4599), .ZN(n3137)
         );
  OAI21_X1 U4018 ( .B1(n3195), .B2(n4604), .A(n3137), .ZN(n3138) );
  AOI21_X1 U4019 ( .B1(n3139), .B2(n4607), .A(n3138), .ZN(n4920) );
  MUX2_X1 U4020 ( .A(n3140), .B(n4920), .S(n4585), .Z(n3145) );
  INV_X1 U4021 ( .A(n3141), .ZN(n3142) );
  AOI21_X1 U4022 ( .B1(n3211), .B2(n3143), .A(n3142), .ZN(n4923) );
  AOI22_X1 U4023 ( .A1(n4923), .A2(n4576), .B1(n3209), .B2(n4574), .ZN(n3144)
         );
  OAI211_X1 U4024 ( .C1(n4588), .C2(n4919), .A(n3145), .B(n3144), .ZN(U3285)
         );
  INV_X1 U4025 ( .A(n3146), .ZN(n3148) );
  NAND2_X1 U4026 ( .A1(n3554), .A2(n3211), .ZN(n3153) );
  XNOR2_X1 U4027 ( .A(n3154), .B(n3612), .ZN(n3156) );
  OAI22_X1 U4028 ( .A1(n3218), .A2(n3615), .B1(n2824), .B2(n2124), .ZN(n3155)
         );
  XOR2_X1 U4029 ( .A(n3156), .B(n3155), .Z(n3208) );
  NAND2_X1 U4030 ( .A1(n3597), .A2(n3961), .ZN(n3158) );
  NAND2_X1 U4031 ( .A1(n3554), .A2(n3220), .ZN(n3157) );
  NAND2_X1 U4032 ( .A1(n3158), .A2(n3157), .ZN(n3159) );
  XNOR2_X1 U4033 ( .A(n3159), .B(n3589), .ZN(n3162) );
  INV_X1 U4034 ( .A(n3162), .ZN(n3161) );
  AOI22_X1 U4035 ( .A1(n3602), .A2(n3961), .B1(n3597), .B2(n3220), .ZN(n3163)
         );
  INV_X1 U4036 ( .A(n3163), .ZN(n3160) );
  NAND2_X1 U4037 ( .A1(n3161), .A2(n3160), .ZN(n3215) );
  OAI22_X1 U4038 ( .A1(n3330), .A2(n3615), .B1(n3194), .B2(n2124), .ZN(n3322)
         );
  OAI22_X1 U4039 ( .A1(n3330), .A2(n2123), .B1(n3194), .B2(n3611), .ZN(n3164)
         );
  XNOR2_X1 U4040 ( .A(n3164), .B(n3612), .ZN(n3323) );
  XOR2_X1 U4041 ( .A(n3322), .B(n3323), .Z(n3165) );
  OAI211_X1 U4042 ( .C1(n3166), .C2(n3165), .A(n3324), .B(n2401), .ZN(n3173)
         );
  INV_X1 U40430 ( .A(n3167), .ZN(n3168) );
  OAI21_X1 U4044 ( .B1(n3780), .B2(n3195), .A(n3168), .ZN(n3171) );
  INV_X1 U4045 ( .A(n3169), .ZN(n3202) );
  OAI22_X1 U4046 ( .A1(n3778), .A2(n3202), .B1(n3769), .B2(n3369), .ZN(n3170)
         );
  AOI211_X1 U4047 ( .C1(n3201), .C2(n3772), .A(n3171), .B(n3170), .ZN(n3172)
         );
  NAND2_X1 U4048 ( .A1(n3173), .A2(n3172), .ZN(U3210) );
  AOI21_X1 U4049 ( .B1(n3189), .B2(n2486), .A(n3293), .ZN(n4898) );
  OR2_X1 U4050 ( .A1(n2753), .A2(n3174), .ZN(n3175) );
  NAND2_X1 U4051 ( .A1(n3176), .A2(n3175), .ZN(n4895) );
  INV_X1 U4052 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3177) );
  OAI22_X1 U4053 ( .A1(n4511), .A2(n4895), .B1(n3177), .B2(n4592), .ZN(n3185)
         );
  NAND2_X1 U4054 ( .A1(n2486), .A2(n4599), .ZN(n3179) );
  NAND2_X1 U4055 ( .A1(n3226), .A2(n4601), .ZN(n3178) );
  OAI211_X1 U4056 ( .C1(n3246), .C2(n4604), .A(n3179), .B(n3178), .ZN(n3180)
         );
  INV_X1 U4057 ( .A(n3180), .ZN(n3183) );
  XNOR2_X1 U4058 ( .A(n2753), .B(n3819), .ZN(n3181) );
  NAND2_X1 U4059 ( .A1(n3181), .A2(n4607), .ZN(n3182) );
  OAI211_X1 U4060 ( .C1(n4895), .C2(n4502), .A(n3183), .B(n3182), .ZN(n4896)
         );
  MUX2_X1 U4061 ( .A(n4896), .B(REG2_REG_1__SCAN_IN), .S(n4609), .Z(n3184) );
  AOI211_X1 U4062 ( .C1(n4576), .C2(n4898), .A(n3185), .B(n3184), .ZN(n3186)
         );
  INV_X1 U4063 ( .A(n3186), .ZN(U3289) );
  NAND2_X1 U4064 ( .A1(n3188), .A2(n3187), .ZN(n3757) );
  AOI22_X1 U4065 ( .A1(n3791), .A2(n3758), .B1(REG3_REG_0__SCAN_IN), .B2(n3757), .ZN(n3191) );
  NAND2_X1 U4066 ( .A1(n3759), .A2(n3189), .ZN(n3190) );
  OAI211_X1 U4067 ( .C1(n3192), .C2(n3801), .A(n3191), .B(n3190), .ZN(U3229)
         );
  XNOR2_X1 U4068 ( .A(n3193), .B(n3899), .ZN(n3198) );
  OAI22_X1 U4069 ( .A1(n3195), .A2(n4545), .B1(n3194), .B2(n4565), .ZN(n3196)
         );
  AOI21_X1 U4070 ( .B1(n4559), .B2(n3263), .A(n3196), .ZN(n3197) );
  OAI21_X1 U4071 ( .B1(n3198), .B2(n4496), .A(n3197), .ZN(n4926) );
  INV_X1 U4072 ( .A(n4926), .ZN(n3206) );
  XOR2_X1 U4073 ( .A(n3199), .B(n3899), .Z(n4929) );
  NAND2_X1 U4074 ( .A1(n4929), .A2(n4613), .ZN(n3205) );
  INV_X1 U4075 ( .A(n4924), .ZN(n4900) );
  AOI211_X1 U4076 ( .C1(n3201), .C2(n3200), .A(n4900), .B(n3313), .ZN(n4927)
         );
  OAI22_X1 U4077 ( .A1(n4585), .A2(n2878), .B1(n3202), .B2(n4592), .ZN(n3203)
         );
  AOI21_X1 U4078 ( .B1(n4927), .B2(n4539), .A(n3203), .ZN(n3204) );
  OAI211_X1 U4079 ( .C1(n3206), .C2(n4609), .A(n3205), .B(n3204), .ZN(U3283)
         );
  XNOR2_X1 U4080 ( .A(n3207), .B(n3208), .ZN(n3214) );
  AOI22_X1 U4081 ( .A1(n3793), .A2(n3209), .B1(n3791), .B2(n3961), .ZN(n3213)
         );
  NAND2_X1 U4082 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3980) );
  OAI21_X1 U4083 ( .B1(n3780), .B2(n3247), .A(n3980), .ZN(n3210) );
  AOI21_X1 U4084 ( .B1(n3211), .B2(n3759), .A(n3210), .ZN(n3212) );
  OAI211_X1 U4085 ( .C1(n3214), .C2(n3801), .A(n3213), .B(n3212), .ZN(U3224)
         );
  NAND2_X1 U4086 ( .A1(n2181), .A2(n3215), .ZN(n3216) );
  XNOR2_X1 U4087 ( .A(n2179), .B(n3216), .ZN(n3223) );
  AOI22_X1 U4088 ( .A1(n3793), .A2(n3301), .B1(n3791), .B2(n3960), .ZN(n3222)
         );
  OAI21_X1 U4089 ( .B1(n3780), .B2(n3218), .A(n3217), .ZN(n3219) );
  AOI21_X1 U4090 ( .B1(n3220), .B2(n3759), .A(n3219), .ZN(n3221) );
  OAI211_X1 U4091 ( .C1(n3223), .C2(n3801), .A(n3222), .B(n3221), .ZN(U3236)
         );
  XNOR2_X1 U4092 ( .A(n3225), .B(n3224), .ZN(n3229) );
  AOI22_X1 U4093 ( .A1(n3798), .A2(n3226), .B1(REG3_REG_1__SCAN_IN), .B2(n3757), .ZN(n3228) );
  AOI22_X1 U4094 ( .A1(n2486), .A2(n3759), .B1(n3791), .B2(n3964), .ZN(n3227)
         );
  OAI211_X1 U4095 ( .C1(n3229), .C2(n3801), .A(n3228), .B(n3227), .ZN(U3219)
         );
  INV_X1 U4096 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n4419) );
  NAND2_X1 U4097 ( .A1(n4098), .A2(U4043), .ZN(n3230) );
  OAI21_X1 U4098 ( .B1(U4043), .B2(n4419), .A(n3230), .ZN(U3577) );
  XNOR2_X1 U4099 ( .A(n3232), .B(n3231), .ZN(n3241) );
  NOR2_X1 U4100 ( .A1(STATE_REG_SCAN_IN), .A2(n3233), .ZN(n3367) );
  AOI21_X1 U4101 ( .B1(n4851), .B2(ADDR_REG_9__SCAN_IN), .A(n3367), .ZN(n3234)
         );
  INV_X1 U4102 ( .A(n3234), .ZN(n3239) );
  AOI211_X1 U4103 ( .C1(n3237), .C2(n3236), .A(n4845), .B(n3235), .ZN(n3238)
         );
  AOI211_X1 U4104 ( .C1(n3998), .C2(n4777), .A(n3239), .B(n3238), .ZN(n3240)
         );
  OAI21_X1 U4105 ( .B1(n3241), .B2(n4838), .A(n3240), .ZN(U3249) );
  INV_X1 U4106 ( .A(n3243), .ZN(n3898) );
  XNOR2_X1 U4107 ( .A(n3242), .B(n3898), .ZN(n4908) );
  NAND2_X1 U4108 ( .A1(n4908), .A2(n3495), .ZN(n3253) );
  XNOR2_X1 U4109 ( .A(n3244), .B(n3243), .ZN(n3251) );
  OAI22_X1 U4110 ( .A1(n3246), .A2(n4545), .B1(n3245), .B2(n4565), .ZN(n3249)
         );
  NOR2_X1 U4111 ( .A1(n3247), .A2(n4604), .ZN(n3248) );
  OR2_X1 U4112 ( .A1(n3249), .A2(n3248), .ZN(n3250) );
  AOI21_X1 U4113 ( .B1(n3251), .B2(n4607), .A(n3250), .ZN(n3252) );
  AND2_X1 U4114 ( .A1(n3253), .A2(n3252), .ZN(n4910) );
  AND2_X1 U4115 ( .A1(n3291), .A2(n3254), .ZN(n3255) );
  NOR2_X1 U4116 ( .A1(n3256), .A2(n3255), .ZN(n4907) );
  INV_X1 U4117 ( .A(n4907), .ZN(n3258) );
  AOI22_X1 U4118 ( .A1(n4609), .A2(REG2_REG_3__SCAN_IN), .B1(n4574), .B2(n4237), .ZN(n3257) );
  OAI21_X1 U4119 ( .B1(n4594), .B2(n3258), .A(n3257), .ZN(n3259) );
  AOI21_X1 U4120 ( .B1(n3499), .B2(n4908), .A(n3259), .ZN(n3260) );
  OAI21_X1 U4121 ( .B1(n4609), .B2(n4910), .A(n3260), .ZN(U3287) );
  INV_X1 U4122 ( .A(n3849), .ZN(n3261) );
  NAND2_X1 U4123 ( .A1(n3261), .A2(n3841), .ZN(n3901) );
  XNOR2_X1 U4124 ( .A(n3262), .B(n3901), .ZN(n3266) );
  AOI22_X1 U4125 ( .A1(n3263), .A2(n4601), .B1(n3373), .B2(n4599), .ZN(n3264)
         );
  OAI21_X1 U4126 ( .B1(n3443), .B2(n4604), .A(n3264), .ZN(n3265) );
  AOI21_X1 U4127 ( .B1(n3266), .B2(n4607), .A(n3265), .ZN(n3278) );
  INV_X1 U4128 ( .A(n3347), .ZN(n3267) );
  AOI21_X1 U4129 ( .B1(n3373), .B2(n3314), .A(n3267), .ZN(n3274) );
  AOI22_X1 U4130 ( .A1(n3274), .A2(n4755), .B1(REG0_REG_9__SCAN_IN), .B2(n4930), .ZN(n3269) );
  XNOR2_X1 U4131 ( .A(n2176), .B(n3901), .ZN(n3275) );
  NAND2_X1 U4132 ( .A1(n4932), .A2(n4928), .ZN(n4758) );
  INV_X1 U4133 ( .A(n4758), .ZN(n4760) );
  NAND2_X1 U4134 ( .A1(n3275), .A2(n4760), .ZN(n3268) );
  OAI211_X1 U4135 ( .C1(n3278), .C2(n4930), .A(n3269), .B(n3268), .ZN(U3485)
         );
  AOI22_X1 U4136 ( .A1(n3274), .A2(n4667), .B1(REG1_REG_9__SCAN_IN), .B2(n4939), .ZN(n3271) );
  NAND2_X1 U4137 ( .A1(n4941), .A2(n4928), .ZN(n4670) );
  INV_X1 U4138 ( .A(n4670), .ZN(n4671) );
  NAND2_X1 U4139 ( .A1(n3275), .A2(n4671), .ZN(n3270) );
  OAI211_X1 U4140 ( .C1(n3278), .C2(n4939), .A(n3271), .B(n3270), .ZN(U3527)
         );
  OAI22_X1 U4141 ( .A1(n4585), .A2(n3272), .B1(n3370), .B2(n4592), .ZN(n3273)
         );
  AOI21_X1 U4142 ( .B1(n3274), .B2(n4576), .A(n3273), .ZN(n3277) );
  NAND2_X1 U4143 ( .A1(n3275), .A2(n4613), .ZN(n3276) );
  OAI211_X1 U4144 ( .C1(n3278), .C2(n4609), .A(n3277), .B(n3276), .ZN(U3281)
         );
  XNOR2_X1 U4145 ( .A(n3279), .B(n2755), .ZN(n3290) );
  CLKBUF_X1 U4146 ( .A(n3281), .Z(n3283) );
  NAND2_X1 U4147 ( .A1(n3283), .A2(n3282), .ZN(n3284) );
  NAND2_X1 U4148 ( .A1(n3280), .A2(n3284), .ZN(n4905) );
  NAND2_X1 U4149 ( .A1(n4905), .A2(n3495), .ZN(n3289) );
  NAND2_X1 U4150 ( .A1(n3760), .A2(n4599), .ZN(n3286) );
  NAND2_X1 U4151 ( .A1(n3963), .A2(n4559), .ZN(n3285) );
  OAI211_X1 U4152 ( .C1(n2478), .C2(n4545), .A(n3286), .B(n3285), .ZN(n3287)
         );
  INV_X1 U4153 ( .A(n3287), .ZN(n3288) );
  OAI211_X1 U4154 ( .C1(n3290), .C2(n4496), .A(n3289), .B(n3288), .ZN(n4903)
         );
  MUX2_X1 U4155 ( .A(n4903), .B(REG2_REG_2__SCAN_IN), .S(n4609), .Z(n3298) );
  INV_X1 U4156 ( .A(n3291), .ZN(n4901) );
  NOR2_X1 U4157 ( .A1(n3293), .A2(n3292), .ZN(n4902) );
  NOR3_X1 U4158 ( .A1(n4594), .A2(n4901), .A3(n4902), .ZN(n3297) );
  INV_X1 U4159 ( .A(n4905), .ZN(n3295) );
  INV_X1 U4160 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3294) );
  OAI22_X1 U4161 ( .A1(n3295), .A2(n4511), .B1(n3294), .B2(n4592), .ZN(n3296)
         );
  OR3_X1 U4162 ( .A1(n3298), .A2(n3297), .A3(n3296), .ZN(U3288) );
  INV_X1 U4163 ( .A(n3299), .ZN(n3307) );
  INV_X1 U4164 ( .A(n3300), .ZN(n3303) );
  AOI22_X1 U4165 ( .A1(n4609), .A2(REG2_REG_6__SCAN_IN), .B1(n3301), .B2(n4574), .ZN(n3302) );
  OAI21_X1 U4166 ( .B1(n3303), .B2(n4594), .A(n3302), .ZN(n3304) );
  AOI21_X1 U4167 ( .B1(n3305), .B2(n4613), .A(n3304), .ZN(n3306) );
  OAI21_X1 U4168 ( .B1(n3307), .B2(n4609), .A(n3306), .ZN(U3284) );
  NAND2_X1 U4169 ( .A1(n3840), .A2(n3838), .ZN(n3890) );
  XOR2_X1 U4170 ( .A(n3308), .B(n3890), .Z(n3311) );
  OAI22_X1 U4171 ( .A1(n3359), .A2(n4604), .B1(n3330), .B2(n4545), .ZN(n3309)
         );
  AOI21_X1 U4172 ( .B1(n3332), .B2(n4599), .A(n3309), .ZN(n3310) );
  OAI21_X1 U4173 ( .B1(n3311), .B2(n4496), .A(n3310), .ZN(n3336) );
  INV_X1 U4174 ( .A(n3336), .ZN(n3321) );
  XOR2_X1 U4175 ( .A(n3890), .B(n3312), .Z(n3337) );
  INV_X1 U4176 ( .A(n3313), .ZN(n3316) );
  INV_X1 U4177 ( .A(n3314), .ZN(n3315) );
  AOI21_X1 U4178 ( .B1(n3332), .B2(n3316), .A(n3315), .ZN(n3339) );
  INV_X1 U4179 ( .A(n3339), .ZN(n3318) );
  AOI22_X1 U4180 ( .A1(n4609), .A2(REG2_REG_8__SCAN_IN), .B1(n3328), .B2(n4574), .ZN(n3317) );
  OAI21_X1 U4181 ( .B1(n3318), .B2(n4594), .A(n3317), .ZN(n3319) );
  AOI21_X1 U4182 ( .B1(n3337), .B2(n4613), .A(n3319), .ZN(n3320) );
  OAI21_X1 U4183 ( .B1(n3321), .B2(n4609), .A(n3320), .ZN(U3282) );
  OAI22_X1 U4184 ( .A1(n3369), .A2(n3615), .B1(n3325), .B2(n2124), .ZN(n3361)
         );
  OAI22_X1 U4185 ( .A1(n3369), .A2(n2124), .B1(n3325), .B2(n3611), .ZN(n3326)
         );
  XNOR2_X1 U4186 ( .A(n3326), .B(n3612), .ZN(n3360) );
  XOR2_X1 U4187 ( .A(n3361), .B(n3360), .Z(n3327) );
  XNOR2_X1 U4188 ( .A(n3362), .B(n3327), .ZN(n3335) );
  AOI22_X1 U4189 ( .A1(n3793), .A2(n3328), .B1(n3791), .B2(n3959), .ZN(n3334)
         );
  OAI21_X1 U4190 ( .B1(n3780), .B2(n3330), .A(n3329), .ZN(n3331) );
  AOI21_X1 U4191 ( .B1(n3332), .B2(n3759), .A(n3331), .ZN(n3333) );
  OAI211_X1 U4192 ( .C1(n3335), .C2(n3801), .A(n3334), .B(n3333), .ZN(U3218)
         );
  AOI21_X1 U4193 ( .B1(n3337), .B2(n4928), .A(n3336), .ZN(n3341) );
  AOI22_X1 U4194 ( .A1(n3339), .A2(n4667), .B1(REG1_REG_8__SCAN_IN), .B2(n4939), .ZN(n3338) );
  OAI21_X1 U4195 ( .B1(n3341), .B2(n4939), .A(n3338), .ZN(U3526) );
  AOI22_X1 U4196 ( .A1(n3339), .A2(n4755), .B1(REG0_REG_8__SCAN_IN), .B2(n4930), .ZN(n3340) );
  OAI21_X1 U4197 ( .B1(n3341), .B2(n4930), .A(n3340), .ZN(U3483) );
  NAND2_X1 U4198 ( .A1(n3844), .A2(n3816), .ZN(n3896) );
  XNOR2_X1 U4199 ( .A(n3342), .B(n3896), .ZN(n3345) );
  OAI22_X1 U4200 ( .A1(n3359), .A2(n4545), .B1(n3457), .B2(n4604), .ZN(n3343)
         );
  AOI21_X1 U4201 ( .B1(n3419), .B2(n4599), .A(n3343), .ZN(n3344) );
  OAI21_X1 U4202 ( .B1(n3345), .B2(n4496), .A(n3344), .ZN(n3386) );
  INV_X1 U4203 ( .A(n3386), .ZN(n3354) );
  XOR2_X1 U4204 ( .A(n3346), .B(n3896), .Z(n3387) );
  NAND2_X1 U4205 ( .A1(n3387), .A2(n4613), .ZN(n3353) );
  AND2_X1 U4206 ( .A1(n3347), .A2(n3419), .ZN(n3348) );
  NOR2_X1 U4207 ( .A1(n3381), .A2(n3348), .ZN(n3389) );
  INV_X1 U4208 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3350) );
  INV_X1 U4209 ( .A(n3349), .ZN(n3427) );
  OAI22_X1 U4210 ( .A1(n4585), .A2(n3350), .B1(n3427), .B2(n4592), .ZN(n3351)
         );
  AOI21_X1 U4211 ( .B1(n3389), .B2(n4576), .A(n3351), .ZN(n3352) );
  OAI211_X1 U4212 ( .C1(n4609), .C2(n3354), .A(n3353), .B(n3352), .ZN(U3280)
         );
  NAND2_X1 U4213 ( .A1(n3597), .A2(n3959), .ZN(n3356) );
  NAND2_X1 U4214 ( .A1(n3554), .A2(n3373), .ZN(n3355) );
  NAND2_X1 U4215 ( .A1(n3356), .A2(n3355), .ZN(n3357) );
  XNOR2_X1 U4216 ( .A(n3357), .B(n3612), .ZN(n3422) );
  OAI22_X1 U4217 ( .A1(n3359), .A2(n3615), .B1(n3358), .B2(n2124), .ZN(n3421)
         );
  XNOR2_X1 U4218 ( .A(n3422), .B(n3421), .ZN(n3366) );
  NAND2_X1 U4219 ( .A1(n3362), .A2(n3361), .ZN(n3363) );
  NAND2_X1 U4220 ( .A1(n3364), .A2(n3363), .ZN(n3365) );
  AOI21_X1 U4221 ( .B1(n3366), .B2(n3365), .A(n3424), .ZN(n3375) );
  INV_X1 U4222 ( .A(n3367), .ZN(n3368) );
  OAI21_X1 U4223 ( .B1(n3780), .B2(n3369), .A(n3368), .ZN(n3372) );
  OAI22_X1 U4224 ( .A1(n3778), .A2(n3370), .B1(n3769), .B2(n3443), .ZN(n3371)
         );
  AOI211_X1 U4225 ( .C1(n3373), .C2(n3772), .A(n3372), .B(n3371), .ZN(n3374)
         );
  OAI21_X1 U4226 ( .B1(n3375), .B2(n3801), .A(n3374), .ZN(U3228) );
  XOR2_X1 U4227 ( .A(n3376), .B(n3902), .Z(n3379) );
  AOI22_X1 U4228 ( .A1(n3448), .A2(n4599), .B1(n4601), .B2(n3415), .ZN(n3377)
         );
  OAI21_X1 U4229 ( .B1(n3738), .B2(n4604), .A(n3377), .ZN(n3378) );
  AOI21_X1 U4230 ( .B1(n3379), .B2(n4607), .A(n3378), .ZN(n4688) );
  XNOR2_X1 U4231 ( .A(n3380), .B(n3902), .ZN(n4686) );
  NOR2_X1 U4232 ( .A1(n3381), .A2(n3437), .ZN(n3382) );
  OR2_X1 U4233 ( .A1(n3410), .A2(n3382), .ZN(n4689) );
  AOI22_X1 U4234 ( .A1(n4609), .A2(REG2_REG_11__SCAN_IN), .B1(n3444), .B2(
        n4574), .ZN(n3383) );
  OAI21_X1 U4235 ( .B1(n4689), .B2(n4594), .A(n3383), .ZN(n3384) );
  AOI21_X1 U4236 ( .B1(n4686), .B2(n4613), .A(n3384), .ZN(n3385) );
  OAI21_X1 U4237 ( .B1(n4688), .B2(n4609), .A(n3385), .ZN(U3279) );
  AOI21_X1 U4238 ( .B1(n3387), .B2(n4928), .A(n3386), .ZN(n3392) );
  AOI22_X1 U4239 ( .A1(n3389), .A2(n4755), .B1(REG0_REG_10__SCAN_IN), .B2(
        n4930), .ZN(n3388) );
  OAI21_X1 U4240 ( .B1(n3392), .B2(n4930), .A(n3388), .ZN(U3487) );
  NAND2_X1 U4241 ( .A1(n4939), .A2(REG1_REG_10__SCAN_IN), .ZN(n3391) );
  NAND2_X1 U4242 ( .A1(n3389), .A2(n4667), .ZN(n3390) );
  OAI211_X1 U4243 ( .C1(n3392), .C2(n4939), .A(n3391), .B(n3390), .ZN(U3528)
         );
  XNOR2_X1 U4244 ( .A(n3394), .B(n3393), .ZN(n3401) );
  OAI211_X1 U4245 ( .C1(n3397), .C2(n3396), .A(n3395), .B(n2901), .ZN(n3399)
         );
  INV_X1 U4246 ( .A(REG3_REG_11__SCAN_IN), .ZN(n4235) );
  NOR2_X1 U4247 ( .A1(STATE_REG_SCAN_IN), .A2(n4235), .ZN(n3441) );
  AOI21_X1 U4248 ( .B1(n4851), .B2(ADDR_REG_11__SCAN_IN), .A(n3441), .ZN(n3398) );
  OAI211_X1 U4249 ( .C1(n4858), .C2(n4776), .A(n3399), .B(n3398), .ZN(n3400)
         );
  AOI21_X1 U4250 ( .B1(n3401), .B2(n4852), .A(n3400), .ZN(n3402) );
  INV_X1 U4251 ( .A(n3402), .ZN(U3251) );
  NAND2_X1 U4252 ( .A1(n3404), .A2(n3403), .ZN(n3479) );
  NAND2_X1 U4253 ( .A1(n3476), .A2(n3477), .ZN(n3881) );
  INV_X1 U4254 ( .A(n3881), .ZN(n3408) );
  XNOR2_X1 U4255 ( .A(n3479), .B(n3408), .ZN(n3407) );
  AOI22_X1 U4256 ( .A1(n3958), .A2(n4601), .B1(n3636), .B2(n4559), .ZN(n3405)
         );
  OAI21_X1 U4257 ( .B1(n3454), .B2(n4565), .A(n3405), .ZN(n3406) );
  AOI21_X1 U4258 ( .B1(n3407), .B2(n4607), .A(n3406), .ZN(n3464) );
  XNOR2_X1 U4259 ( .A(n3409), .B(n3408), .ZN(n3463) );
  OR2_X1 U4260 ( .A1(n3410), .A2(n3454), .ZN(n3411) );
  NAND2_X1 U4261 ( .A1(n3485), .A2(n3411), .ZN(n3471) );
  AOI22_X1 U4262 ( .A1(n4609), .A2(REG2_REG_12__SCAN_IN), .B1(n3456), .B2(
        n4574), .ZN(n3412) );
  OAI21_X1 U4263 ( .B1(n3471), .B2(n4594), .A(n3412), .ZN(n3413) );
  AOI21_X1 U4264 ( .B1(n3463), .B2(n4613), .A(n3413), .ZN(n3414) );
  OAI21_X1 U4265 ( .B1(n4609), .B2(n3464), .A(n3414), .ZN(U3278) );
  NAND2_X1 U4266 ( .A1(n3597), .A2(n3415), .ZN(n3417) );
  NAND2_X1 U4267 ( .A1(n3554), .A2(n3419), .ZN(n3416) );
  NAND2_X1 U4268 ( .A1(n3417), .A2(n3416), .ZN(n3418) );
  XNOR2_X1 U4269 ( .A(n3418), .B(n3612), .ZN(n3434) );
  NAND2_X1 U4270 ( .A1(n3597), .A2(n3419), .ZN(n3420) );
  OAI21_X1 U4271 ( .B1(n3443), .B2(n3615), .A(n3420), .ZN(n3435) );
  XNOR2_X1 U4272 ( .A(n3434), .B(n3435), .ZN(n3426) );
  NOR2_X1 U4273 ( .A1(n3422), .A2(n3421), .ZN(n3423) );
  OR2_X1 U4274 ( .A1(n3424), .A2(n3423), .ZN(n3425) );
  AOI211_X1 U4275 ( .C1(n3426), .C2(n3425), .A(n3801), .B(n3433), .ZN(n3432)
         );
  OAI22_X1 U4276 ( .A1(n3778), .A2(n3427), .B1(n3769), .B2(n3457), .ZN(n3431)
         );
  NOR2_X1 U4277 ( .A1(STATE_REG_SCAN_IN), .A2(n2569), .ZN(n4797) );
  AOI21_X1 U4278 ( .B1(n3798), .B2(n3959), .A(n4797), .ZN(n3428) );
  OAI21_X1 U4279 ( .B1(n3796), .B2(n3429), .A(n3428), .ZN(n3430) );
  OR3_X1 U4280 ( .A1(n3432), .A2(n3431), .A3(n3430), .ZN(U3214) );
  OAI22_X1 U4281 ( .A1(n3457), .A2(n2124), .B1(n3437), .B2(n3611), .ZN(n3436)
         );
  XNOR2_X1 U4282 ( .A(n3436), .B(n3612), .ZN(n3439) );
  OAI22_X1 U4283 ( .A1(n3457), .A2(n3615), .B1(n3437), .B2(n2124), .ZN(n3438)
         );
  NOR2_X1 U4284 ( .A1(n3439), .A2(n3438), .ZN(n3452) );
  NAND2_X1 U4285 ( .A1(n3439), .A2(n3438), .ZN(n3451) );
  NAND2_X1 U4286 ( .A1(n2426), .A2(n3451), .ZN(n3440) );
  XNOR2_X1 U4287 ( .A(n2178), .B(n3440), .ZN(n3450) );
  INV_X1 U4288 ( .A(n3441), .ZN(n3442) );
  OAI21_X1 U4289 ( .B1(n3780), .B2(n3443), .A(n3442), .ZN(n3447) );
  INV_X1 U4290 ( .A(n3444), .ZN(n3445) );
  OAI22_X1 U4291 ( .A1(n3778), .A2(n3445), .B1(n3769), .B2(n3738), .ZN(n3446)
         );
  AOI211_X1 U4292 ( .C1(n3448), .C2(n3759), .A(n3447), .B(n3446), .ZN(n3449)
         );
  OAI21_X1 U4293 ( .B1(n3450), .B2(n3801), .A(n3449), .ZN(U3233) );
  OAI22_X1 U4294 ( .A1(n3454), .A2(n3611), .B1(n3738), .B2(n2124), .ZN(n3453)
         );
  OAI22_X1 U4295 ( .A1(n3454), .A2(n2124), .B1(n3738), .B2(n3615), .ZN(n3504)
         );
  XNOR2_X1 U4296 ( .A(n2135), .B(n3504), .ZN(n3455) );
  XNOR2_X1 U4297 ( .A(n3505), .B(n3455), .ZN(n3462) );
  AOI22_X1 U4298 ( .A1(n3793), .A2(n3456), .B1(n3791), .B2(n3636), .ZN(n3461)
         );
  NAND2_X1 U4299 ( .A1(U3149), .A2(REG3_REG_12__SCAN_IN), .ZN(n4804) );
  OAI21_X1 U4300 ( .B1(n3780), .B2(n3457), .A(n4804), .ZN(n3458) );
  AOI21_X1 U4301 ( .B1(n3459), .B2(n3759), .A(n3458), .ZN(n3460) );
  OAI211_X1 U4302 ( .C1(n3462), .C2(n3801), .A(n3461), .B(n3460), .ZN(U3221)
         );
  NAND2_X1 U4303 ( .A1(n3463), .A2(n4928), .ZN(n3465) );
  AND2_X1 U4304 ( .A1(n3465), .A2(n3464), .ZN(n3468) );
  MUX2_X1 U4305 ( .A(n3466), .B(n3468), .S(n4941), .Z(n3467) );
  OAI21_X1 U4306 ( .B1(n4675), .B2(n3471), .A(n3467), .ZN(U3530) );
  INV_X1 U4307 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3469) );
  MUX2_X1 U4308 ( .A(n3469), .B(n3468), .S(n4932), .Z(n3470) );
  OAI21_X1 U4309 ( .B1(n3471), .B2(n4766), .A(n3470), .ZN(U3491) );
  OAI22_X1 U4310 ( .A1(n3738), .A2(n4545), .B1(n3472), .B2(n4565), .ZN(n3483)
         );
  INV_X1 U4311 ( .A(n3473), .ZN(n3475) );
  OR2_X1 U4312 ( .A1(n3475), .A2(n3474), .ZN(n3892) );
  INV_X1 U4313 ( .A(n3476), .ZN(n3478) );
  OAI21_X1 U4314 ( .B1(n3479), .B2(n3478), .A(n3477), .ZN(n3480) );
  XOR2_X1 U4315 ( .A(n3892), .B(n3480), .Z(n3481) );
  NOR2_X1 U4316 ( .A1(n3481), .A2(n4496), .ZN(n3482) );
  AOI211_X1 U4317 ( .C1(n4559), .C2(n4602), .A(n3483), .B(n3482), .ZN(n4684)
         );
  XNOR2_X1 U4318 ( .A(n3484), .B(n3892), .ZN(n4682) );
  NAND2_X1 U4319 ( .A1(n3485), .A2(n3740), .ZN(n3486) );
  NAND2_X1 U4320 ( .A1(n3496), .A2(n3486), .ZN(n4685) );
  AOI22_X1 U4321 ( .A1(n4609), .A2(REG2_REG_13__SCAN_IN), .B1(n3737), .B2(
        n4574), .ZN(n3487) );
  OAI21_X1 U4322 ( .B1(n4685), .B2(n4594), .A(n3487), .ZN(n3488) );
  AOI21_X1 U4323 ( .B1(n4682), .B2(n4613), .A(n3488), .ZN(n3489) );
  OAI21_X1 U4324 ( .B1(n4684), .B2(n4609), .A(n3489), .ZN(U3277) );
  XNOR2_X1 U4325 ( .A(n3490), .B(n3903), .ZN(n4676) );
  OAI21_X1 U4326 ( .B1(n3903), .B2(n3918), .A(n4596), .ZN(n3491) );
  NAND2_X1 U4327 ( .A1(n3491), .A2(n4607), .ZN(n3493) );
  AOI22_X1 U4328 ( .A1(n3636), .A2(n4601), .B1(n3641), .B2(n4599), .ZN(n3492)
         );
  OAI211_X1 U4329 ( .C1(n3692), .C2(n4604), .A(n3493), .B(n3492), .ZN(n3494)
         );
  AOI21_X1 U4330 ( .B1(n4676), .B2(n3495), .A(n3494), .ZN(n4680) );
  NAND2_X1 U4331 ( .A1(n3496), .A2(n3641), .ZN(n4677) );
  AND3_X1 U4332 ( .A1(n4678), .A2(n4576), .A3(n4677), .ZN(n3498) );
  OAI22_X1 U4333 ( .A1(n4585), .A2(n4826), .B1(n3638), .B2(n4592), .ZN(n3497)
         );
  AOI211_X1 U4334 ( .C1(n4676), .C2(n3499), .A(n3498), .B(n3497), .ZN(n3500)
         );
  OAI21_X1 U4335 ( .B1(n4680), .B2(n4609), .A(n3500), .ZN(U3276) );
  INV_X1 U4336 ( .A(D_REG_0__SCAN_IN), .ZN(n3503) );
  AND2_X1 U4337 ( .A1(n4877), .A2(n3501), .ZN(n3502) );
  AOI22_X1 U4338 ( .A1(n4876), .A2(n3503), .B1(n3502), .B2(n2808), .ZN(U3458)
         );
  INV_X1 U4339 ( .A(n3505), .ZN(n3507) );
  NAND2_X1 U4340 ( .A1(n3636), .A2(n3597), .ZN(n3509) );
  NAND2_X1 U4341 ( .A1(n3554), .A2(n3740), .ZN(n3508) );
  NAND2_X1 U4342 ( .A1(n3509), .A2(n3508), .ZN(n3510) );
  XNOR2_X1 U4343 ( .A(n3510), .B(n3589), .ZN(n3512) );
  AOI22_X1 U4344 ( .A1(n3602), .A2(n3636), .B1(n3597), .B2(n3740), .ZN(n3511)
         );
  NOR2_X1 U4345 ( .A1(n3512), .A2(n3511), .ZN(n3735) );
  NAND2_X1 U4346 ( .A1(n3512), .A2(n3511), .ZN(n3733) );
  NAND2_X1 U4347 ( .A1(n4602), .A2(n3597), .ZN(n3514) );
  NAND2_X1 U4348 ( .A1(n3641), .A2(n3554), .ZN(n3513) );
  NAND2_X1 U4349 ( .A1(n3514), .A2(n3513), .ZN(n3515) );
  XNOR2_X1 U4350 ( .A(n3515), .B(n3589), .ZN(n3681) );
  NAND2_X1 U4351 ( .A1(n3602), .A2(n4602), .ZN(n3517) );
  NAND2_X1 U4352 ( .A1(n3641), .A2(n3597), .ZN(n3516) );
  NAND2_X1 U4353 ( .A1(n4561), .A2(n3597), .ZN(n3519) );
  NAND2_X1 U4354 ( .A1(n4579), .A2(n3554), .ZN(n3518) );
  NAND2_X1 U4355 ( .A1(n3519), .A2(n3518), .ZN(n3520) );
  XNOR2_X1 U4356 ( .A(n3520), .B(n3612), .ZN(n3689) );
  NAND2_X1 U4357 ( .A1(n4561), .A2(n3602), .ZN(n3522) );
  NAND2_X1 U4358 ( .A1(n4579), .A2(n3597), .ZN(n3521) );
  NAND2_X1 U4359 ( .A1(n3522), .A2(n3521), .ZN(n3688) );
  NAND2_X1 U4360 ( .A1(n3689), .A2(n3688), .ZN(n3534) );
  NAND2_X1 U4361 ( .A1(n4580), .A2(n3597), .ZN(n3524) );
  NAND2_X1 U4362 ( .A1(n3554), .A2(n4600), .ZN(n3523) );
  NAND2_X1 U4363 ( .A1(n3524), .A2(n3523), .ZN(n3525) );
  XNOR2_X1 U4364 ( .A(n3525), .B(n3612), .ZN(n3532) );
  NAND2_X1 U4365 ( .A1(n4580), .A2(n3602), .ZN(n3527) );
  NAND2_X1 U4366 ( .A1(n3597), .A2(n4600), .ZN(n3526) );
  NAND2_X1 U4367 ( .A1(n3527), .A2(n3526), .ZN(n3789) );
  NAND2_X1 U4368 ( .A1(n3532), .A2(n3789), .ZN(n3528) );
  NAND2_X1 U4369 ( .A1(n3634), .A2(n3530), .ZN(n3543) );
  INV_X1 U4370 ( .A(n3680), .ZN(n3531) );
  INV_X1 U4371 ( .A(n3681), .ZN(n3684) );
  INV_X1 U4372 ( .A(n3789), .ZN(n3533) );
  INV_X1 U4373 ( .A(n3532), .ZN(n3686) );
  NAND3_X1 U4374 ( .A1(n3534), .A2(n3533), .A3(n3686), .ZN(n3541) );
  OAI22_X1 U4375 ( .A1(n4582), .A2(n2124), .B1(n4564), .B2(n3611), .ZN(n3535)
         );
  XNOR2_X1 U4376 ( .A(n3535), .B(n3589), .ZN(n3700) );
  OR2_X1 U4377 ( .A1(n4582), .A2(n3615), .ZN(n3537) );
  NAND2_X1 U4378 ( .A1(n4555), .A2(n3597), .ZN(n3536) );
  INV_X1 U4379 ( .A(n3689), .ZN(n3539) );
  INV_X1 U4380 ( .A(n3688), .ZN(n3538) );
  AND2_X1 U4381 ( .A1(n3539), .A2(n3538), .ZN(n3698) );
  AOI21_X1 U4382 ( .B1(n3700), .B2(n3701), .A(n3698), .ZN(n3540) );
  INV_X1 U4383 ( .A(n3700), .ZN(n3545) );
  NAND2_X1 U4384 ( .A1(n4560), .A2(n3597), .ZN(n3549) );
  NAND2_X1 U4385 ( .A1(n2666), .A2(n3554), .ZN(n3548) );
  NAND2_X1 U4386 ( .A1(n3549), .A2(n3548), .ZN(n3550) );
  XNOR2_X1 U4387 ( .A(n3550), .B(n3589), .ZN(n3553) );
  NOR2_X1 U4388 ( .A1(n2124), .A2(n4544), .ZN(n3551) );
  AOI21_X1 U4389 ( .B1(n4560), .B2(n3602), .A(n3551), .ZN(n3552) );
  NOR2_X1 U4390 ( .A1(n3553), .A2(n3552), .ZN(n3765) );
  NAND2_X1 U4391 ( .A1(n3553), .A2(n3552), .ZN(n3764) );
  NAND2_X1 U4392 ( .A1(n4547), .A2(n3597), .ZN(n3556) );
  NAND2_X1 U4393 ( .A1(n3554), .A2(n4525), .ZN(n3555) );
  NAND2_X1 U4394 ( .A1(n3556), .A2(n3555), .ZN(n3557) );
  XNOR2_X1 U4395 ( .A(n3557), .B(n3612), .ZN(n3559) );
  OAI22_X1 U4396 ( .A1(n4490), .A2(n3615), .B1(n3880), .B2(n2124), .ZN(n3558)
         );
  XOR2_X1 U4397 ( .A(n3559), .B(n3558), .Z(n3655) );
  OAI22_X1 U4398 ( .A1(n4527), .A2(n2124), .B1(n4504), .B2(n3611), .ZN(n3560)
         );
  XNOR2_X1 U4399 ( .A(n3560), .B(n3612), .ZN(n3561) );
  OAI22_X1 U4400 ( .A1(n4527), .A2(n3615), .B1(n4504), .B2(n2124), .ZN(n3562)
         );
  NAND2_X1 U4401 ( .A1(n3561), .A2(n3562), .ZN(n3723) );
  NAND2_X1 U4402 ( .A1(n3722), .A2(n3723), .ZN(n3721) );
  INV_X1 U4403 ( .A(n3561), .ZN(n3564) );
  INV_X1 U4404 ( .A(n3562), .ZN(n3563) );
  NAND2_X1 U4405 ( .A1(n3564), .A2(n3563), .ZN(n3725) );
  NAND2_X1 U4406 ( .A1(n4500), .A2(n3597), .ZN(n3566) );
  OR2_X1 U4407 ( .A1(n3611), .A2(n3568), .ZN(n3565) );
  NAND2_X1 U4408 ( .A1(n3566), .A2(n3565), .ZN(n3567) );
  XNOR2_X1 U4409 ( .A(n3567), .B(n3612), .ZN(n3661) );
  NAND2_X1 U4410 ( .A1(n4500), .A2(n3602), .ZN(n3570) );
  OR2_X1 U4411 ( .A1(n2124), .A2(n3568), .ZN(n3569) );
  NAND2_X1 U4412 ( .A1(n3570), .A2(n3569), .ZN(n3660) );
  NAND2_X1 U4413 ( .A1(n3661), .A2(n3660), .ZN(n3571) );
  OAI22_X1 U4414 ( .A1(n4483), .A2(n2124), .B1(n4469), .B2(n3611), .ZN(n3573)
         );
  XNOR2_X1 U4415 ( .A(n3573), .B(n3612), .ZN(n3576) );
  OAI22_X1 U4416 ( .A1(n4483), .A2(n3615), .B1(n4469), .B2(n2124), .ZN(n3575)
         );
  XNOR2_X1 U4417 ( .A(n3576), .B(n3575), .ZN(n3746) );
  OAI22_X1 U4418 ( .A1(n4465), .A2(n2124), .B1(n4449), .B2(n3611), .ZN(n3574)
         );
  XNOR2_X1 U4419 ( .A(n3574), .B(n3612), .ZN(n3579) );
  OAI22_X1 U4420 ( .A1(n4465), .A2(n3615), .B1(n4449), .B2(n2124), .ZN(n3578)
         );
  XNOR2_X1 U4421 ( .A(n3579), .B(n3578), .ZN(n3645) );
  NOR2_X1 U4422 ( .A1(n3576), .A2(n3575), .ZN(n3646) );
  NOR2_X1 U4423 ( .A1(n3645), .A2(n3646), .ZN(n3577) );
  NAND2_X1 U4424 ( .A1(n3579), .A2(n3578), .ZN(n3582) );
  NOR2_X1 U4425 ( .A1(n2124), .A2(n4135), .ZN(n3580) );
  AOI21_X1 U4426 ( .B1(n3956), .B2(n3602), .A(n3580), .ZN(n3583) );
  OAI22_X1 U4427 ( .A1(n4448), .A2(n2124), .B1(n4135), .B2(n3611), .ZN(n3581)
         );
  XNOR2_X1 U4428 ( .A(n3581), .B(n3612), .ZN(n3714) );
  NAND2_X1 U4429 ( .A1(n3711), .A2(n3714), .ZN(n3586) );
  INV_X1 U4430 ( .A(n3583), .ZN(n3584) );
  NAND2_X1 U4431 ( .A1(n3585), .A2(n3584), .ZN(n3712) );
  NAND2_X1 U4432 ( .A1(n4137), .A2(n3597), .ZN(n3588) );
  OR2_X1 U4433 ( .A1(n3611), .A2(n4120), .ZN(n3587) );
  NAND2_X1 U4434 ( .A1(n3588), .A2(n3587), .ZN(n3590) );
  XNOR2_X1 U4435 ( .A(n3590), .B(n3589), .ZN(n3593) );
  NOR2_X1 U4436 ( .A1(n2124), .A2(n4120), .ZN(n3591) );
  AOI21_X1 U4437 ( .B1(n4137), .B2(n3602), .A(n3591), .ZN(n3592) );
  NAND2_X1 U4438 ( .A1(n3593), .A2(n3592), .ZN(n3670) );
  NOR2_X1 U4439 ( .A1(n3593), .A2(n3592), .ZN(n3671) );
  OAI22_X1 U4440 ( .A1(n4119), .A2(n2124), .B1(n4099), .B2(n3611), .ZN(n3594)
         );
  XNOR2_X1 U4441 ( .A(n3594), .B(n3612), .ZN(n3596) );
  OAI22_X1 U4442 ( .A1(n4119), .A2(n3615), .B1(n4099), .B2(n2124), .ZN(n3595)
         );
  NAND2_X1 U4443 ( .A1(n3596), .A2(n3595), .ZN(n3775) );
  NAND2_X1 U4444 ( .A1(n4098), .A2(n3597), .ZN(n3599) );
  OR2_X1 U4445 ( .A1(n3611), .A2(n4077), .ZN(n3598) );
  NAND2_X1 U4446 ( .A1(n3599), .A2(n3598), .ZN(n3600) );
  XNOR2_X1 U4447 ( .A(n3600), .B(n3612), .ZN(n3618) );
  NOR2_X1 U4448 ( .A1(n2124), .A2(n4077), .ZN(n3601) );
  AOI21_X1 U4449 ( .B1(n4098), .B2(n3602), .A(n3601), .ZN(n3619) );
  XNOR2_X1 U4450 ( .A(n3618), .B(n3619), .ZN(n3609) );
  OAI22_X1 U4451 ( .A1(n4119), .A2(n3780), .B1(STATE_REG_SCAN_IN), .B2(n3603), 
        .ZN(n3606) );
  INV_X1 U4452 ( .A(n4080), .ZN(n3604) );
  OAI22_X1 U4453 ( .A1(n4074), .A2(n3769), .B1(n3778), .B2(n3604), .ZN(n3605)
         );
  AOI211_X1 U4454 ( .C1(n3607), .C2(n3772), .A(n3606), .B(n3605), .ZN(n3608)
         );
  NAND2_X1 U4455 ( .A1(n3610), .A2(n3609), .ZN(n3633) );
  OAI22_X1 U4456 ( .A1(n4074), .A2(n2124), .B1(n3614), .B2(n3611), .ZN(n3613)
         );
  XNOR2_X1 U4457 ( .A(n3613), .B(n3612), .ZN(n3617) );
  OAI22_X1 U4458 ( .A1(n4074), .A2(n3615), .B1(n3614), .B2(n2124), .ZN(n3616)
         );
  XNOR2_X1 U4459 ( .A(n3617), .B(n3616), .ZN(n3624) );
  NAND2_X1 U4460 ( .A1(n3624), .A2(n2401), .ZN(n3632) );
  INV_X1 U4461 ( .A(n3618), .ZN(n3620) );
  NOR2_X1 U4462 ( .A1(n3620), .A2(n3619), .ZN(n3625) );
  NOR3_X1 U4463 ( .A1(n3624), .A2(n3625), .A3(n3801), .ZN(n3621) );
  NAND2_X1 U4464 ( .A1(n3633), .A2(n3621), .ZN(n3631) );
  AOI22_X1 U4465 ( .A1(n4059), .A2(n3793), .B1(n4030), .B2(n3759), .ZN(n3623)
         );
  NAND2_X1 U4466 ( .A1(U3149), .A2(REG3_REG_28__SCAN_IN), .ZN(n3622) );
  OAI211_X1 U4467 ( .C1(n3877), .C2(n3769), .A(n3623), .B(n3622), .ZN(n3629)
         );
  INV_X1 U4468 ( .A(n3624), .ZN(n3627) );
  INV_X1 U4469 ( .A(n3625), .ZN(n3626) );
  NOR3_X1 U4470 ( .A1(n3627), .A2(n3801), .A3(n3626), .ZN(n3628) );
  AOI211_X1 U4471 ( .C1(n3798), .C2(n4098), .A(n3629), .B(n3628), .ZN(n3630)
         );
  OAI211_X1 U4472 ( .C1(n3633), .C2(n3632), .A(n3631), .B(n3630), .ZN(U3217)
         );
  XNOR2_X1 U4473 ( .A(n3681), .B(n3680), .ZN(n3635) );
  XNOR2_X1 U4474 ( .A(n3682), .B(n3635), .ZN(n3643) );
  INV_X1 U4475 ( .A(n3636), .ZN(n3637) );
  NAND2_X1 U4476 ( .A1(U3149), .A2(REG3_REG_14__SCAN_IN), .ZN(n4823) );
  OAI21_X1 U4477 ( .B1(n3780), .B2(n3637), .A(n4823), .ZN(n3640) );
  OAI22_X1 U4478 ( .A1(n3778), .A2(n3638), .B1(n3769), .B2(n3692), .ZN(n3639)
         );
  AOI211_X1 U4479 ( .C1(n3641), .C2(n3772), .A(n3640), .B(n3639), .ZN(n3642)
         );
  OAI21_X1 U4480 ( .B1(n3643), .B2(n3801), .A(n3642), .ZN(U3212) );
  INV_X1 U4481 ( .A(n3644), .ZN(n3744) );
  OAI21_X1 U4482 ( .B1(n3744), .B2(n3646), .A(n3645), .ZN(n3648) );
  NAND3_X1 U4483 ( .A1(n3648), .A2(n2401), .A3(n3647), .ZN(n3653) );
  AOI22_X1 U4484 ( .A1(n3664), .A2(n3798), .B1(n4442), .B2(n3793), .ZN(n3652)
         );
  OAI22_X1 U4485 ( .A1(n4448), .A2(n3769), .B1(STATE_REG_SCAN_IN), .B2(n3649), 
        .ZN(n3650) );
  AOI21_X1 U4486 ( .B1(n2369), .B2(n3772), .A(n3650), .ZN(n3651) );
  NAND3_X1 U4487 ( .A1(n3653), .A2(n3652), .A3(n3651), .ZN(U3213) );
  XOR2_X1 U4488 ( .A(n3655), .B(n3654), .Z(n3659) );
  AOI22_X1 U4489 ( .A1(n4481), .A2(n3791), .B1(n3793), .B2(n4515), .ZN(n3658)
         );
  NAND2_X1 U4490 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4011) );
  OAI21_X1 U4491 ( .B1(n3780), .B2(n3705), .A(n4011), .ZN(n3656) );
  AOI21_X1 U4492 ( .B1(n4525), .B2(n3759), .A(n3656), .ZN(n3657) );
  OAI211_X1 U4493 ( .C1(n3659), .C2(n3801), .A(n3658), .B(n3657), .ZN(U3216)
         );
  XNOR2_X1 U4494 ( .A(n3661), .B(n3660), .ZN(n3662) );
  XNOR2_X1 U4495 ( .A(n3663), .B(n3662), .ZN(n3669) );
  AOI22_X1 U4496 ( .A1(n3664), .A2(n3791), .B1(n4477), .B2(n3793), .ZN(n3668)
         );
  OAI22_X1 U4497 ( .A1(n4527), .A2(n3780), .B1(STATE_REG_SCAN_IN), .B2(n3665), 
        .ZN(n3666) );
  AOI21_X1 U4498 ( .B1(n4480), .B2(n3759), .A(n3666), .ZN(n3667) );
  OAI211_X1 U4499 ( .C1(n3669), .C2(n3801), .A(n3668), .B(n3667), .ZN(U3220)
         );
  NOR2_X1 U4500 ( .A1(n3671), .A2(n2399), .ZN(n3672) );
  XNOR2_X1 U4501 ( .A(n3673), .B(n3672), .ZN(n3679) );
  INV_X1 U4502 ( .A(n3674), .ZN(n4114) );
  INV_X1 U4503 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3675) );
  OAI22_X1 U4504 ( .A1(n4448), .A2(n3780), .B1(STATE_REG_SCAN_IN), .B2(n3675), 
        .ZN(n3677) );
  OAI22_X1 U4505 ( .A1(n4119), .A2(n3769), .B1(n3796), .B2(n4120), .ZN(n3676)
         );
  AOI211_X1 U4506 ( .C1(n4114), .C2(n3793), .A(n3677), .B(n3676), .ZN(n3678)
         );
  OAI21_X1 U4507 ( .B1(n3679), .B2(n3801), .A(n3678), .ZN(U3222) );
  INV_X1 U4508 ( .A(n3682), .ZN(n3685) );
  AOI21_X1 U4509 ( .B1(n3682), .B2(n3681), .A(n3680), .ZN(n3683) );
  AOI21_X1 U4510 ( .B1(n3685), .B2(n3684), .A(n3683), .ZN(n3687) );
  NOR2_X1 U4511 ( .A1(n3687), .A2(n3686), .ZN(n3788) );
  NAND2_X1 U4512 ( .A1(n3687), .A2(n3686), .ZN(n3786) );
  OAI21_X1 U4513 ( .B1(n3788), .B2(n3789), .A(n3786), .ZN(n3690) );
  XNOR2_X1 U4514 ( .A(n3689), .B(n3688), .ZN(n3697) );
  XNOR2_X1 U4515 ( .A(n3690), .B(n3697), .ZN(n3696) );
  AOI22_X1 U4516 ( .A1(n3793), .A2(n4575), .B1(n3791), .B2(n3691), .ZN(n3695)
         );
  NAND2_X1 U4517 ( .A1(U3149), .A2(REG3_REG_16__SCAN_IN), .ZN(n4842) );
  OAI21_X1 U4518 ( .B1(n3780), .B2(n3692), .A(n4842), .ZN(n3693) );
  AOI21_X1 U4519 ( .B1(n4579), .B2(n3759), .A(n3693), .ZN(n3694) );
  OAI211_X1 U4520 ( .C1(n3696), .C2(n3801), .A(n3695), .B(n3694), .ZN(U3223)
         );
  AOI211_X1 U4521 ( .C1(n3789), .C2(n3786), .A(n3697), .B(n3788), .ZN(n3699)
         );
  NOR2_X1 U4522 ( .A1(n3699), .A2(n3698), .ZN(n3703) );
  XOR2_X1 U4523 ( .A(n3701), .B(n3700), .Z(n3702) );
  XNOR2_X1 U4524 ( .A(n3703), .B(n3702), .ZN(n3710) );
  INV_X1 U4525 ( .A(n4561), .ZN(n4605) );
  INV_X1 U4526 ( .A(REG3_REG_17__SCAN_IN), .ZN(n4259) );
  NOR2_X1 U4527 ( .A1(n4259), .A2(STATE_REG_SCAN_IN), .ZN(n4850) );
  INV_X1 U4528 ( .A(n4850), .ZN(n3704) );
  OAI21_X1 U4529 ( .B1(n3780), .B2(n4605), .A(n3704), .ZN(n3708) );
  OAI22_X1 U4530 ( .A1(n3778), .A2(n3706), .B1(n3769), .B2(n3705), .ZN(n3707)
         );
  AOI211_X1 U4531 ( .C1(n4555), .C2(n3772), .A(n3708), .B(n3707), .ZN(n3709)
         );
  OAI21_X1 U4532 ( .B1(n3710), .B2(n3801), .A(n3709), .ZN(U3225) );
  NAND2_X1 U4533 ( .A1(n3712), .A2(n3711), .ZN(n3713) );
  XOR2_X1 U4534 ( .A(n3714), .B(n3713), .Z(n3720) );
  OAI22_X1 U4535 ( .A1(n4465), .A2(n3780), .B1(n3715), .B2(n3778), .ZN(n3718)
         );
  INV_X1 U4536 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3716) );
  OAI22_X1 U4537 ( .A1(n3781), .A2(n3769), .B1(STATE_REG_SCAN_IN), .B2(n3716), 
        .ZN(n3717) );
  AOI211_X1 U4538 ( .C1(n4128), .C2(n3772), .A(n3718), .B(n3717), .ZN(n3719)
         );
  OAI21_X1 U4539 ( .B1(n3720), .B2(n3801), .A(n3719), .ZN(U3226) );
  INV_X1 U4540 ( .A(n3721), .ZN(n3726) );
  AOI21_X1 U4541 ( .B1(n3725), .B2(n3723), .A(n3722), .ZN(n3724) );
  AOI21_X1 U4542 ( .B1(n3726), .B2(n3725), .A(n3724), .ZN(n3731) );
  OAI22_X1 U4543 ( .A1(n4490), .A2(n3780), .B1(STATE_REG_SCAN_IN), .B2(n3727), 
        .ZN(n3729) );
  INV_X1 U4544 ( .A(n4500), .ZN(n3748) );
  OAI22_X1 U4545 ( .A1(n3748), .A2(n3769), .B1(n3778), .B2(n4506), .ZN(n3728)
         );
  AOI211_X1 U4546 ( .C1(n3879), .C2(n3772), .A(n3729), .B(n3728), .ZN(n3730)
         );
  OAI21_X1 U4547 ( .B1(n3731), .B2(n3801), .A(n3730), .ZN(U3230) );
  INV_X1 U4548 ( .A(n3733), .ZN(n3734) );
  NOR2_X1 U4549 ( .A1(n3735), .A2(n3734), .ZN(n3736) );
  XNOR2_X1 U4550 ( .A(n3732), .B(n3736), .ZN(n3743) );
  AOI22_X1 U4551 ( .A1(n3793), .A2(n3737), .B1(n3791), .B2(n4602), .ZN(n3742)
         );
  NAND2_X1 U4552 ( .A1(U3149), .A2(REG3_REG_13__SCAN_IN), .ZN(n4811) );
  OAI21_X1 U4553 ( .B1(n3780), .B2(n3738), .A(n4811), .ZN(n3739) );
  AOI21_X1 U4554 ( .B1(n3740), .B2(n3759), .A(n3739), .ZN(n3741) );
  OAI211_X1 U4555 ( .C1(n3743), .C2(n3801), .A(n3742), .B(n3741), .ZN(U3231)
         );
  AOI21_X1 U4556 ( .B1(n3746), .B2(n3745), .A(n3744), .ZN(n3752) );
  AOI22_X1 U4557 ( .A1(n3957), .A2(n3791), .B1(n3793), .B2(n4470), .ZN(n3751)
         );
  OAI22_X1 U4558 ( .A1(n3748), .A2(n3780), .B1(STATE_REG_SCAN_IN), .B2(n3747), 
        .ZN(n3749) );
  AOI21_X1 U4559 ( .B1(n4462), .B2(n3759), .A(n3749), .ZN(n3750) );
  OAI211_X1 U4560 ( .C1(n3752), .C2(n3801), .A(n3751), .B(n3750), .ZN(U3232)
         );
  OAI21_X1 U4561 ( .B1(n3755), .B2(n3754), .A(n3753), .ZN(n3756) );
  NAND2_X1 U4562 ( .A1(n3756), .A2(n2401), .ZN(n3763) );
  AOI22_X1 U4563 ( .A1(n3798), .A2(n3758), .B1(REG3_REG_2__SCAN_IN), .B2(n3757), .ZN(n3762) );
  AOI22_X1 U4564 ( .A1(n3760), .A2(n3759), .B1(n3791), .B2(n3963), .ZN(n3761)
         );
  NAND3_X1 U4565 ( .A1(n3763), .A2(n3762), .A3(n3761), .ZN(U3234) );
  NOR2_X1 U4566 ( .A1(n3765), .A2(n2385), .ZN(n3766) );
  XNOR2_X1 U4567 ( .A(n3767), .B(n3766), .ZN(n3774) );
  OAI21_X1 U4568 ( .B1(n3780), .B2(n4582), .A(n3768), .ZN(n3771) );
  OAI22_X1 U4569 ( .A1(n3778), .A2(n4537), .B1(n4490), .B2(n3769), .ZN(n3770)
         );
  AOI211_X1 U4570 ( .C1(n2666), .C2(n3772), .A(n3771), .B(n3770), .ZN(n3773)
         );
  OAI21_X1 U4571 ( .B1(n3774), .B2(n3801), .A(n3773), .ZN(U3235) );
  NAND2_X1 U4572 ( .A1(n2396), .A2(n3775), .ZN(n3776) );
  XNOR2_X1 U4573 ( .A(n3777), .B(n3776), .ZN(n3785) );
  INV_X1 U4574 ( .A(n4105), .ZN(n3779) );
  OAI22_X1 U4575 ( .A1(n3779), .A2(n3778), .B1(n3796), .B2(n4099), .ZN(n3783)
         );
  INV_X1 U4576 ( .A(REG3_REG_26__SCAN_IN), .ZN(n4147) );
  OAI22_X1 U4577 ( .A1(n3781), .A2(n3780), .B1(STATE_REG_SCAN_IN), .B2(n4147), 
        .ZN(n3782) );
  AOI211_X1 U4578 ( .C1(n3791), .C2(n4098), .A(n3783), .B(n3782), .ZN(n3784)
         );
  OAI21_X1 U4579 ( .B1(n3785), .B2(n3801), .A(n3784), .ZN(U3237) );
  INV_X1 U4580 ( .A(n3786), .ZN(n3787) );
  NOR2_X1 U4581 ( .A1(n3788), .A2(n3787), .ZN(n3790) );
  XNOR2_X1 U4582 ( .A(n3790), .B(n3789), .ZN(n3802) );
  INV_X1 U4583 ( .A(n4593), .ZN(n3792) );
  AOI22_X1 U4584 ( .A1(n3793), .A2(n3792), .B1(n3791), .B2(n4561), .ZN(n3800)
         );
  NOR2_X1 U4585 ( .A1(n3794), .A2(STATE_REG_SCAN_IN), .ZN(n3996) );
  NOR2_X1 U4586 ( .A1(n3796), .A2(n3795), .ZN(n3797) );
  AOI211_X1 U4587 ( .C1(n3798), .C2(n4602), .A(n3996), .B(n3797), .ZN(n3799)
         );
  OAI211_X1 U4588 ( .C1(n3802), .C2(n3801), .A(n3800), .B(n3799), .ZN(U3238)
         );
  NAND2_X1 U4589 ( .A1(n2126), .A2(DATAI_29_), .ZN(n4049) );
  INV_X1 U4590 ( .A(n4049), .ZN(n4034) );
  NAND2_X1 U4591 ( .A1(n2125), .A2(DATAI_31_), .ZN(n4020) );
  NAND2_X1 U4592 ( .A1(n4019), .A2(n4020), .ZN(n3874) );
  INV_X1 U4593 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4309) );
  NAND2_X1 U4594 ( .A1(n2941), .A2(REG2_REG_30__SCAN_IN), .ZN(n3805) );
  NAND2_X1 U4595 ( .A1(n3803), .A2(REG0_REG_30__SCAN_IN), .ZN(n3804) );
  OAI211_X1 U4596 ( .C1(n3806), .C2(n4309), .A(n3805), .B(n3804), .ZN(n4047)
         );
  AND2_X1 U4597 ( .A1(n2126), .A2(DATAI_30_), .ZN(n4024) );
  INV_X1 U4598 ( .A(n4024), .ZN(n3872) );
  OR2_X1 U4599 ( .A1(n4047), .A2(n3872), .ZN(n3808) );
  NAND2_X1 U4600 ( .A1(n3874), .A2(n3808), .ZN(n3888) );
  AOI21_X1 U4601 ( .B1(n3877), .B2(n4034), .A(n3888), .ZN(n3811) );
  OR2_X1 U4602 ( .A1(n3877), .A2(n4034), .ZN(n3809) );
  NAND2_X1 U4603 ( .A1(n4039), .A2(n3809), .ZN(n3914) );
  AND3_X1 U4604 ( .A1(n3811), .A2(n4041), .A3(n3810), .ZN(n3930) );
  AOI21_X1 U4605 ( .B1(n3811), .B2(n3914), .A(n3930), .ZN(n3935) );
  INV_X1 U4606 ( .A(n3935), .ZN(n3876) );
  INV_X1 U4607 ( .A(n3914), .ZN(n3870) );
  INV_X1 U4608 ( .A(n3812), .ZN(n3862) );
  NAND2_X1 U4609 ( .A1(n3815), .A2(n3814), .ZN(n3843) );
  NAND3_X1 U4610 ( .A1(n3818), .A2(n3817), .A3(n3816), .ZN(n3855) );
  NOR3_X1 U4611 ( .A1(n3849), .A2(n3843), .A3(n3855), .ZN(n3859) );
  INV_X1 U4612 ( .A(n3899), .ZN(n3837) );
  OAI211_X1 U4613 ( .C1(n2127), .C2(n3822), .A(n3821), .B(n3820), .ZN(n3823)
         );
  NAND3_X1 U4614 ( .A1(n3825), .A2(n3824), .A3(n3823), .ZN(n3826) );
  NAND3_X1 U4615 ( .A1(n3828), .A2(n3827), .A3(n3826), .ZN(n3829) );
  NAND3_X1 U4616 ( .A1(n3831), .A2(n3830), .A3(n3829), .ZN(n3832) );
  NAND4_X1 U4617 ( .A1(n3834), .A2(n3833), .A3(n3845), .A4(n3832), .ZN(n3835)
         );
  AND3_X1 U4618 ( .A1(n3837), .A2(n3836), .A3(n3835), .ZN(n3842) );
  NAND2_X1 U4619 ( .A1(n3839), .A2(n3838), .ZN(n3846) );
  OAI211_X1 U4620 ( .C1(n3842), .C2(n3846), .A(n3841), .B(n3840), .ZN(n3858)
         );
  NAND2_X1 U4621 ( .A1(n3843), .A2(n3852), .ZN(n3916) );
  INV_X1 U4622 ( .A(n3844), .ZN(n3851) );
  INV_X1 U4623 ( .A(n3845), .ZN(n3848) );
  NOR4_X1 U4624 ( .A1(n3849), .A2(n3848), .A3(n3847), .A4(n3846), .ZN(n3850)
         );
  NOR2_X1 U4625 ( .A1(n3851), .A2(n3850), .ZN(n3856) );
  NAND2_X1 U4626 ( .A1(n3852), .A2(n4595), .ZN(n3917) );
  INV_X1 U4627 ( .A(n3917), .ZN(n3854) );
  OAI211_X1 U4628 ( .C1(n3856), .C2(n3855), .A(n3854), .B(n3853), .ZN(n3857)
         );
  AOI22_X1 U4629 ( .A1(n3859), .A2(n3858), .B1(n3916), .B2(n3857), .ZN(n3860)
         );
  OAI21_X1 U4630 ( .B1(n2355), .B2(n3860), .A(n3920), .ZN(n3861) );
  AOI21_X1 U4631 ( .B1(n3862), .B2(n3861), .A(n2172), .ZN(n3863) );
  OAI21_X1 U4632 ( .B1(n4444), .B2(n3863), .A(n3925), .ZN(n3864) );
  INV_X1 U4633 ( .A(n3864), .ZN(n3866) );
  OAI211_X1 U4634 ( .C1(n3867), .C2(n3866), .A(n3931), .B(n3865), .ZN(n3868)
         );
  NAND4_X1 U4635 ( .A1(n3871), .A2(n3870), .A3(n3869), .A4(n3868), .ZN(n3875)
         );
  NAND2_X1 U4636 ( .A1(n4047), .A2(n3872), .ZN(n3937) );
  OR2_X1 U4637 ( .A1(n4019), .A2(n4020), .ZN(n3873) );
  NAND2_X1 U4638 ( .A1(n3937), .A2(n3873), .ZN(n3891) );
  AOI22_X1 U4639 ( .A1(n3876), .A2(n3875), .B1(n3874), .B2(n3891), .ZN(n3946)
         );
  XNOR2_X1 U4640 ( .A(n3877), .B(n4049), .ZN(n4043) );
  NAND2_X1 U4641 ( .A1(n3878), .A2(n4115), .ZN(n4133) );
  XNOR2_X1 U4642 ( .A(n4527), .B(n3879), .ZN(n4493) );
  XNOR2_X1 U4643 ( .A(n4547), .B(n3880), .ZN(n4523) );
  NOR4_X1 U4644 ( .A1(n4133), .A2(n4493), .A3(n4523), .A4(n3881), .ZN(n3913)
         );
  INV_X1 U4645 ( .A(n4444), .ZN(n3882) );
  NAND2_X1 U4646 ( .A1(n3882), .A2(n4443), .ZN(n4478) );
  INV_X1 U4647 ( .A(n4478), .ZN(n3912) );
  NAND2_X1 U4648 ( .A1(n4131), .A2(n3883), .ZN(n4447) );
  INV_X1 U4649 ( .A(n4516), .ZN(n3884) );
  INV_X1 U4650 ( .A(n3915), .ZN(n3886) );
  AND2_X1 U4651 ( .A1(n4093), .A2(n3887), .ZN(n4118) );
  NOR3_X1 U4652 ( .A1(n3890), .A2(n3889), .A3(n3888), .ZN(n3894) );
  NOR2_X1 U4653 ( .A1(n3892), .A2(n3891), .ZN(n3893) );
  NAND4_X1 U4654 ( .A1(n4557), .A2(n3895), .A3(n3894), .A4(n3893), .ZN(n3910)
         );
  NOR2_X1 U4655 ( .A1(n4540), .A2(n3896), .ZN(n3908) );
  NOR4_X1 U4656 ( .A1(n2755), .A2(n3898), .A3(n2753), .A4(n3897), .ZN(n3907)
         );
  NOR4_X1 U4657 ( .A1(n3902), .A2(n3901), .A3(n3900), .A4(n3899), .ZN(n3906)
         );
  NOR4_X1 U4658 ( .A1(n2286), .A2(n4597), .A3(n3904), .A4(n4892), .ZN(n3905)
         );
  NAND4_X1 U4659 ( .A1(n3908), .A2(n3907), .A3(n3906), .A4(n3905), .ZN(n3909)
         );
  NOR4_X1 U4660 ( .A1(n4447), .A2(n4456), .A3(n3910), .A4(n3909), .ZN(n3911)
         );
  AND4_X1 U4661 ( .A1(n4043), .A2(n3913), .A3(n3912), .A4(n3911), .ZN(n3943)
         );
  NOR3_X1 U4662 ( .A1(n4068), .A2(n3915), .A3(n3914), .ZN(n3934) );
  OAI21_X1 U4663 ( .B1(n3918), .B2(n3917), .A(n3916), .ZN(n3921) );
  INV_X1 U4664 ( .A(n4492), .ZN(n3919) );
  AOI211_X1 U4665 ( .C1(n3921), .C2(n3920), .A(n2355), .B(n3919), .ZN(n3924)
         );
  OAI21_X1 U4666 ( .B1(n3924), .B2(n3923), .A(n3922), .ZN(n3926) );
  NAND2_X1 U4667 ( .A1(n3926), .A2(n3925), .ZN(n3929) );
  AOI21_X1 U4668 ( .B1(n3929), .B2(n3928), .A(n3927), .ZN(n3932) );
  OAI211_X1 U4669 ( .C1(n3932), .C2(n4091), .A(n3931), .B(n3930), .ZN(n3933)
         );
  OAI21_X1 U4670 ( .B1(n3935), .B2(n3934), .A(n3933), .ZN(n3940) );
  INV_X1 U4671 ( .A(n4019), .ZN(n3936) );
  NAND2_X1 U4672 ( .A1(n3936), .A2(n4024), .ZN(n3939) );
  AOI21_X1 U4673 ( .B1(n3937), .B2(n4019), .A(n4020), .ZN(n3938) );
  AOI21_X1 U4674 ( .B1(n3940), .B2(n3939), .A(n3938), .ZN(n3942) );
  MUX2_X1 U4675 ( .A(n3943), .B(n3942), .S(n2127), .Z(n3945) );
  XNOR2_X1 U4676 ( .A(n3947), .B(n4004), .ZN(n3954) );
  NOR2_X1 U4677 ( .A1(n3949), .A2(n3948), .ZN(n3952) );
  OAI21_X1 U4678 ( .B1(n3953), .B2(n3950), .A(B_REG_SCAN_IN), .ZN(n3951) );
  OAI22_X1 U4679 ( .A1(n3954), .A2(n3953), .B1(n3952), .B2(n3951), .ZN(U3239)
         );
  MUX2_X1 U4680 ( .A(n4047), .B(DATAO_REG_30__SCAN_IN), .S(n3962), .Z(U3580)
         );
  MUX2_X1 U4681 ( .A(n4051), .B(DATAO_REG_28__SCAN_IN), .S(n3962), .Z(U3578)
         );
  MUX2_X1 U4682 ( .A(n3955), .B(DATAO_REG_26__SCAN_IN), .S(n3962), .Z(U3576)
         );
  MUX2_X1 U4683 ( .A(n4137), .B(DATAO_REG_25__SCAN_IN), .S(n3962), .Z(U3575)
         );
  MUX2_X1 U4684 ( .A(n3956), .B(DATAO_REG_24__SCAN_IN), .S(n3962), .Z(U3574)
         );
  MUX2_X1 U4685 ( .A(DATAO_REG_23__SCAN_IN), .B(n3957), .S(U4043), .Z(U3573)
         );
  MUX2_X1 U4686 ( .A(n4602), .B(DATAO_REG_14__SCAN_IN), .S(n3962), .Z(U3564)
         );
  MUX2_X1 U4687 ( .A(DATAO_REG_11__SCAN_IN), .B(n3958), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4688 ( .A(n3959), .B(DATAO_REG_9__SCAN_IN), .S(n3962), .Z(U3559) );
  MUX2_X1 U4689 ( .A(DATAO_REG_7__SCAN_IN), .B(n3960), .S(U4043), .Z(U3557) );
  MUX2_X1 U4690 ( .A(n3961), .B(DATAO_REG_6__SCAN_IN), .S(n3962), .Z(U3556) );
  MUX2_X1 U4691 ( .A(n3963), .B(DATAO_REG_3__SCAN_IN), .S(n3962), .Z(U3553) );
  MUX2_X1 U4692 ( .A(DATAO_REG_2__SCAN_IN), .B(n3964), .S(U4043), .Z(U3552) );
  NOR2_X1 U4693 ( .A1(STATE_REG_SCAN_IN), .A2(n3177), .ZN(n3967) );
  NOR2_X1 U4694 ( .A1(n4858), .A2(n3965), .ZN(n3966) );
  AOI211_X1 U4695 ( .C1(n4851), .C2(ADDR_REG_1__SCAN_IN), .A(n3967), .B(n3966), 
        .ZN(n3976) );
  OAI211_X1 U4696 ( .C1(n3970), .C2(n3969), .A(n4852), .B(n3968), .ZN(n3975)
         );
  OAI211_X1 U4697 ( .C1(n2861), .C2(n3973), .A(n2901), .B(n3972), .ZN(n3974)
         );
  NAND3_X1 U4698 ( .A1(n3976), .A2(n3975), .A3(n3974), .ZN(U3241) );
  OAI211_X1 U4699 ( .C1(n3979), .C2(n3978), .A(n3977), .B(n4852), .ZN(n3988)
         );
  INV_X1 U4700 ( .A(n4851), .ZN(n4844) );
  INV_X1 U4701 ( .A(ADDR_REG_5__SCAN_IN), .ZN(n3981) );
  OAI21_X1 U4702 ( .B1(n4844), .B2(n3981), .A(n3980), .ZN(n3982) );
  AOI21_X1 U4703 ( .B1(n4779), .B2(n3998), .A(n3982), .ZN(n3987) );
  OAI211_X1 U4704 ( .C1(n3985), .C2(n3984), .A(n2901), .B(n3983), .ZN(n3986)
         );
  NAND3_X1 U4705 ( .A1(n3988), .A2(n3987), .A3(n3986), .ZN(U3245) );
  XOR2_X1 U4706 ( .A(n3990), .B(n3989), .Z(n4001) );
  INV_X1 U4707 ( .A(n3991), .ZN(n3992) );
  AOI211_X1 U4708 ( .C1(n3994), .C2(n3993), .A(n3992), .B(n4845), .ZN(n3995)
         );
  AOI211_X1 U4709 ( .C1(n4851), .C2(ADDR_REG_15__SCAN_IN), .A(n3996), .B(n3995), .ZN(n4000) );
  NAND2_X1 U4710 ( .A1(n3998), .A2(n3997), .ZN(n3999) );
  OAI211_X1 U4711 ( .C1(n4001), .C2(n4838), .A(n4000), .B(n3999), .ZN(U3255)
         );
  XNOR2_X1 U4712 ( .A(n4004), .B(REG1_REG_19__SCAN_IN), .ZN(n4005) );
  XNOR2_X1 U4713 ( .A(n4006), .B(n4005), .ZN(n4016) );
  AOI21_X1 U4714 ( .B1(n4775), .B2(REG2_REG_18__SCAN_IN), .A(n4007), .ZN(n4009) );
  MUX2_X1 U4715 ( .A(n4530), .B(REG2_REG_19__SCAN_IN), .S(n4012), .Z(n4008) );
  XNOR2_X1 U4716 ( .A(n4009), .B(n4008), .ZN(n4014) );
  NAND2_X1 U4717 ( .A1(n4851), .A2(ADDR_REG_19__SCAN_IN), .ZN(n4010) );
  OAI211_X1 U4718 ( .C1(n4858), .C2(n4012), .A(n4011), .B(n4010), .ZN(n4013)
         );
  OAI21_X1 U4719 ( .B1(n4016), .B2(n4838), .A(n4015), .ZN(U3259) );
  AND2_X1 U4720 ( .A1(n4784), .A2(B_REG_SCAN_IN), .ZN(n4018) );
  NOR2_X1 U4721 ( .A1(n4604), .A2(n4018), .ZN(n4046) );
  NAND2_X1 U4722 ( .A1(n4019), .A2(n4046), .ZN(n4026) );
  OAI21_X1 U4723 ( .B1(n4020), .B2(n4565), .A(n4026), .ZN(n4690) );
  NAND2_X1 U4724 ( .A1(n4585), .A2(n4690), .ZN(n4022) );
  NAND2_X1 U4725 ( .A1(n4609), .A2(REG2_REG_31__SCAN_IN), .ZN(n4021) );
  OAI211_X1 U4726 ( .C1(n4693), .C2(n4594), .A(n4022), .B(n4021), .ZN(U3260)
         );
  AOI21_X1 U4727 ( .B1(n4024), .B2(n4037), .A(n4023), .ZN(n4618) );
  INV_X1 U4728 ( .A(n4618), .ZN(n4697) );
  INV_X1 U4729 ( .A(REG2_REG_30__SCAN_IN), .ZN(n4027) );
  NAND2_X1 U4730 ( .A1(n4024), .A2(n4599), .ZN(n4025) );
  AND2_X1 U4731 ( .A1(n4026), .A2(n4025), .ZN(n4694) );
  MUX2_X1 U4732 ( .A(n4027), .B(n4694), .S(n4585), .Z(n4028) );
  OAI21_X1 U4733 ( .B1(n4697), .B2(n4594), .A(n4028), .ZN(U3261) );
  INV_X1 U4734 ( .A(n4029), .ZN(n4031) );
  AOI22_X1 U4735 ( .A1(n4032), .A2(n4031), .B1(n4051), .B2(n4030), .ZN(n4033)
         );
  XNOR2_X1 U4736 ( .A(n4033), .B(n4043), .ZN(n4699) );
  NAND2_X1 U4737 ( .A1(n4035), .A2(n4034), .ZN(n4036) );
  NAND2_X1 U4738 ( .A1(n4037), .A2(n4036), .ZN(n4621) );
  INV_X1 U4739 ( .A(n4621), .ZN(n4038) );
  AOI22_X1 U4740 ( .A1(n4038), .A2(n4576), .B1(REG2_REG_29__SCAN_IN), .B2(
        n4609), .ZN(n4057) );
  NAND2_X1 U4741 ( .A1(n4042), .A2(n4041), .ZN(n4044) );
  XNOR2_X1 U4742 ( .A(n4044), .B(n4043), .ZN(n4045) );
  NAND2_X1 U4743 ( .A1(n4045), .A2(n4607), .ZN(n4053) );
  NAND2_X1 U4744 ( .A1(n4047), .A2(n4046), .ZN(n4048) );
  OAI21_X1 U4745 ( .B1(n4049), .B2(n4565), .A(n4048), .ZN(n4050) );
  AOI21_X1 U4746 ( .B1(n4051), .B2(n4601), .A(n4050), .ZN(n4052) );
  NAND2_X1 U4747 ( .A1(n4053), .A2(n4052), .ZN(n4622) );
  NOR2_X1 U4748 ( .A1(n4054), .A2(n4592), .ZN(n4055) );
  OAI21_X1 U4749 ( .B1(n4622), .B2(n4055), .A(n4585), .ZN(n4056) );
  INV_X1 U4750 ( .A(n4058), .ZN(n4065) );
  AOI22_X1 U4751 ( .A1(n4059), .A2(n4574), .B1(REG2_REG_28__SCAN_IN), .B2(
        n4609), .ZN(n4060) );
  OAI21_X1 U4752 ( .B1(n4061), .B2(n4594), .A(n4060), .ZN(n4062) );
  AOI21_X1 U4753 ( .B1(n4063), .B2(n4585), .A(n4062), .ZN(n4064) );
  OAI21_X1 U4754 ( .B1(n4065), .B2(n4588), .A(n4064), .ZN(U3262) );
  XNOR2_X1 U4755 ( .A(n4067), .B(n4066), .ZN(n4703) );
  INV_X1 U4756 ( .A(n4703), .ZN(n4084) );
  NAND2_X1 U4757 ( .A1(n4069), .A2(n4068), .ZN(n4070) );
  NAND2_X1 U4758 ( .A1(n4071), .A2(n4070), .ZN(n4076) );
  OAI22_X1 U4759 ( .A1(n4119), .A2(n4545), .B1(n4077), .B2(n4565), .ZN(n4072)
         );
  INV_X1 U4760 ( .A(n4072), .ZN(n4073) );
  OAI21_X1 U4761 ( .B1(n4074), .B2(n4604), .A(n4073), .ZN(n4075) );
  NOR2_X1 U4762 ( .A1(n4624), .A2(n4609), .ZN(n4083) );
  OR2_X1 U4763 ( .A1(n4087), .A2(n4077), .ZN(n4078) );
  NAND2_X1 U4764 ( .A1(n4079), .A2(n4078), .ZN(n4625) );
  AOI22_X1 U4765 ( .A1(n4080), .A2(n4574), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4609), .ZN(n4081) );
  OAI21_X1 U4766 ( .B1(n4625), .B2(n4594), .A(n4081), .ZN(n4082) );
  AOI211_X1 U4767 ( .C1(n4084), .C2(n4613), .A(n4083), .B(n4082), .ZN(n4085)
         );
  INV_X1 U4768 ( .A(n4085), .ZN(U3263) );
  XNOR2_X1 U4769 ( .A(n4086), .B(n4095), .ZN(n4629) );
  INV_X1 U4770 ( .A(n4087), .ZN(n4090) );
  NAND2_X1 U4771 ( .A1(n4111), .A2(n4088), .ZN(n4089) );
  NAND2_X1 U4772 ( .A1(n4090), .A2(n4089), .ZN(n4707) );
  INV_X1 U4773 ( .A(n4091), .ZN(n4092) );
  NAND2_X1 U4774 ( .A1(n4116), .A2(n4092), .ZN(n4094) );
  NAND2_X1 U4775 ( .A1(n4094), .A2(n4093), .ZN(n4096) );
  XNOR2_X1 U4776 ( .A(n4096), .B(n4095), .ZN(n4097) );
  NAND2_X1 U4777 ( .A1(n4097), .A2(n4607), .ZN(n4104) );
  NAND2_X1 U4778 ( .A1(n4098), .A2(n4559), .ZN(n4102) );
  NOR2_X1 U4779 ( .A1(n4099), .A2(n4565), .ZN(n4100) );
  AOI21_X1 U4780 ( .B1(n4137), .B2(n4601), .A(n4100), .ZN(n4101) );
  AND2_X1 U4781 ( .A1(n4102), .A2(n4101), .ZN(n4103) );
  NAND2_X1 U4782 ( .A1(n4104), .A2(n4103), .ZN(n4628) );
  NAND2_X1 U4783 ( .A1(n4628), .A2(n4585), .ZN(n4107) );
  AOI22_X1 U4784 ( .A1(n4105), .A2(n4574), .B1(REG2_REG_26__SCAN_IN), .B2(
        n4609), .ZN(n4106) );
  OAI211_X1 U4785 ( .C1(n4707), .C2(n4594), .A(n4107), .B(n4106), .ZN(n4108)
         );
  AOI21_X1 U4786 ( .B1(n4629), .B2(n4613), .A(n4108), .ZN(n4109) );
  INV_X1 U4787 ( .A(n4109), .ZN(U3264) );
  XNOR2_X1 U4788 ( .A(n4110), .B(n4118), .ZN(n4712) );
  INV_X1 U4789 ( .A(n4111), .ZN(n4112) );
  AOI21_X1 U4790 ( .B1(n4113), .B2(n4130), .A(n4112), .ZN(n4710) );
  AOI22_X1 U4791 ( .A1(n4710), .A2(n4576), .B1(n4114), .B2(n4574), .ZN(n4126)
         );
  INV_X1 U4792 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4124) );
  NAND2_X1 U4793 ( .A1(n4116), .A2(n4115), .ZN(n4117) );
  XOR2_X1 U4794 ( .A(n4118), .B(n4117), .Z(n4123) );
  NOR2_X1 U4795 ( .A1(n4119), .A2(n4604), .ZN(n4122) );
  OAI22_X1 U4796 ( .A1(n4448), .A2(n4545), .B1(n4120), .B2(n4565), .ZN(n4121)
         );
  MUX2_X1 U4797 ( .A(n4124), .B(n4632), .S(n4585), .Z(n4125) );
  OAI211_X1 U4798 ( .C1(n4712), .C2(n4588), .A(n4126), .B(n4125), .ZN(U3265)
         );
  XOR2_X1 U4799 ( .A(n4133), .B(n4127), .Z(n4636) );
  NAND2_X1 U4800 ( .A1(n4439), .A2(n4128), .ZN(n4129) );
  NAND2_X1 U4801 ( .A1(n4130), .A2(n4129), .ZN(n4716) );
  NAND2_X1 U4802 ( .A1(n4132), .A2(n4131), .ZN(n4134) );
  XNOR2_X1 U4803 ( .A(n4134), .B(n4133), .ZN(n4139) );
  OAI22_X1 U4804 ( .A1(n4465), .A2(n4545), .B1(n4135), .B2(n4565), .ZN(n4136)
         );
  AOI21_X1 U4805 ( .B1(n4137), .B2(n4559), .A(n4136), .ZN(n4138) );
  OAI21_X1 U4806 ( .B1(n4139), .B2(n4496), .A(n4138), .ZN(n4635) );
  NAND2_X1 U4807 ( .A1(n4635), .A2(n4585), .ZN(n4142) );
  AOI22_X1 U4808 ( .A1(n4140), .A2(n4574), .B1(REG2_REG_24__SCAN_IN), .B2(
        n4609), .ZN(n4141) );
  OAI211_X1 U4809 ( .C1(n4716), .C2(n4594), .A(n4142), .B(n4141), .ZN(n4143)
         );
  AOI21_X1 U4810 ( .B1(n4636), .B2(n4613), .A(n4143), .ZN(n4435) );
  NAND2_X1 U4811 ( .A1(REG3_REG_19__SCAN_IN), .A2(n4378), .ZN(n4145) );
  NAND4_X1 U4812 ( .A1(IR_REG_12__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        DATAI_11_), .A4(DATAI_23_), .ZN(n4144) );
  NOR4_X1 U4813 ( .A1(REG1_REG_14__SCAN_IN), .A2(DATAO_REG_10__SCAN_IN), .A3(
        n4145), .A4(n4144), .ZN(n4159) );
  INV_X1 U4814 ( .A(REG0_REG_8__SCAN_IN), .ZN(n4394) );
  NOR4_X1 U4815 ( .A1(DATAI_9_), .A2(REG1_REG_8__SCAN_IN), .A3(
        DATAO_REG_4__SCAN_IN), .A4(n4394), .ZN(n4158) );
  INV_X1 U4816 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4733) );
  NAND4_X1 U4817 ( .A1(REG3_REG_17__SCAN_IN), .A2(DATAI_30_), .A3(
        DATAO_REG_12__SCAN_IN), .A4(n4733), .ZN(n4146) );
  NOR3_X1 U4818 ( .A1(IR_REG_2__SCAN_IN), .A2(DATAO_REG_5__SCAN_IN), .A3(n4146), .ZN(n4157) );
  NOR4_X1 U4819 ( .A1(IR_REG_4__SCAN_IN), .A2(REG0_REG_24__SCAN_IN), .A3(
        REG0_REG_30__SCAN_IN), .A4(DATAO_REG_15__SCAN_IN), .ZN(n4155) );
  NOR4_X1 U4820 ( .A1(REG0_REG_29__SCAN_IN), .A2(REG0_REG_28__SCAN_IN), .A3(
        REG1_REG_28__SCAN_IN), .A4(REG1_REG_30__SCAN_IN), .ZN(n4154) );
  INV_X1 U4821 ( .A(IR_REG_14__SCAN_IN), .ZN(n4280) );
  NAND4_X1 U4822 ( .A1(IR_REG_22__SCAN_IN), .A2(REG2_REG_24__SCAN_IN), .A3(
        DATAI_22_), .A4(n4280), .ZN(n4152) );
  NAND4_X1 U4823 ( .A1(REG0_REG_11__SCAN_IN), .A2(DATAO_REG_21__SCAN_IN), .A3(
        DATAO_REG_27__SCAN_IN), .A4(n4666), .ZN(n4151) );
  NAND4_X1 U4824 ( .A1(D_REG_6__SCAN_IN), .A2(D_REG_10__SCAN_IN), .A3(
        D_REG_30__SCAN_IN), .A4(n4337), .ZN(n4150) );
  INV_X1 U4825 ( .A(IR_REG_10__SCAN_IN), .ZN(n4148) );
  NAND4_X1 U4826 ( .A1(n4148), .A2(n4147), .A3(IR_REG_16__SCAN_IN), .A4(
        REG0_REG_2__SCAN_IN), .ZN(n4149) );
  NOR4_X1 U4827 ( .A1(n4152), .A2(n4151), .A3(n4150), .A4(n4149), .ZN(n4153)
         );
  AND3_X1 U4828 ( .A1(n4155), .A2(n4154), .A3(n4153), .ZN(n4156) );
  AND4_X1 U4829 ( .A1(n4159), .A2(n4158), .A3(n4157), .A4(n4156), .ZN(n4193)
         );
  NOR4_X1 U4830 ( .A1(DATAI_12_), .A2(REG0_REG_18__SCAN_IN), .A3(
        DATAO_REG_19__SCAN_IN), .A4(n2741), .ZN(n4192) );
  NAND4_X1 U4831 ( .A1(D_REG_5__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(
        REG0_REG_21__SCAN_IN), .A4(DATAO_REG_18__SCAN_IN), .ZN(n4169) );
  NAND4_X1 U4832 ( .A1(n4161), .A2(n4160), .A3(IR_REG_13__SCAN_IN), .A4(
        IR_REG_23__SCAN_IN), .ZN(n4168) );
  NAND4_X1 U4833 ( .A1(REG1_REG_13__SCAN_IN), .A2(REG1_REG_7__SCAN_IN), .A3(
        n4219), .A4(n4221), .ZN(n4163) );
  NAND4_X1 U4834 ( .A1(REG2_REG_13__SCAN_IN), .A2(REG2_REG_5__SCAN_IN), .A3(
        n4306), .A4(n2840), .ZN(n4162) );
  NOR2_X1 U4835 ( .A1(n4163), .A2(n4162), .ZN(n4166) );
  INV_X1 U4836 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4925) );
  NOR2_X1 U4837 ( .A1(n4925), .A2(n4164), .ZN(n4165) );
  NAND4_X1 U4838 ( .A1(n4217), .A2(DATAI_14_), .A3(n4166), .A4(n4165), .ZN(
        n4167) );
  NOR3_X1 U4839 ( .A1(n4169), .A2(n4168), .A3(n4167), .ZN(n4182) );
  NAND4_X1 U4840 ( .A1(D_REG_24__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .A3(
        DATAO_REG_1__SCAN_IN), .A4(n2569), .ZN(n4171) );
  NAND4_X1 U4841 ( .A1(D_REG_16__SCAN_IN), .A2(REG0_REG_19__SCAN_IN), .A3(
        n4637), .A4(n4295), .ZN(n4170) );
  NOR2_X1 U4842 ( .A1(n4171), .A2(n4170), .ZN(n4181) );
  INV_X1 U4843 ( .A(ADDR_REG_16__SCAN_IN), .ZN(n4173) );
  INV_X1 U4844 ( .A(DATAO_REG_0__SCAN_IN), .ZN(n4172) );
  INV_X1 U4845 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4747) );
  NAND4_X1 U4846 ( .A1(n4173), .A2(n4172), .A3(n4269), .A4(n4747), .ZN(n4175)
         );
  NAND4_X1 U4847 ( .A1(n4654), .A2(REG1_REG_25__SCAN_IN), .A3(
        IR_REG_29__SCAN_IN), .A4(DATAI_5_), .ZN(n4174) );
  NOR2_X1 U4848 ( .A1(n4175), .A2(n4174), .ZN(n4180) );
  NAND4_X1 U4849 ( .A1(REG0_REG_10__SCAN_IN), .A2(DATAI_2_), .A3(
        ADDR_REG_0__SCAN_IN), .A4(DATAO_REG_31__SCAN_IN), .ZN(n4178) );
  NAND2_X1 U4850 ( .A1(DATAO_REG_17__SCAN_IN), .A2(D_REG_1__SCAN_IN), .ZN(
        n4176) );
  NOR3_X1 U4851 ( .A1(n4178), .A2(n4177), .A3(n4176), .ZN(n4179) );
  NAND4_X1 U4852 ( .A1(n4182), .A2(n4181), .A3(n4180), .A4(n4179), .ZN(n4185)
         );
  NOR4_X1 U4853 ( .A1(REG1_REG_17__SCAN_IN), .A2(REG1_REG_15__SCAN_IN), .A3(
        ADDR_REG_6__SCAN_IN), .A4(ADDR_REG_7__SCAN_IN), .ZN(n4183) );
  NAND3_X1 U4854 ( .A1(REG2_REG_8__SCAN_IN), .A2(ADDR_REG_10__SCAN_IN), .A3(
        n4183), .ZN(n4184) );
  NOR2_X1 U4855 ( .A1(n4185), .A2(n4184), .ZN(n4191) );
  NOR4_X1 U4856 ( .A1(REG3_REG_6__SCAN_IN), .A2(DATAI_18_), .A3(
        DATAO_REG_16__SCAN_IN), .A4(n4403), .ZN(n4186) );
  INV_X1 U4857 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4405) );
  NAND3_X1 U4858 ( .A1(D_REG_25__SCAN_IN), .A2(n4186), .A3(n4405), .ZN(n4189)
         );
  INV_X1 U4859 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4899) );
  NAND4_X1 U4860 ( .A1(n4187), .A2(D_REG_9__SCAN_IN), .A3(DATAO_REG_8__SCAN_IN), .A4(n4899), .ZN(n4188) );
  NOR2_X1 U4861 ( .A1(n4189), .A2(n4188), .ZN(n4190) );
  AND4_X1 U4862 ( .A1(n4193), .A2(n4192), .A3(n4191), .A4(n4190), .ZN(n4199)
         );
  INV_X1 U4863 ( .A(REG2_REG_31__SCAN_IN), .ZN(n4208) );
  NAND4_X1 U4864 ( .A1(REG1_REG_3__SCAN_IN), .A2(B_REG_SCAN_IN), .A3(
        REG2_REG_23__SCAN_IN), .A4(n4208), .ZN(n4197) );
  INV_X1 U4865 ( .A(REG2_REG_28__SCAN_IN), .ZN(n4206) );
  INV_X1 U4866 ( .A(ADDR_REG_19__SCAN_IN), .ZN(n4201) );
  NAND4_X1 U4867 ( .A1(REG1_REG_19__SCAN_IN), .A2(REG2_REG_17__SCAN_IN), .A3(
        n4206), .A4(n4201), .ZN(n4196) );
  NAND4_X1 U4868 ( .A1(REG3_REG_11__SCAN_IN), .A2(REG3_REG_1__SCAN_IN), .A3(
        ADDR_REG_4__SCAN_IN), .A4(ADDR_REG_5__SCAN_IN), .ZN(n4195) );
  INV_X1 U4869 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4232) );
  NAND4_X1 U4870 ( .A1(DATAI_26_), .A2(DATAI_27_), .A3(REG2_REG_16__SCAN_IN), 
        .A4(n4232), .ZN(n4194) );
  NOR4_X1 U4871 ( .A1(n4197), .A2(n4196), .A3(n4195), .A4(n4194), .ZN(n4198)
         );
  AOI21_X1 U4872 ( .B1(n4199), .B2(n4198), .A(IR_REG_25__SCAN_IN), .ZN(n4200)
         );
  NOR2_X1 U4873 ( .A1(n4200), .A2(keyinput5), .ZN(n4433) );
  INV_X1 U4874 ( .A(keyinput5), .ZN(n4203) );
  XOR2_X1 U4875 ( .A(n4201), .B(keyinput31), .Z(n4202) );
  OAI21_X1 U4876 ( .B1(IR_REG_25__SCAN_IN), .B2(n4203), .A(n4202), .ZN(n4214)
         );
  AOI22_X1 U4877 ( .A1(n4206), .A2(keyinput20), .B1(keyinput40), .B2(n4205), 
        .ZN(n4204) );
  OAI221_X1 U4878 ( .B1(n4206), .B2(keyinput20), .C1(n4205), .C2(keyinput40), 
        .A(n4204), .ZN(n4213) );
  INV_X1 U4879 ( .A(B_REG_SCAN_IN), .ZN(n4209) );
  AOI22_X1 U4880 ( .A1(n4209), .A2(keyinput71), .B1(keyinput111), .B2(n4208), 
        .ZN(n4207) );
  OAI221_X1 U4881 ( .B1(n4209), .B2(keyinput71), .C1(n4208), .C2(keyinput111), 
        .A(n4207), .ZN(n4212) );
  AOI22_X1 U4882 ( .A1(n4656), .A2(keyinput90), .B1(keyinput119), .B2(n2494), 
        .ZN(n4210) );
  OAI221_X1 U4883 ( .B1(n4656), .B2(keyinput90), .C1(n2494), .C2(keyinput119), 
        .A(n4210), .ZN(n4211) );
  NOR4_X1 U4884 ( .A1(n4214), .A2(n4213), .A3(n4212), .A4(n4211), .ZN(n4228)
         );
  AOI22_X1 U4885 ( .A1(n4663), .A2(keyinput7), .B1(keyinput82), .B2(n4672), 
        .ZN(n4215) );
  OAI221_X1 U4886 ( .B1(n4663), .B2(keyinput7), .C1(n4672), .C2(keyinput82), 
        .A(n4215), .ZN(n4226) );
  AOI22_X1 U4887 ( .A1(n4217), .A2(keyinput51), .B1(keyinput102), .B2(n4173), 
        .ZN(n4216) );
  OAI221_X1 U4888 ( .B1(n4217), .B2(keyinput51), .C1(n4173), .C2(keyinput102), 
        .A(n4216), .ZN(n4225) );
  AOI22_X1 U4889 ( .A1(n4219), .A2(keyinput100), .B1(keyinput33), .B2(n3005), 
        .ZN(n4218) );
  OAI221_X1 U4890 ( .B1(n4219), .B2(keyinput100), .C1(n3005), .C2(keyinput33), 
        .A(n4218), .ZN(n4224) );
  AOI22_X1 U4891 ( .A1(n4222), .A2(keyinput26), .B1(keyinput8), .B2(n4221), 
        .ZN(n4220) );
  OAI221_X1 U4892 ( .B1(n4222), .B2(keyinput26), .C1(n4221), .C2(keyinput8), 
        .A(n4220), .ZN(n4223) );
  NOR4_X1 U4893 ( .A1(n4226), .A2(n4225), .A3(n4224), .A4(n4223), .ZN(n4227)
         );
  NAND2_X1 U4894 ( .A1(n4228), .A2(n4227), .ZN(n4432) );
  AOI22_X1 U4895 ( .A1(n4834), .A2(keyinput17), .B1(n4230), .B2(keyinput30), 
        .ZN(n4229) );
  OAI221_X1 U4896 ( .B1(n4834), .B2(keyinput17), .C1(n4230), .C2(keyinput30), 
        .A(n4229), .ZN(n4242) );
  INV_X1 U4897 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4233) );
  AOI22_X1 U4898 ( .A1(n4233), .A2(keyinput81), .B1(keyinput86), .B2(n4232), 
        .ZN(n4231) );
  OAI221_X1 U4899 ( .B1(n4233), .B2(keyinput81), .C1(n4232), .C2(keyinput86), 
        .A(n4231), .ZN(n4241) );
  AOI22_X1 U4900 ( .A1(n3177), .A2(keyinput32), .B1(n4235), .B2(keyinput116), 
        .ZN(n4234) );
  OAI221_X1 U4901 ( .B1(n3177), .B2(keyinput32), .C1(n4235), .C2(keyinput116), 
        .A(n4234), .ZN(n4240) );
  INV_X1 U4902 ( .A(DATAI_26_), .ZN(n4238) );
  AOI22_X1 U4903 ( .A1(n4238), .A2(keyinput2), .B1(n4237), .B2(keyinput125), 
        .ZN(n4236) );
  OAI221_X1 U4904 ( .B1(n4238), .B2(keyinput2), .C1(n4237), .C2(keyinput125), 
        .A(n4236), .ZN(n4239) );
  NOR4_X1 U4905 ( .A1(n4242), .A2(n4241), .A3(n4240), .A4(n4239), .ZN(n4375)
         );
  INV_X1 U4906 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4244) );
  AOI22_X1 U4907 ( .A1(n4637), .A2(keyinput50), .B1(keyinput53), .B2(n4244), 
        .ZN(n4243) );
  OAI221_X1 U4908 ( .B1(n4637), .B2(keyinput50), .C1(n4244), .C2(keyinput53), 
        .A(n4243), .ZN(n4245) );
  INV_X1 U4909 ( .A(n4245), .ZN(n4250) );
  XNOR2_X1 U4910 ( .A(keyinput62), .B(n2450), .ZN(n4248) );
  XNOR2_X1 U4911 ( .A(keyinput15), .B(n4246), .ZN(n4247) );
  NOR2_X1 U4912 ( .A1(n4248), .A2(n4247), .ZN(n4249) );
  NAND2_X1 U4913 ( .A1(n4250), .A2(n4249), .ZN(n4254) );
  AOI22_X1 U4914 ( .A1(n4882), .A2(keyinput37), .B1(n4252), .B2(keyinput6), 
        .ZN(n4251) );
  OAI221_X1 U4915 ( .B1(n4882), .B2(keyinput37), .C1(n4252), .C2(keyinput6), 
        .A(n4251), .ZN(n4253) );
  NOR2_X1 U4916 ( .A1(n4254), .A2(n4253), .ZN(n4275) );
  AOI22_X1 U4917 ( .A1(n4899), .A2(keyinput49), .B1(keyinput48), .B2(n4256), 
        .ZN(n4255) );
  OAI221_X1 U4918 ( .B1(n4899), .B2(keyinput49), .C1(n4256), .C2(keyinput48), 
        .A(n4255), .ZN(n4261) );
  AOI22_X1 U4919 ( .A1(n4259), .A2(keyinput122), .B1(keyinput121), .B2(n4258), 
        .ZN(n4257) );
  OAI221_X1 U4920 ( .B1(n4259), .B2(keyinput122), .C1(n4258), .C2(keyinput121), 
        .A(n4257), .ZN(n4260) );
  NOR2_X1 U4921 ( .A1(n4261), .A2(n4260), .ZN(n4274) );
  INV_X1 U4922 ( .A(D_REG_10__SCAN_IN), .ZN(n4870) );
  INV_X1 U4923 ( .A(D_REG_6__SCAN_IN), .ZN(n4872) );
  AOI22_X1 U4924 ( .A1(n4870), .A2(keyinput63), .B1(keyinput55), .B2(n4872), 
        .ZN(n4262) );
  OAI221_X1 U4925 ( .B1(n4870), .B2(keyinput63), .C1(n4872), .C2(keyinput55), 
        .A(n4262), .ZN(n4266) );
  AOI22_X1 U4926 ( .A1(n4733), .A2(keyinput124), .B1(keyinput126), .B2(n4264), 
        .ZN(n4263) );
  OAI221_X1 U4927 ( .B1(n4733), .B2(keyinput124), .C1(n4264), .C2(keyinput126), 
        .A(n4263), .ZN(n4265) );
  NOR2_X1 U4928 ( .A1(n4266), .A2(n4265), .ZN(n4273) );
  INV_X1 U4929 ( .A(ADDR_REG_10__SCAN_IN), .ZN(n4795) );
  AOI22_X1 U4930 ( .A1(n2265), .A2(keyinput28), .B1(keyinput99), .B2(n4795), 
        .ZN(n4267) );
  OAI221_X1 U4931 ( .B1(n2265), .B2(keyinput28), .C1(n4795), .C2(keyinput99), 
        .A(n4267), .ZN(n4271) );
  AOI22_X1 U4932 ( .A1(n4269), .A2(keyinput42), .B1(n4925), .B2(keyinput45), 
        .ZN(n4268) );
  OAI221_X1 U4933 ( .B1(n4269), .B2(keyinput42), .C1(n4925), .C2(keyinput45), 
        .A(n4268), .ZN(n4270) );
  NOR2_X1 U4934 ( .A1(n4271), .A2(n4270), .ZN(n4272) );
  NAND4_X1 U4935 ( .A1(n4275), .A2(n4274), .A3(n4273), .A4(n4272), .ZN(n4304)
         );
  INV_X1 U4936 ( .A(ADDR_REG_6__SCAN_IN), .ZN(n4278) );
  INV_X1 U4937 ( .A(ADDR_REG_7__SCAN_IN), .ZN(n4277) );
  AOI22_X1 U4938 ( .A1(n4278), .A2(keyinput74), .B1(keyinput1), .B2(n4277), 
        .ZN(n4276) );
  OAI221_X1 U4939 ( .B1(n4278), .B2(keyinput74), .C1(n4277), .C2(keyinput1), 
        .A(n4276), .ZN(n4283) );
  INV_X1 U4940 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4281) );
  AOI22_X1 U4941 ( .A1(n4281), .A2(keyinput115), .B1(n4280), .B2(keyinput123), 
        .ZN(n4279) );
  OAI221_X1 U4942 ( .B1(n4281), .B2(keyinput115), .C1(n4280), .C2(keyinput123), 
        .A(n4279), .ZN(n4282) );
  NOR2_X1 U4943 ( .A1(n4283), .A2(n4282), .ZN(n4302) );
  AOI22_X1 U4944 ( .A1(n4654), .A2(keyinput61), .B1(n4866), .B2(keyinput57), 
        .ZN(n4284) );
  OAI221_X1 U4945 ( .B1(n4654), .B2(keyinput61), .C1(n4866), .C2(keyinput57), 
        .A(n4284), .ZN(n4288) );
  INV_X1 U4946 ( .A(ADDR_REG_4__SCAN_IN), .ZN(n4286) );
  AOI22_X1 U4947 ( .A1(n4286), .A2(keyinput76), .B1(keyinput98), .B2(n3981), 
        .ZN(n4285) );
  OAI221_X1 U4948 ( .B1(n4286), .B2(keyinput76), .C1(n3981), .C2(keyinput98), 
        .A(n4285), .ZN(n4287) );
  NOR2_X1 U4949 ( .A1(n4288), .A2(n4287), .ZN(n4301) );
  INV_X1 U4950 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4290) );
  INV_X1 U4951 ( .A(D_REG_3__SCAN_IN), .ZN(n4874) );
  AOI22_X1 U4952 ( .A1(n4290), .A2(keyinput21), .B1(n4874), .B2(keyinput13), 
        .ZN(n4289) );
  OAI221_X1 U4953 ( .B1(n4290), .B2(keyinput21), .C1(n4874), .C2(keyinput13), 
        .A(n4289), .ZN(n4293) );
  INV_X1 U4954 ( .A(D_REG_24__SCAN_IN), .ZN(n4863) );
  AOI22_X1 U4955 ( .A1(n2569), .A2(keyinput25), .B1(n4863), .B2(keyinput24), 
        .ZN(n4291) );
  OAI221_X1 U4956 ( .B1(n2569), .B2(keyinput25), .C1(n4863), .C2(keyinput24), 
        .A(n4291), .ZN(n4292) );
  NOR2_X1 U4957 ( .A1(n4293), .A2(n4292), .ZN(n4300) );
  INV_X1 U4958 ( .A(D_REG_16__SCAN_IN), .ZN(n4868) );
  AOI22_X1 U4959 ( .A1(n4295), .A2(keyinput56), .B1(n4868), .B2(keyinput54), 
        .ZN(n4294) );
  OAI221_X1 U4960 ( .B1(n4295), .B2(keyinput56), .C1(n4868), .C2(keyinput54), 
        .A(n4294), .ZN(n4298) );
  INV_X1 U4961 ( .A(ADDR_REG_0__SCAN_IN), .ZN(n4296) );
  XNOR2_X1 U4962 ( .A(n4296), .B(keyinput75), .ZN(n4297) );
  NOR2_X1 U4963 ( .A1(n4298), .A2(n4297), .ZN(n4299) );
  NAND4_X1 U4964 ( .A1(n4302), .A2(n4301), .A3(n4300), .A4(n4299), .ZN(n4303)
         );
  NOR2_X1 U4965 ( .A1(n4304), .A2(n4303), .ZN(n4374) );
  AOI22_X1 U4966 ( .A1(n3140), .A2(keyinput80), .B1(n4306), .B2(keyinput66), 
        .ZN(n4305) );
  OAI221_X1 U4967 ( .B1(n3140), .B2(keyinput80), .C1(n4306), .C2(keyinput66), 
        .A(n4305), .ZN(n4317) );
  AOI22_X1 U4968 ( .A1(n2840), .A2(keyinput16), .B1(n2612), .B2(keyinput10), 
        .ZN(n4307) );
  OAI221_X1 U4969 ( .B1(n2840), .B2(keyinput16), .C1(n2612), .C2(keyinput10), 
        .A(n4307), .ZN(n4316) );
  INV_X1 U4970 ( .A(REG0_REG_29__SCAN_IN), .ZN(n4310) );
  AOI22_X1 U4971 ( .A1(n4310), .A2(keyinput59), .B1(keyinput91), .B2(n4309), 
        .ZN(n4308) );
  OAI221_X1 U4972 ( .B1(n4310), .B2(keyinput59), .C1(n4309), .C2(keyinput91), 
        .A(n4308), .ZN(n4315) );
  AOI22_X1 U4973 ( .A1(n4313), .A2(keyinput0), .B1(n4312), .B2(keyinput52), 
        .ZN(n4311) );
  OAI221_X1 U4974 ( .B1(n4313), .B2(keyinput0), .C1(n4312), .C2(keyinput52), 
        .A(n4311), .ZN(n4314) );
  NOR4_X1 U4975 ( .A1(n4317), .A2(n4316), .A3(n4315), .A4(n4314), .ZN(n4373)
         );
  INV_X1 U4976 ( .A(REG0_REG_10__SCAN_IN), .ZN(n4319) );
  AOI22_X1 U4977 ( .A1(n4320), .A2(keyinput29), .B1(n4319), .B2(keyinput22), 
        .ZN(n4318) );
  OAI221_X1 U4978 ( .B1(n4320), .B2(keyinput29), .C1(n4319), .C2(keyinput22), 
        .A(n4318), .ZN(n4325) );
  AOI22_X1 U4979 ( .A1(n4323), .A2(keyinput64), .B1(n4322), .B2(keyinput60), 
        .ZN(n4321) );
  OAI221_X1 U4980 ( .B1(n4323), .B2(keyinput64), .C1(n4322), .C2(keyinput60), 
        .A(n4321), .ZN(n4324) );
  NOR2_X1 U4981 ( .A1(n4325), .A2(n4324), .ZN(n4347) );
  AOI22_X1 U4982 ( .A1(n4328), .A2(keyinput114), .B1(n4327), .B2(keyinput117), 
        .ZN(n4326) );
  OAI221_X1 U4983 ( .B1(n4328), .B2(keyinput114), .C1(n4327), .C2(keyinput117), 
        .A(n4326), .ZN(n4333) );
  INV_X1 U4984 ( .A(DATAI_30_), .ZN(n4330) );
  AOI22_X1 U4985 ( .A1(n4331), .A2(keyinput12), .B1(keyinput14), .B2(n4330), 
        .ZN(n4329) );
  OAI221_X1 U4986 ( .B1(n4331), .B2(keyinput12), .C1(n4330), .C2(keyinput14), 
        .A(n4329), .ZN(n4332) );
  NOR2_X1 U4987 ( .A1(n4333), .A2(n4332), .ZN(n4346) );
  INV_X1 U4988 ( .A(keyinput38), .ZN(n4334) );
  XNOR2_X1 U4989 ( .A(n4335), .B(n4334), .ZN(n4345) );
  INV_X1 U4990 ( .A(D_REG_30__SCAN_IN), .ZN(n4860) );
  AOI22_X1 U4991 ( .A1(n4860), .A2(keyinput43), .B1(keyinput3), .B2(n4337), 
        .ZN(n4336) );
  OAI221_X1 U4992 ( .B1(n4860), .B2(keyinput43), .C1(n4337), .C2(keyinput3), 
        .A(n4336), .ZN(n4343) );
  XNOR2_X1 U4993 ( .A(DATAI_2_), .B(keyinput67), .ZN(n4341) );
  XNOR2_X1 U4994 ( .A(IR_REG_1__SCAN_IN), .B(keyinput36), .ZN(n4340) );
  XNOR2_X1 U4995 ( .A(IR_REG_0__SCAN_IN), .B(keyinput4), .ZN(n4339) );
  XNOR2_X1 U4996 ( .A(IR_REG_10__SCAN_IN), .B(keyinput87), .ZN(n4338) );
  NAND4_X1 U4997 ( .A1(n4341), .A2(n4340), .A3(n4339), .A4(n4338), .ZN(n4342)
         );
  NOR2_X1 U4998 ( .A1(n4343), .A2(n4342), .ZN(n4344) );
  NAND4_X1 U4999 ( .A1(n4347), .A2(n4346), .A3(n4345), .A4(n4344), .ZN(n4371)
         );
  AOI22_X1 U5000 ( .A1(n4865), .A2(keyinput41), .B1(keyinput34), .B2(n4747), 
        .ZN(n4348) );
  OAI221_X1 U5001 ( .B1(n4865), .B2(keyinput41), .C1(n4747), .C2(keyinput34), 
        .A(n4348), .ZN(n4354) );
  XNOR2_X1 U5002 ( .A(keyinput103), .B(REG1_REG_0__SCAN_IN), .ZN(n4352) );
  XNOR2_X1 U5003 ( .A(IR_REG_7__SCAN_IN), .B(keyinput9), .ZN(n4351) );
  XNOR2_X1 U5004 ( .A(keyinput120), .B(IR_REG_23__SCAN_IN), .ZN(n4350) );
  INV_X1 U5005 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4906) );
  XNOR2_X1 U5006 ( .A(keyinput79), .B(REG0_REG_2__SCAN_IN), .ZN(n4349) );
  NAND4_X1 U5007 ( .A1(n4352), .A2(n4351), .A3(n4350), .A4(n4349), .ZN(n4353)
         );
  NOR2_X1 U5008 ( .A1(n4354), .A2(n4353), .ZN(n4369) );
  INV_X1 U5009 ( .A(D_REG_9__SCAN_IN), .ZN(n4871) );
  XNOR2_X1 U5010 ( .A(n4871), .B(keyinput44), .ZN(n4356) );
  INV_X1 U5011 ( .A(D_REG_5__SCAN_IN), .ZN(n4873) );
  XNOR2_X1 U5012 ( .A(n4873), .B(keyinput18), .ZN(n4355) );
  NOR2_X1 U5013 ( .A1(n4356), .A2(n4355), .ZN(n4368) );
  XNOR2_X1 U5014 ( .A(IR_REG_2__SCAN_IN), .B(keyinput118), .ZN(n4360) );
  XNOR2_X1 U5015 ( .A(IR_REG_16__SCAN_IN), .B(keyinput95), .ZN(n4359) );
  XNOR2_X1 U5016 ( .A(REG3_REG_26__SCAN_IN), .B(keyinput83), .ZN(n4358) );
  XNOR2_X1 U5017 ( .A(IR_REG_22__SCAN_IN), .B(keyinput107), .ZN(n4357) );
  NAND4_X1 U5018 ( .A1(n4360), .A2(n4359), .A3(n4358), .A4(n4357), .ZN(n4366)
         );
  XNOR2_X1 U5019 ( .A(REG3_REG_6__SCAN_IN), .B(keyinput113), .ZN(n4364) );
  XNOR2_X1 U5020 ( .A(IR_REG_28__SCAN_IN), .B(keyinput58), .ZN(n4363) );
  XNOR2_X1 U5021 ( .A(IR_REG_13__SCAN_IN), .B(keyinput112), .ZN(n4362) );
  XNOR2_X1 U5022 ( .A(DATAI_5_), .B(keyinput46), .ZN(n4361) );
  NAND4_X1 U5023 ( .A1(n4364), .A2(n4363), .A3(n4362), .A4(n4361), .ZN(n4365)
         );
  NOR2_X1 U5024 ( .A1(n4366), .A2(n4365), .ZN(n4367) );
  NAND3_X1 U5025 ( .A1(n4369), .A2(n4368), .A3(n4367), .ZN(n4370) );
  NOR2_X1 U5026 ( .A1(n4371), .A2(n4370), .ZN(n4372) );
  NAND4_X1 U5027 ( .A1(n4375), .A2(n4374), .A3(n4373), .A4(n4372), .ZN(n4431)
         );
  INV_X1 U5028 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4377) );
  AOI22_X1 U5029 ( .A1(n4378), .A2(keyinput96), .B1(n4377), .B2(keyinput92), 
        .ZN(n4376) );
  OAI221_X1 U5030 ( .B1(n4378), .B2(keyinput96), .C1(n4377), .C2(keyinput92), 
        .A(n4376), .ZN(n4386) );
  INV_X1 U5031 ( .A(D_REG_27__SCAN_IN), .ZN(n4861) );
  AOI22_X1 U5032 ( .A1(n4861), .A2(keyinput94), .B1(keyinput93), .B2(n4380), 
        .ZN(n4379) );
  OAI221_X1 U5033 ( .B1(n4861), .B2(keyinput94), .C1(n4380), .C2(keyinput93), 
        .A(n4379), .ZN(n4385) );
  INV_X1 U5034 ( .A(DATAI_23_), .ZN(n4878) );
  AOI22_X1 U5035 ( .A1(n2594), .A2(keyinput89), .B1(keyinput88), .B2(n4878), 
        .ZN(n4381) );
  OAI221_X1 U5036 ( .B1(n2594), .B2(keyinput89), .C1(n4878), .C2(keyinput88), 
        .A(n4381), .ZN(n4384) );
  INV_X1 U5037 ( .A(D_REG_31__SCAN_IN), .ZN(n4859) );
  AOI22_X1 U5038 ( .A1(n4859), .A2(keyinput84), .B1(n2741), .B2(keyinput85), 
        .ZN(n4382) );
  OAI221_X1 U5039 ( .B1(n4859), .B2(keyinput84), .C1(n2741), .C2(keyinput85), 
        .A(n4382), .ZN(n4383) );
  NOR4_X1 U5040 ( .A1(n4386), .A2(n4385), .A3(n4384), .A4(n4383), .ZN(n4429)
         );
  INV_X1 U5041 ( .A(REG0_REG_18__SCAN_IN), .ZN(n4742) );
  AOI22_X1 U5042 ( .A1(n2596), .A2(keyinput78), .B1(n4742), .B2(keyinput77), 
        .ZN(n4387) );
  OAI221_X1 U5043 ( .B1(n2596), .B2(keyinput78), .C1(n4742), .C2(keyinput77), 
        .A(n4387), .ZN(n4399) );
  AOI22_X1 U5044 ( .A1(n4389), .A2(keyinput73), .B1(n4869), .B2(keyinput72), 
        .ZN(n4388) );
  OAI221_X1 U5045 ( .B1(n4389), .B2(keyinput73), .C1(n4869), .C2(keyinput72), 
        .A(n4388), .ZN(n4398) );
  INV_X1 U5046 ( .A(DATAI_9_), .ZN(n4392) );
  AOI22_X1 U5047 ( .A1(n4392), .A2(keyinput68), .B1(n4391), .B2(keyinput70), 
        .ZN(n4390) );
  OAI221_X1 U5048 ( .B1(n4392), .B2(keyinput68), .C1(n4391), .C2(keyinput70), 
        .A(n4390), .ZN(n4397) );
  AOI22_X1 U5049 ( .A1(n4395), .A2(keyinput69), .B1(n4394), .B2(keyinput65), 
        .ZN(n4393) );
  OAI221_X1 U5050 ( .B1(n4395), .B2(keyinput69), .C1(n4394), .C2(keyinput65), 
        .A(n4393), .ZN(n4396) );
  NOR4_X1 U5051 ( .A1(n4399), .A2(n4398), .A3(n4397), .A4(n4396), .ZN(n4428)
         );
  AOI22_X1 U5052 ( .A1(n4172), .A2(keyinput108), .B1(n4867), .B2(keyinput110), 
        .ZN(n4400) );
  OAI221_X1 U5053 ( .B1(n4172), .B2(keyinput108), .C1(n4867), .C2(keyinput110), 
        .A(n4400), .ZN(n4412) );
  AOI22_X1 U5054 ( .A1(n4403), .A2(keyinput106), .B1(keyinput109), .B2(n4402), 
        .ZN(n4401) );
  OAI221_X1 U5055 ( .B1(n4403), .B2(keyinput106), .C1(n4402), .C2(keyinput109), 
        .A(n4401), .ZN(n4411) );
  INV_X1 U5056 ( .A(D_REG_25__SCAN_IN), .ZN(n4862) );
  AOI22_X1 U5057 ( .A1(n4862), .A2(keyinput105), .B1(keyinput104), .B2(n4405), 
        .ZN(n4404) );
  OAI221_X1 U5058 ( .B1(n4862), .B2(keyinput105), .C1(n4405), .C2(keyinput104), 
        .A(n4404), .ZN(n4410) );
  INV_X1 U5059 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4407) );
  AOI22_X1 U5060 ( .A1(n4408), .A2(keyinput101), .B1(n4407), .B2(keyinput97), 
        .ZN(n4406) );
  OAI221_X1 U5061 ( .B1(n4408), .B2(keyinput101), .C1(n4407), .C2(keyinput97), 
        .A(n4406), .ZN(n4409) );
  NOR4_X1 U5062 ( .A1(n4412), .A2(n4411), .A3(n4410), .A4(n4409), .ZN(n4427)
         );
  INV_X1 U5063 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4714) );
  INV_X1 U5064 ( .A(IR_REG_4__SCAN_IN), .ZN(n4414) );
  AOI22_X1 U5065 ( .A1(n4714), .A2(keyinput19), .B1(n4414), .B2(keyinput23), 
        .ZN(n4413) );
  OAI221_X1 U5066 ( .B1(n4714), .B2(keyinput19), .C1(n4414), .C2(keyinput23), 
        .A(n4413), .ZN(n4425) );
  INV_X1 U5067 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4695) );
  AOI22_X1 U5068 ( .A1(n4695), .A2(keyinput47), .B1(keyinput27), .B2(n4416), 
        .ZN(n4415) );
  OAI221_X1 U5069 ( .B1(n4695), .B2(keyinput47), .C1(n4416), .C2(keyinput27), 
        .A(n4415), .ZN(n4424) );
  INV_X1 U5070 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4418) );
  AOI22_X1 U5071 ( .A1(n4419), .A2(keyinput39), .B1(n4418), .B2(keyinput127), 
        .ZN(n4417) );
  OAI221_X1 U5072 ( .B1(n4419), .B2(keyinput39), .C1(n4418), .C2(keyinput127), 
        .A(n4417), .ZN(n4423) );
  AOI22_X1 U5073 ( .A1(n4421), .A2(keyinput11), .B1(n4666), .B2(keyinput35), 
        .ZN(n4420) );
  OAI221_X1 U5074 ( .B1(n4421), .B2(keyinput11), .C1(n4666), .C2(keyinput35), 
        .A(n4420), .ZN(n4422) );
  NOR4_X1 U5075 ( .A1(n4425), .A2(n4424), .A3(n4423), .A4(n4422), .ZN(n4426)
         );
  NAND4_X1 U5076 ( .A1(n4429), .A2(n4428), .A3(n4427), .A4(n4426), .ZN(n4430)
         );
  NOR4_X1 U5077 ( .A1(n4433), .A2(n4432), .A3(n4431), .A4(n4430), .ZN(n4434)
         );
  XNOR2_X1 U5078 ( .A(n4435), .B(n4434), .ZN(U3266) );
  NAND2_X1 U5079 ( .A1(n4457), .A2(n4456), .ZN(n4455) );
  NAND2_X1 U5080 ( .A1(n4455), .A2(n4437), .ZN(n4438) );
  XNOR2_X1 U5081 ( .A(n4438), .B(n4447), .ZN(n4721) );
  INV_X1 U5082 ( .A(n4642), .ZN(n4441) );
  INV_X1 U5083 ( .A(n4439), .ZN(n4440) );
  AOI21_X1 U5084 ( .B1(n2369), .B2(n4441), .A(n4440), .ZN(n4719) );
  AOI22_X1 U5085 ( .A1(n4719), .A2(n4576), .B1(n4442), .B2(n4574), .ZN(n4454)
         );
  INV_X1 U5086 ( .A(n4456), .ZN(n4460) );
  NAND2_X1 U5087 ( .A1(n4459), .A2(n4460), .ZN(n4458) );
  NAND2_X1 U5088 ( .A1(n4458), .A2(n4445), .ZN(n4446) );
  XOR2_X1 U5089 ( .A(n4447), .B(n4446), .Z(n4452) );
  NOR2_X1 U5090 ( .A1(n4448), .A2(n4604), .ZN(n4451) );
  OAI22_X1 U5091 ( .A1(n4483), .A2(n4545), .B1(n4449), .B2(n4565), .ZN(n4450)
         );
  MUX2_X1 U5092 ( .A(n4233), .B(n4639), .S(n4585), .Z(n4453) );
  OAI211_X1 U5093 ( .C1(n4721), .C2(n4588), .A(n4454), .B(n4453), .ZN(U3267)
         );
  OAI21_X1 U5094 ( .B1(n4457), .B2(n4456), .A(n4455), .ZN(n4725) );
  OAI21_X1 U5095 ( .B1(n4460), .B2(n4459), .A(n4458), .ZN(n4461) );
  NAND2_X1 U5096 ( .A1(n4461), .A2(n4607), .ZN(n4468) );
  NAND2_X1 U5097 ( .A1(n4462), .A2(n4599), .ZN(n4464) );
  NAND2_X1 U5098 ( .A1(n4500), .A2(n4601), .ZN(n4463) );
  OAI211_X1 U5099 ( .C1(n4465), .C2(n4604), .A(n4464), .B(n4463), .ZN(n4466)
         );
  INV_X1 U5100 ( .A(n4466), .ZN(n4467) );
  NAND2_X1 U5101 ( .A1(n4468), .A2(n4467), .ZN(n4645) );
  NOR2_X1 U5102 ( .A1(n4476), .A2(n4469), .ZN(n4643) );
  OR3_X1 U5103 ( .A1(n4642), .A2(n4643), .A3(n4594), .ZN(n4472) );
  AOI22_X1 U5104 ( .A1(n4470), .A2(n4574), .B1(REG2_REG_22__SCAN_IN), .B2(
        n4609), .ZN(n4471) );
  NAND2_X1 U5105 ( .A1(n4472), .A2(n4471), .ZN(n4473) );
  AOI21_X1 U5106 ( .B1(n4645), .B2(n4585), .A(n4473), .ZN(n4474) );
  OAI21_X1 U5107 ( .B1(n4725), .B2(n4588), .A(n4474), .ZN(U3268) );
  XOR2_X1 U5108 ( .A(n4478), .B(n4475), .Z(n4731) );
  AOI21_X1 U5109 ( .B1(n4480), .B2(n2143), .A(n4476), .ZN(n4729) );
  AOI22_X1 U5110 ( .A1(n4729), .A2(n4576), .B1(n4477), .B2(n4574), .ZN(n4488)
         );
  INV_X1 U5111 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4486) );
  XNOR2_X1 U5112 ( .A(n4479), .B(n4478), .ZN(n4485) );
  AOI22_X1 U5113 ( .A1(n4481), .A2(n4601), .B1(n4480), .B2(n4599), .ZN(n4482)
         );
  OAI21_X1 U5114 ( .B1(n4483), .B2(n4604), .A(n4482), .ZN(n4484) );
  AOI21_X1 U5115 ( .B1(n4485), .B2(n4607), .A(n4484), .ZN(n4726) );
  MUX2_X1 U5116 ( .A(n4486), .B(n4726), .S(n4585), .Z(n4487) );
  OAI211_X1 U5117 ( .C1(n4731), .C2(n4588), .A(n4488), .B(n4487), .ZN(U3269)
         );
  XNOR2_X1 U5118 ( .A(n4489), .B(n4493), .ZN(n4651) );
  OAI22_X1 U5119 ( .A1(n4490), .A2(n4545), .B1(n4565), .B2(n4504), .ZN(n4499)
         );
  INV_X1 U5120 ( .A(n4517), .ZN(n4558) );
  AOI21_X1 U5121 ( .B1(n4558), .B2(n4492), .A(n4491), .ZN(n4495) );
  INV_X1 U5122 ( .A(n4493), .ZN(n4494) );
  XNOR2_X1 U5123 ( .A(n4495), .B(n4494), .ZN(n4497) );
  NOR2_X1 U5124 ( .A1(n4497), .A2(n4496), .ZN(n4498) );
  AOI211_X1 U5125 ( .C1(n4559), .C2(n4500), .A(n4499), .B(n4498), .ZN(n4501)
         );
  OAI21_X1 U5126 ( .B1(n4651), .B2(n4502), .A(n4501), .ZN(n4652) );
  NAND2_X1 U5127 ( .A1(n4652), .A2(n4585), .ZN(n4510) );
  INV_X1 U5128 ( .A(n4503), .ZN(n4513) );
  OAI21_X1 U5129 ( .B1(n4513), .B2(n4504), .A(n2143), .ZN(n4735) );
  INV_X1 U5130 ( .A(n4735), .ZN(n4508) );
  INV_X1 U5131 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4505) );
  OAI22_X1 U5132 ( .A1(n4506), .A2(n4592), .B1(n4585), .B2(n4505), .ZN(n4507)
         );
  AOI21_X1 U5133 ( .B1(n4508), .B2(n4576), .A(n4507), .ZN(n4509) );
  OAI211_X1 U5134 ( .C1(n4651), .C2(n4511), .A(n4510), .B(n4509), .ZN(U3270)
         );
  XNOR2_X1 U5135 ( .A(n4512), .B(n4523), .ZN(n4741) );
  INV_X1 U5136 ( .A(n4536), .ZN(n4514) );
  AOI21_X1 U5137 ( .B1(n4525), .B2(n4514), .A(n4513), .ZN(n4739) );
  AOI22_X1 U5138 ( .A1(n4739), .A2(n4576), .B1(n4515), .B2(n4574), .ZN(n4532)
         );
  INV_X1 U5139 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4530) );
  OR2_X1 U5140 ( .A1(n4517), .A2(n4516), .ZN(n4519) );
  NAND2_X1 U5141 ( .A1(n4519), .A2(n4518), .ZN(n4542) );
  INV_X1 U5142 ( .A(n4520), .ZN(n4522) );
  OAI21_X1 U5143 ( .B1(n4542), .B2(n4522), .A(n4521), .ZN(n4524) );
  XNOR2_X1 U5144 ( .A(n4524), .B(n4523), .ZN(n4529) );
  AOI22_X1 U5145 ( .A1(n4560), .A2(n4601), .B1(n4525), .B2(n4599), .ZN(n4526)
         );
  OAI21_X1 U5146 ( .B1(n4527), .B2(n4604), .A(n4526), .ZN(n4528) );
  AOI21_X1 U5147 ( .B1(n4529), .B2(n4607), .A(n4528), .ZN(n4736) );
  MUX2_X1 U5148 ( .A(n4530), .B(n4736), .S(n4585), .Z(n4531) );
  OAI211_X1 U5149 ( .C1(n4741), .C2(n4588), .A(n4532), .B(n4531), .ZN(U3271)
         );
  XOR2_X1 U5150 ( .A(n4540), .B(n4533), .Z(n4745) );
  NAND2_X1 U5151 ( .A1(n4553), .A2(n2666), .ZN(n4534) );
  NAND2_X1 U5152 ( .A1(n4534), .A2(n4924), .ZN(n4535) );
  NOR2_X1 U5153 ( .A1(n4536), .A2(n4535), .ZN(n4659) );
  OAI22_X1 U5154 ( .A1(n4585), .A2(n2898), .B1(n4537), .B2(n4592), .ZN(n4538)
         );
  AOI21_X1 U5155 ( .B1(n4659), .B2(n4539), .A(n4538), .ZN(n4551) );
  INV_X1 U5156 ( .A(n4540), .ZN(n4541) );
  XNOR2_X1 U5157 ( .A(n4542), .B(n4541), .ZN(n4543) );
  NAND2_X1 U5158 ( .A1(n4543), .A2(n4607), .ZN(n4549) );
  OAI22_X1 U5159 ( .A1(n4582), .A2(n4545), .B1(n4544), .B2(n4565), .ZN(n4546)
         );
  AOI21_X1 U5160 ( .B1(n4559), .B2(n4547), .A(n4546), .ZN(n4548) );
  NAND2_X1 U5161 ( .A1(n4549), .A2(n4548), .ZN(n4660) );
  NAND2_X1 U5162 ( .A1(n4660), .A2(n4585), .ZN(n4550) );
  OAI211_X1 U5163 ( .C1(n4745), .C2(n4588), .A(n4551), .B(n4550), .ZN(U3272)
         );
  XNOR2_X1 U5164 ( .A(n4552), .B(n4557), .ZN(n4751) );
  INV_X1 U5165 ( .A(n4553), .ZN(n4554) );
  AOI21_X1 U5166 ( .B1(n4555), .B2(n4572), .A(n4554), .ZN(n4748) );
  AOI22_X1 U5167 ( .A1(n4748), .A2(n4576), .B1(n4556), .B2(n4574), .ZN(n4569)
         );
  XNOR2_X1 U5168 ( .A(n4558), .B(n4557), .ZN(n4567) );
  NAND2_X1 U5169 ( .A1(n4560), .A2(n4559), .ZN(n4563) );
  NAND2_X1 U5170 ( .A1(n4561), .A2(n4601), .ZN(n4562) );
  OAI211_X1 U5171 ( .C1(n4565), .C2(n4564), .A(n4563), .B(n4562), .ZN(n4566)
         );
  AOI21_X1 U5172 ( .B1(n4567), .B2(n4607), .A(n4566), .ZN(n4746) );
  MUX2_X1 U5173 ( .A(n4205), .B(n4746), .S(n4585), .Z(n4568) );
  OAI211_X1 U5174 ( .C1(n4751), .C2(n4588), .A(n4569), .B(n4568), .ZN(U3273)
         );
  XNOR2_X1 U5175 ( .A(n4570), .B(n4577), .ZN(n4759) );
  INV_X1 U5176 ( .A(n4571), .ZN(n4591) );
  INV_X1 U5177 ( .A(n4572), .ZN(n4573) );
  AOI21_X1 U5178 ( .B1(n4579), .B2(n4591), .A(n4573), .ZN(n4756) );
  AOI22_X1 U5179 ( .A1(n4756), .A2(n4576), .B1(n4575), .B2(n4574), .ZN(n4587)
         );
  XNOR2_X1 U5180 ( .A(n4578), .B(n4577), .ZN(n4584) );
  AOI22_X1 U5181 ( .A1(n4580), .A2(n4601), .B1(n4579), .B2(n4599), .ZN(n4581)
         );
  OAI21_X1 U5182 ( .B1(n4582), .B2(n4604), .A(n4581), .ZN(n4583) );
  AOI21_X1 U5183 ( .B1(n4584), .B2(n4607), .A(n4583), .ZN(n4752) );
  MUX2_X1 U5184 ( .A(n4834), .B(n4752), .S(n4585), .Z(n4586) );
  OAI211_X1 U5185 ( .C1(n4759), .C2(n4588), .A(n4587), .B(n4586), .ZN(U3274)
         );
  XNOR2_X1 U5186 ( .A(n4589), .B(n4597), .ZN(n4761) );
  NAND2_X1 U5187 ( .A1(n4678), .A2(n4600), .ZN(n4590) );
  NAND2_X1 U5188 ( .A1(n4591), .A2(n4590), .ZN(n4767) );
  OAI22_X1 U5189 ( .A1(n4767), .A2(n4594), .B1(n4593), .B2(n4592), .ZN(n4612)
         );
  NAND2_X1 U5190 ( .A1(n4596), .A2(n4595), .ZN(n4598) );
  XOR2_X1 U5191 ( .A(n4598), .B(n4597), .Z(n4608) );
  AOI22_X1 U5192 ( .A1(n4602), .A2(n4601), .B1(n4600), .B2(n4599), .ZN(n4603)
         );
  OAI21_X1 U5193 ( .B1(n4605), .B2(n4604), .A(n4603), .ZN(n4606) );
  AOI21_X1 U5194 ( .B1(n4608), .B2(n4607), .A(n4606), .ZN(n4763) );
  INV_X1 U5195 ( .A(n4763), .ZN(n4610) );
  MUX2_X1 U5196 ( .A(n4610), .B(REG2_REG_15__SCAN_IN), .S(n4609), .Z(n4611) );
  AOI211_X1 U5197 ( .C1(n4613), .C2(n4761), .A(n4612), .B(n4611), .ZN(n4614)
         );
  INV_X1 U5198 ( .A(n4614), .ZN(U3275) );
  NOR2_X1 U5199 ( .A1(n4941), .A2(n4615), .ZN(n4616) );
  AOI21_X1 U5200 ( .B1(n4941), .B2(n4690), .A(n4616), .ZN(n4617) );
  OAI21_X1 U5201 ( .B1(n4693), .B2(n4675), .A(n4617), .ZN(U3549) );
  NAND2_X1 U5202 ( .A1(n4618), .A2(n4667), .ZN(n4620) );
  NAND2_X1 U5203 ( .A1(n4939), .A2(REG1_REG_30__SCAN_IN), .ZN(n4619) );
  OAI211_X1 U5204 ( .C1(n4694), .C2(n4939), .A(n4620), .B(n4619), .ZN(U3548)
         );
  INV_X1 U5205 ( .A(n4622), .ZN(n4623) );
  OAI21_X1 U5206 ( .B1(n4625), .B2(n4900), .A(n4624), .ZN(n4700) );
  MUX2_X1 U5207 ( .A(REG1_REG_27__SCAN_IN), .B(n4700), .S(n4941), .Z(n4626) );
  INV_X1 U5208 ( .A(n4626), .ZN(n4627) );
  AOI21_X1 U5209 ( .B1(n4629), .B2(n4928), .A(n4628), .ZN(n4704) );
  MUX2_X1 U5210 ( .A(n4630), .B(n4704), .S(n4941), .Z(n4631) );
  OAI21_X1 U5211 ( .B1(n4675), .B2(n4707), .A(n4631), .ZN(U3544) );
  MUX2_X1 U5212 ( .A(REG1_REG_25__SCAN_IN), .B(n4708), .S(n4941), .Z(n4633) );
  AOI21_X1 U5213 ( .B1(n4710), .B2(n4667), .A(n4633), .ZN(n4634) );
  OAI21_X1 U5214 ( .B1(n4712), .B2(n4670), .A(n4634), .ZN(U3543) );
  AOI21_X1 U5215 ( .B1(n4636), .B2(n4928), .A(n4635), .ZN(n4713) );
  MUX2_X1 U5216 ( .A(n4637), .B(n4713), .S(n4941), .Z(n4638) );
  OAI21_X1 U5217 ( .B1(n4675), .B2(n4716), .A(n4638), .ZN(U3542) );
  AOI21_X1 U5218 ( .B1(n4719), .B2(n4667), .A(n4640), .ZN(n4641) );
  OAI21_X1 U5219 ( .B1(n4721), .B2(n4670), .A(n4641), .ZN(U3541) );
  NOR3_X1 U5220 ( .A1(n4643), .A2(n4642), .A3(n4900), .ZN(n4644) );
  NOR2_X1 U5221 ( .A1(n4645), .A2(n4644), .ZN(n4722) );
  MUX2_X1 U5222 ( .A(n4646), .B(n4722), .S(n4941), .Z(n4647) );
  OAI21_X1 U5223 ( .B1(n4725), .B2(n4670), .A(n4647), .ZN(U3540) );
  MUX2_X1 U5224 ( .A(n4648), .B(n4726), .S(n4941), .Z(n4650) );
  NAND2_X1 U5225 ( .A1(n4729), .A2(n4667), .ZN(n4649) );
  OAI211_X1 U5226 ( .C1(n4731), .C2(n4670), .A(n4650), .B(n4649), .ZN(U3539)
         );
  INV_X1 U5227 ( .A(n4894), .ZN(n4915) );
  INV_X1 U5228 ( .A(n4651), .ZN(n4653) );
  AOI21_X1 U5229 ( .B1(n4915), .B2(n4653), .A(n4652), .ZN(n4732) );
  MUX2_X1 U5230 ( .A(n4654), .B(n4732), .S(n4941), .Z(n4655) );
  OAI21_X1 U5231 ( .B1(n4675), .B2(n4735), .A(n4655), .ZN(U3538) );
  MUX2_X1 U5232 ( .A(n4656), .B(n4736), .S(n4941), .Z(n4658) );
  NAND2_X1 U5233 ( .A1(n4739), .A2(n4667), .ZN(n4657) );
  OAI211_X1 U5234 ( .C1(n4741), .C2(n4670), .A(n4658), .B(n4657), .ZN(U3537)
         );
  NOR2_X1 U5235 ( .A1(n4660), .A2(n4659), .ZN(n4743) );
  MUX2_X1 U5236 ( .A(n4743), .B(n4661), .S(n4939), .Z(n4662) );
  OAI21_X1 U5237 ( .B1(n4745), .B2(n4670), .A(n4662), .ZN(U3536) );
  MUX2_X1 U5238 ( .A(n4663), .B(n4746), .S(n4941), .Z(n4665) );
  NAND2_X1 U5239 ( .A1(n4748), .A2(n4667), .ZN(n4664) );
  OAI211_X1 U5240 ( .C1(n4751), .C2(n4670), .A(n4665), .B(n4664), .ZN(U3535)
         );
  MUX2_X1 U5241 ( .A(n4666), .B(n4752), .S(n4941), .Z(n4669) );
  NAND2_X1 U5242 ( .A1(n4756), .A2(n4667), .ZN(n4668) );
  OAI211_X1 U5243 ( .C1(n4759), .C2(n4670), .A(n4669), .B(n4668), .ZN(U3534)
         );
  NAND2_X1 U5244 ( .A1(n4761), .A2(n4671), .ZN(n4674) );
  MUX2_X1 U5245 ( .A(n4763), .B(n4672), .S(n4939), .Z(n4673) );
  OAI211_X1 U5246 ( .C1(n4675), .C2(n4767), .A(n4674), .B(n4673), .ZN(U3533)
         );
  INV_X1 U5247 ( .A(n4676), .ZN(n4681) );
  NAND3_X1 U5248 ( .A1(n4678), .A2(n4924), .A3(n4677), .ZN(n4679) );
  OAI211_X1 U5249 ( .C1(n4681), .C2(n4894), .A(n4680), .B(n4679), .ZN(n4768)
         );
  MUX2_X1 U5250 ( .A(REG1_REG_14__SCAN_IN), .B(n4768), .S(n4941), .Z(U3532) );
  NAND2_X1 U5251 ( .A1(n4682), .A2(n4928), .ZN(n4683) );
  OAI211_X1 U5252 ( .C1(n4900), .C2(n4685), .A(n4684), .B(n4683), .ZN(n4769)
         );
  MUX2_X1 U5253 ( .A(REG1_REG_13__SCAN_IN), .B(n4769), .S(n4941), .Z(U3531) );
  NAND2_X1 U5254 ( .A1(n4686), .A2(n4928), .ZN(n4687) );
  OAI211_X1 U5255 ( .C1(n4900), .C2(n4689), .A(n4688), .B(n4687), .ZN(n4770)
         );
  MUX2_X1 U5256 ( .A(n4770), .B(REG1_REG_11__SCAN_IN), .S(n4939), .Z(U3529) );
  NAND2_X1 U5257 ( .A1(n4932), .A2(n4690), .ZN(n4692) );
  NAND2_X1 U5258 ( .A1(n4930), .A2(REG0_REG_31__SCAN_IN), .ZN(n4691) );
  OAI211_X1 U5259 ( .C1(n4693), .C2(n4766), .A(n4692), .B(n4691), .ZN(U3517)
         );
  MUX2_X1 U5260 ( .A(n4695), .B(n4694), .S(n4932), .Z(n4696) );
  OAI21_X1 U5261 ( .B1(n4697), .B2(n4766), .A(n4696), .ZN(U3516) );
  MUX2_X1 U5262 ( .A(REG0_REG_27__SCAN_IN), .B(n4700), .S(n4932), .Z(n4701) );
  INV_X1 U5263 ( .A(n4701), .ZN(n4702) );
  OAI21_X1 U5264 ( .B1(n4703), .B2(n4758), .A(n4702), .ZN(U3513) );
  INV_X1 U5265 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4705) );
  MUX2_X1 U5266 ( .A(n4705), .B(n4704), .S(n4932), .Z(n4706) );
  MUX2_X1 U5267 ( .A(REG0_REG_25__SCAN_IN), .B(n4708), .S(n4932), .Z(n4709) );
  AOI21_X1 U5268 ( .B1(n4710), .B2(n4755), .A(n4709), .ZN(n4711) );
  OAI21_X1 U5269 ( .B1(n4712), .B2(n4758), .A(n4711), .ZN(U3511) );
  MUX2_X1 U5270 ( .A(n4714), .B(n4713), .S(n4932), .Z(n4715) );
  OAI21_X1 U5271 ( .B1(n4716), .B2(n4766), .A(n4715), .ZN(U3510) );
  MUX2_X1 U5272 ( .A(REG0_REG_23__SCAN_IN), .B(n4717), .S(n4932), .Z(n4718) );
  AOI21_X1 U5273 ( .B1(n4719), .B2(n4755), .A(n4718), .ZN(n4720) );
  OAI21_X1 U5274 ( .B1(n4721), .B2(n4758), .A(n4720), .ZN(U3509) );
  INV_X1 U5275 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4723) );
  MUX2_X1 U5276 ( .A(n4723), .B(n4722), .S(n4932), .Z(n4724) );
  OAI21_X1 U5277 ( .B1(n4725), .B2(n4758), .A(n4724), .ZN(U3508) );
  INV_X1 U5278 ( .A(n4726), .ZN(n4727) );
  MUX2_X1 U5279 ( .A(REG0_REG_21__SCAN_IN), .B(n4727), .S(n4932), .Z(n4728) );
  AOI21_X1 U5280 ( .B1(n4729), .B2(n4755), .A(n4728), .ZN(n4730) );
  OAI21_X1 U5281 ( .B1(n4731), .B2(n4758), .A(n4730), .ZN(U3507) );
  MUX2_X1 U5282 ( .A(n4733), .B(n4732), .S(n4932), .Z(n4734) );
  OAI21_X1 U5283 ( .B1(n4735), .B2(n4766), .A(n4734), .ZN(U3506) );
  INV_X1 U5284 ( .A(n4736), .ZN(n4737) );
  MUX2_X1 U5285 ( .A(REG0_REG_19__SCAN_IN), .B(n4737), .S(n4932), .Z(n4738) );
  AOI21_X1 U5286 ( .B1(n4739), .B2(n4755), .A(n4738), .ZN(n4740) );
  OAI21_X1 U5287 ( .B1(n4741), .B2(n4758), .A(n4740), .ZN(U3505) );
  MUX2_X1 U5288 ( .A(n4743), .B(n4742), .S(n4930), .Z(n4744) );
  OAI21_X1 U5289 ( .B1(n4745), .B2(n4758), .A(n4744), .ZN(U3503) );
  MUX2_X1 U5290 ( .A(n4747), .B(n4746), .S(n4932), .Z(n4750) );
  NAND2_X1 U5291 ( .A1(n4748), .A2(n4755), .ZN(n4749) );
  OAI211_X1 U5292 ( .C1(n4751), .C2(n4758), .A(n4750), .B(n4749), .ZN(U3501)
         );
  INV_X1 U5293 ( .A(n4752), .ZN(n4753) );
  MUX2_X1 U5294 ( .A(REG0_REG_16__SCAN_IN), .B(n4753), .S(n4932), .Z(n4754) );
  AOI21_X1 U5295 ( .B1(n4756), .B2(n4755), .A(n4754), .ZN(n4757) );
  OAI21_X1 U5296 ( .B1(n4759), .B2(n4758), .A(n4757), .ZN(U3499) );
  NAND2_X1 U5297 ( .A1(n4761), .A2(n4760), .ZN(n4765) );
  INV_X1 U5298 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4762) );
  MUX2_X1 U5299 ( .A(n4763), .B(n4762), .S(n4930), .Z(n4764) );
  OAI211_X1 U5300 ( .C1(n4767), .C2(n4766), .A(n4765), .B(n4764), .ZN(U3497)
         );
  MUX2_X1 U5301 ( .A(REG0_REG_14__SCAN_IN), .B(n4768), .S(n4932), .Z(U3495) );
  MUX2_X1 U5302 ( .A(REG0_REG_13__SCAN_IN), .B(n4769), .S(n4932), .Z(U3493) );
  MUX2_X1 U5303 ( .A(REG0_REG_11__SCAN_IN), .B(n4770), .S(n4932), .Z(U3489) );
  MUX2_X1 U5304 ( .A(n4771), .B(DATAI_30_), .S(U3149), .Z(U3322) );
  MUX2_X1 U5305 ( .A(n4772), .B(DATAI_29_), .S(U3149), .Z(U3323) );
  MUX2_X1 U5306 ( .A(n4773), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U5307 ( .A(DATAI_25_), .B(n4774), .S(STATE_REG_SCAN_IN), .Z(U3327)
         );
  MUX2_X1 U5308 ( .A(n2818), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U5309 ( .A(DATAI_18_), .B(n4775), .S(STATE_REG_SCAN_IN), .Z(U3334)
         );
  MUX2_X1 U5310 ( .A(n2210), .B(DATAI_11_), .S(U3149), .Z(U3341) );
  MUX2_X1 U5311 ( .A(DATAI_9_), .B(n4777), .S(STATE_REG_SCAN_IN), .Z(U3343) );
  MUX2_X1 U5312 ( .A(DATAI_8_), .B(n4778), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U5313 ( .A(DATAI_5_), .B(n4779), .S(STATE_REG_SCAN_IN), .Z(U3347) );
  MUX2_X1 U5314 ( .A(n4780), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5315 ( .A(n4781), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  MUX2_X1 U5316 ( .A(DATAI_0_), .B(IR_REG_0__SCAN_IN), .S(STATE_REG_SCAN_IN), 
        .Z(U3352) );
  INV_X1 U5317 ( .A(DATAI_28_), .ZN(n4782) );
  AOI22_X1 U5318 ( .A1(STATE_REG_SCAN_IN), .A2(n4783), .B1(n4782), .B2(U3149), 
        .ZN(U3324) );
  INV_X1 U5319 ( .A(n4784), .ZN(n4787) );
  INV_X1 U5320 ( .A(n4785), .ZN(n4786) );
  AOI21_X1 U5321 ( .B1(n2963), .B2(n4787), .A(n4786), .ZN(n4788) );
  XNOR2_X1 U5322 ( .A(n4788), .B(IR_REG_0__SCAN_IN), .ZN(n4790) );
  AOI22_X1 U5323 ( .A1(n4851), .A2(ADDR_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4789) );
  OAI21_X1 U5324 ( .B1(n4791), .B2(n4790), .A(n4789), .ZN(U3240) );
  OAI211_X1 U5325 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4793), .A(n2901), .B(n4792), .ZN(n4794) );
  OAI21_X1 U5326 ( .B1(n4844), .B2(n4795), .A(n4794), .ZN(n4796) );
  NOR2_X1 U5327 ( .A1(n4797), .A2(n4796), .ZN(n4801) );
  OAI211_X1 U5328 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4799), .A(n4852), .B(n4798), .ZN(n4800) );
  OAI211_X1 U5329 ( .C1(n4858), .C2(n2359), .A(n4801), .B(n4800), .ZN(U3250)
         );
  OAI211_X1 U5330 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4803), .A(n2901), .B(n4802), .ZN(n4805) );
  NAND2_X1 U5331 ( .A1(n4805), .A2(n4804), .ZN(n4806) );
  AOI21_X1 U5332 ( .B1(n4851), .B2(ADDR_REG_12__SCAN_IN), .A(n4806), .ZN(n4810) );
  OAI211_X1 U5333 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4808), .A(n4852), .B(n4807), .ZN(n4809) );
  OAI211_X1 U5334 ( .C1(n4858), .C2(n4886), .A(n4810), .B(n4809), .ZN(U3252)
         );
  INV_X1 U5335 ( .A(n4811), .ZN(n4817) );
  AOI21_X1 U5336 ( .B1(n4885), .B2(n2612), .A(n4812), .ZN(n4815) );
  OAI21_X1 U5337 ( .B1(n4815), .B2(n4814), .A(n2901), .ZN(n4813) );
  AOI21_X1 U5338 ( .B1(n4815), .B2(n4814), .A(n4813), .ZN(n4816) );
  AOI211_X1 U5339 ( .C1(n4851), .C2(ADDR_REG_13__SCAN_IN), .A(n4817), .B(n4816), .ZN(n4822) );
  OAI211_X1 U5340 ( .C1(n4820), .C2(n4819), .A(n4852), .B(n4818), .ZN(n4821)
         );
  OAI211_X1 U5341 ( .C1(n4858), .C2(n4885), .A(n4822), .B(n4821), .ZN(U3253)
         );
  INV_X1 U5342 ( .A(n4823), .ZN(n4828) );
  AOI211_X1 U5343 ( .C1(n4826), .C2(n4825), .A(n4824), .B(n4845), .ZN(n4827)
         );
  AOI211_X1 U5344 ( .C1(n4851), .C2(ADDR_REG_14__SCAN_IN), .A(n4828), .B(n4827), .ZN(n4832) );
  OAI211_X1 U5345 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4830), .A(n4852), .B(n4829), .ZN(n4831) );
  OAI211_X1 U5346 ( .C1(n4858), .C2(n4883), .A(n4832), .B(n4831), .ZN(U3254)
         );
  OAI21_X1 U5347 ( .B1(n4835), .B2(n4834), .A(n4833), .ZN(n4841) );
  AOI21_X1 U5348 ( .B1(REG1_REG_16__SCAN_IN), .B2(n4837), .A(n4836), .ZN(n4839) );
  OAI22_X1 U5349 ( .A1(n4839), .A2(n4838), .B1(n4881), .B2(n4858), .ZN(n4840)
         );
  AOI21_X1 U5350 ( .B1(n2901), .B2(n4841), .A(n4840), .ZN(n4843) );
  OAI211_X1 U5351 ( .C1(n4173), .C2(n4844), .A(n4843), .B(n4842), .ZN(U3256)
         );
  AOI221_X1 U5352 ( .B1(n4848), .B2(n4847), .C1(n4846), .C2(n4847), .A(n4845), 
        .ZN(n4849) );
  AOI211_X1 U5353 ( .C1(n4851), .C2(ADDR_REG_17__SCAN_IN), .A(n4850), .B(n4849), .ZN(n4857) );
  OAI221_X1 U5354 ( .B1(n4855), .B2(n4854), .C1(n4855), .C2(n4853), .A(n4852), 
        .ZN(n4856) );
  OAI211_X1 U5355 ( .C1(n4858), .C2(n4880), .A(n4857), .B(n4856), .ZN(U3257)
         );
  NOR2_X1 U5356 ( .A1(n4875), .A2(n4859), .ZN(U3291) );
  NOR2_X1 U5357 ( .A1(n4875), .A2(n4860), .ZN(U3292) );
  AND2_X1 U5358 ( .A1(D_REG_29__SCAN_IN), .A2(n4876), .ZN(U3293) );
  AND2_X1 U5359 ( .A1(D_REG_28__SCAN_IN), .A2(n4876), .ZN(U3294) );
  NOR2_X1 U5360 ( .A1(n4875), .A2(n4861), .ZN(U3295) );
  AND2_X1 U5361 ( .A1(D_REG_26__SCAN_IN), .A2(n4876), .ZN(U3296) );
  NOR2_X1 U5362 ( .A1(n4875), .A2(n4862), .ZN(U3297) );
  NOR2_X1 U5363 ( .A1(n4875), .A2(n4863), .ZN(U3298) );
  NOR2_X1 U5364 ( .A1(n4875), .A2(n4864), .ZN(U3299) );
  NOR2_X1 U5365 ( .A1(n4875), .A2(n4865), .ZN(U3300) );
  NOR2_X1 U5366 ( .A1(n4875), .A2(n4866), .ZN(U3301) );
  AND2_X1 U5367 ( .A1(D_REG_20__SCAN_IN), .A2(n4876), .ZN(U3302) );
  AND2_X1 U5368 ( .A1(D_REG_19__SCAN_IN), .A2(n4876), .ZN(U3303) );
  NOR2_X1 U5369 ( .A1(n4875), .A2(n4867), .ZN(U3304) );
  AND2_X1 U5370 ( .A1(D_REG_17__SCAN_IN), .A2(n4876), .ZN(U3305) );
  NOR2_X1 U5371 ( .A1(n4875), .A2(n4868), .ZN(U3306) );
  NOR2_X1 U5372 ( .A1(n4875), .A2(n4869), .ZN(U3307) );
  AND2_X1 U5373 ( .A1(D_REG_14__SCAN_IN), .A2(n4876), .ZN(U3308) );
  AND2_X1 U5374 ( .A1(D_REG_13__SCAN_IN), .A2(n4876), .ZN(U3309) );
  AND2_X1 U5375 ( .A1(D_REG_12__SCAN_IN), .A2(n4876), .ZN(U3310) );
  AND2_X1 U5376 ( .A1(D_REG_11__SCAN_IN), .A2(n4876), .ZN(U3311) );
  NOR2_X1 U5377 ( .A1(n4875), .A2(n4870), .ZN(U3312) );
  NOR2_X1 U5378 ( .A1(n4875), .A2(n4871), .ZN(U3313) );
  AND2_X1 U5379 ( .A1(D_REG_8__SCAN_IN), .A2(n4876), .ZN(U3314) );
  AND2_X1 U5380 ( .A1(D_REG_7__SCAN_IN), .A2(n4876), .ZN(U3315) );
  NOR2_X1 U5381 ( .A1(n4875), .A2(n4872), .ZN(U3316) );
  NOR2_X1 U5382 ( .A1(n4875), .A2(n4873), .ZN(U3317) );
  AND2_X1 U5383 ( .A1(D_REG_4__SCAN_IN), .A2(n4876), .ZN(U3318) );
  NOR2_X1 U5384 ( .A1(n4875), .A2(n4874), .ZN(U3319) );
  AND2_X1 U5385 ( .A1(D_REG_2__SCAN_IN), .A2(n4876), .ZN(U3320) );
  AOI21_X1 U5386 ( .B1(U3149), .B2(n4878), .A(n4877), .ZN(U3329) );
  AOI22_X1 U5387 ( .A1(STATE_REG_SCAN_IN), .A2(n4880), .B1(n4879), .B2(U3149), 
        .ZN(U3335) );
  AOI22_X1 U5388 ( .A1(STATE_REG_SCAN_IN), .A2(n4881), .B1(n2641), .B2(U3149), 
        .ZN(U3336) );
  AOI22_X1 U5389 ( .A1(STATE_REG_SCAN_IN), .A2(n4883), .B1(n4882), .B2(U3149), 
        .ZN(U3338) );
  INV_X1 U5390 ( .A(DATAI_13_), .ZN(n4884) );
  AOI22_X1 U5391 ( .A1(STATE_REG_SCAN_IN), .A2(n4885), .B1(n4884), .B2(U3149), 
        .ZN(U3339) );
  AOI22_X1 U5392 ( .A1(STATE_REG_SCAN_IN), .A2(n4886), .B1(n2596), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U5393 ( .A(DATAI_10_), .ZN(n4887) );
  AOI22_X1 U5394 ( .A1(STATE_REG_SCAN_IN), .A2(n2359), .B1(n4887), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5395 ( .A(n4888), .ZN(n4891) );
  INV_X1 U5396 ( .A(n4889), .ZN(n4890) );
  AOI211_X1 U5397 ( .C1(n4915), .C2(n4892), .A(n4891), .B(n4890), .ZN(n4933)
         );
  INV_X1 U5398 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4893) );
  AOI22_X1 U5399 ( .A1(n4932), .A2(n4933), .B1(n4893), .B2(n4930), .ZN(U3467)
         );
  NOR2_X1 U5400 ( .A1(n4895), .A2(n4894), .ZN(n4897) );
  AOI211_X1 U5401 ( .C1(n4924), .C2(n4898), .A(n4897), .B(n4896), .ZN(n4934)
         );
  AOI22_X1 U5402 ( .A1(n4932), .A2(n4934), .B1(n4899), .B2(n4930), .ZN(U3469)
         );
  NOR3_X1 U5403 ( .A1(n4902), .A2(n4901), .A3(n4900), .ZN(n4904) );
  AOI211_X1 U5404 ( .C1(n4915), .C2(n4905), .A(n4904), .B(n4903), .ZN(n4935)
         );
  AOI22_X1 U5405 ( .A1(n4932), .A2(n4935), .B1(n4906), .B2(n4930), .ZN(U3471)
         );
  AOI22_X1 U5406 ( .A1(n4908), .A2(n4915), .B1(n4924), .B2(n4907), .ZN(n4909)
         );
  AND2_X1 U5407 ( .A1(n4910), .A2(n4909), .ZN(n4936) );
  INV_X1 U5408 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4911) );
  AOI22_X1 U5409 ( .A1(n4932), .A2(n4936), .B1(n4911), .B2(n4930), .ZN(U3473)
         );
  INV_X1 U5410 ( .A(n4912), .ZN(n4914) );
  AOI211_X1 U5411 ( .C1(n4916), .C2(n4915), .A(n4914), .B(n4913), .ZN(n4937)
         );
  INV_X1 U5412 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4917) );
  AOI22_X1 U5413 ( .A1(n4932), .A2(n4937), .B1(n4917), .B2(n4930), .ZN(U3475)
         );
  INV_X1 U5414 ( .A(n4928), .ZN(n4918) );
  NOR2_X1 U5415 ( .A1(n4919), .A2(n4918), .ZN(n4922) );
  INV_X1 U5416 ( .A(n4920), .ZN(n4921) );
  AOI211_X1 U5417 ( .C1(n4924), .C2(n4923), .A(n4922), .B(n4921), .ZN(n4938)
         );
  AOI22_X1 U5418 ( .A1(n4932), .A2(n4938), .B1(n4925), .B2(n4930), .ZN(U3477)
         );
  AOI211_X1 U5419 ( .C1(n4929), .C2(n4928), .A(n4927), .B(n4926), .ZN(n4940)
         );
  INV_X1 U5420 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4931) );
  AOI22_X1 U5421 ( .A1(n4932), .A2(n4940), .B1(n4931), .B2(n4930), .ZN(U3481)
         );
  AOI22_X1 U5422 ( .A1(n4941), .A2(n4933), .B1(n2963), .B2(n4939), .ZN(U3518)
         );
  AOI22_X1 U5423 ( .A1(n4941), .A2(n4934), .B1(n2838), .B2(n4939), .ZN(U3519)
         );
  AOI22_X1 U5424 ( .A1(n4941), .A2(n4935), .B1(n2840), .B2(n4939), .ZN(U3520)
         );
  AOI22_X1 U5425 ( .A1(n4941), .A2(n4936), .B1(n2494), .B2(n4939), .ZN(U3521)
         );
  AOI22_X1 U5426 ( .A1(n4941), .A2(n4937), .B1(n2503), .B2(n4939), .ZN(U3522)
         );
  AOI22_X1 U5427 ( .A1(n4941), .A2(n4938), .B1(n2842), .B2(n4939), .ZN(U3523)
         );
  AOI22_X1 U5428 ( .A1(n4941), .A2(n4940), .B1(n3005), .B2(n4939), .ZN(U3525)
         );
  NAND2_X1 U2986 ( .A1(n2147), .A2(n2498), .ZN(n3963) );
  CLKBUF_X1 U2455 ( .A(n2479), .Z(n2495) );
  CLKBUF_X1 U2730 ( .A(n3634), .Z(n3682) );
endmodule

