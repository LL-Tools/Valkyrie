

module b15_C_gen_AntiSAT_k_128_3 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, 
        U3209, U3208, U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, 
        U3199, U3198, U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, 
        U3189, U3188, U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, 
        U3452, U3180, U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, 
        U3171, U3170, U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, 
        U3161, U3160, U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, 
        U3151, U3453, U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, 
        U3142, U3141, U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, 
        U3132, U3131, U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, 
        U3122, U3121, U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, 
        U3112, U3111, U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, 
        U3102, U3101, U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, 
        U3092, U3091, U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, 
        U3082, U3081, U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, 
        U3072, U3071, U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, 
        U3062, U3061, U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, 
        U3052, U3051, U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, 
        U3042, U3041, U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, 
        U3032, U3031, U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, 
        U3022, U3021, U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, 
        U3463, U3464, U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, 
        U3011, U3010, U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, 
        U3001, U3000, U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, 
        U2991, U2990, U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, 
        U2981, U2980, U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, 
        U2971, U2970, U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, 
        U2961, U2960, U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, 
        U2951, U2950, U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, 
        U2941, U2940, U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, 
        U2931, U2930, U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, 
        U2921, U2920, U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, 
        U2911, U2910, U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, 
        U2901, U2900, U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, 
        U2891, U2890, U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, 
        U2881, U2880, U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, 
        U2871, U2870, U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, 
        U2861, U2860, U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, 
        U2851, U2850, U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, 
        U2841, U2840, U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, 
        U2831, U2830, U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, 
        U2821, U2820, U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, 
        U2811, U2810, U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, 
        U2801, U2800, U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, 
        U3470, U2793, U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, 
        U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1,
         keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6,
         keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11,
         keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16,
         keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21,
         keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26,
         keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31,
         keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36,
         keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41,
         keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46,
         keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51,
         keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56,
         keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61,
         keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823;

  AND2_X1 U3434 ( .A1(n5987), .A2(n5749), .ZN(n4158) );
  INV_X1 U3435 ( .A(n3789), .ZN(n6249) );
  OR2_X1 U3436 ( .A1(n3817), .A2(n4297), .ZN(n4324) );
  AND2_X1 U3437 ( .A1(n4295), .A2(n4294), .ZN(n4297) );
  CLKBUF_X1 U3439 ( .A(n5342), .Z(n3011) );
  CLKBUF_X2 U3440 ( .A(n3180), .Z(n5326) );
  CLKBUF_X2 U3441 ( .A(n3323), .Z(n5340) );
  CLKBUF_X2 U3442 ( .A(n3213), .Z(n4108) );
  CLKBUF_X1 U3443 ( .A(n4234), .Z(n3006) );
  AND4_X1 U3444 ( .A1(n3110), .A2(n3109), .A3(n3108), .A4(n3107), .ZN(n3121)
         );
  AND4_X1 U34450 ( .A1(n3114), .A2(n3113), .A3(n3112), .A4(n3111), .ZN(n3120)
         );
  AND4_X1 U34460 ( .A1(n3118), .A2(n3117), .A3(n3116), .A4(n3115), .ZN(n3119)
         );
  AND2_X1 U34470 ( .A1(n3094), .A2(n3048), .ZN(n3323) );
  AND2_X2 U34480 ( .A1(n3077), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3048) );
  NOR2_X2 U3449 ( .A1(n3796), .A2(n6498), .ZN(n3985) );
  INV_X1 U34510 ( .A(n6823), .ZN(n2986) );
  BUF_X1 U34530 ( .A(n3224), .Z(n4232) );
  INV_X1 U34550 ( .A(n3789), .ZN(n2988) );
  AND2_X1 U34560 ( .A1(n3013), .A2(n3230), .ZN(n3261) );
  OR2_X1 U3457 ( .A1(n5609), .A2(n5808), .ZN(n5806) );
  INV_X1 U3458 ( .A(n3513), .ZN(n3789) );
  INV_X1 U34590 ( .A(n6187), .ZN(n6160) );
  AND2_X1 U34600 ( .A1(n5593), .A2(n5497), .ZN(n5513) );
  AOI21_X1 U34610 ( .B1(n5514), .B2(n5595), .A(n5513), .ZN(n5704) );
  CLKBUF_X1 U34620 ( .A(n3017), .Z(n2990) );
  NAND2_X2 U34630 ( .A1(n4319), .A2(n4320), .ZN(n4446) );
  NAND2_X2 U34640 ( .A1(n3819), .A2(n3818), .ZN(n4319) );
  NAND2_X2 U34650 ( .A1(n3444), .A2(n3443), .ZN(n4975) );
  NAND2_X4 U3466 ( .A1(n3074), .A2(n3185), .ZN(n3222) );
  AND4_X2 U3467 ( .A1(n3184), .A2(n3183), .A3(n3182), .A4(n3181), .ZN(n3185)
         );
  NOR2_X2 U34680 ( .A1(n3724), .A2(n5452), .ZN(n3611) );
  OAI21_X2 U34690 ( .B1(n3711), .B2(EBX_REG_1__SCAN_IN), .A(n3622), .ZN(n3040)
         );
  AND2_X1 U34700 ( .A1(n3048), .A2(n4248), .ZN(n2987) );
  AND2_X1 U34710 ( .A1(n3048), .A2(n4248), .ZN(n3213) );
  OAI21_X2 U34730 ( .B1(n5513), .B2(n5499), .A(n5498), .ZN(n5587) );
  INV_X2 U34740 ( .A(n3223), .ZN(n3796) );
  OAI21_X2 U3476 ( .B1(n5484), .B2(n5431), .A(n5430), .ZN(n5669) );
  AND2_X1 U3477 ( .A1(n2992), .A2(n2993), .ZN(n5677) );
  CLKBUF_X1 U3478 ( .A(n3786), .Z(n5735) );
  NAND2_X1 U3479 ( .A1(n5047), .A2(n5048), .ZN(n5049) );
  NAND2_X1 U3480 ( .A1(n3496), .A2(n3419), .ZN(n3513) );
  NAND2_X1 U3481 ( .A1(n3376), .A2(n3375), .ZN(n4334) );
  NAND2_X1 U3482 ( .A1(n3736), .A2(n3615), .ZN(n6283) );
  NAND2_X1 U3483 ( .A1(n5640), .A2(n4305), .ZN(n5983) );
  INV_X2 U3484 ( .A(n4975), .ZN(n3446) );
  AND3_X1 U3485 ( .A1(n3206), .A2(n3205), .A3(n3204), .ZN(n3258) );
  OR2_X1 U3486 ( .A1(n4524), .A2(n6499), .ZN(n3364) );
  INV_X1 U3487 ( .A(n4232), .ZN(n4524) );
  INV_X2 U3488 ( .A(n3221), .ZN(n3239) );
  NAND4_X1 U3489 ( .A1(n3099), .A2(n3100), .A3(n3101), .A4(n3102), .ZN(n4441)
         );
  AND4_X1 U3490 ( .A1(n3167), .A2(n3166), .A3(n3165), .A4(n3164), .ZN(n3173)
         );
  AND4_X1 U3491 ( .A1(n3092), .A2(n3091), .A3(n3090), .A4(n3089), .ZN(n3100)
         );
  AND4_X1 U3492 ( .A1(n3217), .A2(n3216), .A3(n3215), .A4(n3214), .ZN(n3218)
         );
  BUF_X2 U3493 ( .A(n3008), .Z(n3391) );
  CLKBUF_X2 U3494 ( .A(n3324), .Z(n5349) );
  CLKBUF_X2 U3495 ( .A(n3283), .Z(n5258) );
  BUF_X2 U3497 ( .A(n3207), .Z(n3012) );
  BUF_X2 U3498 ( .A(n3190), .Z(n3005) );
  NAND2_X1 U3499 ( .A1(n6592), .A2(n6498), .ZN(n5875) );
  XNOR2_X1 U3500 ( .A(n4164), .B(n4163), .ZN(n4172) );
  OAI22_X1 U3501 ( .A1(n4162), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .B1(n5714), .B2(n3792), .ZN(n3793) );
  INV_X1 U3502 ( .A(n5426), .ZN(n5647) );
  INV_X1 U3503 ( .A(n5676), .ZN(n5700) );
  OAI21_X1 U3504 ( .B1(n5658), .B2(n6267), .A(n4177), .ZN(n4178) );
  XNOR2_X1 U3505 ( .A(n5415), .B(n5414), .ZN(n5642) );
  AND2_X1 U3506 ( .A1(n5595), .A2(n5594), .ZN(n5984) );
  XNOR2_X1 U3507 ( .A(n5430), .B(n3075), .ZN(n5426) );
  AND2_X1 U3508 ( .A1(n5593), .A2(n5412), .ZN(n5415) );
  AND2_X1 U3509 ( .A1(n5593), .A2(n5429), .ZN(n5484) );
  NAND2_X1 U3510 ( .A1(n5593), .A2(n5411), .ZN(n5430) );
  OAI21_X1 U3511 ( .B1(n5744), .B2(n3521), .A(n3522), .ZN(n3523) );
  NAND2_X1 U3512 ( .A1(n5234), .A2(n3946), .ZN(n5635) );
  OAI21_X1 U3513 ( .B1(n6247), .B2(n3052), .A(n3050), .ZN(n3056) );
  NAND2_X1 U3514 ( .A1(n3061), .A2(n3064), .ZN(n5177) );
  NAND2_X1 U3515 ( .A1(n3932), .A2(n3931), .ZN(n3946) );
  INV_X1 U3516 ( .A(n3051), .ZN(n3050) );
  OAI21_X1 U3517 ( .B1(n5194), .B2(n3053), .A(n5192), .ZN(n3052) );
  NAND2_X1 U3518 ( .A1(n5489), .A2(n3628), .ZN(n3774) );
  AND2_X1 U3519 ( .A1(n3698), .A2(n3043), .ZN(n5596) );
  NAND2_X1 U3520 ( .A1(n3417), .A2(n3482), .ZN(n3496) );
  NAND2_X1 U3521 ( .A1(n3404), .A2(n3473), .ZN(n3483) );
  NAND2_X1 U3522 ( .A1(n3377), .A2(n3021), .ZN(n3474) );
  NOR2_X1 U3523 ( .A1(n6243), .A2(n6221), .ZN(n6242) );
  CLKBUF_X1 U3524 ( .A(n4337), .Z(n6167) );
  NAND2_X2 U3525 ( .A1(n4775), .A2(n4289), .ZN(n4422) );
  NAND2_X1 U3526 ( .A1(n3291), .A2(n3290), .ZN(n3295) );
  NOR2_X1 U3527 ( .A1(n5015), .A2(n5016), .ZN(n5134) );
  NAND2_X1 U3528 ( .A1(n3362), .A2(n3361), .ZN(n4614) );
  OAI21_X1 U3529 ( .B1(n3272), .B2(n4256), .A(n3276), .ZN(n3355) );
  CLKBUF_X1 U3530 ( .A(n3271), .Z(n3272) );
  AND2_X1 U3531 ( .A1(n3340), .A2(n3440), .ZN(n3341) );
  AND2_X1 U3532 ( .A1(n3188), .A2(n3538), .ZN(n3220) );
  AND2_X1 U3533 ( .A1(n3202), .A2(n3201), .ZN(n3267) );
  XNOR2_X1 U3534 ( .A(n3040), .B(n4230), .ZN(n6196) );
  NAND2_X1 U3535 ( .A1(n3562), .A2(n4524), .ZN(n3578) );
  NAND2_X2 U3536 ( .A1(n3796), .A2(n3222), .ZN(n5452) );
  NAND2_X1 U3537 ( .A1(n3241), .A2(n3174), .ZN(n3186) );
  INV_X1 U3538 ( .A(n4441), .ZN(n3013) );
  OR2_X1 U3539 ( .A1(n3307), .A2(n3306), .ZN(n3435) );
  AND3_X2 U3540 ( .A1(n3173), .A2(n3172), .A3(n3171), .ZN(n3223) );
  NAND2_X2 U3541 ( .A1(n3219), .A2(n3218), .ZN(n4431) );
  OR2_X1 U3542 ( .A1(n3335), .A2(n3334), .ZN(n3505) );
  AND4_X1 U3543 ( .A1(n3134), .A2(n3133), .A3(n3132), .A4(n3131), .ZN(n3140)
         );
  AND4_X1 U3544 ( .A1(n3155), .A2(n3154), .A3(n3153), .A4(n3152), .ZN(n3161)
         );
  AND4_X1 U3545 ( .A1(n3098), .A2(n3097), .A3(n3096), .A4(n3095), .ZN(n3099)
         );
  AND4_X1 U3546 ( .A1(n3130), .A2(n3129), .A3(n3128), .A4(n3127), .ZN(n3141)
         );
  AND4_X1 U3547 ( .A1(n3211), .A2(n3210), .A3(n3209), .A4(n3208), .ZN(n3219)
         );
  AND3_X1 U3548 ( .A1(n3170), .A2(n3169), .A3(n3168), .ZN(n3172) );
  AND2_X1 U3549 ( .A1(n3147), .A2(n3020), .ZN(n3163) );
  AND4_X1 U3550 ( .A1(n3106), .A2(n3105), .A3(n3104), .A4(n3103), .ZN(n3122)
         );
  AND4_X1 U3551 ( .A1(n3138), .A2(n3137), .A3(n3136), .A4(n3135), .ZN(n3139)
         );
  AND4_X1 U3552 ( .A1(n3151), .A2(n3150), .A3(n3149), .A4(n3148), .ZN(n3162)
         );
  AND4_X1 U3553 ( .A1(n3126), .A2(n3125), .A3(n3124), .A4(n3123), .ZN(n3142)
         );
  AND4_X1 U3554 ( .A1(n3087), .A2(n3086), .A3(n3085), .A4(n3084), .ZN(n3101)
         );
  AND4_X1 U3555 ( .A1(n3083), .A2(n3082), .A3(n3081), .A4(n3080), .ZN(n3102)
         );
  AND4_X1 U3556 ( .A1(n3159), .A2(n3158), .A3(n3157), .A4(n3156), .ZN(n3160)
         );
  INV_X2 U3557 ( .A(n6267), .ZN(n5749) );
  BUF_X2 U3558 ( .A(n3189), .Z(n4119) );
  BUF_X2 U3559 ( .A(n3175), .Z(n5348) );
  AND2_X4 U3560 ( .A1(n3094), .A2(n4473), .ZN(n3207) );
  AND2_X2 U3561 ( .A1(n3078), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3093)
         );
  AND2_X2 U3562 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4473) );
  INV_X1 U3563 ( .A(n3226), .ZN(n2991) );
  NAND2_X1 U3564 ( .A1(n3786), .A2(n2995), .ZN(n2992) );
  OR2_X1 U3565 ( .A1(n2994), .A2(n3527), .ZN(n2993) );
  INV_X1 U3566 ( .A(n3529), .ZN(n2994) );
  AND2_X1 U3567 ( .A1(n3525), .A2(n3529), .ZN(n2995) );
  BUF_X1 U3568 ( .A(n3354), .Z(n2996) );
  INV_X1 U3569 ( .A(n2991), .ZN(n2997) );
  NAND2_X1 U3570 ( .A1(n3786), .A2(n3525), .ZN(n5736) );
  INV_X2 U3571 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3078) );
  NOR2_X2 U3572 ( .A1(n3726), .A2(n3224), .ZN(n3263) );
  INV_X2 U3573 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3079) );
  NAND2_X1 U3574 ( .A1(n3223), .A2(n3222), .ZN(n3726) );
  NAND2_X1 U3575 ( .A1(n3238), .A2(n3014), .ZN(n2998) );
  AND2_X2 U3576 ( .A1(n3258), .A2(n3227), .ZN(n3535) );
  INV_X1 U3577 ( .A(n3230), .ZN(n2999) );
  INV_X1 U3578 ( .A(n3230), .ZN(n3000) );
  OAI21_X2 U3579 ( .B1(n3235), .B2(n3805), .A(n4431), .ZN(n3228) );
  NAND2_X2 U3580 ( .A1(n3343), .A2(n3342), .ZN(n3352) );
  NOR2_X4 U3581 ( .A1(n5532), .A2(n5608), .ZN(n5606) );
  AND2_X1 U3582 ( .A1(n4473), .A2(n4248), .ZN(n3001) );
  AND2_X2 U3583 ( .A1(n4473), .A2(n4248), .ZN(n3002) );
  NAND2_X1 U3584 ( .A1(n3616), .A2(n3230), .ZN(n3707) );
  AND2_X2 U3585 ( .A1(n3230), .A2(n3014), .ZN(n4233) );
  OAI211_X2 U3586 ( .C1(n3229), .C2(n4431), .A(n3262), .B(n3228), .ZN(n3255)
         );
  AND2_X2 U3587 ( .A1(n3079), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3088)
         );
  OR2_X2 U3588 ( .A1(n5677), .A2(n5707), .ZN(n3765) );
  NAND2_X2 U3589 ( .A1(n3221), .A2(n3224), .ZN(n3241) );
  AND2_X4 U3590 ( .A1(n4476), .A2(n4473), .ZN(n3003) );
  BUF_X2 U3591 ( .A(n3281), .Z(n3007) );
  BUF_X4 U3592 ( .A(n3281), .Z(n3008) );
  AND2_X1 U3593 ( .A1(n3094), .A2(n3048), .ZN(n3009) );
  AND2_X2 U3594 ( .A1(n4461), .A2(n4248), .ZN(n3180) );
  AND2_X2 U3595 ( .A1(n3077), .A2(n3079), .ZN(n4461) );
  AND2_X2 U3596 ( .A1(n3094), .A2(n3088), .ZN(n5342) );
  NAND2_X2 U3597 ( .A1(n3237), .A2(n3236), .ZN(n3605) );
  NAND2_X2 U3598 ( .A1(n3353), .A2(n3426), .ZN(n3420) );
  NOR2_X2 U3599 ( .A1(n4446), .A2(n4447), .ZN(n4445) );
  NAND2_X1 U3600 ( .A1(n3765), .A2(n3530), .ZN(n5676) );
  OR2_X1 U3601 ( .A1(n4174), .A2(n4173), .ZN(n5658) );
  INV_X2 U3602 ( .A(n3523), .ZN(n5386) );
  NOR2_X4 U3603 ( .A1(n5393), .A2(n3992), .ZN(n5395) );
  NAND2_X2 U3604 ( .A1(n5177), .A2(n5178), .ZN(n6247) );
  NOR2_X2 U3605 ( .A1(n4452), .A2(n4605), .ZN(n4604) );
  NAND2_X1 U3606 ( .A1(n3310), .A2(n3311), .ZN(n3296) );
  BUF_X4 U3607 ( .A(n4441), .Z(n3014) );
  OAI21_X2 U3608 ( .B1(n5218), .B2(n3520), .A(n3519), .ZN(n5744) );
  NOR2_X2 U3609 ( .A1(n5542), .A2(n5543), .ZN(n5531) );
  NOR2_X2 U3610 ( .A1(n5124), .A2(n3044), .ZN(n4196) );
  NOR2_X2 U3611 ( .A1(n5128), .A2(n5185), .ZN(n5183) );
  NAND2_X2 U3612 ( .A1(n5635), .A2(n5634), .ZN(n5393) );
  AND2_X1 U3613 ( .A1(n3088), .A2(n4248), .ZN(n3015) );
  CLKBUF_X1 U3614 ( .A(n3015), .Z(n3016) );
  CLKBUF_X1 U3615 ( .A(n5341), .Z(n3017) );
  AND2_X1 U3616 ( .A1(n3088), .A2(n4248), .ZN(n5341) );
  AND2_X1 U3617 ( .A1(n6507), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3603) );
  OAI21_X1 U3618 ( .B1(n3578), .B2(n3390), .A(n3389), .ZN(n3464) );
  NAND2_X1 U3619 ( .A1(n3238), .A2(n3014), .ZN(n3628) );
  NAND2_X1 U3620 ( .A1(n5531), .A2(n5533), .ZN(n5532) );
  NAND2_X1 U3621 ( .A1(n4233), .A2(n3770), .ZN(n3712) );
  AND4_X2 U3622 ( .A1(n3163), .A2(n3162), .A3(n3161), .A4(n3160), .ZN(n3224)
         );
  NAND2_X1 U3623 ( .A1(n4337), .A2(n6499), .ZN(n3376) );
  INV_X1 U3624 ( .A(n5489), .ZN(n5434) );
  NOR2_X1 U3625 ( .A1(n3238), .A2(n4431), .ZN(n4234) );
  OR2_X1 U3626 ( .A1(n5486), .A2(n5487), .ZN(n5489) );
  NAND2_X1 U3627 ( .A1(n3608), .A2(n3607), .ZN(n3736) );
  AND2_X1 U3628 ( .A1(n3603), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4301) );
  AND2_X1 U3629 ( .A1(n3238), .A2(n3222), .ZN(n3206) );
  AND3_X1 U3630 ( .A1(n3351), .A2(n3350), .A3(n3349), .ZN(n3432) );
  NAND2_X1 U3631 ( .A1(n3226), .A2(n3238), .ZN(n3262) );
  AOI22_X1 U3632 ( .A1(n3329), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n5341), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3169) );
  AOI22_X1 U3633 ( .A1(n3324), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3167) );
  AOI22_X1 U3634 ( .A1(n3009), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3213), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3165) );
  XNOR2_X1 U3635 ( .A(n3496), .B(n3495), .ZN(n3795) );
  NAND2_X1 U3636 ( .A1(n3377), .A2(n4334), .ZN(n3465) );
  INV_X1 U3637 ( .A(n3726), .ZN(n3805) );
  INV_X1 U3638 ( .A(n5723), .ZN(n3790) );
  AND2_X1 U3639 ( .A1(n3732), .A2(n4312), .ZN(n5196) );
  AND2_X1 U3640 ( .A1(n5224), .A2(n4284), .ZN(n5200) );
  OAI21_X1 U3641 ( .B1(n3271), .B2(n3078), .A(n3254), .ZN(n3310) );
  INV_X1 U3642 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4838) );
  INV_X1 U3643 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6364) );
  INV_X1 U3644 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6471) );
  XNOR2_X1 U3645 ( .A(n4478), .B(n4614), .ZN(n4337) );
  INV_X1 U3646 ( .A(n6609), .ZN(n4194) );
  OR2_X1 U3647 ( .A1(n6609), .A2(n4187), .ZN(n6159) );
  OR2_X1 U3648 ( .A1(n5337), .A2(n5335), .ZN(n5368) );
  NAND2_X1 U3649 ( .A1(n5240), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5337)
         );
  NAND2_X1 U3650 ( .A1(n5606), .A2(n4103), .ZN(n5239) );
  OR2_X1 U3651 ( .A1(n3932), .A2(n3931), .ZN(n3933) );
  NAND2_X1 U3652 ( .A1(n3046), .A2(n3933), .ZN(n5234) );
  AND2_X1 U3653 ( .A1(n3946), .A2(n3945), .ZN(n3046) );
  INV_X1 U3654 ( .A(n5231), .ZN(n3945) );
  NAND2_X1 U3655 ( .A1(n3045), .A2(n4198), .ZN(n3044) );
  INV_X1 U3656 ( .A(n5123), .ZN(n3045) );
  AND2_X1 U3657 ( .A1(n3859), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3864)
         );
  NOR2_X1 U3658 ( .A1(n3844), .A2(n6137), .ZN(n3859) );
  AND2_X1 U3659 ( .A1(n5596), .A2(n5515), .ZN(n5517) );
  NOR2_X1 U3660 ( .A1(n5535), .A2(n3686), .ZN(n5611) );
  NAND2_X1 U3661 ( .A1(n5620), .A2(n5549), .ZN(n5535) );
  AND2_X1 U3662 ( .A1(n3677), .A2(n3676), .ZN(n5559) );
  OR2_X1 U3663 ( .A1(n5225), .A2(n3670), .ZN(n5627) );
  NOR2_X1 U3664 ( .A1(n5194), .A2(n3055), .ZN(n3054) );
  INV_X1 U3665 ( .A(n3515), .ZN(n3055) );
  NAND2_X1 U3666 ( .A1(n3516), .A2(n3515), .ZN(n3053) );
  AOI21_X1 U3667 ( .B1(n3511), .B2(n3065), .A(n3022), .ZN(n3064) );
  INV_X1 U3668 ( .A(n3510), .ZN(n3065) );
  AND2_X1 U3669 ( .A1(n5200), .A2(n4285), .ZN(n6296) );
  NAND2_X1 U3670 ( .A1(n3459), .A2(n3458), .ZN(n3460) );
  INV_X1 U3671 ( .A(n3039), .ZN(n4328) );
  OAI21_X1 U3672 ( .B1(n6196), .B2(n4298), .A(n3040), .ZN(n3039) );
  NAND2_X1 U3673 ( .A1(n3707), .A2(n3770), .ZN(n4229) );
  INV_X1 U3674 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4256) );
  NOR2_X1 U3675 ( .A1(n3820), .A2(n4837), .ZN(n4884) );
  NAND2_X1 U3676 ( .A1(n4574), .A2(n3820), .ZN(n4809) );
  AND2_X1 U3677 ( .A1(n4836), .A2(n4612), .ZN(n4705) );
  INV_X1 U3678 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6478) );
  AND2_X1 U3679 ( .A1(n3593), .A2(n3592), .ZN(n4262) );
  INV_X1 U3680 ( .A(n3591), .ZN(n3592) );
  INV_X2 U3681 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6498) );
  OR2_X1 U3682 ( .A1(n4221), .A2(n6505), .ZN(n4212) );
  NAND2_X1 U3683 ( .A1(n4291), .A2(n4212), .ZN(n6609) );
  INV_X1 U3684 ( .A(n6193), .ZN(n6176) );
  INV_X1 U3685 ( .A(n6122), .ZN(n6197) );
  OAI211_X1 U3686 ( .C1(n3033), .C2(n3032), .A(n3031), .B(n3030), .ZN(n5583)
         );
  NAND2_X1 U3687 ( .A1(n5434), .A2(n3024), .ZN(n3030) );
  NAND2_X1 U3688 ( .A1(n3033), .A2(n3029), .ZN(n3031) );
  NAND2_X1 U3689 ( .A1(n4353), .A2(n4304), .ZN(n5640) );
  AOI21_X1 U3690 ( .B1(n3531), .B2(n5676), .A(n3768), .ZN(n3533) );
  OR2_X1 U3691 ( .A1(n5790), .A2(n5769), .ZN(n5776) );
  AND2_X1 U3692 ( .A1(n3736), .A2(n3719), .ZN(n6353) );
  INV_X1 U3693 ( .A(n6167), .ZN(n6368) );
  NAND2_X1 U3694 ( .A1(n6471), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3546) );
  NAND2_X1 U3695 ( .A1(n3013), .A2(n3595), .ZN(n3240) );
  AND2_X2 U3696 ( .A1(n3234), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3094)
         );
  AND2_X1 U3697 ( .A1(n3230), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3562) );
  AND2_X1 U3698 ( .A1(n3553), .A2(n3554), .ZN(n3551) );
  OR2_X1 U3699 ( .A1(n3559), .A2(n3560), .ZN(n3543) );
  INV_X1 U3700 ( .A(n3364), .ZN(n3336) );
  OR2_X1 U3701 ( .A1(n3414), .A2(n3413), .ZN(n3498) );
  OR2_X1 U3702 ( .A1(n3289), .A2(n3288), .ZN(n3292) );
  OR2_X1 U3703 ( .A1(n3241), .A2(n2998), .ZN(n3201) );
  OR2_X1 U3704 ( .A1(n3374), .A2(n3373), .ZN(n3466) );
  OR2_X1 U3705 ( .A1(n3230), .A2(n6499), .ZN(n3363) );
  INV_X1 U3706 ( .A(n3578), .ZN(n3586) );
  INV_X1 U3707 ( .A(n3557), .ZN(n3596) );
  AND2_X1 U3708 ( .A1(n5319), .A2(n5483), .ZN(n5429) );
  NOR2_X1 U3709 ( .A1(n4024), .A2(n5563), .ZN(n4025) );
  NAND2_X1 U3710 ( .A1(n4196), .A2(n5129), .ZN(n5128) );
  INV_X1 U3711 ( .A(n3821), .ZN(n3833) );
  NAND2_X1 U3712 ( .A1(n5386), .A2(n3067), .ZN(n3786) );
  NOR2_X1 U3713 ( .A1(n3068), .A2(n3019), .ZN(n3067) );
  INV_X1 U3714 ( .A(n5387), .ZN(n3068) );
  INV_X1 U3715 ( .A(n3707), .ZN(n3699) );
  OAI21_X1 U3716 ( .B1(n3052), .B2(n3054), .A(n6008), .ZN(n3051) );
  NAND2_X1 U3717 ( .A1(n3648), .A2(n3034), .ZN(n3036) );
  NOR2_X1 U3718 ( .A1(n3656), .A2(n4195), .ZN(n3034) );
  NOR2_X1 U3719 ( .A1(n3066), .A2(n3063), .ZN(n3062) );
  INV_X1 U3720 ( .A(n5149), .ZN(n3063) );
  INV_X1 U3721 ( .A(n3511), .ZN(n3066) );
  AND2_X1 U3722 ( .A1(n3641), .A2(n3640), .ZN(n4607) );
  INV_X1 U3723 ( .A(n3292), .ZN(n3427) );
  OR2_X1 U3724 ( .A1(n3249), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3250)
         );
  INV_X1 U3725 ( .A(n3241), .ZN(n3612) );
  AND3_X1 U3726 ( .A1(n3239), .A2(n3227), .A3(n3238), .ZN(n3237) );
  INV_X1 U3727 ( .A(n4151), .ZN(n3360) );
  AND2_X1 U3728 ( .A1(n3246), .A2(n3274), .ZN(n4715) );
  OAI21_X1 U3729 ( .B1(n6613), .B2(n4779), .A(n6594), .ZN(n4343) );
  NAND2_X1 U3730 ( .A1(n3364), .A2(n3363), .ZN(n3590) );
  INV_X1 U3731 ( .A(n5029), .ZN(n4222) );
  AOI21_X1 U3732 ( .B1(n5434), .B2(n3027), .A(n3778), .ZN(n3029) );
  NOR2_X1 U3733 ( .A1(n3028), .A2(n3775), .ZN(n3027) );
  AND2_X1 U3734 ( .A1(n3774), .A2(n3773), .ZN(n3033) );
  NOR2_X1 U3735 ( .A1(n3028), .A2(n3025), .ZN(n3024) );
  NAND2_X1 U3736 ( .A1(n3778), .A2(n3026), .ZN(n3025) );
  INV_X1 U3737 ( .A(n3775), .ZN(n3026) );
  AND2_X1 U3738 ( .A1(n4778), .A2(n4777), .ZN(n6221) );
  AND2_X1 U3739 ( .A1(n5429), .A2(n5431), .ZN(n5411) );
  AND2_X1 U3740 ( .A1(n4201), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5240)
         );
  AND2_X1 U3741 ( .A1(n5314), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5297)
         );
  NOR2_X1 U3742 ( .A1(n5238), .A2(n5717), .ZN(n3047) );
  OR2_X1 U3743 ( .A1(n3076), .A2(n5237), .ZN(n5238) );
  AND2_X1 U3744 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n4099), .ZN(n4100)
         );
  INV_X1 U3745 ( .A(n4098), .ZN(n4099) );
  NAND2_X1 U3746 ( .A1(n4100), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4145)
         );
  AND2_X1 U3747 ( .A1(n4062), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4063)
         );
  AND2_X1 U3748 ( .A1(PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n4025), .ZN(n4062)
         );
  INV_X1 U3749 ( .A(n5623), .ZN(n4032) );
  NAND2_X1 U3750 ( .A1(n3993), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4024)
         );
  NOR2_X1 U3751 ( .A1(n3976), .A2(n5573), .ZN(n3993) );
  AND2_X1 U3752 ( .A1(n3927), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3928)
         );
  NAND2_X1 U3753 ( .A1(n3928), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3947)
         );
  NOR2_X1 U3754 ( .A1(n3908), .A2(n3907), .ZN(n3927) );
  NAND2_X1 U3755 ( .A1(n3891), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3908)
         );
  INV_X1 U3756 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3907) );
  NOR2_X1 U3757 ( .A1(n3878), .A2(n4188), .ZN(n3891) );
  CLKBUF_X1 U3758 ( .A(n5128), .Z(n5184) );
  NAND2_X1 U3759 ( .A1(n3864), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3878)
         );
  AND4_X1 U3760 ( .A1(n3863), .A2(n3862), .A3(n3861), .A4(n3860), .ZN(n5123)
         );
  AOI21_X1 U3761 ( .B1(n3795), .B2(n3985), .A(n3799), .ZN(n5014) );
  AOI21_X1 U3762 ( .B1(n3843), .B2(n3985), .A(n3847), .ZN(n4605) );
  NAND2_X1 U3763 ( .A1(n3842), .A2(n3841), .ZN(n4453) );
  AOI21_X1 U3764 ( .B1(n3829), .B2(n3985), .A(n3837), .ZN(n4447) );
  CLKBUF_X1 U3765 ( .A(n4445), .Z(n4454) );
  INV_X1 U3766 ( .A(n3814), .ZN(n3822) );
  NAND2_X1 U3767 ( .A1(n3822), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3821)
         );
  NAND2_X1 U3768 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3814) );
  NOR2_X1 U3769 ( .A1(n5697), .A2(n3071), .ZN(n3070) );
  INV_X1 U3770 ( .A(n3530), .ZN(n3071) );
  OR2_X1 U3771 ( .A1(n6339), .A2(n3747), .ZN(n5827) );
  OR2_X1 U3772 ( .A1(n5406), .A2(n3760), .ZN(n5790) );
  AOI21_X1 U3773 ( .B1(n4160), .B2(n3060), .A(n3018), .ZN(n3058) );
  NOR2_X1 U3774 ( .A1(n5729), .A2(n5840), .ZN(n3060) );
  NOR2_X1 U3775 ( .A1(n5729), .A2(n6249), .ZN(n3059) );
  AND2_X1 U3776 ( .A1(n3683), .A2(n5545), .ZN(n5548) );
  AND3_X1 U3777 ( .A1(n3741), .A2(n5196), .A3(n3740), .ZN(n5863) );
  NAND2_X1 U3778 ( .A1(n3038), .A2(n5559), .ZN(n3037) );
  INV_X1 U3779 ( .A(n5628), .ZN(n3038) );
  NOR2_X1 U3780 ( .A1(n5627), .A2(n5628), .ZN(n5626) );
  AND2_X1 U3781 ( .A1(n3662), .A2(n3661), .ZN(n6029) );
  NOR2_X2 U3782 ( .A1(n3036), .A2(n3035), .ZN(n6030) );
  INV_X1 U3783 ( .A(n5204), .ZN(n3035) );
  NAND2_X1 U3784 ( .A1(n3648), .A2(n3647), .ZN(n5131) );
  NAND2_X1 U3785 ( .A1(n5147), .A2(n5149), .ZN(n5148) );
  NAND2_X1 U3786 ( .A1(n5134), .A2(n5133), .ZN(n5136) );
  NAND2_X1 U3787 ( .A1(n3636), .A2(n3041), .ZN(n5015) );
  AND2_X1 U3788 ( .A1(n3042), .A2(n3635), .ZN(n3041) );
  INV_X1 U3789 ( .A(n4607), .ZN(n3042) );
  NAND2_X1 U3790 ( .A1(n3636), .A2(n3635), .ZN(n4608) );
  NAND2_X1 U3791 ( .A1(n4328), .A2(n4327), .ZN(n4326) );
  INV_X2 U3792 ( .A(n4233), .ZN(n4298) );
  NAND2_X1 U3793 ( .A1(n4332), .A2(n3445), .ZN(n3069) );
  AND2_X1 U3794 ( .A1(n3624), .A2(n3623), .ZN(n4230) );
  XNOR2_X1 U3795 ( .A(n3312), .B(n3311), .ZN(n3807) );
  CLKBUF_X1 U3796 ( .A(n3609), .Z(n3610) );
  NAND2_X1 U3797 ( .A1(n3356), .A2(n3355), .ZN(n4478) );
  AND2_X1 U3798 ( .A1(n6368), .A2(n4666), .ZN(n5888) );
  AND2_X1 U3799 ( .A1(n4666), .A2(n6167), .ZN(n5079) );
  INV_X1 U3800 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6137) );
  NAND2_X1 U3801 ( .A1(n6159), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6138) );
  INV_X1 U3802 ( .A(n6138), .ZN(n6184) );
  NOR2_X2 U3803 ( .A1(n4194), .A2(n4183), .ZN(n6193) );
  INV_X1 U3804 ( .A(n6182), .ZN(n6140) );
  NOR2_X2 U3805 ( .A1(n4194), .A2(n4193), .ZN(n6122) );
  AND2_X1 U3806 ( .A1(n5030), .A2(n6129), .ZN(n6188) );
  NAND2_X1 U3807 ( .A1(n5434), .A2(n5433), .ZN(n5432) );
  INV_X1 U3808 ( .A(n5637), .ZN(n6203) );
  INV_X1 U3809 ( .A(n6207), .ZN(n5617) );
  AND2_X2 U3810 ( .A1(n4237), .A2(n4301), .ZN(n6207) );
  NAND2_X1 U3811 ( .A1(n6207), .A2(n5641), .ZN(n5637) );
  INV_X1 U3812 ( .A(n5983), .ZN(n6215) );
  AND2_X1 U3813 ( .A1(n5640), .A2(n5453), .ZN(n6214) );
  INV_X1 U3814 ( .A(n5640), .ZN(n6217) );
  AND2_X1 U3815 ( .A1(n5640), .A2(n4306), .ZN(n5663) );
  INV_X2 U3817 ( .A(n4352), .ZN(n4418) );
  OR2_X1 U3818 ( .A1(n4291), .A2(n4290), .ZN(n4353) );
  XNOR2_X1 U3819 ( .A(n4204), .B(n4203), .ZN(n5418) );
  AOI21_X1 U3820 ( .B1(n5717), .B2(n5716), .A(n5715), .ZN(n5990) );
  NAND2_X1 U3821 ( .A1(n3933), .A2(n3946), .ZN(n5232) );
  INV_X1 U3822 ( .A(n6281), .ZN(n6253) );
  CLKBUF_X1 U3823 ( .A(n5067), .Z(n5068) );
  CLKBUF_X1 U3824 ( .A(n5055), .Z(n5056) );
  AND2_X1 U3825 ( .A1(n5489), .A2(n5488), .ZN(n5773) );
  NOR2_X1 U3826 ( .A1(n5847), .A2(n3759), .ZN(n5824) );
  INV_X1 U3827 ( .A(n3049), .ZN(n6007) );
  AOI21_X1 U3828 ( .B1(n6247), .B2(n3054), .A(n3052), .ZN(n3049) );
  INV_X1 U3829 ( .A(n6283), .ZN(n6355) );
  INV_X1 U3830 ( .A(n6353), .ZN(n6342) );
  AND2_X1 U3831 ( .A1(n3736), .A2(n4216), .ZN(n6339) );
  CLKBUF_X1 U3832 ( .A(n4338), .Z(n4339) );
  CLKBUF_X1 U3833 ( .A(n4243), .Z(n6170) );
  NOR2_X1 U3834 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n6593) );
  OAI21_X1 U3835 ( .B1(n4842), .B2(n4841), .A(n4840), .ZN(n4867) );
  INV_X1 U3836 ( .A(n6455), .ZN(n4603) );
  OR2_X1 U3837 ( .A1(n4618), .A2(n4617), .ZN(n4645) );
  AND3_X1 U3838 ( .A1(n4757), .A2(n4879), .A3(n4756), .ZN(n4802) );
  INV_X1 U3839 ( .A(n6384), .ZN(n5894) );
  INV_X1 U3840 ( .A(n6390), .ZN(n5901) );
  INV_X1 U3841 ( .A(n6433), .ZN(n5908) );
  INV_X1 U3842 ( .A(n6443), .ZN(n5913) );
  INV_X1 U3843 ( .A(n6404), .ZN(n5918) );
  INV_X1 U3844 ( .A(n6410), .ZN(n5925) );
  AND2_X1 U3845 ( .A1(n4342), .A2(n4341), .ZN(n4556) );
  CLKBUF_X1 U3846 ( .A(n4335), .Z(n4743) );
  INV_X1 U3847 ( .A(n4301), .ZN(n6505) );
  INV_X1 U3848 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6592) );
  AND3_X1 U3849 ( .A1(n3784), .A2(n3783), .A3(n3782), .ZN(n3785) );
  AND2_X1 U3850 ( .A1(n3763), .A2(n3762), .ZN(n3764) );
  NAND2_X1 U3851 ( .A1(n5395), .A2(n5558), .ZN(n5557) );
  NAND2_X1 U3852 ( .A1(n3058), .A2(n3057), .ZN(n5721) );
  NAND2_X1 U3853 ( .A1(n5395), .A2(n3023), .ZN(n5542) );
  AND2_X1 U3854 ( .A1(n3789), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3018)
         );
  AND2_X1 U3855 ( .A1(n5386), .A2(n5387), .ZN(n5385) );
  INV_X1 U3856 ( .A(n4431), .ZN(n3227) );
  AOI22_X1 U3857 ( .A1(n3788), .A2(n3789), .B1(n4160), .B2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5728) );
  AND2_X1 U3858 ( .A1(n6249), .A2(n3742), .ZN(n3019) );
  AND3_X1 U3859 ( .A1(n3146), .A2(n3145), .A3(n3144), .ZN(n3020) );
  NAND2_X1 U3860 ( .A1(n3424), .A2(n3423), .ZN(n3462) );
  XNOR2_X1 U3861 ( .A(n3474), .B(n3473), .ZN(n3838) );
  AND2_X1 U3862 ( .A1(n4334), .A2(n3464), .ZN(n3021) );
  AND2_X1 U3863 ( .A1(n3789), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n3022)
         );
  INV_X1 U3864 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3234) );
  NOR2_X1 U3865 ( .A1(n5124), .A2(n5123), .ZN(n4197) );
  OAI21_X1 U3866 ( .B1(n6247), .B2(n3516), .A(n3515), .ZN(n5191) );
  NAND2_X1 U3867 ( .A1(n5148), .A2(n3510), .ZN(n5139) );
  NAND2_X1 U3868 ( .A1(n6030), .A2(n6029), .ZN(n5225) );
  INV_X1 U3869 ( .A(n4195), .ZN(n3647) );
  INV_X1 U3870 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6499) );
  AND2_X1 U3871 ( .A1(n4775), .A2(n3794), .ZN(n6276) );
  NOR2_X1 U3872 ( .A1(n4326), .A2(n4318), .ZN(n4317) );
  AND2_X1 U3873 ( .A1(n4032), .A2(n5558), .ZN(n3023) );
  OAI21_X1 U3874 ( .B1(n3255), .B2(n3256), .A(n3257), .ZN(n3720) );
  INV_X1 U3875 ( .A(n5717), .ZN(n4103) );
  INV_X1 U3876 ( .A(n5433), .ZN(n3028) );
  INV_X1 U3877 ( .A(n3778), .ZN(n3032) );
  AND2_X4 U3878 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4248) );
  INV_X1 U3879 ( .A(n3036), .ZN(n6115) );
  NOR2_X2 U3880 ( .A1(n5627), .A2(n3037), .ZN(n5620) );
  NAND2_X1 U3881 ( .A1(n2999), .A2(n3014), .ZN(n4225) );
  INV_X1 U3882 ( .A(n3698), .ZN(n5597) );
  NAND2_X1 U3883 ( .A1(n5517), .A2(n5501), .ZN(n5486) );
  INV_X1 U3884 ( .A(n5598), .ZN(n3043) );
  INV_X1 U3885 ( .A(n3474), .ZN(n3404) );
  NOR2_X4 U3886 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4476) );
  AND2_X2 U3887 ( .A1(n5606), .A2(n3047), .ZN(n5593) );
  AND2_X2 U3888 ( .A1(n3093), .A2(n3048), .ZN(n3324) );
  AND2_X4 U3889 ( .A1(n4476), .A2(n3048), .ZN(n3329) );
  NAND2_X1 U3890 ( .A1(n3056), .A2(n3518), .ZN(n5218) );
  NAND3_X1 U3891 ( .A1(n3058), .A2(n3057), .A3(n3790), .ZN(n3791) );
  NAND2_X1 U3892 ( .A1(n3788), .A2(n3059), .ZN(n3057) );
  NAND2_X1 U3893 ( .A1(n5147), .A2(n3062), .ZN(n3061) );
  INV_X1 U3894 ( .A(n5736), .ZN(n3787) );
  NAND2_X1 U3895 ( .A1(n3069), .A2(n3439), .ZN(n4308) );
  XNOR2_X1 U3896 ( .A(n3431), .B(n3433), .ZN(n4332) );
  AND2_X2 U3897 ( .A1(n3765), .A2(n3070), .ZN(n5690) );
  CLKBUF_X1 U3898 ( .A(n4332), .Z(n4835) );
  NAND2_X1 U3899 ( .A1(n3470), .A2(n3469), .ZN(n3471) );
  XNOR2_X1 U3900 ( .A(n3297), .B(n3296), .ZN(n4338) );
  AOI21_X2 U3901 ( .B1(n3807), .B2(n6499), .A(n3341), .ZN(n3444) );
  NAND2_X1 U3902 ( .A1(n3223), .A2(n3221), .ZN(n3226) );
  OR2_X2 U3903 ( .A1(n3200), .A2(n3199), .ZN(n3238) );
  CLKBUF_X1 U3904 ( .A(n4331), .Z(n4836) );
  XNOR2_X1 U3905 ( .A(n3426), .B(n3425), .ZN(n4331) );
  AOI21_X1 U3906 ( .B1(n4308), .B2(n4307), .A(n3456), .ZN(n4562) );
  OR2_X1 U3907 ( .A1(n3789), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3072)
         );
  AND2_X1 U3908 ( .A1(n6249), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3073)
         );
  AND4_X1 U3909 ( .A1(n3179), .A2(n3178), .A3(n3177), .A4(n3176), .ZN(n3074)
         );
  INV_X1 U3910 ( .A(n3809), .ZN(n4006) );
  INV_X1 U3911 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5840) );
  INV_X1 U3912 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6040) );
  INV_X1 U3913 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4188) );
  BUF_X1 U3914 ( .A(n3329), .Z(n3382) );
  AND2_X1 U3915 ( .A1(n5371), .A2(n5370), .ZN(n3075) );
  AND2_X1 U3916 ( .A1(n4150), .A2(n4149), .ZN(n3076) );
  INV_X1 U3917 ( .A(n5606), .ZN(n5716) );
  OR2_X1 U3918 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n5362) );
  NAND2_X1 U3919 ( .A1(n5055), .A2(n5057), .ZN(n5058) );
  AND2_X1 U3920 ( .A1(n3143), .A2(n4225), .ZN(n3188) );
  OR2_X1 U3921 ( .A1(n3388), .A2(n3387), .ZN(n3485) );
  NAND2_X1 U3922 ( .A1(n3796), .A2(n3239), .ZN(n3204) );
  AOI22_X1 U3923 ( .A1(n3213), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3190), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3178) );
  BUF_X1 U3924 ( .A(n3004), .Z(n5350) );
  OR2_X1 U3925 ( .A1(n3401), .A2(n3400), .ZN(n3484) );
  OAI21_X1 U3926 ( .B1(n3578), .B2(n3403), .A(n3402), .ZN(n3473) );
  OAI21_X1 U3927 ( .B1(n3578), .B2(n3416), .A(n3415), .ZN(n3482) );
  OR2_X1 U3928 ( .A1(n3556), .A2(n3555), .ZN(n3557) );
  AND2_X1 U3929 ( .A1(n6249), .A2(n5219), .ZN(n3520) );
  XNOR2_X1 U3930 ( .A(n3483), .B(n3482), .ZN(n3843) );
  INV_X1 U3931 ( .A(n3603), .ZN(n3359) );
  NAND2_X1 U3932 ( .A1(n3336), .A2(n3505), .ZN(n3418) );
  INV_X1 U3933 ( .A(n3712), .ZN(n3674) );
  AOI21_X1 U3934 ( .B1(n3590), .B2(n3601), .A(n3589), .ZN(n3591) );
  NOR2_X1 U3935 ( .A1(n3578), .A2(n3548), .ZN(n3575) );
  AND2_X1 U3936 ( .A1(n4200), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5314)
         );
  OR2_X1 U3937 ( .A1(n6071), .A2(n5362), .ZN(n4030) );
  INV_X1 U3938 ( .A(n5014), .ZN(n3848) );
  XNOR2_X1 U3939 ( .A(n3465), .B(n3464), .ZN(n3829) );
  INV_X1 U3940 ( .A(n4457), .ZN(n3635) );
  AND2_X1 U3941 ( .A1(n3358), .A2(n4557), .ZN(n4615) );
  OR2_X1 U3942 ( .A1(n3322), .A2(n3321), .ZN(n3449) );
  AOI21_X1 U3943 ( .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n6478), .A(n3551), 
        .ZN(n3549) );
  NOR2_X1 U3944 ( .A1(n6176), .A2(n5437), .ZN(n6072) );
  OR2_X1 U3945 ( .A1(n6463), .A2(n6499), .ZN(n5366) );
  OR2_X1 U3946 ( .A1(n5394), .A2(n5571), .ZN(n3992) );
  OR2_X1 U3947 ( .A1(n5368), .A2(n4202), .ZN(n4204) );
  NAND2_X1 U3948 ( .A1(n5297), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5301)
         );
  NAND2_X1 U3949 ( .A1(n4063), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4098)
         );
  NAND2_X1 U3950 ( .A1(n3961), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3976)
         );
  INV_X1 U3951 ( .A(n4146), .ZN(n5413) );
  AND2_X1 U3952 ( .A1(n3535), .A2(n3536), .ZN(n3613) );
  AND2_X1 U3953 ( .A1(n4336), .A2(n4343), .ZN(n4539) );
  NOR2_X1 U3954 ( .A1(n4145), .A2(n5527), .ZN(n4200) );
  INV_X1 U3955 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5573) );
  AND2_X1 U3956 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n3833), .ZN(n3839)
         );
  INV_X1 U3957 ( .A(n5362), .ZN(n5369) );
  INV_X1 U3958 ( .A(n3947), .ZN(n3961) );
  NAND2_X1 U3959 ( .A1(n3839), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3844)
         );
  NAND2_X1 U3960 ( .A1(n5700), .A2(n3073), .ZN(n5681) );
  OR2_X1 U3961 ( .A1(n4508), .A2(n4835), .ZN(n4976) );
  OR2_X1 U3962 ( .A1(n4508), .A2(n4580), .ZN(n6438) );
  NAND2_X1 U3963 ( .A1(n4815), .A2(n3446), .ZN(n5084) );
  AND2_X1 U3964 ( .A1(n4623), .A2(n4622), .ZN(n4646) );
  AND2_X1 U3965 ( .A1(n4717), .A2(n4716), .ZN(n4740) );
  AOI21_X1 U3966 ( .B1(n6364), .B2(STATE2_REG_3__SCAN_IN), .A(n4616), .ZN(
        n4879) );
  NOR2_X1 U3967 ( .A1(n6592), .A2(n4262), .ZN(n6497) );
  INV_X1 U3968 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6507) );
  NOR2_X1 U3969 ( .A1(n3255), .A2(n3534), .ZN(n4220) );
  NOR2_X1 U3970 ( .A1(n5524), .A2(n6660), .ZN(n5944) );
  NOR2_X1 U3971 ( .A1(n5440), .A2(n6065), .ZN(n5971) );
  OR2_X1 U3972 ( .A1(n6084), .A2(n6183), .ZN(n6082) );
  INV_X1 U3973 ( .A(n6129), .ZN(n6146) );
  AND2_X1 U3974 ( .A1(n5418), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4206) );
  AND2_X1 U3976 ( .A1(n5640), .A2(n5455), .ZN(n6218) );
  NOR2_X1 U3977 ( .A1(n4262), .A2(n6505), .ZN(n4775) );
  INV_X1 U3978 ( .A(n4353), .ZN(n4410) );
  INV_X1 U3979 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3532) );
  NAND2_X1 U3980 ( .A1(n3791), .A2(n3072), .ZN(n5714) );
  AND2_X1 U3981 ( .A1(n6023), .A2(n3757), .ZN(n5868) );
  NOR2_X1 U3982 ( .A1(n6288), .A2(n6011), .ZN(n6023) );
  AND2_X1 U3983 ( .A1(n3454), .A2(n3455), .ZN(n4307) );
  NAND2_X1 U3984 ( .A1(n6499), .A2(n4343), .ZN(n4616) );
  INV_X1 U3985 ( .A(n6497), .ZN(n6594) );
  INV_X1 U3986 ( .A(n4843), .ZN(n4871) );
  OAI221_X1 U3987 ( .B1(n5885), .B2(n6592), .C1(n5885), .C2(n5884), .A(n5883), 
        .ZN(n5932) );
  OAI21_X1 U3988 ( .B1(n4677), .B2(n4676), .A(n4675), .ZN(n4701) );
  INV_X1 U3989 ( .A(n4699), .ZN(n4543) );
  OAI21_X1 U3990 ( .B1(n4974), .B2(n4512), .A(n4511), .ZN(n4538) );
  NOR2_X1 U3991 ( .A1(n4809), .A2(n4835), .ZN(n4815) );
  INV_X1 U3992 ( .A(n4920), .ZN(n4962) );
  INV_X1 U3993 ( .A(n5084), .ZN(n5109) );
  INV_X1 U3994 ( .A(n4800), .ZN(n4649) );
  AND2_X1 U3995 ( .A1(n4705), .A2(n3446), .ZN(n4706) );
  NAND2_X1 U3996 ( .A1(n4215), .A2(n4775), .ZN(n4291) );
  NAND2_X1 U3997 ( .A1(n6159), .A2(n4205), .ZN(n6129) );
  NAND2_X1 U3998 ( .A1(n6159), .A2(n4206), .ZN(n6187) );
  INV_X1 U3999 ( .A(n5686), .ZN(n5650) );
  INV_X1 U4000 ( .A(n5663), .ZN(n5039) );
  INV_X1 U4001 ( .A(n6221), .ZN(n6245) );
  INV_X1 U4002 ( .A(n4178), .ZN(n4179) );
  OR2_X1 U4003 ( .A1(n6517), .A2(n5875), .ZN(n6267) );
  OR2_X1 U4004 ( .A1(n6263), .A2(n4550), .ZN(n6281) );
  AND2_X1 U4005 ( .A1(n4169), .A2(n4168), .ZN(n4170) );
  NAND2_X1 U4006 ( .A1(n5868), .A2(n3758), .ZN(n5847) );
  NOR2_X1 U4007 ( .A1(n6028), .A2(n3756), .ZN(n6288) );
  INV_X1 U4008 ( .A(n6598), .ZN(n5384) );
  NAND2_X1 U4009 ( .A1(n4884), .A2(n4975), .ZN(n4913) );
  NAND2_X1 U4010 ( .A1(n4884), .A2(n3446), .ZN(n5943) );
  NAND2_X1 U4011 ( .A1(n4509), .A2(n4975), .ZN(n5007) );
  OR2_X1 U4012 ( .A1(n4508), .A2(n4671), .ZN(n6447) );
  AOI21_X1 U4013 ( .B1(n4926), .B2(n4929), .A(n4925), .ZN(n4965) );
  OR2_X1 U4014 ( .A1(n4809), .A2(n4671), .ZN(n6460) );
  INV_X1 U4015 ( .A(n6417), .ZN(n5933) );
  OR2_X1 U4016 ( .A1(n4809), .A2(n4580), .ZN(n6453) );
  INV_X1 U4017 ( .A(n4706), .ZN(n4808) );
  OR2_X1 U4018 ( .A1(n4345), .A2(n4975), .ZN(n4843) );
  INV_X1 U4019 ( .A(n6588), .ZN(n6518) );
  INV_X1 U4020 ( .A(n6576), .ZN(n6584) );
  INV_X1 U4021 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3077) );
  NAND2_X1 U4022 ( .A1(n2987), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3083)
         );
  AND2_X4 U4023 ( .A1(n3093), .A2(n4473), .ZN(n3190) );
  NAND2_X1 U4024 ( .A1(n3190), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3082)
         );
  NAND2_X1 U4025 ( .A1(n3323), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3081) );
  AND2_X2 U4026 ( .A1(n3088), .A2(n4476), .ZN(n3175) );
  NAND2_X1 U4027 ( .A1(n3175), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3080) );
  AND2_X2 U4028 ( .A1(n3093), .A2(n3088), .ZN(n3189) );
  NAND2_X1 U4029 ( .A1(n3189), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3087) );
  NAND2_X1 U4030 ( .A1(n3324), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3086)
         );
  NAND2_X1 U4031 ( .A1(n3207), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3085)
         );
  AND2_X4 U4032 ( .A1(n4476), .A2(n4473), .ZN(n5343) );
  NAND2_X1 U4033 ( .A1(n5343), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3084)
         );
  NAND2_X1 U4034 ( .A1(n3329), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3092) );
  NAND2_X1 U4035 ( .A1(n5342), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3091) );
  NAND2_X1 U4036 ( .A1(n3015), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3090) );
  AND2_X4 U4037 ( .A1(n4473), .A2(n4248), .ZN(n3212) );
  NAND2_X1 U4038 ( .A1(n3212), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3089)
         );
  AND2_X2 U4039 ( .A1(n3093), .A2(n4461), .ZN(n3281) );
  NAND2_X1 U4040 ( .A1(n3008), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3098) );
  AND2_X2 U4041 ( .A1(n3094), .A2(n4461), .ZN(n3283) );
  NAND2_X1 U4042 ( .A1(n3283), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3097) );
  AND2_X2 U4043 ( .A1(n4476), .A2(n4461), .ZN(n3282) );
  NAND2_X1 U4044 ( .A1(n3282), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3096) );
  NAND2_X1 U4045 ( .A1(n3180), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3095) );
  NAND2_X1 U4046 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_1__SCAN_IN), .ZN(
        n6534) );
  OAI21_X1 U4047 ( .B1(STATE_REG_2__SCAN_IN), .B2(STATE_REG_1__SCAN_IN), .A(
        n6534), .ZN(n3595) );
  NAND2_X1 U4048 ( .A1(n3189), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3106) );
  NAND2_X1 U4049 ( .A1(n3324), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3105)
         );
  NAND2_X1 U4050 ( .A1(n3207), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3104)
         );
  NAND2_X1 U4051 ( .A1(n5343), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3103)
         );
  NAND2_X1 U4052 ( .A1(n3213), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3110)
         );
  NAND2_X1 U4053 ( .A1(n3190), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3109)
         );
  NAND2_X1 U4054 ( .A1(n3009), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3108) );
  NAND2_X1 U4055 ( .A1(n3175), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3107) );
  NAND2_X1 U4056 ( .A1(n5342), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3114) );
  NAND2_X1 U4057 ( .A1(n3329), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3113) );
  NAND2_X1 U4058 ( .A1(n5341), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3112) );
  NAND2_X1 U4059 ( .A1(n3212), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3111)
         );
  NAND2_X1 U4060 ( .A1(n3008), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3118) );
  NAND2_X1 U4061 ( .A1(n3283), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3117) );
  NAND2_X1 U4062 ( .A1(n3282), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3116) );
  NAND2_X1 U4063 ( .A1(n3180), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3115) );
  NAND4_X4 U4064 ( .A1(n3122), .A2(n3121), .A3(n3120), .A4(n3119), .ZN(n3221)
         );
  NAND2_X1 U4065 ( .A1(n3240), .A2(n3239), .ZN(n3143) );
  NAND2_X1 U4066 ( .A1(n3009), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3126) );
  NAND2_X1 U4067 ( .A1(n3190), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3125)
         );
  NAND2_X1 U4068 ( .A1(n3189), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3124) );
  NAND2_X1 U4069 ( .A1(n3175), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3123) );
  NAND2_X1 U4070 ( .A1(n3207), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3130)
         );
  NAND2_X1 U4071 ( .A1(n3213), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3129)
         );
  NAND2_X1 U4072 ( .A1(n5341), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3128) );
  NAND2_X1 U4073 ( .A1(n3329), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3127) );
  NAND2_X1 U4074 ( .A1(n3007), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3134) );
  NAND2_X1 U4075 ( .A1(n5342), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3133) );
  NAND2_X1 U4076 ( .A1(n3283), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3132) );
  NAND2_X1 U4077 ( .A1(n3180), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3131) );
  NAND2_X1 U4078 ( .A1(n3324), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3138)
         );
  NAND2_X1 U4079 ( .A1(n5343), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3137)
         );
  NAND2_X1 U4080 ( .A1(n3282), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3136) );
  NAND2_X1 U4081 ( .A1(n3002), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3135)
         );
  NAND4_X4 U4082 ( .A1(n3142), .A2(n3141), .A3(n3140), .A4(n3139), .ZN(n3230)
         );
  NAND2_X1 U4083 ( .A1(n3175), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3147) );
  NAND2_X1 U4084 ( .A1(n3323), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3146) );
  NAND2_X1 U4085 ( .A1(n3190), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3145)
         );
  NAND2_X1 U4086 ( .A1(n2987), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3144)
         );
  NAND2_X1 U4087 ( .A1(n5342), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3151) );
  NAND2_X1 U4088 ( .A1(n3329), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3150) );
  NAND2_X1 U4089 ( .A1(n5341), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3149) );
  NAND2_X1 U4090 ( .A1(n3212), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3148)
         );
  NAND2_X1 U4091 ( .A1(n3008), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3155) );
  NAND2_X1 U4092 ( .A1(n3283), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3154) );
  NAND2_X1 U4093 ( .A1(n3282), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3153) );
  NAND2_X1 U4094 ( .A1(n3180), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3152) );
  NAND2_X1 U4095 ( .A1(n3189), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3159) );
  NAND2_X1 U4096 ( .A1(n3324), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3158)
         );
  NAND2_X1 U4097 ( .A1(n3207), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3157)
         );
  NAND2_X1 U4098 ( .A1(n5343), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3156)
         );
  AOI22_X1 U4099 ( .A1(n3282), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3166) );
  AOI22_X1 U4100 ( .A1(n3007), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3180), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3164) );
  AOI22_X1 U4101 ( .A1(n5342), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3283), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3170) );
  AOI22_X1 U4102 ( .A1(n3189), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n5343), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3168) );
  AOI22_X1 U4103 ( .A1(n3190), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3175), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3171) );
  NAND2_X1 U4104 ( .A1(n3223), .A2(n3224), .ZN(n3174) );
  AOI22_X1 U4105 ( .A1(n3189), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3179) );
  AOI22_X1 U4106 ( .A1(n3009), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3175), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3177) );
  AOI22_X1 U4107 ( .A1(n3324), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3003), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3176) );
  AOI22_X1 U4108 ( .A1(n5342), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3015), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3184) );
  AOI22_X1 U4109 ( .A1(n3007), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3183) );
  AOI22_X1 U4110 ( .A1(n3283), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3180), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3182) );
  AOI22_X1 U4111 ( .A1(n3329), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3002), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3181) );
  NAND2_X2 U4112 ( .A1(n3186), .A2(n3222), .ZN(n3235) );
  AND2_X1 U4113 ( .A1(n3226), .A2(n3230), .ZN(n3187) );
  NAND2_X1 U4114 ( .A1(n3235), .A2(n3187), .ZN(n3538) );
  NAND2_X1 U4115 ( .A1(n3235), .A2(n3261), .ZN(n3202) );
  AOI22_X1 U4116 ( .A1(n3189), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3194) );
  AOI22_X1 U4117 ( .A1(n3009), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3175), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3193) );
  AOI22_X1 U4118 ( .A1(n3190), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        INSTQUEUE_REG_11__3__SCAN_IN), .B2(n2987), .ZN(n3192) );
  AOI22_X1 U4119 ( .A1(n3324), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n5343), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3191) );
  NAND4_X1 U4120 ( .A1(n3194), .A2(n3193), .A3(n3192), .A4(n3191), .ZN(n3200)
         );
  AOI22_X1 U4121 ( .A1(n5342), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3015), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3198) );
  AOI22_X1 U4122 ( .A1(n3007), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3197) );
  AOI22_X1 U4123 ( .A1(n3283), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3180), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3196) );
  AOI22_X1 U4124 ( .A1(n3329), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3212), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3195) );
  NAND4_X1 U4125 ( .A1(n3198), .A2(n3197), .A3(n3196), .A4(n3195), .ZN(n3199)
         );
  INV_X1 U4126 ( .A(n3226), .ZN(n3203) );
  NAND2_X1 U4127 ( .A1(n3203), .A2(n4232), .ZN(n3205) );
  AOI22_X1 U4128 ( .A1(n3175), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3211) );
  AOI22_X1 U4129 ( .A1(n5342), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n5341), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3210) );
  AOI22_X1 U4130 ( .A1(n3007), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3283), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3209) );
  AOI22_X1 U4131 ( .A1(n3324), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n5343), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3208) );
  AOI22_X1 U4132 ( .A1(n3329), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3002), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3217) );
  AOI22_X1 U4133 ( .A1(n3323), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3216) );
  AOI22_X1 U4134 ( .A1(n2987), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3190), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3215) );
  AOI22_X1 U4135 ( .A1(n3282), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3180), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3214) );
  AND3_X2 U4136 ( .A1(n3220), .A2(n3267), .A3(n3535), .ZN(n3232) );
  INV_X1 U4137 ( .A(n3263), .ZN(n3225) );
  OAI21_X1 U4138 ( .B1(n3221), .B2(n5452), .A(n3225), .ZN(n3229) );
  NAND2_X1 U4139 ( .A1(n3255), .A2(n3000), .ZN(n3231) );
  NAND2_X1 U4140 ( .A1(n3232), .A2(n3231), .ZN(n3233) );
  NAND2_X1 U4141 ( .A1(n3233), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3271) );
  INV_X1 U4142 ( .A(n3235), .ZN(n3236) );
  NOR2_X2 U4143 ( .A1(n3605), .A2(n3000), .ZN(n4215) );
  AND2_X2 U4144 ( .A1(n3013), .A2(n2999), .ZN(n5029) );
  NAND3_X1 U4145 ( .A1(n3006), .A2(n5029), .A3(n3239), .ZN(n3724) );
  AOI21_X1 U4146 ( .B1(n4215), .B2(n3240), .A(n3611), .ZN(n3244) );
  INV_X1 U4147 ( .A(n3255), .ZN(n3243) );
  NOR2_X1 U4148 ( .A1(n4222), .A2(n3241), .ZN(n3242) );
  NAND2_X1 U4149 ( .A1(n3243), .A2(n3242), .ZN(n3609) );
  NAND2_X1 U4150 ( .A1(n3244), .A2(n3609), .ZN(n3245) );
  NAND2_X1 U4151 ( .A1(n3245), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3247) );
  NAND2_X1 U4152 ( .A1(n6593), .A2(n6499), .ZN(n4151) );
  NAND2_X1 U4153 ( .A1(n6364), .A2(n4838), .ZN(n3246) );
  NAND2_X1 U4154 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3274) );
  AOI22_X1 U4155 ( .A1(n3360), .A2(n4715), .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n3359), .ZN(n3248) );
  OAI211_X1 U4156 ( .C1(n3271), .C2(n3234), .A(n3247), .B(n3248), .ZN(n3269)
         );
  INV_X1 U4157 ( .A(n3247), .ZN(n3251) );
  INV_X1 U4158 ( .A(n3248), .ZN(n3249) );
  NAND2_X1 U4159 ( .A1(n3251), .A2(n3250), .ZN(n3252) );
  AND2_X2 U4160 ( .A1(n3269), .A2(n3252), .ZN(n3297) );
  MUX2_X1 U4161 ( .A(n3360), .B(n3359), .S(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), 
        .Z(n3253) );
  INV_X1 U4162 ( .A(n3253), .ZN(n3254) );
  AND2_X1 U4163 ( .A1(n3241), .A2(n3014), .ZN(n3256) );
  NAND2_X1 U4164 ( .A1(n3227), .A2(n3230), .ZN(n3257) );
  INV_X1 U4165 ( .A(n3258), .ZN(n3260) );
  AND2_X1 U4166 ( .A1(n2997), .A2(n4524), .ZN(n3259) );
  OAI21_X1 U4167 ( .B1(n3260), .B2(n3259), .A(n3014), .ZN(n3266) );
  NAND2_X1 U4168 ( .A1(n6593), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6506) );
  AOI21_X1 U4169 ( .B1(n3262), .B2(n2989), .A(n6506), .ZN(n3265) );
  NAND2_X1 U4170 ( .A1(n3263), .A2(n3006), .ZN(n3264) );
  AND4_X1 U4171 ( .A1(n3267), .A2(n3266), .A3(n3265), .A4(n3264), .ZN(n3268)
         );
  NAND2_X1 U4172 ( .A1(n3720), .A2(n3268), .ZN(n3311) );
  NAND2_X1 U4173 ( .A1(n3297), .A2(n3296), .ZN(n3270) );
  NAND2_X1 U4174 ( .A1(n3270), .A2(n3269), .ZN(n3354) );
  INV_X1 U4175 ( .A(n3274), .ZN(n3273) );
  NAND2_X1 U4176 ( .A1(n3273), .A2(n6471), .ZN(n4667) );
  NAND2_X1 U4177 ( .A1(n3274), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3275) );
  NAND2_X1 U4178 ( .A1(n4667), .A2(n3275), .ZN(n4514) );
  AOI22_X1 U4179 ( .A1(n3360), .A2(n4514), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3359), .ZN(n3276) );
  XNOR2_X1 U4180 ( .A(n3354), .B(n3355), .ZN(n4243) );
  NAND2_X1 U4181 ( .A1(n4243), .A2(n6499), .ZN(n3291) );
  AOI22_X1 U4182 ( .A1(n4108), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3005), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3280) );
  AOI22_X1 U4183 ( .A1(n5340), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n5348), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3279) );
  AOI22_X1 U4184 ( .A1(n4119), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3012), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3278) );
  AOI22_X1 U4185 ( .A1(n5349), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3003), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3277) );
  NAND4_X1 U4186 ( .A1(n3280), .A2(n3279), .A3(n3278), .A4(n3277), .ZN(n3289)
         );
  AOI22_X1 U4187 ( .A1(n3010), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3017), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3287) );
  AOI22_X1 U4188 ( .A1(n3391), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n5350), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3286) );
  AOI22_X1 U4189 ( .A1(n5258), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n5326), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3285) );
  AOI22_X1 U4190 ( .A1(n3382), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3002), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3284) );
  NAND4_X1 U4191 ( .A1(n3287), .A2(n3286), .A3(n3285), .A4(n3284), .ZN(n3288)
         );
  NAND2_X1 U4192 ( .A1(n3336), .A2(n3292), .ZN(n3290) );
  INV_X1 U4193 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3293) );
  OAI22_X1 U4194 ( .A1(n3578), .A2(n3293), .B1(n3427), .B2(n3363), .ZN(n3294)
         );
  XNOR2_X2 U4195 ( .A(n3295), .B(n3294), .ZN(n3425) );
  INV_X1 U4196 ( .A(n3425), .ZN(n3353) );
  AOI22_X1 U4197 ( .A1(n4108), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3005), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3301) );
  AOI22_X1 U4198 ( .A1(n5340), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5348), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3300) );
  AOI22_X1 U4199 ( .A1(n4119), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3012), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3299) );
  AOI22_X1 U4200 ( .A1(n3324), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n5343), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3298) );
  NAND4_X1 U4201 ( .A1(n3301), .A2(n3300), .A3(n3299), .A4(n3298), .ZN(n3307)
         );
  AOI22_X1 U4202 ( .A1(n3011), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3305) );
  AOI22_X1 U4203 ( .A1(n3391), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n5350), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3304) );
  AOI22_X1 U4204 ( .A1(n5258), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n5326), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3303) );
  AOI22_X1 U4205 ( .A1(n3382), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3212), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3302) );
  NAND4_X1 U4206 ( .A1(n3305), .A2(n3304), .A3(n3303), .A4(n3302), .ZN(n3306)
         );
  INV_X1 U4207 ( .A(n3435), .ZN(n3308) );
  NOR2_X1 U4208 ( .A1(n3308), .A2(n3364), .ZN(n3309) );
  AOI21_X2 U4209 ( .B1(n4338), .B2(n6499), .A(n3309), .ZN(n3344) );
  INV_X1 U4210 ( .A(n3344), .ZN(n3343) );
  INV_X1 U4211 ( .A(n3310), .ZN(n3312) );
  AOI22_X1 U4212 ( .A1(n5340), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3316) );
  AOI22_X1 U4213 ( .A1(n3324), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3012), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3315) );
  AOI22_X1 U4214 ( .A1(n3016), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3002), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3314) );
  AOI22_X1 U4215 ( .A1(n3391), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n5326), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3313) );
  NAND4_X1 U4216 ( .A1(n3316), .A2(n3315), .A3(n3314), .A4(n3313), .ZN(n3322)
         );
  AOI22_X1 U4217 ( .A1(n4108), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3005), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3320) );
  AOI22_X1 U4218 ( .A1(n3011), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3329), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3319) );
  AOI22_X1 U4219 ( .A1(n5348), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n5343), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3318) );
  AOI22_X1 U4220 ( .A1(n3283), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3004), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3317) );
  NAND4_X1 U4221 ( .A1(n3320), .A2(n3319), .A3(n3318), .A4(n3317), .ZN(n3321)
         );
  AOI22_X1 U4222 ( .A1(n4108), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3005), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3328) );
  AOI22_X1 U4223 ( .A1(n5340), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n5348), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3327) );
  AOI22_X1 U4224 ( .A1(n4119), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3326) );
  AOI22_X1 U4225 ( .A1(n3324), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n5343), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3325) );
  NAND4_X1 U4226 ( .A1(n3328), .A2(n3327), .A3(n3326), .A4(n3325), .ZN(n3335)
         );
  AOI22_X1 U4227 ( .A1(n3010), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3333) );
  AOI22_X1 U4228 ( .A1(n3008), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3332) );
  AOI22_X1 U4229 ( .A1(n3283), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n5326), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3331) );
  AOI22_X1 U4230 ( .A1(n3329), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3212), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3330) );
  NAND4_X1 U4231 ( .A1(n3333), .A2(n3332), .A3(n3331), .A4(n3330), .ZN(n3334)
         );
  NOR2_X1 U4232 ( .A1(n3364), .A2(n3505), .ZN(n3347) );
  NAND2_X1 U4233 ( .A1(n3347), .A2(n3449), .ZN(n3441) );
  OAI21_X1 U4234 ( .B1(n3449), .B2(n3418), .A(n3441), .ZN(n3340) );
  INV_X1 U4235 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3339) );
  AOI21_X1 U4236 ( .B1(n4232), .B2(n3505), .A(n6499), .ZN(n3338) );
  NAND2_X1 U4237 ( .A1(n3000), .A2(n3449), .ZN(n3337) );
  OAI211_X1 U4238 ( .C1(n3578), .C2(n3339), .A(n3338), .B(n3337), .ZN(n3440)
         );
  NAND2_X1 U4239 ( .A1(n3444), .A2(n3418), .ZN(n3342) );
  AND2_X1 U4240 ( .A1(n3444), .A2(n3418), .ZN(n3345) );
  NAND2_X1 U4241 ( .A1(n3345), .A2(n3344), .ZN(n3346) );
  NAND2_X1 U4242 ( .A1(n3352), .A2(n3346), .ZN(n3431) );
  NAND2_X1 U4243 ( .A1(n3586), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3351) );
  INV_X1 U4244 ( .A(n3347), .ZN(n3350) );
  INV_X1 U4245 ( .A(n3363), .ZN(n3348) );
  NAND2_X1 U4246 ( .A1(n3348), .A2(n3435), .ZN(n3349) );
  OAI21_X2 U4247 ( .B1(n3431), .B2(n3432), .A(n3352), .ZN(n3426) );
  INV_X1 U4248 ( .A(n3420), .ZN(n3377) );
  INV_X1 U4249 ( .A(n2996), .ZN(n3356) );
  INV_X1 U4250 ( .A(n3272), .ZN(n3357) );
  NAND2_X1 U4251 ( .A1(n3357), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3362) );
  NOR3_X1 U4252 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6471), .A3(n4838), 
        .ZN(n6363) );
  NAND2_X1 U4253 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6363), .ZN(n6439) );
  NAND2_X1 U4254 ( .A1(n6478), .A2(n6439), .ZN(n3358) );
  NOR3_X1 U4255 ( .A1(n6478), .A2(n6471), .A3(n4838), .ZN(n4710) );
  NAND2_X1 U4256 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4710), .ZN(n4557) );
  AOI22_X1 U4257 ( .A1(n3360), .A2(n4615), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3359), .ZN(n3361) );
  AOI22_X1 U4258 ( .A1(n5340), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3005), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3368) );
  AOI22_X1 U4259 ( .A1(n4119), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n5348), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3367) );
  AOI22_X1 U4260 ( .A1(n5349), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3382), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3366) );
  AOI22_X1 U4261 ( .A1(n5258), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n5350), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3365) );
  NAND4_X1 U4262 ( .A1(n3368), .A2(n3367), .A3(n3366), .A4(n3365), .ZN(n3374)
         );
  AOI22_X1 U4263 ( .A1(n4108), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3012), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3372) );
  AOI22_X1 U4264 ( .A1(n3011), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3017), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3371) );
  AOI22_X1 U4265 ( .A1(n5343), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3002), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3370) );
  AOI22_X1 U4266 ( .A1(n3391), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n5326), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3369) );
  NAND4_X1 U4267 ( .A1(n3372), .A2(n3371), .A3(n3370), .A4(n3369), .ZN(n3373)
         );
  AOI22_X1 U4268 ( .A1(n3586), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3590), 
        .B2(n3466), .ZN(n3375) );
  INV_X1 U4269 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3390) );
  AOI22_X1 U4270 ( .A1(n4108), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3005), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3381) );
  AOI22_X1 U4271 ( .A1(n5340), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n5348), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3380) );
  AOI22_X1 U4272 ( .A1(n4119), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3012), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3379) );
  AOI22_X1 U4273 ( .A1(n5349), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3003), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3378) );
  NAND4_X1 U4274 ( .A1(n3381), .A2(n3380), .A3(n3379), .A4(n3378), .ZN(n3388)
         );
  AOI22_X1 U4275 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n3011), .B1(n3016), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3386) );
  AOI22_X1 U4276 ( .A1(n3391), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n5350), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3385) );
  AOI22_X1 U4277 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n5258), .B1(n5326), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3384) );
  AOI22_X1 U4278 ( .A1(n3382), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3212), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3383) );
  NAND4_X1 U4279 ( .A1(n3386), .A2(n3385), .A3(n3384), .A4(n3383), .ZN(n3387)
         );
  NAND2_X1 U4280 ( .A1(n3590), .A2(n3485), .ZN(n3389) );
  INV_X1 U4281 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3403) );
  AOI22_X1 U4282 ( .A1(n4108), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3005), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3395) );
  AOI22_X1 U4283 ( .A1(n5340), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3382), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3394) );
  AOI22_X1 U4284 ( .A1(n3391), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n5258), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3393) );
  AOI22_X1 U4285 ( .A1(n3010), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n5350), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3392) );
  NAND4_X1 U4286 ( .A1(n3395), .A2(n3394), .A3(n3393), .A4(n3392), .ZN(n3401)
         );
  AOI22_X1 U4287 ( .A1(n4119), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n5348), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3399) );
  AOI22_X1 U4288 ( .A1(n5349), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3012), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3398) );
  AOI22_X1 U4289 ( .A1(n5343), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3002), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3397) );
  AOI22_X1 U4290 ( .A1(n2990), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n5326), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3396) );
  NAND4_X1 U4291 ( .A1(n3399), .A2(n3398), .A3(n3397), .A4(n3396), .ZN(n3400)
         );
  NAND2_X1 U4292 ( .A1(n3590), .A2(n3484), .ZN(n3402) );
  INV_X1 U4293 ( .A(n3483), .ZN(n3417) );
  INV_X1 U4294 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3416) );
  AOI22_X1 U4295 ( .A1(n4108), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3005), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3408) );
  AOI22_X1 U4296 ( .A1(n5340), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n5348), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3407) );
  AOI22_X1 U4297 ( .A1(n4119), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3012), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3406) );
  AOI22_X1 U4298 ( .A1(n5349), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3003), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3405) );
  NAND4_X1 U4299 ( .A1(n3408), .A2(n3407), .A3(n3406), .A4(n3405), .ZN(n3414)
         );
  AOI22_X1 U4300 ( .A1(n3011), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3412) );
  AOI22_X1 U4301 ( .A1(n3391), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n5350), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3411) );
  AOI22_X1 U4302 ( .A1(n5258), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n5326), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3410) );
  AOI22_X1 U4303 ( .A1(n3382), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3212), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3409) );
  NAND4_X1 U4304 ( .A1(n3412), .A2(n3411), .A3(n3410), .A4(n3409), .ZN(n3413)
         );
  NAND2_X1 U4305 ( .A1(n3590), .A2(n3498), .ZN(n3415) );
  NAND2_X1 U4306 ( .A1(n3221), .A2(n3014), .ZN(n3548) );
  NOR2_X1 U4307 ( .A1(n3418), .A2(n3548), .ZN(n3419) );
  NOR2_X1 U4308 ( .A1(n6249), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5678)
         );
  NOR2_X1 U4309 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5775) );
  AND2_X1 U4310 ( .A1(n5678), .A2(n5775), .ZN(n5665) );
  INV_X1 U4311 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5764) );
  NAND2_X1 U4312 ( .A1(n5665), .A2(n5764), .ZN(n3766) );
  INV_X1 U4313 ( .A(n3766), .ZN(n3531) );
  XNOR2_X2 U4314 ( .A(n3420), .B(n4334), .ZN(n3820) );
  NAND2_X1 U4315 ( .A1(n3820), .A2(n3445), .ZN(n3424) );
  NAND2_X1 U4316 ( .A1(n3435), .A2(n3449), .ZN(n3434) );
  NAND2_X1 U4317 ( .A1(n3434), .A2(n3427), .ZN(n3467) );
  INV_X1 U4318 ( .A(n3466), .ZN(n3421) );
  XNOR2_X1 U4319 ( .A(n3467), .B(n3421), .ZN(n3422) );
  NAND2_X1 U4320 ( .A1(n3422), .A2(n2989), .ZN(n3423) );
  INV_X1 U4321 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6360) );
  XNOR2_X1 U4322 ( .A(n3462), .B(n6360), .ZN(n6264) );
  NAND2_X1 U4323 ( .A1(n4331), .A2(n3445), .ZN(n3430) );
  XNOR2_X1 U4324 ( .A(n3434), .B(n3427), .ZN(n3428) );
  AND2_X1 U4325 ( .A1(n3000), .A2(n3238), .ZN(n3447) );
  AOI21_X1 U4326 ( .B1(n3428), .B2(n2989), .A(n3447), .ZN(n3429) );
  NAND2_X1 U4327 ( .A1(n3430), .A2(n3429), .ZN(n4563) );
  NAND2_X1 U4328 ( .A1(n4563), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3457)
         );
  INV_X1 U4329 ( .A(n3432), .ZN(n3433) );
  OAI21_X1 U4330 ( .B1(n3435), .B2(n3449), .A(n3434), .ZN(n3436) );
  INV_X1 U4331 ( .A(n3436), .ZN(n3438) );
  NAND3_X1 U4332 ( .A1(n3227), .A2(n3221), .A3(n3238), .ZN(n3437) );
  AOI21_X1 U4333 ( .B1(n3438), .B2(n2989), .A(n3437), .ZN(n3439) );
  INV_X1 U4334 ( .A(n3440), .ZN(n3442) );
  NAND2_X1 U4335 ( .A1(n3442), .A2(n3441), .ZN(n3443) );
  INV_X1 U4336 ( .A(n3548), .ZN(n3445) );
  NAND2_X1 U4337 ( .A1(n3446), .A2(n3445), .ZN(n3452) );
  INV_X1 U4338 ( .A(n2989), .ZN(n6612) );
  INV_X1 U4339 ( .A(n3447), .ZN(n3448) );
  OAI21_X1 U4340 ( .B1(n6612), .B2(n3449), .A(n3448), .ZN(n3450) );
  INV_X1 U4341 ( .A(n3450), .ZN(n3451) );
  NAND2_X1 U4342 ( .A1(n3452), .A2(n3451), .ZN(n4282) );
  NAND2_X1 U4343 ( .A1(n4282), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3453)
         );
  INV_X1 U4344 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4566) );
  NAND2_X1 U4345 ( .A1(n3453), .A2(n4566), .ZN(n3454) );
  AND2_X1 U4346 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4567) );
  NAND2_X1 U4347 ( .A1(n4282), .A2(n4567), .ZN(n3455) );
  INV_X1 U4348 ( .A(n3455), .ZN(n3456) );
  NAND2_X1 U4349 ( .A1(n3457), .A2(n4562), .ZN(n3461) );
  INV_X1 U4350 ( .A(n4563), .ZN(n3459) );
  INV_X1 U4351 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3458) );
  AND2_X1 U4352 ( .A1(n3461), .A2(n3460), .ZN(n6266) );
  NAND2_X1 U4353 ( .A1(n6264), .A2(n6266), .ZN(n6265) );
  NAND2_X1 U4354 ( .A1(n3462), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3463)
         );
  NAND2_X1 U4355 ( .A1(n6265), .A2(n3463), .ZN(n5047) );
  NAND2_X1 U4356 ( .A1(n3829), .A2(n3445), .ZN(n3470) );
  NAND2_X1 U4357 ( .A1(n3467), .A2(n3466), .ZN(n3487) );
  XNOR2_X1 U4358 ( .A(n3487), .B(n3485), .ZN(n3468) );
  NAND2_X1 U4359 ( .A1(n3468), .A2(n2989), .ZN(n3469) );
  INV_X1 U4360 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6350) );
  XNOR2_X1 U4361 ( .A(n3471), .B(n6350), .ZN(n5048) );
  NAND2_X1 U4362 ( .A1(n3471), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3472)
         );
  NAND2_X1 U4363 ( .A1(n5049), .A2(n3472), .ZN(n5055) );
  NAND2_X1 U4364 ( .A1(n3838), .A2(n3445), .ZN(n3479) );
  INV_X1 U4365 ( .A(n3485), .ZN(n3475) );
  OR2_X1 U4366 ( .A1(n3487), .A2(n3475), .ZN(n3476) );
  XNOR2_X1 U4367 ( .A(n3476), .B(n3484), .ZN(n3477) );
  NAND2_X1 U4368 ( .A1(n3477), .A2(n2989), .ZN(n3478) );
  NAND2_X1 U4369 ( .A1(n3479), .A2(n3478), .ZN(n3480) );
  INV_X1 U4370 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n6326) );
  XNOR2_X1 U4371 ( .A(n3480), .B(n6326), .ZN(n5057) );
  NAND2_X1 U4372 ( .A1(n3480), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3481)
         );
  NAND2_X1 U4373 ( .A1(n5058), .A2(n3481), .ZN(n4652) );
  NAND2_X1 U4374 ( .A1(n3843), .A2(n3445), .ZN(n3490) );
  NAND2_X1 U4375 ( .A1(n3485), .A2(n3484), .ZN(n3486) );
  OR2_X1 U4376 ( .A1(n3487), .A2(n3486), .ZN(n3497) );
  XNOR2_X1 U4377 ( .A(n3497), .B(n3498), .ZN(n3488) );
  NAND2_X1 U4378 ( .A1(n3488), .A2(n2989), .ZN(n3489) );
  NAND2_X1 U4379 ( .A1(n3490), .A2(n3489), .ZN(n3491) );
  INV_X1 U4380 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3637) );
  XNOR2_X1 U4381 ( .A(n3491), .B(n3637), .ZN(n4653) );
  NAND2_X1 U4382 ( .A1(n4652), .A2(n4653), .ZN(n4654) );
  NAND2_X1 U4383 ( .A1(n3491), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3492)
         );
  NAND2_X1 U4384 ( .A1(n4654), .A2(n3492), .ZN(n5066) );
  INV_X1 U4385 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3494) );
  NAND2_X1 U4386 ( .A1(n3590), .A2(n3505), .ZN(n3493) );
  OAI21_X1 U4387 ( .B1(n3578), .B2(n3494), .A(n3493), .ZN(n3495) );
  NAND2_X1 U4388 ( .A1(n3795), .A2(n3445), .ZN(n3502) );
  INV_X1 U4389 ( .A(n3497), .ZN(n3499) );
  NAND2_X1 U4390 ( .A1(n3499), .A2(n3498), .ZN(n3507) );
  XNOR2_X1 U4391 ( .A(n3507), .B(n3505), .ZN(n3500) );
  NAND2_X1 U4392 ( .A1(n3500), .A2(n2989), .ZN(n3501) );
  NAND2_X1 U4393 ( .A1(n3502), .A2(n3501), .ZN(n3503) );
  INV_X1 U4394 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6324) );
  XNOR2_X1 U4395 ( .A(n3503), .B(n6324), .ZN(n5069) );
  NAND2_X1 U4396 ( .A1(n5066), .A2(n5069), .ZN(n5067) );
  NAND2_X1 U4397 ( .A1(n3503), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3504)
         );
  NAND2_X1 U4398 ( .A1(n5067), .A2(n3504), .ZN(n5147) );
  INV_X1 U4399 ( .A(n3505), .ZN(n3506) );
  OR3_X1 U4400 ( .A1(n3507), .A2(n3506), .A3(n6612), .ZN(n3508) );
  NAND2_X1 U4401 ( .A1(n3513), .A2(n3508), .ZN(n3509) );
  INV_X1 U4402 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6315) );
  XNOR2_X1 U4403 ( .A(n3509), .B(n6315), .ZN(n5149) );
  NAND2_X1 U4404 ( .A1(n3509), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3510)
         );
  INV_X1 U4405 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5140) );
  NAND2_X1 U4406 ( .A1(n3513), .A2(n5140), .ZN(n3511) );
  NAND2_X1 U4407 ( .A1(n2988), .A2(n6290), .ZN(n5178) );
  INV_X1 U4408 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3512) );
  AND2_X1 U4409 ( .A1(n3513), .A2(n3512), .ZN(n3516) );
  NAND2_X1 U4410 ( .A1(n3789), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6248) );
  NAND2_X1 U4411 ( .A1(n3789), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3514) );
  AND2_X1 U4412 ( .A1(n6248), .A2(n3514), .ZN(n3515) );
  INV_X1 U4413 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5202) );
  NOR2_X1 U4414 ( .A1(n3513), .A2(n5202), .ZN(n5194) );
  NAND2_X1 U4415 ( .A1(n2988), .A2(n5202), .ZN(n5192) );
  XNOR2_X1 U4416 ( .A(n2988), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6008)
         );
  INV_X1 U4417 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3517) );
  NAND2_X1 U4418 ( .A1(n6249), .A2(n3517), .ZN(n3518) );
  INV_X1 U4419 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5219) );
  NAND2_X1 U4420 ( .A1(n3789), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3519) );
  INV_X1 U4421 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6022) );
  NOR2_X1 U4422 ( .A1(n6249), .A2(n6022), .ZN(n3521) );
  NAND2_X1 U4423 ( .A1(n6249), .A2(n6022), .ZN(n3522) );
  INV_X1 U4424 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5858) );
  NAND2_X1 U4425 ( .A1(n6249), .A2(n5858), .ZN(n5387) );
  NAND2_X1 U4426 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3742) );
  INV_X1 U4427 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5861) );
  INV_X1 U4428 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5854) );
  NAND3_X1 U4429 ( .A1(n5861), .A2(n5858), .A3(n5854), .ZN(n3524) );
  NAND2_X1 U4430 ( .A1(n3789), .A2(n3524), .ZN(n3525) );
  AND2_X1 U4431 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5813) );
  AND2_X1 U4432 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5833) );
  AND2_X1 U4433 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3748) );
  NAND3_X1 U4434 ( .A1(n5813), .A2(n5833), .A3(n3748), .ZN(n3526) );
  NAND2_X1 U4435 ( .A1(n6249), .A2(n3526), .ZN(n3527) );
  NOR2_X1 U4436 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5812) );
  NOR2_X1 U4437 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5403) );
  NOR2_X1 U4438 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5832) );
  NAND3_X1 U4439 ( .A1(n5812), .A2(n5403), .A3(n5832), .ZN(n3528) );
  NAND2_X1 U4440 ( .A1(n3789), .A2(n3528), .ZN(n3529) );
  INV_X1 U4441 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5802) );
  XNOR2_X1 U4442 ( .A(n6249), .B(n5802), .ZN(n5707) );
  NAND2_X1 U4443 ( .A1(n6249), .A2(n5802), .ZN(n3530) );
  NAND2_X1 U4444 ( .A1(n6249), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5697) );
  AND2_X1 U4445 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5774) );
  NAND2_X1 U4446 ( .A1(n5690), .A2(n5774), .ZN(n5667) );
  NOR2_X2 U4447 ( .A1(n5667), .A2(n5764), .ZN(n3768) );
  XNOR2_X1 U4448 ( .A(n3533), .B(n3532), .ZN(n5428) );
  NAND2_X1 U4449 ( .A1(n3612), .A2(n3000), .ZN(n3534) );
  INV_X1 U4450 ( .A(n4220), .ZN(n3540) );
  NAND2_X1 U4451 ( .A1(n3263), .A2(n3221), .ZN(n6463) );
  NAND2_X1 U4452 ( .A1(n6463), .A2(n3000), .ZN(n3536) );
  NAND2_X1 U4453 ( .A1(n2991), .A2(n2989), .ZN(n3537) );
  AND2_X1 U4454 ( .A1(n3538), .A2(n3537), .ZN(n3721) );
  NAND2_X1 U4455 ( .A1(n3613), .A2(n3721), .ZN(n3539) );
  NAND2_X1 U4456 ( .A1(n3540), .A2(n3539), .ZN(n3735) );
  NAND2_X1 U4457 ( .A1(n4838), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3542) );
  NAND2_X1 U4458 ( .A1(n3234), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3541) );
  NAND2_X1 U4459 ( .A1(n3542), .A2(n3541), .ZN(n3559) );
  NAND2_X1 U4460 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6364), .ZN(n3560) );
  NAND2_X1 U4461 ( .A1(n3543), .A2(n3542), .ZN(n3577) );
  NAND2_X1 U4462 ( .A1(n4256), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3544) );
  NAND2_X1 U4463 ( .A1(n3546), .A2(n3544), .ZN(n3576) );
  INV_X1 U4464 ( .A(n3576), .ZN(n3545) );
  NAND2_X1 U4465 ( .A1(n3577), .A2(n3545), .ZN(n3547) );
  NAND2_X1 U4466 ( .A1(n3547), .A2(n3546), .ZN(n3553) );
  XNOR2_X1 U4467 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3554) );
  OAI222_X1 U4468 ( .A1(n6040), .A2(n3549), .B1(n6040), .B2(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C1(n3549), .C2(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n3601) );
  NAND2_X1 U4469 ( .A1(n3601), .A2(n3575), .ZN(n3593) );
  NAND2_X1 U4470 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n3549), .ZN(n3550) );
  NOR2_X1 U4471 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n3550), .ZN(n3556)
         );
  INV_X1 U4472 ( .A(n3551), .ZN(n3552) );
  OAI21_X1 U4473 ( .B1(n3554), .B2(n3553), .A(n3552), .ZN(n3555) );
  AOI22_X1 U4474 ( .A1(n3575), .A2(n3557), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6499), .ZN(n3588) );
  INV_X1 U4475 ( .A(n3560), .ZN(n3558) );
  XNOR2_X1 U4476 ( .A(n3559), .B(n3558), .ZN(n3597) );
  AOI21_X1 U4477 ( .B1(n3590), .B2(n3014), .A(n3239), .ZN(n3572) );
  NAND2_X1 U4478 ( .A1(n3597), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3571) );
  NAND2_X1 U4479 ( .A1(n3572), .A2(n3571), .ZN(n3566) );
  NAND2_X1 U4480 ( .A1(n3078), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3561) );
  NAND2_X1 U4481 ( .A1(n3561), .A2(n3560), .ZN(n3567) );
  OAI21_X1 U4482 ( .B1(n3612), .B2(n3567), .A(n3562), .ZN(n3564) );
  NAND2_X1 U4483 ( .A1(n3239), .A2(n3230), .ZN(n3563) );
  NAND2_X1 U4484 ( .A1(n3563), .A2(n3013), .ZN(n3579) );
  NAND2_X1 U4485 ( .A1(n3564), .A2(n3579), .ZN(n3565) );
  NAND2_X1 U4486 ( .A1(n3566), .A2(n3565), .ZN(n3569) );
  NAND2_X1 U4487 ( .A1(n3597), .A2(n3569), .ZN(n3574) );
  INV_X1 U4488 ( .A(n3567), .ZN(n3568) );
  NAND2_X1 U4489 ( .A1(n3568), .A2(n3590), .ZN(n3570) );
  OAI22_X1 U4490 ( .A1(n3572), .A2(n3571), .B1(n3570), .B2(n3569), .ZN(n3573)
         );
  AOI21_X1 U4491 ( .B1(n3575), .B2(n3574), .A(n3573), .ZN(n3584) );
  XNOR2_X1 U4492 ( .A(n3577), .B(n3576), .ZN(n3599) );
  NOR2_X1 U4493 ( .A1(n3578), .A2(n3599), .ZN(n3580) );
  INV_X1 U4494 ( .A(n3579), .ZN(n3581) );
  AOI211_X1 U4495 ( .C1(n3590), .C2(n3599), .A(n3580), .B(n3581), .ZN(n3583)
         );
  NAND3_X1 U4496 ( .A1(n3581), .A2(n3590), .A3(n3599), .ZN(n3582) );
  OAI21_X1 U4497 ( .B1(n3584), .B2(n3583), .A(n3582), .ZN(n3585) );
  OAI21_X1 U4498 ( .B1(n3586), .B2(n3596), .A(n3585), .ZN(n3587) );
  NAND2_X1 U4499 ( .A1(n3588), .A2(n3587), .ZN(n3589) );
  INV_X1 U4500 ( .A(n6463), .ZN(n5375) );
  NAND3_X1 U4501 ( .A1(n4262), .A2(n5375), .A3(n3014), .ZN(n3594) );
  NAND2_X1 U4502 ( .A1(n3735), .A2(n3594), .ZN(n4260) );
  OR2_X1 U4503 ( .A1(n3595), .A2(STATE_REG_0__SCAN_IN), .ZN(n6523) );
  NAND2_X1 U4504 ( .A1(n3014), .A2(n6523), .ZN(n3602) );
  AND2_X1 U4505 ( .A1(n3597), .A2(n3596), .ZN(n3598) );
  AND2_X1 U4506 ( .A1(n3599), .A2(n3598), .ZN(n3600) );
  OR2_X1 U4507 ( .A1(n3601), .A2(n3600), .ZN(n4219) );
  NOR2_X1 U4508 ( .A1(READY_N), .A2(n4219), .ZN(n4261) );
  AND3_X1 U4509 ( .A1(n3602), .A2(n4261), .A3(n4431), .ZN(n3604) );
  OAI21_X1 U4510 ( .B1(n4260), .B2(n3604), .A(n4301), .ZN(n3608) );
  NAND2_X1 U4511 ( .A1(n3013), .A2(n6523), .ZN(n4182) );
  INV_X1 U4512 ( .A(READY_N), .ZN(n6735) );
  NAND2_X1 U4513 ( .A1(n4182), .A2(n6735), .ZN(n4268) );
  OAI211_X1 U4514 ( .C1(n3605), .C2(n4268), .A(n3230), .B(n5452), .ZN(n3606)
         );
  NAND3_X1 U4515 ( .A1(n4775), .A2(n3227), .A3(n3606), .ZN(n3607) );
  INV_X1 U4516 ( .A(n3605), .ZN(n4272) );
  AOI22_X1 U4517 ( .A1(n3611), .A2(n4524), .B1(n4272), .B2(n4233), .ZN(n3614)
         );
  AND2_X1 U4518 ( .A1(n3613), .A2(n3612), .ZN(n3794) );
  INV_X1 U4519 ( .A(n3794), .ZN(n6483) );
  NAND2_X1 U4520 ( .A1(n3613), .A2(n5029), .ZN(n4263) );
  NAND4_X1 U4521 ( .A1(n3610), .A2(n3614), .A3(n6483), .A4(n4263), .ZN(n3615)
         );
  INV_X1 U4522 ( .A(n3238), .ZN(n3616) );
  OR2_X1 U4523 ( .A1(n4229), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3618)
         );
  INV_X1 U4524 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5459) );
  NAND2_X1 U4525 ( .A1(n4233), .A2(n5459), .ZN(n3617) );
  NAND2_X1 U4526 ( .A1(n3618), .A2(n3617), .ZN(n3771) );
  INV_X1 U4527 ( .A(n3771), .ZN(n3714) );
  OR2_X2 U4528 ( .A1(n3628), .A2(n4298), .ZN(n3711) );
  NAND2_X1 U4529 ( .A1(n3707), .A2(n4566), .ZN(n3621) );
  INV_X1 U4530 ( .A(EBX_REG_1__SCAN_IN), .ZN(n3619) );
  NAND2_X1 U4531 ( .A1(n4233), .A2(n3619), .ZN(n3620) );
  NAND3_X1 U4532 ( .A1(n3621), .A2(n3770), .A3(n3620), .ZN(n3622) );
  NAND2_X1 U4533 ( .A1(n3707), .A2(EBX_REG_0__SCAN_IN), .ZN(n3624) );
  INV_X1 U4534 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5116) );
  NAND2_X1 U4535 ( .A1(n3770), .A2(n5116), .ZN(n3623) );
  MUX2_X1 U4536 ( .A(n3711), .B(n3707), .S(EBX_REG_2__SCAN_IN), .Z(n3627) );
  NAND2_X1 U4537 ( .A1(n3699), .A2(n4298), .ZN(n3702) );
  NAND2_X1 U4538 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n4298), .ZN(n3625)
         );
  AND2_X1 U4539 ( .A1(n3702), .A2(n3625), .ZN(n3626) );
  NAND2_X1 U4540 ( .A1(n3627), .A2(n3626), .ZN(n4327) );
  MUX2_X1 U4541 ( .A(n3712), .B(n3770), .S(EBX_REG_3__SCAN_IN), .Z(n3629) );
  OAI21_X1 U4542 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n4229), .A(n3629), 
        .ZN(n4318) );
  NAND2_X1 U4543 ( .A1(n3707), .A2(n6350), .ZN(n3632) );
  INV_X1 U4544 ( .A(EBX_REG_4__SCAN_IN), .ZN(n3630) );
  NAND2_X1 U4545 ( .A1(n4233), .A2(n3630), .ZN(n3631) );
  NAND3_X1 U4546 ( .A1(n3632), .A2(n3770), .A3(n3631), .ZN(n3633) );
  OAI21_X1 U4547 ( .B1(EBX_REG_4__SCAN_IN), .B2(n3711), .A(n3633), .ZN(n4448)
         );
  NAND2_X1 U4548 ( .A1(n4317), .A2(n4448), .ZN(n4456) );
  INV_X1 U4549 ( .A(n4456), .ZN(n3636) );
  MUX2_X1 U4550 ( .A(n3712), .B(n3770), .S(EBX_REG_5__SCAN_IN), .Z(n3634) );
  OAI21_X1 U4551 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n4229), .A(n3634), 
        .ZN(n4457) );
  INV_X1 U4552 ( .A(n3711), .ZN(n3700) );
  INV_X1 U4553 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6141) );
  NAND2_X1 U4554 ( .A1(n3700), .A2(n6141), .ZN(n3641) );
  NAND2_X1 U4555 ( .A1(n3707), .A2(n3637), .ZN(n3639) );
  NAND2_X1 U4556 ( .A1(n4233), .A2(n6141), .ZN(n3638) );
  NAND3_X1 U4557 ( .A1(n3639), .A2(n3770), .A3(n3638), .ZN(n3640) );
  MUX2_X1 U4558 ( .A(n3712), .B(n3770), .S(EBX_REG_7__SCAN_IN), .Z(n3642) );
  OAI21_X1 U4559 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n4229), .A(n3642), 
        .ZN(n5016) );
  NAND2_X1 U4560 ( .A1(n3707), .A2(n6315), .ZN(n3644) );
  INV_X1 U4561 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5157) );
  NAND2_X1 U4562 ( .A1(n4233), .A2(n5157), .ZN(n3643) );
  NAND3_X1 U4563 ( .A1(n3644), .A2(n3770), .A3(n3643), .ZN(n3645) );
  OAI21_X1 U4564 ( .B1(EBX_REG_8__SCAN_IN), .B2(n3711), .A(n3645), .ZN(n5133)
         );
  INV_X1 U4565 ( .A(n5136), .ZN(n3648) );
  MUX2_X1 U4566 ( .A(n3712), .B(n3770), .S(EBX_REG_9__SCAN_IN), .Z(n3646) );
  OAI21_X1 U4567 ( .B1(n4229), .B2(INSTADDRPOINTER_REG_9__SCAN_IN), .A(n3646), 
        .ZN(n4195) );
  MUX2_X1 U4568 ( .A(n3711), .B(n3707), .S(EBX_REG_10__SCAN_IN), .Z(n3651) );
  NAND2_X1 U4569 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n4298), .ZN(n3649) );
  AND2_X1 U4570 ( .A1(n3702), .A2(n3649), .ZN(n3650) );
  NAND2_X1 U4571 ( .A1(n3651), .A2(n3650), .ZN(n6113) );
  INV_X1 U4572 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6206) );
  NAND2_X1 U4573 ( .A1(n3674), .A2(n6206), .ZN(n3655) );
  NAND2_X1 U4574 ( .A1(n4233), .A2(n6206), .ZN(n3653) );
  NAND2_X1 U4575 ( .A1(n3770), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3652) );
  NAND3_X1 U4576 ( .A1(n3653), .A2(n3707), .A3(n3652), .ZN(n3654) );
  AND2_X1 U4577 ( .A1(n3655), .A2(n3654), .ZN(n6112) );
  NAND2_X1 U4578 ( .A1(n6113), .A2(n6112), .ZN(n3656) );
  MUX2_X1 U4579 ( .A(n3711), .B(n3707), .S(EBX_REG_12__SCAN_IN), .Z(n3659) );
  NAND2_X1 U4580 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n4298), .ZN(n3657) );
  AND2_X1 U4581 ( .A1(n3702), .A2(n3657), .ZN(n3658) );
  NAND2_X1 U4582 ( .A1(n3659), .A2(n3658), .ZN(n5204) );
  INV_X1 U4583 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6201) );
  NAND2_X1 U4584 ( .A1(n3674), .A2(n6201), .ZN(n3662) );
  NAND2_X1 U4585 ( .A1(n3770), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3660) );
  OAI211_X1 U4586 ( .C1(n4298), .C2(EBX_REG_13__SCAN_IN), .A(n3707), .B(n3660), 
        .ZN(n3661) );
  MUX2_X1 U4587 ( .A(n3711), .B(n3707), .S(EBX_REG_14__SCAN_IN), .Z(n3665) );
  NAND2_X1 U4588 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n4298), .ZN(n3663) );
  AND2_X1 U4589 ( .A1(n3702), .A2(n3663), .ZN(n3664) );
  NAND2_X1 U4590 ( .A1(n3665), .A2(n3664), .ZN(n5575) );
  INV_X1 U4591 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5631) );
  NAND2_X1 U4592 ( .A1(n3674), .A2(n5631), .ZN(n3669) );
  NAND2_X1 U4593 ( .A1(n4233), .A2(n5631), .ZN(n3667) );
  NAND2_X1 U4594 ( .A1(n3770), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3666) );
  NAND3_X1 U4595 ( .A1(n3667), .A2(n3707), .A3(n3666), .ZN(n3668) );
  AND2_X1 U4596 ( .A1(n3669), .A2(n3668), .ZN(n5576) );
  NAND2_X1 U4597 ( .A1(n5575), .A2(n5576), .ZN(n3670) );
  MUX2_X1 U4598 ( .A(n3700), .B(n3699), .S(EBX_REG_16__SCAN_IN), .Z(n3673) );
  NAND2_X1 U4599 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n4298), .ZN(n3671) );
  NAND2_X1 U4600 ( .A1(n3702), .A2(n3671), .ZN(n3672) );
  NOR2_X1 U4601 ( .A1(n3673), .A2(n3672), .ZN(n5628) );
  INV_X1 U4602 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5625) );
  NAND2_X1 U4603 ( .A1(n3674), .A2(n5625), .ZN(n3677) );
  NAND2_X1 U4604 ( .A1(n3628), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3675) );
  OAI211_X1 U4605 ( .C1(EBX_REG_17__SCAN_IN), .C2(n4298), .A(n3707), .B(n3675), 
        .ZN(n3676) );
  NAND2_X1 U4606 ( .A1(n3707), .A2(n5840), .ZN(n3680) );
  INV_X1 U4607 ( .A(EBX_REG_19__SCAN_IN), .ZN(n3678) );
  NAND2_X1 U4608 ( .A1(n4233), .A2(n3678), .ZN(n3679) );
  NAND3_X1 U4609 ( .A1(n3680), .A2(n3628), .A3(n3679), .ZN(n3681) );
  OAI21_X1 U4610 ( .B1(EBX_REG_19__SCAN_IN), .B2(n3711), .A(n3681), .ZN(n5549)
         );
  OR2_X1 U4611 ( .A1(n4229), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3683)
         );
  INV_X1 U4612 ( .A(EBX_REG_18__SCAN_IN), .ZN(n3682) );
  NAND2_X1 U4613 ( .A1(n4233), .A2(n3682), .ZN(n5545) );
  INV_X1 U4614 ( .A(n3770), .ZN(n5546) );
  OAI22_X1 U4615 ( .A1(n4229), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .B1(n4298), .B2(EBX_REG_20__SCAN_IN), .ZN(n5536) );
  NAND2_X1 U4616 ( .A1(n5548), .A2(n5536), .ZN(n3685) );
  NAND2_X1 U4617 ( .A1(n5546), .A2(EBX_REG_20__SCAN_IN), .ZN(n3684) );
  OAI211_X1 U4618 ( .C1(n5548), .C2(n5546), .A(n3685), .B(n3684), .ZN(n3686)
         );
  INV_X1 U4619 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5823) );
  NAND2_X1 U4620 ( .A1(n3707), .A2(n5823), .ZN(n3688) );
  INV_X1 U4621 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5976) );
  NAND2_X1 U4622 ( .A1(n4233), .A2(n5976), .ZN(n3687) );
  NAND3_X1 U4623 ( .A1(n3688), .A2(n3628), .A3(n3687), .ZN(n3689) );
  OAI21_X1 U4624 ( .B1(EBX_REG_21__SCAN_IN), .B2(n3711), .A(n3689), .ZN(n5610)
         );
  NAND2_X1 U4625 ( .A1(n5611), .A2(n5610), .ZN(n5609) );
  NAND2_X1 U4626 ( .A1(n3628), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3690) );
  OAI211_X1 U4627 ( .C1(n4298), .C2(EBX_REG_22__SCAN_IN), .A(n3707), .B(n3690), 
        .ZN(n3691) );
  OAI21_X1 U4628 ( .B1(n3712), .B2(EBX_REG_22__SCAN_IN), .A(n3691), .ZN(n5808)
         );
  MUX2_X1 U4629 ( .A(n3700), .B(n3699), .S(EBX_REG_23__SCAN_IN), .Z(n3694) );
  NAND2_X1 U4630 ( .A1(n4298), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3692) );
  NAND2_X1 U4631 ( .A1(n3702), .A2(n3692), .ZN(n3693) );
  NOR2_X1 U4632 ( .A1(n3694), .A2(n3693), .ZN(n5401) );
  INV_X1 U4633 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5956) );
  NAND2_X1 U4634 ( .A1(n4233), .A2(n5956), .ZN(n3696) );
  NAND2_X1 U4635 ( .A1(n3628), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3695) );
  NAND3_X1 U4636 ( .A1(n3696), .A2(n3707), .A3(n3695), .ZN(n3697) );
  OAI21_X1 U4637 ( .B1(n3712), .B2(EBX_REG_24__SCAN_IN), .A(n3697), .ZN(n5400)
         );
  NOR3_X2 U4638 ( .A1(n5806), .A2(n5401), .A3(n5400), .ZN(n3698) );
  MUX2_X1 U4639 ( .A(n3700), .B(n3699), .S(EBX_REG_25__SCAN_IN), .Z(n3704) );
  NAND2_X1 U4640 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n4298), .ZN(n3701) );
  NAND2_X1 U4641 ( .A1(n3702), .A2(n3701), .ZN(n3703) );
  NOR2_X1 U4642 ( .A1(n3704), .A2(n3703), .ZN(n5598) );
  MUX2_X1 U4643 ( .A(n3712), .B(n3628), .S(EBX_REG_26__SCAN_IN), .Z(n3706) );
  OR2_X1 U4644 ( .A1(n4229), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3705)
         );
  AND2_X1 U4645 ( .A1(n3706), .A2(n3705), .ZN(n5515) );
  INV_X1 U4646 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5785) );
  NAND2_X1 U4647 ( .A1(n3707), .A2(n5785), .ZN(n3709) );
  INV_X1 U4648 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U4649 ( .A1(n4233), .A2(n5588), .ZN(n3708) );
  NAND3_X1 U4650 ( .A1(n3709), .A2(n3628), .A3(n3708), .ZN(n3710) );
  OAI21_X1 U4651 ( .B1(EBX_REG_27__SCAN_IN), .B2(n3711), .A(n3710), .ZN(n5501)
         );
  MUX2_X1 U4652 ( .A(n3712), .B(n3628), .S(EBX_REG_28__SCAN_IN), .Z(n3713) );
  OAI21_X1 U4653 ( .B1(INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n4229), .A(n3713), 
        .ZN(n5487) );
  OAI21_X1 U4654 ( .B1(n3714), .B2(n5489), .A(n3774), .ZN(n3717) );
  NAND2_X1 U4655 ( .A1(n4229), .A2(EBX_REG_30__SCAN_IN), .ZN(n3716) );
  NAND2_X1 U4656 ( .A1(n4298), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3715) );
  NAND2_X1 U4657 ( .A1(n3716), .A2(n3715), .ZN(n3775) );
  XNOR2_X1 U4658 ( .A(n3717), .B(n3775), .ZN(n5479) );
  NAND2_X1 U4659 ( .A1(n4272), .A2(n2989), .ZN(n6495) );
  NAND2_X1 U4660 ( .A1(n3611), .A2(n4232), .ZN(n3718) );
  NAND2_X1 U4661 ( .A1(n6495), .A2(n3718), .ZN(n3719) );
  OR2_X2 U4662 ( .A1(n4151), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6341) );
  INV_X1 U4663 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6716) );
  NOR2_X1 U4664 ( .A1(n6341), .A2(n6716), .ZN(n5422) );
  AND2_X1 U4665 ( .A1(n4220), .A2(n3014), .ZN(n4774) );
  NAND2_X1 U4666 ( .A1(n3736), .A2(n4774), .ZN(n5224) );
  INV_X1 U4667 ( .A(n4229), .ZN(n3777) );
  OAI21_X1 U4668 ( .B1(n3535), .B2(n3777), .A(n3721), .ZN(n3722) );
  INV_X1 U4669 ( .A(n3722), .ZN(n3723) );
  NAND2_X1 U4670 ( .A1(n3720), .A2(n3723), .ZN(n4244) );
  INV_X1 U4671 ( .A(n3006), .ZN(n3725) );
  OR2_X1 U4672 ( .A1(n6463), .A2(n3725), .ZN(n4466) );
  OAI21_X1 U4673 ( .B1(n3724), .B2(n3726), .A(n4466), .ZN(n3727) );
  OR2_X1 U4674 ( .A1(n4244), .A2(n3727), .ZN(n3728) );
  NAND2_X1 U4675 ( .A1(n3736), .A2(n3728), .ZN(n4284) );
  NAND4_X1 U4676 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .A3(INSTADDRPOINTER_REG_3__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6328) );
  NAND2_X1 U4677 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3729) );
  NOR2_X1 U4678 ( .A1(n6328), .A2(n3729), .ZN(n5199) );
  INV_X1 U4679 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6290) );
  NAND2_X1 U4680 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6312) );
  NOR3_X1 U4681 ( .A1(n5140), .A2(n6290), .A3(n6312), .ZN(n3737) );
  NAND2_X1 U4682 ( .A1(n5199), .A2(n3737), .ZN(n3753) );
  NAND2_X1 U4683 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6026) );
  NOR2_X1 U4684 ( .A1(n3517), .A2(n6026), .ZN(n5226) );
  NAND2_X1 U4685 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5226), .ZN(n6011) );
  NAND2_X1 U4686 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6015) );
  NOR2_X1 U4687 ( .A1(n6011), .A2(n6015), .ZN(n3738) );
  INV_X1 U4688 ( .A(n3738), .ZN(n3730) );
  NOR2_X1 U4689 ( .A1(n3753), .A2(n3730), .ZN(n3731) );
  OR2_X1 U4690 ( .A1(n5200), .A2(n3731), .ZN(n3741) );
  OR2_X1 U4691 ( .A1(n4284), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3732)
         );
  INV_X2 U4692 ( .A(n6341), .ZN(n6351) );
  OR2_X1 U4693 ( .A1(n3736), .A2(n6351), .ZN(n4312) );
  OR2_X1 U4694 ( .A1(n4225), .A2(n4431), .ZN(n4266) );
  NAND2_X1 U4695 ( .A1(n4266), .A2(n3014), .ZN(n3733) );
  NOR2_X1 U4696 ( .A1(n6463), .A2(n3733), .ZN(n3734) );
  NAND2_X1 U4697 ( .A1(n3735), .A2(n3734), .ZN(n4247) );
  INV_X1 U4698 ( .A(n4247), .ZN(n4216) );
  INV_X1 U4699 ( .A(n3737), .ZN(n5201) );
  AOI21_X1 U4700 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6346) );
  NAND2_X1 U4701 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6347) );
  NOR2_X1 U4702 ( .A1(n6346), .A2(n6347), .ZN(n6330) );
  NAND3_X1 U4703 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n6330), .ZN(n6289) );
  NOR2_X1 U4704 ( .A1(n5201), .A2(n6289), .ZN(n3755) );
  NAND2_X1 U4705 ( .A1(n3755), .A2(n3738), .ZN(n3739) );
  NAND2_X1 U4706 ( .A1(n6339), .A2(n3739), .ZN(n3740) );
  INV_X1 U4707 ( .A(n6339), .ZN(n4285) );
  INV_X1 U4708 ( .A(n3742), .ZN(n3758) );
  AND2_X1 U4709 ( .A1(n3758), .A2(n5833), .ZN(n3743) );
  OR2_X1 U4710 ( .A1(n6296), .A2(n3743), .ZN(n3744) );
  NAND2_X1 U4711 ( .A1(n5863), .A2(n3744), .ZN(n5819) );
  NOR2_X1 U4712 ( .A1(n6296), .A2(n5813), .ZN(n3745) );
  NOR2_X1 U4713 ( .A1(n5819), .A2(n3745), .ZN(n4165) );
  INV_X1 U4714 ( .A(n5200), .ZN(n3746) );
  INV_X1 U4715 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4286) );
  NAND2_X1 U4716 ( .A1(n5224), .A2(n4286), .ZN(n4309) );
  NAND2_X1 U4717 ( .A1(n3746), .A2(n4309), .ZN(n6327) );
  INV_X1 U4718 ( .A(n6327), .ZN(n3747) );
  INV_X1 U4719 ( .A(n3748), .ZN(n3760) );
  NAND2_X1 U4720 ( .A1(n5827), .A2(n3760), .ZN(n3749) );
  NAND2_X1 U4721 ( .A1(n4165), .A2(n3749), .ZN(n5799) );
  INV_X1 U4722 ( .A(n5774), .ZN(n3750) );
  NAND2_X1 U4723 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5769) );
  OR3_X1 U4724 ( .A1(n5799), .A2(n3750), .A3(n5769), .ZN(n3751) );
  NAND2_X1 U4725 ( .A1(n6296), .A2(n5196), .ZN(n5768) );
  NAND2_X1 U4726 ( .A1(n3751), .A2(n5768), .ZN(n5760) );
  INV_X1 U4727 ( .A(n5768), .ZN(n5203) );
  AOI211_X1 U4728 ( .C1(n5760), .C2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5203), .B(n3532), .ZN(n3752) );
  AOI211_X1 U4729 ( .C1(n5479), .C2(n6353), .A(n5422), .B(n3752), .ZN(n3763)
         );
  NOR2_X1 U4730 ( .A1(n5224), .A2(n3753), .ZN(n6028) );
  NOR3_X1 U4731 ( .A1(n4284), .A2(n3753), .A3(n4286), .ZN(n3754) );
  AOI21_X1 U4732 ( .B1(n3755), .B2(n6339), .A(n3754), .ZN(n5221) );
  INV_X1 U4733 ( .A(n5221), .ZN(n3756) );
  AND2_X1 U4734 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3757) );
  INV_X1 U4735 ( .A(n5833), .ZN(n3759) );
  NAND2_X1 U4736 ( .A1(n5824), .A2(n5813), .ZN(n5406) );
  NAND2_X1 U4737 ( .A1(n5774), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3761) );
  NOR2_X1 U4738 ( .A1(n5776), .A2(n3761), .ZN(n3779) );
  NAND2_X1 U4739 ( .A1(n3779), .A2(n3532), .ZN(n3762) );
  OAI21_X1 U4740 ( .B1(n5428), .B2(n6283), .A(n3764), .ZN(U2988) );
  INV_X1 U4741 ( .A(n3765), .ZN(n5706) );
  NOR2_X1 U4742 ( .A1(n3766), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3767)
         );
  AOI22_X1 U4743 ( .A1(n3768), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .B1(n5706), .B2(n3767), .ZN(n3769) );
  INV_X1 U4744 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4255) );
  XNOR2_X1 U4745 ( .A(n3769), .B(n4255), .ZN(n5421) );
  NAND2_X1 U4746 ( .A1(n3771), .A2(n3628), .ZN(n3773) );
  NAND2_X1 U4747 ( .A1(n5546), .A2(EBX_REG_29__SCAN_IN), .ZN(n3772) );
  AND2_X1 U4748 ( .A1(n3773), .A2(n3772), .ZN(n5433) );
  NOR2_X1 U4749 ( .A1(n4298), .A2(EBX_REG_31__SCAN_IN), .ZN(n3776) );
  AOI21_X1 U4750 ( .B1(n3777), .B2(n4255), .A(n3776), .ZN(n3778) );
  NAND2_X1 U4751 ( .A1(n5583), .A2(n6353), .ZN(n3784) );
  NAND3_X1 U4752 ( .A1(n3779), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n4255), .ZN(n3783) );
  AND2_X1 U4753 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3780) );
  OAI21_X1 U4754 ( .B1(n6296), .B2(n3780), .A(n5760), .ZN(n3781) );
  INV_X1 U4755 ( .A(REIP_REG_31__SCAN_IN), .ZN(n5469) );
  NOR2_X1 U4756 ( .A1(n6341), .A2(n5469), .ZN(n5416) );
  AOI21_X1 U4757 ( .B1(n3781), .B2(INSTADDRPOINTER_REG_31__SCAN_IN), .A(n5416), 
        .ZN(n3782) );
  OAI21_X1 U4758 ( .B1(n5421), .B2(n6283), .A(n3785), .ZN(U2987) );
  INV_X1 U4759 ( .A(n5735), .ZN(n4160) );
  NAND2_X1 U4760 ( .A1(n3787), .A2(n5840), .ZN(n3788) );
  XNOR2_X1 U4761 ( .A(n3789), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5729)
         );
  INV_X1 U4762 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5831) );
  XNOR2_X1 U4763 ( .A(n6249), .B(n5823), .ZN(n5723) );
  INV_X1 U4764 ( .A(n3791), .ZN(n5722) );
  NOR2_X1 U4765 ( .A1(n6249), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5712)
         );
  NAND2_X1 U4766 ( .A1(n5722), .A2(n5712), .ZN(n4162) );
  NAND3_X1 U4767 ( .A1(n6249), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3792) );
  XNOR2_X1 U4768 ( .A(n3793), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5410)
         );
  INV_X2 U4769 ( .A(n6276), .ZN(n6269) );
  CLKBUF_X1 U4770 ( .A(n3222), .Z(n5454) );
  NOR2_X2 U4771 ( .A1(n5454), .A2(n6498), .ZN(n3809) );
  INV_X1 U4772 ( .A(EAX_REG_7__SCAN_IN), .ZN(n4388) );
  XNOR2_X1 U4773 ( .A(n3859), .B(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5071) );
  NAND2_X1 U4774 ( .A1(n6498), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4146) );
  INV_X1 U4775 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5019) );
  NOR2_X1 U4776 ( .A1(n4146), .A2(n5019), .ZN(n3797) );
  AOI21_X1 U4777 ( .B1(n5071), .B2(n5369), .A(n3797), .ZN(n3798) );
  OAI21_X1 U4778 ( .B1(n4006), .B2(n4388), .A(n3798), .ZN(n3799) );
  NAND2_X1 U4779 ( .A1(n4331), .A2(n3985), .ZN(n3800) );
  NAND2_X1 U4780 ( .A1(n3800), .A2(n4146), .ZN(n3817) );
  NAND2_X1 U4781 ( .A1(n4332), .A2(n3985), .ZN(n3804) );
  INV_X1 U4782 ( .A(n4006), .ZN(n5364) );
  AOI22_X1 U4783 ( .A1(n5364), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6498), .ZN(n3802) );
  NOR2_X1 U4784 ( .A1(n5452), .A2(n6498), .ZN(n3830) );
  NAND2_X1 U4785 ( .A1(n3830), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3801) );
  AND2_X1 U4786 ( .A1(n3802), .A2(n3801), .ZN(n3803) );
  NAND2_X1 U4787 ( .A1(n3804), .A2(n3803), .ZN(n4295) );
  NAND2_X1 U4788 ( .A1(n4975), .A2(n3805), .ZN(n3806) );
  NAND2_X1 U4789 ( .A1(n3806), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4240) );
  INV_X1 U4791 ( .A(n3830), .ZN(n3825) );
  NAND2_X1 U4792 ( .A1(PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n6498), .ZN(n3811)
         );
  NAND2_X1 U4793 ( .A1(n3809), .A2(EAX_REG_0__SCAN_IN), .ZN(n3810) );
  OAI211_X1 U4794 ( .C1(n3825), .C2(n3078), .A(n3811), .B(n3810), .ZN(n3812)
         );
  AOI21_X1 U4795 ( .B1(n3808), .B2(n3985), .A(n3812), .ZN(n4241) );
  OR2_X1 U4796 ( .A1(n4240), .A2(n4241), .ZN(n4238) );
  NAND2_X1 U4797 ( .A1(n4241), .A2(n5369), .ZN(n3813) );
  NAND2_X1 U4798 ( .A1(n4238), .A2(n3813), .ZN(n4294) );
  OAI21_X1 U4799 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3814), .ZN(n6280) );
  AOI22_X1 U4800 ( .A1(n5413), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n5369), 
        .B2(n6280), .ZN(n3816) );
  NAND2_X1 U4801 ( .A1(n5364), .A2(EAX_REG_2__SCAN_IN), .ZN(n3815) );
  OAI211_X1 U4802 ( .C1(n3825), .C2(n4256), .A(n3816), .B(n3815), .ZN(n4323)
         );
  NAND2_X1 U4803 ( .A1(n4324), .A2(n4323), .ZN(n3819) );
  NAND2_X1 U4804 ( .A1(n3817), .A2(n4297), .ZN(n3818) );
  NAND2_X1 U4805 ( .A1(n3820), .A2(n3985), .ZN(n3828) );
  OAI21_X1 U4806 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3822), .A(n3821), 
        .ZN(n6273) );
  AOI22_X1 U4807 ( .A1(n5369), .A2(n6273), .B1(n5413), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3824) );
  NAND2_X1 U4808 ( .A1(n5364), .A2(EAX_REG_3__SCAN_IN), .ZN(n3823) );
  OAI211_X1 U4809 ( .C1(n3825), .C2(n3079), .A(n3824), .B(n3823), .ZN(n3826)
         );
  INV_X1 U4810 ( .A(n3826), .ZN(n3827) );
  NAND2_X1 U4811 ( .A1(n3828), .A2(n3827), .ZN(n4320) );
  NAND2_X1 U4812 ( .A1(n3830), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3836) );
  INV_X1 U4813 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3831) );
  AOI21_X1 U4814 ( .B1(n3831), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3832) );
  AOI21_X1 U4815 ( .B1(n5364), .B2(EAX_REG_4__SCAN_IN), .A(n3832), .ZN(n3835)
         );
  NOR2_X1 U4816 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n3833), .ZN(n3834)
         );
  NOR2_X1 U4817 ( .A1(n3839), .A2(n3834), .ZN(n5050) );
  AOI22_X1 U4818 ( .A1(n3836), .A2(n3835), .B1(n5369), .B2(n5050), .ZN(n3837)
         );
  NAND2_X1 U4819 ( .A1(n3838), .A2(n3985), .ZN(n3842) );
  INV_X1 U4820 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5035) );
  XNOR2_X1 U4821 ( .A(n3839), .B(n5035), .ZN(n5060) );
  OAI22_X1 U4822 ( .A1(n5060), .A2(n5362), .B1(n4146), .B2(n5035), .ZN(n3840)
         );
  AOI21_X1 U4823 ( .B1(n5364), .B2(EAX_REG_5__SCAN_IN), .A(n3840), .ZN(n3841)
         );
  NAND2_X1 U4824 ( .A1(n4445), .A2(n4453), .ZN(n4452) );
  AND2_X1 U4825 ( .A1(n3844), .A2(n6137), .ZN(n3845) );
  OR2_X1 U4826 ( .A1(n3845), .A2(n3859), .ZN(n6262) );
  INV_X1 U4827 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4364) );
  OAI22_X1 U4828 ( .A1(n4006), .A2(n4364), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6137), .ZN(n3846) );
  MUX2_X1 U4829 ( .A(n6262), .B(n3846), .S(n5362), .Z(n3847) );
  NAND2_X1 U4830 ( .A1(n3848), .A2(n4604), .ZN(n5124) );
  AOI22_X1 U4831 ( .A1(n3190), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n5348), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3852) );
  AOI22_X1 U4832 ( .A1(n4119), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3003), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3851) );
  AOI22_X1 U4833 ( .A1(n3391), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n5326), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3850) );
  AOI22_X1 U4834 ( .A1(n3382), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3212), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3849) );
  NAND4_X1 U4835 ( .A1(n3852), .A2(n3851), .A3(n3850), .A4(n3849), .ZN(n3858)
         );
  AOI22_X1 U4836 ( .A1(n5340), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3856) );
  AOI22_X1 U4837 ( .A1(n5349), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3012), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4838 ( .A1(n3010), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3017), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3854) );
  AOI22_X1 U4839 ( .A1(n5258), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n5350), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3853) );
  NAND4_X1 U4840 ( .A1(n3856), .A2(n3855), .A3(n3854), .A4(n3853), .ZN(n3857)
         );
  OAI21_X1 U4841 ( .B1(n3858), .B2(n3857), .A(n3985), .ZN(n3863) );
  NAND2_X1 U4842 ( .A1(n3809), .A2(EAX_REG_8__SCAN_IN), .ZN(n3862) );
  XNOR2_X1 U4843 ( .A(n3864), .B(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5159) );
  NAND2_X1 U4844 ( .A1(n5159), .A2(n5369), .ZN(n3861) );
  NAND2_X1 U4845 ( .A1(n5413), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3860)
         );
  XOR2_X1 U4846 ( .A(n4188), .B(n3878), .Z(n5143) );
  AOI22_X1 U4847 ( .A1(n4108), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n5348), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3868) );
  AOI22_X1 U4848 ( .A1(n4119), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3012), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3867) );
  AOI22_X1 U4849 ( .A1(n5349), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3003), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3866) );
  AOI22_X1 U4850 ( .A1(n3382), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3212), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3865) );
  NAND4_X1 U4851 ( .A1(n3868), .A2(n3867), .A3(n3866), .A4(n3865), .ZN(n3874)
         );
  AOI22_X1 U4852 ( .A1(n5340), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3005), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3872) );
  AOI22_X1 U4853 ( .A1(n3011), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3871) );
  AOI22_X1 U4854 ( .A1(n3391), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n5350), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3870) );
  AOI22_X1 U4855 ( .A1(n5258), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n5326), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3869) );
  NAND4_X1 U4856 ( .A1(n3872), .A2(n3871), .A3(n3870), .A4(n3869), .ZN(n3873)
         );
  OR2_X1 U4857 ( .A1(n3874), .A2(n3873), .ZN(n3875) );
  AOI22_X1 U4858 ( .A1(n3985), .A2(n3875), .B1(n5413), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3877) );
  NAND2_X1 U4859 ( .A1(n3809), .A2(EAX_REG_9__SCAN_IN), .ZN(n3876) );
  OAI211_X1 U4860 ( .C1(n5143), .C2(n5362), .A(n3877), .B(n3876), .ZN(n4198)
         );
  INV_X1 U4861 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n6124) );
  XNOR2_X1 U4862 ( .A(n3891), .B(n6124), .ZN(n6132) );
  AOI22_X1 U4863 ( .A1(n3809), .A2(EAX_REG_10__SCAN_IN), .B1(n5413), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4864 ( .A1(n4108), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n5348), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3882) );
  AOI22_X1 U4865 ( .A1(n3011), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3382), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3881) );
  AOI22_X1 U4866 ( .A1(n4119), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3880) );
  AOI22_X1 U4867 ( .A1(n5258), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n5350), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3879) );
  NAND4_X1 U4868 ( .A1(n3882), .A2(n3881), .A3(n3880), .A4(n3879), .ZN(n3888)
         );
  AOI22_X1 U4869 ( .A1(n5340), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3005), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3886) );
  AOI22_X1 U4870 ( .A1(n5349), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3012), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3885) );
  AOI22_X1 U4871 ( .A1(n2990), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3003), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3884) );
  AOI22_X1 U4872 ( .A1(n3391), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n5326), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3883) );
  NAND4_X1 U4873 ( .A1(n3886), .A2(n3885), .A3(n3884), .A4(n3883), .ZN(n3887)
         );
  OAI21_X1 U4874 ( .B1(n3888), .B2(n3887), .A(n3985), .ZN(n3889) );
  OAI211_X1 U4875 ( .C1(n6132), .C2(n5362), .A(n3890), .B(n3889), .ZN(n5129)
         );
  XOR2_X1 U4876 ( .A(n3907), .B(n3908), .Z(n6252) );
  INV_X1 U4877 ( .A(n6252), .ZN(n3906) );
  AOI22_X1 U4878 ( .A1(n5348), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3012), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3895) );
  AOI22_X1 U4879 ( .A1(n3011), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n2990), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3894) );
  AOI22_X1 U4880 ( .A1(n3382), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3212), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3893) );
  AOI22_X1 U4881 ( .A1(n5350), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n5326), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3892) );
  NAND4_X1 U4882 ( .A1(n3895), .A2(n3894), .A3(n3893), .A4(n3892), .ZN(n3901)
         );
  AOI22_X1 U4883 ( .A1(n4108), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3005), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3899) );
  AOI22_X1 U4884 ( .A1(n5340), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4119), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3898) );
  AOI22_X1 U4885 ( .A1(n3391), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n5258), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3897) );
  AOI22_X1 U4886 ( .A1(n5349), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n5343), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3896) );
  NAND4_X1 U4887 ( .A1(n3899), .A2(n3898), .A3(n3897), .A4(n3896), .ZN(n3900)
         );
  OAI21_X1 U4888 ( .B1(n3901), .B2(n3900), .A(n3985), .ZN(n3904) );
  NAND2_X1 U4889 ( .A1(n3809), .A2(EAX_REG_11__SCAN_IN), .ZN(n3903) );
  NAND2_X1 U4890 ( .A1(n5413), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3902)
         );
  NAND3_X1 U4891 ( .A1(n3904), .A2(n3903), .A3(n3902), .ZN(n3905) );
  AOI21_X1 U4892 ( .B1(n3906), .B2(n5369), .A(n3905), .ZN(n5185) );
  INV_X1 U4893 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3909) );
  XNOR2_X1 U4894 ( .A(n3927), .B(n3909), .ZN(n6107) );
  NAND2_X1 U4895 ( .A1(n6107), .A2(n5369), .ZN(n3925) );
  INV_X1 U4896 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6226) );
  INV_X1 U4897 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6728) );
  OAI21_X1 U4898 ( .B1(n6728), .B2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n6498), 
        .ZN(n3910) );
  OAI21_X1 U4899 ( .B1(n4006), .B2(n6226), .A(n3910), .ZN(n3924) );
  INV_X1 U4900 ( .A(n3985), .ZN(n3922) );
  AOI22_X1 U4901 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n5340), .B1(n5348), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3914) );
  AOI22_X1 U4902 ( .A1(n4119), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3913) );
  AOI22_X1 U4903 ( .A1(n3010), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3002), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3912) );
  AOI22_X1 U4904 ( .A1(n5258), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n5350), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3911) );
  NAND4_X1 U4905 ( .A1(n3914), .A2(n3913), .A3(n3912), .A4(n3911), .ZN(n3920)
         );
  AOI22_X1 U4906 ( .A1(n4108), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3005), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3918) );
  AOI22_X1 U4907 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n2990), .B1(n3382), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3917) );
  AOI22_X1 U4908 ( .A1(n5349), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n5343), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3916) );
  AOI22_X1 U4909 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(n3391), .B1(n5326), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3915) );
  NAND4_X1 U4910 ( .A1(n3918), .A2(n3917), .A3(n3916), .A4(n3915), .ZN(n3919)
         );
  NOR2_X1 U4911 ( .A1(n3920), .A2(n3919), .ZN(n3921) );
  NOR2_X1 U4912 ( .A1(n3922), .A2(n3921), .ZN(n3923) );
  AOI21_X1 U4913 ( .B1(n3925), .B2(n3924), .A(n3923), .ZN(n5189) );
  INV_X1 U4914 ( .A(n5189), .ZN(n3926) );
  AND2_X2 U4915 ( .A1(n5183), .A2(n3926), .ZN(n3932) );
  NAND2_X1 U4916 ( .A1(n3809), .A2(EAX_REG_13__SCAN_IN), .ZN(n3930) );
  OAI21_X1 U4917 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n3928), .A(n3947), 
        .ZN(n6101) );
  AOI22_X1 U4918 ( .A1(n5369), .A2(n6101), .B1(n5413), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3929) );
  NAND2_X1 U4919 ( .A1(n3930), .A2(n3929), .ZN(n3931) );
  AOI22_X1 U4920 ( .A1(n3190), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n5348), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3937) );
  AOI22_X1 U4921 ( .A1(n4119), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3012), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3936) );
  AOI22_X1 U4922 ( .A1(n5349), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3011), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3935) );
  AOI22_X1 U4923 ( .A1(n3391), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n5258), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3934) );
  NAND4_X1 U4924 ( .A1(n3937), .A2(n3936), .A3(n3935), .A4(n3934), .ZN(n3943)
         );
  AOI22_X1 U4925 ( .A1(n5340), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3941) );
  AOI22_X1 U4926 ( .A1(n3382), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3017), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3940) );
  AOI22_X1 U4927 ( .A1(n3003), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3212), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3939) );
  AOI22_X1 U4928 ( .A1(n5350), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n5326), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3938) );
  NAND4_X1 U4929 ( .A1(n3941), .A2(n3940), .A3(n3939), .A4(n3938), .ZN(n3942)
         );
  OR2_X1 U4930 ( .A1(n3943), .A2(n3942), .ZN(n3944) );
  NAND2_X1 U4931 ( .A1(n3985), .A2(n3944), .ZN(n5231) );
  XOR2_X1 U4932 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3961), .Z(n6087) );
  AOI22_X1 U4933 ( .A1(n4108), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n5348), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3951) );
  AOI22_X1 U4934 ( .A1(n3382), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n2990), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3950) );
  AOI22_X1 U4935 ( .A1(n3391), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n5258), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3949) );
  AOI22_X1 U4936 ( .A1(n4119), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n5343), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3948) );
  NAND4_X1 U4937 ( .A1(n3951), .A2(n3950), .A3(n3949), .A4(n3948), .ZN(n3957)
         );
  AOI22_X1 U4938 ( .A1(n5340), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3005), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3955) );
  AOI22_X1 U4939 ( .A1(n5349), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3012), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3954) );
  AOI22_X1 U4940 ( .A1(n3011), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3002), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3953) );
  AOI22_X1 U4941 ( .A1(n5350), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n5326), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3952) );
  NAND4_X1 U4942 ( .A1(n3955), .A2(n3954), .A3(n3953), .A4(n3952), .ZN(n3956)
         );
  OR2_X1 U4943 ( .A1(n3957), .A2(n3956), .ZN(n3958) );
  AOI22_X1 U4944 ( .A1(n3985), .A2(n3958), .B1(n5413), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3960) );
  NAND2_X1 U4945 ( .A1(n3809), .A2(EAX_REG_14__SCAN_IN), .ZN(n3959) );
  OAI211_X1 U4946 ( .C1(n6087), .C2(n5362), .A(n3960), .B(n3959), .ZN(n5634)
         );
  XOR2_X1 U4947 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n3993), .Z(n6078) );
  INV_X1 U4948 ( .A(n6078), .ZN(n3975) );
  AOI22_X1 U4949 ( .A1(n4119), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3965) );
  AOI22_X1 U4950 ( .A1(n3382), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n2990), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3964) );
  AOI22_X1 U4951 ( .A1(n3012), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3002), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3963) );
  AOI22_X1 U4952 ( .A1(n3391), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3004), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3962) );
  NAND4_X1 U4953 ( .A1(n3965), .A2(n3964), .A3(n3963), .A4(n3962), .ZN(n3971)
         );
  AOI22_X1 U4954 ( .A1(n5340), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3005), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3969) );
  AOI22_X1 U4955 ( .A1(n5349), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n5348), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3968) );
  AOI22_X1 U4956 ( .A1(n3010), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n5343), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3967) );
  AOI22_X1 U4957 ( .A1(n5258), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n5326), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3966) );
  NAND4_X1 U4958 ( .A1(n3969), .A2(n3968), .A3(n3967), .A4(n3966), .ZN(n3970)
         );
  NOR2_X1 U4959 ( .A1(n3971), .A2(n3970), .ZN(n3973) );
  AOI22_X1 U4960 ( .A1(n3809), .A2(EAX_REG_16__SCAN_IN), .B1(n5413), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3972) );
  OAI21_X1 U4961 ( .B1(n5366), .B2(n3973), .A(n3972), .ZN(n3974) );
  AOI21_X1 U4962 ( .B1(n3975), .B2(n5369), .A(n3974), .ZN(n5394) );
  XNOR2_X1 U4963 ( .A(n3976), .B(n5573), .ZN(n5747) );
  AOI22_X1 U4964 ( .A1(n4108), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3005), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3980) );
  AOI22_X1 U4965 ( .A1(n3011), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3382), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3979) );
  AOI22_X1 U4966 ( .A1(n3391), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n5258), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U4967 ( .A1(n3012), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3003), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3977) );
  NAND4_X1 U4968 ( .A1(n3980), .A2(n3979), .A3(n3978), .A4(n3977), .ZN(n3987)
         );
  AOI22_X1 U4969 ( .A1(n4119), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n5349), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3984) );
  AOI22_X1 U4970 ( .A1(n5340), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n5348), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3983) );
  AOI22_X1 U4971 ( .A1(n2990), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3982) );
  AOI22_X1 U4972 ( .A1(n3004), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n5326), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3981) );
  NAND4_X1 U4973 ( .A1(n3984), .A2(n3983), .A3(n3982), .A4(n3981), .ZN(n3986)
         );
  OAI21_X1 U4974 ( .B1(n3987), .B2(n3986), .A(n3985), .ZN(n3990) );
  NAND2_X1 U4975 ( .A1(n3809), .A2(EAX_REG_15__SCAN_IN), .ZN(n3989) );
  NAND2_X1 U4976 ( .A1(n5413), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3988)
         );
  NAND3_X1 U4977 ( .A1(n3990), .A2(n3989), .A3(n3988), .ZN(n3991) );
  AOI21_X1 U4978 ( .B1(n5747), .B2(n5369), .A(n3991), .ZN(n5571) );
  XNOR2_X1 U4979 ( .A(n4024), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6003)
         );
  NAND2_X1 U4980 ( .A1(n5366), .A2(n5362), .ZN(n4077) );
  AOI22_X1 U4981 ( .A1(n3005), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3012), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3999) );
  AOI22_X1 U4982 ( .A1(n4119), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3382), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3998) );
  NAND2_X1 U4983 ( .A1(n5348), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3995) );
  NAND2_X1 U4984 ( .A1(n3004), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3994) );
  AND3_X1 U4985 ( .A1(n3995), .A2(n5362), .A3(n3994), .ZN(n3997) );
  AOI22_X1 U4986 ( .A1(n3017), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3996) );
  NAND4_X1 U4987 ( .A1(n3999), .A2(n3998), .A3(n3997), .A4(n3996), .ZN(n4005)
         );
  AOI22_X1 U4988 ( .A1(n5349), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4003) );
  AOI22_X1 U4989 ( .A1(n3011), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n5258), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4002) );
  AOI22_X1 U4990 ( .A1(n5340), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3003), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4001) );
  AOI22_X1 U4991 ( .A1(n4108), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n5326), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4000) );
  NAND4_X1 U4992 ( .A1(n4003), .A2(n4002), .A3(n4001), .A4(n4000), .ZN(n4004)
         );
  OR2_X1 U4993 ( .A1(n4005), .A2(n4004), .ZN(n4008) );
  INV_X1 U4994 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4421) );
  INV_X1 U4995 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5563) );
  OAI22_X1 U4996 ( .A1(n4006), .A2(n4421), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5563), .ZN(n4007) );
  AOI21_X1 U4997 ( .B1(n4077), .B2(n4008), .A(n4007), .ZN(n4009) );
  AOI21_X1 U4998 ( .B1(n6003), .B2(n5369), .A(n4009), .ZN(n5558) );
  AOI22_X1 U4999 ( .A1(n4108), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3005), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4013) );
  AOI22_X1 U5000 ( .A1(n5340), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4012) );
  AOI22_X1 U5001 ( .A1(n5349), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4011) );
  AOI22_X1 U5002 ( .A1(n3011), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3003), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4010) );
  NAND4_X1 U5003 ( .A1(n4013), .A2(n4012), .A3(n4011), .A4(n4010), .ZN(n4019)
         );
  AOI22_X1 U5004 ( .A1(n3329), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n2990), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4017) );
  AOI22_X1 U5005 ( .A1(n3391), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3004), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4016) );
  AOI22_X1 U5006 ( .A1(n5258), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n5326), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4015) );
  AOI22_X1 U5007 ( .A1(n5348), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3002), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4014) );
  NAND4_X1 U5008 ( .A1(n4017), .A2(n4016), .A3(n4015), .A4(n4014), .ZN(n4018)
         );
  NOR2_X1 U5009 ( .A1(n4019), .A2(n4018), .ZN(n4023) );
  NAND2_X1 U5010 ( .A1(n6498), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4020)
         );
  NAND2_X1 U5011 ( .A1(n5362), .A2(n4020), .ZN(n4021) );
  AOI21_X1 U5012 ( .B1(n3809), .B2(EAX_REG_18__SCAN_IN), .A(n4021), .ZN(n4022)
         );
  OAI21_X1 U5013 ( .B1(n5366), .B2(n4023), .A(n4022), .ZN(n4031) );
  INV_X1 U5014 ( .A(n4062), .ZN(n4029) );
  INV_X1 U5015 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4027) );
  INV_X1 U5016 ( .A(n4025), .ZN(n4026) );
  NAND2_X1 U5017 ( .A1(n4027), .A2(n4026), .ZN(n4028) );
  NAND2_X1 U5018 ( .A1(n4029), .A2(n4028), .ZN(n6071) );
  NAND2_X1 U5019 ( .A1(n4031), .A2(n4030), .ZN(n5623) );
  AOI22_X1 U5020 ( .A1(n4108), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3012), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4036) );
  AOI22_X1 U5021 ( .A1(n5340), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3008), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4035) );
  AOI22_X1 U5022 ( .A1(n4119), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3002), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4034) );
  AOI22_X1 U5023 ( .A1(n3003), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n5326), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4033) );
  NAND4_X1 U5024 ( .A1(n4036), .A2(n4035), .A3(n4034), .A4(n4033), .ZN(n4044)
         );
  AOI22_X1 U5025 ( .A1(n3190), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3329), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4042) );
  AOI22_X1 U5026 ( .A1(n5349), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3011), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4041) );
  NAND2_X1 U5027 ( .A1(n5258), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4038) );
  NAND2_X1 U5028 ( .A1(n5348), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4037) );
  AND3_X1 U5029 ( .A1(n4038), .A2(n4037), .A3(n5362), .ZN(n4040) );
  AOI22_X1 U5030 ( .A1(n2990), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3004), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4039) );
  NAND4_X1 U5031 ( .A1(n4042), .A2(n4041), .A3(n4040), .A4(n4039), .ZN(n4043)
         );
  OAI21_X1 U5032 ( .B1(n4044), .B2(n4043), .A(n4077), .ZN(n4046) );
  AOI22_X1 U5033 ( .A1(n3809), .A2(EAX_REG_19__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6498), .ZN(n4045) );
  NAND2_X1 U5034 ( .A1(n4046), .A2(n4045), .ZN(n4048) );
  INV_X1 U5035 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5738) );
  XNOR2_X1 U5036 ( .A(n4062), .B(n5738), .ZN(n5740) );
  NAND2_X1 U5037 ( .A1(n5740), .A2(n5369), .ZN(n4047) );
  NAND2_X1 U5038 ( .A1(n4048), .A2(n4047), .ZN(n5543) );
  AOI22_X1 U5039 ( .A1(n4108), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3005), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4052) );
  AOI22_X1 U5040 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4119), .B1(n5349), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4051) );
  AOI22_X1 U5041 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n3329), .B1(n3017), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4050) );
  AOI22_X1 U5042 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(n5258), .B1(n3004), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4049) );
  NAND4_X1 U5043 ( .A1(n4052), .A2(n4051), .A3(n4050), .A4(n4049), .ZN(n4058)
         );
  AOI22_X1 U5044 ( .A1(n5340), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n5348), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4056) );
  AOI22_X1 U5045 ( .A1(n3012), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n5343), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4055) );
  AOI22_X1 U5046 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n3008), .B1(n5326), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4054) );
  AOI22_X1 U5047 ( .A1(n3011), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3212), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4053) );
  NAND4_X1 U5048 ( .A1(n4056), .A2(n4055), .A3(n4054), .A4(n4053), .ZN(n4057)
         );
  NOR2_X1 U5049 ( .A1(n4058), .A2(n4057), .ZN(n4059) );
  OR2_X1 U5050 ( .A1(n5366), .A2(n4059), .ZN(n4066) );
  NAND2_X1 U5051 ( .A1(n6498), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4060)
         );
  NAND2_X1 U5052 ( .A1(n5362), .A2(n4060), .ZN(n4061) );
  AOI21_X1 U5053 ( .B1(n3809), .B2(EAX_REG_20__SCAN_IN), .A(n4061), .ZN(n4065)
         );
  OAI21_X1 U5054 ( .B1(n4063), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n4098), 
        .ZN(n5732) );
  NOR2_X1 U5055 ( .A1(n5732), .A2(n5362), .ZN(n4064) );
  AOI21_X1 U5056 ( .B1(n4066), .B2(n4065), .A(n4064), .ZN(n5533) );
  AOI22_X1 U5057 ( .A1(n3012), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3017), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4070) );
  AOI22_X1 U5058 ( .A1(n3011), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n5348), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4069) );
  AOI22_X1 U5059 ( .A1(n4108), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n5343), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4068) );
  AOI22_X1 U5060 ( .A1(n3008), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3002), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4067) );
  NAND4_X1 U5061 ( .A1(n4070), .A2(n4069), .A3(n4068), .A4(n4067), .ZN(n4079)
         );
  AOI22_X1 U5062 ( .A1(n5349), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3190), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4076) );
  NAND2_X1 U5063 ( .A1(n5340), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4072)
         );
  NAND2_X1 U5064 ( .A1(n5258), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4071) );
  AND3_X1 U5065 ( .A1(n4072), .A2(n4071), .A3(n5362), .ZN(n4075) );
  AOI22_X1 U5066 ( .A1(n4119), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3004), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4074) );
  AOI22_X1 U5067 ( .A1(n3329), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n5326), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4073) );
  NAND4_X1 U5068 ( .A1(n4076), .A2(n4075), .A3(n4074), .A4(n4073), .ZN(n4078)
         );
  OAI21_X1 U5069 ( .B1(n4079), .B2(n4078), .A(n4077), .ZN(n4081) );
  AOI22_X1 U5070 ( .A1(n3809), .A2(EAX_REG_21__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6498), .ZN(n4080) );
  NAND2_X1 U5071 ( .A1(n4081), .A2(n4080), .ZN(n4083) );
  XNOR2_X1 U5072 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .B(n4098), .ZN(n5973)
         );
  NAND2_X1 U5073 ( .A1(n5973), .A2(n5369), .ZN(n4082) );
  NAND2_X1 U5074 ( .A1(n4083), .A2(n4082), .ZN(n5608) );
  AOI22_X1 U5075 ( .A1(n5340), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3005), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4087) );
  AOI22_X1 U5076 ( .A1(n3329), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n2990), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4086) );
  AOI22_X1 U5077 ( .A1(n3008), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n5258), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4085) );
  AOI22_X1 U5078 ( .A1(n3011), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3004), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4084) );
  NAND4_X1 U5079 ( .A1(n4087), .A2(n4086), .A3(n4085), .A4(n4084), .ZN(n4093)
         );
  AOI22_X1 U5080 ( .A1(n4108), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n5348), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4091) );
  AOI22_X1 U5081 ( .A1(n4119), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3012), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4090) );
  AOI22_X1 U5082 ( .A1(n5349), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3003), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4089) );
  AOI22_X1 U5083 ( .A1(n5326), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3212), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4088) );
  NAND4_X1 U5084 ( .A1(n4091), .A2(n4090), .A3(n4089), .A4(n4088), .ZN(n4092)
         );
  NOR2_X1 U5085 ( .A1(n4093), .A2(n4092), .ZN(n4097) );
  OAI21_X1 U5086 ( .B1(PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6728), .A(n6498), 
        .ZN(n4094) );
  INV_X1 U5087 ( .A(n4094), .ZN(n4095) );
  AOI21_X1 U5088 ( .B1(n3809), .B2(EAX_REG_22__SCAN_IN), .A(n4095), .ZN(n4096)
         );
  OAI21_X1 U5089 ( .B1(n5366), .B2(n4097), .A(n4096), .ZN(n4102) );
  OAI21_X1 U5090 ( .B1(n4100), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n4145), 
        .ZN(n5964) );
  OR2_X1 U5091 ( .A1(n5964), .A2(n5362), .ZN(n4101) );
  NAND2_X1 U5092 ( .A1(n4102), .A2(n4101), .ZN(n5717) );
  AOI22_X1 U5093 ( .A1(n5340), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3005), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4107) );
  AOI22_X1 U5094 ( .A1(n4119), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3012), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4106) );
  AOI22_X1 U5095 ( .A1(n3382), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3003), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4105) );
  AOI22_X1 U5096 ( .A1(n5350), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n5326), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4104) );
  NAND4_X1 U5097 ( .A1(n4107), .A2(n4106), .A3(n4105), .A4(n4104), .ZN(n4114)
         );
  AOI22_X1 U5098 ( .A1(n4108), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n5348), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4112) );
  AOI22_X1 U5099 ( .A1(n3011), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n2990), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4111) );
  AOI22_X1 U5100 ( .A1(n3391), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n5258), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4110) );
  AOI22_X1 U5101 ( .A1(n5349), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3002), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4109) );
  NAND4_X1 U5102 ( .A1(n4112), .A2(n4111), .A3(n4110), .A4(n4109), .ZN(n4113)
         );
  NOR2_X1 U5103 ( .A1(n4114), .A2(n4113), .ZN(n4132) );
  AOI22_X1 U5104 ( .A1(n5340), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5348), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4118) );
  AOI22_X1 U5105 ( .A1(n5349), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3012), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4117) );
  AOI22_X1 U5106 ( .A1(n3011), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3017), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4116) );
  AOI22_X1 U5107 ( .A1(n5258), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n5350), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4115) );
  NAND4_X1 U5108 ( .A1(n4118), .A2(n4117), .A3(n4116), .A4(n4115), .ZN(n4125)
         );
  AOI22_X1 U5109 ( .A1(n4108), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3005), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4123) );
  AOI22_X1 U5110 ( .A1(n4119), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3003), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4122) );
  AOI22_X1 U5111 ( .A1(n3391), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n5326), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4121) );
  AOI22_X1 U5112 ( .A1(n3382), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3002), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4120) );
  NAND4_X1 U5113 ( .A1(n4123), .A2(n4122), .A3(n4121), .A4(n4120), .ZN(n4124)
         );
  NOR2_X1 U5114 ( .A1(n4125), .A2(n4124), .ZN(n4131) );
  XNOR2_X1 U5115 ( .A(n4132), .B(n4131), .ZN(n4128) );
  INV_X1 U5116 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5527) );
  AOI21_X1 U5117 ( .B1(n5527), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4126) );
  AOI21_X1 U5118 ( .B1(n3809), .B2(EAX_REG_23__SCAN_IN), .A(n4126), .ZN(n4127)
         );
  OAI21_X1 U5119 ( .B1(n5366), .B2(n4128), .A(n4127), .ZN(n4130) );
  XNOR2_X1 U5120 ( .A(n4145), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5525)
         );
  NAND2_X1 U5121 ( .A1(n5525), .A2(n5369), .ZN(n4129) );
  NAND2_X1 U5122 ( .A1(n4130), .A2(n4129), .ZN(n5237) );
  NOR2_X2 U5123 ( .A1(n5239), .A2(n5237), .ZN(n4173) );
  NOR2_X1 U5124 ( .A1(n4132), .A2(n4131), .ZN(n5266) );
  AOI22_X1 U5125 ( .A1(n4108), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3005), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4136) );
  AOI22_X1 U5126 ( .A1(n5340), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n5348), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4135) );
  AOI22_X1 U5127 ( .A1(n4119), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4134) );
  AOI22_X1 U5128 ( .A1(n5349), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3003), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4133) );
  NAND4_X1 U5129 ( .A1(n4136), .A2(n4135), .A3(n4134), .A4(n4133), .ZN(n4142)
         );
  AOI22_X1 U5130 ( .A1(n3011), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n2990), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4140) );
  AOI22_X1 U5131 ( .A1(n3391), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n5350), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4139) );
  AOI22_X1 U5132 ( .A1(n5258), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n5326), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4138) );
  AOI22_X1 U5133 ( .A1(n3382), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3002), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4137) );
  NAND4_X1 U5134 ( .A1(n4140), .A2(n4139), .A3(n4138), .A4(n4137), .ZN(n4141)
         );
  OR2_X1 U5135 ( .A1(n4142), .A2(n4141), .ZN(n5265) );
  INV_X1 U5136 ( .A(n5265), .ZN(n4143) );
  XNOR2_X1 U5137 ( .A(n5266), .B(n4143), .ZN(n4144) );
  INV_X1 U5138 ( .A(n5366), .ZN(n5333) );
  NAND2_X1 U5139 ( .A1(n4144), .A2(n5333), .ZN(n4150) );
  INV_X1 U5140 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5955) );
  XNOR2_X1 U5141 ( .A(n4200), .B(n5955), .ZN(n5959) );
  NOR2_X1 U5142 ( .A1(n5959), .A2(n5362), .ZN(n4148) );
  NOR2_X1 U5143 ( .A1(n4146), .A2(n5955), .ZN(n4147) );
  AOI211_X1 U5144 ( .C1(n5364), .C2(EAX_REG_24__SCAN_IN), .A(n4148), .B(n4147), 
        .ZN(n4149) );
  XNOR2_X2 U5145 ( .A(n4173), .B(n3076), .ZN(n5987) );
  AND2_X1 U5146 ( .A1(n6499), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4184) );
  NAND2_X1 U5147 ( .A1(n4184), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6517) );
  NAND2_X1 U5148 ( .A1(n4151), .A2(n5875), .ZN(n6610) );
  NAND2_X1 U5149 ( .A1(n6610), .A2(n6499), .ZN(n4152) );
  AND2_X2 U5150 ( .A1(n6269), .A2(n4152), .ZN(n6263) );
  NAND2_X1 U5151 ( .A1(n6499), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4154) );
  NAND2_X1 U5152 ( .A1(n6728), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4153) );
  AND2_X1 U5153 ( .A1(n4154), .A2(n4153), .ZN(n4550) );
  AND2_X1 U5154 ( .A1(n6351), .A2(REIP_REG_24__SCAN_IN), .ZN(n5408) );
  INV_X1 U5155 ( .A(n6263), .ZN(n5755) );
  NOR2_X1 U5156 ( .A1(n5755), .A2(n5955), .ZN(n4155) );
  AOI211_X1 U5157 ( .C1(n6253), .C2(n5959), .A(n5408), .B(n4155), .ZN(n4156)
         );
  INV_X1 U5158 ( .A(n4156), .ZN(n4157) );
  NOR2_X1 U5159 ( .A1(n4158), .A2(n4157), .ZN(n4159) );
  OAI21_X1 U5160 ( .B1(n5410), .B2(n6269), .A(n4159), .ZN(U2962) );
  NAND4_X1 U5161 ( .A1(n4160), .A2(n5813), .A3(n5833), .A4(n2988), .ZN(n4161)
         );
  NAND2_X1 U5162 ( .A1(n4162), .A2(n4161), .ZN(n4164) );
  INV_X1 U5163 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4163) );
  NAND2_X1 U5164 ( .A1(n4172), .A2(n6355), .ZN(n4171) );
  XOR2_X1 U5165 ( .A(n5401), .B(n5806), .Z(n5604) );
  INV_X1 U5166 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6660) );
  NOR2_X1 U5167 ( .A1(n6341), .A2(n6660), .ZN(n4176) );
  NOR2_X1 U5168 ( .A1(n4165), .A2(n4163), .ZN(n4166) );
  AOI211_X1 U5169 ( .C1(n5604), .C2(n6353), .A(n4176), .B(n4166), .ZN(n4169)
         );
  INV_X1 U5170 ( .A(n5406), .ZN(n4167) );
  NAND2_X1 U5171 ( .A1(n4167), .A2(n4163), .ZN(n4168) );
  NAND2_X1 U5172 ( .A1(n4171), .A2(n4170), .ZN(U2995) );
  NAND2_X1 U5173 ( .A1(n4172), .A2(n6276), .ZN(n4180) );
  AND2_X1 U5174 ( .A1(n5239), .A2(n5237), .ZN(n4174) );
  NOR2_X1 U5175 ( .A1(n5755), .A2(n5527), .ZN(n4175) );
  AOI211_X1 U5176 ( .C1(n6253), .C2(n5525), .A(n4176), .B(n4175), .ZN(n4177)
         );
  NAND2_X1 U5177 ( .A1(n4180), .A2(n4179), .ZN(U2963) );
  INV_X1 U5178 ( .A(n4219), .ZN(n4181) );
  NAND2_X1 U5179 ( .A1(n4220), .A2(n4181), .ZN(n4221) );
  NAND2_X1 U5180 ( .A1(n6735), .A2(n6728), .ZN(n4192) );
  INV_X1 U5181 ( .A(n4192), .ZN(n4189) );
  NAND3_X1 U5182 ( .A1(n4182), .A2(n4189), .A3(n3230), .ZN(n4183) );
  INV_X1 U5183 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6548) );
  INV_X1 U5184 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6545) );
  INV_X1 U5185 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6542) );
  NAND3_X1 U5186 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n6150) );
  NOR2_X1 U5187 ( .A1(n6542), .A2(n6150), .ZN(n5031) );
  NAND2_X1 U5188 ( .A1(REIP_REG_5__SCAN_IN), .A2(n5031), .ZN(n5020) );
  NOR2_X1 U5189 ( .A1(n6545), .A2(n5020), .ZN(n5022) );
  NAND2_X1 U5190 ( .A1(REIP_REG_7__SCAN_IN), .A2(n5022), .ZN(n5155) );
  NOR2_X1 U5191 ( .A1(n6548), .A2(n5155), .ZN(n5436) );
  NAND2_X1 U5192 ( .A1(n6193), .A2(n5436), .ZN(n6123) );
  NOR2_X1 U5193 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6613) );
  INV_X1 U5194 ( .A(n6613), .ZN(n6514) );
  NOR3_X1 U5195 ( .A1(n6499), .A2(n6592), .A3(n6514), .ZN(n6489) );
  AND2_X1 U5196 ( .A1(n4184), .A2(n5369), .ZN(n6509) );
  INV_X1 U5197 ( .A(n6509), .ZN(n4185) );
  NAND2_X1 U5198 ( .A1(n4185), .A2(n6341), .ZN(n4186) );
  OR2_X1 U5199 ( .A1(n6489), .A2(n4186), .ZN(n4187) );
  OAI22_X1 U5200 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6123), .B1(n4188), .B2(n6138), .ZN(n4211) );
  NAND2_X1 U5201 ( .A1(n6176), .A2(n6159), .ZN(n6178) );
  NAND2_X1 U5202 ( .A1(n6159), .A2(n5436), .ZN(n5154) );
  NAND2_X1 U5203 ( .A1(n6178), .A2(n5154), .ZN(n6136) );
  INV_X1 U5204 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6550) );
  INV_X1 U5205 ( .A(n6523), .ZN(n4777) );
  NAND2_X1 U5206 ( .A1(n4777), .A2(n4189), .ZN(n6496) );
  AND2_X1 U5207 ( .A1(n2989), .A2(n6496), .ZN(n5464) );
  INV_X1 U5208 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5584) );
  AND3_X1 U5209 ( .A1(n3230), .A2(n5584), .A3(n4192), .ZN(n4190) );
  NOR2_X1 U5210 ( .A1(n5464), .A2(n4190), .ZN(n4191) );
  NOR2_X4 U5211 ( .A1(n4194), .A2(n4191), .ZN(n6182) );
  NAND3_X1 U5212 ( .A1(n4233), .A2(EBX_REG_31__SCAN_IN), .A3(n4192), .ZN(n4193) );
  INV_X1 U5213 ( .A(n5131), .ZN(n6114) );
  AOI21_X1 U5214 ( .B1(n4195), .B2(n5136), .A(n6114), .ZN(n6303) );
  AOI22_X1 U5215 ( .A1(EBX_REG_9__SCAN_IN), .A2(n6182), .B1(n6122), .B2(n6303), 
        .ZN(n4209) );
  NOR2_X1 U5216 ( .A1(n4197), .A2(n4198), .ZN(n4199) );
  OR2_X1 U5217 ( .A1(n4196), .A2(n4199), .ZN(n5146) );
  INV_X1 U5218 ( .A(n5146), .ZN(n4207) );
  INV_X1 U5219 ( .A(n5301), .ZN(n4201) );
  INV_X1 U5220 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5335) );
  INV_X1 U5221 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4202) );
  INV_X1 U5222 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4203) );
  NOR2_X1 U5223 ( .A1(n5418), .A2(n6507), .ZN(n4205) );
  AOI22_X1 U5224 ( .A1(n4207), .A2(n6146), .B1(n6160), .B2(n5143), .ZN(n4208)
         );
  OAI211_X1 U5225 ( .C1(n6136), .C2(n6550), .A(n4209), .B(n4208), .ZN(n4210)
         );
  OR3_X1 U5226 ( .A1(n6351), .A2(n4211), .A3(n4210), .ZN(U2818) );
  INV_X1 U5227 ( .A(n4212), .ZN(n4214) );
  INV_X1 U5228 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n4213) );
  OR2_X1 U5229 ( .A1(n5875), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5460) );
  OAI211_X1 U5230 ( .C1(n4214), .C2(n4213), .A(n4291), .B(n5460), .ZN(U2788)
         );
  INV_X1 U5231 ( .A(n4215), .ZN(n4269) );
  NAND3_X1 U5232 ( .A1(n6483), .A2(n4269), .A3(n4263), .ZN(n4217) );
  INV_X1 U5233 ( .A(n4262), .ZN(n4270) );
  MUX2_X1 U5234 ( .A(n4217), .B(n4216), .S(n4270), .Z(n4218) );
  AOI21_X1 U5235 ( .B1(n4220), .B2(n4219), .A(n4218), .ZN(n6484) );
  NAND2_X1 U5236 ( .A1(n4221), .A2(n4269), .ZN(n4224) );
  NAND2_X1 U5237 ( .A1(n4262), .A2(n4222), .ZN(n4223) );
  NAND2_X1 U5238 ( .A1(n4224), .A2(n4223), .ZN(n6043) );
  INV_X1 U5239 ( .A(n4225), .ZN(n5119) );
  OR2_X1 U5240 ( .A1(n2989), .A2(n5119), .ZN(n5461) );
  AOI21_X1 U5241 ( .B1(n5461), .B2(n6523), .A(READY_N), .ZN(n6611) );
  NOR2_X1 U5242 ( .A1(n6043), .A2(n6611), .ZN(n6481) );
  OR2_X1 U5243 ( .A1(n6481), .A2(n6505), .ZN(n4228) );
  INV_X1 U5244 ( .A(n4228), .ZN(n6049) );
  INV_X1 U5245 ( .A(MORE_REG_SCAN_IN), .ZN(n4226) );
  OR2_X1 U5246 ( .A1(n6049), .A2(n4226), .ZN(n4227) );
  OAI21_X1 U5247 ( .B1(n6484), .B2(n4228), .A(n4227), .ZN(U3471) );
  NOR2_X1 U5248 ( .A1(n4229), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4231)
         );
  NOR2_X1 U5249 ( .A1(n4231), .A2(n4230), .ZN(n5118) );
  INV_X1 U5250 ( .A(n5118), .ZN(n4242) );
  INV_X1 U5251 ( .A(n5454), .ZN(n5641) );
  NAND3_X1 U5252 ( .A1(n5641), .A2(n4232), .A3(n3796), .ZN(n4300) );
  INV_X1 U5253 ( .A(n4300), .ZN(n4235) );
  NAND4_X1 U5254 ( .A1(n4235), .A2(n3239), .A3(n3006), .A4(n4233), .ZN(n4236)
         );
  OAI21_X1 U5255 ( .B1(n4247), .B2(n4270), .A(n4236), .ZN(n4237) );
  INV_X1 U5256 ( .A(n4238), .ZN(n4239) );
  AOI21_X1 U5257 ( .B1(n4241), .B2(n4240), .A(n4239), .ZN(n4553) );
  INV_X1 U5258 ( .A(n4553), .ZN(n5122) );
  NAND2_X2 U5259 ( .A1(n6207), .A2(n5454), .ZN(n5639) );
  OAI222_X1 U5260 ( .A1(n4242), .A2(n5637), .B1(n5116), .B2(n6207), .C1(n5122), 
        .C2(n5639), .ZN(U2859) );
  INV_X1 U5261 ( .A(n4244), .ZN(n4246) );
  AND3_X1 U5262 ( .A1(n3610), .A2(n3724), .A3(n3605), .ZN(n4245) );
  NAND2_X1 U5263 ( .A1(n4246), .A2(n4245), .ZN(n5373) );
  NAND2_X1 U5264 ( .A1(n6170), .A2(n5373), .ZN(n4254) );
  NAND2_X1 U5265 ( .A1(n4247), .A2(n4263), .ZN(n4464) );
  XNOR2_X1 U5266 ( .A(n4248), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4252)
         );
  XNOR2_X1 U5267 ( .A(n3234), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4249)
         );
  NAND2_X1 U5268 ( .A1(n4774), .A2(n4249), .ZN(n4250) );
  OAI21_X1 U5269 ( .B1(n4252), .B2(n4466), .A(n4250), .ZN(n4251) );
  AOI21_X1 U5270 ( .B1(n4464), .B2(n4252), .A(n4251), .ZN(n4253) );
  NAND2_X1 U5271 ( .A1(n4254), .A2(n4253), .ZN(n4471) );
  NOR2_X1 U5272 ( .A1(n6507), .A2(n4286), .ZN(n5380) );
  INV_X1 U5273 ( .A(n5380), .ZN(n4258) );
  AOI22_X1 U5274 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4255), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4566), .ZN(n5381) );
  NAND3_X1 U5275 ( .A1(n4248), .A2(n6497), .A3(n4256), .ZN(n4257) );
  OAI21_X1 U5276 ( .B1(n4258), .B2(n5381), .A(n4257), .ZN(n4259) );
  AOI21_X1 U5277 ( .B1(n4471), .B2(n6593), .A(n4259), .ZN(n4277) );
  INV_X1 U5278 ( .A(n4260), .ZN(n4275) );
  INV_X1 U5279 ( .A(n4261), .ZN(n4265) );
  OR2_X1 U5280 ( .A1(n4263), .A2(n4262), .ZN(n4264) );
  OAI21_X1 U5281 ( .B1(n3610), .B2(n4265), .A(n4264), .ZN(n4303) );
  INV_X1 U5282 ( .A(n4266), .ZN(n4267) );
  NOR2_X1 U5283 ( .A1(n4303), .A2(n4267), .ZN(n4274) );
  AOI21_X1 U5284 ( .B1(n4269), .B2(n6523), .A(n4268), .ZN(n4271) );
  OAI211_X1 U5285 ( .C1(n4774), .C2(n4272), .A(n4271), .B(n4270), .ZN(n4273)
         );
  NAND3_X1 U5286 ( .A1(n4275), .A2(n4274), .A3(n4273), .ZN(n6467) );
  NOR2_X1 U5287 ( .A1(n6507), .A2(n6498), .ZN(n4779) );
  NAND2_X1 U5288 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4779), .ZN(n6589) );
  INV_X1 U5289 ( .A(n6589), .ZN(n6490) );
  AOI22_X1 U5290 ( .A1(n4301), .A2(n6467), .B1(FLUSH_REG_SCAN_IN), .B2(n6490), 
        .ZN(n6042) );
  NAND2_X1 U5291 ( .A1(n6499), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6590) );
  NAND2_X1 U5292 ( .A1(n6042), .A2(n6590), .ZN(n6598) );
  NOR2_X1 U5293 ( .A1(n4248), .A2(n6594), .ZN(n5378) );
  OAI21_X1 U5294 ( .B1(n5384), .B2(n5378), .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), 
        .ZN(n4276) );
  OAI21_X1 U5295 ( .B1(n4277), .B2(n5384), .A(n4276), .ZN(U3459) );
  AOI21_X1 U5296 ( .B1(n6593), .B2(n4774), .A(n5384), .ZN(n4281) );
  NAND2_X1 U5297 ( .A1(n3808), .A2(n5373), .ZN(n6465) );
  OAI21_X1 U5298 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6463), .A(n6465), 
        .ZN(n4279) );
  OAI22_X1 U5299 ( .A1(n6507), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6594), .ZN(n4278) );
  AOI21_X1 U5300 ( .B1(n4279), .B2(n6593), .A(n4278), .ZN(n4280) );
  OAI22_X1 U5301 ( .A1(n4281), .A2(n3078), .B1(n4280), .B2(n5384), .ZN(U3461)
         );
  XNOR2_X1 U5302 ( .A(n4282), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4555)
         );
  INV_X1 U5303 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6605) );
  NOR2_X1 U5304 ( .A1(n6341), .A2(n6605), .ZN(n4552) );
  AOI21_X1 U5305 ( .B1(n4312), .B2(n5224), .A(n4286), .ZN(n4283) );
  AOI211_X1 U5306 ( .C1(n6353), .C2(n5118), .A(n4552), .B(n4283), .ZN(n4288)
         );
  NAND2_X1 U5307 ( .A1(n4285), .A2(n4284), .ZN(n5222) );
  AND2_X1 U5308 ( .A1(n5222), .A2(n4286), .ZN(n4314) );
  INV_X1 U5309 ( .A(n4314), .ZN(n4287) );
  OAI211_X1 U5310 ( .C1(n4555), .C2(n6283), .A(n4288), .B(n4287), .ZN(U3018)
         );
  INV_X1 U5311 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n4293) );
  INV_X1 U5312 ( .A(n6495), .ZN(n4289) );
  OAI21_X1 U5313 ( .B1(n4291), .B2(READY_N), .A(n4422), .ZN(n4352) );
  NAND2_X1 U5314 ( .A1(n3014), .A2(n6735), .ZN(n4290) );
  INV_X1 U5315 ( .A(DATAI_15_), .ZN(n6686) );
  INV_X1 U5316 ( .A(EAX_REG_15__SCAN_IN), .ZN(n4292) );
  OAI222_X1 U5317 ( .A1(n4293), .A2(n4352), .B1(n4353), .B2(n6686), .C1(n4292), 
        .C2(n4422), .ZN(U2954) );
  NOR2_X1 U5318 ( .A1(n4295), .A2(n4294), .ZN(n4296) );
  OR2_X1 U5319 ( .A1(n4297), .A2(n4296), .ZN(n6189) );
  XNOR2_X1 U5320 ( .A(n6196), .B(n4298), .ZN(n4311) );
  AOI22_X1 U5321 ( .A1(n6203), .A2(n4311), .B1(EBX_REG_1__SCAN_IN), .B2(n5617), 
        .ZN(n4299) );
  OAI21_X1 U5322 ( .B1(n6189), .B2(n5639), .A(n4299), .ZN(U2858) );
  NOR2_X1 U5323 ( .A1(n3724), .A2(n4300), .ZN(n4302) );
  OAI21_X1 U5324 ( .B1(n4303), .B2(n4302), .A(n4301), .ZN(n4304) );
  NAND2_X1 U5325 ( .A1(n2997), .A2(n5454), .ZN(n4305) );
  INV_X1 U5326 ( .A(n4305), .ZN(n4306) );
  INV_X1 U5327 ( .A(DATAI_1_), .ZN(n6712) );
  INV_X1 U5328 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6241) );
  OAI222_X1 U5329 ( .A1(n6189), .A2(n5983), .B1(n5039), .B2(n6712), .C1(n5640), 
        .C2(n6241), .ZN(U2890) );
  XNOR2_X1 U5330 ( .A(n4308), .B(n4307), .ZN(n5046) );
  INV_X1 U5331 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6600) );
  NOR2_X1 U5332 ( .A1(n6341), .A2(n6600), .ZN(n5041) );
  INV_X1 U5333 ( .A(n6296), .ZN(n5829) );
  AND3_X1 U5334 ( .A1(n5829), .A2(n4309), .A3(n4566), .ZN(n4310) );
  AOI211_X1 U5335 ( .C1(n6353), .C2(n4311), .A(n5041), .B(n4310), .ZN(n4316)
         );
  INV_X1 U5336 ( .A(n4312), .ZN(n4313) );
  OAI21_X1 U5337 ( .B1(n4314), .B2(n4313), .A(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .ZN(n4315) );
  OAI211_X1 U5338 ( .C1(n5046), .C2(n6283), .A(n4316), .B(n4315), .ZN(U3017)
         );
  AOI21_X1 U5339 ( .B1(n4318), .B2(n4326), .A(n4317), .ZN(n6352) );
  INV_X1 U5340 ( .A(n6352), .ZN(n6164) );
  INV_X1 U5341 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4322) );
  OR2_X1 U5342 ( .A1(n4319), .A2(n4320), .ZN(n4321) );
  NAND2_X1 U5343 ( .A1(n4321), .A2(n4446), .ZN(n6268) );
  OAI222_X1 U5344 ( .A1(n6164), .A2(n5637), .B1(n4322), .B2(n6207), .C1(n6268), 
        .C2(n5639), .ZN(U2856) );
  NOR2_X1 U5345 ( .A1(n4324), .A2(n4323), .ZN(n4325) );
  NOR2_X1 U5346 ( .A1(n4319), .A2(n4325), .ZN(n6275) );
  INV_X1 U5347 ( .A(n6275), .ZN(n4329) );
  INV_X1 U5348 ( .A(DATAI_2_), .ZN(n4430) );
  INV_X1 U5349 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6239) );
  OAI222_X1 U5350 ( .A1(n4329), .A2(n5983), .B1(n5039), .B2(n4430), .C1(n5640), 
        .C2(n6239), .ZN(U2889) );
  OAI21_X1 U5351 ( .B1(n4328), .B2(n4327), .A(n4326), .ZN(n6173) );
  INV_X1 U5352 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4330) );
  OAI222_X1 U5353 ( .A1(n6173), .A2(n5637), .B1(n6207), .B2(n4330), .C1(n4329), 
        .C2(n5639), .ZN(U2857) );
  AND2_X1 U5354 ( .A1(n4835), .A2(n4334), .ZN(n4333) );
  NAND2_X1 U5355 ( .A1(n4836), .A2(n4333), .ZN(n4345) );
  NAND2_X1 U5356 ( .A1(n5749), .A2(DATAI_16_), .ZN(n6452) );
  NAND2_X1 U5357 ( .A1(n5749), .A2(DATAI_24_), .ZN(n6461) );
  INV_X1 U5358 ( .A(n6461), .ZN(n6381) );
  INV_X1 U5359 ( .A(n4836), .ZN(n4574) );
  INV_X1 U5360 ( .A(n4334), .ZN(n4611) );
  NAND2_X1 U5361 ( .A1(n4835), .A2(n4975), .ZN(n4671) );
  NOR3_X1 U5362 ( .A1(n4574), .A2(n4611), .A3(n4671), .ZN(n4335) );
  INV_X1 U5363 ( .A(n6590), .ZN(n4336) );
  NAND2_X1 U5364 ( .A1(n4539), .A2(n3230), .ZN(n6451) );
  NAND2_X1 U5365 ( .A1(n6167), .A2(n3808), .ZN(n4746) );
  INV_X1 U5366 ( .A(n4339), .ZN(n4575) );
  NAND2_X1 U5367 ( .A1(n6170), .A2(n4339), .ZN(n4707) );
  OR2_X1 U5368 ( .A1(n4746), .A2(n4707), .ZN(n4340) );
  NAND2_X1 U5369 ( .A1(n4340), .A2(n4557), .ZN(n4346) );
  INV_X1 U5370 ( .A(n5875), .ZN(n6367) );
  NAND2_X1 U5371 ( .A1(n4346), .A2(n6367), .ZN(n4342) );
  NAND2_X1 U5372 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n4710), .ZN(n4341) );
  INV_X1 U5373 ( .A(DATAI_0_), .ZN(n6787) );
  NOR2_X1 U5374 ( .A1(n6787), .A2(n4616), .ZN(n6456) );
  INV_X1 U5375 ( .A(n6456), .ZN(n5889) );
  OAI22_X1 U5376 ( .A1(n6451), .A2(n4557), .B1(n4556), .B2(n5889), .ZN(n4344)
         );
  AOI21_X1 U5377 ( .B1(n6381), .B2(n4743), .A(n4344), .ZN(n4351) );
  AND2_X1 U5378 ( .A1(n4345), .A2(n5749), .ZN(n4348) );
  NOR2_X1 U5379 ( .A1(n5875), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6375) );
  INV_X1 U5380 ( .A(n4346), .ZN(n4347) );
  OAI21_X1 U5381 ( .B1(n4348), .B2(n6375), .A(n4347), .ZN(n4349) );
  OAI211_X1 U5382 ( .C1(n4710), .C2(n6367), .A(n4349), .B(n4879), .ZN(n4559)
         );
  NAND2_X1 U5383 ( .A1(n4559), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4350)
         );
  OAI211_X1 U5384 ( .C1(n4843), .C2(n6452), .A(n4351), .B(n4350), .ZN(U3140)
         );
  INV_X1 U5385 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4355) );
  NAND2_X1 U5386 ( .A1(n4418), .A2(UWORD_REG_10__SCAN_IN), .ZN(n4354) );
  NAND2_X1 U5387 ( .A1(n4410), .A2(DATAI_10_), .ZN(n4356) );
  OAI211_X1 U5388 ( .C1(n4422), .C2(n4355), .A(n4354), .B(n4356), .ZN(U2934)
         );
  INV_X1 U5389 ( .A(EAX_REG_10__SCAN_IN), .ZN(n4358) );
  NAND2_X1 U5390 ( .A1(n4418), .A2(LWORD_REG_10__SCAN_IN), .ZN(n4357) );
  OAI211_X1 U5391 ( .C1(n4422), .C2(n4358), .A(n4357), .B(n4356), .ZN(U2949)
         );
  INV_X1 U5392 ( .A(EAX_REG_14__SCAN_IN), .ZN(n4360) );
  NAND2_X1 U5393 ( .A1(n4418), .A2(LWORD_REG_14__SCAN_IN), .ZN(n4359) );
  NAND2_X1 U5394 ( .A1(n4410), .A2(DATAI_14_), .ZN(n4389) );
  OAI211_X1 U5395 ( .C1(n4422), .C2(n4360), .A(n4359), .B(n4389), .ZN(U2953)
         );
  INV_X1 U5396 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4362) );
  NAND2_X1 U5397 ( .A1(n4418), .A2(UWORD_REG_11__SCAN_IN), .ZN(n4361) );
  NAND2_X1 U5398 ( .A1(n4410), .A2(DATAI_11_), .ZN(n4377) );
  OAI211_X1 U5399 ( .C1(n4422), .C2(n4362), .A(n4361), .B(n4377), .ZN(U2935)
         );
  NAND2_X1 U5400 ( .A1(n4418), .A2(LWORD_REG_6__SCAN_IN), .ZN(n4363) );
  NAND2_X1 U5401 ( .A1(n4410), .A2(DATAI_6_), .ZN(n4394) );
  OAI211_X1 U5402 ( .C1(n4422), .C2(n4364), .A(n4363), .B(n4394), .ZN(U2945)
         );
  INV_X1 U5403 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4366) );
  NAND2_X1 U5404 ( .A1(n4418), .A2(UWORD_REG_9__SCAN_IN), .ZN(n4365) );
  NAND2_X1 U5405 ( .A1(n4410), .A2(DATAI_9_), .ZN(n4381) );
  OAI211_X1 U5406 ( .C1(n4422), .C2(n4366), .A(n4365), .B(n4381), .ZN(U2933)
         );
  INV_X1 U5407 ( .A(EAX_REG_4__SCAN_IN), .ZN(n4368) );
  NAND2_X1 U5408 ( .A1(n4418), .A2(LWORD_REG_4__SCAN_IN), .ZN(n4367) );
  NAND2_X1 U5409 ( .A1(n4410), .A2(DATAI_4_), .ZN(n4405) );
  OAI211_X1 U5410 ( .C1(n4422), .C2(n4368), .A(n4367), .B(n4405), .ZN(U2943)
         );
  NAND2_X1 U5411 ( .A1(n4418), .A2(LWORD_REG_5__SCAN_IN), .ZN(n4369) );
  NAND2_X1 U5412 ( .A1(n4410), .A2(DATAI_5_), .ZN(n4384) );
  OAI211_X1 U5413 ( .C1(n4422), .C2(n6234), .A(n4369), .B(n4384), .ZN(U2944)
         );
  INV_X1 U5414 ( .A(EAX_REG_8__SCAN_IN), .ZN(n4371) );
  NAND2_X1 U5415 ( .A1(n4418), .A2(LWORD_REG_8__SCAN_IN), .ZN(n4370) );
  NAND2_X1 U5416 ( .A1(n4410), .A2(DATAI_8_), .ZN(n4392) );
  OAI211_X1 U5417 ( .C1(n4422), .C2(n4371), .A(n4370), .B(n4392), .ZN(U2947)
         );
  NAND2_X1 U5418 ( .A1(n4418), .A2(LWORD_REG_1__SCAN_IN), .ZN(n4372) );
  NAND2_X1 U5419 ( .A1(n4410), .A2(DATAI_1_), .ZN(n4419) );
  OAI211_X1 U5420 ( .C1(n4422), .C2(n6241), .A(n4372), .B(n4419), .ZN(U2940)
         );
  NAND2_X1 U5421 ( .A1(n4418), .A2(LWORD_REG_0__SCAN_IN), .ZN(n4373) );
  NAND2_X1 U5422 ( .A1(n4410), .A2(DATAI_0_), .ZN(n4408) );
  OAI211_X1 U5423 ( .C1(n4422), .C2(n6246), .A(n4373), .B(n4408), .ZN(U2939)
         );
  INV_X1 U5424 ( .A(EAX_REG_13__SCAN_IN), .ZN(n4375) );
  NAND2_X1 U5425 ( .A1(n4418), .A2(LWORD_REG_13__SCAN_IN), .ZN(n4374) );
  NAND2_X1 U5426 ( .A1(n4410), .A2(DATAI_13_), .ZN(n4399) );
  OAI211_X1 U5427 ( .C1(n4422), .C2(n4375), .A(n4374), .B(n4399), .ZN(U2952)
         );
  NAND2_X1 U5428 ( .A1(n4418), .A2(LWORD_REG_12__SCAN_IN), .ZN(n4376) );
  NAND2_X1 U5429 ( .A1(n4410), .A2(DATAI_12_), .ZN(n4402) );
  OAI211_X1 U5430 ( .C1(n4422), .C2(n6226), .A(n4376), .B(n4402), .ZN(U2951)
         );
  INV_X1 U5431 ( .A(EAX_REG_11__SCAN_IN), .ZN(n4379) );
  NAND2_X1 U5432 ( .A1(n4418), .A2(LWORD_REG_11__SCAN_IN), .ZN(n4378) );
  OAI211_X1 U5433 ( .C1(n4422), .C2(n4379), .A(n4378), .B(n4377), .ZN(U2950)
         );
  NAND2_X1 U5434 ( .A1(n4418), .A2(UWORD_REG_3__SCAN_IN), .ZN(n4380) );
  NAND2_X1 U5435 ( .A1(n4410), .A2(DATAI_3_), .ZN(n4415) );
  OAI211_X1 U5436 ( .C1(n4422), .C2(n5172), .A(n4380), .B(n4415), .ZN(U2927)
         );
  INV_X1 U5437 ( .A(EAX_REG_9__SCAN_IN), .ZN(n4383) );
  NAND2_X1 U5438 ( .A1(n4418), .A2(LWORD_REG_9__SCAN_IN), .ZN(n4382) );
  OAI211_X1 U5439 ( .C1(n4422), .C2(n4383), .A(n4382), .B(n4381), .ZN(U2948)
         );
  INV_X1 U5440 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4386) );
  NAND2_X1 U5441 ( .A1(n4418), .A2(UWORD_REG_5__SCAN_IN), .ZN(n4385) );
  OAI211_X1 U5442 ( .C1(n4422), .C2(n4386), .A(n4385), .B(n4384), .ZN(U2929)
         );
  NAND2_X1 U5443 ( .A1(n4418), .A2(LWORD_REG_7__SCAN_IN), .ZN(n4387) );
  NAND2_X1 U5444 ( .A1(n4410), .A2(DATAI_7_), .ZN(n4396) );
  OAI211_X1 U5445 ( .C1(n4422), .C2(n4388), .A(n4387), .B(n4396), .ZN(U2946)
         );
  INV_X1 U5446 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4391) );
  NAND2_X1 U5447 ( .A1(n4418), .A2(UWORD_REG_14__SCAN_IN), .ZN(n4390) );
  OAI211_X1 U5448 ( .C1(n4422), .C2(n4391), .A(n4390), .B(n4389), .ZN(U2938)
         );
  NAND2_X1 U5449 ( .A1(n4418), .A2(UWORD_REG_8__SCAN_IN), .ZN(n4393) );
  OAI211_X1 U5450 ( .C1(n4422), .C2(n4784), .A(n4393), .B(n4392), .ZN(U2932)
         );
  INV_X1 U5451 ( .A(EAX_REG_22__SCAN_IN), .ZN(n5174) );
  NAND2_X1 U5452 ( .A1(n4418), .A2(UWORD_REG_6__SCAN_IN), .ZN(n4395) );
  OAI211_X1 U5453 ( .C1(n4422), .C2(n5174), .A(n4395), .B(n4394), .ZN(U2930)
         );
  INV_X1 U5454 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4398) );
  NAND2_X1 U5455 ( .A1(n4418), .A2(UWORD_REG_7__SCAN_IN), .ZN(n4397) );
  OAI211_X1 U5456 ( .C1(n4422), .C2(n4398), .A(n4397), .B(n4396), .ZN(U2931)
         );
  INV_X1 U5457 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4401) );
  NAND2_X1 U5458 ( .A1(n4418), .A2(UWORD_REG_13__SCAN_IN), .ZN(n4400) );
  OAI211_X1 U5459 ( .C1(n4422), .C2(n4401), .A(n4400), .B(n4399), .ZN(U2937)
         );
  INV_X1 U5460 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4404) );
  NAND2_X1 U5461 ( .A1(n4418), .A2(UWORD_REG_12__SCAN_IN), .ZN(n4403) );
  OAI211_X1 U5462 ( .C1(n4422), .C2(n4404), .A(n4403), .B(n4402), .ZN(U2936)
         );
  INV_X1 U5463 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4407) );
  NAND2_X1 U5464 ( .A1(n4418), .A2(UWORD_REG_4__SCAN_IN), .ZN(n4406) );
  OAI211_X1 U5465 ( .C1(n4422), .C2(n4407), .A(n4406), .B(n4405), .ZN(U2928)
         );
  NAND2_X1 U5466 ( .A1(n4418), .A2(UWORD_REG_0__SCAN_IN), .ZN(n4409) );
  OAI211_X1 U5467 ( .C1(n4422), .C2(n5169), .A(n4409), .B(n4408), .ZN(U2924)
         );
  INV_X1 U5468 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4412) );
  NAND2_X1 U5469 ( .A1(n4418), .A2(UWORD_REG_2__SCAN_IN), .ZN(n4411) );
  NAND2_X1 U5470 ( .A1(n4410), .A2(DATAI_2_), .ZN(n4413) );
  OAI211_X1 U5471 ( .C1(n4422), .C2(n4412), .A(n4411), .B(n4413), .ZN(U2926)
         );
  NAND2_X1 U5472 ( .A1(n4418), .A2(LWORD_REG_2__SCAN_IN), .ZN(n4414) );
  OAI211_X1 U5473 ( .C1(n4422), .C2(n6239), .A(n4414), .B(n4413), .ZN(U2941)
         );
  INV_X1 U5474 ( .A(EAX_REG_3__SCAN_IN), .ZN(n4417) );
  NAND2_X1 U5475 ( .A1(n4418), .A2(LWORD_REG_3__SCAN_IN), .ZN(n4416) );
  OAI211_X1 U5476 ( .C1(n4422), .C2(n4417), .A(n4416), .B(n4415), .ZN(U2942)
         );
  NAND2_X1 U5477 ( .A1(n4418), .A2(UWORD_REG_1__SCAN_IN), .ZN(n4420) );
  OAI211_X1 U5478 ( .C1(n4422), .C2(n4421), .A(n4420), .B(n4419), .ZN(U2925)
         );
  NAND2_X1 U5479 ( .A1(n4836), .A2(n4611), .ZN(n4508) );
  NAND2_X1 U5480 ( .A1(n4835), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4664) );
  NOR2_X1 U5481 ( .A1(n4508), .A2(n4664), .ZN(n5870) );
  NOR2_X1 U5482 ( .A1(n5870), .A2(n5875), .ZN(n4425) );
  OR2_X1 U5483 ( .A1(n4707), .A2(n4614), .ZN(n6374) );
  INV_X1 U5484 ( .A(n3808), .ZN(n4967) );
  OAI21_X1 U5485 ( .B1(n6374), .B2(n4967), .A(n6439), .ZN(n4423) );
  AOI22_X1 U5486 ( .A1(n4425), .A2(n4423), .B1(n6363), .B2(
        STATE2_REG_2__SCAN_IN), .ZN(n6427) );
  INV_X1 U5487 ( .A(DATAI_5_), .ZN(n6733) );
  NOR2_X1 U5488 ( .A1(n6733), .A2(n4616), .ZN(n6404) );
  INV_X1 U5489 ( .A(n4423), .ZN(n4424) );
  NAND2_X1 U5490 ( .A1(n4425), .A2(n4424), .ZN(n4426) );
  OAI211_X1 U5491 ( .C1(n6363), .C2(n6367), .A(n4426), .B(n4879), .ZN(n6444)
         );
  INV_X1 U5492 ( .A(DATAI_29_), .ZN(n6746) );
  NOR2_X1 U5493 ( .A1(n6267), .A2(n6746), .ZN(n6406) );
  INV_X1 U5494 ( .A(n6406), .ZN(n5924) );
  NOR2_X1 U5495 ( .A1(n6447), .A2(n5924), .ZN(n4428) );
  NAND2_X1 U5496 ( .A1(n4539), .A2(n3221), .ZN(n5919) );
  AND2_X1 U5497 ( .A1(n4835), .A2(n3446), .ZN(n4510) );
  INV_X1 U5498 ( .A(n4510), .ZN(n4580) );
  NAND2_X1 U5499 ( .A1(n5749), .A2(DATAI_21_), .ZN(n6409) );
  OAI22_X1 U5500 ( .A1(n5919), .A2(n6439), .B1(n6438), .B2(n6409), .ZN(n4427)
         );
  AOI211_X1 U5501 ( .C1(n6444), .C2(INSTQUEUE_REG_7__5__SCAN_IN), .A(n4428), 
        .B(n4427), .ZN(n4429) );
  OAI21_X1 U5502 ( .B1(n6427), .B2(n5918), .A(n4429), .ZN(U3081) );
  NOR2_X1 U5503 ( .A1(n4430), .A2(n4616), .ZN(n6390) );
  INV_X1 U5504 ( .A(DATAI_26_), .ZN(n6684) );
  NOR2_X1 U5505 ( .A1(n6267), .A2(n6684), .ZN(n6392) );
  INV_X1 U5506 ( .A(n6392), .ZN(n5907) );
  NOR2_X1 U5507 ( .A1(n6447), .A2(n5907), .ZN(n4433) );
  NAND2_X1 U5508 ( .A1(n4539), .A2(n4431), .ZN(n5902) );
  NAND2_X1 U5509 ( .A1(n5749), .A2(DATAI_18_), .ZN(n6395) );
  OAI22_X1 U5510 ( .A1(n5902), .A2(n6439), .B1(n6438), .B2(n6395), .ZN(n4432)
         );
  AOI211_X1 U5511 ( .C1(n6444), .C2(INSTQUEUE_REG_7__2__SCAN_IN), .A(n4433), 
        .B(n4432), .ZN(n4434) );
  OAI21_X1 U5512 ( .B1(n6427), .B2(n5901), .A(n4434), .ZN(U3078) );
  INV_X1 U5513 ( .A(DATAI_7_), .ZN(n6818) );
  NOR2_X1 U5514 ( .A1(n6818), .A2(n4616), .ZN(n6417) );
  INV_X1 U5515 ( .A(DATAI_31_), .ZN(n6745) );
  NOR2_X1 U5516 ( .A1(n6267), .A2(n6745), .ZN(n6421) );
  INV_X1 U5517 ( .A(n6421), .ZN(n5942) );
  NOR2_X1 U5518 ( .A1(n6447), .A2(n5942), .ZN(n4436) );
  NAND2_X1 U5519 ( .A1(n4539), .A2(n5454), .ZN(n5936) );
  NAND2_X1 U5520 ( .A1(n5749), .A2(DATAI_23_), .ZN(n6425) );
  OAI22_X1 U5521 ( .A1(n5936), .A2(n6439), .B1(n6438), .B2(n6425), .ZN(n4435)
         );
  AOI211_X1 U5522 ( .C1(n6444), .C2(INSTQUEUE_REG_7__7__SCAN_IN), .A(n4436), 
        .B(n4435), .ZN(n4437) );
  OAI21_X1 U5523 ( .B1(n6427), .B2(n5933), .A(n4437), .ZN(U3083) );
  INV_X1 U5524 ( .A(DATAI_6_), .ZN(n6621) );
  NOR2_X1 U5525 ( .A1(n6621), .A2(n4616), .ZN(n6410) );
  INV_X1 U5526 ( .A(DATAI_30_), .ZN(n6675) );
  NOR2_X1 U5527 ( .A1(n6267), .A2(n6675), .ZN(n6412) );
  INV_X1 U5528 ( .A(n6412), .ZN(n5931) );
  NOR2_X1 U5529 ( .A1(n6447), .A2(n5931), .ZN(n4439) );
  NAND2_X1 U5530 ( .A1(n4539), .A2(n3796), .ZN(n5926) );
  NAND2_X1 U5531 ( .A1(n5749), .A2(DATAI_22_), .ZN(n6415) );
  OAI22_X1 U5532 ( .A1(n5926), .A2(n6439), .B1(n6438), .B2(n6415), .ZN(n4438)
         );
  AOI211_X1 U5533 ( .C1(n6444), .C2(INSTQUEUE_REG_7__6__SCAN_IN), .A(n4439), 
        .B(n4438), .ZN(n4440) );
  OAI21_X1 U5534 ( .B1(n6427), .B2(n5925), .A(n4440), .ZN(U3082) );
  NOR2_X1 U5535 ( .A1(n6712), .A2(n4616), .ZN(n6384) );
  INV_X1 U5536 ( .A(DATAI_25_), .ZN(n6758) );
  NOR2_X1 U5537 ( .A1(n6267), .A2(n6758), .ZN(n6386) );
  INV_X1 U5538 ( .A(n6386), .ZN(n5900) );
  NOR2_X1 U5539 ( .A1(n6447), .A2(n5900), .ZN(n4443) );
  NAND2_X1 U5540 ( .A1(n4539), .A2(n3014), .ZN(n5895) );
  NAND2_X1 U5541 ( .A1(n5749), .A2(DATAI_17_), .ZN(n6389) );
  OAI22_X1 U5542 ( .A1(n5895), .A2(n6439), .B1(n6438), .B2(n6389), .ZN(n4442)
         );
  AOI211_X1 U5543 ( .C1(n6444), .C2(INSTQUEUE_REG_7__1__SCAN_IN), .A(n4443), 
        .B(n4442), .ZN(n4444) );
  OAI21_X1 U5544 ( .B1(n6427), .B2(n5894), .A(n4444), .ZN(U3077) );
  AOI21_X1 U5545 ( .B1(n4447), .B2(n4446), .A(n4454), .ZN(n5053) );
  INV_X1 U5546 ( .A(n5053), .ZN(n6154) );
  OR2_X1 U5547 ( .A1(n4317), .A2(n4448), .ZN(n4449) );
  NAND2_X1 U5548 ( .A1(n4456), .A2(n4449), .ZN(n6343) );
  INV_X1 U5549 ( .A(n6343), .ZN(n4450) );
  AOI22_X1 U5550 ( .A1(n6203), .A2(n4450), .B1(EBX_REG_4__SCAN_IN), .B2(n5617), 
        .ZN(n4451) );
  OAI21_X1 U5551 ( .B1(n6154), .B2(n5639), .A(n4451), .ZN(U2855) );
  OAI21_X1 U5552 ( .B1(n4454), .B2(n4453), .A(n4452), .ZN(n5059) );
  INV_X1 U5553 ( .A(n4608), .ZN(n4455) );
  AOI21_X1 U5554 ( .B1(n4457), .B2(n4456), .A(n4455), .ZN(n6332) );
  AOI22_X1 U5555 ( .A1(n6332), .A2(n6203), .B1(EBX_REG_5__SCAN_IN), .B2(n5617), 
        .ZN(n4458) );
  OAI21_X1 U5556 ( .B1(n5059), .B2(n5639), .A(n4458), .ZN(U2854) );
  INV_X1 U5557 ( .A(DATAI_4_), .ZN(n4525) );
  OAI222_X1 U5558 ( .A1(n6154), .A2(n5983), .B1(n5039), .B2(n4525), .C1(n5640), 
        .C2(n4368), .ZN(U2887) );
  INV_X1 U5559 ( .A(DATAI_3_), .ZN(n6721) );
  OAI222_X1 U5560 ( .A1(n6268), .A2(n5983), .B1(n5039), .B2(n6721), .C1(n5640), 
        .C2(n4417), .ZN(U2888) );
  INV_X1 U5561 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6246) );
  OAI222_X1 U5562 ( .A1(n5122), .A2(n5983), .B1(n5039), .B2(n6787), .C1(n5640), 
        .C2(n6246), .ZN(U2891) );
  NAND2_X1 U5563 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4460) );
  INV_X1 U5564 ( .A(n4460), .ZN(n4459) );
  MUX2_X1 U5565 ( .A(n4460), .B(n4459), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4469) );
  INV_X1 U5566 ( .A(n4774), .ZN(n6462) );
  MUX2_X1 U5567 ( .A(n4461), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4248), 
        .Z(n4462) );
  NOR2_X1 U5568 ( .A1(n4462), .A2(n4473), .ZN(n4463) );
  NAND2_X1 U5569 ( .A1(n4464), .A2(n4463), .ZN(n4468) );
  AOI21_X1 U5570 ( .B1(n4248), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3079), 
        .ZN(n4465) );
  NOR2_X1 U5571 ( .A1(n3017), .A2(n4465), .ZN(n6595) );
  OR2_X1 U5572 ( .A1(n4466), .A2(n6595), .ZN(n4467) );
  OAI211_X1 U5573 ( .C1(n4469), .C2(n6462), .A(n4468), .B(n4467), .ZN(n4470)
         );
  AOI21_X1 U5574 ( .B1(n6167), .B2(n5373), .A(n4470), .ZN(n6597) );
  MUX2_X1 U5575 ( .A(n3079), .B(n6597), .S(n6467), .Z(n6473) );
  INV_X1 U5576 ( .A(n6473), .ZN(n6479) );
  MUX2_X1 U5577 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n4471), .S(n6467), 
        .Z(n6470) );
  NAND3_X1 U5578 ( .A1(n6479), .A2(n6470), .A3(n6507), .ZN(n4475) );
  INV_X1 U5579 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6718) );
  AND2_X1 U5580 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6718), .ZN(n4472) );
  NAND2_X1 U5581 ( .A1(n4473), .A2(n4472), .ZN(n4474) );
  NAND2_X1 U5582 ( .A1(n4475), .A2(n4474), .ZN(n6487) );
  INV_X1 U5583 ( .A(n4476), .ZN(n5379) );
  INV_X1 U5584 ( .A(n4614), .ZN(n4477) );
  OR2_X1 U5585 ( .A1(n4478), .A2(n4477), .ZN(n4479) );
  XNOR2_X1 U5586 ( .A(n4479), .B(n6040), .ZN(n6152) );
  INV_X1 U5587 ( .A(n3610), .ZN(n6038) );
  NAND2_X1 U5588 ( .A1(n6038), .A2(n6507), .ZN(n4481) );
  MUX2_X1 U5589 ( .A(n6467), .B(FLUSH_REG_SCAN_IN), .S(STATE2_REG_1__SCAN_IN), 
        .Z(n4480) );
  OAI22_X1 U5590 ( .A1(n6152), .A2(n4481), .B1(n4480), .B2(n6040), .ZN(n6486)
         );
  AOI21_X1 U5591 ( .B1(n6487), .B2(n5379), .A(n6486), .ZN(n6491) );
  AND2_X1 U5592 ( .A1(n6491), .A2(n6718), .ZN(n4482) );
  OAI21_X1 U5593 ( .B1(n4482), .B2(n6589), .A(n4616), .ZN(n6362) );
  INV_X1 U5594 ( .A(n6362), .ZN(n4492) );
  INV_X1 U5595 ( .A(n4835), .ZN(n4483) );
  AOI21_X1 U5596 ( .B1(n4483), .B2(n6728), .A(n5875), .ZN(n4484) );
  NAND2_X1 U5597 ( .A1(n6592), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5872) );
  AOI22_X1 U5598 ( .A1(n4484), .A2(n4664), .B1(n4339), .B2(n5872), .ZN(n4486)
         );
  NAND2_X1 U5599 ( .A1(n4492), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4485) );
  OAI21_X1 U5600 ( .B1(n4492), .B2(n4486), .A(n4485), .ZN(U3464) );
  XNOR2_X1 U5601 ( .A(n4836), .B(n4664), .ZN(n4487) );
  AOI22_X1 U5602 ( .A1(n4487), .A2(n6367), .B1(n5872), .B2(n6170), .ZN(n4489)
         );
  NAND2_X1 U5603 ( .A1(n4492), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4488) );
  OAI21_X1 U5604 ( .B1(n4492), .B2(n4489), .A(n4488), .ZN(U3463) );
  AOI222_X1 U5605 ( .A1(n6491), .A2(n4779), .B1(n3808), .B2(n5872), .C1(n3446), 
        .C2(n6367), .ZN(n4491) );
  NAND2_X1 U5606 ( .A1(n4492), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4490) );
  OAI21_X1 U5607 ( .B1(n4492), .B2(n4491), .A(n4490), .ZN(U3465) );
  OAI22_X1 U5608 ( .A1(n5895), .A2(n4557), .B1(n4556), .B2(n5894), .ZN(n4493)
         );
  AOI21_X1 U5609 ( .B1(n6386), .B2(n4743), .A(n4493), .ZN(n4495) );
  NAND2_X1 U5610 ( .A1(n4559), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4494)
         );
  OAI211_X1 U5611 ( .C1(n4843), .C2(n6389), .A(n4495), .B(n4494), .ZN(U3141)
         );
  OAI22_X1 U5612 ( .A1(n5936), .A2(n4557), .B1(n4556), .B2(n5933), .ZN(n4496)
         );
  AOI21_X1 U5613 ( .B1(n6421), .B2(n4743), .A(n4496), .ZN(n4498) );
  NAND2_X1 U5614 ( .A1(n4559), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4497)
         );
  OAI211_X1 U5615 ( .C1(n4843), .C2(n6425), .A(n4498), .B(n4497), .ZN(U3147)
         );
  OAI22_X1 U5616 ( .A1(n5919), .A2(n4557), .B1(n4556), .B2(n5918), .ZN(n4499)
         );
  AOI21_X1 U5617 ( .B1(n6406), .B2(n4743), .A(n4499), .ZN(n4501) );
  NAND2_X1 U5618 ( .A1(n4559), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4500)
         );
  OAI211_X1 U5619 ( .C1(n4843), .C2(n6409), .A(n4501), .B(n4500), .ZN(U3145)
         );
  OAI22_X1 U5620 ( .A1(n5926), .A2(n4557), .B1(n4556), .B2(n5925), .ZN(n4502)
         );
  AOI21_X1 U5621 ( .B1(n6412), .B2(n4743), .A(n4502), .ZN(n4504) );
  NAND2_X1 U5622 ( .A1(n4559), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4503)
         );
  OAI211_X1 U5623 ( .C1(n4843), .C2(n6415), .A(n4504), .B(n4503), .ZN(U3146)
         );
  OAI22_X1 U5624 ( .A1(n5902), .A2(n4557), .B1(n4556), .B2(n5901), .ZN(n4505)
         );
  AOI21_X1 U5625 ( .B1(n6392), .B2(n4743), .A(n4505), .ZN(n4507) );
  NAND2_X1 U5626 ( .A1(n4559), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4506)
         );
  OAI211_X1 U5627 ( .C1(n4843), .C2(n6395), .A(n4507), .B(n4506), .ZN(U3142)
         );
  INV_X1 U5628 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6234) );
  OAI222_X1 U5629 ( .A1(n5059), .A2(n5983), .B1(n5039), .B2(n6733), .C1(n5640), 
        .C2(n6234), .ZN(U2886) );
  INV_X1 U5630 ( .A(n4976), .ZN(n4509) );
  OAI21_X1 U5631 ( .B1(n4976), .B2(n6728), .A(n6367), .ZN(n4974) );
  INV_X1 U5632 ( .A(n3820), .ZN(n5876) );
  NAND3_X1 U5633 ( .A1(n5876), .A2(n4574), .A3(n4510), .ZN(n4699) );
  NAND2_X1 U5634 ( .A1(n6170), .A2(n4575), .ZN(n4513) );
  OR2_X1 U5635 ( .A1(n4513), .A2(n4614), .ZN(n4968) );
  OAI21_X1 U5636 ( .B1(n4699), .B2(n6375), .A(n4968), .ZN(n4512) );
  NAND2_X1 U5637 ( .A1(n4838), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4748) );
  OR2_X1 U5638 ( .A1(n4748), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4972)
         );
  OR2_X1 U5639 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4972), .ZN(n4541)
         );
  NOR2_X1 U5640 ( .A1(n4514), .A2(n6498), .ZN(n5887) );
  NOR2_X1 U5641 ( .A1(n4715), .A2(n4615), .ZN(n4845) );
  INV_X1 U5642 ( .A(n4616), .ZN(n4709) );
  OAI21_X1 U5643 ( .B1(n4845), .B2(n6498), .A(n4709), .ZN(n4839) );
  AOI211_X1 U5644 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4541), .A(n5887), .B(
        n4839), .ZN(n4511) );
  NAND2_X1 U5645 ( .A1(n4538), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4517) );
  INV_X1 U5646 ( .A(n4513), .ZN(n4747) );
  AND2_X1 U5647 ( .A1(n4747), .A2(n6367), .ZN(n4620) );
  AND2_X1 U5648 ( .A1(n4514), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5078) );
  AOI22_X1 U5649 ( .A1(n4620), .A2(n6368), .B1(n5078), .B2(n4845), .ZN(n4540)
         );
  OAI22_X1 U5650 ( .A1(n5936), .A2(n4541), .B1(n4540), .B2(n5933), .ZN(n4515)
         );
  AOI21_X1 U5651 ( .B1(n6421), .B2(n4543), .A(n4515), .ZN(n4516) );
  OAI211_X1 U5652 ( .C1(n5007), .C2(n6425), .A(n4517), .B(n4516), .ZN(U3059)
         );
  NAND2_X1 U5653 ( .A1(n4538), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4520) );
  OAI22_X1 U5654 ( .A1(n5926), .A2(n4541), .B1(n4540), .B2(n5925), .ZN(n4518)
         );
  AOI21_X1 U5655 ( .B1(n6412), .B2(n4543), .A(n4518), .ZN(n4519) );
  OAI211_X1 U5656 ( .C1(n5007), .C2(n6415), .A(n4520), .B(n4519), .ZN(U3058)
         );
  NAND2_X1 U5657 ( .A1(n4538), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4523) );
  OAI22_X1 U5658 ( .A1(n5919), .A2(n4541), .B1(n4540), .B2(n5918), .ZN(n4521)
         );
  AOI21_X1 U5659 ( .B1(n6406), .B2(n4543), .A(n4521), .ZN(n4522) );
  OAI211_X1 U5660 ( .C1(n5007), .C2(n6409), .A(n4523), .B(n4522), .ZN(U3057)
         );
  NAND2_X1 U5661 ( .A1(n5749), .A2(DATAI_20_), .ZN(n6437) );
  NAND2_X1 U5662 ( .A1(n4538), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4528) );
  NAND2_X1 U5663 ( .A1(n5749), .A2(DATAI_28_), .ZN(n6448) );
  INV_X1 U5664 ( .A(n6448), .ZN(n6401) );
  NAND2_X1 U5665 ( .A1(n4539), .A2(n4524), .ZN(n6440) );
  NOR2_X1 U5666 ( .A1(n4525), .A2(n4616), .ZN(n6443) );
  OAI22_X1 U5667 ( .A1(n6440), .A2(n4541), .B1(n4540), .B2(n5913), .ZN(n4526)
         );
  AOI21_X1 U5668 ( .B1(n6401), .B2(n4543), .A(n4526), .ZN(n4527) );
  OAI211_X1 U5669 ( .C1(n5007), .C2(n6437), .A(n4528), .B(n4527), .ZN(U3056)
         );
  NAND2_X1 U5670 ( .A1(n4538), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4531) );
  OAI22_X1 U5671 ( .A1(n5902), .A2(n4541), .B1(n4540), .B2(n5901), .ZN(n4529)
         );
  AOI21_X1 U5672 ( .B1(n6392), .B2(n4543), .A(n4529), .ZN(n4530) );
  OAI211_X1 U5673 ( .C1(n5007), .C2(n6395), .A(n4531), .B(n4530), .ZN(U3054)
         );
  NAND2_X1 U5674 ( .A1(n4538), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4534) );
  OAI22_X1 U5675 ( .A1(n5895), .A2(n4541), .B1(n4540), .B2(n5894), .ZN(n4532)
         );
  AOI21_X1 U5676 ( .B1(n6386), .B2(n4543), .A(n4532), .ZN(n4533) );
  OAI211_X1 U5677 ( .C1(n5007), .C2(n6389), .A(n4534), .B(n4533), .ZN(U3053)
         );
  NAND2_X1 U5678 ( .A1(n4538), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4537) );
  OAI22_X1 U5679 ( .A1(n6451), .A2(n4541), .B1(n4540), .B2(n5889), .ZN(n4535)
         );
  AOI21_X1 U5680 ( .B1(n6381), .B2(n4543), .A(n4535), .ZN(n4536) );
  OAI211_X1 U5681 ( .C1(n5007), .C2(n6452), .A(n4537), .B(n4536), .ZN(U3052)
         );
  NAND2_X1 U5682 ( .A1(n5749), .A2(DATAI_19_), .ZN(n6430) );
  NAND2_X1 U5683 ( .A1(n4538), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4545) );
  NAND2_X1 U5684 ( .A1(n5749), .A2(DATAI_27_), .ZN(n6436) );
  INV_X1 U5685 ( .A(n6436), .ZN(n6397) );
  NAND2_X1 U5686 ( .A1(n4539), .A2(n3238), .ZN(n6431) );
  NOR2_X1 U5687 ( .A1(n6721), .A2(n4616), .ZN(n6433) );
  OAI22_X1 U5688 ( .A1(n6431), .A2(n4541), .B1(n4540), .B2(n5908), .ZN(n4542)
         );
  AOI21_X1 U5689 ( .B1(n6397), .B2(n4543), .A(n4542), .ZN(n4544) );
  OAI211_X1 U5690 ( .C1(n5007), .C2(n6430), .A(n4545), .B(n4544), .ZN(U3055)
         );
  OAI22_X1 U5691 ( .A1(n6440), .A2(n4557), .B1(n4556), .B2(n5913), .ZN(n4546)
         );
  AOI21_X1 U5692 ( .B1(n6401), .B2(n4743), .A(n4546), .ZN(n4548) );
  NAND2_X1 U5693 ( .A1(n4559), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4547)
         );
  OAI211_X1 U5694 ( .C1(n4843), .C2(n6437), .A(n4548), .B(n4547), .ZN(U3144)
         );
  INV_X1 U5695 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n4549) );
  AOI21_X1 U5696 ( .B1(n5755), .B2(n4550), .A(n4549), .ZN(n4551) );
  AOI211_X1 U5697 ( .C1(n4553), .C2(n5749), .A(n4552), .B(n4551), .ZN(n4554)
         );
  OAI21_X1 U5698 ( .B1(n4555), .B2(n6269), .A(n4554), .ZN(U2986) );
  OAI22_X1 U5699 ( .A1(n6431), .A2(n4557), .B1(n4556), .B2(n5908), .ZN(n4558)
         );
  AOI21_X1 U5700 ( .B1(n6397), .B2(n4743), .A(n4558), .ZN(n4561) );
  NAND2_X1 U5701 ( .A1(n4559), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4560)
         );
  OAI211_X1 U5702 ( .C1(n4843), .C2(n6430), .A(n4561), .B(n4560), .ZN(U3143)
         );
  XNOR2_X1 U5703 ( .A(n4562), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4564)
         );
  XNOR2_X1 U5704 ( .A(n4564), .B(n4563), .ZN(n6274) );
  INV_X1 U5705 ( .A(REIP_REG_2__SCAN_IN), .ZN(n4565) );
  OAI22_X1 U5706 ( .A1(n6342), .A2(n6173), .B1(n6341), .B2(n4565), .ZN(n4572)
         );
  NOR2_X1 U5707 ( .A1(n4566), .A2(n6327), .ZN(n4570) );
  NOR2_X1 U5708 ( .A1(n3458), .A2(n4566), .ZN(n4655) );
  OAI21_X1 U5709 ( .B1(n5200), .B2(n4655), .A(n5196), .ZN(n6338) );
  AOI21_X1 U5710 ( .B1(n6339), .B2(n4567), .A(n6338), .ZN(n4568) );
  INV_X1 U5711 ( .A(n4568), .ZN(n4569) );
  MUX2_X1 U5712 ( .A(n4570), .B(n4569), .S(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .Z(n4571) );
  AOI211_X1 U5713 ( .C1(n6339), .C2(n6346), .A(n4572), .B(n4571), .ZN(n4573)
         );
  OAI21_X1 U5714 ( .B1(n6283), .B2(n6274), .A(n4573), .ZN(U3016) );
  OAI21_X1 U5715 ( .B1(n4809), .B2(n4664), .A(n6367), .ZN(n4579) );
  NOR2_X1 U5716 ( .A1(n6170), .A2(n4575), .ZN(n4666) );
  NOR2_X1 U5717 ( .A1(n4667), .A2(n6478), .ZN(n6449) );
  AOI21_X1 U5718 ( .B1(n5079), .B2(n3808), .A(n6449), .ZN(n4576) );
  NAND3_X1 U5719 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6471), .ZN(n5080) );
  OAI22_X1 U5720 ( .A1(n4579), .A2(n4576), .B1(n5080), .B2(n6498), .ZN(n6455)
         );
  INV_X1 U5721 ( .A(n4576), .ZN(n4578) );
  INV_X1 U5722 ( .A(n4879), .ZN(n4970) );
  AOI21_X1 U5723 ( .B1(n5875), .B2(n5080), .A(n4970), .ZN(n4577) );
  OAI21_X1 U5724 ( .B1(n4579), .B2(n4578), .A(n4577), .ZN(n6457) );
  INV_X1 U5725 ( .A(n6453), .ZN(n4599) );
  INV_X1 U5726 ( .A(n6437), .ZN(n5915) );
  INV_X1 U5727 ( .A(n6440), .ZN(n6400) );
  AOI22_X1 U5728 ( .A1(n4599), .A2(n5915), .B1(n6400), .B2(n6449), .ZN(n4581)
         );
  OAI21_X1 U5729 ( .B1(n6460), .B2(n6448), .A(n4581), .ZN(n4582) );
  AOI21_X1 U5730 ( .B1(INSTQUEUE_REG_11__4__SCAN_IN), .B2(n6457), .A(n4582), 
        .ZN(n4583) );
  OAI21_X1 U5731 ( .B1(n4603), .B2(n5913), .A(n4583), .ZN(U3112) );
  INV_X1 U5732 ( .A(n6425), .ZN(n5939) );
  INV_X1 U5733 ( .A(n5936), .ZN(n6419) );
  AOI22_X1 U5734 ( .A1(n4599), .A2(n5939), .B1(n6419), .B2(n6449), .ZN(n4584)
         );
  OAI21_X1 U5735 ( .B1(n6460), .B2(n5942), .A(n4584), .ZN(n4585) );
  AOI21_X1 U5736 ( .B1(INSTQUEUE_REG_11__7__SCAN_IN), .B2(n6457), .A(n4585), 
        .ZN(n4586) );
  OAI21_X1 U5737 ( .B1(n4603), .B2(n5933), .A(n4586), .ZN(U3115) );
  INV_X1 U5738 ( .A(n6415), .ZN(n5928) );
  INV_X1 U5739 ( .A(n5926), .ZN(n6411) );
  AOI22_X1 U5740 ( .A1(n4599), .A2(n5928), .B1(n6411), .B2(n6449), .ZN(n4587)
         );
  OAI21_X1 U5741 ( .B1(n6460), .B2(n5931), .A(n4587), .ZN(n4588) );
  AOI21_X1 U5742 ( .B1(INSTQUEUE_REG_11__6__SCAN_IN), .B2(n6457), .A(n4588), 
        .ZN(n4589) );
  OAI21_X1 U5743 ( .B1(n4603), .B2(n5925), .A(n4589), .ZN(U3114) );
  INV_X1 U5744 ( .A(n6409), .ZN(n5921) );
  INV_X1 U5745 ( .A(n5919), .ZN(n6405) );
  AOI22_X1 U5746 ( .A1(n4599), .A2(n5921), .B1(n6405), .B2(n6449), .ZN(n4590)
         );
  OAI21_X1 U5747 ( .B1(n6460), .B2(n5924), .A(n4590), .ZN(n4591) );
  AOI21_X1 U5748 ( .B1(INSTQUEUE_REG_11__5__SCAN_IN), .B2(n6457), .A(n4591), 
        .ZN(n4592) );
  OAI21_X1 U5749 ( .B1(n4603), .B2(n5918), .A(n4592), .ZN(U3113) );
  INV_X1 U5750 ( .A(n6389), .ZN(n5897) );
  INV_X1 U5751 ( .A(n5895), .ZN(n6385) );
  AOI22_X1 U5752 ( .A1(n4599), .A2(n5897), .B1(n6385), .B2(n6449), .ZN(n4593)
         );
  OAI21_X1 U5753 ( .B1(n6460), .B2(n5900), .A(n4593), .ZN(n4594) );
  AOI21_X1 U5754 ( .B1(INSTQUEUE_REG_11__1__SCAN_IN), .B2(n6457), .A(n4594), 
        .ZN(n4595) );
  OAI21_X1 U5755 ( .B1(n4603), .B2(n5894), .A(n4595), .ZN(U3109) );
  INV_X1 U5756 ( .A(n6430), .ZN(n5910) );
  INV_X1 U5757 ( .A(n6431), .ZN(n6396) );
  AOI22_X1 U5758 ( .A1(n4599), .A2(n5910), .B1(n6396), .B2(n6449), .ZN(n4596)
         );
  OAI21_X1 U5759 ( .B1(n6460), .B2(n6436), .A(n4596), .ZN(n4597) );
  AOI21_X1 U5760 ( .B1(INSTQUEUE_REG_11__3__SCAN_IN), .B2(n6457), .A(n4597), 
        .ZN(n4598) );
  OAI21_X1 U5761 ( .B1(n4603), .B2(n5908), .A(n4598), .ZN(U3111) );
  INV_X1 U5762 ( .A(n6395), .ZN(n5904) );
  INV_X1 U5763 ( .A(n5902), .ZN(n6391) );
  AOI22_X1 U5764 ( .A1(n4599), .A2(n5904), .B1(n6391), .B2(n6449), .ZN(n4600)
         );
  OAI21_X1 U5765 ( .B1(n6460), .B2(n5907), .A(n4600), .ZN(n4601) );
  AOI21_X1 U5766 ( .B1(INSTQUEUE_REG_11__2__SCAN_IN), .B2(n6457), .A(n4601), 
        .ZN(n4602) );
  OAI21_X1 U5767 ( .B1(n4603), .B2(n5901), .A(n4602), .ZN(U3110) );
  INV_X1 U5768 ( .A(n4604), .ZN(n5013) );
  NAND2_X1 U5769 ( .A1(n4452), .A2(n4605), .ZN(n4606) );
  AND2_X1 U5770 ( .A1(n5013), .A2(n4606), .ZN(n6258) );
  INV_X1 U5771 ( .A(n6258), .ZN(n4663) );
  NAND2_X1 U5772 ( .A1(n4608), .A2(n4607), .ZN(n4609) );
  NAND2_X1 U5773 ( .A1(n5015), .A2(n4609), .ZN(n6139) );
  INV_X1 U5774 ( .A(n6139), .ZN(n4660) );
  AOI22_X1 U5775 ( .A1(n4660), .A2(n6203), .B1(EBX_REG_6__SCAN_IN), .B2(n5617), 
        .ZN(n4610) );
  OAI21_X1 U5776 ( .B1(n4663), .B2(n5639), .A(n4610), .ZN(U2853) );
  NOR2_X1 U5777 ( .A1(n4835), .A2(n4611), .ZN(n4612) );
  NAND2_X1 U5778 ( .A1(n4705), .A2(n4975), .ZN(n4800) );
  AOI21_X1 U5779 ( .B1(n6453), .B2(n4800), .A(n6728), .ZN(n4613) );
  AOI211_X1 U5780 ( .C1(n4747), .C2(n4614), .A(n5875), .B(n4613), .ZN(n4618)
         );
  NOR2_X1 U5781 ( .A1(n6478), .A2(n4748), .ZN(n4754) );
  AND2_X1 U5782 ( .A1(n6364), .A2(n4754), .ZN(n4619) );
  INV_X1 U5783 ( .A(n5887), .ZN(n4928) );
  INV_X1 U5784 ( .A(n4715), .ZN(n5886) );
  NAND2_X1 U5785 ( .A1(n5886), .A2(n4615), .ZN(n4927) );
  AOI21_X1 U5786 ( .B1(n4927), .B2(STATE2_REG_2__SCAN_IN), .A(n4616), .ZN(
        n4924) );
  OAI211_X1 U5787 ( .C1(n6592), .C2(n4619), .A(n4928), .B(n4924), .ZN(n4617)
         );
  NAND2_X1 U5788 ( .A1(n4645), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4626)
         );
  INV_X1 U5789 ( .A(n4619), .ZN(n4647) );
  NAND2_X1 U5790 ( .A1(n4620), .A2(n6167), .ZN(n4623) );
  INV_X1 U5791 ( .A(n4927), .ZN(n4621) );
  NAND2_X1 U5792 ( .A1(n4621), .A2(n5078), .ZN(n4622) );
  OAI22_X1 U5793 ( .A1(n6440), .A2(n4647), .B1(n4646), .B2(n5913), .ZN(n4624)
         );
  AOI21_X1 U5794 ( .B1(n5915), .B2(n4649), .A(n4624), .ZN(n4625) );
  OAI211_X1 U5795 ( .C1(n6453), .C2(n6448), .A(n4626), .B(n4625), .ZN(U3120)
         );
  NAND2_X1 U5796 ( .A1(n4645), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4629)
         );
  OAI22_X1 U5797 ( .A1(n5895), .A2(n4647), .B1(n4646), .B2(n5894), .ZN(n4627)
         );
  AOI21_X1 U5798 ( .B1(n5897), .B2(n4649), .A(n4627), .ZN(n4628) );
  OAI211_X1 U5799 ( .C1(n6453), .C2(n5900), .A(n4629), .B(n4628), .ZN(U3117)
         );
  NAND2_X1 U5800 ( .A1(n4645), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4632)
         );
  OAI22_X1 U5801 ( .A1(n5926), .A2(n4647), .B1(n4646), .B2(n5925), .ZN(n4630)
         );
  AOI21_X1 U5802 ( .B1(n5928), .B2(n4649), .A(n4630), .ZN(n4631) );
  OAI211_X1 U5803 ( .C1(n6453), .C2(n5931), .A(n4632), .B(n4631), .ZN(U3122)
         );
  NAND2_X1 U5804 ( .A1(n4645), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4635)
         );
  OAI22_X1 U5805 ( .A1(n5902), .A2(n4647), .B1(n4646), .B2(n5901), .ZN(n4633)
         );
  AOI21_X1 U5806 ( .B1(n5904), .B2(n4649), .A(n4633), .ZN(n4634) );
  OAI211_X1 U5807 ( .C1(n6453), .C2(n5907), .A(n4635), .B(n4634), .ZN(U3118)
         );
  NAND2_X1 U5808 ( .A1(n4645), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4638)
         );
  OAI22_X1 U5809 ( .A1(n5936), .A2(n4647), .B1(n4646), .B2(n5933), .ZN(n4636)
         );
  AOI21_X1 U5810 ( .B1(n5939), .B2(n4649), .A(n4636), .ZN(n4637) );
  OAI211_X1 U5811 ( .C1(n6453), .C2(n5942), .A(n4638), .B(n4637), .ZN(U3123)
         );
  NAND2_X1 U5812 ( .A1(n4645), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4641)
         );
  INV_X1 U5813 ( .A(n6452), .ZN(n5891) );
  OAI22_X1 U5814 ( .A1(n6451), .A2(n4647), .B1(n4646), .B2(n5889), .ZN(n4639)
         );
  AOI21_X1 U5815 ( .B1(n5891), .B2(n4649), .A(n4639), .ZN(n4640) );
  OAI211_X1 U5816 ( .C1(n6453), .C2(n6461), .A(n4641), .B(n4640), .ZN(U3116)
         );
  NAND2_X1 U5817 ( .A1(n4645), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4644)
         );
  OAI22_X1 U5818 ( .A1(n6431), .A2(n4647), .B1(n4646), .B2(n5908), .ZN(n4642)
         );
  AOI21_X1 U5819 ( .B1(n5910), .B2(n4649), .A(n4642), .ZN(n4643) );
  OAI211_X1 U5820 ( .C1(n6453), .C2(n6436), .A(n4644), .B(n4643), .ZN(U3119)
         );
  NAND2_X1 U5821 ( .A1(n4645), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4651)
         );
  OAI22_X1 U5822 ( .A1(n5919), .A2(n4647), .B1(n4646), .B2(n5918), .ZN(n4648)
         );
  AOI21_X1 U5823 ( .B1(n5921), .B2(n4649), .A(n4648), .ZN(n4650) );
  OAI211_X1 U5824 ( .C1(n6453), .C2(n5924), .A(n4651), .B(n4650), .ZN(U3121)
         );
  OAI21_X1 U5825 ( .B1(n4652), .B2(n4653), .A(n4654), .ZN(n6257) );
  OAI21_X1 U5826 ( .B1(n6339), .B2(n4655), .A(n5827), .ZN(n6345) );
  NAND2_X1 U5827 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6330), .ZN(n4656)
         );
  NOR2_X1 U5828 ( .A1(n6345), .A2(n4656), .ZN(n4658) );
  AOI21_X1 U5829 ( .B1(n5829), .B2(n4656), .A(n6338), .ZN(n6337) );
  INV_X1 U5830 ( .A(n6337), .ZN(n4657) );
  MUX2_X1 U5831 ( .A(n4658), .B(n4657), .S(INSTADDRPOINTER_REG_6__SCAN_IN), 
        .Z(n4659) );
  INV_X1 U5832 ( .A(n4659), .ZN(n4662) );
  AOI22_X1 U5833 ( .A1(n4660), .A2(n6353), .B1(n6351), .B2(REIP_REG_6__SCAN_IN), .ZN(n4661) );
  OAI211_X1 U5834 ( .C1(n6257), .C2(n6283), .A(n4662), .B(n4661), .ZN(U3012)
         );
  OAI222_X1 U5835 ( .A1(n4663), .A2(n5983), .B1(n5039), .B2(n6621), .C1(n5640), 
        .C2(n4364), .ZN(U2885) );
  NAND2_X1 U5836 ( .A1(n4705), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4751) );
  NAND2_X1 U5837 ( .A1(n4751), .A2(n4809), .ZN(n5871) );
  NOR3_X1 U5838 ( .A1(n5871), .A2(n4836), .A3(n4664), .ZN(n4665) );
  NOR2_X1 U5839 ( .A1(n4665), .A2(n5875), .ZN(n4674) );
  NAND2_X1 U5840 ( .A1(n5888), .A2(n3808), .ZN(n4669) );
  INV_X1 U5841 ( .A(n4667), .ZN(n4668) );
  NAND2_X1 U5842 ( .A1(n4668), .A2(n6478), .ZN(n4698) );
  NAND2_X1 U5843 ( .A1(n4669), .A2(n4698), .ZN(n4676) );
  NAND3_X1 U5844 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6478), .A3(n6471), .ZN(n5878) );
  INV_X1 U5845 ( .A(n5878), .ZN(n4670) );
  AOI22_X1 U5846 ( .A1(n4674), .A2(n4676), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4670), .ZN(n4704) );
  OR2_X1 U5847 ( .A1(n4836), .A2(n4671), .ZN(n4672) );
  OAI22_X1 U5848 ( .A1(n4699), .A2(n6409), .B1(n5919), .B2(n4698), .ZN(n4673)
         );
  AOI21_X1 U5849 ( .B1(n6406), .B2(n2986), .A(n4673), .ZN(n4679) );
  INV_X1 U5850 ( .A(n4674), .ZN(n4677) );
  AOI21_X1 U5851 ( .B1(n5875), .B2(n5878), .A(n4970), .ZN(n4675) );
  NAND2_X1 U5852 ( .A1(n4701), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4678) );
  OAI211_X1 U5853 ( .C1(n4704), .C2(n5918), .A(n4679), .B(n4678), .ZN(U3049)
         );
  OAI22_X1 U5854 ( .A1(n4699), .A2(n6425), .B1(n5936), .B2(n4698), .ZN(n4680)
         );
  AOI21_X1 U5855 ( .B1(n6421), .B2(n2986), .A(n4680), .ZN(n4682) );
  NAND2_X1 U5856 ( .A1(n4701), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4681) );
  OAI211_X1 U5857 ( .C1(n4704), .C2(n5933), .A(n4682), .B(n4681), .ZN(U3051)
         );
  OAI22_X1 U5858 ( .A1(n4699), .A2(n6415), .B1(n5926), .B2(n4698), .ZN(n4683)
         );
  AOI21_X1 U5859 ( .B1(n6412), .B2(n2986), .A(n4683), .ZN(n4685) );
  NAND2_X1 U5860 ( .A1(n4701), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4684) );
  OAI211_X1 U5861 ( .C1(n4704), .C2(n5925), .A(n4685), .B(n4684), .ZN(U3050)
         );
  OAI22_X1 U5862 ( .A1(n4699), .A2(n6452), .B1(n6451), .B2(n4698), .ZN(n4686)
         );
  AOI21_X1 U5863 ( .B1(n6381), .B2(n2986), .A(n4686), .ZN(n4688) );
  NAND2_X1 U5864 ( .A1(n4701), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4687) );
  OAI211_X1 U5865 ( .C1(n4704), .C2(n5889), .A(n4688), .B(n4687), .ZN(U3044)
         );
  OAI22_X1 U5866 ( .A1(n4699), .A2(n6389), .B1(n5895), .B2(n4698), .ZN(n4689)
         );
  AOI21_X1 U5867 ( .B1(n6386), .B2(n2986), .A(n4689), .ZN(n4691) );
  NAND2_X1 U5868 ( .A1(n4701), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4690) );
  OAI211_X1 U5869 ( .C1(n4704), .C2(n5894), .A(n4691), .B(n4690), .ZN(U3045)
         );
  OAI22_X1 U5870 ( .A1(n4699), .A2(n6430), .B1(n6431), .B2(n4698), .ZN(n4692)
         );
  AOI21_X1 U5871 ( .B1(n6397), .B2(n2986), .A(n4692), .ZN(n4694) );
  NAND2_X1 U5872 ( .A1(n4701), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4693) );
  OAI211_X1 U5873 ( .C1(n4704), .C2(n5908), .A(n4694), .B(n4693), .ZN(U3047)
         );
  OAI22_X1 U5874 ( .A1(n4699), .A2(n6437), .B1(n6440), .B2(n4698), .ZN(n4695)
         );
  AOI21_X1 U5875 ( .B1(n6401), .B2(n2986), .A(n4695), .ZN(n4697) );
  NAND2_X1 U5876 ( .A1(n4701), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4696) );
  OAI211_X1 U5877 ( .C1(n4704), .C2(n5913), .A(n4697), .B(n4696), .ZN(U3048)
         );
  OAI22_X1 U5878 ( .A1(n4699), .A2(n6395), .B1(n5902), .B2(n4698), .ZN(n4700)
         );
  AOI21_X1 U5879 ( .B1(n6392), .B2(n2986), .A(n4700), .ZN(n4703) );
  NAND2_X1 U5880 ( .A1(n4701), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4702) );
  OAI211_X1 U5881 ( .C1(n4704), .C2(n5901), .A(n4703), .B(n4702), .ZN(U3046)
         );
  NOR3_X1 U5882 ( .A1(n4743), .A2(n4706), .A3(n5875), .ZN(n4708) );
  INV_X1 U5883 ( .A(n4707), .ZN(n6366) );
  NAND2_X1 U5884 ( .A1(n6366), .A2(n6167), .ZN(n4714) );
  OAI21_X1 U5885 ( .B1(n4708), .B2(n6375), .A(n4714), .ZN(n4713) );
  OAI21_X1 U5886 ( .B1(n4715), .B2(n6498), .A(n4709), .ZN(n5077) );
  NOR2_X1 U5887 ( .A1(n5887), .A2(n5077), .ZN(n6379) );
  INV_X1 U5888 ( .A(n4710), .ZN(n4711) );
  OR2_X1 U5889 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4711), .ZN(n4741)
         );
  AOI21_X1 U5890 ( .B1(n4741), .B2(STATE2_REG_3__SCAN_IN), .A(n6478), .ZN(
        n4712) );
  NAND3_X1 U5891 ( .A1(n4713), .A2(n6379), .A3(n4712), .ZN(n4739) );
  NAND2_X1 U5892 ( .A1(n4739), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4720)
         );
  OR2_X1 U5893 ( .A1(n4714), .A2(n5875), .ZN(n4717) );
  AND2_X1 U5894 ( .A1(n4715), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5076)
         );
  NAND2_X1 U5895 ( .A1(n5078), .A2(n5076), .ZN(n4716) );
  OAI22_X1 U5896 ( .A1(n6440), .A2(n4741), .B1(n4740), .B2(n5913), .ZN(n4718)
         );
  AOI21_X1 U5897 ( .B1(n5915), .B2(n4743), .A(n4718), .ZN(n4719) );
  OAI211_X1 U5898 ( .C1(n4808), .C2(n6448), .A(n4720), .B(n4719), .ZN(U3136)
         );
  NAND2_X1 U5899 ( .A1(n4739), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4723)
         );
  OAI22_X1 U5900 ( .A1(n5936), .A2(n4741), .B1(n4740), .B2(n5933), .ZN(n4721)
         );
  AOI21_X1 U5901 ( .B1(n5939), .B2(n4743), .A(n4721), .ZN(n4722) );
  OAI211_X1 U5902 ( .C1(n4808), .C2(n5942), .A(n4723), .B(n4722), .ZN(U3139)
         );
  NAND2_X1 U5903 ( .A1(n4739), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4726)
         );
  OAI22_X1 U5904 ( .A1(n6431), .A2(n4741), .B1(n4740), .B2(n5908), .ZN(n4724)
         );
  AOI21_X1 U5905 ( .B1(n5910), .B2(n4743), .A(n4724), .ZN(n4725) );
  OAI211_X1 U5906 ( .C1(n4808), .C2(n6436), .A(n4726), .B(n4725), .ZN(U3135)
         );
  NAND2_X1 U5907 ( .A1(n4739), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4729)
         );
  OAI22_X1 U5908 ( .A1(n5902), .A2(n4741), .B1(n4740), .B2(n5901), .ZN(n4727)
         );
  AOI21_X1 U5909 ( .B1(n5904), .B2(n4743), .A(n4727), .ZN(n4728) );
  OAI211_X1 U5910 ( .C1(n4808), .C2(n5907), .A(n4729), .B(n4728), .ZN(U3134)
         );
  NAND2_X1 U5911 ( .A1(n4739), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4732)
         );
  OAI22_X1 U5912 ( .A1(n5895), .A2(n4741), .B1(n4740), .B2(n5894), .ZN(n4730)
         );
  AOI21_X1 U5913 ( .B1(n5897), .B2(n4743), .A(n4730), .ZN(n4731) );
  OAI211_X1 U5914 ( .C1(n4808), .C2(n5900), .A(n4732), .B(n4731), .ZN(U3133)
         );
  NAND2_X1 U5915 ( .A1(n4739), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4735)
         );
  OAI22_X1 U5916 ( .A1(n5926), .A2(n4741), .B1(n4740), .B2(n5925), .ZN(n4733)
         );
  AOI21_X1 U5917 ( .B1(n5928), .B2(n4743), .A(n4733), .ZN(n4734) );
  OAI211_X1 U5918 ( .C1(n4808), .C2(n5931), .A(n4735), .B(n4734), .ZN(U3138)
         );
  NAND2_X1 U5919 ( .A1(n4739), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4738)
         );
  OAI22_X1 U5920 ( .A1(n6451), .A2(n4741), .B1(n4740), .B2(n5889), .ZN(n4736)
         );
  AOI21_X1 U5921 ( .B1(n5891), .B2(n4743), .A(n4736), .ZN(n4737) );
  OAI211_X1 U5922 ( .C1(n4808), .C2(n6461), .A(n4738), .B(n4737), .ZN(U3132)
         );
  NAND2_X1 U5923 ( .A1(n4739), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4745)
         );
  OAI22_X1 U5924 ( .A1(n5919), .A2(n4741), .B1(n4740), .B2(n5918), .ZN(n4742)
         );
  AOI21_X1 U5925 ( .B1(n5921), .B2(n4743), .A(n4742), .ZN(n4744) );
  OAI211_X1 U5926 ( .C1(n4808), .C2(n5924), .A(n4745), .B(n4744), .ZN(U3137)
         );
  INV_X1 U5927 ( .A(n4746), .ZN(n4810) );
  AND2_X1 U5928 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4754), .ZN(n4750)
         );
  AOI21_X1 U5929 ( .B1(n4810), .B2(n4747), .A(n4750), .ZN(n4752) );
  NAND2_X1 U5930 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4749) );
  OAI22_X1 U5931 ( .A1(n4752), .A2(n5875), .B1(n4749), .B2(n4748), .ZN(n4806)
         );
  NOR2_X1 U5932 ( .A1(n4800), .A2(n5942), .ZN(n4760) );
  INV_X1 U5933 ( .A(n4750), .ZN(n4803) );
  NAND2_X1 U5934 ( .A1(n4752), .A2(n4751), .ZN(n4753) );
  OR2_X1 U5935 ( .A1(n5875), .A2(n4753), .ZN(n4757) );
  INV_X1 U5936 ( .A(n4754), .ZN(n4755) );
  NAND2_X1 U5937 ( .A1(n5875), .A2(n4755), .ZN(n4756) );
  INV_X1 U5938 ( .A(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4758) );
  OAI22_X1 U5939 ( .A1(n5936), .A2(n4803), .B1(n4802), .B2(n4758), .ZN(n4759)
         );
  AOI211_X1 U5940 ( .C1(n6417), .C2(n4806), .A(n4760), .B(n4759), .ZN(n4761)
         );
  OAI21_X1 U5941 ( .B1(n6425), .B2(n4808), .A(n4761), .ZN(U3131) );
  NOR2_X1 U5942 ( .A1(n4800), .A2(n6436), .ZN(n4764) );
  INV_X1 U5943 ( .A(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4762) );
  OAI22_X1 U5944 ( .A1(n6431), .A2(n4803), .B1(n4802), .B2(n4762), .ZN(n4763)
         );
  AOI211_X1 U5945 ( .C1(n6433), .C2(n4806), .A(n4764), .B(n4763), .ZN(n4765)
         );
  OAI21_X1 U5946 ( .B1(n6430), .B2(n4808), .A(n4765), .ZN(U3127) );
  NOR2_X1 U5947 ( .A1(n4800), .A2(n5907), .ZN(n4768) );
  INV_X1 U5948 ( .A(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4766) );
  OAI22_X1 U5949 ( .A1(n5902), .A2(n4803), .B1(n4802), .B2(n4766), .ZN(n4767)
         );
  AOI211_X1 U5950 ( .C1(n6390), .C2(n4806), .A(n4768), .B(n4767), .ZN(n4769)
         );
  OAI21_X1 U5951 ( .B1(n6395), .B2(n4808), .A(n4769), .ZN(U3126) );
  NOR2_X1 U5952 ( .A1(n4800), .A2(n6461), .ZN(n4772) );
  INV_X1 U5953 ( .A(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4770) );
  OAI22_X1 U5954 ( .A1(n6451), .A2(n4803), .B1(n4802), .B2(n4770), .ZN(n4771)
         );
  AOI211_X1 U5955 ( .C1(n6456), .C2(n4806), .A(n4772), .B(n4771), .ZN(n4773)
         );
  OAI21_X1 U5956 ( .B1(n6452), .B2(n4808), .A(n4773), .ZN(U3124) );
  NAND2_X1 U5957 ( .A1(n4775), .A2(n4774), .ZN(n4776) );
  NAND2_X1 U5958 ( .A1(n4422), .A2(n4776), .ZN(n4778) );
  NAND2_X1 U5959 ( .A1(n6221), .A2(n3230), .ZN(n5176) );
  AND2_X2 U5960 ( .A1(n4779), .A2(n6499), .ZN(n6243) );
  INV_X1 U5961 ( .A(n6243), .ZN(n6492) );
  AOI22_X1 U5962 ( .A1(n6243), .A2(UWORD_REG_12__SCAN_IN), .B1(n6242), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4780) );
  OAI21_X1 U5963 ( .B1(n4404), .B2(n5176), .A(n4780), .ZN(U2895) );
  AOI22_X1 U5964 ( .A1(n6243), .A2(UWORD_REG_11__SCAN_IN), .B1(n6242), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4781) );
  OAI21_X1 U5965 ( .B1(n4362), .B2(n5176), .A(n4781), .ZN(U2896) );
  AOI22_X1 U5966 ( .A1(n6243), .A2(UWORD_REG_9__SCAN_IN), .B1(n6242), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4782) );
  OAI21_X1 U5967 ( .B1(n4366), .B2(n5176), .A(n4782), .ZN(U2898) );
  INV_X1 U5968 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4784) );
  AOI22_X1 U5969 ( .A1(n6243), .A2(UWORD_REG_8__SCAN_IN), .B1(n6242), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4783) );
  OAI21_X1 U5970 ( .B1(n4784), .B2(n5176), .A(n4783), .ZN(U2899) );
  AOI22_X1 U5971 ( .A1(n6243), .A2(UWORD_REG_14__SCAN_IN), .B1(n6242), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4785) );
  OAI21_X1 U5972 ( .B1(n4391), .B2(n5176), .A(n4785), .ZN(U2893) );
  AOI22_X1 U5973 ( .A1(n6243), .A2(UWORD_REG_13__SCAN_IN), .B1(n6242), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4786) );
  OAI21_X1 U5974 ( .B1(n4401), .B2(n5176), .A(n4786), .ZN(U2894) );
  AOI22_X1 U5975 ( .A1(n6243), .A2(UWORD_REG_10__SCAN_IN), .B1(n6242), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4787) );
  OAI21_X1 U5976 ( .B1(n4355), .B2(n5176), .A(n4787), .ZN(U2897) );
  NOR2_X1 U5977 ( .A1(n4800), .A2(n5900), .ZN(n4790) );
  INV_X1 U5978 ( .A(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4788) );
  OAI22_X1 U5979 ( .A1(n5895), .A2(n4803), .B1(n4802), .B2(n4788), .ZN(n4789)
         );
  AOI211_X1 U5980 ( .C1(n6384), .C2(n4806), .A(n4790), .B(n4789), .ZN(n4791)
         );
  OAI21_X1 U5981 ( .B1(n6389), .B2(n4808), .A(n4791), .ZN(U3125) );
  NOR2_X1 U5982 ( .A1(n4800), .A2(n6448), .ZN(n4794) );
  INV_X1 U5983 ( .A(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4792) );
  OAI22_X1 U5984 ( .A1(n6440), .A2(n4803), .B1(n4802), .B2(n4792), .ZN(n4793)
         );
  AOI211_X1 U5985 ( .C1(n6443), .C2(n4806), .A(n4794), .B(n4793), .ZN(n4795)
         );
  OAI21_X1 U5986 ( .B1(n6437), .B2(n4808), .A(n4795), .ZN(U3128) );
  NOR2_X1 U5987 ( .A1(n4800), .A2(n5931), .ZN(n4798) );
  INV_X1 U5988 ( .A(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4796) );
  OAI22_X1 U5989 ( .A1(n5926), .A2(n4803), .B1(n4802), .B2(n4796), .ZN(n4797)
         );
  AOI211_X1 U5990 ( .C1(n6410), .C2(n4806), .A(n4798), .B(n4797), .ZN(n4799)
         );
  OAI21_X1 U5991 ( .B1(n6415), .B2(n4808), .A(n4799), .ZN(U3130) );
  NOR2_X1 U5992 ( .A1(n4800), .A2(n5924), .ZN(n4805) );
  INV_X1 U5993 ( .A(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4801) );
  OAI22_X1 U5994 ( .A1(n5919), .A2(n4803), .B1(n4802), .B2(n4801), .ZN(n4804)
         );
  AOI211_X1 U5995 ( .C1(n6404), .C2(n4806), .A(n4805), .B(n4804), .ZN(n4807)
         );
  OAI21_X1 U5996 ( .B1(n6409), .B2(n4808), .A(n4807), .ZN(U3129) );
  AOI21_X1 U5997 ( .B1(n4815), .B2(STATEBS16_REG_SCAN_IN), .A(n5875), .ZN(
        n4812) );
  NOR2_X1 U5998 ( .A1(n6170), .A2(n4339), .ZN(n4922) );
  NAND3_X1 U5999 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6471), .A3(n4838), .ZN(n4923) );
  NOR2_X1 U6000 ( .A1(n6364), .A2(n4923), .ZN(n4816) );
  AOI21_X1 U6001 ( .B1(n4810), .B2(n4922), .A(n4816), .ZN(n4814) );
  AOI22_X1 U6002 ( .A1(n4812), .A2(n4814), .B1(n5875), .B2(n4923), .ZN(n4811)
         );
  NAND2_X1 U6003 ( .A1(n4879), .A2(n4811), .ZN(n4915) );
  INV_X1 U6004 ( .A(n4812), .ZN(n4813) );
  OAI22_X1 U6005 ( .A1(n4814), .A2(n4813), .B1(n6498), .B2(n4923), .ZN(n4914)
         );
  AOI22_X1 U6006 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4915), .B1(n6417), 
        .B2(n4914), .ZN(n4819) );
  NAND2_X1 U6007 ( .A1(n4815), .A2(n4975), .ZN(n4920) );
  INV_X1 U6008 ( .A(n4816), .ZN(n4916) );
  OAI22_X1 U6009 ( .A1(n5084), .A2(n6425), .B1(n5936), .B2(n4916), .ZN(n4817)
         );
  AOI21_X1 U6010 ( .B1(n6421), .B2(n4962), .A(n4817), .ZN(n4818) );
  NAND2_X1 U6011 ( .A1(n4819), .A2(n4818), .ZN(U3099) );
  AOI22_X1 U6012 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4915), .B1(n6384), 
        .B2(n4914), .ZN(n4822) );
  OAI22_X1 U6013 ( .A1(n5084), .A2(n6389), .B1(n5895), .B2(n4916), .ZN(n4820)
         );
  AOI21_X1 U6014 ( .B1(n6386), .B2(n4962), .A(n4820), .ZN(n4821) );
  NAND2_X1 U6015 ( .A1(n4822), .A2(n4821), .ZN(U3093) );
  AOI22_X1 U6016 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4915), .B1(n6410), 
        .B2(n4914), .ZN(n4825) );
  OAI22_X1 U6017 ( .A1(n5084), .A2(n6415), .B1(n5926), .B2(n4916), .ZN(n4823)
         );
  AOI21_X1 U6018 ( .B1(n6412), .B2(n4962), .A(n4823), .ZN(n4824) );
  NAND2_X1 U6019 ( .A1(n4825), .A2(n4824), .ZN(U3098) );
  AOI22_X1 U6020 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4915), .B1(n6390), 
        .B2(n4914), .ZN(n4828) );
  OAI22_X1 U6021 ( .A1(n5084), .A2(n6395), .B1(n5902), .B2(n4916), .ZN(n4826)
         );
  AOI21_X1 U6022 ( .B1(n6392), .B2(n4962), .A(n4826), .ZN(n4827) );
  NAND2_X1 U6023 ( .A1(n4828), .A2(n4827), .ZN(U3094) );
  AOI22_X1 U6024 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4915), .B1(n6404), 
        .B2(n4914), .ZN(n4831) );
  OAI22_X1 U6025 ( .A1(n5084), .A2(n6409), .B1(n5919), .B2(n4916), .ZN(n4829)
         );
  AOI21_X1 U6026 ( .B1(n6406), .B2(n4962), .A(n4829), .ZN(n4830) );
  NAND2_X1 U6027 ( .A1(n4831), .A2(n4830), .ZN(U3097) );
  AOI22_X1 U6028 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4915), .B1(n6433), 
        .B2(n4914), .ZN(n4834) );
  OAI22_X1 U6029 ( .A1(n5084), .A2(n6430), .B1(n6431), .B2(n4916), .ZN(n4832)
         );
  AOI21_X1 U6030 ( .B1(n6397), .B2(n4962), .A(n4832), .ZN(n4833) );
  NAND2_X1 U6031 ( .A1(n4834), .A2(n4833), .ZN(U3095) );
  OR2_X1 U6032 ( .A1(n4836), .A2(n4835), .ZN(n4837) );
  AOI21_X1 U6033 ( .B1(n4913), .B2(n4843), .A(n6728), .ZN(n4842) );
  NAND2_X1 U6034 ( .A1(n6368), .A2(n4922), .ZN(n4844) );
  NAND2_X1 U6035 ( .A1(n4844), .A2(n6367), .ZN(n4841) );
  NAND3_X1 U6036 ( .A1(n6478), .A2(n6471), .A3(n4838), .ZN(n4881) );
  OR2_X1 U6037 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4881), .ZN(n4869)
         );
  AOI211_X1 U6038 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4869), .A(n5078), .B(
        n4839), .ZN(n4840) );
  NAND2_X1 U6039 ( .A1(n4867), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4848) );
  INV_X1 U6040 ( .A(n4844), .ZN(n4877) );
  AOI22_X1 U6041 ( .A1(n4877), .A2(n6367), .B1(n5887), .B2(n4845), .ZN(n4868)
         );
  OAI22_X1 U6042 ( .A1(n5919), .A2(n4869), .B1(n4868), .B2(n5918), .ZN(n4846)
         );
  AOI21_X1 U6043 ( .B1(n6406), .B2(n4871), .A(n4846), .ZN(n4847) );
  OAI211_X1 U6044 ( .C1(n4913), .C2(n6409), .A(n4848), .B(n4847), .ZN(U3025)
         );
  NAND2_X1 U6045 ( .A1(n4867), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4851) );
  OAI22_X1 U6046 ( .A1(n5936), .A2(n4869), .B1(n4868), .B2(n5933), .ZN(n4849)
         );
  AOI21_X1 U6047 ( .B1(n6421), .B2(n4871), .A(n4849), .ZN(n4850) );
  OAI211_X1 U6048 ( .C1(n4913), .C2(n6425), .A(n4851), .B(n4850), .ZN(U3027)
         );
  NAND2_X1 U6049 ( .A1(n4867), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4854) );
  OAI22_X1 U6050 ( .A1(n5926), .A2(n4869), .B1(n4868), .B2(n5925), .ZN(n4852)
         );
  AOI21_X1 U6051 ( .B1(n6412), .B2(n4871), .A(n4852), .ZN(n4853) );
  OAI211_X1 U6052 ( .C1(n4913), .C2(n6415), .A(n4854), .B(n4853), .ZN(U3026)
         );
  NAND2_X1 U6053 ( .A1(n4867), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4857) );
  OAI22_X1 U6054 ( .A1(n5902), .A2(n4869), .B1(n4868), .B2(n5901), .ZN(n4855)
         );
  AOI21_X1 U6055 ( .B1(n6392), .B2(n4871), .A(n4855), .ZN(n4856) );
  OAI211_X1 U6056 ( .C1(n4913), .C2(n6395), .A(n4857), .B(n4856), .ZN(U3022)
         );
  NAND2_X1 U6057 ( .A1(n4867), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4860) );
  OAI22_X1 U6058 ( .A1(n5895), .A2(n4869), .B1(n4868), .B2(n5894), .ZN(n4858)
         );
  AOI21_X1 U6059 ( .B1(n6386), .B2(n4871), .A(n4858), .ZN(n4859) );
  OAI211_X1 U6060 ( .C1(n4913), .C2(n6389), .A(n4860), .B(n4859), .ZN(U3021)
         );
  NAND2_X1 U6061 ( .A1(n4867), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4863) );
  OAI22_X1 U6062 ( .A1(n6440), .A2(n4869), .B1(n4868), .B2(n5913), .ZN(n4861)
         );
  AOI21_X1 U6063 ( .B1(n6401), .B2(n4871), .A(n4861), .ZN(n4862) );
  OAI211_X1 U6064 ( .C1(n4913), .C2(n6437), .A(n4863), .B(n4862), .ZN(U3024)
         );
  NAND2_X1 U6065 ( .A1(n4867), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4866) );
  OAI22_X1 U6066 ( .A1(n6451), .A2(n4869), .B1(n4868), .B2(n5889), .ZN(n4864)
         );
  AOI21_X1 U6067 ( .B1(n6381), .B2(n4871), .A(n4864), .ZN(n4865) );
  OAI211_X1 U6068 ( .C1(n4913), .C2(n6452), .A(n4866), .B(n4865), .ZN(U3020)
         );
  NAND2_X1 U6069 ( .A1(n4867), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4873) );
  OAI22_X1 U6070 ( .A1(n6431), .A2(n4869), .B1(n4868), .B2(n5908), .ZN(n4870)
         );
  AOI21_X1 U6071 ( .B1(n6397), .B2(n4871), .A(n4870), .ZN(n4872) );
  OAI211_X1 U6072 ( .C1(n4913), .C2(n6430), .A(n4873), .B(n4872), .ZN(U3023)
         );
  AOI22_X1 U6073 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4915), .B1(n6443), 
        .B2(n4914), .ZN(n4876) );
  OAI22_X1 U6074 ( .A1(n5084), .A2(n6437), .B1(n6440), .B2(n4916), .ZN(n4874)
         );
  AOI21_X1 U6075 ( .B1(n6401), .B2(n4962), .A(n4874), .ZN(n4875) );
  NAND2_X1 U6076 ( .A1(n4876), .A2(n4875), .ZN(U3096) );
  NOR2_X1 U6077 ( .A1(n6364), .A2(n4881), .ZN(n4885) );
  AOI21_X1 U6078 ( .B1(n4877), .B2(n3808), .A(n4885), .ZN(n4883) );
  AOI21_X1 U6079 ( .B1(n4884), .B2(STATEBS16_REG_SCAN_IN), .A(n5875), .ZN(
        n4880) );
  AOI22_X1 U6080 ( .A1(n4883), .A2(n4880), .B1(n5875), .B2(n4881), .ZN(n4878)
         );
  NAND2_X1 U6081 ( .A1(n4879), .A2(n4878), .ZN(n4908) );
  INV_X1 U6082 ( .A(n4880), .ZN(n4882) );
  OAI22_X1 U6083 ( .A1(n4883), .A2(n4882), .B1(n6498), .B2(n4881), .ZN(n4907)
         );
  AOI22_X1 U6084 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4908), .B1(n6433), 
        .B2(n4907), .ZN(n4888) );
  INV_X1 U6085 ( .A(n4885), .ZN(n4909) );
  OAI22_X1 U6086 ( .A1(n5943), .A2(n6430), .B1(n6431), .B2(n4909), .ZN(n4886)
         );
  INV_X1 U6087 ( .A(n4886), .ZN(n4887) );
  OAI211_X1 U6088 ( .C1(n6436), .C2(n4913), .A(n4888), .B(n4887), .ZN(U3031)
         );
  AOI22_X1 U6089 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4908), .B1(n6384), 
        .B2(n4907), .ZN(n4891) );
  OAI22_X1 U6090 ( .A1(n5943), .A2(n6389), .B1(n5895), .B2(n4909), .ZN(n4889)
         );
  INV_X1 U6091 ( .A(n4889), .ZN(n4890) );
  OAI211_X1 U6092 ( .C1(n5900), .C2(n4913), .A(n4891), .B(n4890), .ZN(U3029)
         );
  AOI22_X1 U6093 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4908), .B1(n6456), 
        .B2(n4907), .ZN(n4894) );
  OAI22_X1 U6094 ( .A1(n5943), .A2(n6452), .B1(n6451), .B2(n4909), .ZN(n4892)
         );
  INV_X1 U6095 ( .A(n4892), .ZN(n4893) );
  OAI211_X1 U6096 ( .C1(n6461), .C2(n4913), .A(n4894), .B(n4893), .ZN(U3028)
         );
  AOI22_X1 U6097 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4908), .B1(n6390), 
        .B2(n4907), .ZN(n4897) );
  OAI22_X1 U6098 ( .A1(n5943), .A2(n6395), .B1(n5902), .B2(n4909), .ZN(n4895)
         );
  INV_X1 U6099 ( .A(n4895), .ZN(n4896) );
  OAI211_X1 U6100 ( .C1(n5907), .C2(n4913), .A(n4897), .B(n4896), .ZN(U3030)
         );
  AOI22_X1 U6101 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4908), .B1(n6417), 
        .B2(n4907), .ZN(n4900) );
  OAI22_X1 U6102 ( .A1(n5943), .A2(n6425), .B1(n5936), .B2(n4909), .ZN(n4898)
         );
  INV_X1 U6103 ( .A(n4898), .ZN(n4899) );
  OAI211_X1 U6104 ( .C1(n5942), .C2(n4913), .A(n4900), .B(n4899), .ZN(U3035)
         );
  AOI22_X1 U6105 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4908), .B1(n6410), 
        .B2(n4907), .ZN(n4903) );
  OAI22_X1 U6106 ( .A1(n5943), .A2(n6415), .B1(n5926), .B2(n4909), .ZN(n4901)
         );
  INV_X1 U6107 ( .A(n4901), .ZN(n4902) );
  OAI211_X1 U6108 ( .C1(n5931), .C2(n4913), .A(n4903), .B(n4902), .ZN(U3034)
         );
  AOI22_X1 U6109 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4908), .B1(n6404), 
        .B2(n4907), .ZN(n4906) );
  OAI22_X1 U6110 ( .A1(n5943), .A2(n6409), .B1(n5919), .B2(n4909), .ZN(n4904)
         );
  INV_X1 U6111 ( .A(n4904), .ZN(n4905) );
  OAI211_X1 U6112 ( .C1(n5924), .C2(n4913), .A(n4906), .B(n4905), .ZN(U3033)
         );
  AOI22_X1 U6113 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4908), .B1(n6443), 
        .B2(n4907), .ZN(n4912) );
  OAI22_X1 U6114 ( .A1(n5943), .A2(n6437), .B1(n6440), .B2(n4909), .ZN(n4910)
         );
  INV_X1 U6115 ( .A(n4910), .ZN(n4911) );
  OAI211_X1 U6116 ( .C1(n6448), .C2(n4913), .A(n4912), .B(n4911), .ZN(U3032)
         );
  AOI22_X1 U6117 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4915), .B1(n6456), 
        .B2(n4914), .ZN(n4919) );
  OAI22_X1 U6118 ( .A1(n5084), .A2(n6452), .B1(n6451), .B2(n4916), .ZN(n4917)
         );
  INV_X1 U6119 ( .A(n4917), .ZN(n4918) );
  OAI211_X1 U6120 ( .C1(n6461), .C2(n4920), .A(n4919), .B(n4918), .ZN(U3092)
         );
  NAND3_X1 U6121 ( .A1(n4920), .A2(n6367), .A3(n6438), .ZN(n4921) );
  INV_X1 U6122 ( .A(n6375), .ZN(n5879) );
  NAND2_X1 U6123 ( .A1(n4921), .A2(n5879), .ZN(n4926) );
  NAND2_X1 U6124 ( .A1(n4922), .A2(n6167), .ZN(n4929) );
  NOR2_X1 U6125 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4923), .ZN(n4959)
         );
  INV_X1 U6126 ( .A(n5078), .ZN(n6371) );
  OAI211_X1 U6127 ( .C1(n6592), .C2(n4959), .A(n6371), .B(n4924), .ZN(n4925)
         );
  INV_X1 U6128 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4933) );
  OAI22_X1 U6129 ( .A1(n4929), .A2(n5875), .B1(n4928), .B2(n4927), .ZN(n4958)
         );
  AOI22_X1 U6130 ( .A1(n6411), .A2(n4959), .B1(n6410), .B2(n4958), .ZN(n4930)
         );
  OAI21_X1 U6131 ( .B1(n5931), .B2(n6438), .A(n4930), .ZN(n4931) );
  AOI21_X1 U6132 ( .B1(n5928), .B2(n4962), .A(n4931), .ZN(n4932) );
  OAI21_X1 U6133 ( .B1(n4965), .B2(n4933), .A(n4932), .ZN(U3090) );
  INV_X1 U6134 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4937) );
  AOI22_X1 U6135 ( .A1(n6419), .A2(n4959), .B1(n6417), .B2(n4958), .ZN(n4934)
         );
  OAI21_X1 U6136 ( .B1(n5942), .B2(n6438), .A(n4934), .ZN(n4935) );
  AOI21_X1 U6137 ( .B1(n5939), .B2(n4962), .A(n4935), .ZN(n4936) );
  OAI21_X1 U6138 ( .B1(n4965), .B2(n4937), .A(n4936), .ZN(U3091) );
  INV_X1 U6139 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4941) );
  INV_X1 U6140 ( .A(n6451), .ZN(n6372) );
  AOI22_X1 U6141 ( .A1(n6372), .A2(n4959), .B1(n6456), .B2(n4958), .ZN(n4938)
         );
  OAI21_X1 U6142 ( .B1(n6461), .B2(n6438), .A(n4938), .ZN(n4939) );
  AOI21_X1 U6143 ( .B1(n5891), .B2(n4962), .A(n4939), .ZN(n4940) );
  OAI21_X1 U6144 ( .B1(n4965), .B2(n4941), .A(n4940), .ZN(U3084) );
  INV_X1 U6145 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4945) );
  AOI22_X1 U6146 ( .A1(n6385), .A2(n4959), .B1(n6384), .B2(n4958), .ZN(n4942)
         );
  OAI21_X1 U6147 ( .B1(n5900), .B2(n6438), .A(n4942), .ZN(n4943) );
  AOI21_X1 U6148 ( .B1(n5897), .B2(n4962), .A(n4943), .ZN(n4944) );
  OAI21_X1 U6149 ( .B1(n4965), .B2(n4945), .A(n4944), .ZN(U3085) );
  INV_X1 U6150 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4949) );
  AOI22_X1 U6151 ( .A1(n6391), .A2(n4959), .B1(n6390), .B2(n4958), .ZN(n4946)
         );
  OAI21_X1 U6152 ( .B1(n5907), .B2(n6438), .A(n4946), .ZN(n4947) );
  AOI21_X1 U6153 ( .B1(n5904), .B2(n4962), .A(n4947), .ZN(n4948) );
  OAI21_X1 U6154 ( .B1(n4965), .B2(n4949), .A(n4948), .ZN(U3086) );
  INV_X1 U6155 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4953) );
  AOI22_X1 U6156 ( .A1(n6396), .A2(n4959), .B1(n6433), .B2(n4958), .ZN(n4950)
         );
  OAI21_X1 U6157 ( .B1(n6436), .B2(n6438), .A(n4950), .ZN(n4951) );
  AOI21_X1 U6158 ( .B1(n5910), .B2(n4962), .A(n4951), .ZN(n4952) );
  OAI21_X1 U6159 ( .B1(n4965), .B2(n4953), .A(n4952), .ZN(U3087) );
  INV_X1 U6160 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4957) );
  AOI22_X1 U6161 ( .A1(n6400), .A2(n4959), .B1(n6443), .B2(n4958), .ZN(n4954)
         );
  OAI21_X1 U6162 ( .B1(n6448), .B2(n6438), .A(n4954), .ZN(n4955) );
  AOI21_X1 U6163 ( .B1(n5915), .B2(n4962), .A(n4955), .ZN(n4956) );
  OAI21_X1 U6164 ( .B1(n4965), .B2(n4957), .A(n4956), .ZN(U3088) );
  INV_X1 U6165 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4964) );
  AOI22_X1 U6166 ( .A1(n6405), .A2(n4959), .B1(n6404), .B2(n4958), .ZN(n4960)
         );
  OAI21_X1 U6167 ( .B1(n5924), .B2(n6438), .A(n4960), .ZN(n4961) );
  AOI21_X1 U6168 ( .B1(n5921), .B2(n4962), .A(n4961), .ZN(n4963) );
  OAI21_X1 U6169 ( .B1(n4965), .B2(n4964), .A(n4963), .ZN(U3089) );
  NOR2_X1 U6170 ( .A1(n6364), .A2(n4972), .ZN(n5005) );
  INV_X1 U6171 ( .A(n5005), .ZN(n4966) );
  OAI21_X1 U6172 ( .B1(n4968), .B2(n4967), .A(n4966), .ZN(n4971) );
  NOR2_X1 U6173 ( .A1(n4974), .A2(n4971), .ZN(n4969) );
  INV_X1 U6174 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4980) );
  INV_X1 U6175 ( .A(n4971), .ZN(n4973) );
  OAI22_X1 U6176 ( .A1(n4974), .A2(n4973), .B1(n4972), .B2(n6498), .ZN(n5009)
         );
  NOR2_X2 U6177 ( .A1(n4976), .A2(n4975), .ZN(n6420) );
  AOI22_X1 U6178 ( .A1(n6420), .A2(n5915), .B1(n6400), .B2(n5005), .ZN(n4977)
         );
  OAI21_X1 U6179 ( .B1(n6448), .B2(n5007), .A(n4977), .ZN(n4978) );
  AOI21_X1 U6180 ( .B1(n6443), .B2(n5009), .A(n4978), .ZN(n4979) );
  OAI21_X1 U6181 ( .B1(n5012), .B2(n4980), .A(n4979), .ZN(U3064) );
  INV_X1 U6182 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4984) );
  AOI22_X1 U6183 ( .A1(n6420), .A2(n5910), .B1(n6396), .B2(n5005), .ZN(n4981)
         );
  OAI21_X1 U6184 ( .B1(n6436), .B2(n5007), .A(n4981), .ZN(n4982) );
  AOI21_X1 U6185 ( .B1(n6433), .B2(n5009), .A(n4982), .ZN(n4983) );
  OAI21_X1 U6186 ( .B1(n5012), .B2(n4984), .A(n4983), .ZN(U3063) );
  INV_X1 U6187 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4988) );
  AOI22_X1 U6188 ( .A1(n6420), .A2(n5928), .B1(n6411), .B2(n5005), .ZN(n4985)
         );
  OAI21_X1 U6189 ( .B1(n5931), .B2(n5007), .A(n4985), .ZN(n4986) );
  AOI21_X1 U6190 ( .B1(n6410), .B2(n5009), .A(n4986), .ZN(n4987) );
  OAI21_X1 U6191 ( .B1(n5012), .B2(n4988), .A(n4987), .ZN(U3066) );
  INV_X1 U6192 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4992) );
  AOI22_X1 U6193 ( .A1(n6420), .A2(n5939), .B1(n6419), .B2(n5005), .ZN(n4989)
         );
  OAI21_X1 U6194 ( .B1(n5942), .B2(n5007), .A(n4989), .ZN(n4990) );
  AOI21_X1 U6195 ( .B1(n6417), .B2(n5009), .A(n4990), .ZN(n4991) );
  OAI21_X1 U6196 ( .B1(n5012), .B2(n4992), .A(n4991), .ZN(U3067) );
  INV_X1 U6197 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4996) );
  AOI22_X1 U6198 ( .A1(n6420), .A2(n5891), .B1(n6372), .B2(n5005), .ZN(n4993)
         );
  OAI21_X1 U6199 ( .B1(n6461), .B2(n5007), .A(n4993), .ZN(n4994) );
  AOI21_X1 U6200 ( .B1(n6456), .B2(n5009), .A(n4994), .ZN(n4995) );
  OAI21_X1 U6201 ( .B1(n5012), .B2(n4996), .A(n4995), .ZN(U3060) );
  INV_X1 U6202 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n5000) );
  AOI22_X1 U6203 ( .A1(n6420), .A2(n5897), .B1(n6385), .B2(n5005), .ZN(n4997)
         );
  OAI21_X1 U6204 ( .B1(n5900), .B2(n5007), .A(n4997), .ZN(n4998) );
  AOI21_X1 U6205 ( .B1(n6384), .B2(n5009), .A(n4998), .ZN(n4999) );
  OAI21_X1 U6206 ( .B1(n5012), .B2(n5000), .A(n4999), .ZN(U3061) );
  INV_X1 U6207 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n5004) );
  AOI22_X1 U6208 ( .A1(n6420), .A2(n5904), .B1(n6391), .B2(n5005), .ZN(n5001)
         );
  OAI21_X1 U6209 ( .B1(n5907), .B2(n5007), .A(n5001), .ZN(n5002) );
  AOI21_X1 U6210 ( .B1(n6390), .B2(n5009), .A(n5002), .ZN(n5003) );
  OAI21_X1 U6211 ( .B1(n5012), .B2(n5004), .A(n5003), .ZN(U3062) );
  INV_X1 U6212 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n5011) );
  AOI22_X1 U6213 ( .A1(n6420), .A2(n5921), .B1(n6405), .B2(n5005), .ZN(n5006)
         );
  OAI21_X1 U6214 ( .B1(n5924), .B2(n5007), .A(n5006), .ZN(n5008) );
  AOI21_X1 U6215 ( .B1(n6404), .B2(n5009), .A(n5008), .ZN(n5010) );
  OAI21_X1 U6216 ( .B1(n5012), .B2(n5011), .A(n5010), .ZN(U3065) );
  XOR2_X1 U6217 ( .A(n5014), .B(n5013), .Z(n5073) );
  INV_X1 U6218 ( .A(n5073), .ZN(n5040) );
  AOI21_X1 U6219 ( .B1(n5016), .B2(n5015), .A(n5134), .ZN(n6318) );
  AOI22_X1 U6220 ( .A1(n6318), .A2(n6203), .B1(EBX_REG_7__SCAN_IN), .B2(n5617), 
        .ZN(n5017) );
  OAI21_X1 U6221 ( .B1(n5040), .B2(n5639), .A(n5017), .ZN(U2852) );
  AOI22_X1 U6222 ( .A1(EBX_REG_7__SCAN_IN), .A2(n6182), .B1(n6122), .B2(n6318), 
        .ZN(n5018) );
  OAI211_X1 U6223 ( .C1(n6138), .C2(n5019), .A(n5018), .B(n6341), .ZN(n5027)
         );
  NOR3_X1 U6224 ( .A1(n6176), .A2(REIP_REG_6__SCAN_IN), .A3(n5020), .ZN(n6144)
         );
  NAND2_X1 U6225 ( .A1(n6193), .A2(n5020), .ZN(n5021) );
  NAND2_X1 U6226 ( .A1(n5021), .A2(n6159), .ZN(n6145) );
  OAI21_X1 U6227 ( .B1(n6144), .B2(n6145), .A(REIP_REG_7__SCAN_IN), .ZN(n5025)
         );
  INV_X1 U6228 ( .A(n5022), .ZN(n5023) );
  OR3_X1 U6229 ( .A1(n6176), .A2(REIP_REG_7__SCAN_IN), .A3(n5023), .ZN(n5024)
         );
  OAI211_X1 U6230 ( .C1(n6187), .C2(n5071), .A(n5025), .B(n5024), .ZN(n5026)
         );
  AOI211_X1 U6231 ( .C1(n5073), .C2(n6146), .A(n5027), .B(n5026), .ZN(n5028)
         );
  INV_X1 U6232 ( .A(n5028), .ZN(U2820) );
  NAND2_X1 U6233 ( .A1(n6609), .A2(n5029), .ZN(n5030) );
  INV_X1 U6234 ( .A(n6145), .ZN(n5033) );
  AOI21_X1 U6235 ( .B1(n6193), .B2(n5031), .A(REIP_REG_5__SCAN_IN), .ZN(n5032)
         );
  NOR2_X1 U6236 ( .A1(n5033), .A2(n5032), .ZN(n5037) );
  AOI22_X1 U6237 ( .A1(EBX_REG_5__SCAN_IN), .A2(n6182), .B1(n6122), .B2(n6332), 
        .ZN(n5034) );
  OAI211_X1 U6238 ( .C1(n6138), .C2(n5035), .A(n5034), .B(n6341), .ZN(n5036)
         );
  AOI211_X1 U6239 ( .C1(n6160), .C2(n5060), .A(n5037), .B(n5036), .ZN(n5038)
         );
  OAI21_X1 U6240 ( .B1(n6188), .B2(n5059), .A(n5038), .ZN(U2822) );
  OAI222_X1 U6241 ( .A1(n5983), .A2(n5040), .B1(n5039), .B2(n6818), .C1(n5640), 
        .C2(n4388), .ZN(U2884) );
  INV_X1 U6242 ( .A(n6189), .ZN(n5044) );
  AOI21_X1 U6243 ( .B1(n6263), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n5041), 
        .ZN(n5042) );
  OAI21_X1 U6244 ( .B1(n6281), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n5042), 
        .ZN(n5043) );
  AOI21_X1 U6245 ( .B1(n5044), .B2(n5749), .A(n5043), .ZN(n5045) );
  OAI21_X1 U6246 ( .B1(n5046), .B2(n6269), .A(n5045), .ZN(U2985) );
  OAI21_X1 U6247 ( .B1(n5047), .B2(n5048), .A(n5049), .ZN(n6340) );
  INV_X1 U6248 ( .A(n5050), .ZN(n6153) );
  AOI22_X1 U6249 ( .A1(n6263), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .B1(n6351), 
        .B2(REIP_REG_4__SCAN_IN), .ZN(n5051) );
  OAI21_X1 U6250 ( .B1(n6281), .B2(n6153), .A(n5051), .ZN(n5052) );
  AOI21_X1 U6251 ( .B1(n5053), .B2(n5749), .A(n5052), .ZN(n5054) );
  OAI21_X1 U6252 ( .B1(n6269), .B2(n6340), .A(n5054), .ZN(U2982) );
  OAI21_X1 U6253 ( .B1(n5056), .B2(n5057), .A(n5058), .ZN(n6331) );
  INV_X1 U6254 ( .A(n5059), .ZN(n5064) );
  INV_X1 U6255 ( .A(n5060), .ZN(n5062) );
  AOI22_X1 U6256 ( .A1(n6263), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .B1(n6351), 
        .B2(REIP_REG_5__SCAN_IN), .ZN(n5061) );
  OAI21_X1 U6257 ( .B1(n6281), .B2(n5062), .A(n5061), .ZN(n5063) );
  AOI21_X1 U6258 ( .B1(n5064), .B2(n5749), .A(n5063), .ZN(n5065) );
  OAI21_X1 U6259 ( .B1(n6269), .B2(n6331), .A(n5065), .ZN(U2981) );
  OAI21_X1 U6260 ( .B1(n5066), .B2(n5069), .A(n5068), .ZN(n6319) );
  NAND2_X1 U6261 ( .A1(n6351), .A2(REIP_REG_7__SCAN_IN), .ZN(n6316) );
  NAND2_X1 U6262 ( .A1(n6263), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5070)
         );
  OAI211_X1 U6263 ( .C1(n6281), .C2(n5071), .A(n6316), .B(n5070), .ZN(n5072)
         );
  AOI21_X1 U6264 ( .B1(n5073), .B2(n5749), .A(n5072), .ZN(n5074) );
  OAI21_X1 U6265 ( .B1(n6319), .B2(n6269), .A(n5074), .ZN(U2979) );
  NAND2_X1 U6266 ( .A1(n5084), .A2(n6460), .ZN(n5075) );
  AOI21_X1 U6267 ( .B1(n5075), .B2(STATEBS16_REG_SCAN_IN), .A(n5875), .ZN(
        n5082) );
  AOI22_X1 U6268 ( .A1(n5082), .A2(n5079), .B1(n5887), .B2(n5076), .ZN(n5112)
         );
  NOR2_X1 U6269 ( .A1(n5078), .A2(n5077), .ZN(n5883) );
  INV_X1 U6270 ( .A(n5079), .ZN(n5081) );
  OR2_X1 U6271 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5080), .ZN(n5107)
         );
  AOI22_X1 U6272 ( .A1(n5082), .A2(n5081), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n5107), .ZN(n5083) );
  OAI211_X1 U6273 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6498), .A(n5883), .B(n5083), .ZN(n5106) );
  NAND2_X1 U6274 ( .A1(n5106), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n5087)
         );
  OAI22_X1 U6275 ( .A1(n6460), .A2(n6437), .B1(n6440), .B2(n5107), .ZN(n5085)
         );
  AOI21_X1 U6276 ( .B1(n5109), .B2(n6401), .A(n5085), .ZN(n5086) );
  OAI211_X1 U6277 ( .C1(n5112), .C2(n5913), .A(n5087), .B(n5086), .ZN(U3104)
         );
  NAND2_X1 U6278 ( .A1(n5106), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n5090)
         );
  OAI22_X1 U6279 ( .A1(n6460), .A2(n6409), .B1(n5919), .B2(n5107), .ZN(n5088)
         );
  AOI21_X1 U6280 ( .B1(n5109), .B2(n6406), .A(n5088), .ZN(n5089) );
  OAI211_X1 U6281 ( .C1(n5112), .C2(n5918), .A(n5090), .B(n5089), .ZN(U3105)
         );
  NAND2_X1 U6282 ( .A1(n5106), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5093)
         );
  OAI22_X1 U6283 ( .A1(n6460), .A2(n6415), .B1(n5926), .B2(n5107), .ZN(n5091)
         );
  AOI21_X1 U6284 ( .B1(n5109), .B2(n6412), .A(n5091), .ZN(n5092) );
  OAI211_X1 U6285 ( .C1(n5112), .C2(n5925), .A(n5093), .B(n5092), .ZN(U3106)
         );
  NAND2_X1 U6286 ( .A1(n5106), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n5096)
         );
  OAI22_X1 U6287 ( .A1(n6460), .A2(n6425), .B1(n5936), .B2(n5107), .ZN(n5094)
         );
  AOI21_X1 U6288 ( .B1(n5109), .B2(n6421), .A(n5094), .ZN(n5095) );
  OAI211_X1 U6289 ( .C1(n5112), .C2(n5933), .A(n5096), .B(n5095), .ZN(U3107)
         );
  NAND2_X1 U6290 ( .A1(n5106), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n5099)
         );
  OAI22_X1 U6291 ( .A1(n6460), .A2(n6430), .B1(n6431), .B2(n5107), .ZN(n5097)
         );
  AOI21_X1 U6292 ( .B1(n5109), .B2(n6397), .A(n5097), .ZN(n5098) );
  OAI211_X1 U6293 ( .C1(n5112), .C2(n5908), .A(n5099), .B(n5098), .ZN(U3103)
         );
  NAND2_X1 U6294 ( .A1(n5106), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n5102)
         );
  OAI22_X1 U6295 ( .A1(n6460), .A2(n6452), .B1(n6451), .B2(n5107), .ZN(n5100)
         );
  AOI21_X1 U6296 ( .B1(n5109), .B2(n6381), .A(n5100), .ZN(n5101) );
  OAI211_X1 U6297 ( .C1(n5112), .C2(n5889), .A(n5102), .B(n5101), .ZN(U3100)
         );
  NAND2_X1 U6298 ( .A1(n5106), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n5105)
         );
  OAI22_X1 U6299 ( .A1(n6460), .A2(n6389), .B1(n5895), .B2(n5107), .ZN(n5103)
         );
  AOI21_X1 U6300 ( .B1(n5109), .B2(n6386), .A(n5103), .ZN(n5104) );
  OAI211_X1 U6301 ( .C1(n5112), .C2(n5894), .A(n5105), .B(n5104), .ZN(U3101)
         );
  NAND2_X1 U6302 ( .A1(n5106), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5111)
         );
  OAI22_X1 U6303 ( .A1(n6460), .A2(n6395), .B1(n5902), .B2(n5107), .ZN(n5108)
         );
  AOI21_X1 U6304 ( .B1(n5109), .B2(n6392), .A(n5108), .ZN(n5110) );
  OAI211_X1 U6305 ( .C1(n5112), .C2(n5901), .A(n5111), .B(n5110), .ZN(U3102)
         );
  AOI22_X1 U6306 ( .A1(n6303), .A2(n6203), .B1(EBX_REG_9__SCAN_IN), .B2(n5617), 
        .ZN(n5113) );
  OAI21_X1 U6307 ( .B1(n5146), .B2(n5639), .A(n5113), .ZN(U2850) );
  AOI22_X1 U6308 ( .A1(n5663), .A2(DATAI_9_), .B1(n6217), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n5114) );
  OAI21_X1 U6309 ( .B1(n5146), .B2(n5983), .A(n5114), .ZN(U2882) );
  OAI21_X1 U6310 ( .B1(n6184), .B2(n6160), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5115) );
  OAI21_X1 U6311 ( .B1(n6140), .B2(n5116), .A(n5115), .ZN(n5117) );
  AOI21_X1 U6312 ( .B1(n6122), .B2(n5118), .A(n5117), .ZN(n5121) );
  NAND2_X1 U6313 ( .A1(n6609), .A2(n5119), .ZN(n6151) );
  INV_X1 U6314 ( .A(n6151), .ZN(n6192) );
  AOI22_X1 U6315 ( .A1(n3808), .A2(n6192), .B1(n6178), .B2(REIP_REG_0__SCAN_IN), .ZN(n5120) );
  OAI211_X1 U6316 ( .C1(n5122), .C2(n6188), .A(n5121), .B(n5120), .ZN(U2827)
         );
  AND2_X1 U6317 ( .A1(n5124), .A2(n5123), .ZN(n5125) );
  NOR2_X1 U6318 ( .A1(n4197), .A2(n5125), .ZN(n5153) );
  INV_X1 U6319 ( .A(n5153), .ZN(n5127) );
  AOI22_X1 U6320 ( .A1(n5663), .A2(DATAI_8_), .B1(n6217), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n5126) );
  OAI21_X1 U6321 ( .B1(n5127), .B2(n5983), .A(n5126), .ZN(U2883) );
  OAI21_X1 U6322 ( .B1(n4196), .B2(n5129), .A(n5184), .ZN(n6130) );
  AOI22_X1 U6323 ( .A1(n5663), .A2(DATAI_10_), .B1(n6217), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n5130) );
  OAI21_X1 U6324 ( .B1(n6130), .B2(n5983), .A(n5130), .ZN(U2881) );
  XNOR2_X1 U6325 ( .A(n5131), .B(n6113), .ZN(n6293) );
  AOI22_X1 U6326 ( .A1(n6293), .A2(n6203), .B1(EBX_REG_10__SCAN_IN), .B2(n5617), .ZN(n5132) );
  OAI21_X1 U6327 ( .B1(n6130), .B2(n5639), .A(n5132), .ZN(U2849) );
  INV_X1 U6328 ( .A(n5639), .ZN(n6204) );
  OR2_X1 U6329 ( .A1(n5134), .A2(n5133), .ZN(n5135) );
  NAND2_X1 U6330 ( .A1(n5136), .A2(n5135), .ZN(n6310) );
  OAI22_X1 U6331 ( .A1(n6310), .A2(n5637), .B1(n5157), .B2(n6207), .ZN(n5137)
         );
  AOI21_X1 U6332 ( .B1(n5153), .B2(n6204), .A(n5137), .ZN(n5138) );
  INV_X1 U6333 ( .A(n5138), .ZN(U2851) );
  XNOR2_X1 U6334 ( .A(n6249), .B(n5140), .ZN(n5141) );
  XNOR2_X1 U6335 ( .A(n5139), .B(n5141), .ZN(n6305) );
  NAND2_X1 U6336 ( .A1(n6305), .A2(n6276), .ZN(n5145) );
  NAND2_X1 U6337 ( .A1(n6351), .A2(REIP_REG_9__SCAN_IN), .ZN(n6301) );
  OAI21_X1 U6338 ( .B1(n5755), .B2(n4188), .A(n6301), .ZN(n5142) );
  AOI21_X1 U6339 ( .B1(n6253), .B2(n5143), .A(n5142), .ZN(n5144) );
  OAI211_X1 U6340 ( .C1(n6267), .C2(n5146), .A(n5145), .B(n5144), .ZN(U2977)
         );
  OAI21_X1 U6341 ( .B1(n5147), .B2(n5149), .A(n5148), .ZN(n6309) );
  AOI22_X1 U6342 ( .A1(n6263), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n6351), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n5150) );
  OAI21_X1 U6343 ( .B1(n6281), .B2(n5159), .A(n5150), .ZN(n5151) );
  AOI21_X1 U6344 ( .B1(n5153), .B2(n5749), .A(n5151), .ZN(n5152) );
  OAI21_X1 U6345 ( .B1(n6309), .B2(n6269), .A(n5152), .ZN(U2978) );
  NAND2_X1 U6346 ( .A1(n5153), .A2(n6146), .ZN(n5164) );
  INV_X1 U6347 ( .A(n5154), .ZN(n5156) );
  NOR3_X1 U6348 ( .A1(n6176), .A2(n5156), .A3(n5155), .ZN(n5162) );
  OAI22_X1 U6349 ( .A1(n5157), .A2(n6140), .B1(n6197), .B2(n6310), .ZN(n5161)
         );
  INV_X1 U6350 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5158) );
  OAI22_X1 U6351 ( .A1(n5159), .A2(n6187), .B1(n6138), .B2(n5158), .ZN(n5160)
         );
  NOR4_X1 U6352 ( .A1(n5162), .A2(n6351), .A3(n5161), .A4(n5160), .ZN(n5163)
         );
  OAI211_X1 U6353 ( .C1(n6548), .C2(n6136), .A(n5164), .B(n5163), .ZN(U2819)
         );
  AOI22_X1 U6354 ( .A1(n6243), .A2(UWORD_REG_7__SCAN_IN), .B1(n6235), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n5165) );
  OAI21_X1 U6355 ( .B1(n4398), .B2(n5176), .A(n5165), .ZN(U2900) );
  AOI22_X1 U6356 ( .A1(n6243), .A2(UWORD_REG_2__SCAN_IN), .B1(n6235), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n5166) );
  OAI21_X1 U6357 ( .B1(n4412), .B2(n5176), .A(n5166), .ZN(U2905) );
  AOI22_X1 U6358 ( .A1(n6243), .A2(UWORD_REG_1__SCAN_IN), .B1(n6235), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n5167) );
  OAI21_X1 U6359 ( .B1(n4421), .B2(n5176), .A(n5167), .ZN(U2906) );
  INV_X1 U6360 ( .A(EAX_REG_16__SCAN_IN), .ZN(n5169) );
  AOI22_X1 U6361 ( .A1(n6243), .A2(UWORD_REG_0__SCAN_IN), .B1(n6235), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n5168) );
  OAI21_X1 U6362 ( .B1(n5169), .B2(n5176), .A(n5168), .ZN(U2907) );
  AOI22_X1 U6363 ( .A1(n6243), .A2(UWORD_REG_4__SCAN_IN), .B1(n6235), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n5170) );
  OAI21_X1 U6364 ( .B1(n4407), .B2(n5176), .A(n5170), .ZN(U2903) );
  INV_X1 U6365 ( .A(EAX_REG_19__SCAN_IN), .ZN(n5172) );
  AOI22_X1 U6366 ( .A1(n6243), .A2(UWORD_REG_3__SCAN_IN), .B1(n6235), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n5171) );
  OAI21_X1 U6367 ( .B1(n5172), .B2(n5176), .A(n5171), .ZN(U2904) );
  AOI22_X1 U6368 ( .A1(n6243), .A2(UWORD_REG_6__SCAN_IN), .B1(n6235), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n5173) );
  OAI21_X1 U6369 ( .B1(n5174), .B2(n5176), .A(n5173), .ZN(U2901) );
  AOI22_X1 U6370 ( .A1(n6243), .A2(UWORD_REG_5__SCAN_IN), .B1(n6235), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n5175) );
  OAI21_X1 U6371 ( .B1(n4386), .B2(n5176), .A(n5175), .ZN(U2902) );
  NAND2_X1 U6372 ( .A1(n6248), .A2(n5178), .ZN(n5179) );
  XNOR2_X1 U6373 ( .A(n5177), .B(n5179), .ZN(n6297) );
  NAND2_X1 U6374 ( .A1(n6297), .A2(n6276), .ZN(n5182) );
  NAND2_X1 U6375 ( .A1(n6351), .A2(REIP_REG_10__SCAN_IN), .ZN(n6291) );
  OAI21_X1 U6376 ( .B1(n5755), .B2(n6124), .A(n6291), .ZN(n5180) );
  AOI21_X1 U6377 ( .B1(n6132), .B2(n6253), .A(n5180), .ZN(n5181) );
  OAI211_X1 U6378 ( .C1(n6267), .C2(n6130), .A(n5182), .B(n5181), .ZN(U2976)
         );
  INV_X1 U6379 ( .A(n5183), .ZN(n5188) );
  AOI21_X1 U6380 ( .B1(n5185), .B2(n5184), .A(n5183), .ZN(n6254) );
  INV_X1 U6381 ( .A(n6254), .ZN(n5187) );
  AOI22_X1 U6382 ( .A1(n5663), .A2(DATAI_11_), .B1(n6217), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n5186) );
  OAI21_X1 U6383 ( .B1(n5187), .B2(n5983), .A(n5186), .ZN(U2880) );
  XOR2_X1 U6384 ( .A(n5189), .B(n5188), .Z(n5214) );
  INV_X1 U6385 ( .A(n5214), .ZN(n6105) );
  AOI22_X1 U6386 ( .A1(n5663), .A2(DATAI_12_), .B1(n6217), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n5190) );
  OAI21_X1 U6387 ( .B1(n6105), .B2(n5983), .A(n5190), .ZN(U2879) );
  INV_X1 U6388 ( .A(n5192), .ZN(n5193) );
  NOR2_X1 U6389 ( .A1(n5194), .A2(n5193), .ZN(n5195) );
  XNOR2_X1 U6390 ( .A(n5191), .B(n5195), .ZN(n5216) );
  INV_X1 U6391 ( .A(n5196), .ZN(n5197) );
  AOI21_X1 U6392 ( .B1(n6339), .B2(n6289), .A(n5197), .ZN(n5198) );
  OAI21_X1 U6393 ( .B1(n5200), .B2(n5199), .A(n5198), .ZN(n6294) );
  AOI21_X1 U6394 ( .B1(n5829), .B2(n5201), .A(n6294), .ZN(n6287) );
  AOI211_X1 U6395 ( .C1(n6287), .C2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(n5203), .B(n5202), .ZN(n5208) );
  NOR3_X1 U6396 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n6288), .A3(n3512), 
        .ZN(n5207) );
  NOR2_X1 U6397 ( .A1(n6115), .A2(n5204), .ZN(n5205) );
  OR2_X1 U6398 ( .A1(n6030), .A2(n5205), .ZN(n6110) );
  NAND2_X1 U6399 ( .A1(n6351), .A2(REIP_REG_12__SCAN_IN), .ZN(n5211) );
  OAI21_X1 U6400 ( .B1(n6110), .B2(n6342), .A(n5211), .ZN(n5206) );
  NOR3_X1 U6401 ( .A1(n5208), .A2(n5207), .A3(n5206), .ZN(n5209) );
  OAI21_X1 U6402 ( .B1(n5216), .B2(n6283), .A(n5209), .ZN(U3006) );
  INV_X1 U6403 ( .A(n6107), .ZN(n5212) );
  NAND2_X1 U6404 ( .A1(n6263), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5210)
         );
  OAI211_X1 U6405 ( .C1(n6281), .C2(n5212), .A(n5211), .B(n5210), .ZN(n5213)
         );
  AOI21_X1 U6406 ( .B1(n5214), .B2(n5749), .A(n5213), .ZN(n5215) );
  OAI21_X1 U6407 ( .B1(n5216), .B2(n6269), .A(n5215), .ZN(U2974) );
  INV_X1 U6408 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5217) );
  OAI222_X1 U6409 ( .A1(n6110), .A2(n5637), .B1(n6207), .B2(n5217), .C1(n5639), 
        .C2(n6105), .ZN(U2847) );
  XNOR2_X1 U6410 ( .A(n6249), .B(n5219), .ZN(n5220) );
  XNOR2_X1 U6411 ( .A(n5218), .B(n5220), .ZN(n5759) );
  NOR3_X1 U6412 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5221), .A3(n6026), 
        .ZN(n6034) );
  AOI21_X1 U6413 ( .B1(n5222), .B2(n6026), .A(n6034), .ZN(n5223) );
  OAI211_X1 U6414 ( .C1(n5226), .C2(n5224), .A(n6287), .B(n5223), .ZN(n6033)
         );
  XNOR2_X1 U6415 ( .A(n5225), .B(n5575), .ZN(n6083) );
  INV_X1 U6416 ( .A(n6083), .ZN(n5636) );
  NOR2_X1 U6417 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n6288), .ZN(n5227)
         );
  NAND2_X1 U6418 ( .A1(n5227), .A2(n5226), .ZN(n5228) );
  NAND2_X1 U6419 ( .A1(n6351), .A2(REIP_REG_14__SCAN_IN), .ZN(n5753) );
  OAI211_X1 U6420 ( .C1(n5636), .C2(n6342), .A(n5228), .B(n5753), .ZN(n5229)
         );
  AOI21_X1 U6421 ( .B1(n6033), .B2(INSTADDRPOINTER_REG_14__SCAN_IN), .A(n5229), 
        .ZN(n5230) );
  OAI21_X1 U6422 ( .B1(n5759), .B2(n6283), .A(n5230), .ZN(U3004) );
  NAND2_X1 U6423 ( .A1(n5232), .A2(n5231), .ZN(n5233) );
  AND2_X1 U6424 ( .A1(n5234), .A2(n5233), .ZN(n6199) );
  INV_X1 U6425 ( .A(n6199), .ZN(n5236) );
  AOI22_X1 U6426 ( .A1(n5663), .A2(DATAI_13_), .B1(n6217), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n5235) );
  OAI21_X1 U6427 ( .B1(n5236), .B2(n5983), .A(n5235), .ZN(U2878) );
  INV_X1 U6428 ( .A(n5240), .ZN(n5242) );
  INV_X1 U6429 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5241) );
  NAND2_X1 U6430 ( .A1(n5242), .A2(n5241), .ZN(n5243) );
  NAND2_X1 U6431 ( .A1(n5337), .A2(n5243), .ZN(n5684) );
  AOI22_X1 U6432 ( .A1(n5340), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n5247) );
  AOI22_X1 U6433 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n5349), .B1(n5348), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5246) );
  AOI22_X1 U6434 ( .A1(n5343), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3212), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n5245) );
  AOI22_X1 U6435 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n2990), .B1(n3004), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5244) );
  NAND4_X1 U6436 ( .A1(n5247), .A2(n5246), .A3(n5245), .A4(n5244), .ZN(n5253)
         );
  AOI22_X1 U6437 ( .A1(n4119), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3005), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5251) );
  AOI22_X1 U6438 ( .A1(n3207), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3329), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5250) );
  AOI22_X1 U6439 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n3011), .B1(n3391), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n5249) );
  AOI22_X1 U6440 ( .A1(n5258), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n5326), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n5248) );
  NAND4_X1 U6441 ( .A1(n5251), .A2(n5250), .A3(n5249), .A4(n5248), .ZN(n5252)
         );
  NOR2_X1 U6442 ( .A1(n5253), .A2(n5252), .ZN(n5291) );
  AOI22_X1 U6443 ( .A1(n4108), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3190), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5257) );
  AOI22_X1 U6444 ( .A1(n5340), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n5348), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5256) );
  AOI22_X1 U6445 ( .A1(n4119), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3012), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n5255) );
  AOI22_X1 U6446 ( .A1(n5349), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3003), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5254) );
  NAND4_X1 U6447 ( .A1(n5257), .A2(n5256), .A3(n5255), .A4(n5254), .ZN(n5264)
         );
  AOI22_X1 U6448 ( .A1(n3010), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3017), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n5262) );
  AOI22_X1 U6449 ( .A1(n3391), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n5350), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5261) );
  AOI22_X1 U6450 ( .A1(n5258), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n5326), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n5260) );
  AOI22_X1 U6451 ( .A1(n3382), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n5259) );
  NAND4_X1 U6452 ( .A1(n5262), .A2(n5261), .A3(n5260), .A4(n5259), .ZN(n5263)
         );
  NOR2_X1 U6453 ( .A1(n5264), .A2(n5263), .ZN(n5309) );
  NAND2_X1 U6454 ( .A1(n5266), .A2(n5265), .ZN(n5308) );
  NOR2_X1 U6455 ( .A1(n5309), .A2(n5308), .ZN(n5303) );
  AOI22_X1 U6456 ( .A1(n4108), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3005), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5270) );
  AOI22_X1 U6457 ( .A1(n5340), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n5348), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5269) );
  AOI22_X1 U6458 ( .A1(n4119), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n5268) );
  AOI22_X1 U6459 ( .A1(n5349), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3003), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5267) );
  NAND4_X1 U6460 ( .A1(n5270), .A2(n5269), .A3(n5268), .A4(n5267), .ZN(n5276)
         );
  AOI22_X1 U6461 ( .A1(n3011), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3017), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n5274) );
  AOI22_X1 U6462 ( .A1(n3391), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n5350), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n5273) );
  AOI22_X1 U6463 ( .A1(n5258), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n5326), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n5272) );
  AOI22_X1 U6464 ( .A1(n3329), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3212), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n5271) );
  NAND4_X1 U6465 ( .A1(n5274), .A2(n5273), .A3(n5272), .A4(n5271), .ZN(n5275)
         );
  OR2_X1 U6466 ( .A1(n5276), .A2(n5275), .ZN(n5302) );
  NAND2_X1 U6467 ( .A1(n5303), .A2(n5302), .ZN(n5292) );
  NOR2_X1 U6468 ( .A1(n5291), .A2(n5292), .ZN(n5321) );
  AOI22_X1 U6469 ( .A1(n4108), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3005), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5280) );
  AOI22_X1 U6470 ( .A1(n5340), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n5348), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5279) );
  AOI22_X1 U6471 ( .A1(n4119), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3012), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n5278) );
  AOI22_X1 U6472 ( .A1(n5349), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3003), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5277) );
  NAND4_X1 U6473 ( .A1(n5280), .A2(n5279), .A3(n5278), .A4(n5277), .ZN(n5286)
         );
  AOI22_X1 U6474 ( .A1(n3010), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3017), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n5284) );
  AOI22_X1 U6475 ( .A1(n3008), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3004), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5283) );
  AOI22_X1 U6476 ( .A1(n5258), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n5326), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n5282) );
  AOI22_X1 U6477 ( .A1(n3329), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3212), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n5281) );
  NAND4_X1 U6478 ( .A1(n5284), .A2(n5283), .A3(n5282), .A4(n5281), .ZN(n5285)
         );
  OR2_X1 U6479 ( .A1(n5286), .A2(n5285), .ZN(n5320) );
  XNOR2_X1 U6480 ( .A(n5321), .B(n5320), .ZN(n5289) );
  AOI21_X1 U6481 ( .B1(PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6498), .A(n5369), 
        .ZN(n5288) );
  NAND2_X1 U6482 ( .A1(n5364), .A2(EAX_REG_28__SCAN_IN), .ZN(n5287) );
  OAI211_X1 U6483 ( .C1(n5289), .C2(n5366), .A(n5288), .B(n5287), .ZN(n5290)
         );
  OAI21_X1 U6484 ( .B1(n5362), .B2(n5684), .A(n5290), .ZN(n5485) );
  INV_X1 U6485 ( .A(n5485), .ZN(n5319) );
  XOR2_X1 U6486 ( .A(n5292), .B(n5291), .Z(n5293) );
  NAND2_X1 U6487 ( .A1(n5293), .A2(n5333), .ZN(n5296) );
  INV_X1 U6488 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5504) );
  NOR2_X1 U6489 ( .A1(n5504), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5294) );
  AOI211_X1 U6490 ( .C1(n5364), .C2(EAX_REG_27__SCAN_IN), .A(n5369), .B(n5294), 
        .ZN(n5295) );
  XNOR2_X1 U6491 ( .A(n5301), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5503)
         );
  AOI22_X1 U6492 ( .A1(n5296), .A2(n5295), .B1(n5369), .B2(n5503), .ZN(n5499)
         );
  INV_X1 U6493 ( .A(n5297), .ZN(n5299) );
  INV_X1 U6494 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5298) );
  NAND2_X1 U6495 ( .A1(n5299), .A2(n5298), .ZN(n5300) );
  NAND2_X1 U6496 ( .A1(n5301), .A2(n5300), .ZN(n5702) );
  XNOR2_X1 U6497 ( .A(n5303), .B(n5302), .ZN(n5306) );
  AOI21_X1 U6498 ( .B1(PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n6498), .A(n5369), 
        .ZN(n5305) );
  NAND2_X1 U6499 ( .A1(n3809), .A2(EAX_REG_26__SCAN_IN), .ZN(n5304) );
  OAI211_X1 U6500 ( .C1(n5306), .C2(n5366), .A(n5305), .B(n5304), .ZN(n5307)
         );
  OAI21_X1 U6501 ( .B1(n5362), .B2(n5702), .A(n5307), .ZN(n5514) );
  INV_X1 U6502 ( .A(n5514), .ZN(n5318) );
  XOR2_X1 U6503 ( .A(n5309), .B(n5308), .Z(n5310) );
  NAND2_X1 U6504 ( .A1(n5310), .A2(n5333), .ZN(n5317) );
  NAND2_X1 U6505 ( .A1(n6498), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5311)
         );
  NAND2_X1 U6506 ( .A1(n5362), .A2(n5311), .ZN(n5312) );
  AOI21_X1 U6507 ( .B1(n3809), .B2(EAX_REG_25__SCAN_IN), .A(n5312), .ZN(n5316)
         );
  INV_X1 U6508 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5313) );
  XNOR2_X1 U6509 ( .A(n5314), .B(n5313), .ZN(n5945) );
  AND2_X1 U6510 ( .A1(n5945), .A2(n5369), .ZN(n5315) );
  AOI21_X1 U6511 ( .B1(n5317), .B2(n5316), .A(n5315), .ZN(n5592) );
  AND2_X1 U6512 ( .A1(n5318), .A2(n5592), .ZN(n5497) );
  AND2_X1 U6513 ( .A1(n5499), .A2(n5497), .ZN(n5483) );
  NAND2_X1 U6514 ( .A1(n5321), .A2(n5320), .ZN(n5357) );
  AOI22_X1 U6515 ( .A1(n4108), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3005), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5325) );
  AOI22_X1 U6516 ( .A1(n5348), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3012), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n5324) );
  AOI22_X1 U6517 ( .A1(n5349), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3003), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5323) );
  AOI22_X1 U6518 ( .A1(n3011), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n5322) );
  NAND4_X1 U6519 ( .A1(n5325), .A2(n5324), .A3(n5323), .A4(n5322), .ZN(n5332)
         );
  AOI22_X1 U6520 ( .A1(n5340), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5330) );
  AOI22_X1 U6521 ( .A1(n3329), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n2990), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n5329) );
  AOI22_X1 U6522 ( .A1(n3008), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3004), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5328) );
  AOI22_X1 U6523 ( .A1(n5258), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n5326), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n5327) );
  NAND4_X1 U6524 ( .A1(n5330), .A2(n5329), .A3(n5328), .A4(n5327), .ZN(n5331)
         );
  NOR2_X1 U6525 ( .A1(n5332), .A2(n5331), .ZN(n5358) );
  XOR2_X1 U6526 ( .A(n5357), .B(n5358), .Z(n5334) );
  NAND2_X1 U6527 ( .A1(n5334), .A2(n5333), .ZN(n5339) );
  NOR2_X1 U6528 ( .A1(n5335), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5336) );
  AOI211_X1 U6529 ( .C1(n5364), .C2(EAX_REG_29__SCAN_IN), .A(n5369), .B(n5336), 
        .ZN(n5338) );
  XNOR2_X1 U6530 ( .A(n5337), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5670)
         );
  AOI22_X1 U6531 ( .A1(n5339), .A2(n5338), .B1(n5369), .B2(n5670), .ZN(n5431)
         );
  AOI22_X1 U6532 ( .A1(n5340), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n5347) );
  AOI22_X1 U6533 ( .A1(n3010), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n2990), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n5346) );
  AOI22_X1 U6534 ( .A1(n3008), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n5258), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n5345) );
  AOI22_X1 U6535 ( .A1(n3329), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5343), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5344) );
  NAND4_X1 U6536 ( .A1(n5347), .A2(n5346), .A3(n5345), .A4(n5344), .ZN(n5356)
         );
  AOI22_X1 U6537 ( .A1(n3190), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n5348), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5354) );
  AOI22_X1 U6538 ( .A1(n4119), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3012), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n5353) );
  AOI22_X1 U6539 ( .A1(n5349), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n5352) );
  AOI22_X1 U6540 ( .A1(n3004), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n5326), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n5351) );
  NAND4_X1 U6541 ( .A1(n5354), .A2(n5353), .A3(n5352), .A4(n5351), .ZN(n5355)
         );
  NOR2_X1 U6542 ( .A1(n5356), .A2(n5355), .ZN(n5360) );
  NOR2_X1 U6543 ( .A1(n5358), .A2(n5357), .ZN(n5359) );
  XOR2_X1 U6544 ( .A(n5360), .B(n5359), .Z(n5367) );
  NAND2_X1 U6545 ( .A1(n6498), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5361)
         );
  NAND2_X1 U6546 ( .A1(n5362), .A2(n5361), .ZN(n5363) );
  AOI21_X1 U6547 ( .B1(n5364), .B2(EAX_REG_30__SCAN_IN), .A(n5363), .ZN(n5365)
         );
  OAI21_X1 U6548 ( .B1(n5367), .B2(n5366), .A(n5365), .ZN(n5371) );
  XNOR2_X1 U6549 ( .A(n5368), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5474)
         );
  NAND2_X1 U6550 ( .A1(n5474), .A2(n5369), .ZN(n5370) );
  INV_X1 U6551 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5477) );
  INV_X1 U6552 ( .A(n5479), .ZN(n5372) );
  OAI222_X1 U6553 ( .A1(n5639), .A2(n5647), .B1(n5477), .B2(n6207), .C1(n5637), 
        .C2(n5372), .ZN(U2829) );
  NAND2_X1 U6554 ( .A1(n4339), .A2(n5373), .ZN(n5377) );
  INV_X1 U6555 ( .A(n4248), .ZN(n5374) );
  NAND3_X1 U6556 ( .A1(n5375), .A2(n5374), .A3(n5379), .ZN(n5376) );
  OAI211_X1 U6557 ( .C1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n6462), .A(n5377), .B(n5376), .ZN(n6466) );
  AOI222_X1 U6558 ( .A1(n6466), .A2(n6593), .B1(n5381), .B2(n5380), .C1(n5379), 
        .C2(n5378), .ZN(n5383) );
  NAND2_X1 U6559 ( .A1(n5384), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5382) );
  OAI21_X1 U6560 ( .B1(n5384), .B2(n5383), .A(n5382), .ZN(U3460) );
  INV_X1 U6561 ( .A(n5385), .ZN(n5391) );
  NAND2_X1 U6562 ( .A1(n3789), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5388) );
  INV_X1 U6563 ( .A(n5388), .ZN(n5390) );
  AND2_X1 U6564 ( .A1(n5388), .A2(n5387), .ZN(n5389) );
  OAI22_X1 U6565 ( .A1(n5391), .A2(n5390), .B1(n5386), .B2(n5389), .ZN(n6013)
         );
  INV_X1 U6566 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5392) );
  OAI22_X1 U6567 ( .A1(n5755), .A2(n5392), .B1(n6341), .B2(n6562), .ZN(n5398)
         );
  OR2_X1 U6568 ( .A1(n5393), .A2(n5571), .ZN(n5569) );
  AND2_X1 U6569 ( .A1(n5569), .A2(n5394), .ZN(n5396) );
  OR2_X1 U6570 ( .A1(n5396), .A2(n5395), .ZN(n6077) );
  NOR2_X1 U6571 ( .A1(n6077), .A2(n6267), .ZN(n5397) );
  AOI211_X1 U6572 ( .C1(n6253), .C2(n6078), .A(n5398), .B(n5397), .ZN(n5399)
         );
  OAI21_X1 U6573 ( .B1(n6013), .B2(n6269), .A(n5399), .ZN(U2970) );
  OAI21_X1 U6574 ( .B1(n5806), .B2(n5401), .A(n5400), .ZN(n5402) );
  AND2_X1 U6575 ( .A1(n5402), .A2(n5597), .ZN(n5960) );
  INV_X1 U6576 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5405) );
  INV_X1 U6577 ( .A(n5799), .ZN(n5404) );
  AOI211_X1 U6578 ( .C1(n5406), .C2(n5405), .A(n5404), .B(n5403), .ZN(n5407)
         );
  AOI211_X1 U6579 ( .C1(n6353), .C2(n5960), .A(n5408), .B(n5407), .ZN(n5409)
         );
  OAI21_X1 U6580 ( .B1(n5410), .B2(n6283), .A(n5409), .ZN(U2994) );
  AND2_X1 U6581 ( .A1(n3075), .A2(n5411), .ZN(n5412) );
  AOI22_X1 U6582 ( .A1(n3809), .A2(EAX_REG_31__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n5413), .ZN(n5414) );
  AOI21_X1 U6583 ( .B1(n6263), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5416), 
        .ZN(n5417) );
  OAI21_X1 U6584 ( .B1(n6281), .B2(n5418), .A(n5417), .ZN(n5419) );
  AOI21_X1 U6585 ( .B1(n5642), .B2(n5749), .A(n5419), .ZN(n5420) );
  OAI21_X1 U6586 ( .B1(n5421), .B2(n6269), .A(n5420), .ZN(U2955) );
  INV_X1 U6587 ( .A(n5474), .ZN(n5424) );
  AOI21_X1 U6588 ( .B1(n6263), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n5422), 
        .ZN(n5423) );
  OAI21_X1 U6589 ( .B1(n6281), .B2(n5424), .A(n5423), .ZN(n5425) );
  AOI21_X1 U6590 ( .B1(n5426), .B2(n5749), .A(n5425), .ZN(n5427) );
  OAI21_X1 U6591 ( .B1(n5428), .B2(n6269), .A(n5427), .ZN(U2956) );
  OAI21_X1 U6592 ( .B1(n5434), .B2(n5433), .A(n5432), .ZN(n5458) );
  INV_X1 U6593 ( .A(n5458), .ZN(n5763) );
  AOI22_X1 U6594 ( .A1(PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n6184), .B1(n6160), 
        .B2(n5670), .ZN(n5435) );
  OAI21_X1 U6595 ( .B1(n6140), .B2(n5459), .A(n5435), .ZN(n5450) );
  INV_X1 U6596 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6713) );
  INV_X1 U6597 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6682) );
  INV_X1 U6598 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6565) );
  OR3_X1 U6599 ( .A1(n6713), .A2(n6682), .A3(n6565), .ZN(n5440) );
  NAND4_X1 U6600 ( .A1(REIP_REG_11__SCAN_IN), .A2(n5436), .A3(
        REIP_REG_10__SCAN_IN), .A4(REIP_REG_9__SCAN_IN), .ZN(n6095) );
  NAND2_X1 U6601 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .ZN(
        n6093) );
  NOR2_X1 U6602 ( .A1(n6095), .A2(n6093), .ZN(n6085) );
  NAND2_X1 U6603 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6085), .ZN(n5437) );
  NAND4_X1 U6604 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .A4(n6072), .ZN(n6065) );
  NAND3_X1 U6605 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .A3(
        n5971), .ZN(n5524) );
  NAND4_X1 U6606 ( .A1(n5944), .A2(REIP_REG_24__SCAN_IN), .A3(
        REIP_REG_26__SCAN_IN), .A4(REIP_REG_25__SCAN_IN), .ZN(n5500) );
  NAND2_X1 U6607 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n5447) );
  NOR2_X1 U6608 ( .A1(n5500), .A2(n5447), .ZN(n5480) );
  AND2_X1 U6609 ( .A1(n6193), .A2(n5437), .ZN(n6084) );
  INV_X1 U6610 ( .A(n6159), .ZN(n6183) );
  NAND3_X1 U6611 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .ZN(n5438) );
  AND2_X1 U6612 ( .A1(n6193), .A2(n5438), .ZN(n5439) );
  NOR2_X1 U6613 ( .A1(n6082), .A2(n5439), .ZN(n6064) );
  NAND2_X1 U6614 ( .A1(n6193), .A2(n5440), .ZN(n5441) );
  NAND2_X1 U6615 ( .A1(n6064), .A2(n5441), .ZN(n5972) );
  NAND2_X1 U6616 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n5966) );
  INV_X1 U6617 ( .A(n5966), .ZN(n5442) );
  NAND2_X1 U6618 ( .A1(REIP_REG_23__SCAN_IN), .A2(n5442), .ZN(n5443) );
  AND2_X1 U6619 ( .A1(n6178), .A2(n5443), .ZN(n5444) );
  NOR2_X1 U6620 ( .A1(n5972), .A2(n5444), .ZN(n5963) );
  INV_X1 U6621 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6715) );
  INV_X1 U6622 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6650) );
  INV_X1 U6623 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6573) );
  OR3_X1 U6624 ( .A1(n6715), .A2(n6650), .A3(n6573), .ZN(n5445) );
  NAND2_X1 U6625 ( .A1(n6178), .A2(n5445), .ZN(n5446) );
  NAND2_X1 U6626 ( .A1(n5963), .A2(n5446), .ZN(n5511) );
  AND2_X1 U6627 ( .A1(n6193), .A2(n5447), .ZN(n5448) );
  OR2_X1 U6628 ( .A1(n5511), .A2(n5448), .ZN(n5492) );
  MUX2_X1 U6629 ( .A(n5480), .B(n5492), .S(REIP_REG_29__SCAN_IN), .Z(n5449) );
  AOI211_X1 U6630 ( .C1(n6122), .C2(n5763), .A(n5450), .B(n5449), .ZN(n5451)
         );
  OAI21_X1 U6631 ( .B1(n5669), .B2(n6129), .A(n5451), .ZN(U2798) );
  INV_X1 U6632 ( .A(n5452), .ZN(n5453) );
  AOI22_X1 U6633 ( .A1(n6214), .A2(DATAI_29_), .B1(n6217), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5457) );
  AND2_X1 U6634 ( .A1(n3239), .A2(n5454), .ZN(n5455) );
  NAND2_X1 U6635 ( .A1(n6218), .A2(DATAI_13_), .ZN(n5456) );
  OAI211_X1 U6636 ( .C1(n5669), .C2(n5983), .A(n5457), .B(n5456), .ZN(U2862)
         );
  OAI222_X1 U6637 ( .A1(n5639), .A2(n5669), .B1(n5459), .B2(n6207), .C1(n5458), 
        .C2(n5637), .ZN(U2830) );
  INV_X1 U6638 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n6657) );
  NAND2_X1 U6639 ( .A1(n6657), .A2(n5460), .ZN(n5463) );
  INV_X1 U6640 ( .A(n5461), .ZN(n5462) );
  MUX2_X1 U6641 ( .A(n5463), .B(n5462), .S(n6609), .Z(U3474) );
  INV_X1 U6642 ( .A(n5642), .ZN(n5472) );
  INV_X1 U6643 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6767) );
  OR2_X1 U6644 ( .A1(n5492), .A2(n6767), .ZN(n5473) );
  OAI211_X1 U6645 ( .C1(n5473), .C2(n6716), .A(REIP_REG_31__SCAN_IN), .B(n6178), .ZN(n5467) );
  NAND2_X1 U6646 ( .A1(n6184), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5466)
         );
  NAND3_X1 U6647 ( .A1(n6609), .A2(EBX_REG_31__SCAN_IN), .A3(n5464), .ZN(n5465) );
  NAND3_X1 U6648 ( .A1(n5467), .A2(n5466), .A3(n5465), .ZN(n5468) );
  AOI21_X1 U6649 ( .B1(n5583), .B2(n6122), .A(n5468), .ZN(n5471) );
  NAND4_X1 U6650 ( .A1(n5480), .A2(REIP_REG_30__SCAN_IN), .A3(
        REIP_REG_29__SCAN_IN), .A4(n5469), .ZN(n5470) );
  OAI211_X1 U6651 ( .C1(n5472), .C2(n6129), .A(n5471), .B(n5470), .ZN(U2796)
         );
  NAND3_X1 U6652 ( .A1(n5473), .A2(REIP_REG_30__SCAN_IN), .A3(n6178), .ZN(
        n5476) );
  AOI22_X1 U6653 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n6184), .B1(n6160), 
        .B2(n5474), .ZN(n5475) );
  OAI211_X1 U6654 ( .C1(n5477), .C2(n6140), .A(n5476), .B(n5475), .ZN(n5478)
         );
  AOI21_X1 U6655 ( .B1(n5479), .B2(n6122), .A(n5478), .ZN(n5482) );
  NAND3_X1 U6656 ( .A1(n5480), .A2(REIP_REG_29__SCAN_IN), .A3(n6716), .ZN(
        n5481) );
  OAI211_X1 U6657 ( .C1(n5647), .C2(n6129), .A(n5482), .B(n5481), .ZN(U2797)
         );
  NAND2_X1 U6658 ( .A1(n5593), .A2(n5483), .ZN(n5498) );
  AOI21_X1 U6659 ( .B1(n5485), .B2(n5498), .A(n5484), .ZN(n5686) );
  NAND2_X1 U6660 ( .A1(n5486), .A2(n5487), .ZN(n5488) );
  NAND2_X1 U6661 ( .A1(n6182), .A2(EBX_REG_28__SCAN_IN), .ZN(n5491) );
  NAND2_X1 U6662 ( .A1(n6184), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5490)
         );
  OAI211_X1 U6663 ( .C1(n6187), .C2(n5684), .A(n5491), .B(n5490), .ZN(n5495)
         );
  INV_X1 U6664 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6692) );
  NOR2_X1 U6665 ( .A1(n5500), .A2(n6692), .ZN(n5493) );
  MUX2_X1 U6666 ( .A(n5493), .B(n5492), .S(REIP_REG_28__SCAN_IN), .Z(n5494) );
  AOI211_X1 U6667 ( .C1(n6122), .C2(n5773), .A(n5495), .B(n5494), .ZN(n5496)
         );
  OAI21_X1 U6668 ( .B1(n5650), .B2(n6129), .A(n5496), .ZN(U2799) );
  INV_X1 U6669 ( .A(n5500), .ZN(n5509) );
  OR2_X1 U6670 ( .A1(n5517), .A2(n5501), .ZN(n5502) );
  NAND2_X1 U6671 ( .A1(n5486), .A2(n5502), .ZN(n5780) );
  INV_X1 U6672 ( .A(n5503), .ZN(n5693) );
  OAI22_X1 U6673 ( .A1(n5504), .A2(n6138), .B1(n6187), .B2(n5693), .ZN(n5505)
         );
  AOI21_X1 U6674 ( .B1(n6182), .B2(EBX_REG_27__SCAN_IN), .A(n5505), .ZN(n5507)
         );
  NAND2_X1 U6675 ( .A1(n5511), .A2(REIP_REG_27__SCAN_IN), .ZN(n5506) );
  OAI211_X1 U6676 ( .C1(n5780), .C2(n6197), .A(n5507), .B(n5506), .ZN(n5508)
         );
  AOI21_X1 U6677 ( .B1(n5509), .B2(n6692), .A(n5508), .ZN(n5510) );
  OAI21_X1 U6678 ( .B1(n5587), .B2(n6129), .A(n5510), .ZN(U2800) );
  INV_X1 U6679 ( .A(n5511), .ZN(n5523) );
  NOR2_X1 U6680 ( .A1(n6715), .A2(n6573), .ZN(n5512) );
  AOI21_X1 U6681 ( .B1(n5944), .B2(n5512), .A(REIP_REG_26__SCAN_IN), .ZN(n5522) );
  NAND2_X1 U6682 ( .A1(n5593), .A2(n5592), .ZN(n5595) );
  NAND2_X1 U6683 ( .A1(n5704), .A2(n6146), .ZN(n5521) );
  OAI22_X1 U6684 ( .A1(n5298), .A2(n6138), .B1(n5702), .B2(n6187), .ZN(n5519)
         );
  NOR2_X1 U6685 ( .A1(n5596), .A2(n5515), .ZN(n5516) );
  OR2_X1 U6686 ( .A1(n5517), .A2(n5516), .ZN(n5793) );
  NOR2_X1 U6687 ( .A1(n5793), .A2(n6197), .ZN(n5518) );
  AOI211_X1 U6688 ( .C1(n6182), .C2(EBX_REG_26__SCAN_IN), .A(n5519), .B(n5518), 
        .ZN(n5520) );
  OAI211_X1 U6689 ( .C1(n5523), .C2(n5522), .A(n5521), .B(n5520), .ZN(U2801)
         );
  AOI21_X1 U6690 ( .B1(n6660), .B2(n5524), .A(n5963), .ZN(n5529) );
  AOI22_X1 U6691 ( .A1(EBX_REG_23__SCAN_IN), .A2(n6182), .B1(n5525), .B2(n6160), .ZN(n5526) );
  OAI21_X1 U6692 ( .B1(n5527), .B2(n6138), .A(n5526), .ZN(n5528) );
  AOI211_X1 U6693 ( .C1(n5604), .C2(n6122), .A(n5529), .B(n5528), .ZN(n5530)
         );
  OAI21_X1 U6694 ( .B1(n5658), .B2(n6129), .A(n5530), .ZN(U2804) );
  OAI21_X1 U6695 ( .B1(n5531), .B2(n5533), .A(n5607), .ZN(n5730) );
  NAND2_X1 U6696 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5552) );
  OAI21_X1 U6697 ( .B1(n5552), .B2(n6065), .A(n6713), .ZN(n5540) );
  INV_X1 U6698 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5534) );
  OAI22_X1 U6699 ( .A1(n5534), .A2(n6138), .B1(n5732), .B2(n6187), .ZN(n5539)
         );
  MUX2_X1 U6700 ( .A(n5548), .B(n5546), .S(n5535), .Z(n5537) );
  XNOR2_X1 U6701 ( .A(n5537), .B(n5536), .ZN(n5836) );
  INV_X1 U6702 ( .A(n5836), .ZN(n5615) );
  INV_X1 U6703 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5616) );
  OAI22_X1 U6704 ( .A1(n5615), .A2(n6197), .B1(n5616), .B2(n6140), .ZN(n5538)
         );
  AOI211_X1 U6705 ( .C1(n5540), .C2(n5972), .A(n5539), .B(n5538), .ZN(n5541)
         );
  OAI21_X1 U6706 ( .B1(n5730), .B2(n6129), .A(n5541), .ZN(U2807) );
  AND2_X1 U6707 ( .A1(n5542), .A2(n5543), .ZN(n5544) );
  OR2_X1 U6708 ( .A1(n5531), .A2(n5544), .ZN(n5743) );
  INV_X1 U6709 ( .A(n5545), .ZN(n5547) );
  MUX2_X1 U6710 ( .A(n5548), .B(n5547), .S(n5546), .Z(n5619) );
  NAND2_X1 U6711 ( .A1(n5620), .A2(n5619), .ZN(n5622) );
  XNOR2_X1 U6712 ( .A(n5622), .B(n5549), .ZN(n5844) );
  OAI21_X1 U6713 ( .B1(n6138), .B2(n5738), .A(n6341), .ZN(n5550) );
  AOI21_X1 U6714 ( .B1(n6160), .B2(n5740), .A(n5550), .ZN(n5551) );
  OAI21_X1 U6715 ( .B1(n6140), .B2(n3678), .A(n5551), .ZN(n5555) );
  OAI21_X1 U6716 ( .B1(REIP_REG_19__SCAN_IN), .B2(REIP_REG_18__SCAN_IN), .A(
        n5552), .ZN(n5553) );
  OAI22_X1 U6717 ( .A1(n6064), .A2(n6682), .B1(n5553), .B2(n6065), .ZN(n5554)
         );
  AOI211_X1 U6718 ( .C1(n6122), .C2(n5844), .A(n5555), .B(n5554), .ZN(n5556)
         );
  OAI21_X1 U6719 ( .B1(n5743), .B2(n6129), .A(n5556), .ZN(U2808) );
  OAI21_X1 U6720 ( .B1(n5395), .B2(n5558), .A(n5557), .ZN(n6002) );
  NOR2_X1 U6721 ( .A1(n5626), .A2(n5559), .ZN(n5560) );
  OR2_X1 U6722 ( .A1(n5620), .A2(n5560), .ZN(n5866) );
  INV_X1 U6723 ( .A(n5866), .ZN(n5567) );
  INV_X1 U6724 ( .A(n6003), .ZN(n5562) );
  AOI21_X1 U6725 ( .B1(n6182), .B2(EBX_REG_17__SCAN_IN), .A(n6351), .ZN(n5561)
         );
  OAI21_X1 U6726 ( .B1(n5562), .B2(n6187), .A(n5561), .ZN(n5566) );
  INV_X1 U6727 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6562) );
  INV_X1 U6728 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6560) );
  NOR2_X1 U6729 ( .A1(n6562), .A2(n6560), .ZN(n6075) );
  AOI21_X1 U6730 ( .B1(n6075), .B2(n6072), .A(REIP_REG_17__SCAN_IN), .ZN(n5564) );
  OAI22_X1 U6731 ( .A1(n6064), .A2(n5564), .B1(n5563), .B2(n6138), .ZN(n5565)
         );
  AOI211_X1 U6732 ( .C1(n5567), .C2(n6122), .A(n5566), .B(n5565), .ZN(n5568)
         );
  OAI21_X1 U6733 ( .B1(n6002), .B2(n6129), .A(n5568), .ZN(U2810) );
  INV_X1 U6734 ( .A(n5569), .ZN(n5570) );
  AOI21_X1 U6735 ( .B1(n5571), .B2(n5393), .A(n5570), .ZN(n5750) );
  INV_X1 U6736 ( .A(n5750), .ZN(n5662) );
  AOI22_X1 U6737 ( .A1(EBX_REG_15__SCAN_IN), .A2(n6182), .B1(n6072), .B2(n6560), .ZN(n5572) );
  OAI211_X1 U6738 ( .C1(n6138), .C2(n5573), .A(n5572), .B(n6341), .ZN(n5574)
         );
  AOI21_X1 U6739 ( .B1(REIP_REG_15__SCAN_IN), .B2(n6082), .A(n5574), .ZN(n5582) );
  INV_X1 U6740 ( .A(n5575), .ZN(n5578) );
  INV_X1 U6741 ( .A(n5576), .ZN(n5577) );
  OAI21_X1 U6742 ( .B1(n5225), .B2(n5578), .A(n5577), .ZN(n5579) );
  AND2_X1 U6743 ( .A1(n5579), .A2(n5627), .ZN(n6018) );
  NOR2_X1 U6744 ( .A1(n6187), .A2(n5747), .ZN(n5580) );
  AOI21_X1 U6745 ( .B1(n6018), .B2(n6122), .A(n5580), .ZN(n5581) );
  OAI211_X1 U6746 ( .C1(n5662), .C2(n6129), .A(n5582), .B(n5581), .ZN(U2812)
         );
  INV_X1 U6747 ( .A(n5583), .ZN(n5585) );
  OAI22_X1 U6748 ( .A1(n5585), .A2(n5637), .B1(n6207), .B2(n5584), .ZN(U2828)
         );
  AOI22_X1 U6749 ( .A1(n5773), .A2(n6203), .B1(EBX_REG_28__SCAN_IN), .B2(n5617), .ZN(n5586) );
  OAI21_X1 U6750 ( .B1(n5650), .B2(n5639), .A(n5586), .ZN(U2831) );
  INV_X1 U6751 ( .A(n5587), .ZN(n5695) );
  OAI22_X1 U6752 ( .A1(n5780), .A2(n5637), .B1(n5588), .B2(n6207), .ZN(n5589)
         );
  AOI21_X1 U6753 ( .B1(n5695), .B2(n6204), .A(n5589), .ZN(n5590) );
  INV_X1 U6754 ( .A(n5590), .ZN(U2832) );
  INV_X1 U6755 ( .A(n5704), .ZN(n5655) );
  INV_X1 U6756 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5591) );
  OAI222_X1 U6757 ( .A1(n5639), .A2(n5655), .B1(n5591), .B2(n6207), .C1(n5793), 
        .C2(n5637), .ZN(U2833) );
  OR2_X1 U6758 ( .A1(n5593), .A2(n5592), .ZN(n5594) );
  INV_X1 U6759 ( .A(n5984), .ZN(n5601) );
  INV_X1 U6760 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5600) );
  AOI21_X1 U6761 ( .B1(n5598), .B2(n5597), .A(n5596), .ZN(n5599) );
  INV_X1 U6762 ( .A(n5599), .ZN(n5953) );
  OAI222_X1 U6763 ( .A1(n5601), .A2(n5639), .B1(n6207), .B2(n5600), .C1(n5953), 
        .C2(n5637), .ZN(U2834) );
  INV_X1 U6764 ( .A(n5987), .ZN(n5603) );
  AOI22_X1 U6765 ( .A1(n5960), .A2(n6203), .B1(EBX_REG_24__SCAN_IN), .B2(n5617), .ZN(n5602) );
  OAI21_X1 U6766 ( .B1(n5603), .B2(n5639), .A(n5602), .ZN(U2835) );
  AOI22_X1 U6767 ( .A1(n5604), .A2(n6203), .B1(EBX_REG_23__SCAN_IN), .B2(n5617), .ZN(n5605) );
  OAI21_X1 U6768 ( .B1(n5658), .B2(n5639), .A(n5605), .ZN(U2836) );
  AOI21_X1 U6769 ( .B1(n5608), .B2(n5607), .A(n5606), .ZN(n5993) );
  OR2_X1 U6770 ( .A1(n5611), .A2(n5610), .ZN(n5612) );
  NAND2_X1 U6771 ( .A1(n5609), .A2(n5612), .ZN(n5979) );
  OAI22_X1 U6772 ( .A1(n5979), .A2(n5637), .B1(n5976), .B2(n6207), .ZN(n5613)
         );
  AOI21_X1 U6773 ( .B1(n5993), .B2(n6204), .A(n5613), .ZN(n5614) );
  INV_X1 U6774 ( .A(n5614), .ZN(U2838) );
  OAI222_X1 U6775 ( .A1(n5639), .A2(n5730), .B1(n5616), .B2(n6207), .C1(n5615), 
        .C2(n5637), .ZN(U2839) );
  AOI22_X1 U6776 ( .A1(n5844), .A2(n6203), .B1(EBX_REG_19__SCAN_IN), .B2(n5617), .ZN(n5618) );
  OAI21_X1 U6777 ( .B1(n5743), .B2(n5639), .A(n5618), .ZN(U2840) );
  OR2_X1 U6778 ( .A1(n5620), .A2(n5619), .ZN(n5621) );
  AND2_X1 U6779 ( .A1(n5622), .A2(n5621), .ZN(n5853) );
  INV_X1 U6780 ( .A(n5853), .ZN(n6066) );
  NAND2_X1 U6781 ( .A1(n5557), .A2(n5623), .ZN(n5624) );
  AND2_X1 U6782 ( .A1(n5542), .A2(n5624), .ZN(n6208) );
  INV_X1 U6783 ( .A(n6208), .ZN(n6067) );
  OAI222_X1 U6784 ( .A1(n6066), .A2(n5637), .B1(n6207), .B2(n3682), .C1(n6067), 
        .C2(n5639), .ZN(U2841) );
  OAI222_X1 U6785 ( .A1(n6002), .A2(n5639), .B1(n5625), .B2(n6207), .C1(n5866), 
        .C2(n5637), .ZN(U2842) );
  INV_X1 U6786 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5630) );
  AOI21_X1 U6787 ( .B1(n5628), .B2(n5627), .A(n5626), .ZN(n5629) );
  INV_X1 U6788 ( .A(n5629), .ZN(n6081) );
  OAI222_X1 U6789 ( .A1(n6077), .A2(n5639), .B1(n5630), .B2(n6207), .C1(n5637), 
        .C2(n6081), .ZN(U2843) );
  NOR2_X1 U6790 ( .A1(n6207), .A2(n5631), .ZN(n5632) );
  AOI21_X1 U6791 ( .B1(n6018), .B2(n6203), .A(n5632), .ZN(n5633) );
  OAI21_X1 U6792 ( .B1(n5662), .B2(n5639), .A(n5633), .ZN(U2844) );
  OAI21_X1 U6793 ( .B1(n5635), .B2(n5634), .A(n5393), .ZN(n6086) );
  INV_X1 U6794 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5638) );
  OAI222_X1 U6795 ( .A1(n6086), .A2(n5639), .B1(n5638), .B2(n6207), .C1(n5637), 
        .C2(n5636), .ZN(U2845) );
  NAND3_X1 U6796 ( .A1(n5642), .A2(n5641), .A3(n5640), .ZN(n5644) );
  AOI22_X1 U6797 ( .A1(n6214), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6217), .ZN(n5643) );
  NAND2_X1 U6798 ( .A1(n5644), .A2(n5643), .ZN(U2860) );
  AOI22_X1 U6799 ( .A1(n6214), .A2(DATAI_30_), .B1(n6217), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5646) );
  NAND2_X1 U6800 ( .A1(n6218), .A2(DATAI_14_), .ZN(n5645) );
  OAI211_X1 U6801 ( .C1(n5647), .C2(n5983), .A(n5646), .B(n5645), .ZN(U2861)
         );
  AOI22_X1 U6802 ( .A1(n6214), .A2(DATAI_28_), .B1(n6217), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5649) );
  NAND2_X1 U6803 ( .A1(n6218), .A2(DATAI_12_), .ZN(n5648) );
  OAI211_X1 U6804 ( .C1(n5650), .C2(n5983), .A(n5649), .B(n5648), .ZN(U2863)
         );
  AOI22_X1 U6805 ( .A1(n6214), .A2(DATAI_27_), .B1(n6217), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5652) );
  NAND2_X1 U6806 ( .A1(n6218), .A2(DATAI_11_), .ZN(n5651) );
  OAI211_X1 U6807 ( .C1(n5587), .C2(n5983), .A(n5652), .B(n5651), .ZN(U2864)
         );
  AOI22_X1 U6808 ( .A1(n6214), .A2(DATAI_26_), .B1(n6217), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5654) );
  NAND2_X1 U6809 ( .A1(n6218), .A2(DATAI_10_), .ZN(n5653) );
  OAI211_X1 U6810 ( .C1(n5655), .C2(n5983), .A(n5654), .B(n5653), .ZN(U2865)
         );
  AOI22_X1 U6811 ( .A1(n6214), .A2(DATAI_23_), .B1(n6217), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5657) );
  NAND2_X1 U6812 ( .A1(n6218), .A2(DATAI_7_), .ZN(n5656) );
  OAI211_X1 U6813 ( .C1(n5658), .C2(n5983), .A(n5657), .B(n5656), .ZN(U2868)
         );
  AOI22_X1 U6814 ( .A1(n6214), .A2(DATAI_19_), .B1(n6217), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5660) );
  NAND2_X1 U6815 ( .A1(n6218), .A2(DATAI_3_), .ZN(n5659) );
  OAI211_X1 U6816 ( .C1(n5743), .C2(n5983), .A(n5660), .B(n5659), .ZN(U2872)
         );
  AOI22_X1 U6817 ( .A1(n5663), .A2(DATAI_15_), .B1(n6217), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5661) );
  OAI21_X1 U6818 ( .B1(n5662), .B2(n5983), .A(n5661), .ZN(U2876) );
  AOI22_X1 U6819 ( .A1(n5663), .A2(DATAI_14_), .B1(n6217), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5664) );
  OAI21_X1 U6820 ( .B1(n6086), .B2(n5983), .A(n5664), .ZN(U2877) );
  NAND2_X1 U6821 ( .A1(n5676), .A2(n5665), .ZN(n5666) );
  NAND2_X1 U6822 ( .A1(n5667), .A2(n5666), .ZN(n5668) );
  XNOR2_X1 U6823 ( .A(n5668), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5767)
         );
  INV_X1 U6824 ( .A(n5669), .ZN(n5674) );
  INV_X1 U6825 ( .A(n5670), .ZN(n5672) );
  NOR2_X1 U6826 ( .A1(n6341), .A2(n6767), .ZN(n5762) );
  AOI21_X1 U6827 ( .B1(n6263), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5762), 
        .ZN(n5671) );
  OAI21_X1 U6828 ( .B1(n6281), .B2(n5672), .A(n5671), .ZN(n5673) );
  AOI21_X1 U6829 ( .B1(n5674), .B2(n5749), .A(n5673), .ZN(n5675) );
  OAI21_X1 U6830 ( .B1(n5767), .B2(n6269), .A(n5675), .ZN(U2957) );
  INV_X1 U6831 ( .A(n5678), .ZN(n5698) );
  OR3_X1 U6832 ( .A1(n5677), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .A3(n5698), 
        .ZN(n5688) );
  INV_X1 U6833 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5679) );
  AND2_X1 U6834 ( .A1(n5679), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5680)
         );
  XNOR2_X1 U6835 ( .A(n5682), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5779)
         );
  INV_X1 U6836 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6580) );
  NOR2_X1 U6837 ( .A1(n6341), .A2(n6580), .ZN(n5772) );
  AOI21_X1 U6838 ( .B1(n6263), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5772), 
        .ZN(n5683) );
  OAI21_X1 U6839 ( .B1(n6281), .B2(n5684), .A(n5683), .ZN(n5685) );
  AOI21_X1 U6840 ( .B1(n5686), .B2(n5749), .A(n5685), .ZN(n5687) );
  OAI21_X1 U6841 ( .B1(n6269), .B2(n5779), .A(n5687), .ZN(U2958) );
  INV_X1 U6842 ( .A(n5688), .ZN(n5689) );
  OR2_X1 U6843 ( .A1(n5690), .A2(n5689), .ZN(n5691) );
  XNOR2_X1 U6844 ( .A(n5691), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5789)
         );
  NOR2_X1 U6845 ( .A1(n6341), .A2(n6692), .ZN(n5783) );
  AOI21_X1 U6846 ( .B1(n6263), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5783), 
        .ZN(n5692) );
  OAI21_X1 U6847 ( .B1(n6281), .B2(n5693), .A(n5692), .ZN(n5694) );
  AOI21_X1 U6848 ( .B1(n5695), .B2(n5749), .A(n5694), .ZN(n5696) );
  OAI21_X1 U6849 ( .B1(n5789), .B2(n6269), .A(n5696), .ZN(U2959) );
  NAND2_X1 U6850 ( .A1(n5698), .A2(n5697), .ZN(n5699) );
  XNOR2_X1 U6851 ( .A(n5700), .B(n5699), .ZN(n5797) );
  NOR2_X1 U6852 ( .A1(n6341), .A2(n6650), .ZN(n5791) );
  AOI21_X1 U6853 ( .B1(n6263), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5791), 
        .ZN(n5701) );
  OAI21_X1 U6854 ( .B1(n6281), .B2(n5702), .A(n5701), .ZN(n5703) );
  AOI21_X1 U6855 ( .B1(n5704), .B2(n5749), .A(n5703), .ZN(n5705) );
  OAI21_X1 U6856 ( .B1(n5797), .B2(n6269), .A(n5705), .ZN(U2960) );
  AOI21_X1 U6857 ( .B1(n5707), .B2(n5677), .A(n5706), .ZN(n5805) );
  INV_X1 U6858 ( .A(n5945), .ZN(n5709) );
  NOR2_X1 U6859 ( .A1(n6341), .A2(n6573), .ZN(n5798) );
  AOI21_X1 U6860 ( .B1(n6263), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n5798), 
        .ZN(n5708) );
  OAI21_X1 U6861 ( .B1(n6281), .B2(n5709), .A(n5708), .ZN(n5710) );
  AOI21_X1 U6862 ( .B1(n5984), .B2(n5749), .A(n5710), .ZN(n5711) );
  OAI21_X1 U6863 ( .B1(n5805), .B2(n6269), .A(n5711), .ZN(U2961) );
  AOI21_X1 U6864 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n6249), .A(n5712), 
        .ZN(n5713) );
  XNOR2_X1 U6865 ( .A(n5714), .B(n5713), .ZN(n5818) );
  INV_X1 U6866 ( .A(n5239), .ZN(n5715) );
  NAND2_X1 U6867 ( .A1(n6351), .A2(REIP_REG_22__SCAN_IN), .ZN(n5809) );
  NAND2_X1 U6868 ( .A1(n6263), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5718)
         );
  OAI211_X1 U6869 ( .C1(n6281), .C2(n5964), .A(n5809), .B(n5718), .ZN(n5719)
         );
  AOI21_X1 U6870 ( .B1(n5990), .B2(n5749), .A(n5719), .ZN(n5720) );
  OAI21_X1 U6871 ( .B1(n5818), .B2(n6269), .A(n5720), .ZN(U2964) );
  AOI21_X1 U6872 ( .B1(n5723), .B2(n5721), .A(n5722), .ZN(n5826) );
  INV_X1 U6873 ( .A(n5973), .ZN(n5725) );
  NAND2_X1 U6874 ( .A1(n6263), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5724)
         );
  NAND2_X1 U6875 ( .A1(n6351), .A2(REIP_REG_21__SCAN_IN), .ZN(n5821) );
  OAI211_X1 U6876 ( .C1(n6281), .C2(n5725), .A(n5724), .B(n5821), .ZN(n5726)
         );
  AOI21_X1 U6877 ( .B1(n5993), .B2(n5749), .A(n5726), .ZN(n5727) );
  OAI21_X1 U6878 ( .B1(n5826), .B2(n6269), .A(n5727), .ZN(U2965) );
  XNOR2_X1 U6879 ( .A(n5728), .B(n5729), .ZN(n5838) );
  INV_X1 U6880 ( .A(n5730), .ZN(n5996) );
  OR2_X1 U6881 ( .A1(n6341), .A2(n6713), .ZN(n5830) );
  NAND2_X1 U6882 ( .A1(n6263), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5731)
         );
  OAI211_X1 U6883 ( .C1(n6281), .C2(n5732), .A(n5830), .B(n5731), .ZN(n5733)
         );
  AOI21_X1 U6884 ( .B1(n5996), .B2(n5749), .A(n5733), .ZN(n5734) );
  OAI21_X1 U6885 ( .B1(n5838), .B2(n6269), .A(n5734), .ZN(U2966) );
  MUX2_X1 U6886 ( .A(n5736), .B(n5735), .S(n6249), .Z(n5737) );
  XNOR2_X1 U6887 ( .A(n5737), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5839)
         );
  NAND2_X1 U6888 ( .A1(n5839), .A2(n6276), .ZN(n5742) );
  NOR2_X1 U6889 ( .A1(n6341), .A2(n6682), .ZN(n5843) );
  NOR2_X1 U6890 ( .A1(n5755), .A2(n5738), .ZN(n5739) );
  AOI211_X1 U6891 ( .C1(n6253), .C2(n5740), .A(n5843), .B(n5739), .ZN(n5741)
         );
  OAI211_X1 U6892 ( .C1(n6267), .C2(n5743), .A(n5742), .B(n5741), .ZN(U2967)
         );
  XNOR2_X1 U6893 ( .A(n6249), .B(n6022), .ZN(n5745) );
  XNOR2_X1 U6894 ( .A(n5744), .B(n5745), .ZN(n6019) );
  INV_X1 U6895 ( .A(n6019), .ZN(n5752) );
  AOI22_X1 U6896 ( .A1(n6263), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n6351), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n5746) );
  OAI21_X1 U6897 ( .B1(n6281), .B2(n5747), .A(n5746), .ZN(n5748) );
  AOI21_X1 U6898 ( .B1(n5750), .B2(n5749), .A(n5748), .ZN(n5751) );
  OAI21_X1 U6899 ( .B1(n5752), .B2(n6269), .A(n5751), .ZN(U2971) );
  INV_X1 U6900 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5754) );
  OAI21_X1 U6901 ( .B1(n5755), .B2(n5754), .A(n5753), .ZN(n5757) );
  NOR2_X1 U6902 ( .A1(n6086), .A2(n6267), .ZN(n5756) );
  AOI211_X1 U6903 ( .C1(n6253), .C2(n6087), .A(n5757), .B(n5756), .ZN(n5758)
         );
  OAI21_X1 U6904 ( .B1(n6269), .B2(n5759), .A(n5758), .ZN(U2972) );
  NOR2_X1 U6905 ( .A1(n5760), .A2(n5764), .ZN(n5761) );
  AOI211_X1 U6906 ( .C1(n5763), .C2(n6353), .A(n5762), .B(n5761), .ZN(n5766)
         );
  INV_X1 U6907 ( .A(n5776), .ZN(n5786) );
  NAND3_X1 U6908 ( .A1(n5786), .A2(n5774), .A3(n5764), .ZN(n5765) );
  OAI211_X1 U6909 ( .C1(n5767), .C2(n6283), .A(n5766), .B(n5765), .ZN(U2989)
         );
  OAI21_X1 U6910 ( .B1(n5799), .B2(n5769), .A(n5768), .ZN(n5781) );
  INV_X1 U6911 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5770) );
  NOR2_X1 U6912 ( .A1(n5781), .A2(n5770), .ZN(n5771) );
  AOI211_X1 U6913 ( .C1(n5773), .C2(n6353), .A(n5772), .B(n5771), .ZN(n5778)
         );
  OR3_X1 U6914 ( .A1(n5776), .A2(n5775), .A3(n5774), .ZN(n5777) );
  OAI211_X1 U6915 ( .C1(n5779), .C2(n6283), .A(n5778), .B(n5777), .ZN(U2990)
         );
  INV_X1 U6916 ( .A(n5780), .ZN(n5784) );
  NOR2_X1 U6917 ( .A1(n5781), .A2(n5785), .ZN(n5782) );
  AOI211_X1 U6918 ( .C1(n5784), .C2(n6353), .A(n5783), .B(n5782), .ZN(n5788)
         );
  NAND2_X1 U6919 ( .A1(n5786), .A2(n5785), .ZN(n5787) );
  OAI211_X1 U6920 ( .C1(n5789), .C2(n6283), .A(n5788), .B(n5787), .ZN(U2991)
         );
  INV_X1 U6921 ( .A(n5790), .ZN(n5803) );
  XNOR2_X1 U6922 ( .A(n5802), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5795)
         );
  AOI21_X1 U6923 ( .B1(n5799), .B2(INSTADDRPOINTER_REG_26__SCAN_IN), .A(n5791), 
        .ZN(n5792) );
  OAI21_X1 U6924 ( .B1(n5793), .B2(n6342), .A(n5792), .ZN(n5794) );
  AOI21_X1 U6925 ( .B1(n5803), .B2(n5795), .A(n5794), .ZN(n5796) );
  OAI21_X1 U6926 ( .B1(n5797), .B2(n6283), .A(n5796), .ZN(U2992) );
  AOI21_X1 U6927 ( .B1(n5799), .B2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5798), 
        .ZN(n5800) );
  OAI21_X1 U6928 ( .B1(n5953), .B2(n6342), .A(n5800), .ZN(n5801) );
  AOI21_X1 U6929 ( .B1(n5803), .B2(n5802), .A(n5801), .ZN(n5804) );
  OAI21_X1 U6930 ( .B1(n5805), .B2(n6283), .A(n5804), .ZN(U2993) );
  INV_X1 U6931 ( .A(n5806), .ZN(n5807) );
  AOI21_X1 U6932 ( .B1(n5808), .B2(n5609), .A(n5807), .ZN(n5980) );
  INV_X1 U6933 ( .A(n5819), .ZN(n5811) );
  INV_X1 U6934 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5810) );
  OAI21_X1 U6935 ( .B1(n5811), .B2(n5810), .A(n5809), .ZN(n5816) );
  INV_X1 U6936 ( .A(n5824), .ZN(n5814) );
  NOR3_X1 U6937 ( .A1(n5814), .A2(n5813), .A3(n5812), .ZN(n5815) );
  AOI211_X1 U6938 ( .C1(n6353), .C2(n5980), .A(n5816), .B(n5815), .ZN(n5817)
         );
  OAI21_X1 U6939 ( .B1(n5818), .B2(n6283), .A(n5817), .ZN(U2996) );
  NAND2_X1 U6940 ( .A1(n5819), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5820) );
  OAI211_X1 U6941 ( .C1(n5979), .C2(n6342), .A(n5821), .B(n5820), .ZN(n5822)
         );
  AOI21_X1 U6942 ( .B1(n5824), .B2(n5823), .A(n5822), .ZN(n5825) );
  OAI21_X1 U6943 ( .B1(n5826), .B2(n6283), .A(n5825), .ZN(U2997) );
  INV_X1 U6944 ( .A(n5827), .ZN(n5828) );
  OAI21_X1 U6945 ( .B1(n5828), .B2(INSTADDRPOINTER_REG_17__SCAN_IN), .A(n5863), 
        .ZN(n5850) );
  AOI21_X1 U6946 ( .B1(n5854), .B2(n5829), .A(n5850), .ZN(n5841) );
  OAI21_X1 U6947 ( .B1(n5841), .B2(n5831), .A(n5830), .ZN(n5835) );
  NOR3_X1 U6948 ( .A1(n5847), .A2(n5833), .A3(n5832), .ZN(n5834) );
  AOI211_X1 U6949 ( .C1(n6353), .C2(n5836), .A(n5835), .B(n5834), .ZN(n5837)
         );
  OAI21_X1 U6950 ( .B1(n5838), .B2(n6283), .A(n5837), .ZN(U2998) );
  NAND2_X1 U6951 ( .A1(n5839), .A2(n6355), .ZN(n5846) );
  NOR2_X1 U6952 ( .A1(n5841), .A2(n5840), .ZN(n5842) );
  AOI211_X1 U6953 ( .C1(n5844), .C2(n6353), .A(n5843), .B(n5842), .ZN(n5845)
         );
  OAI211_X1 U6954 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n5847), .A(n5846), .B(n5845), .ZN(U2999) );
  NOR3_X1 U6955 ( .A1(n5386), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n6249), 
        .ZN(n5859) );
  NOR2_X1 U6956 ( .A1(n3789), .A2(n5861), .ZN(n5848) );
  AOI22_X1 U6957 ( .A1(n5859), .A2(n5861), .B1(n5848), .B2(n5385), .ZN(n5849)
         );
  XNOR2_X1 U6958 ( .A(n5849), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5999)
         );
  INV_X1 U6959 ( .A(n5999), .ZN(n5857) );
  INV_X1 U6960 ( .A(n5850), .ZN(n5851) );
  OAI22_X1 U6961 ( .A1(n5851), .A2(n5854), .B1(n6565), .B2(n6341), .ZN(n5852)
         );
  AOI21_X1 U6962 ( .B1(n5853), .B2(n6353), .A(n5852), .ZN(n5856) );
  NAND3_X1 U6963 ( .A1(n5868), .A2(n5854), .A3(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5855) );
  OAI211_X1 U6964 ( .C1(n5857), .C2(n6283), .A(n5856), .B(n5855), .ZN(U3000)
         );
  NOR2_X1 U6965 ( .A1(n3789), .A2(n5858), .ZN(n5860) );
  AOI21_X1 U6966 ( .B1(n5386), .B2(n5860), .A(n5859), .ZN(n5862) );
  XNOR2_X1 U6967 ( .A(n5862), .B(n5861), .ZN(n6006) );
  INV_X1 U6968 ( .A(n5863), .ZN(n5864) );
  AOI22_X1 U6969 ( .A1(n5864), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .B1(n6351), .B2(REIP_REG_17__SCAN_IN), .ZN(n5865) );
  OAI21_X1 U6970 ( .B1(n5866), .B2(n6342), .A(n5865), .ZN(n5867) );
  AOI21_X1 U6971 ( .B1(n5868), .B2(n5861), .A(n5867), .ZN(n5869) );
  OAI21_X1 U6972 ( .B1(n6006), .B2(n6283), .A(n5869), .ZN(U3001) );
  NOR2_X1 U6973 ( .A1(n5871), .A2(n5870), .ZN(n5874) );
  INV_X1 U6974 ( .A(n5872), .ZN(n5873) );
  OAI222_X1 U6975 ( .A1(n5879), .A2(n5876), .B1(n5875), .B2(n5874), .C1(n5873), 
        .C2(n6368), .ZN(n5877) );
  MUX2_X1 U6976 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n5877), .S(n6362), 
        .Z(U3462) );
  NOR2_X1 U6977 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5878), .ZN(n5885)
         );
  INV_X1 U6978 ( .A(n5943), .ZN(n5880) );
  OAI21_X1 U6979 ( .B1(n5880), .B2(n2986), .A(n5879), .ZN(n5882) );
  INV_X1 U6980 ( .A(n5888), .ZN(n5881) );
  NAND2_X1 U6981 ( .A1(n5882), .A2(n5881), .ZN(n5884) );
  NAND2_X1 U6982 ( .A1(n5932), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5893) );
  INV_X1 U6983 ( .A(n5885), .ZN(n5935) );
  NOR2_X1 U6984 ( .A1(n5886), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6365)
         );
  AOI22_X1 U6985 ( .A1(n5888), .A2(n6367), .B1(n5887), .B2(n6365), .ZN(n5934)
         );
  OAI22_X1 U6986 ( .A1(n6451), .A2(n5935), .B1(n5934), .B2(n5889), .ZN(n5890)
         );
  AOI21_X1 U6987 ( .B1(n5891), .B2(n2986), .A(n5890), .ZN(n5892) );
  OAI211_X1 U6988 ( .C1(n6461), .C2(n5943), .A(n5893), .B(n5892), .ZN(U3036)
         );
  NAND2_X1 U6989 ( .A1(n5932), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5899) );
  OAI22_X1 U6990 ( .A1(n5895), .A2(n5935), .B1(n5934), .B2(n5894), .ZN(n5896)
         );
  AOI21_X1 U6991 ( .B1(n5897), .B2(n2986), .A(n5896), .ZN(n5898) );
  OAI211_X1 U6992 ( .C1(n5943), .C2(n5900), .A(n5899), .B(n5898), .ZN(U3037)
         );
  NAND2_X1 U6993 ( .A1(n5932), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5906) );
  OAI22_X1 U6994 ( .A1(n5902), .A2(n5935), .B1(n5934), .B2(n5901), .ZN(n5903)
         );
  AOI21_X1 U6995 ( .B1(n5904), .B2(n2986), .A(n5903), .ZN(n5905) );
  OAI211_X1 U6996 ( .C1(n5943), .C2(n5907), .A(n5906), .B(n5905), .ZN(U3038)
         );
  NAND2_X1 U6997 ( .A1(n5932), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5912) );
  OAI22_X1 U6998 ( .A1(n6431), .A2(n5935), .B1(n5934), .B2(n5908), .ZN(n5909)
         );
  AOI21_X1 U6999 ( .B1(n5910), .B2(n2986), .A(n5909), .ZN(n5911) );
  OAI211_X1 U7000 ( .C1(n5943), .C2(n6436), .A(n5912), .B(n5911), .ZN(U3039)
         );
  NAND2_X1 U7001 ( .A1(n5932), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5917) );
  OAI22_X1 U7002 ( .A1(n6440), .A2(n5935), .B1(n5934), .B2(n5913), .ZN(n5914)
         );
  AOI21_X1 U7003 ( .B1(n5915), .B2(n2986), .A(n5914), .ZN(n5916) );
  OAI211_X1 U7004 ( .C1(n5943), .C2(n6448), .A(n5917), .B(n5916), .ZN(U3040)
         );
  NAND2_X1 U7005 ( .A1(n5932), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5923) );
  OAI22_X1 U7006 ( .A1(n5919), .A2(n5935), .B1(n5934), .B2(n5918), .ZN(n5920)
         );
  AOI21_X1 U7007 ( .B1(n5921), .B2(n2986), .A(n5920), .ZN(n5922) );
  OAI211_X1 U7008 ( .C1(n5943), .C2(n5924), .A(n5923), .B(n5922), .ZN(U3041)
         );
  NAND2_X1 U7009 ( .A1(n5932), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5930) );
  OAI22_X1 U7010 ( .A1(n5926), .A2(n5935), .B1(n5934), .B2(n5925), .ZN(n5927)
         );
  AOI21_X1 U7011 ( .B1(n5928), .B2(n2986), .A(n5927), .ZN(n5929) );
  OAI211_X1 U7012 ( .C1(n5943), .C2(n5931), .A(n5930), .B(n5929), .ZN(U3042)
         );
  NAND2_X1 U7013 ( .A1(n5932), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5941) );
  OAI22_X1 U7014 ( .A1(n5936), .A2(n5935), .B1(n5934), .B2(n5933), .ZN(n5937)
         );
  AOI21_X1 U7015 ( .B1(n5939), .B2(n2986), .A(n5937), .ZN(n5940) );
  OAI211_X1 U7016 ( .C1(n5943), .C2(n5942), .A(n5941), .B(n5940), .ZN(U3043)
         );
  AND2_X1 U7017 ( .A1(n6235), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  NAND2_X1 U7018 ( .A1(n5944), .A2(n6715), .ZN(n5954) );
  AOI21_X1 U7019 ( .B1(n5963), .B2(n5954), .A(n6573), .ZN(n5950) );
  NAND3_X1 U7020 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5944), .A3(n6573), .ZN(
        n5948) );
  AOI22_X1 U7021 ( .A1(EBX_REG_25__SCAN_IN), .A2(n6182), .B1(n5945), .B2(n6160), .ZN(n5947) );
  NAND2_X1 U7022 ( .A1(n6184), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5946)
         );
  NAND3_X1 U7023 ( .A1(n5948), .A2(n5947), .A3(n5946), .ZN(n5949) );
  OR2_X1 U7024 ( .A1(n5950), .A2(n5949), .ZN(n5951) );
  AOI21_X1 U7025 ( .B1(n5984), .B2(n6146), .A(n5951), .ZN(n5952) );
  OAI21_X1 U7026 ( .B1(n6197), .B2(n5953), .A(n5952), .ZN(U2802) );
  INV_X1 U7027 ( .A(n5954), .ZN(n5958) );
  OAI22_X1 U7028 ( .A1(n5956), .A2(n6140), .B1(n5955), .B2(n6138), .ZN(n5957)
         );
  AOI211_X1 U7029 ( .C1(n6160), .C2(n5959), .A(n5958), .B(n5957), .ZN(n5962)
         );
  AOI22_X1 U7030 ( .A1(n5987), .A2(n6146), .B1(n5960), .B2(n6122), .ZN(n5961)
         );
  OAI211_X1 U7031 ( .C1(n5963), .C2(n6715), .A(n5962), .B(n5961), .ZN(U2803)
         );
  INV_X1 U7032 ( .A(n5964), .ZN(n5965) );
  AOI22_X1 U7033 ( .A1(n5965), .A2(n6160), .B1(REIP_REG_22__SCAN_IN), .B2(
        n5972), .ZN(n5970) );
  AOI22_X1 U7034 ( .A1(EBX_REG_22__SCAN_IN), .A2(n6182), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6184), .ZN(n5969) );
  AOI22_X1 U7035 ( .A1(n5990), .A2(n6146), .B1(n5980), .B2(n6122), .ZN(n5968)
         );
  OAI211_X1 U7036 ( .C1(REIP_REG_22__SCAN_IN), .C2(REIP_REG_21__SCAN_IN), .A(
        n5971), .B(n5966), .ZN(n5967) );
  NAND4_X1 U7037 ( .A1(n5970), .A2(n5969), .A3(n5968), .A4(n5967), .ZN(U2805)
         );
  INV_X1 U7038 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6569) );
  AOI22_X1 U7039 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n6184), .B1(n5971), 
        .B2(n6569), .ZN(n5975) );
  AOI22_X1 U7040 ( .A1(n5973), .A2(n6160), .B1(REIP_REG_21__SCAN_IN), .B2(
        n5972), .ZN(n5974) );
  OAI211_X1 U7041 ( .C1(n5976), .C2(n6140), .A(n5975), .B(n5974), .ZN(n5977)
         );
  AOI21_X1 U7042 ( .B1(n5993), .B2(n6146), .A(n5977), .ZN(n5978) );
  OAI21_X1 U7043 ( .B1(n5979), .B2(n6197), .A(n5978), .ZN(U2806) );
  INV_X1 U7044 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5982) );
  AOI22_X1 U7045 ( .A1(n5990), .A2(n6204), .B1(n5980), .B2(n6203), .ZN(n5981)
         );
  OAI21_X1 U7046 ( .B1(n6207), .B2(n5982), .A(n5981), .ZN(U2837) );
  AOI22_X1 U7047 ( .A1(n5984), .A2(n6215), .B1(n6214), .B2(DATAI_25_), .ZN(
        n5986) );
  AOI22_X1 U7048 ( .A1(n6218), .A2(DATAI_9_), .B1(n6217), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5985) );
  NAND2_X1 U7049 ( .A1(n5986), .A2(n5985), .ZN(U2866) );
  AOI22_X1 U7050 ( .A1(n5987), .A2(n6215), .B1(DATAI_24_), .B2(n6214), .ZN(
        n5989) );
  AOI22_X1 U7051 ( .A1(n6218), .A2(DATAI_8_), .B1(n6217), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5988) );
  NAND2_X1 U7052 ( .A1(n5989), .A2(n5988), .ZN(U2867) );
  AOI22_X1 U7053 ( .A1(n5990), .A2(n6215), .B1(n6214), .B2(DATAI_22_), .ZN(
        n5992) );
  AOI22_X1 U7054 ( .A1(n6218), .A2(DATAI_6_), .B1(n6217), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5991) );
  NAND2_X1 U7055 ( .A1(n5992), .A2(n5991), .ZN(U2869) );
  AOI22_X1 U7056 ( .A1(n5993), .A2(n6215), .B1(n6214), .B2(DATAI_21_), .ZN(
        n5995) );
  AOI22_X1 U7057 ( .A1(n6218), .A2(DATAI_5_), .B1(n6217), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5994) );
  NAND2_X1 U7058 ( .A1(n5995), .A2(n5994), .ZN(U2870) );
  AOI22_X1 U7059 ( .A1(n5996), .A2(n6215), .B1(n6214), .B2(DATAI_20_), .ZN(
        n5998) );
  AOI22_X1 U7060 ( .A1(n6218), .A2(DATAI_4_), .B1(n6217), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5997) );
  NAND2_X1 U7061 ( .A1(n5998), .A2(n5997), .ZN(U2871) );
  AOI22_X1 U7062 ( .A1(n6351), .A2(REIP_REG_18__SCAN_IN), .B1(n6263), .B2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n6001) );
  AOI22_X1 U7063 ( .A1(n5999), .A2(n6276), .B1(n5749), .B2(n6208), .ZN(n6000)
         );
  OAI211_X1 U7064 ( .C1(n6281), .C2(n6071), .A(n6001), .B(n6000), .ZN(U2968)
         );
  AOI22_X1 U7065 ( .A1(n6351), .A2(REIP_REG_17__SCAN_IN), .B1(n6263), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6005) );
  INV_X1 U7066 ( .A(n6002), .ZN(n6211) );
  AOI22_X1 U7067 ( .A1(n6211), .A2(n5749), .B1(n6253), .B2(n6003), .ZN(n6004)
         );
  OAI211_X1 U7068 ( .C1(n6006), .C2(n6269), .A(n6005), .B(n6004), .ZN(U2969)
         );
  AOI22_X1 U7069 ( .A1(n6351), .A2(REIP_REG_13__SCAN_IN), .B1(n6263), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6010) );
  XNOR2_X1 U7070 ( .A(n6007), .B(n6008), .ZN(n6032) );
  AOI22_X1 U7071 ( .A1(n6032), .A2(n6276), .B1(n5749), .B2(n6199), .ZN(n6009)
         );
  OAI211_X1 U7072 ( .C1(n6281), .C2(n6101), .A(n6010), .B(n6009), .ZN(U2973)
         );
  INV_X1 U7073 ( .A(n6011), .ZN(n6012) );
  OAI21_X1 U7074 ( .B1(n6296), .B2(n6012), .A(n6287), .ZN(n6021) );
  OAI22_X1 U7075 ( .A1(n6013), .A2(n6283), .B1(n6342), .B2(n6081), .ZN(n6014)
         );
  AOI21_X1 U7076 ( .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n6021), .A(n6014), 
        .ZN(n6017) );
  OAI211_X1 U7077 ( .C1(INSTADDRPOINTER_REG_15__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A(n6023), .B(n6015), .ZN(n6016) );
  OAI211_X1 U7078 ( .C1(n6562), .C2(n6341), .A(n6017), .B(n6016), .ZN(U3002)
         );
  AOI22_X1 U7079 ( .A1(n6019), .A2(n6355), .B1(n6353), .B2(n6018), .ZN(n6025)
         );
  NOR2_X1 U7080 ( .A1(n6341), .A2(n6560), .ZN(n6020) );
  AOI221_X1 U7081 ( .B1(n6023), .B2(n6022), .C1(n6021), .C2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .A(n6020), .ZN(n6024) );
  NAND2_X1 U7082 ( .A1(n6025), .A2(n6024), .ZN(U3003) );
  NOR2_X1 U7083 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n6026), .ZN(n6027)
         );
  AOI22_X1 U7084 ( .A1(n6351), .A2(REIP_REG_13__SCAN_IN), .B1(n6028), .B2(
        n6027), .ZN(n6037) );
  OR2_X1 U7085 ( .A1(n6030), .A2(n6029), .ZN(n6031) );
  AND2_X1 U7086 ( .A1(n5225), .A2(n6031), .ZN(n6198) );
  AOI22_X1 U7087 ( .A1(n6032), .A2(n6355), .B1(n6353), .B2(n6198), .ZN(n6036)
         );
  OAI21_X1 U7088 ( .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n6034), .A(n6033), 
        .ZN(n6035) );
  NAND3_X1 U7089 ( .A1(n6037), .A2(n6036), .A3(n6035), .ZN(U3005) );
  INV_X1 U7090 ( .A(n6152), .ZN(n6039) );
  NAND3_X1 U7091 ( .A1(n6039), .A2(n6038), .A3(n6593), .ZN(n6041) );
  OAI22_X1 U7092 ( .A1(n6042), .A2(n6041), .B1(n6040), .B2(n6598), .ZN(U3455)
         );
  INV_X1 U7093 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6536) );
  INV_X1 U7094 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6530) );
  AOI21_X1 U7095 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6536), .A(n6530), .ZN(n6047) );
  INV_X1 U7096 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6752) );
  AND2_X1 U7097 ( .A1(n6530), .A2(STATE_REG_1__SCAN_IN), .ZN(n6820) );
  AOI21_X1 U7098 ( .B1(n6047), .B2(n6752), .A(n6820), .ZN(U2789) );
  NAND2_X1 U7099 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6613), .ZN(n6045) );
  OAI21_X1 U7100 ( .B1(n6043), .B2(n6505), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6044) );
  OAI21_X1 U7101 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6045), .A(n6044), .ZN(
        U2790) );
  INV_X2 U7102 ( .A(n6820), .ZN(n6819) );
  NOR2_X1 U7103 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6048) );
  OAI21_X1 U7104 ( .B1(n6048), .B2(D_C_N_REG_SCAN_IN), .A(n6819), .ZN(n6046)
         );
  OAI21_X1 U7105 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6819), .A(n6046), .ZN(
        U2791) );
  NOR2_X1 U7106 ( .A1(n6820), .A2(n6047), .ZN(n6588) );
  OAI21_X1 U7107 ( .B1(BS16_N), .B2(n6048), .A(n6588), .ZN(n6586) );
  OAI21_X1 U7108 ( .B1(n6588), .B2(n6728), .A(n6586), .ZN(U2792) );
  OAI21_X1 U7109 ( .B1(n6049), .B2(n6718), .A(n6269), .ZN(U2793) );
  NOR4_X1 U7110 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(
        DATAWIDTH_REG_21__SCAN_IN), .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n6053) );
  NOR4_X1 U7111 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .A3(DATAWIDTH_REG_18__SCAN_IN), .A4(
        DATAWIDTH_REG_19__SCAN_IN), .ZN(n6052) );
  NOR4_X1 U7112 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6051) );
  NOR4_X1 U7113 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n6050) );
  NAND4_X1 U7114 ( .A1(n6053), .A2(n6052), .A3(n6051), .A4(n6050), .ZN(n6059)
         );
  NOR4_X1 U7115 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), 
        .A3(DATAWIDTH_REG_6__SCAN_IN), .A4(DATAWIDTH_REG_7__SCAN_IN), .ZN(
        n6057) );
  AOI211_X1 U7116 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_2__SCAN_IN), .B(
        DATAWIDTH_REG_3__SCAN_IN), .ZN(n6056) );
  NOR4_X1 U7117 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(
        DATAWIDTH_REG_13__SCAN_IN), .A3(DATAWIDTH_REG_14__SCAN_IN), .A4(
        DATAWIDTH_REG_15__SCAN_IN), .ZN(n6055) );
  NOR4_X1 U7118 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(DATAWIDTH_REG_9__SCAN_IN), 
        .A3(DATAWIDTH_REG_10__SCAN_IN), .A4(DATAWIDTH_REG_11__SCAN_IN), .ZN(
        n6054) );
  NAND4_X1 U7119 ( .A1(n6057), .A2(n6056), .A3(n6055), .A4(n6054), .ZN(n6058)
         );
  NOR2_X1 U7120 ( .A1(n6059), .A2(n6058), .ZN(n6603) );
  INV_X1 U7121 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6729) );
  NOR3_X1 U7122 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6061) );
  OAI21_X1 U7123 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6061), .A(n6603), .ZN(n6060)
         );
  OAI21_X1 U7124 ( .B1(n6603), .B2(n6729), .A(n6060), .ZN(U2794) );
  INV_X1 U7125 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6587) );
  AOI21_X1 U7126 ( .B1(n6600), .B2(n6587), .A(n6061), .ZN(n6062) );
  INV_X1 U7127 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6751) );
  INV_X1 U7128 ( .A(n6603), .ZN(n6606) );
  AOI22_X1 U7129 ( .A1(n6603), .A2(n6062), .B1(n6751), .B2(n6606), .ZN(U2795)
         );
  AOI21_X1 U7130 ( .B1(n6184), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6351), 
        .ZN(n6063) );
  OAI221_X1 U7131 ( .B1(REIP_REG_18__SCAN_IN), .B2(n6065), .C1(n6565), .C2(
        n6064), .A(n6063), .ZN(n6069) );
  OAI22_X1 U7132 ( .A1(n6067), .A2(n6129), .B1(n6197), .B2(n6066), .ZN(n6068)
         );
  AOI211_X1 U7133 ( .C1(EBX_REG_18__SCAN_IN), .C2(n6182), .A(n6069), .B(n6068), 
        .ZN(n6070) );
  OAI21_X1 U7134 ( .B1(n6071), .B2(n6187), .A(n6070), .ZN(U2809) );
  OAI21_X1 U7135 ( .B1(REIP_REG_16__SCAN_IN), .B2(REIP_REG_15__SCAN_IN), .A(
        n6072), .ZN(n6074) );
  AOI22_X1 U7136 ( .A1(EBX_REG_16__SCAN_IN), .A2(n6182), .B1(
        REIP_REG_16__SCAN_IN), .B2(n6082), .ZN(n6073) );
  OAI21_X1 U7137 ( .B1(n6075), .B2(n6074), .A(n6073), .ZN(n6076) );
  AOI211_X1 U7138 ( .C1(n6184), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6351), 
        .B(n6076), .ZN(n6080) );
  INV_X1 U7139 ( .A(n6077), .ZN(n6216) );
  AOI22_X1 U7140 ( .A1(n6216), .A2(n6146), .B1(n6160), .B2(n6078), .ZN(n6079)
         );
  OAI211_X1 U7141 ( .C1(n6197), .C2(n6081), .A(n6080), .B(n6079), .ZN(U2811)
         );
  AOI22_X1 U7142 ( .A1(n6122), .A2(n6083), .B1(REIP_REG_14__SCAN_IN), .B2(
        n6082), .ZN(n6092) );
  AOI22_X1 U7143 ( .A1(PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n6184), .B1(n6085), 
        .B2(n6084), .ZN(n6091) );
  AOI21_X1 U7144 ( .B1(n6182), .B2(EBX_REG_14__SCAN_IN), .A(n6351), .ZN(n6090)
         );
  INV_X1 U7145 ( .A(n6086), .ZN(n6088) );
  AOI22_X1 U7146 ( .A1(n6088), .A2(n6146), .B1(n6160), .B2(n6087), .ZN(n6089)
         );
  NAND4_X1 U7147 ( .A1(n6092), .A2(n6091), .A3(n6090), .A4(n6089), .ZN(U2813)
         );
  INV_X1 U7148 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6555) );
  INV_X1 U7149 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6557) );
  AOI211_X1 U7150 ( .C1(n6555), .C2(n6557), .A(n6095), .B(n6176), .ZN(n6094)
         );
  AOI22_X1 U7151 ( .A1(n6122), .A2(n6198), .B1(n6094), .B2(n6093), .ZN(n6100)
         );
  INV_X1 U7152 ( .A(n6095), .ZN(n6102) );
  OAI21_X1 U7153 ( .B1(n6176), .B2(n6102), .A(n6159), .ZN(n6117) );
  AOI22_X1 U7154 ( .A1(PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n6184), .B1(
        REIP_REG_13__SCAN_IN), .B2(n6117), .ZN(n6097) );
  NAND2_X1 U7155 ( .A1(n6182), .A2(EBX_REG_13__SCAN_IN), .ZN(n6096) );
  NAND3_X1 U7156 ( .A1(n6097), .A2(n6341), .A3(n6096), .ZN(n6098) );
  AOI21_X1 U7157 ( .B1(n6199), .B2(n6146), .A(n6098), .ZN(n6099) );
  OAI211_X1 U7158 ( .C1(n6101), .C2(n6187), .A(n6100), .B(n6099), .ZN(U2814)
         );
  AOI22_X1 U7159 ( .A1(EBX_REG_12__SCAN_IN), .A2(n6182), .B1(
        REIP_REG_12__SCAN_IN), .B2(n6117), .ZN(n6109) );
  AOI21_X1 U7160 ( .B1(PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n6184), .A(n6351), 
        .ZN(n6104) );
  NAND3_X1 U7161 ( .A1(n6193), .A2(n6555), .A3(n6102), .ZN(n6103) );
  OAI211_X1 U7162 ( .C1(n6105), .C2(n6129), .A(n6104), .B(n6103), .ZN(n6106)
         );
  AOI21_X1 U7163 ( .B1(n6107), .B2(n6160), .A(n6106), .ZN(n6108) );
  OAI211_X1 U7164 ( .C1(n6197), .C2(n6110), .A(n6109), .B(n6108), .ZN(U2815)
         );
  NAND2_X1 U7165 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .ZN(
        n6126) );
  NOR3_X1 U7166 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6126), .A3(n6123), .ZN(n6111) );
  AOI211_X1 U7167 ( .C1(n6184), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6351), 
        .B(n6111), .ZN(n6121) );
  AOI21_X1 U7168 ( .B1(n6114), .B2(n6113), .A(n6112), .ZN(n6116) );
  OR2_X1 U7169 ( .A1(n6116), .A2(n6115), .ZN(n6284) );
  INV_X1 U7170 ( .A(n6284), .ZN(n6202) );
  AOI22_X1 U7171 ( .A1(EBX_REG_11__SCAN_IN), .A2(n6182), .B1(n6122), .B2(n6202), .ZN(n6120) );
  AOI22_X1 U7172 ( .A1(n6254), .A2(n6146), .B1(n6160), .B2(n6252), .ZN(n6119)
         );
  NAND2_X1 U7173 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6117), .ZN(n6118) );
  NAND4_X1 U7174 ( .A1(n6121), .A2(n6120), .A3(n6119), .A4(n6118), .ZN(U2816)
         );
  INV_X1 U7175 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6135) );
  AOI22_X1 U7176 ( .A1(EBX_REG_10__SCAN_IN), .A2(n6182), .B1(n6122), .B2(n6293), .ZN(n6134) );
  AOI21_X1 U7177 ( .B1(n6135), .B2(n6550), .A(n6123), .ZN(n6127) );
  OAI21_X1 U7178 ( .B1(n6138), .B2(n6124), .A(n6341), .ZN(n6125) );
  AOI21_X1 U7179 ( .B1(n6127), .B2(n6126), .A(n6125), .ZN(n6128) );
  OAI21_X1 U7180 ( .B1(n6130), .B2(n6129), .A(n6128), .ZN(n6131) );
  AOI21_X1 U7181 ( .B1(n6132), .B2(n6160), .A(n6131), .ZN(n6133) );
  OAI211_X1 U7182 ( .C1(n6136), .C2(n6135), .A(n6134), .B(n6133), .ZN(U2817)
         );
  OAI21_X1 U7183 ( .B1(n6138), .B2(n6137), .A(n6341), .ZN(n6143) );
  OAI22_X1 U7184 ( .A1(n6141), .A2(n6140), .B1(n6197), .B2(n6139), .ZN(n6142)
         );
  NOR3_X1 U7185 ( .A1(n6144), .A2(n6143), .A3(n6142), .ZN(n6148) );
  AOI22_X1 U7186 ( .A1(n6258), .A2(n6146), .B1(REIP_REG_6__SCAN_IN), .B2(n6145), .ZN(n6147) );
  OAI211_X1 U7187 ( .C1(n6262), .C2(n6187), .A(n6148), .B(n6147), .ZN(U2821)
         );
  NOR3_X1 U7188 ( .A1(n6176), .A2(REIP_REG_4__SCAN_IN), .A3(n6150), .ZN(n6149)
         );
  AOI211_X1 U7189 ( .C1(n6184), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6351), 
        .B(n6149), .ZN(n6158) );
  OAI21_X1 U7190 ( .B1(n6183), .B2(n6150), .A(n6178), .ZN(n6169) );
  OAI22_X1 U7191 ( .A1(n6169), .A2(n6542), .B1(n6152), .B2(n6151), .ZN(n6156)
         );
  OAI22_X1 U7192 ( .A1(n6154), .A2(n6188), .B1(n6153), .B2(n6187), .ZN(n6155)
         );
  AOI211_X1 U7193 ( .C1(EBX_REG_4__SCAN_IN), .C2(n6182), .A(n6156), .B(n6155), 
        .ZN(n6157) );
  OAI211_X1 U7194 ( .C1(n6197), .C2(n6343), .A(n6158), .B(n6157), .ZN(U2823)
         );
  INV_X1 U7195 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6539) );
  NAND3_X1 U7196 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6159), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n6177) );
  INV_X1 U7197 ( .A(n6273), .ZN(n6161) );
  AOI22_X1 U7198 ( .A1(n6161), .A2(n6160), .B1(n6184), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6163) );
  NAND2_X1 U7199 ( .A1(n6182), .A2(EBX_REG_3__SCAN_IN), .ZN(n6162) );
  OAI211_X1 U7200 ( .C1(n6197), .C2(n6164), .A(n6163), .B(n6162), .ZN(n6166)
         );
  NOR2_X1 U7201 ( .A1(n6268), .A2(n6188), .ZN(n6165) );
  AOI211_X1 U7202 ( .C1(n6192), .C2(n6167), .A(n6166), .B(n6165), .ZN(n6168)
         );
  OAI221_X1 U7203 ( .B1(n6169), .B2(n6539), .C1(n6169), .C2(n6177), .A(n6168), 
        .ZN(U2824) );
  INV_X1 U7204 ( .A(n6188), .ZN(n6175) );
  AOI22_X1 U7205 ( .A1(n6182), .A2(EBX_REG_2__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n6184), .ZN(n6172) );
  NAND2_X1 U7206 ( .A1(n6192), .A2(n6170), .ZN(n6171) );
  OAI211_X1 U7207 ( .C1(n6197), .C2(n6173), .A(n6172), .B(n6171), .ZN(n6174)
         );
  AOI21_X1 U7208 ( .B1(n6275), .B2(n6175), .A(n6174), .ZN(n6181) );
  NOR2_X1 U7209 ( .A1(n6176), .A2(n6600), .ZN(n6179) );
  OAI211_X1 U7210 ( .C1(n6179), .C2(REIP_REG_2__SCAN_IN), .A(n6178), .B(n6177), 
        .ZN(n6180) );
  OAI211_X1 U7211 ( .C1(n6187), .C2(n6280), .A(n6181), .B(n6180), .ZN(U2825)
         );
  NAND2_X1 U7212 ( .A1(n6182), .A2(EBX_REG_1__SCAN_IN), .ZN(n6186) );
  AOI22_X1 U7213 ( .A1(n6184), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6183), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n6185) );
  OAI211_X1 U7214 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n6187), .A(n6186), 
        .B(n6185), .ZN(n6191) );
  NOR2_X1 U7215 ( .A1(n6189), .A2(n6188), .ZN(n6190) );
  AOI211_X1 U7216 ( .C1(n6192), .C2(n4339), .A(n6191), .B(n6190), .ZN(n6195)
         );
  NAND2_X1 U7217 ( .A1(n6193), .A2(n6600), .ZN(n6194) );
  OAI211_X1 U7218 ( .C1(n6197), .C2(n6196), .A(n6195), .B(n6194), .ZN(U2826)
         );
  AOI22_X1 U7219 ( .A1(n6199), .A2(n6204), .B1(n6203), .B2(n6198), .ZN(n6200)
         );
  OAI21_X1 U7220 ( .B1(n6207), .B2(n6201), .A(n6200), .ZN(U2846) );
  AOI22_X1 U7221 ( .A1(n6254), .A2(n6204), .B1(n6203), .B2(n6202), .ZN(n6205)
         );
  OAI21_X1 U7222 ( .B1(n6207), .B2(n6206), .A(n6205), .ZN(U2848) );
  AOI22_X1 U7223 ( .A1(n6208), .A2(n6215), .B1(n6214), .B2(DATAI_18_), .ZN(
        n6210) );
  AOI22_X1 U7224 ( .A1(n6218), .A2(DATAI_2_), .B1(n6217), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6209) );
  NAND2_X1 U7225 ( .A1(n6210), .A2(n6209), .ZN(U2873) );
  AOI22_X1 U7226 ( .A1(n6211), .A2(n6215), .B1(n6214), .B2(DATAI_17_), .ZN(
        n6213) );
  AOI22_X1 U7227 ( .A1(n6218), .A2(DATAI_1_), .B1(n6217), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6212) );
  NAND2_X1 U7228 ( .A1(n6213), .A2(n6212), .ZN(U2874) );
  AOI22_X1 U7229 ( .A1(n6216), .A2(n6215), .B1(n6214), .B2(DATAI_16_), .ZN(
        n6220) );
  AOI22_X1 U7230 ( .A1(n6218), .A2(DATAI_0_), .B1(n6217), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6219) );
  NAND2_X1 U7231 ( .A1(n6220), .A2(n6219), .ZN(U2875) );
  AOI22_X1 U7232 ( .A1(n6243), .A2(LWORD_REG_15__SCAN_IN), .B1(n6235), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6222) );
  OAI21_X1 U7233 ( .B1(n4292), .B2(n6245), .A(n6222), .ZN(U2908) );
  AOI22_X1 U7234 ( .A1(n6243), .A2(LWORD_REG_14__SCAN_IN), .B1(n6235), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6223) );
  OAI21_X1 U7235 ( .B1(n4360), .B2(n6245), .A(n6223), .ZN(U2909) );
  AOI22_X1 U7236 ( .A1(n6243), .A2(LWORD_REG_13__SCAN_IN), .B1(n6235), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6224) );
  OAI21_X1 U7237 ( .B1(n4375), .B2(n6245), .A(n6224), .ZN(U2910) );
  AOI22_X1 U7238 ( .A1(n6243), .A2(LWORD_REG_12__SCAN_IN), .B1(n6235), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6225) );
  OAI21_X1 U7239 ( .B1(n6226), .B2(n6245), .A(n6225), .ZN(U2911) );
  AOI22_X1 U7240 ( .A1(n6243), .A2(LWORD_REG_11__SCAN_IN), .B1(n6235), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6227) );
  OAI21_X1 U7241 ( .B1(n4379), .B2(n6245), .A(n6227), .ZN(U2912) );
  AOI22_X1 U7242 ( .A1(n6243), .A2(LWORD_REG_10__SCAN_IN), .B1(n6235), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6228) );
  OAI21_X1 U7243 ( .B1(n4358), .B2(n6245), .A(n6228), .ZN(U2913) );
  AOI22_X1 U7244 ( .A1(n6243), .A2(LWORD_REG_9__SCAN_IN), .B1(n6235), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6229) );
  OAI21_X1 U7245 ( .B1(n4383), .B2(n6245), .A(n6229), .ZN(U2914) );
  AOI22_X1 U7246 ( .A1(n6243), .A2(LWORD_REG_8__SCAN_IN), .B1(n6235), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6230) );
  OAI21_X1 U7247 ( .B1(n4371), .B2(n6245), .A(n6230), .ZN(U2915) );
  AOI22_X1 U7248 ( .A1(n6243), .A2(LWORD_REG_7__SCAN_IN), .B1(n6235), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6231) );
  OAI21_X1 U7249 ( .B1(n4388), .B2(n6245), .A(n6231), .ZN(U2916) );
  AOI22_X1 U7250 ( .A1(n6243), .A2(LWORD_REG_6__SCAN_IN), .B1(n6235), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6232) );
  OAI21_X1 U7251 ( .B1(n4364), .B2(n6245), .A(n6232), .ZN(U2917) );
  AOI22_X1 U7252 ( .A1(n6243), .A2(LWORD_REG_5__SCAN_IN), .B1(n6235), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6233) );
  OAI21_X1 U7253 ( .B1(n6234), .B2(n6245), .A(n6233), .ZN(U2918) );
  AOI22_X1 U7254 ( .A1(n6243), .A2(LWORD_REG_4__SCAN_IN), .B1(n6235), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6236) );
  OAI21_X1 U7255 ( .B1(n4368), .B2(n6245), .A(n6236), .ZN(U2919) );
  AOI22_X1 U7256 ( .A1(n6243), .A2(LWORD_REG_3__SCAN_IN), .B1(n6242), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6237) );
  OAI21_X1 U7257 ( .B1(n4417), .B2(n6245), .A(n6237), .ZN(U2920) );
  AOI22_X1 U7258 ( .A1(n6243), .A2(LWORD_REG_2__SCAN_IN), .B1(n6242), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6238) );
  OAI21_X1 U7259 ( .B1(n6239), .B2(n6245), .A(n6238), .ZN(U2921) );
  AOI22_X1 U7260 ( .A1(n6243), .A2(LWORD_REG_1__SCAN_IN), .B1(n6242), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6240) );
  OAI21_X1 U7261 ( .B1(n6241), .B2(n6245), .A(n6240), .ZN(U2922) );
  AOI22_X1 U7262 ( .A1(n6243), .A2(LWORD_REG_0__SCAN_IN), .B1(n6242), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6244) );
  OAI21_X1 U7263 ( .B1(n6246), .B2(n6245), .A(n6244), .ZN(U2923) );
  NAND2_X1 U7264 ( .A1(n6247), .A2(n6248), .ZN(n6251) );
  XNOR2_X1 U7265 ( .A(n6249), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6250)
         );
  XNOR2_X1 U7266 ( .A(n6251), .B(n6250), .ZN(n6282) );
  AOI22_X1 U7267 ( .A1(n6351), .A2(REIP_REG_11__SCAN_IN), .B1(n6263), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6256) );
  AOI22_X1 U7268 ( .A1(n6254), .A2(n5749), .B1(n6253), .B2(n6252), .ZN(n6255)
         );
  OAI211_X1 U7269 ( .C1(n6282), .C2(n6269), .A(n6256), .B(n6255), .ZN(U2975)
         );
  AOI22_X1 U7270 ( .A1(n6351), .A2(REIP_REG_6__SCAN_IN), .B1(n6263), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6261) );
  INV_X1 U7271 ( .A(n6257), .ZN(n6259) );
  AOI22_X1 U7272 ( .A1(n6259), .A2(n6276), .B1(n5749), .B2(n6258), .ZN(n6260)
         );
  OAI211_X1 U7273 ( .C1(n6281), .C2(n6262), .A(n6261), .B(n6260), .ZN(U2980)
         );
  AOI22_X1 U7274 ( .A1(n6351), .A2(REIP_REG_3__SCAN_IN), .B1(n6263), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6272) );
  OAI21_X1 U7275 ( .B1(n6264), .B2(n6266), .A(n6265), .ZN(n6354) );
  OAI22_X1 U7276 ( .A1(n6354), .A2(n6269), .B1(n6268), .B2(n6267), .ZN(n6270)
         );
  INV_X1 U7277 ( .A(n6270), .ZN(n6271) );
  OAI211_X1 U7278 ( .C1(n6281), .C2(n6273), .A(n6272), .B(n6271), .ZN(U2983)
         );
  AOI22_X1 U7279 ( .A1(n6351), .A2(REIP_REG_2__SCAN_IN), .B1(n6263), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6279) );
  INV_X1 U7280 ( .A(n6274), .ZN(n6277) );
  AOI22_X1 U7281 ( .A1(n6277), .A2(n6276), .B1(n6275), .B2(n5749), .ZN(n6278)
         );
  OAI211_X1 U7282 ( .C1(n6281), .C2(n6280), .A(n6279), .B(n6278), .ZN(U2984)
         );
  INV_X1 U7283 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6552) );
  OAI222_X1 U7284 ( .A1(n6284), .A2(n6342), .B1(n6341), .B2(n6552), .C1(n6283), 
        .C2(n6282), .ZN(n6285) );
  INV_X1 U7285 ( .A(n6285), .ZN(n6286) );
  OAI221_X1 U7286 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6288), .C1(
        n3512), .C2(n6287), .A(n6286), .ZN(U3007) );
  INV_X1 U7287 ( .A(n6312), .ZN(n6295) );
  NOR2_X1 U7288 ( .A1(n6289), .A2(n6345), .ZN(n6320) );
  NAND2_X1 U7289 ( .A1(n6295), .A2(n6320), .ZN(n6308) );
  AOI22_X1 U7290 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n6290), .B1(
        INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n5140), .ZN(n6300) );
  INV_X1 U7291 ( .A(n6291), .ZN(n6292) );
  AOI21_X1 U7292 ( .B1(n6293), .B2(n6353), .A(n6292), .ZN(n6299) );
  INV_X1 U7293 ( .A(n6294), .ZN(n6325) );
  OAI21_X1 U7294 ( .B1(n6296), .B2(n6295), .A(n6325), .ZN(n6304) );
  AOI22_X1 U7295 ( .A1(n6297), .A2(n6355), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6304), .ZN(n6298) );
  OAI211_X1 U7296 ( .C1(n6308), .C2(n6300), .A(n6299), .B(n6298), .ZN(U3008)
         );
  INV_X1 U7297 ( .A(n6301), .ZN(n6302) );
  AOI21_X1 U7298 ( .B1(n6303), .B2(n6353), .A(n6302), .ZN(n6307) );
  AOI22_X1 U7299 ( .A1(n6305), .A2(n6355), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n6304), .ZN(n6306) );
  OAI211_X1 U7300 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6308), .A(n6307), 
        .B(n6306), .ZN(U3009) );
  OAI222_X1 U7301 ( .A1(n6310), .A2(n6342), .B1(n6341), .B2(n6548), .C1(n6283), 
        .C2(n6309), .ZN(n6311) );
  INV_X1 U7302 ( .A(n6311), .ZN(n6314) );
  OAI211_X1 U7303 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n6320), .B(n6312), .ZN(n6313) );
  OAI211_X1 U7304 ( .C1(n6325), .C2(n6315), .A(n6314), .B(n6313), .ZN(U3010)
         );
  INV_X1 U7305 ( .A(n6316), .ZN(n6317) );
  AOI21_X1 U7306 ( .B1(n6318), .B2(n6353), .A(n6317), .ZN(n6323) );
  INV_X1 U7307 ( .A(n6319), .ZN(n6321) );
  AOI22_X1 U7308 ( .A1(n6321), .A2(n6355), .B1(n6320), .B2(n6324), .ZN(n6322)
         );
  OAI211_X1 U7309 ( .C1(n6325), .C2(n6324), .A(n6323), .B(n6322), .ZN(U3011)
         );
  OAI21_X1 U7310 ( .B1(n6328), .B2(n6327), .A(n6326), .ZN(n6329) );
  AOI21_X1 U7311 ( .B1(n6339), .B2(n6330), .A(n6329), .ZN(n6336) );
  INV_X1 U7312 ( .A(n6331), .ZN(n6333) );
  AOI22_X1 U7313 ( .A1(n6333), .A2(n6355), .B1(n6353), .B2(n6332), .ZN(n6335)
         );
  NAND2_X1 U7314 ( .A1(n6351), .A2(REIP_REG_5__SCAN_IN), .ZN(n6334) );
  OAI211_X1 U7315 ( .C1(n6337), .C2(n6336), .A(n6335), .B(n6334), .ZN(U3013)
         );
  AOI21_X1 U7316 ( .B1(n6339), .B2(n6346), .A(n6338), .ZN(n6361) );
  OAI222_X1 U7317 ( .A1(n6343), .A2(n6342), .B1(n6341), .B2(n6542), .C1(n6283), 
        .C2(n6340), .ZN(n6344) );
  INV_X1 U7318 ( .A(n6344), .ZN(n6349) );
  NOR2_X1 U7319 ( .A1(n6346), .A2(n6345), .ZN(n6357) );
  OAI211_X1 U7320 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n6357), .B(n6347), .ZN(n6348) );
  OAI211_X1 U7321 ( .C1(n6361), .C2(n6350), .A(n6349), .B(n6348), .ZN(U3014)
         );
  AOI22_X1 U7322 ( .A1(n6353), .A2(n6352), .B1(n6351), .B2(REIP_REG_3__SCAN_IN), .ZN(n6359) );
  INV_X1 U7323 ( .A(n6354), .ZN(n6356) );
  AOI22_X1 U7324 ( .A1(n6357), .A2(n6360), .B1(n6356), .B2(n6355), .ZN(n6358)
         );
  OAI211_X1 U7325 ( .C1(n6361), .C2(n6360), .A(n6359), .B(n6358), .ZN(U3015)
         );
  INV_X1 U7326 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6476) );
  NOR2_X1 U7327 ( .A1(n6476), .A2(n6362), .ZN(U3019) );
  NAND2_X1 U7328 ( .A1(n6364), .A2(n6363), .ZN(n6377) );
  INV_X1 U7329 ( .A(n6377), .ZN(n6418) );
  INV_X1 U7330 ( .A(n6365), .ZN(n6370) );
  NAND3_X1 U7331 ( .A1(n6368), .A2(n6367), .A3(n6366), .ZN(n6369) );
  OAI21_X1 U7332 ( .B1(n6371), .B2(n6370), .A(n6369), .ZN(n6416) );
  AOI22_X1 U7333 ( .A1(n6372), .A2(n6418), .B1(n6456), .B2(n6416), .ZN(n6383)
         );
  INV_X1 U7334 ( .A(n6447), .ZN(n6373) );
  NOR3_X1 U7335 ( .A1(n6420), .A2(n6373), .A3(n5875), .ZN(n6376) );
  OAI21_X1 U7336 ( .B1(n6376), .B2(n6375), .A(n6374), .ZN(n6380) );
  AOI21_X1 U7337 ( .B1(n6377), .B2(STATE2_REG_3__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6378) );
  NAND3_X1 U7338 ( .A1(n6380), .A2(n6379), .A3(n6378), .ZN(n6422) );
  AOI22_X1 U7339 ( .A1(n6422), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6381), 
        .B2(n6420), .ZN(n6382) );
  OAI211_X1 U7340 ( .C1(n6452), .C2(n6447), .A(n6383), .B(n6382), .ZN(U3068)
         );
  AOI22_X1 U7341 ( .A1(n6385), .A2(n6418), .B1(n6384), .B2(n6416), .ZN(n6388)
         );
  AOI22_X1 U7342 ( .A1(n6422), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6386), 
        .B2(n6420), .ZN(n6387) );
  OAI211_X1 U7343 ( .C1(n6389), .C2(n6447), .A(n6388), .B(n6387), .ZN(U3069)
         );
  AOI22_X1 U7344 ( .A1(n6391), .A2(n6418), .B1(n6390), .B2(n6416), .ZN(n6394)
         );
  AOI22_X1 U7345 ( .A1(n6422), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6392), 
        .B2(n6420), .ZN(n6393) );
  OAI211_X1 U7346 ( .C1(n6395), .C2(n6447), .A(n6394), .B(n6393), .ZN(U3070)
         );
  AOI22_X1 U7347 ( .A1(n6396), .A2(n6418), .B1(n6433), .B2(n6416), .ZN(n6399)
         );
  AOI22_X1 U7348 ( .A1(n6422), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6397), 
        .B2(n6420), .ZN(n6398) );
  OAI211_X1 U7349 ( .C1(n6430), .C2(n6447), .A(n6399), .B(n6398), .ZN(U3071)
         );
  AOI22_X1 U7350 ( .A1(n6400), .A2(n6418), .B1(n6443), .B2(n6416), .ZN(n6403)
         );
  AOI22_X1 U7351 ( .A1(n6422), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6401), 
        .B2(n6420), .ZN(n6402) );
  OAI211_X1 U7352 ( .C1(n6437), .C2(n6447), .A(n6403), .B(n6402), .ZN(U3072)
         );
  AOI22_X1 U7353 ( .A1(n6405), .A2(n6418), .B1(n6404), .B2(n6416), .ZN(n6408)
         );
  AOI22_X1 U7354 ( .A1(n6422), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6406), 
        .B2(n6420), .ZN(n6407) );
  OAI211_X1 U7355 ( .C1(n6409), .C2(n6447), .A(n6408), .B(n6407), .ZN(U3073)
         );
  AOI22_X1 U7356 ( .A1(n6411), .A2(n6418), .B1(n6410), .B2(n6416), .ZN(n6414)
         );
  AOI22_X1 U7357 ( .A1(n6422), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6412), 
        .B2(n6420), .ZN(n6413) );
  OAI211_X1 U7358 ( .C1(n6415), .C2(n6447), .A(n6414), .B(n6413), .ZN(U3074)
         );
  AOI22_X1 U7359 ( .A1(n6419), .A2(n6418), .B1(n6417), .B2(n6416), .ZN(n6424)
         );
  AOI22_X1 U7360 ( .A1(n6422), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6421), 
        .B2(n6420), .ZN(n6423) );
  OAI211_X1 U7361 ( .C1(n6425), .C2(n6447), .A(n6424), .B(n6423), .ZN(U3075)
         );
  OAI22_X1 U7362 ( .A1(n6451), .A2(n6439), .B1(n6438), .B2(n6452), .ZN(n6426)
         );
  INV_X1 U7363 ( .A(n6426), .ZN(n6429) );
  INV_X1 U7364 ( .A(n6427), .ZN(n6442) );
  AOI22_X1 U7365 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6444), .B1(n6456), 
        .B2(n6442), .ZN(n6428) );
  OAI211_X1 U7366 ( .C1(n6461), .C2(n6447), .A(n6429), .B(n6428), .ZN(U3076)
         );
  OAI22_X1 U7367 ( .A1(n6431), .A2(n6439), .B1(n6438), .B2(n6430), .ZN(n6432)
         );
  INV_X1 U7368 ( .A(n6432), .ZN(n6435) );
  AOI22_X1 U7369 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6444), .B1(n6433), 
        .B2(n6442), .ZN(n6434) );
  OAI211_X1 U7370 ( .C1(n6436), .C2(n6447), .A(n6435), .B(n6434), .ZN(U3079)
         );
  OAI22_X1 U7371 ( .A1(n6440), .A2(n6439), .B1(n6438), .B2(n6437), .ZN(n6441)
         );
  INV_X1 U7372 ( .A(n6441), .ZN(n6446) );
  AOI22_X1 U7373 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6444), .B1(n6443), 
        .B2(n6442), .ZN(n6445) );
  OAI211_X1 U7374 ( .C1(n6448), .C2(n6447), .A(n6446), .B(n6445), .ZN(U3080)
         );
  INV_X1 U7375 ( .A(n6449), .ZN(n6450) );
  OAI22_X1 U7376 ( .A1(n6453), .A2(n6452), .B1(n6451), .B2(n6450), .ZN(n6454)
         );
  INV_X1 U7377 ( .A(n6454), .ZN(n6459) );
  AOI22_X1 U7378 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6457), .B1(n6456), 
        .B2(n6455), .ZN(n6458) );
  OAI211_X1 U7379 ( .C1(n6461), .C2(n6460), .A(n6459), .B(n6458), .ZN(U3108)
         );
  MUX2_X1 U7380 ( .A(n6463), .B(n6462), .S(INSTQUEUERD_ADDR_REG_0__SCAN_IN), 
        .Z(n6464) );
  AND3_X1 U7381 ( .A1(n6465), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n6464), 
        .ZN(n6469) );
  NAND2_X1 U7382 ( .A1(n6467), .A2(n6466), .ZN(n6468) );
  AOI222_X1 U7383 ( .A1(n6469), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n6469), .B2(n6468), .C1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n6468), 
        .ZN(n6472) );
  AOI21_X1 U7384 ( .B1(n6472), .B2(n6471), .A(n6470), .ZN(n6475) );
  NOR2_X1 U7385 ( .A1(n6472), .A2(n6471), .ZN(n6474) );
  OAI22_X1 U7386 ( .A1(n6475), .A2(n6474), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n6473), .ZN(n6477) );
  OAI211_X1 U7387 ( .C1(n6479), .C2(n6478), .A(n6477), .B(n6476), .ZN(n6480)
         );
  INV_X1 U7388 ( .A(n6480), .ZN(n6488) );
  OAI21_X1 U7389 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6481), 
        .ZN(n6482) );
  NAND3_X1 U7390 ( .A1(n6484), .A2(n6483), .A3(n6482), .ZN(n6485) );
  NOR4_X1 U7391 ( .A1(n6488), .A2(n6487), .A3(n6486), .A4(n6485), .ZN(n6504)
         );
  AOI21_X1 U7392 ( .B1(n6491), .B2(n6490), .A(n6489), .ZN(n6503) );
  INV_X1 U7393 ( .A(n6504), .ZN(n6493) );
  OAI22_X1 U7394 ( .A1(n6493), .A2(n6505), .B1(n6735), .B2(n6492), .ZN(n6494)
         );
  OAI21_X1 U7395 ( .B1(n6496), .B2(n6495), .A(n6494), .ZN(n6591) );
  AOI21_X1 U7396 ( .B1(n6613), .B2(n6497), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n6501) );
  NAND2_X1 U7397 ( .A1(READY_N), .A2(n6498), .ZN(n6513) );
  AOI21_X1 U7398 ( .B1(n6513), .B2(n6591), .A(n6499), .ZN(n6500) );
  AOI21_X1 U7399 ( .B1(n6591), .B2(n6501), .A(n6500), .ZN(n6502) );
  OAI211_X1 U7400 ( .C1(n6504), .C2(n6505), .A(n6503), .B(n6502), .ZN(U3148)
         );
  OAI21_X1 U7401 ( .B1(READY_N), .B2(n6506), .A(n6505), .ZN(n6510) );
  NOR2_X1 U7402 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6512) );
  AOI211_X1 U7403 ( .C1(n6591), .C2(n6513), .A(n6512), .B(n6507), .ZN(n6508)
         );
  AOI211_X1 U7404 ( .C1(n6591), .C2(n6510), .A(n6509), .B(n6508), .ZN(n6511)
         );
  INV_X1 U7405 ( .A(n6511), .ZN(U3149) );
  INV_X1 U7406 ( .A(n6512), .ZN(n6515) );
  NAND4_X1 U7407 ( .A1(n6515), .A2(n6514), .A3(n6513), .A4(n6589), .ZN(n6516)
         );
  NAND2_X1 U7408 ( .A1(n6517), .A2(n6516), .ZN(U3150) );
  AND2_X1 U7409 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6518), .ZN(U3151) );
  AND2_X1 U7410 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6518), .ZN(U3152) );
  AND2_X1 U7411 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6518), .ZN(U3153) );
  AND2_X1 U7412 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6518), .ZN(U3154) );
  AND2_X1 U7413 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6518), .ZN(U3155) );
  AND2_X1 U7414 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6518), .ZN(U3156) );
  AND2_X1 U7415 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6518), .ZN(U3157) );
  AND2_X1 U7416 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6518), .ZN(U3158) );
  AND2_X1 U7417 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6518), .ZN(U3159) );
  AND2_X1 U7418 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6518), .ZN(U3160) );
  AND2_X1 U7419 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6518), .ZN(U3161) );
  AND2_X1 U7420 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6518), .ZN(U3162) );
  AND2_X1 U7421 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6518), .ZN(U3163) );
  AND2_X1 U7422 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6518), .ZN(U3164) );
  AND2_X1 U7423 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6518), .ZN(U3165) );
  AND2_X1 U7424 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6518), .ZN(U3166) );
  AND2_X1 U7425 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6518), .ZN(U3167) );
  AND2_X1 U7426 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6518), .ZN(U3168) );
  AND2_X1 U7427 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6518), .ZN(U3169) );
  AND2_X1 U7428 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6518), .ZN(U3170) );
  AND2_X1 U7429 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6518), .ZN(U3171) );
  AND2_X1 U7430 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6518), .ZN(U3172) );
  AND2_X1 U7431 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6518), .ZN(U3173) );
  AND2_X1 U7432 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6518), .ZN(U3174) );
  AND2_X1 U7433 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6518), .ZN(U3175) );
  AND2_X1 U7434 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6518), .ZN(U3176) );
  AND2_X1 U7435 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6518), .ZN(U3177) );
  AND2_X1 U7436 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6518), .ZN(U3178) );
  AND2_X1 U7437 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6518), .ZN(U3179) );
  AND2_X1 U7438 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6518), .ZN(U3180) );
  INV_X1 U7439 ( .A(n6534), .ZN(n6520) );
  NAND2_X1 U7440 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .ZN(n6522) );
  INV_X1 U7441 ( .A(n6522), .ZN(n6531) );
  AOI21_X1 U7442 ( .B1(HOLD), .B2(STATE_REG_2__SCAN_IN), .A(n6531), .ZN(n6535)
         );
  INV_X1 U7443 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6526) );
  INV_X1 U7444 ( .A(HOLD), .ZN(n6742) );
  NOR2_X1 U7445 ( .A1(n6526), .A2(n6742), .ZN(n6521) );
  INV_X1 U7446 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6762) );
  OAI21_X1 U7447 ( .B1(n6521), .B2(n6762), .A(n6819), .ZN(n6519) );
  OAI211_X1 U7448 ( .C1(NA_N), .C2(n6536), .A(n6530), .B(n6534), .ZN(n6528) );
  OAI211_X1 U7449 ( .C1(n6520), .C2(n6535), .A(n6519), .B(n6528), .ZN(U3181)
         );
  NOR2_X1 U7450 ( .A1(n6536), .A2(n6742), .ZN(n6525) );
  AOI21_X1 U7451 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(STATE_REG_0__SCAN_IN), 
        .A(n6521), .ZN(n6524) );
  OAI211_X1 U7452 ( .C1(n6525), .C2(n6524), .A(n6523), .B(n6522), .ZN(U3182)
         );
  INV_X1 U7453 ( .A(NA_N), .ZN(n6749) );
  OAI221_X1 U7454 ( .B1(n6526), .B2(READY_N), .C1(n6526), .C2(n6749), .A(n6762), .ZN(n6527) );
  AOI21_X1 U7455 ( .B1(n6536), .B2(n6527), .A(n6742), .ZN(n6529) );
  OAI21_X1 U7456 ( .B1(n6530), .B2(n6529), .A(n6528), .ZN(n6533) );
  NAND4_X1 U7457 ( .A1(REQUESTPENDING_REG_SCAN_IN), .A2(STATE_REG_0__SCAN_IN), 
        .A3(n6531), .A4(n6749), .ZN(n6532) );
  OAI211_X1 U7458 ( .C1(n6535), .C2(n6534), .A(n6533), .B(n6532), .ZN(U3183)
         );
  NOR2_X2 U7459 ( .A1(n6536), .A2(n6819), .ZN(n6576) );
  NAND2_X1 U7460 ( .A1(n6536), .A2(n6820), .ZN(n6578) );
  INV_X1 U7461 ( .A(n6578), .ZN(n6582) );
  AOI22_X1 U7462 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6582), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6819), .ZN(n6537) );
  OAI21_X1 U7463 ( .B1(n6600), .B2(n6584), .A(n6537), .ZN(U3184) );
  AOI22_X1 U7464 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6576), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6819), .ZN(n6538) );
  OAI21_X1 U7465 ( .B1(n6539), .B2(n6578), .A(n6538), .ZN(U3185) );
  AOI22_X1 U7466 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6576), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6819), .ZN(n6540) );
  OAI21_X1 U7467 ( .B1(n6542), .B2(n6578), .A(n6540), .ZN(U3186) );
  AOI22_X1 U7468 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6582), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6819), .ZN(n6541) );
  OAI21_X1 U7469 ( .B1(n6542), .B2(n6584), .A(n6541), .ZN(U3187) );
  AOI22_X1 U7470 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6576), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6819), .ZN(n6543) );
  OAI21_X1 U7471 ( .B1(n6545), .B2(n6578), .A(n6543), .ZN(U3188) );
  AOI22_X1 U7472 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6582), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6819), .ZN(n6544) );
  OAI21_X1 U7473 ( .B1(n6545), .B2(n6584), .A(n6544), .ZN(U3189) );
  AOI22_X1 U7474 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6576), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6819), .ZN(n6546) );
  OAI21_X1 U7475 ( .B1(n6548), .B2(n6578), .A(n6546), .ZN(U3190) );
  AOI22_X1 U7476 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6582), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6819), .ZN(n6547) );
  OAI21_X1 U7477 ( .B1(n6548), .B2(n6584), .A(n6547), .ZN(U3191) );
  AOI22_X1 U7478 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6582), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6819), .ZN(n6549) );
  OAI21_X1 U7479 ( .B1(n6550), .B2(n6584), .A(n6549), .ZN(U3192) );
  AOI22_X1 U7480 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6576), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6819), .ZN(n6551) );
  OAI21_X1 U7481 ( .B1(n6552), .B2(n6578), .A(n6551), .ZN(U3193) );
  AOI22_X1 U7482 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6576), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6819), .ZN(n6553) );
  OAI21_X1 U7483 ( .B1(n6555), .B2(n6578), .A(n6553), .ZN(U3194) );
  AOI22_X1 U7484 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6582), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6819), .ZN(n6554) );
  OAI21_X1 U7485 ( .B1(n6555), .B2(n6584), .A(n6554), .ZN(U3195) );
  AOI22_X1 U7486 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6582), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6819), .ZN(n6556) );
  OAI21_X1 U7487 ( .B1(n6557), .B2(n6584), .A(n6556), .ZN(U3196) );
  AOI22_X1 U7488 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6576), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6819), .ZN(n6558) );
  OAI21_X1 U7489 ( .B1(n6560), .B2(n6578), .A(n6558), .ZN(U3197) );
  AOI22_X1 U7490 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6582), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6819), .ZN(n6559) );
  OAI21_X1 U7491 ( .B1(n6560), .B2(n6584), .A(n6559), .ZN(U3198) );
  AOI22_X1 U7492 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6582), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6819), .ZN(n6561) );
  OAI21_X1 U7493 ( .B1(n6562), .B2(n6584), .A(n6561), .ZN(U3199) );
  AOI22_X1 U7494 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6576), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6819), .ZN(n6563) );
  OAI21_X1 U7495 ( .B1(n6565), .B2(n6578), .A(n6563), .ZN(U3200) );
  AOI22_X1 U7496 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6582), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6819), .ZN(n6564) );
  OAI21_X1 U7497 ( .B1(n6565), .B2(n6584), .A(n6564), .ZN(U3201) );
  AOI22_X1 U7498 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6576), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6819), .ZN(n6566) );
  OAI21_X1 U7499 ( .B1(n6713), .B2(n6578), .A(n6566), .ZN(U3202) );
  AOI22_X1 U7500 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6582), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6819), .ZN(n6567) );
  OAI21_X1 U7501 ( .B1(n6713), .B2(n6584), .A(n6567), .ZN(U3203) );
  AOI22_X1 U7502 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6582), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6819), .ZN(n6568) );
  OAI21_X1 U7503 ( .B1(n6569), .B2(n6584), .A(n6568), .ZN(U3204) );
  AOI22_X1 U7504 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6576), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6819), .ZN(n6570) );
  OAI21_X1 U7505 ( .B1(n6660), .B2(n6578), .A(n6570), .ZN(U3205) );
  AOI22_X1 U7506 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6582), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6819), .ZN(n6571) );
  OAI21_X1 U7507 ( .B1(n6660), .B2(n6584), .A(n6571), .ZN(U3206) );
  AOI22_X1 U7508 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6576), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6819), .ZN(n6572) );
  OAI21_X1 U7509 ( .B1(n6573), .B2(n6578), .A(n6572), .ZN(U3207) );
  AOI22_X1 U7510 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6576), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6819), .ZN(n6574) );
  OAI21_X1 U7511 ( .B1(n6650), .B2(n6578), .A(n6574), .ZN(U3208) );
  AOI22_X1 U7512 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6582), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6819), .ZN(n6575) );
  OAI21_X1 U7513 ( .B1(n6650), .B2(n6584), .A(n6575), .ZN(U3209) );
  AOI22_X1 U7514 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6576), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6819), .ZN(n6577) );
  OAI21_X1 U7515 ( .B1(n6580), .B2(n6578), .A(n6577), .ZN(U3210) );
  AOI22_X1 U7516 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6582), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6819), .ZN(n6579) );
  OAI21_X1 U7517 ( .B1(n6580), .B2(n6584), .A(n6579), .ZN(U3211) );
  AOI22_X1 U7518 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6582), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6819), .ZN(n6581) );
  OAI21_X1 U7519 ( .B1(n6767), .B2(n6584), .A(n6581), .ZN(U3212) );
  AOI22_X1 U7520 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6582), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6819), .ZN(n6583) );
  OAI21_X1 U7521 ( .B1(n6716), .B2(n6584), .A(n6583), .ZN(U3213) );
  MUX2_X1 U7522 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6819), .Z(U3446) );
  MUX2_X1 U7523 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6819), .Z(U3447) );
  MUX2_X1 U7524 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6819), .Z(U3448) );
  OAI21_X1 U7525 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6588), .A(n6586), .ZN(
        n6585) );
  INV_X1 U7526 ( .A(n6585), .ZN(U3451) );
  OAI21_X1 U7527 ( .B1(n6588), .B2(n6587), .A(n6586), .ZN(U3452) );
  OAI211_X1 U7528 ( .C1(n6592), .C2(n6591), .A(n6590), .B(n6589), .ZN(U3453)
         );
  INV_X1 U7529 ( .A(n6593), .ZN(n6596) );
  OAI22_X1 U7530 ( .A1(n6597), .A2(n6596), .B1(n6595), .B2(n6594), .ZN(n6599)
         );
  MUX2_X1 U7531 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6599), .S(n6598), 
        .Z(U3456) );
  AOI21_X1 U7532 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6601) );
  AOI22_X1 U7533 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6601), .B2(n6600), .ZN(n6602) );
  INV_X1 U7534 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6759) );
  AOI22_X1 U7535 ( .A1(n6603), .A2(n6602), .B1(n6759), .B2(n6606), .ZN(U3468)
         );
  INV_X1 U7536 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6607) );
  NOR2_X1 U7537 ( .A1(n6606), .A2(REIP_REG_1__SCAN_IN), .ZN(n6604) );
  AOI22_X1 U7538 ( .A1(n6607), .A2(n6606), .B1(n6605), .B2(n6604), .ZN(U3469)
         );
  OAI22_X1 U7539 ( .A1(n6819), .A2(n6657), .B1(W_R_N_REG_SCAN_IN), .B2(n6820), 
        .ZN(n6608) );
  INV_X1 U7540 ( .A(n6608), .ZN(U3470) );
  AOI211_X1 U7541 ( .C1(n6243), .C2(n6735), .A(n6610), .B(n6609), .ZN(n6617)
         );
  OAI211_X1 U7542 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6612), .A(n6611), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6614) );
  AOI21_X1 U7543 ( .B1(n6614), .B2(STATE2_REG_0__SCAN_IN), .A(n6613), .ZN(
        n6616) );
  NAND2_X1 U7544 ( .A1(n6617), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6615) );
  OAI21_X1 U7545 ( .B1(n6617), .B2(n6616), .A(n6615), .ZN(U3472) );
  INV_X1 U7546 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n6761) );
  AOI22_X1 U7547 ( .A1(n6820), .A2(n4213), .B1(n6761), .B2(n6819), .ZN(U3473)
         );
  INV_X1 U7548 ( .A(keyinput_f24), .ZN(n6710) );
  AOI22_X1 U7549 ( .A1(DATAI_10_), .A2(keyinput_f21), .B1(REIP_REG_28__SCAN_IN), .B2(keyinput_f54), .ZN(n6618) );
  OAI221_X1 U7550 ( .B1(DATAI_10_), .B2(keyinput_f21), .C1(
        REIP_REG_28__SCAN_IN), .C2(keyinput_f54), .A(n6618), .ZN(n6708) );
  AOI22_X1 U7551 ( .A1(REIP_REG_25__SCAN_IN), .A2(keyinput_f57), .B1(
        REIP_REG_22__SCAN_IN), .B2(keyinput_f60), .ZN(n6619) );
  OAI221_X1 U7552 ( .B1(REIP_REG_25__SCAN_IN), .B2(keyinput_f57), .C1(
        REIP_REG_22__SCAN_IN), .C2(keyinput_f60), .A(n6619), .ZN(n6707) );
  AOI22_X1 U7553 ( .A1(keyinput_f34), .A2(BS16_N), .B1(n6621), .B2(
        keyinput_f25), .ZN(n6620) );
  OAI221_X1 U7554 ( .B1(keyinput_f34), .B2(BS16_N), .C1(n6621), .C2(
        keyinput_f25), .A(n6620), .ZN(n6631) );
  OAI22_X1 U7555 ( .A1(DATAI_2_), .A2(keyinput_f29), .B1(keyinput_f40), .B2(
        M_IO_N_REG_SCAN_IN), .ZN(n6622) );
  AOI221_X1 U7556 ( .B1(DATAI_2_), .B2(keyinput_f29), .C1(M_IO_N_REG_SCAN_IN), 
        .C2(keyinput_f40), .A(n6622), .ZN(n6629) );
  OAI22_X1 U7557 ( .A1(DATAI_23_), .A2(keyinput_f8), .B1(keyinput_f13), .B2(
        DATAI_18_), .ZN(n6623) );
  AOI221_X1 U7558 ( .B1(DATAI_23_), .B2(keyinput_f8), .C1(DATAI_18_), .C2(
        keyinput_f13), .A(n6623), .ZN(n6628) );
  OAI22_X1 U7559 ( .A1(REIP_REG_21__SCAN_IN), .A2(keyinput_f61), .B1(
        keyinput_f10), .B2(DATAI_21_), .ZN(n6624) );
  AOI221_X1 U7560 ( .B1(REIP_REG_21__SCAN_IN), .B2(keyinput_f61), .C1(
        DATAI_21_), .C2(keyinput_f10), .A(n6624), .ZN(n6627) );
  OAI22_X1 U7561 ( .A1(REIP_REG_30__SCAN_IN), .A2(keyinput_f52), .B1(
        REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_f42), .ZN(n6625) );
  AOI221_X1 U7562 ( .B1(REIP_REG_30__SCAN_IN), .B2(keyinput_f52), .C1(
        keyinput_f42), .C2(REQUESTPENDING_REG_SCAN_IN), .A(n6625), .ZN(n6626)
         );
  NAND4_X1 U7563 ( .A1(n6629), .A2(n6628), .A3(n6627), .A4(n6626), .ZN(n6630)
         );
  AOI211_X1 U7564 ( .C1(keyinput_f62), .C2(REIP_REG_20__SCAN_IN), .A(n6631), 
        .B(n6630), .ZN(n6632) );
  OAI21_X1 U7565 ( .B1(keyinput_f62), .B2(REIP_REG_20__SCAN_IN), .A(n6632), 
        .ZN(n6706) );
  AOI22_X1 U7566 ( .A1(keyinput_f46), .A2(W_R_N_REG_SCAN_IN), .B1(
        MORE_REG_SCAN_IN), .B2(keyinput_f44), .ZN(n6633) );
  OAI221_X1 U7567 ( .B1(keyinput_f46), .B2(W_R_N_REG_SCAN_IN), .C1(
        MORE_REG_SCAN_IN), .C2(keyinput_f44), .A(n6633), .ZN(n6640) );
  AOI22_X1 U7568 ( .A1(keyinput_f41), .A2(D_C_N_REG_SCAN_IN), .B1(
        REIP_REG_24__SCAN_IN), .B2(keyinput_f58), .ZN(n6634) );
  OAI221_X1 U7569 ( .B1(keyinput_f41), .B2(D_C_N_REG_SCAN_IN), .C1(
        REIP_REG_24__SCAN_IN), .C2(keyinput_f58), .A(n6634), .ZN(n6639) );
  AOI22_X1 U7570 ( .A1(DATAI_4_), .A2(keyinput_f27), .B1(DATAI_31_), .B2(
        keyinput_f0), .ZN(n6635) );
  OAI221_X1 U7571 ( .B1(DATAI_4_), .B2(keyinput_f27), .C1(DATAI_31_), .C2(
        keyinput_f0), .A(n6635), .ZN(n6638) );
  AOI22_X1 U7572 ( .A1(keyinput_f38), .A2(ADS_N_REG_SCAN_IN), .B1(keyinput_f50), .B2(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6636) );
  OAI221_X1 U7573 ( .B1(keyinput_f38), .B2(ADS_N_REG_SCAN_IN), .C1(
        keyinput_f50), .C2(BYTEENABLE_REG_3__SCAN_IN), .A(n6636), .ZN(n6637)
         );
  NOR4_X1 U7574 ( .A1(n6640), .A2(n6639), .A3(n6638), .A4(n6637), .ZN(n6704)
         );
  AOI22_X1 U7575 ( .A1(DATAI_3_), .A2(keyinput_f28), .B1(REIP_REG_31__SCAN_IN), 
        .B2(keyinput_f51), .ZN(n6641) );
  OAI221_X1 U7576 ( .B1(DATAI_3_), .B2(keyinput_f28), .C1(REIP_REG_31__SCAN_IN), .C2(keyinput_f51), .A(n6641), .ZN(n6648) );
  AOI22_X1 U7577 ( .A1(keyinput_f36), .A2(HOLD), .B1(DATAI_22_), .B2(
        keyinput_f9), .ZN(n6642) );
  OAI221_X1 U7578 ( .B1(keyinput_f36), .B2(HOLD), .C1(DATAI_22_), .C2(
        keyinput_f9), .A(n6642), .ZN(n6647) );
  AOI22_X1 U7579 ( .A1(DATAI_1_), .A2(keyinput_f30), .B1(DATAI_24_), .B2(
        keyinput_f7), .ZN(n6643) );
  OAI221_X1 U7580 ( .B1(DATAI_1_), .B2(keyinput_f30), .C1(DATAI_24_), .C2(
        keyinput_f7), .A(n6643), .ZN(n6646) );
  AOI22_X1 U7581 ( .A1(DATAI_19_), .A2(keyinput_f12), .B1(DATAI_25_), .B2(
        keyinput_f6), .ZN(n6644) );
  OAI221_X1 U7582 ( .B1(DATAI_19_), .B2(keyinput_f12), .C1(DATAI_25_), .C2(
        keyinput_f6), .A(n6644), .ZN(n6645) );
  NOR4_X1 U7583 ( .A1(n6648), .A2(n6647), .A3(n6646), .A4(n6645), .ZN(n6703)
         );
  XNOR2_X1 U7584 ( .A(keyinput_f48), .B(n6729), .ZN(n6652) );
  AOI22_X1 U7585 ( .A1(n6746), .A2(keyinput_f2), .B1(n6650), .B2(keyinput_f56), 
        .ZN(n6649) );
  OAI221_X1 U7586 ( .B1(n6746), .B2(keyinput_f2), .C1(n6650), .C2(keyinput_f56), .A(n6649), .ZN(n6651) );
  AOI211_X1 U7587 ( .C1(n4213), .C2(keyinput_f32), .A(n6652), .B(n6651), .ZN(
        n6653) );
  OAI21_X1 U7588 ( .B1(n4213), .B2(keyinput_f32), .A(n6653), .ZN(n6673) );
  INV_X1 U7589 ( .A(DATAI_11_), .ZN(n6748) );
  AOI22_X1 U7590 ( .A1(n6735), .A2(keyinput_f35), .B1(keyinput_f20), .B2(n6748), .ZN(n6654) );
  OAI221_X1 U7591 ( .B1(n6735), .B2(keyinput_f35), .C1(n6748), .C2(
        keyinput_f20), .A(n6654), .ZN(n6672) );
  INV_X1 U7592 ( .A(DATAI_14_), .ZN(n6656) );
  AOI22_X1 U7593 ( .A1(n6657), .A2(keyinput_f37), .B1(n6656), .B2(keyinput_f17), .ZN(n6655) );
  OAI221_X1 U7594 ( .B1(n6657), .B2(keyinput_f37), .C1(n6656), .C2(
        keyinput_f17), .A(n6655), .ZN(n6671) );
  INV_X1 U7595 ( .A(DATAI_8_), .ZN(n6659) );
  OAI22_X1 U7596 ( .A1(n6660), .A2(keyinput_f59), .B1(n6659), .B2(keyinput_f23), .ZN(n6658) );
  AOI221_X1 U7597 ( .B1(n6660), .B2(keyinput_f59), .C1(keyinput_f23), .C2(
        n6659), .A(n6658), .ZN(n6669) );
  INV_X1 U7598 ( .A(DATAI_13_), .ZN(n6719) );
  OAI22_X1 U7599 ( .A1(n6719), .A2(keyinput_f18), .B1(keyinput_f53), .B2(
        REIP_REG_29__SCAN_IN), .ZN(n6661) );
  AOI221_X1 U7600 ( .B1(n6719), .B2(keyinput_f18), .C1(REIP_REG_29__SCAN_IN), 
        .C2(keyinput_f53), .A(n6661), .ZN(n6668) );
  INV_X1 U7601 ( .A(DATAI_28_), .ZN(n6732) );
  INV_X1 U7602 ( .A(DATAI_9_), .ZN(n6785) );
  OAI22_X1 U7603 ( .A1(n6732), .A2(keyinput_f3), .B1(n6785), .B2(keyinput_f22), 
        .ZN(n6662) );
  AOI221_X1 U7604 ( .B1(n6732), .B2(keyinput_f3), .C1(keyinput_f22), .C2(n6785), .A(n6662), .ZN(n6667) );
  INV_X1 U7605 ( .A(DATAI_17_), .ZN(n6665) );
  INV_X1 U7606 ( .A(keyinput_f47), .ZN(n6664) );
  OAI22_X1 U7607 ( .A1(n6665), .A2(keyinput_f14), .B1(n6664), .B2(
        BYTEENABLE_REG_0__SCAN_IN), .ZN(n6663) );
  AOI221_X1 U7608 ( .B1(n6665), .B2(keyinput_f14), .C1(
        BYTEENABLE_REG_0__SCAN_IN), .C2(n6664), .A(n6663), .ZN(n6666) );
  NAND4_X1 U7609 ( .A1(n6669), .A2(n6668), .A3(n6667), .A4(n6666), .ZN(n6670)
         );
  NOR4_X1 U7610 ( .A1(n6673), .A2(n6672), .A3(n6671), .A4(n6670), .ZN(n6702)
         );
  XNOR2_X1 U7611 ( .A(keyinput_f33), .B(n6749), .ZN(n6677) );
  AOI22_X1 U7612 ( .A1(n6733), .A2(keyinput_f26), .B1(n6675), .B2(keyinput_f1), 
        .ZN(n6674) );
  OAI221_X1 U7613 ( .B1(n6733), .B2(keyinput_f26), .C1(n6675), .C2(keyinput_f1), .A(n6674), .ZN(n6676) );
  AOI211_X1 U7614 ( .C1(n6759), .C2(keyinput_f49), .A(n6677), .B(n6676), .ZN(
        n6678) );
  OAI21_X1 U7615 ( .B1(n6759), .B2(keyinput_f49), .A(n6678), .ZN(n6700) );
  INV_X1 U7616 ( .A(DATAI_16_), .ZN(n6764) );
  AOI22_X1 U7617 ( .A1(n6764), .A2(keyinput_f15), .B1(n6787), .B2(keyinput_f31), .ZN(n6679) );
  OAI221_X1 U7618 ( .B1(n6764), .B2(keyinput_f15), .C1(n6787), .C2(
        keyinput_f31), .A(n6679), .ZN(n6699) );
  INV_X1 U7619 ( .A(DATAI_27_), .ZN(n6681) );
  AOI22_X1 U7620 ( .A1(n6682), .A2(keyinput_f63), .B1(keyinput_f4), .B2(n6681), 
        .ZN(n6680) );
  OAI221_X1 U7621 ( .B1(n6682), .B2(keyinput_f63), .C1(n6681), .C2(keyinput_f4), .A(n6680), .ZN(n6698) );
  OAI22_X1 U7622 ( .A1(n6684), .A2(keyinput_f5), .B1(n6718), .B2(keyinput_f45), 
        .ZN(n6683) );
  AOI221_X1 U7623 ( .B1(n6684), .B2(keyinput_f5), .C1(keyinput_f45), .C2(n6718), .A(n6683), .ZN(n6696) );
  INV_X1 U7624 ( .A(DATAI_12_), .ZN(n6687) );
  OAI22_X1 U7625 ( .A1(n6687), .A2(keyinput_f19), .B1(n6686), .B2(keyinput_f16), .ZN(n6685) );
  AOI221_X1 U7626 ( .B1(n6687), .B2(keyinput_f19), .C1(keyinput_f16), .C2(
        n6686), .A(n6685), .ZN(n6695) );
  INV_X1 U7627 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6689) );
  OAI22_X1 U7628 ( .A1(n6728), .A2(keyinput_f43), .B1(n6689), .B2(keyinput_f39), .ZN(n6688) );
  AOI221_X1 U7629 ( .B1(n6728), .B2(keyinput_f43), .C1(keyinput_f39), .C2(
        n6689), .A(n6688), .ZN(n6694) );
  INV_X1 U7630 ( .A(DATAI_20_), .ZN(n6691) );
  OAI22_X1 U7631 ( .A1(n6692), .A2(keyinput_f55), .B1(n6691), .B2(keyinput_f11), .ZN(n6690) );
  AOI221_X1 U7632 ( .B1(n6692), .B2(keyinput_f55), .C1(keyinput_f11), .C2(
        n6691), .A(n6690), .ZN(n6693) );
  NAND4_X1 U7633 ( .A1(n6696), .A2(n6695), .A3(n6694), .A4(n6693), .ZN(n6697)
         );
  NOR4_X1 U7634 ( .A1(n6700), .A2(n6699), .A3(n6698), .A4(n6697), .ZN(n6701)
         );
  NAND4_X1 U7635 ( .A1(n6704), .A2(n6703), .A3(n6702), .A4(n6701), .ZN(n6705)
         );
  NOR4_X1 U7636 ( .A1(n6708), .A2(n6707), .A3(n6706), .A4(n6705), .ZN(n6709)
         );
  AOI221_X1 U7637 ( .B1(DATAI_7_), .B2(keyinput_f24), .C1(n6818), .C2(n6710), 
        .A(n6709), .ZN(n6817) );
  AOI22_X1 U7638 ( .A1(n6713), .A2(keyinput_g62), .B1(keyinput_g30), .B2(n6712), .ZN(n6711) );
  OAI221_X1 U7639 ( .B1(n6713), .B2(keyinput_g62), .C1(n6712), .C2(
        keyinput_g30), .A(n6711), .ZN(n6726) );
  AOI22_X1 U7640 ( .A1(n6716), .A2(keyinput_g52), .B1(keyinput_g58), .B2(n6715), .ZN(n6714) );
  OAI221_X1 U7641 ( .B1(n6716), .B2(keyinput_g52), .C1(n6715), .C2(
        keyinput_g58), .A(n6714), .ZN(n6725) );
  AOI22_X1 U7642 ( .A1(n6719), .A2(keyinput_g18), .B1(keyinput_g45), .B2(n6718), .ZN(n6717) );
  OAI221_X1 U7643 ( .B1(n6719), .B2(keyinput_g18), .C1(n6718), .C2(
        keyinput_g45), .A(n6717), .ZN(n6724) );
  INV_X1 U7644 ( .A(DATAI_24_), .ZN(n6722) );
  AOI22_X1 U7645 ( .A1(n6722), .A2(keyinput_g7), .B1(keyinput_g28), .B2(n6721), 
        .ZN(n6720) );
  OAI221_X1 U7646 ( .B1(n6722), .B2(keyinput_g7), .C1(n6721), .C2(keyinput_g28), .A(n6720), .ZN(n6723) );
  NOR4_X1 U7647 ( .A1(n6726), .A2(n6725), .A3(n6724), .A4(n6723), .ZN(n6776)
         );
  AOI22_X1 U7648 ( .A1(n6729), .A2(keyinput_g48), .B1(n6728), .B2(keyinput_g43), .ZN(n6727) );
  OAI221_X1 U7649 ( .B1(n6729), .B2(keyinput_g48), .C1(n6728), .C2(
        keyinput_g43), .A(n6727), .ZN(n6740) );
  AOI22_X1 U7650 ( .A1(READREQUEST_REG_SCAN_IN), .A2(keyinput_g37), .B1(
        REIP_REG_22__SCAN_IN), .B2(keyinput_g60), .ZN(n6730) );
  OAI221_X1 U7651 ( .B1(READREQUEST_REG_SCAN_IN), .B2(keyinput_g37), .C1(
        REIP_REG_22__SCAN_IN), .C2(keyinput_g60), .A(n6730), .ZN(n6739) );
  AOI22_X1 U7652 ( .A1(n6733), .A2(keyinput_g26), .B1(n6732), .B2(keyinput_g3), 
        .ZN(n6731) );
  OAI221_X1 U7653 ( .B1(n6733), .B2(keyinput_g26), .C1(n6732), .C2(keyinput_g3), .A(n6731), .ZN(n6738) );
  INV_X1 U7654 ( .A(DATAI_19_), .ZN(n6736) );
  AOI22_X1 U7655 ( .A1(n6736), .A2(keyinput_g12), .B1(n6735), .B2(keyinput_g35), .ZN(n6734) );
  OAI221_X1 U7656 ( .B1(n6736), .B2(keyinput_g12), .C1(n6735), .C2(
        keyinput_g35), .A(n6734), .ZN(n6737) );
  NOR4_X1 U7657 ( .A1(n6740), .A2(n6739), .A3(n6738), .A4(n6737), .ZN(n6775)
         );
  INV_X1 U7658 ( .A(DATAI_10_), .ZN(n6743) );
  AOI22_X1 U7659 ( .A1(n6743), .A2(keyinput_g21), .B1(keyinput_g36), .B2(n6742), .ZN(n6741) );
  OAI221_X1 U7660 ( .B1(n6743), .B2(keyinput_g21), .C1(n6742), .C2(
        keyinput_g36), .A(n6741), .ZN(n6756) );
  AOI22_X1 U7661 ( .A1(n6746), .A2(keyinput_g2), .B1(n6745), .B2(keyinput_g0), 
        .ZN(n6744) );
  OAI221_X1 U7662 ( .B1(n6746), .B2(keyinput_g2), .C1(n6745), .C2(keyinput_g0), 
        .A(n6744), .ZN(n6755) );
  AOI22_X1 U7663 ( .A1(n6749), .A2(keyinput_g33), .B1(n6748), .B2(keyinput_g20), .ZN(n6747) );
  OAI221_X1 U7664 ( .B1(n6749), .B2(keyinput_g33), .C1(n6748), .C2(
        keyinput_g20), .A(n6747), .ZN(n6754) );
  AOI22_X1 U7665 ( .A1(n6752), .A2(keyinput_g38), .B1(n6751), .B2(keyinput_g50), .ZN(n6750) );
  OAI221_X1 U7666 ( .B1(n6752), .B2(keyinput_g38), .C1(n6751), .C2(
        keyinput_g50), .A(n6750), .ZN(n6753) );
  NOR4_X1 U7667 ( .A1(n6756), .A2(n6755), .A3(n6754), .A4(n6753), .ZN(n6774)
         );
  AOI22_X1 U7668 ( .A1(n6759), .A2(keyinput_g49), .B1(n6758), .B2(keyinput_g6), 
        .ZN(n6757) );
  OAI221_X1 U7669 ( .B1(n6759), .B2(keyinput_g49), .C1(n6758), .C2(keyinput_g6), .A(n6757), .ZN(n6772) );
  AOI22_X1 U7670 ( .A1(n6762), .A2(keyinput_g42), .B1(keyinput_g40), .B2(n6761), .ZN(n6760) );
  OAI221_X1 U7671 ( .B1(n6762), .B2(keyinput_g42), .C1(n6761), .C2(
        keyinput_g40), .A(n6760), .ZN(n6771) );
  INV_X1 U7672 ( .A(DATAI_23_), .ZN(n6765) );
  AOI22_X1 U7673 ( .A1(n6765), .A2(keyinput_g8), .B1(keyinput_g15), .B2(n6764), 
        .ZN(n6763) );
  OAI221_X1 U7674 ( .B1(n6765), .B2(keyinput_g8), .C1(n6764), .C2(keyinput_g15), .A(n6763), .ZN(n6770) );
  INV_X1 U7675 ( .A(BS16_N), .ZN(n6768) );
  AOI22_X1 U7676 ( .A1(n6768), .A2(keyinput_g34), .B1(n6767), .B2(keyinput_g53), .ZN(n6766) );
  OAI221_X1 U7677 ( .B1(n6768), .B2(keyinput_g34), .C1(n6767), .C2(
        keyinput_g53), .A(n6766), .ZN(n6769) );
  NOR4_X1 U7678 ( .A1(n6772), .A2(n6771), .A3(n6770), .A4(n6769), .ZN(n6773)
         );
  NAND4_X1 U7679 ( .A1(n6776), .A2(n6775), .A3(n6774), .A4(n6773), .ZN(n6815)
         );
  AOI22_X1 U7680 ( .A1(REIP_REG_27__SCAN_IN), .A2(keyinput_g55), .B1(
        REIP_REG_23__SCAN_IN), .B2(keyinput_g59), .ZN(n6777) );
  OAI221_X1 U7681 ( .B1(REIP_REG_27__SCAN_IN), .B2(keyinput_g55), .C1(
        REIP_REG_23__SCAN_IN), .C2(keyinput_g59), .A(n6777), .ZN(n6784) );
  AOI22_X1 U7682 ( .A1(DATAI_22_), .A2(keyinput_g9), .B1(REIP_REG_19__SCAN_IN), 
        .B2(keyinput_g63), .ZN(n6778) );
  OAI221_X1 U7683 ( .B1(DATAI_22_), .B2(keyinput_g9), .C1(REIP_REG_19__SCAN_IN), .C2(keyinput_g63), .A(n6778), .ZN(n6783) );
  AOI22_X1 U7684 ( .A1(DATAI_6_), .A2(keyinput_g25), .B1(DATAI_27_), .B2(
        keyinput_g4), .ZN(n6779) );
  OAI221_X1 U7685 ( .B1(DATAI_6_), .B2(keyinput_g25), .C1(DATAI_27_), .C2(
        keyinput_g4), .A(n6779), .ZN(n6782) );
  AOI22_X1 U7686 ( .A1(DATAI_14_), .A2(keyinput_g17), .B1(REIP_REG_25__SCAN_IN), .B2(keyinput_g57), .ZN(n6780) );
  OAI221_X1 U7687 ( .B1(DATAI_14_), .B2(keyinput_g17), .C1(
        REIP_REG_25__SCAN_IN), .C2(keyinput_g57), .A(n6780), .ZN(n6781) );
  NOR4_X1 U7688 ( .A1(n6784), .A2(n6783), .A3(n6782), .A4(n6781), .ZN(n6813)
         );
  XOR2_X1 U7689 ( .A(n6785), .B(keyinput_g22), .Z(n6793) );
  AOI22_X1 U7690 ( .A1(D_C_N_REG_SCAN_IN), .A2(keyinput_g41), .B1(n6787), .B2(
        keyinput_g31), .ZN(n6786) );
  OAI221_X1 U7691 ( .B1(D_C_N_REG_SCAN_IN), .B2(keyinput_g41), .C1(n6787), 
        .C2(keyinput_g31), .A(n6786), .ZN(n6792) );
  AOI22_X1 U7692 ( .A1(DATAI_21_), .A2(keyinput_g10), .B1(DATAI_12_), .B2(
        keyinput_g19), .ZN(n6788) );
  OAI221_X1 U7693 ( .B1(DATAI_21_), .B2(keyinput_g10), .C1(DATAI_12_), .C2(
        keyinput_g19), .A(n6788), .ZN(n6791) );
  AOI22_X1 U7694 ( .A1(W_R_N_REG_SCAN_IN), .A2(keyinput_g46), .B1(DATAI_30_), 
        .B2(keyinput_g1), .ZN(n6789) );
  OAI221_X1 U7695 ( .B1(W_R_N_REG_SCAN_IN), .B2(keyinput_g46), .C1(DATAI_30_), 
        .C2(keyinput_g1), .A(n6789), .ZN(n6790) );
  NOR4_X1 U7696 ( .A1(n6793), .A2(n6792), .A3(n6791), .A4(n6790), .ZN(n6812)
         );
  AOI22_X1 U7697 ( .A1(DATAI_20_), .A2(keyinput_g11), .B1(REIP_REG_21__SCAN_IN), .B2(keyinput_g61), .ZN(n6794) );
  OAI221_X1 U7698 ( .B1(DATAI_20_), .B2(keyinput_g11), .C1(
        REIP_REG_21__SCAN_IN), .C2(keyinput_g61), .A(n6794), .ZN(n6801) );
  AOI22_X1 U7699 ( .A1(DATAI_26_), .A2(keyinput_g5), .B1(REIP_REG_31__SCAN_IN), 
        .B2(keyinput_g51), .ZN(n6795) );
  OAI221_X1 U7700 ( .B1(DATAI_26_), .B2(keyinput_g5), .C1(REIP_REG_31__SCAN_IN), .C2(keyinput_g51), .A(n6795), .ZN(n6800) );
  AOI22_X1 U7701 ( .A1(DATAI_18_), .A2(keyinput_g13), .B1(DATAI_2_), .B2(
        keyinput_g29), .ZN(n6796) );
  OAI221_X1 U7702 ( .B1(DATAI_18_), .B2(keyinput_g13), .C1(DATAI_2_), .C2(
        keyinput_g29), .A(n6796), .ZN(n6799) );
  AOI22_X1 U7703 ( .A1(MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_g32), .B1(
        REIP_REG_26__SCAN_IN), .B2(keyinput_g56), .ZN(n6797) );
  OAI221_X1 U7704 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_g32), .C1(
        REIP_REG_26__SCAN_IN), .C2(keyinput_g56), .A(n6797), .ZN(n6798) );
  NOR4_X1 U7705 ( .A1(n6801), .A2(n6800), .A3(n6799), .A4(n6798), .ZN(n6811)
         );
  AOI22_X1 U7706 ( .A1(MORE_REG_SCAN_IN), .A2(keyinput_g44), .B1(DATAI_8_), 
        .B2(keyinput_g23), .ZN(n6802) );
  OAI221_X1 U7707 ( .B1(MORE_REG_SCAN_IN), .B2(keyinput_g44), .C1(DATAI_8_), 
        .C2(keyinput_g23), .A(n6802), .ZN(n6809) );
  AOI22_X1 U7708 ( .A1(BYTEENABLE_REG_0__SCAN_IN), .A2(keyinput_g47), .B1(
        REIP_REG_28__SCAN_IN), .B2(keyinput_g54), .ZN(n6803) );
  OAI221_X1 U7709 ( .B1(BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_g47), .C1(
        REIP_REG_28__SCAN_IN), .C2(keyinput_g54), .A(n6803), .ZN(n6808) );
  AOI22_X1 U7710 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(keyinput_g39), .B1(
        DATAI_15_), .B2(keyinput_g16), .ZN(n6804) );
  OAI221_X1 U7711 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(keyinput_g39), .C1(
        DATAI_15_), .C2(keyinput_g16), .A(n6804), .ZN(n6807) );
  AOI22_X1 U7712 ( .A1(DATAI_17_), .A2(keyinput_g14), .B1(DATAI_4_), .B2(
        keyinput_g27), .ZN(n6805) );
  OAI221_X1 U7713 ( .B1(DATAI_17_), .B2(keyinput_g14), .C1(DATAI_4_), .C2(
        keyinput_g27), .A(n6805), .ZN(n6806) );
  NOR4_X1 U7714 ( .A1(n6809), .A2(n6808), .A3(n6807), .A4(n6806), .ZN(n6810)
         );
  NAND4_X1 U7715 ( .A1(n6813), .A2(n6812), .A3(n6811), .A4(n6810), .ZN(n6814)
         );
  OAI22_X1 U7716 ( .A1(keyinput_g24), .A2(n6818), .B1(n6815), .B2(n6814), .ZN(
        n6816) );
  AOI211_X1 U7717 ( .C1(keyinput_g24), .C2(n6818), .A(n6817), .B(n6816), .ZN(
        n6822) );
  AOI22_X1 U7718 ( .A1(n6820), .A2(BYTEENABLE_REG_3__SCAN_IN), .B1(
        BE_N_REG_3__SCAN_IN), .B2(n6819), .ZN(n6821) );
  XNOR2_X1 U7719 ( .A(n6822), .B(n6821), .ZN(U3445) );
  BUF_X1 U3438 ( .A(n3261), .Z(n2989) );
  AOI211_X2 U3433 ( .C1(n4972), .C2(n5875), .A(n4970), .B(n4969), .ZN(n5012)
         );
  CLKBUF_X1 U3450 ( .A(n5342), .Z(n3010) );
  CLKBUF_X1 U34520 ( .A(n3282), .Z(n3004) );
  CLKBUF_X1 U3454 ( .A(n3628), .Z(n3770) );
  CLKBUF_X1 U34720 ( .A(n5532), .Z(n5607) );
  AOI21_X1 U3475 ( .B1(n5681), .B2(n5688), .A(n5680), .ZN(n5682) );
  CLKBUF_X1 U3496 ( .A(n3807), .Z(n3808) );
  CLKBUF_X1 U3816 ( .A(n6242), .Z(n6235) );
  OR2_X1 U3975 ( .A1(n3820), .A2(n4672), .ZN(n6823) );
endmodule

