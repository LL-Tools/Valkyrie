

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9710, n9711, n9712, n9713, n9714, n9715, n9717, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
         n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642,
         n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
         n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658,
         n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666,
         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
         n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
         n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,
         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,
         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,
         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,
         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,
         n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,
         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,
         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,
         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050,
         n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
         n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
         n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074,
         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
         n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090,
         n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
         n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
         n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
         n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,
         n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
         n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,
         n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146,
         n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
         n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162,
         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
         n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,
         n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
         n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234,
         n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,
         n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,
         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
         n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
         n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
         n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,
         n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
         n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306,
         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
         n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
         n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338,
         n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
         n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
         n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,
         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
         n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
         n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
         n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
         n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,
         n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
         n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
         n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
         n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
         n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,
         n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,
         n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,
         n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546,
         n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554,
         n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562,
         n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,
         n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578,
         n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586,
         n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594,
         n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602,
         n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
         n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618,
         n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626,
         n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634,
         n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642,
         n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650,
         n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658,
         n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666,
         n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674,
         n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682,
         n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690,
         n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698,
         n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706,
         n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714,
         n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722,
         n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730,
         n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738,
         n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746,
         n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754,
         n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762,
         n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770,
         n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778,
         n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786,
         n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794,
         n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802,
         n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810,
         n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818,
         n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826,
         n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834,
         n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842,
         n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850,
         n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858,
         n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866,
         n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874,
         n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882,
         n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890,
         n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898,
         n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906,
         n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914,
         n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922,
         n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930,
         n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938,
         n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946,
         n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954,
         n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962,
         n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970,
         n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978,
         n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986,
         n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994,
         n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002,
         n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010,
         n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018,
         n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026,
         n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034,
         n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042,
         n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050,
         n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058,
         n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066,
         n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074,
         n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082,
         n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090,
         n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098,
         n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106,
         n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114,
         n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122,
         n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130,
         n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138,
         n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146,
         n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154,
         n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162,
         n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170,
         n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178,
         n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186,
         n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194,
         n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202,
         n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210,
         n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218,
         n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226,
         n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234,
         n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242,
         n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250,
         n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258,
         n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266,
         n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274,
         n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282,
         n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290,
         n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298,
         n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306,
         n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314,
         n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322,
         n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330,
         n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338,
         n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346,
         n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354,
         n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362,
         n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370,
         n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378,
         n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386,
         n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394,
         n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402,
         n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410,
         n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418,
         n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426,
         n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434,
         n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442,
         n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450,
         n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458,
         n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466,
         n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474,
         n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482,
         n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490,
         n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498,
         n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506,
         n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514,
         n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
         n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530,
         n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538,
         n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546,
         n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554,
         n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562,
         n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570,
         n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578,
         n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586,
         n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594,
         n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602,
         n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610,
         n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618,
         n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626,
         n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634,
         n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642,
         n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650,
         n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658,
         n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666,
         n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674,
         n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682,
         n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690,
         n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698,
         n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706,
         n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714,
         n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722,
         n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730,
         n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738,
         n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746,
         n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754,
         n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762,
         n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770,
         n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778,
         n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786,
         n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794,
         n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802,
         n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810,
         n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818,
         n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826,
         n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834,
         n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842,
         n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850,
         n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858,
         n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866,
         n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874,
         n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882,
         n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890,
         n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898,
         n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906,
         n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914,
         n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922,
         n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930,
         n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938,
         n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946,
         n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954,
         n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962,
         n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970,
         n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978,
         n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986,
         n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994,
         n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002,
         n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010,
         n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018,
         n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026,
         n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034,
         n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042,
         n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050,
         n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058,
         n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066,
         n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074,
         n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082,
         n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090,
         n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098,
         n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106,
         n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114,
         n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122,
         n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130,
         n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138,
         n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146,
         n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154,
         n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162,
         n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170,
         n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178,
         n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186,
         n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194,
         n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202,
         n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210,
         n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218,
         n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226,
         n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234,
         n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242,
         n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250,
         n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258,
         n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266,
         n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274,
         n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282,
         n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290,
         n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298,
         n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306,
         n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314,
         n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322,
         n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330,
         n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338,
         n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346,
         n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354,
         n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362,
         n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370,
         n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378,
         n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386,
         n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394,
         n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402,
         n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410,
         n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418,
         n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426,
         n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434,
         n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442,
         n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450,
         n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458,
         n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466,
         n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474,
         n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482,
         n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490,
         n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498,
         n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506,
         n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514,
         n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522,
         n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530,
         n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538,
         n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546,
         n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554,
         n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18563,
         n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571,
         n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579,
         n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587,
         n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595,
         n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603,
         n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611,
         n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619,
         n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627,
         n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635,
         n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643,
         n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651,
         n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659,
         n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667,
         n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675,
         n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683,
         n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691,
         n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699,
         n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707,
         n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715,
         n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723,
         n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731,
         n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
         n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747,
         n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755,
         n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763,
         n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771,
         n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779,
         n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787,
         n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795,
         n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803,
         n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811,
         n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819,
         n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827,
         n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835,
         n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843,
         n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851,
         n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859,
         n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867,
         n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875,
         n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883,
         n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891,
         n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899,
         n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907,
         n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915,
         n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923,
         n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931,
         n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939,
         n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947,
         n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955,
         n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963,
         n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971,
         n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979,
         n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987,
         n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995,
         n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003,
         n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011,
         n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019,
         n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027,
         n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035,
         n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043,
         n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051,
         n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059,
         n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067,
         n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075,
         n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083,
         n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091,
         n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099,
         n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107,
         n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115,
         n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123,
         n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131,
         n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139,
         n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147,
         n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155,
         n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163,
         n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171,
         n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179,
         n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187,
         n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195,
         n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203,
         n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211,
         n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219,
         n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227,
         n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235,
         n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243,
         n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251,
         n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259,
         n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267,
         n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275,
         n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283,
         n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291,
         n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299,
         n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307,
         n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315,
         n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323,
         n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331,
         n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339,
         n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347,
         n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355,
         n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363,
         n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371,
         n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379,
         n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387,
         n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395,
         n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403,
         n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411,
         n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419,
         n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427,
         n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435,
         n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443,
         n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451,
         n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459,
         n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467,
         n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475,
         n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483,
         n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491,
         n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499,
         n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507,
         n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515,
         n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523,
         n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531,
         n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539,
         n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547,
         n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555,
         n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563,
         n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571,
         n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579,
         n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587,
         n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595,
         n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603,
         n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611,
         n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619,
         n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627,
         n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635,
         n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643,
         n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651,
         n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659,
         n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667,
         n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675,
         n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683,
         n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691,
         n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699,
         n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707,
         n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715,
         n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723,
         n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731,
         n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739,
         n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747,
         n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755,
         n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763,
         n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771,
         n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779,
         n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787,
         n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795,
         n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803,
         n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811,
         n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819,
         n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827,
         n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835,
         n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843,
         n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851,
         n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859,
         n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867,
         n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875,
         n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883,
         n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891,
         n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899,
         n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907,
         n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915,
         n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923,
         n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931,
         n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939,
         n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947,
         n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955,
         n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963,
         n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971,
         n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979,
         n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987,
         n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995,
         n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003,
         n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011,
         n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019,
         n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027,
         n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035,
         n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043,
         n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051,
         n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059,
         n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067,
         n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075,
         n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083,
         n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091,
         n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099,
         n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107,
         n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115,
         n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123,
         n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131,
         n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139,
         n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147,
         n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155,
         n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163,
         n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171,
         n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179,
         n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187,
         n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195,
         n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203,
         n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211,
         n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219,
         n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227,
         n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235,
         n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243,
         n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251,
         n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259,
         n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267,
         n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275,
         n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283,
         n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291,
         n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299,
         n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307,
         n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315,
         n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323,
         n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331,
         n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339,
         n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347,
         n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355,
         n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363,
         n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371,
         n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379,
         n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387,
         n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395,
         n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403,
         n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411,
         n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419,
         n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427,
         n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435,
         n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443,
         n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451,
         n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459,
         n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467,
         n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475,
         n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483,
         n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491,
         n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499,
         n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507,
         n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515,
         n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523,
         n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531,
         n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539,
         n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547,
         n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555,
         n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563,
         n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571,
         n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579,
         n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587,
         n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595,
         n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603,
         n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611,
         n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619,
         n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627,
         n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635,
         n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643,
         n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651,
         n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659,
         n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667,
         n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675,
         n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683,
         n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691,
         n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699,
         n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707,
         n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715,
         n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723,
         n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731,
         n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739,
         n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747,
         n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755,
         n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763,
         n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771,
         n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779,
         n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787,
         n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795,
         n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803,
         n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811,
         n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819,
         n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827,
         n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835,
         n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843,
         n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851,
         n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859,
         n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867,
         n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875,
         n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883,
         n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891,
         n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899,
         n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907,
         n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915,
         n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923,
         n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931,
         n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939,
         n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947,
         n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955,
         n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963,
         n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971,
         n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979,
         n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987,
         n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995,
         n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003,
         n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011,
         n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019,
         n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027,
         n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035,
         n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043,
         n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051,
         n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059,
         n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067,
         n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075,
         n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083,
         n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091,
         n21092, n21093, n21095, n21096, n21097, n21098, n21099, n21100,
         n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108,
         n21109, n21110, n21111, n21112, n21113, n21114, n21115, n21116,
         n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124,
         n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132,
         n21133, n21134, n21135, n21136, n21137, n21138, n21139, n21140,
         n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148,
         n21149, n21150, n21151, n21152, n21153, n21154, n21155, n21156,
         n21157, n21158, n21159, n21160, n21161, n21162, n21163, n21164,
         n21165, n21166, n21167, n21168, n21169, n21170, n21171, n21172,
         n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180,
         n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188,
         n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196,
         n21197, n21198, n21199, n21200, n21201, n21202, n21203, n21204,
         n21205, n21206, n21207, n21208, n21209, n21210, n21211, n21212,
         n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220,
         n21221, n21222, n21223, n21224, n21225, n21226, n21227, n21228,
         n21229, n21230, n21231, n21232, n21233, n21234, n21235, n21236,
         n21237, n21238, n21239, n21240, n21241, n21242, n21243, n21244,
         n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252,
         n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260,
         n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268,
         n21269, n21270, n21271, n21272, n21273, n21274, n21275, n21276,
         n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21284,
         n21285, n21286, n21287, n21288, n21289, n21290, n21291, n21292,
         n21293, n21294, n21295, n21296, n21297, n21298, n21299, n21300,
         n21301, n21302, n21303, n21304, n21305, n21306, n21307, n21308,
         n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316,
         n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324,
         n21325, n21326, n21327, n21328, n21329, n21330, n21331, n21332,
         n21333, n21334, n21335, n21336, n21337, n21338, n21339, n21340,
         n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348,
         n21349, n21350, n21351, n21352, n21353, n21354, n21355, n21356,
         n21357, n21358, n21359, n21360, n21361, n21362, n21363, n21364,
         n21365, n21366, n21367, n21368, n21369, n21370, n21371, n21372,
         n21373, n21374, n21375, n21376, n21377, n21378, n21379, n21380,
         n21381, n21382, n21383, n21384, n21385, n21386, n21387, n21388,
         n21389, n21390, n21391, n21392, n21393, n21394, n21395, n21396,
         n21397, n21398, n21399, n21400, n21401, n21402, n21403, n21404,
         n21405, n21406, n21407, n21408, n21409, n21410, n21411, n21412,
         n21413, n21414, n21415, n21416, n21417, n21418, n21419, n21420,
         n21421, n21422, n21423, n21424, n21425, n21426, n21427, n21428,
         n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21436,
         n21437, n21438, n21439, n21440, n21441, n21442, n21443, n21444,
         n21445, n21446, n21447, n21448, n21449, n21450, n21451, n21452,
         n21453, n21454, n21455, n21456, n21457, n21458, n21459, n21460,
         n21461, n21462, n21463, n21464, n21465, n21466, n21467, n21468,
         n21469, n21470, n21471, n21472, n21473, n21474, n21475, n21476,
         n21477, n21478, n21479, n21480, n21481, n21482, n21483, n21484,
         n21485, n21486, n21487, n21488, n21489, n21490, n21491, n21492,
         n21493, n21494, n21495, n21496, n21497, n21498, n21499, n21500,
         n21501, n21502, n21503, n21504, n21505, n21506, n21507, n21508,
         n21509, n21510, n21511, n21512, n21513, n21514, n21515, n21516,
         n21517, n21518, n21519, n21520, n21521, n21522, n21523, n21524,
         n21525, n21526, n21527, n21528, n21529, n21530, n21531, n21532,
         n21533, n21534, n21535, n21536, n21537, n21538, n21539, n21540,
         n21541, n21542, n21543, n21544, n21545, n21546, n21547, n21548,
         n21549, n21550, n21551, n21552, n21553, n21554, n21555, n21556,
         n21557, n21558, n21559, n21560, n21561, n21562, n21563, n21564,
         n21565, n21566, n21567, n21568, n21569, n21570, n21571, n21572,
         n21573, n21574, n21575, n21576, n21577, n21578, n21579, n21580,
         n21581, n21582, n21583, n21584, n21585, n21586, n21587, n21588,
         n21589, n21590, n21591, n21592, n21593, n21594, n21595, n21596,
         n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604,
         n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612,
         n21613, n21614, n21615, n21616, n21617, n21618, n21619, n21620,
         n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628,
         n21629, n21630, n21631, n21632, n21633, n21634, n21635, n21636,
         n21637, n21638, n21639, n21640, n21641, n21642, n21643, n21644,
         n21645, n21646, n21647, n21648, n21649, n21650, n21651, n21652,
         n21653, n21654, n21655, n21656, n21657, n21658, n21659, n21660,
         n21661, n21662, n21663, n21664, n21665, n21666, n21667, n21668,
         n21669, n21670, n21671, n21672, n21673, n21674, n21675, n21676,
         n21677, n21678, n21679, n21680, n21681, n21682, n21683, n21684,
         n21685, n21686, n21687, n21688, n21689, n21690, n21691, n21692,
         n21693, n21694, n21695, n21696, n21697, n21698, n21699, n21700,
         n21701, n21702, n21703, n21704, n21705, n21706, n21707, n21708,
         n21709, n21710, n21711, n21712, n21713, n21714, n21715, n21716,
         n21717, n21718, n21719, n21720, n21721, n21722, n21723, n21724,
         n21725, n21726, n21727, n21728, n21729, n21730, n21731, n21732,
         n21733, n21734, n21735, n21736, n21737, n21738, n21739, n21740,
         n21741, n21742, n21743, n21744, n21745, n21746, n21747, n21748,
         n21749, n21750, n21751, n21752, n21753, n21754, n21755, n21756,
         n21757, n21758, n21759, n21760, n21761, n21762, n21763, n21764,
         n21765, n21766, n21767, n21768, n21769, n21770, n21771, n21772,
         n21773, n21774, n21775, n21776, n21777, n21778, n21779, n21780,
         n21781, n21782, n21783, n21784, n21785, n21786, n21787, n21788,
         n21789, n21790, n21791, n21792, n21793, n21794, n21795, n21796,
         n21797, n21798, n21799, n21800, n21801, n21802, n21803, n21804,
         n21805, n21806, n21807, n21808, n21809, n21810, n21811, n21812,
         n21813, n21814, n21815, n21816, n21817, n21818, n21819, n21820,
         n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828,
         n21829, n21830, n21831, n21832, n21833, n21834, n21835, n21836,
         n21837, n21838, n21839, n21840, n21841, n21842, n21843, n21844,
         n21845, n21846, n21847, n21848, n21849, n21850, n21851, n21852,
         n21853, n21854, n21855, n21856, n21857, n21858, n21859, n21860,
         n21861, n21862, n21863, n21864, n21865, n21866, n21867, n21868,
         n21869, n21870, n21871, n21872, n21873, n21874, n21875, n21876,
         n21877, n21878, n21879, n21880, n21881, n21882, n21883, n21884,
         n21885, n21886, n21887, n21888, n21889, n21890, n21891, n21892,
         n21893, n21894, n21895, n21896, n21897, n21898, n21899, n21900,
         n21901, n21902, n21903, n21904, n21905, n21906, n21907, n21908,
         n21909, n21910, n21911, n21912, n21913, n21914, n21915, n21916,
         n21917, n21918, n21919, n21920, n21921, n21922, n21923, n21924,
         n21925, n21926, n21927, n21928, n21929, n21930, n21931, n21932,
         n21933, n21934, n21935, n21936, n21937, n21938, n21939, n21940,
         n21941, n21942, n21943, n21944, n21945, n21946, n21947, n21948,
         n21949, n21950, n21951, n21952, n21953, n21954, n21955, n21956,
         n21957, n21958, n21959, n21960, n21961, n21962, n21963, n21964,
         n21965, n21966, n21967, n21968, n21969, n21970, n21971, n21972,
         n21973, n21974, n21975, n21976, n21977, n21978, n21979, n21980,
         n21981, n21982, n21983, n21984, n21985, n21986, n21987, n21988,
         n21989, n21990, n21991, n21992, n21993, n21994, n21995, n21996,
         n21997, n21998, n21999, n22000, n22001, n22002, n22003, n22004,
         n22005, n22006, n22007, n22008, n22009, n22010, n22011, n22012,
         n22013, n22014, n22015, n22016, n22017, n22018, n22019, n22020,
         n22021, n22022, n22023, n22024, n22025, n22026, n22027, n22028,
         n22029, n22030, n22031, n22032, n22033, n22034, n22035, n22036,
         n22037, n22038, n22039, n22040, n22041, n22042, n22043, n22044,
         n22045, n22046, n22047, n22048, n22049, n22050, n22051, n22052,
         n22053, n22054, n22055, n22056, n22057, n22058, n22059, n22060,
         n22061, n22062, n22063, n22064, n22065, n22066, n22067, n22068,
         n22069, n22070, n22071, n22072, n22073, n22074, n22075, n22076,
         n22077, n22078, n22079, n22080, n22081, n22082, n22083, n22084,
         n22085, n22086, n22087, n22088, n22089, n22090, n22091, n22092,
         n22093, n22094, n22095, n22096, n22097, n22098, n22099, n22100,
         n22101, n22102, n22103, n22104, n22105, n22106, n22107, n22108,
         n22109, n22110, n22111, n22112, n22113, n22114, n22115, n22116,
         n22117, n22118, n22119, n22120, n22121, n22122, n22123, n22124,
         n22125, n22126, n22127, n22128, n22129, n22130, n22131, n22132,
         n22133, n22134, n22135, n22136, n22137, n22138, n22139, n22140,
         n22141, n22142, n22143, n22144, n22145, n22146, n22147, n22148,
         n22149;

  INV_X2 U11142 ( .A(n21095), .ZN(n20976) );
  OAI21_X1 U11143 ( .B1(n20688), .B2(n20687), .A(n20686), .ZN(n20704) );
  NOR2_X1 U11144 ( .A1(n20682), .A2(n10370), .ZN(n20683) );
  NOR2_X1 U11145 ( .A1(n20722), .A2(n20721), .ZN(n20755) );
  OR3_X1 U11146 ( .A1(n17992), .A2(n21099), .A3(n18011), .ZN(n21105) );
  AND2_X1 U11147 ( .A1(n11240), .A2(n10050), .ZN(n15391) );
  INV_X2 U11148 ( .A(n20708), .ZN(n20679) );
  NAND2_X1 U11150 ( .A1(n20094), .A2(n20212), .ZN(n18244) );
  NAND2_X1 U11151 ( .A1(n13934), .A2(n13933), .ZN(n20094) );
  XNOR2_X1 U11152 ( .A(n12422), .B(n12423), .ZN(n17234) );
  NAND2_X1 U11153 ( .A1(n14451), .A2(n14522), .ZN(n14521) );
  NAND2_X1 U11154 ( .A1(n10617), .A2(n9991), .ZN(n20757) );
  OR2_X2 U11155 ( .A1(n14219), .A2(n17778), .ZN(n19196) );
  CLKBUF_X1 U11156 ( .A(n10871), .Z(n11434) );
  NAND4_X1 U11157 ( .A1(n12045), .A2(n12044), .A3(n12043), .A4(n12042), .ZN(
        n18917) );
  CLKBUF_X2 U11158 ( .A(n12919), .Z(n13126) );
  CLKBUF_X2 U11160 ( .A(n10756), .Z(n11478) );
  INV_X1 U11161 ( .A(n10877), .ZN(n10893) );
  INV_X1 U11162 ( .A(n18773), .ZN(n18742) );
  CLKBUF_X2 U11163 ( .A(n10775), .Z(n11269) );
  AOI21_X1 U11164 ( .B1(n14713), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10076), 
        .ZN(n10075) );
  NAND2_X1 U11165 ( .A1(n11877), .A2(n10675), .ZN(n11875) );
  CLKBUF_X2 U11166 ( .A(n12901), .Z(n13145) );
  NAND2_X1 U11167 ( .A1(n14189), .A2(n14188), .ZN(n14198) );
  INV_X1 U11168 ( .A(n15177), .ZN(n15145) );
  AND2_X1 U11171 ( .A1(n12577), .A2(n13824), .ZN(n15173) );
  INV_X1 U11172 ( .A(n14112), .ZN(n17695) );
  NAND2_X2 U11173 ( .A1(n14026), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n18775) );
  INV_X4 U11174 ( .A(n9890), .ZN(n9712) );
  AND2_X2 U11175 ( .A1(n10699), .A2(n14351), .ZN(n10943) );
  AND2_X2 U11176 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14351) );
  CLKBUF_X1 U11177 ( .A(n14583), .Z(n9698) );
  NOR2_X1 U11178 ( .A1(n18057), .A2(n14547), .ZN(n14583) );
  OR2_X1 U11179 ( .A1(n21270), .A2(n14561), .ZN(n21271) );
  INV_X1 U11180 ( .A(n21271), .ZN(n9699) );
  INV_X1 U11181 ( .A(n18086), .ZN(n9700) );
  NAND2_X1 U11183 ( .A1(n17093), .A2(n17365), .ZN(n17113) );
  AND2_X4 U11184 ( .A1(n13670), .A2(n13671), .ZN(n17966) );
  INV_X2 U11185 ( .A(n18917), .ZN(n19628) );
  AOI21_X1 U11186 ( .B1(n11716), .B2(n10978), .A(n10913), .ZN(n9702) );
  AOI21_X1 U11187 ( .B1(n11716), .B2(n10978), .A(n10913), .ZN(n10968) );
  NOR2_X2 U11188 ( .A1(n11870), .A2(n19031), .ZN(n11869) );
  NAND2_X1 U11189 ( .A1(n12585), .A2(n9809), .ZN(n10115) );
  AND2_X1 U11190 ( .A1(n10706), .A2(n10705), .ZN(n11111) );
  AND2_X1 U11191 ( .A1(n10574), .A2(n9861), .ZN(n11716) );
  XNOR2_X1 U11192 ( .A(n12798), .B(n12261), .ZN(n12262) );
  INV_X1 U11193 ( .A(n13862), .ZN(n18624) );
  NOR2_X1 U11194 ( .A1(n14879), .A2(n15593), .ZN(n15594) );
  AND2_X2 U11195 ( .A1(n12724), .A2(n12630), .ZN(n12731) );
  OR2_X1 U11196 ( .A1(n12629), .A2(n12692), .ZN(n12696) );
  INV_X1 U11198 ( .A(n12879), .ZN(n13220) );
  OR2_X1 U11199 ( .A1(n10551), .A2(n10283), .ZN(n10282) );
  NAND2_X1 U11200 ( .A1(n10617), .A2(n9962), .ZN(n17579) );
  INV_X2 U11201 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12129) );
  INV_X1 U11202 ( .A(n18715), .ZN(n10682) );
  CLKBUF_X3 U11203 ( .A(n9711), .Z(n9706) );
  AND2_X1 U11204 ( .A1(n19303), .A2(n10320), .ZN(n10319) );
  INV_X1 U11205 ( .A(n9724), .ZN(n13570) );
  CLKBUF_X3 U11206 ( .A(n15028), .Z(n9703) );
  AND2_X1 U11207 ( .A1(n15526), .A2(n10545), .ZN(n15481) );
  AND2_X2 U11208 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13805) );
  INV_X1 U11210 ( .A(n12901), .ZN(n12551) );
  NAND2_X1 U11211 ( .A1(n20713), .A2(n21079), .ZN(n20619) );
  INV_X1 U11212 ( .A(n19560), .ZN(n20058) );
  OAI211_X1 U11213 ( .C1(n14201), .C2(n10321), .A(n10319), .B(1'b1), .ZN(
        n19302) );
  INV_X1 U11214 ( .A(n19236), .ZN(n19183) );
  INV_X1 U11215 ( .A(n19604), .ZN(n19410) );
  INV_X1 U11216 ( .A(n13690), .ZN(n19634) );
  INV_X1 U11217 ( .A(n21203), .ZN(n21190) );
  INV_X1 U11218 ( .A(n21205), .ZN(n21173) );
  INV_X1 U11219 ( .A(n15781), .ZN(n13423) );
  OR2_X1 U11220 ( .A1(n15453), .A2(n15454), .ZN(n10662) );
  NOR2_X1 U11224 ( .A1(n20753), .A2(n20752), .ZN(n20779) );
  INV_X1 U11225 ( .A(n19654), .ZN(n18606) );
  INV_X1 U11226 ( .A(n18973), .ZN(n20217) );
  CLKBUF_X3 U11227 ( .A(n21217), .Z(n9710) );
  INV_X1 U11228 ( .A(n21047), .ZN(n20713) );
  AOI211_X2 U11229 ( .C1(n17565), .C2(n17564), .A(n20623), .B(n17563), .ZN(
        n20459) );
  AND2_X2 U11230 ( .A1(n12312), .A2(n21964), .ZN(n9736) );
  AND2_X2 U11231 ( .A1(n12312), .A2(n21964), .ZN(n9728) );
  AND2_X4 U11232 ( .A1(n9717), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12379) );
  AND2_X2 U11233 ( .A1(n14708), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9720) );
  AND2_X2 U11234 ( .A1(n14708), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9719) );
  OAI21_X2 U11235 ( .B1(n10385), .B2(n10242), .A(n9788), .ZN(n17220) );
  NOR2_X2 U11236 ( .A1(n12674), .A2(n10506), .ZN(n10505) );
  AOI21_X2 U11237 ( .B1(n10185), .B2(n9749), .A(n9828), .ZN(n10183) );
  BUF_X1 U11238 ( .A(n12797), .Z(n14439) );
  NAND2_X2 U11239 ( .A1(n12731), .A2(n10512), .ZN(n12745) );
  AND2_X1 U11240 ( .A1(n14553), .A2(n14561), .ZN(n15028) );
  AND2_X4 U11241 ( .A1(n14684), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9730) );
  AND2_X2 U11242 ( .A1(n14684), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9729) );
  INV_X2 U11243 ( .A(n12202), .ZN(n9940) );
  AND2_X2 U11245 ( .A1(n12901), .A2(n10104), .ZN(n12220) );
  OR2_X2 U11247 ( .A1(n10726), .A2(n10725), .ZN(n10799) );
  NOR2_X4 U11248 ( .A1(n13263), .A2(n18113), .ZN(n13260) );
  NAND2_X2 U11249 ( .A1(n13264), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13263) );
  NOR2_X2 U11250 ( .A1(n10662), .A2(n15444), .ZN(n15428) );
  AND3_X1 U11251 ( .A1(n12239), .A2(n12238), .A3(n12237), .ZN(n12240) );
  AND2_X4 U11252 ( .A1(n14684), .A2(n21964), .ZN(n9721) );
  OR2_X2 U11253 ( .A1(n10755), .A2(n10754), .ZN(n14553) );
  BUF_X4 U11254 ( .A(n12213), .Z(n14870) );
  INV_X2 U11255 ( .A(n12213), .ZN(n9941) );
  XNOR2_X2 U11256 ( .A(n9778), .B(n12793), .ZN(n12794) );
  OR2_X2 U11257 ( .A1(n12783), .A2(n12777), .ZN(n9778) );
  NOR2_X2 U11258 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12313) );
  NOR2_X4 U11259 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10699) );
  NOR2_X2 U11260 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n18437), .ZN(n18419) );
  CLKBUF_X1 U11261 ( .A(n9890), .Z(n9704) );
  NAND2_X1 U11262 ( .A1(n11897), .A2(n13787), .ZN(n9890) );
  BUF_X4 U11263 ( .A(n9711), .Z(n9705) );
  INV_X2 U11264 ( .A(n18755), .ZN(n9711) );
  XNOR2_X1 U11265 ( .A(n10980), .B(n10979), .ZN(n14384) );
  NAND2_X2 U11266 ( .A1(n12120), .A2(n14685), .ZN(n15259) );
  AOI21_X2 U11267 ( .B1(n15215), .B2(n15214), .A(n9877), .ZN(n15235) );
  NAND2_X2 U11268 ( .A1(n9949), .A2(n9948), .ZN(n12600) );
  BUF_X8 U11269 ( .A(n12177), .Z(n9727) );
  NOR2_X1 U11270 ( .A1(n20721), .A2(n20619), .ZN(n20486) );
  AND2_X4 U11271 ( .A1(n10705), .A2(n10170), .ZN(n10889) );
  AND2_X2 U11272 ( .A1(n10144), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10705) );
  XNOR2_X2 U11273 ( .A(n10970), .B(n14389), .ZN(n10047) );
  AOI21_X2 U11275 ( .B1(n10610), .B2(n17193), .A(n9796), .ZN(n10551) );
  NOR2_X2 U11276 ( .A1(n10365), .A2(n12589), .ZN(n10364) );
  NOR2_X2 U11277 ( .A1(n19146), .A2(n18360), .ZN(n18359) );
  AOI211_X2 U11278 ( .C1(n19593), .C2(n19453), .A(n17937), .B(n19451), .ZN(
        n19414) );
  OAI21_X2 U11279 ( .B1(n20703), .B2(n20683), .A(n20896), .ZN(n20705) );
  NOR2_X2 U11280 ( .A1(n15380), .A2(n15382), .ZN(n15381) );
  NAND2_X1 U11281 ( .A1(n15391), .A2(n15392), .ZN(n15380) );
  NAND2_X1 U11282 ( .A1(n17234), .A2(n22037), .ZN(n9984) );
  AOI21_X1 U11283 ( .B1(n10570), .B2(n15909), .A(n9750), .ZN(n10566) );
  OR2_X1 U11284 ( .A1(n19575), .A2(n19422), .ZN(n19478) );
  AND2_X1 U11285 ( .A1(n14619), .A2(n9856), .ZN(n16573) );
  AND2_X1 U11286 ( .A1(n17873), .A2(n17891), .ZN(n19117) );
  NOR2_X2 U11287 ( .A1(n20753), .A2(n20721), .ZN(n20744) );
  INV_X1 U11288 ( .A(n12690), .ZN(n10169) );
  NAND2_X1 U11289 ( .A1(n21047), .A2(n21079), .ZN(n20753) );
  NAND2_X1 U11290 ( .A1(n10346), .A2(n12318), .ZN(n10211) );
  NAND2_X1 U11291 ( .A1(n21047), .A2(n14849), .ZN(n20722) );
  AOI21_X1 U11292 ( .B1(n16003), .B2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n10669), .ZN(n11760) );
  NOR2_X1 U11293 ( .A1(n21047), .A2(n21079), .ZN(n20656) );
  INV_X4 U11294 ( .A(n20350), .ZN(n10160) );
  INV_X2 U11295 ( .A(n9784), .ZN(n15979) );
  AND2_X1 U11296 ( .A1(n11748), .A2(n11747), .ZN(n9784) );
  INV_X1 U11297 ( .A(n12770), .ZN(n12637) );
  AND2_X1 U11298 ( .A1(n14013), .A2(n16186), .ZN(n16252) );
  NAND2_X1 U11299 ( .A1(n9991), .A2(n9990), .ZN(n12429) );
  NAND3_X2 U11300 ( .A1(n9913), .A2(n9944), .A3(n9946), .ZN(n14287) );
  NAND3_X1 U11301 ( .A1(n12797), .A2(n12800), .A3(n10336), .ZN(n9913) );
  NAND2_X1 U11302 ( .A1(n10829), .A2(n10828), .ZN(n10859) );
  NAND2_X1 U11303 ( .A1(n9956), .A2(n12263), .ZN(n12797) );
  NAND2_X1 U11304 ( .A1(n14541), .A2(n10858), .ZN(n16373) );
  AND2_X1 U11305 ( .A1(n12731), .A2(n9805), .ZN(n12734) );
  XNOR2_X1 U11306 ( .A(n14183), .B(n10304), .ZN(n19280) );
  NAND2_X2 U11307 ( .A1(n19438), .A2(n19410), .ZN(n19477) );
  NAND2_X1 U11308 ( .A1(n12214), .A2(n10075), .ZN(n9961) );
  AOI21_X1 U11309 ( .B1(n19569), .B2(n19297), .A(n14180), .ZN(n19290) );
  OR2_X1 U11311 ( .A1(n12629), .A2(n12631), .ZN(n12726) );
  INV_X1 U11312 ( .A(n13136), .ZN(n9926) );
  NOR2_X1 U11313 ( .A1(n14064), .A2(n13562), .ZN(n13420) );
  NOR2_X1 U11314 ( .A1(n13691), .A2(n12069), .ZN(n12086) );
  AND3_X1 U11315 ( .A1(n10344), .A2(n12217), .A3(n12216), .ZN(n9957) );
  NAND2_X1 U11316 ( .A1(n11650), .A2(n9714), .ZN(n11607) );
  AND2_X1 U11317 ( .A1(n12211), .A2(n20433), .ZN(n14420) );
  AND2_X1 U11318 ( .A1(n12206), .A2(n14870), .ZN(n16419) );
  INV_X1 U11319 ( .A(n13685), .ZN(n19650) );
  NAND2_X1 U11320 ( .A1(n9715), .A2(n12898), .ZN(n12900) );
  AND2_X1 U11321 ( .A1(n12210), .A2(n12215), .ZN(n10591) );
  BUF_X2 U11322 ( .A(n11581), .Z(n9734) );
  NAND2_X1 U11323 ( .A1(n10126), .A2(n10130), .ZN(n13148) );
  NAND2_X1 U11325 ( .A1(n12189), .A2(n12188), .ZN(n12206) );
  BUF_X1 U11326 ( .A(n10769), .Z(n14557) );
  NAND2_X1 U11327 ( .A1(n10685), .A2(n10688), .ZN(n14567) );
  INV_X4 U11328 ( .A(n13659), .ZN(n18613) );
  CLKBUF_X3 U11329 ( .A(n9719), .Z(n9717) );
  CLKBUF_X2 U11330 ( .A(n14099), .Z(n14896) );
  BUF_X2 U11331 ( .A(n10845), .Z(n11335) );
  AOI22_X1 U11332 ( .A1(n9728), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(n9726), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12167) );
  BUF_X2 U11333 ( .A(n10741), .Z(n11412) );
  CLKBUF_X2 U11334 ( .A(n11111), .Z(n11304) );
  CLKBUF_X2 U11335 ( .A(n10727), .Z(n11413) );
  AND2_X2 U11336 ( .A1(n14708), .A2(n21964), .ZN(n15157) );
  AND2_X2 U11337 ( .A1(n14708), .A2(n21964), .ZN(n9732) );
  CLKBUF_X1 U11338 ( .A(n9721), .Z(n15158) );
  AND2_X2 U11339 ( .A1(n10170), .A2(n10699), .ZN(n10775) );
  CLKBUF_X2 U11340 ( .A(n10938), .Z(n11324) );
  AND2_X2 U11342 ( .A1(n12312), .A2(n15153), .ZN(n12371) );
  AND2_X1 U11343 ( .A1(n10830), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10707) );
  AND3_X2 U11344 ( .A1(n13824), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12177) );
  INV_X1 U11345 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13824) );
  NOR3_X2 U11346 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n18580) );
  NOR2_X1 U11347 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12120) );
  AND2_X1 U11348 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13261) );
  OAI21_X1 U11349 ( .B1(n10615), .B2(n10253), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10252) );
  AND2_X1 U11350 ( .A1(n13409), .A2(n18118), .ZN(n13410) );
  NAND2_X1 U11351 ( .A1(n9975), .A2(n9811), .ZN(n10615) );
  AOI211_X1 U11352 ( .C1(n17297), .C2(n18126), .A(n17296), .B(n17295), .ZN(
        n17298) );
  AOI211_X1 U11353 ( .C1(n17337), .C2(n18108), .A(n17064), .B(n17063), .ZN(
        n17065) );
  AOI21_X1 U11354 ( .B1(n10436), .B2(n9814), .A(n10433), .ZN(n17074) );
  AOI21_X1 U11355 ( .B1(n15357), .B2(n18105), .A(n10105), .ZN(n10684) );
  XNOR2_X1 U11356 ( .A(n10106), .B(n12795), .ZN(n15357) );
  AND2_X1 U11357 ( .A1(n17011), .A2(n10001), .ZN(n17297) );
  OAI22_X1 U11358 ( .A1(n10378), .A2(n10377), .B1(n10381), .B2(n10382), .ZN(
        n10376) );
  AOI21_X1 U11359 ( .B1(n10043), .B2(n17431), .A(n17158), .ZN(n17424) );
  AOI21_X1 U11360 ( .B1(n17328), .B2(n17094), .A(n17079), .ZN(n17359) );
  NAND2_X1 U11361 ( .A1(n17118), .A2(n17380), .ZN(n9994) );
  AND2_X1 U11362 ( .A1(n17000), .A2(n10343), .ZN(n17286) );
  NOR2_X1 U11363 ( .A1(n13193), .A2(n10679), .ZN(n16986) );
  NOR2_X1 U11364 ( .A1(n17011), .A2(n9973), .ZN(n17001) );
  NOR2_X1 U11365 ( .A1(n17011), .A2(n9739), .ZN(n13193) );
  AND2_X1 U11366 ( .A1(n17364), .A2(n9770), .ZN(n17079) );
  AND2_X1 U11367 ( .A1(n11866), .A2(n11865), .ZN(n10362) );
  NAND2_X1 U11368 ( .A1(n10339), .A2(n9903), .ZN(n16992) );
  NAND2_X1 U11369 ( .A1(n10391), .A2(n13353), .ZN(n17078) );
  NAND2_X1 U11370 ( .A1(n10397), .A2(n10395), .ZN(n10391) );
  AOI211_X1 U11371 ( .C1(n20362), .C2(BUF2_REG_30__SCAN_IN), .A(n15345), .B(
        n15344), .ZN(n15346) );
  NOR2_X1 U11372 ( .A1(n13341), .A2(n13340), .ZN(n13342) );
  NOR2_X1 U11373 ( .A1(n10496), .A2(n10493), .ZN(n10492) );
  AOI21_X1 U11374 ( .B1(n13425), .B2(n18052), .A(n11690), .ZN(n10565) );
  AOI21_X1 U11375 ( .B1(n17027), .B2(n10372), .A(n10064), .ZN(n13199) );
  XNOR2_X1 U11376 ( .A(n11500), .B(n11499), .ZN(n13425) );
  NAND2_X1 U11377 ( .A1(n10247), .A2(n10248), .ZN(n17098) );
  NAND2_X1 U11378 ( .A1(n10247), .A2(n10245), .ZN(n10397) );
  NAND2_X1 U11379 ( .A1(n10598), .A2(n13344), .ZN(n17156) );
  NAND2_X1 U11380 ( .A1(n10171), .A2(n10566), .ZN(n15857) );
  AOI21_X1 U11381 ( .B1(n15382), .B2(n15380), .A(n15381), .ZN(n15802) );
  NAND2_X1 U11382 ( .A1(n17106), .A2(n10600), .ZN(n10247) );
  NAND2_X1 U11383 ( .A1(n10142), .A2(n10296), .ZN(n15836) );
  AND2_X1 U11384 ( .A1(n9979), .A2(n9978), .ZN(n17020) );
  NAND2_X1 U11385 ( .A1(n10021), .A2(n10022), .ZN(n17204) );
  NAND2_X1 U11386 ( .A1(n10184), .A2(n10183), .ZN(n17040) );
  NAND2_X1 U11387 ( .A1(n10023), .A2(n12514), .ZN(n10022) );
  AND2_X1 U11388 ( .A1(n11240), .A2(n10051), .ZN(n15442) );
  OR2_X1 U11389 ( .A1(n16764), .A2(n16763), .ZN(n10637) );
  NAND2_X1 U11390 ( .A1(n15256), .A2(n10672), .ZN(n10664) );
  XNOR2_X1 U11391 ( .A(n10527), .B(n13224), .ZN(n15359) );
  NAND2_X1 U11392 ( .A1(n17178), .A2(n17180), .ZN(n10185) );
  NAND2_X1 U11393 ( .A1(n12684), .A2(n12683), .ZN(n17490) );
  NAND2_X1 U11394 ( .A1(n12691), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17178) );
  AOI21_X1 U11395 ( .B1(n10298), .B2(n10566), .A(n10297), .ZN(n10299) );
  XNOR2_X1 U11396 ( .A(n12691), .B(n17494), .ZN(n17489) );
  AOI21_X1 U11397 ( .B1(n10372), .B2(n10113), .A(n10112), .ZN(n10111) );
  AND2_X1 U11398 ( .A1(n17225), .A2(n12514), .ZN(n9988) );
  NAND3_X1 U11399 ( .A1(n9974), .A2(n10276), .A3(n10369), .ZN(n12691) );
  XNOR2_X1 U11400 ( .A(n12542), .B(n12627), .ZN(n17206) );
  NAND3_X1 U11401 ( .A1(n10235), .A2(n10234), .A3(n12679), .ZN(n17219) );
  XNOR2_X1 U11402 ( .A(n11656), .B(n11655), .ZN(n11797) );
  NAND2_X1 U11403 ( .A1(n12507), .A2(n12506), .ZN(n17223) );
  AOI211_X2 U11404 ( .C1(n19526), .C2(n19424), .A(n19478), .B(n19423), .ZN(
        n19437) );
  XNOR2_X1 U11405 ( .A(n9989), .B(n12685), .ZN(n12514) );
  AND2_X1 U11406 ( .A1(n13202), .A2(n10678), .ZN(n12784) );
  NOR2_X1 U11407 ( .A1(n16443), .A2(n16990), .ZN(n16434) );
  NAND2_X1 U11408 ( .A1(n9915), .A2(n10550), .ZN(n12542) );
  NOR3_X1 U11409 ( .A1(n20744), .A2(n20717), .A3(n20679), .ZN(n20681) );
  NAND2_X1 U11410 ( .A1(n12682), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17225) );
  OR2_X1 U11411 ( .A1(n12791), .A2(n13197), .ZN(n13203) );
  NAND2_X1 U11412 ( .A1(n10291), .A2(n10289), .ZN(n15906) );
  AND2_X1 U11413 ( .A1(n16535), .A2(n10037), .ZN(n16453) );
  AND2_X1 U11414 ( .A1(n12650), .A2(n9838), .ZN(n10372) );
  INV_X1 U11415 ( .A(n19117), .ZN(n19187) );
  INV_X1 U11416 ( .A(n10277), .ZN(n10550) );
  NOR2_X1 U11417 ( .A1(n10277), .A2(n12690), .ZN(n9989) );
  NAND2_X1 U11418 ( .A1(n20656), .A2(n20893), .ZN(n20708) );
  AND2_X1 U11419 ( .A1(n10571), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10570) );
  AND2_X1 U11420 ( .A1(n20656), .A2(n21043), .ZN(n21836) );
  NOR2_X1 U11421 ( .A1(n10999), .A2(n14447), .ZN(n14513) );
  INV_X1 U11422 ( .A(n10212), .ZN(n10210) );
  INV_X1 U11423 ( .A(n10211), .ZN(n10208) );
  NAND2_X1 U11424 ( .A1(n20656), .A2(n20835), .ZN(n20644) );
  NAND2_X2 U11425 ( .A1(n10399), .A2(n10334), .ZN(n10277) );
  AND2_X1 U11426 ( .A1(n10169), .A2(n12515), .ZN(n9915) );
  OR2_X1 U11427 ( .A1(n10572), .A2(n15909), .ZN(n10571) );
  NOR2_X1 U11428 ( .A1(n11766), .A2(n9810), .ZN(n10292) );
  INV_X1 U11429 ( .A(n14617), .ZN(n14618) );
  AND2_X1 U11430 ( .A1(n10402), .A2(n12393), .ZN(n10212) );
  AND2_X1 U11431 ( .A1(n10402), .A2(n9886), .ZN(n10399) );
  OAI21_X1 U11432 ( .B1(n12787), .B2(n12627), .A(n17266), .ZN(n17008) );
  XNOR2_X1 U11433 ( .A(n12641), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16996) );
  NAND2_X1 U11434 ( .A1(n16000), .A2(n11761), .ZN(n10358) );
  AND2_X1 U11435 ( .A1(n12988), .A2(n9857), .ZN(n14617) );
  OAI21_X1 U11436 ( .B1(n11699), .B2(n11082), .A(n10956), .ZN(n14512) );
  AND2_X1 U11437 ( .A1(n15897), .A2(n10573), .ZN(n10572) );
  OR2_X1 U11438 ( .A1(n16485), .A2(n12627), .ZN(n17018) );
  INV_X1 U11439 ( .A(n14646), .ZN(n10036) );
  NAND2_X1 U11440 ( .A1(n14333), .A2(n10638), .ZN(n15063) );
  OAI21_X1 U11441 ( .B1(n11694), .B2(n11820), .A(n11693), .ZN(n11736) );
  NAND2_X1 U11442 ( .A1(n12471), .A2(n12470), .ZN(n12690) );
  OR2_X1 U11443 ( .A1(n11745), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n18050) );
  AND2_X1 U11444 ( .A1(n18044), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10669) );
  INV_X1 U11445 ( .A(n14625), .ZN(n12988) );
  OR2_X1 U11446 ( .A1(n14392), .A2(n11820), .ZN(n11704) );
  OR2_X1 U11447 ( .A1(n15979), .A2(n22124), .ZN(n15931) );
  OR2_X1 U11448 ( .A1(n15979), .A2(n11840), .ZN(n15939) );
  NAND2_X1 U11449 ( .A1(n11759), .A2(n11758), .ZN(n18044) );
  NAND2_X1 U11450 ( .A1(n15993), .A2(n11753), .ZN(n16003) );
  OR2_X1 U11451 ( .A1(n14285), .A2(n9855), .ZN(n14286) );
  INV_X2 U11452 ( .A(n9784), .ZN(n15993) );
  AND2_X1 U11453 ( .A1(n21058), .A2(n21045), .ZN(n20714) );
  OR2_X1 U11454 ( .A1(n14283), .A2(n14284), .ZN(n10641) );
  OAI22_X1 U11455 ( .A1(n12276), .A2(n20580), .B1(n17579), .B2(n20876), .ZN(
        n12277) );
  NAND2_X1 U11456 ( .A1(n11032), .A2(n11024), .ZN(n11738) );
  OR2_X2 U11457 ( .A1(n19342), .A2(n17942), .ZN(n19208) );
  INV_X1 U11458 ( .A(n10957), .ZN(n10935) );
  NAND2_X1 U11459 ( .A1(n13998), .A2(n14282), .ZN(n14283) );
  NOR2_X2 U11460 ( .A1(n14596), .A2(n15020), .ZN(n13436) );
  OR2_X1 U11461 ( .A1(n16529), .A2(n12627), .ZN(n12747) );
  OR2_X1 U11462 ( .A1(n20646), .A2(n12302), .ZN(n10121) );
  NAND2_X1 U11463 ( .A1(n10168), .A2(n10617), .ZN(n20494) );
  NAND2_X1 U11464 ( .A1(n10168), .A2(n9802), .ZN(n20526) );
  NAND2_X1 U11465 ( .A1(n9992), .A2(n9962), .ZN(n14853) );
  NAND2_X1 U11466 ( .A1(n10168), .A2(n9990), .ZN(n20460) );
  NAND2_X2 U11467 ( .A1(n14591), .A2(n15709), .ZN(n15702) );
  NAND2_X2 U11468 ( .A1(n15709), .A2(n14069), .ZN(n15704) );
  CLKBUF_X1 U11469 ( .A(n10969), .Z(n14389) );
  OR2_X1 U11470 ( .A1(n13997), .A2(n13996), .ZN(n13998) );
  NAND2_X1 U11471 ( .A1(n13997), .A2(n13996), .ZN(n14282) );
  NAND2_X1 U11472 ( .A1(n14004), .A2(n14003), .ZN(n14284) );
  NAND2_X1 U11473 ( .A1(n9962), .A2(n9802), .ZN(n12438) );
  INV_X1 U11474 ( .A(n14287), .ZN(n10123) );
  XNOR2_X1 U11475 ( .A(n14000), .B(n13999), .ZN(n21072) );
  NAND2_X1 U11476 ( .A1(n13164), .A2(n12892), .ZN(n17518) );
  NOR2_X2 U11477 ( .A1(n14704), .A2(n14287), .ZN(n10168) );
  XNOR2_X1 U11478 ( .A(n17539), .B(n14001), .ZN(n14000) );
  NAND2_X1 U11479 ( .A1(n13826), .A2(n13825), .ZN(n17539) );
  BUF_X2 U11480 ( .A(n12274), .Z(n14704) );
  XNOR2_X1 U11481 ( .A(n10912), .B(n10910), .ZN(n10978) );
  INV_X2 U11482 ( .A(n16835), .ZN(n9713) );
  NAND2_X1 U11483 ( .A1(n10905), .A2(n10904), .ZN(n10912) );
  NAND2_X1 U11484 ( .A1(n19280), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n19279) );
  OR2_X1 U11485 ( .A1(n16718), .A2(n13822), .ZN(n12291) );
  XNOR2_X1 U11486 ( .A(n10987), .B(n10986), .ZN(n14752) );
  NAND2_X1 U11487 ( .A1(n12252), .A2(n9947), .ZN(n12800) );
  CLKBUF_X1 U11488 ( .A(n10857), .Z(n14541) );
  OAI22_X1 U11489 ( .A1(n10989), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n10900), 
        .B2(n10921), .ZN(n10987) );
  NAND2_X1 U11490 ( .A1(n12719), .A2(n12726), .ZN(n12724) );
  INV_X2 U11491 ( .A(n20432), .ZN(n13533) );
  NAND2_X1 U11492 ( .A1(n10815), .A2(n10814), .ZN(n10989) );
  NAND2_X1 U11493 ( .A1(n12247), .A2(n12246), .ZN(n12253) );
  INV_X1 U11494 ( .A(n12696), .ZN(n10508) );
  NAND2_X1 U11495 ( .A1(n14033), .A2(n13677), .ZN(n19604) );
  AOI21_X1 U11496 ( .B1(n9747), .B2(n10579), .A(n10578), .ZN(n10577) );
  AND2_X1 U11497 ( .A1(n9959), .A2(n9958), .ZN(n12798) );
  INV_X2 U11498 ( .A(n11894), .ZN(n10450) );
  OR2_X2 U11499 ( .A1(n12087), .A2(n12073), .ZN(n10261) );
  NAND2_X2 U11500 ( .A1(n9926), .A2(n12218), .ZN(n14713) );
  CLKBUF_X1 U11501 ( .A(n13136), .Z(n14736) );
  OAI21_X1 U11502 ( .B1(n12879), .B2(n12235), .A(n12234), .ZN(n12236) );
  NAND2_X1 U11503 ( .A1(n12666), .A2(n12665), .ZN(n12664) );
  NAND2_X1 U11504 ( .A1(n11573), .A2(n11572), .ZN(n11575) );
  NAND2_X1 U11505 ( .A1(n10501), .A2(n12621), .ZN(n12665) );
  AND3_X1 U11506 ( .A1(n10665), .A2(n12176), .A3(n12175), .ZN(n13144) );
  NAND2_X1 U11507 ( .A1(n11202), .A2(n11201), .ZN(n11205) );
  OR2_X1 U11508 ( .A1(n12076), .A2(n13680), .ZN(n13676) );
  NAND3_X1 U11509 ( .A1(n9927), .A2(n14420), .A3(n14421), .ZN(n12218) );
  NAND2_X1 U11510 ( .A1(n12611), .A2(n16419), .ZN(n14748) );
  AND2_X1 U11511 ( .A1(n14426), .A2(n12551), .ZN(n12228) );
  NAND3_X1 U11512 ( .A1(n9940), .A2(n10163), .A3(n9929), .ZN(n13621) );
  INV_X1 U11513 ( .A(n11624), .ZN(n11649) );
  CLKBUF_X2 U11514 ( .A(n12918), .Z(n13127) );
  AND2_X1 U11515 ( .A1(n11806), .A2(n11807), .ZN(n10804) );
  AND2_X1 U11516 ( .A1(n12893), .A2(n12908), .ZN(n12920) );
  INV_X1 U11517 ( .A(n21825), .ZN(n11798) );
  NAND2_X1 U11518 ( .A1(n10921), .A2(n10920), .ZN(n11552) );
  CLKBUF_X1 U11519 ( .A(n10802), .Z(n16270) );
  OR2_X1 U11520 ( .A1(n12377), .A2(n12376), .ZN(n12909) );
  INV_X1 U11521 ( .A(n20433), .ZN(n12174) );
  OR2_X1 U11522 ( .A1(n12392), .A2(n12391), .ZN(n12591) );
  INV_X1 U11523 ( .A(n13674), .ZN(n19638) );
  INV_X1 U11524 ( .A(n12079), .ZN(n19642) );
  OR2_X1 U11525 ( .A1(n11557), .A2(n10799), .ZN(n10801) );
  OR2_X1 U11526 ( .A1(n12469), .A2(n12468), .ZN(n12938) );
  AND2_X2 U11527 ( .A1(n10799), .A2(n14591), .ZN(n10792) );
  NAND2_X1 U11528 ( .A1(n10795), .A2(n14577), .ZN(n11557) );
  AND2_X1 U11529 ( .A1(n11781), .A2(n14553), .ZN(n11805) );
  NAND4_X2 U11530 ( .A1(n12068), .A2(n12067), .A3(n12066), .A4(n12065), .ZN(
        n18973) );
  NAND4_X1 U11531 ( .A1(n11942), .A2(n11941), .A3(n11940), .A4(n11939), .ZN(
        n13690) );
  NAND4_X2 U11532 ( .A1(n11963), .A2(n11962), .A3(n11961), .A4(n11960), .ZN(
        n19654) );
  NAND4_X1 U11533 ( .A1(n12025), .A2(n12024), .A3(n12023), .A4(n12022), .ZN(
        n13685) );
  INV_X1 U11534 ( .A(n14238), .ZN(n9714) );
  AND4_X1 U11535 ( .A1(n11924), .A2(n11923), .A3(n11922), .A4(n11921), .ZN(
        n19646) );
  OAI21_X1 U11536 ( .B1(n10133), .B2(n10131), .A(n12129), .ZN(n10130) );
  NOR2_X1 U11537 ( .A1(n16904), .A2(n19863), .ZN(n20039) );
  INV_X1 U11538 ( .A(n10795), .ZN(n11799) );
  INV_X1 U11539 ( .A(n10162), .ZN(n10816) );
  CLKBUF_X3 U11540 ( .A(n14567), .Z(n9724) );
  INV_X2 U11541 ( .A(n14331), .ZN(n9715) );
  INV_X1 U11542 ( .A(n10769), .ZN(n11781) );
  INV_X2 U11543 ( .A(n15181), .ZN(n15148) );
  INV_X2 U11544 ( .A(U214), .ZN(n18189) );
  AND4_X2 U11545 ( .A1(n10715), .A2(n10714), .A3(n10713), .A4(n10712), .ZN(
        n10795) );
  NAND2_X2 U11546 ( .A1(n10736), .A2(n10687), .ZN(n14591) );
  AND4_X1 U11547 ( .A1(n12136), .A2(n12135), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A4(n12134), .ZN(n12138) );
  NAND2_X2 U11548 ( .A1(n20208), .A2(n20133), .ZN(n20185) );
  NAND2_X2 U11549 ( .A1(n20976), .A2(n20977), .ZN(n21033) );
  INV_X1 U11550 ( .A(n15173), .ZN(n13078) );
  AND4_X1 U11551 ( .A1(n10731), .A2(n10730), .A3(n10729), .A4(n10728), .ZN(
        n10736) );
  AND4_X1 U11552 ( .A1(n10693), .A2(n10692), .A3(n10691), .A4(n10690), .ZN(
        n10715) );
  AND4_X1 U11553 ( .A1(n10711), .A2(n10710), .A3(n10709), .A4(n10708), .ZN(
        n10712) );
  INV_X1 U11554 ( .A(n15176), .ZN(n15143) );
  AOI21_X1 U11555 ( .B1(n10780), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n10716), .ZN(n10720) );
  CLKBUF_X1 U11556 ( .A(n9736), .Z(n15320) );
  BUF_X2 U11557 ( .A(n10884), .Z(n10936) );
  INV_X2 U11558 ( .A(n18227), .ZN(U215) );
  AND2_X1 U11559 ( .A1(n10845), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n10716) );
  AND2_X2 U11560 ( .A1(n12577), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15176) );
  AND2_X2 U11562 ( .A1(n11898), .A2(n13787), .ZN(n18652) );
  INV_X1 U11563 ( .A(n15259), .ZN(n9723) );
  NOR2_X2 U11564 ( .A1(n19861), .A2(n19841), .ZN(n19933) );
  NAND2_X1 U11565 ( .A1(n11914), .A2(n11913), .ZN(n11955) );
  AND2_X2 U11566 ( .A1(n10700), .A2(n10707), .ZN(n10845) );
  AND2_X2 U11567 ( .A1(n10700), .A2(n10705), .ZN(n10780) );
  AND2_X2 U11568 ( .A1(n10706), .A2(n10707), .ZN(n10884) );
  INV_X2 U11569 ( .A(n18231), .ZN(n18233) );
  AND2_X1 U11570 ( .A1(n10694), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10706) );
  AND2_X2 U11571 ( .A1(n14351), .A2(n13805), .ZN(n10846) );
  AND3_X1 U11572 ( .A1(n14054), .A2(n13965), .A3(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11897) );
  NAND2_X1 U11573 ( .A1(n13261), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13262) );
  INV_X2 U11574 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n10952) );
  INV_X1 U11575 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10408) );
  INV_X2 U11576 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n21964) );
  NOR2_X4 U11577 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10700) );
  NOR2_X2 U11578 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14019) );
  NAND2_X1 U11579 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14031) );
  INV_X1 U11580 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14054) );
  INV_X1 U11581 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n22115) );
  NOR2_X1 U11582 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15153) );
  NAND2_X1 U11584 ( .A1(n10803), .A2(n10045), .ZN(n13562) );
  NAND3_X1 U11585 ( .A1(n10301), .A2(n15836), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15817) );
  INV_X1 U11586 ( .A(n12600), .ZN(n14866) );
  AOI211_X1 U11587 ( .C1(n17104), .C2(n18107), .A(n17103), .B(n17102), .ZN(
        n17105) );
  AND2_X2 U11588 ( .A1(n15428), .A2(n15430), .ZN(n15416) );
  OR2_X1 U11589 ( .A1(n10766), .A2(n10765), .ZN(n10162) );
  NAND2_X4 U11590 ( .A1(n14026), .A2(n13787), .ZN(n18773) );
  OR2_X1 U11591 ( .A1(n17101), .A2(n9873), .ZN(n9975) );
  INV_X4 U11592 ( .A(n12248), .ZN(n12809) );
  INV_X1 U11593 ( .A(n15158), .ZN(n9722) );
  INV_X2 U11594 ( .A(n15259), .ZN(n15323) );
  NAND2_X2 U11595 ( .A1(n10812), .A2(n10808), .ZN(n10834) );
  INV_X1 U11596 ( .A(n9987), .ZN(n9725) );
  AND2_X4 U11597 ( .A1(n12140), .A2(n12139), .ZN(n12898) );
  AND3_X2 U11598 ( .A1(n14513), .A2(n14827), .A3(n14600), .ZN(n14784) );
  NAND2_X2 U11599 ( .A1(n9992), .A2(n9991), .ZN(n9934) );
  OAI211_X1 U11600 ( .C1(n11042), .C2(n10352), .A(n10351), .B(n10349), .ZN(
        n11754) );
  NOR2_X2 U11601 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n18343), .ZN(n18332) );
  NOR2_X2 U11602 ( .A1(n14075), .A2(n10532), .ZN(n14451) );
  NAND2_X2 U11603 ( .A1(n9925), .A2(n9924), .ZN(n10172) );
  NAND2_X1 U11604 ( .A1(n10177), .A2(n14509), .ZN(n10176) );
  NAND2_X2 U11605 ( .A1(n11602), .A2(n11601), .ZN(n14875) );
  AND2_X1 U11606 ( .A1(n14684), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12310) );
  AND2_X1 U11607 ( .A1(n14708), .A2(n21964), .ZN(n9731) );
  XNOR2_X1 U11608 ( .A(n11887), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9733) );
  NOR2_X2 U11609 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n18326), .ZN(n18312) );
  NAND2_X1 U11610 ( .A1(n11569), .A2(n9724), .ZN(n11581) );
  NAND2_X1 U11611 ( .A1(n15035), .A2(n15034), .ZN(n21217) );
  INV_X1 U11612 ( .A(n12206), .ZN(n9735) );
  XNOR2_X2 U11613 ( .A(n15381), .B(n11856), .ZN(n15043) );
  NOR2_X2 U11614 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n18305), .ZN(n18290) );
  NOR2_X1 U11615 ( .A1(n10611), .A2(n10553), .ZN(n10552) );
  AOI21_X1 U11616 ( .B1(n16718), .B2(n14275), .A(n13837), .ZN(n13999) );
  INV_X2 U11617 ( .A(n9987), .ZN(n12631) );
  NOR2_X2 U11618 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n18284), .ZN(n18270) );
  NOR2_X2 U11619 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n18512), .ZN(n18491) );
  NAND2_X1 U11620 ( .A1(n11532), .A2(n11531), .ZN(n11537) );
  AND3_X1 U11621 ( .A1(n11799), .A2(n9724), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11509) );
  AND2_X1 U11622 ( .A1(n10052), .A2(n15457), .ZN(n10051) );
  INV_X1 U11623 ( .A(n11780), .ZN(n10098) );
  NAND2_X1 U11624 ( .A1(n14866), .A2(n20433), .ZN(n10365) );
  AND2_X1 U11625 ( .A1(n13835), .A2(n9715), .ZN(n15275) );
  NOR2_X1 U11626 ( .A1(n12551), .A2(n17596), .ZN(n13835) );
  NAND2_X1 U11627 ( .A1(n15063), .A2(n9875), .ZN(n16773) );
  NAND2_X1 U11628 ( .A1(n17490), .A2(n17489), .ZN(n17179) );
  AND2_X1 U11629 ( .A1(n15275), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n14280) );
  NAND2_X1 U11630 ( .A1(n9953), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9951) );
  INV_X1 U11631 ( .A(n10012), .ZN(n17767) );
  NAND2_X1 U11632 ( .A1(n13777), .A2(n18243), .ZN(n12087) );
  OR2_X1 U11633 ( .A1(n13694), .A2(n12102), .ZN(n13697) );
  INV_X1 U11634 ( .A(n18975), .ZN(n18243) );
  NOR2_X1 U11635 ( .A1(n10290), .A2(n11770), .ZN(n10143) );
  AND2_X1 U11636 ( .A1(n12619), .A2(n20237), .ZN(n13164) );
  NAND2_X1 U11637 ( .A1(n9832), .A2(n12220), .ZN(n9971) );
  INV_X1 U11638 ( .A(n10353), .ZN(n11032) );
  NAND2_X1 U11639 ( .A1(n10935), .A2(n9936), .ZN(n10180) );
  AND2_X1 U11640 ( .A1(n9967), .A2(n9760), .ZN(n9936) );
  NAND2_X1 U11641 ( .A1(n10968), .A2(n10969), .ZN(n10957) );
  AOI21_X1 U11642 ( .B1(n11537), .B2(n11536), .A(n11535), .ZN(n11546) );
  NOR2_X1 U11643 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n21303), .ZN(
        n11549) );
  NAND2_X1 U11644 ( .A1(n10595), .A2(n10594), .ZN(n10593) );
  INV_X1 U11645 ( .A(n10599), .ZN(n10594) );
  AND2_X1 U11646 ( .A1(n12905), .A2(n20834), .ZN(n12908) );
  AND2_X2 U11647 ( .A1(n14287), .A2(n14704), .ZN(n9962) );
  NAND2_X1 U11648 ( .A1(n14196), .A2(n14195), .ZN(n14207) );
  AND2_X1 U11649 ( .A1(n11409), .A2(n10635), .ZN(n10634) );
  NOR2_X1 U11650 ( .A1(n15433), .A2(n10636), .ZN(n10635) );
  INV_X1 U11651 ( .A(n15443), .ZN(n10636) );
  INV_X1 U11652 ( .A(n11472), .ZN(n11494) );
  NOR2_X1 U11653 ( .A1(n10625), .A2(n15529), .ZN(n10052) );
  NAND2_X1 U11654 ( .A1(n11318), .A2(n10626), .ZN(n10625) );
  AND2_X1 U11655 ( .A1(n10618), .A2(n11099), .ZN(n10048) );
  NOR2_X1 U11656 ( .A1(n10621), .A2(n10619), .ZN(n10618) );
  INV_X1 U11657 ( .A(n15538), .ZN(n10619) );
  INV_X1 U11658 ( .A(n14845), .ZN(n10049) );
  NAND2_X1 U11659 ( .A1(n10821), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11082) );
  INV_X1 U11660 ( .A(n15959), .ZN(n10293) );
  NAND2_X1 U11661 ( .A1(n9830), .A2(n11590), .ZN(n10536) );
  OR2_X1 U11662 ( .A1(n10353), .A2(n10352), .ZN(n10351) );
  AND2_X1 U11663 ( .A1(n11654), .A2(n14238), .ZN(n11624) );
  NAND2_X1 U11664 ( .A1(n11722), .A2(n11721), .ZN(n11729) );
  AND3_X1 U11665 ( .A1(n11684), .A2(n11805), .A3(n11685), .ZN(n13414) );
  AND2_X1 U11666 ( .A1(n14577), .A2(n14561), .ZN(n11784) );
  AND4_X1 U11667 ( .A1(n10824), .A2(n10823), .A3(n10822), .A4(n11816), .ZN(
        n10826) );
  AND3_X1 U11668 ( .A1(n10909), .A2(n10908), .A3(n10907), .ZN(n10910) );
  NAND2_X1 U11669 ( .A1(n10989), .A2(n10990), .ZN(n10858) );
  INV_X1 U11670 ( .A(n11509), .ZN(n11541) );
  AOI21_X1 U11671 ( .B1(n12565), .B2(n12563), .A(n12562), .ZN(n12569) );
  NOR2_X1 U11672 ( .A1(n12129), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12562) );
  INV_X1 U11673 ( .A(n12927), .ZN(n12919) );
  NAND2_X1 U11674 ( .A1(n10637), .A2(n10664), .ZN(n10222) );
  AND2_X1 U11675 ( .A1(n17076), .A2(n17066), .ZN(n10609) );
  NAND2_X1 U11676 ( .A1(n10337), .A2(n16695), .ZN(n10243) );
  INV_X1 U11677 ( .A(n12260), .ZN(n9959) );
  NOR2_X1 U11678 ( .A1(n12804), .A2(n14440), .ZN(n12805) );
  INV_X1 U11679 ( .A(n12253), .ZN(n9947) );
  NAND2_X1 U11680 ( .A1(n13995), .A2(n13994), .ZN(n13997) );
  AND2_X1 U11681 ( .A1(n15275), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n13996) );
  NAND2_X1 U11682 ( .A1(n13621), .A2(n9928), .ZN(n13136) );
  AND2_X1 U11683 ( .A1(n14428), .A2(n12215), .ZN(n9927) );
  AND2_X2 U11684 ( .A1(n10591), .A2(n9920), .ZN(n12611) );
  AND3_X1 U11685 ( .A1(n14032), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11898) );
  INV_X1 U11686 ( .A(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14943) );
  NOR2_X1 U11687 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11917) );
  INV_X1 U11688 ( .A(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17689) );
  NAND2_X1 U11689 ( .A1(n9836), .A2(n10333), .ZN(n10012) );
  NAND2_X1 U11690 ( .A1(n10007), .A2(n10429), .ZN(n17759) );
  AND2_X1 U11691 ( .A1(n10426), .A2(n19464), .ZN(n10007) );
  NAND2_X1 U11692 ( .A1(n19267), .A2(n14224), .ZN(n14225) );
  NAND2_X1 U11693 ( .A1(n19289), .A2(n14181), .ZN(n14183) );
  AND4_X1 U11694 ( .A1(n12008), .A2(n12007), .A3(n12006), .A4(n12005), .ZN(
        n12025) );
  AND4_X1 U11695 ( .A1(n12017), .A2(n12016), .A3(n12015), .A4(n12014), .ZN(
        n12023) );
  INV_X1 U11696 ( .A(n9703), .ZN(n11654) );
  AND2_X1 U11697 ( .A1(n15818), .A2(n10146), .ZN(n11860) );
  NOR2_X1 U11698 ( .A1(n10556), .A2(n10147), .ZN(n10146) );
  INV_X1 U11699 ( .A(n10667), .ZN(n10556) );
  NAND2_X1 U11700 ( .A1(n15818), .A2(n16029), .ZN(n10145) );
  NAND2_X1 U11701 ( .A1(n15827), .A2(n15817), .ZN(n15818) );
  NAND2_X1 U11702 ( .A1(n11791), .A2(n13800), .ZN(n11824) );
  AND2_X1 U11703 ( .A1(n18034), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13800) );
  AND4_X1 U11704 ( .A1(n10698), .A2(n10697), .A3(n10696), .A4(n10695), .ZN(
        n10714) );
  AND4_X1 U11705 ( .A1(n10704), .A2(n10703), .A3(n10702), .A4(n10701), .ZN(
        n10713) );
  NAND2_X1 U11706 ( .A1(n9707), .A2(n16317), .ZN(n21410) );
  NOR2_X1 U11707 ( .A1(n14335), .A2(n10639), .ZN(n10638) );
  INV_X1 U11708 ( .A(n14332), .ZN(n10639) );
  INV_X1 U11709 ( .A(n13210), .ZN(n10581) );
  AND2_X1 U11710 ( .A1(n13315), .A2(n13314), .ZN(n16990) );
  NAND2_X1 U11711 ( .A1(n16453), .A2(n12878), .ZN(n16441) );
  NAND2_X1 U11712 ( .A1(n10191), .A2(n10190), .ZN(n17010) );
  INV_X1 U11713 ( .A(n10339), .ZN(n17021) );
  NOR2_X1 U11714 ( .A1(n13355), .A2(n10607), .ZN(n10606) );
  INV_X1 U11715 ( .A(n17058), .ZN(n10607) );
  NAND2_X1 U11716 ( .A1(n12704), .A2(n10599), .ZN(n10598) );
  AND2_X1 U11717 ( .A1(n17364), .A2(n10398), .ZN(n17158) );
  INV_X1 U11718 ( .A(n14280), .ZN(n10225) );
  NAND2_X1 U11719 ( .A1(n10201), .A2(n9818), .ZN(n14854) );
  INV_X1 U11720 ( .A(n12575), .ZN(n10201) );
  AND4_X1 U11721 ( .A1(n11928), .A2(n11927), .A3(n11926), .A4(n11925), .ZN(
        n11942) );
  AND4_X1 U11722 ( .A1(n11938), .A2(n11937), .A3(n11936), .A4(n11935), .ZN(
        n11939) );
  AND4_X1 U11723 ( .A1(n12000), .A2(n11999), .A3(n11998), .A4(n11997), .ZN(
        n12001) );
  AND4_X1 U11724 ( .A1(n11989), .A2(n11988), .A3(n11987), .A4(n11986), .ZN(
        n12004) );
  AND4_X1 U11725 ( .A1(n11993), .A2(n11992), .A3(n11991), .A4(n11990), .ZN(
        n12003) );
  NAND2_X1 U11726 ( .A1(n9829), .A2(n9741), .ZN(n10471) );
  AND4_X1 U11727 ( .A1(n14136), .A2(n14135), .A3(n14134), .A4(n14133), .ZN(
        n14145) );
  NAND2_X1 U11728 ( .A1(n10261), .A2(n9740), .ZN(n10260) );
  AOI21_X1 U11729 ( .B1(n13677), .B2(n9740), .A(n9878), .ZN(n10257) );
  NOR2_X1 U11730 ( .A1(n10473), .A2(n10472), .ZN(n13872) );
  INV_X1 U11731 ( .A(n20059), .ZN(n10472) );
  NAND2_X1 U11732 ( .A1(n9834), .A2(n10015), .ZN(n17764) );
  NAND2_X1 U11733 ( .A1(n17760), .A2(n19073), .ZN(n10015) );
  OAI21_X1 U11734 ( .B1(n19302), .B2(n10011), .A(n10009), .ZN(n14214) );
  INV_X1 U11735 ( .A(n10010), .ZN(n10009) );
  OAI21_X1 U11736 ( .B1(n14205), .B2(n10011), .A(n19286), .ZN(n10010) );
  AND2_X1 U11737 ( .A1(n14205), .A2(n10011), .ZN(n10008) );
  AND4_X1 U11738 ( .A1(n11906), .A2(n11905), .A3(n11904), .A4(n11903), .ZN(
        n11923) );
  AND4_X1 U11739 ( .A1(n11902), .A2(n11901), .A3(n11900), .A4(n11899), .ZN(
        n11924) );
  NOR2_X1 U11740 ( .A1(n20109), .A2(n20107), .ZN(n20212) );
  AND2_X1 U11741 ( .A1(n15373), .A2(n15371), .ZN(n21820) );
  OR2_X1 U11742 ( .A1(n16429), .A2(n10494), .ZN(n10493) );
  NAND2_X1 U11743 ( .A1(n10495), .A2(n16428), .ZN(n10494) );
  OR2_X1 U11744 ( .A1(n16984), .A2(n20345), .ZN(n10159) );
  INV_X1 U11745 ( .A(n10194), .ZN(n10044) );
  OAI21_X1 U11746 ( .B1(n15343), .B2(n18123), .A(n15354), .ZN(n10194) );
  OAI21_X1 U11747 ( .B1(n17370), .B2(n17518), .A(n17369), .ZN(n10255) );
  INV_X1 U11748 ( .A(n17375), .ZN(n10613) );
  INV_X1 U11749 ( .A(n17505), .ZN(n18123) );
  NAND2_X1 U11750 ( .A1(n13881), .A2(P3_EAX_REG_0__SCAN_IN), .ZN(n13882) );
  OAI22_X1 U11751 ( .A1(n20494), .A2(n15142), .B1(n13058), .B2(n9934), .ZN(
        n12482) );
  NAND2_X1 U11752 ( .A1(n11011), .A2(n11010), .ZN(n11030) );
  INV_X1 U11753 ( .A(n10221), .ZN(n10220) );
  OAI21_X1 U11754 ( .B1(n10217), .B2(n12291), .A(n13145), .ZN(n10221) );
  NAND2_X1 U11755 ( .A1(n10219), .A2(n10218), .ZN(n10217) );
  NOR2_X1 U11756 ( .A1(n12280), .A2(n12281), .ZN(n10231) );
  NAND2_X1 U11757 ( .A1(n9787), .A2(n9752), .ZN(n9970) );
  AND2_X1 U11758 ( .A1(n15157), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n9914) );
  NAND2_X1 U11759 ( .A1(n10568), .A2(n15979), .ZN(n10567) );
  INV_X1 U11760 ( .A(n10570), .ZN(n10568) );
  NAND2_X1 U11761 ( .A1(n14557), .A2(n11557), .ZN(n9932) );
  NAND2_X1 U11762 ( .A1(n10802), .A2(n14553), .ZN(n10770) );
  AOI21_X1 U11763 ( .B1(n10079), .B2(n11528), .A(n9816), .ZN(n10082) );
  INV_X1 U11764 ( .A(n11523), .ZN(n10079) );
  INV_X1 U11765 ( .A(n11528), .ZN(n10083) );
  NOR2_X1 U11766 ( .A1(n13279), .A2(n10500), .ZN(n10499) );
  AND2_X1 U11767 ( .A1(n17058), .A2(n12703), .ZN(n10070) );
  NAND2_X1 U11768 ( .A1(n12205), .A2(n12204), .ZN(n12230) );
  NAND2_X1 U11769 ( .A1(n14422), .A2(n12211), .ZN(n12204) );
  OAI21_X1 U11770 ( .B1(n12557), .B2(n10198), .A(n10197), .ZN(n12572) );
  NAND2_X1 U11771 ( .A1(n12207), .A2(n12594), .ZN(n10197) );
  OAI21_X1 U11772 ( .B1(n15209), .B2(n10200), .A(n10199), .ZN(n10198) );
  NOR2_X1 U11773 ( .A1(n10323), .A2(n10326), .ZN(n10325) );
  INV_X1 U11774 ( .A(n17762), .ZN(n10326) );
  AND2_X1 U11775 ( .A1(n13771), .A2(n19650), .ZN(n12076) );
  INV_X1 U11776 ( .A(n11555), .ZN(n13792) );
  AND3_X1 U11777 ( .A1(n10821), .A2(n10795), .A3(n10816), .ZN(n10796) );
  NOR2_X1 U11778 ( .A1(n10627), .A2(n15480), .ZN(n10626) );
  INV_X1 U11779 ( .A(n10629), .ZN(n10627) );
  NOR2_X1 U11780 ( .A1(n10630), .A2(n15505), .ZN(n10629) );
  INV_X1 U11781 ( .A(n15493), .ZN(n10630) );
  INV_X1 U11782 ( .A(n15504), .ZN(n10628) );
  NAND2_X1 U11783 ( .A1(n11186), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11472) );
  INV_X1 U11784 ( .A(n11082), .ZN(n11174) );
  INV_X1 U11785 ( .A(n15399), .ZN(n10537) );
  NOR2_X1 U11786 ( .A1(n10539), .A2(n15403), .ZN(n10538) );
  INV_X1 U11787 ( .A(n15417), .ZN(n10539) );
  INV_X1 U11788 ( .A(n10567), .ZN(n10298) );
  AOI21_X1 U11789 ( .B1(n10570), .B2(n15909), .A(n15909), .ZN(n10296) );
  NAND2_X1 U11790 ( .A1(n15898), .A2(n10570), .ZN(n10142) );
  NAND2_X1 U11791 ( .A1(n10567), .A2(n15898), .ZN(n10171) );
  INV_X1 U11792 ( .A(n16093), .ZN(n10573) );
  NAND2_X1 U11793 ( .A1(n10674), .A2(n10544), .ZN(n10543) );
  INV_X1 U11794 ( .A(n15616), .ZN(n10544) );
  NAND2_X1 U11795 ( .A1(n10172), .A2(n11763), .ZN(n15952) );
  NAND2_X1 U11796 ( .A1(n11762), .A2(n9922), .ZN(n9921) );
  INV_X1 U11797 ( .A(n15705), .ZN(n10535) );
  MUX2_X1 U11798 ( .A(n11576), .B(n9734), .S(P1_EBX_REG_1__SCAN_IN), .Z(n11573) );
  OR2_X1 U11799 ( .A1(n10899), .A2(n10898), .ZN(n11724) );
  OR2_X1 U11800 ( .A1(n10883), .A2(n10882), .ZN(n11755) );
  INV_X1 U11801 ( .A(n10812), .ZN(n10833) );
  INV_X1 U11802 ( .A(n11557), .ZN(n11808) );
  INV_X1 U11803 ( .A(n14752), .ZN(n16317) );
  INV_X1 U11804 ( .A(n10934), .ZN(n9968) );
  XNOR2_X1 U11805 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12563) );
  NAND2_X1 U11806 ( .A1(n12561), .A2(n12560), .ZN(n12565) );
  INV_X1 U11807 ( .A(n12687), .ZN(n10506) );
  INV_X1 U11808 ( .A(n12938), .ZN(n12624) );
  NAND2_X1 U11809 ( .A1(n12656), .A2(n10059), .ZN(n10058) );
  INV_X1 U11810 ( .A(n12657), .ZN(n10059) );
  AND2_X1 U11811 ( .A1(n9717), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10065) );
  CLKBUF_X1 U11812 ( .A(n12311), .Z(n15326) );
  INV_X1 U11813 ( .A(n16753), .ZN(n10648) );
  NOR2_X1 U11814 ( .A1(n16748), .A2(n10644), .ZN(n10643) );
  INV_X1 U11815 ( .A(n10650), .ZN(n10644) );
  OR2_X1 U11816 ( .A1(n15235), .A2(n15236), .ZN(n10661) );
  AND2_X1 U11817 ( .A1(n9746), .A2(n10228), .ZN(n10227) );
  INV_X1 U11818 ( .A(n16792), .ZN(n10228) );
  AND2_X1 U11819 ( .A1(n9795), .A2(n10590), .ZN(n10589) );
  INV_X1 U11820 ( .A(n16591), .ZN(n10590) );
  INV_X1 U11821 ( .A(n14639), .ZN(n10582) );
  INV_X1 U11822 ( .A(n14631), .ZN(n12987) );
  AND3_X1 U11823 ( .A1(n10676), .A2(n12361), .A3(n12360), .ZN(n12904) );
  INV_X1 U11824 ( .A(n12359), .ZN(n12360) );
  AND2_X1 U11825 ( .A1(n10485), .A2(n13233), .ZN(n10483) );
  AND4_X1 U11826 ( .A1(n12519), .A2(n12518), .A3(n12517), .A4(n12516), .ZN(
        n12538) );
  INV_X1 U11827 ( .A(n12776), .ZN(n10112) );
  AND2_X1 U11828 ( .A1(n9849), .A2(n16537), .ZN(n10039) );
  AND2_X1 U11829 ( .A1(n10586), .A2(n9898), .ZN(n10585) );
  AND2_X1 U11830 ( .A1(n9869), .A2(n16512), .ZN(n10586) );
  INV_X1 U11831 ( .A(n13362), .ZN(n10196) );
  AOI21_X1 U11832 ( .B1(n10600), .B2(n17107), .A(n10249), .ZN(n10248) );
  INV_X1 U11833 ( .A(n17110), .ZN(n10249) );
  INV_X1 U11834 ( .A(n10393), .ZN(n10392) );
  OAI21_X1 U11835 ( .B1(n10395), .B2(n10394), .A(n10609), .ZN(n10393) );
  NOR2_X1 U11836 ( .A1(n17097), .A2(n10394), .ZN(n10390) );
  NAND2_X1 U11837 ( .A1(n10383), .A2(n10592), .ZN(n17106) );
  AND2_X1 U11838 ( .A1(n10593), .A2(n10601), .ZN(n10592) );
  AND2_X1 U11839 ( .A1(n13346), .A2(n17132), .ZN(n10601) );
  AND2_X1 U11840 ( .A1(n10516), .A2(n14822), .ZN(n10042) );
  AND2_X1 U11841 ( .A1(n10518), .A2(n10517), .ZN(n10516) );
  INV_X1 U11842 ( .A(n16614), .ZN(n10517) );
  INV_X1 U11843 ( .A(n14647), .ZN(n12840) );
  INV_X1 U11844 ( .A(n14337), .ZN(n10515) );
  AOI21_X1 U11845 ( .B1(n9819), .B2(n12690), .A(n16682), .ZN(n10369) );
  NAND2_X1 U11846 ( .A1(n10550), .A2(n9742), .ZN(n9974) );
  NAND2_X1 U11847 ( .A1(n12242), .A2(n9960), .ZN(n12243) );
  INV_X1 U11848 ( .A(n14420), .ZN(n10125) );
  INV_X1 U11849 ( .A(n12597), .ZN(n12574) );
  NOR2_X1 U11850 ( .A1(n12300), .A2(n12129), .ZN(n12577) );
  NAND2_X1 U11851 ( .A1(n9991), .A2(n9802), .ZN(n12426) );
  NOR2_X1 U11852 ( .A1(n9848), .A2(n10024), .ZN(n10137) );
  AOI21_X1 U11853 ( .B1(n9730), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A(
        n12129), .ZN(n10025) );
  NAND2_X1 U11854 ( .A1(n9719), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n10136) );
  NAND2_X1 U11855 ( .A1(n9729), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n9997) );
  NAND2_X1 U11856 ( .A1(n9955), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9949) );
  INV_X1 U11857 ( .A(n12013), .ZN(n17608) );
  AND4_X1 U11858 ( .A1(n13947), .A2(n13946), .A3(n13945), .A4(n13944), .ZN(
        n13961) );
  AND4_X1 U11859 ( .A1(n13891), .A2(n13890), .A3(n13889), .A4(n13888), .ZN(
        n13907) );
  NAND2_X1 U11860 ( .A1(n14209), .A2(n14208), .ZN(n14218) );
  INV_X1 U11861 ( .A(n17766), .ZN(n10333) );
  AND2_X1 U11862 ( .A1(n19476), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17891) );
  OR2_X1 U11863 ( .A1(n17856), .A2(n19174), .ZN(n19403) );
  INV_X1 U11864 ( .A(n14401), .ZN(n10303) );
  OR2_X1 U11865 ( .A1(n19650), .A2(n19646), .ZN(n13691) );
  NOR2_X1 U11866 ( .A1(n13775), .A2(n13787), .ZN(n13840) );
  NAND4_X1 U11867 ( .A1(n11985), .A2(n11984), .A3(n11983), .A4(n11982), .ZN(
        n12079) );
  AND4_X1 U11868 ( .A1(n11981), .A2(n11980), .A3(n11979), .A4(n11978), .ZN(
        n11982) );
  AND4_X1 U11869 ( .A1(n11967), .A2(n11966), .A3(n11965), .A4(n11964), .ZN(
        n11985) );
  AND2_X1 U11870 ( .A1(n13575), .A2(n13573), .ZN(n13563) );
  AND2_X1 U11871 ( .A1(n11614), .A2(n11613), .ZN(n15599) );
  NAND2_X1 U11872 ( .A1(n10794), .A2(n10793), .ZN(n14064) );
  INV_X1 U11873 ( .A(n14577), .ZN(n10793) );
  OR2_X1 U11874 ( .A1(n13794), .A2(n11819), .ZN(n14063) );
  NAND2_X1 U11875 ( .A1(n13419), .A2(n13418), .ZN(n13798) );
  OR2_X1 U11876 ( .A1(n17992), .A2(n13416), .ZN(n13419) );
  AND2_X1 U11877 ( .A1(n13806), .A2(n13415), .ZN(n13416) );
  AND2_X1 U11878 ( .A1(n10632), .A2(n10051), .ZN(n10050) );
  NOR2_X1 U11879 ( .A1(n10633), .A2(n15407), .ZN(n10632) );
  INV_X1 U11880 ( .A(n10634), .ZN(n10633) );
  NAND2_X1 U11881 ( .A1(n11388), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11410) );
  INV_X1 U11882 ( .A(n11389), .ZN(n11388) );
  NAND2_X1 U11883 ( .A1(n11281), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11319) );
  AND2_X1 U11884 ( .A1(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11201) );
  INV_X1 U11885 ( .A(n11200), .ZN(n11202) );
  AND2_X1 U11886 ( .A1(n10624), .A2(n14846), .ZN(n10623) );
  NAND2_X1 U11887 ( .A1(n16061), .A2(n16137), .ZN(n11837) );
  AND2_X1 U11888 ( .A1(n9868), .A2(n10546), .ZN(n10545) );
  INV_X1 U11889 ( .A(n15482), .ZN(n10546) );
  NAND2_X1 U11890 ( .A1(n9800), .A2(n10290), .ZN(n10289) );
  AND2_X1 U11891 ( .A1(n16088), .A2(n16087), .ZN(n16190) );
  AOI22_X1 U11892 ( .A1(n10176), .A2(n11707), .B1(n14507), .B2(n9904), .ZN(
        n10175) );
  OR2_X1 U11893 ( .A1(n11824), .A2(n17995), .ZN(n16186) );
  OR2_X1 U11894 ( .A1(n11824), .A2(n13807), .ZN(n16203) );
  INV_X1 U11895 ( .A(n10858), .ZN(n10828) );
  AOI21_X1 U11896 ( .B1(n10834), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n10835), .ZN(n10839) );
  INV_X1 U11897 ( .A(n14754), .ZN(n21564) );
  OR2_X1 U11898 ( .A1(n14391), .A2(n14390), .ZN(n21455) );
  NOR2_X1 U11899 ( .A1(n14608), .A2(n21309), .ZN(n21565) );
  NOR2_X1 U11900 ( .A1(n14757), .A2(n16325), .ZN(n21457) );
  INV_X1 U11901 ( .A(n16321), .ZN(n14757) );
  AOI21_X1 U11902 ( .B1(n21561), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n14757), 
        .ZN(n21677) );
  OR2_X1 U11903 ( .A1(n10103), .A2(n11534), .ZN(n10102) );
  NAND2_X1 U11904 ( .A1(n9833), .A2(n9753), .ZN(n10099) );
  NAND2_X1 U11905 ( .A1(n10101), .A2(n11554), .ZN(n10100) );
  INV_X1 U11906 ( .A(n11545), .ZN(n10101) );
  NAND2_X1 U11907 ( .A1(n9941), .A2(n12206), .ZN(n10406) );
  NOR2_X1 U11908 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n16421) );
  NAND2_X1 U11909 ( .A1(n13312), .A2(n10487), .ZN(n13319) );
  NAND2_X1 U11910 ( .A1(n13312), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13317) );
  AND2_X1 U11911 ( .A1(n9805), .A2(n12634), .ZN(n10512) );
  NAND2_X1 U11912 ( .A1(n16577), .A2(n17090), .ZN(n16559) );
  OR2_X1 U11913 ( .A1(n20313), .A2(n17174), .ZN(n16635) );
  NAND2_X1 U11914 ( .A1(n9799), .A2(n20324), .ZN(n16681) );
  INV_X1 U11915 ( .A(n16722), .ZN(n10153) );
  AND2_X1 U11916 ( .A1(n10154), .A2(n17243), .ZN(n10152) );
  INV_X1 U11917 ( .A(n16742), .ZN(n16692) );
  OR2_X1 U11918 ( .A1(n13053), .A2(n13052), .ZN(n15056) );
  OR2_X1 U11919 ( .A1(n12983), .A2(n12982), .ZN(n14820) );
  AND2_X1 U11920 ( .A1(n10651), .A2(n16753), .ZN(n10650) );
  NAND2_X2 U11921 ( .A1(n10222), .A2(n15277), .ZN(n16752) );
  XNOR2_X1 U11922 ( .A(n15256), .B(n10672), .ZN(n16764) );
  AND3_X1 U11923 ( .A1(n13005), .A2(n13004), .A3(n13003), .ZN(n14603) );
  AND3_X1 U11924 ( .A1(n12966), .A2(n12965), .A3(n12964), .ZN(n14627) );
  OAI21_X1 U11925 ( .B1(n12152), .B2(n12151), .A(n12129), .ZN(n12159) );
  NAND2_X1 U11926 ( .A1(n14854), .A2(n13145), .ZN(n13627) );
  INV_X1 U11927 ( .A(n13238), .ZN(n10420) );
  NAND2_X1 U11928 ( .A1(n10165), .A2(n10167), .ZN(n13215) );
  INV_X1 U11929 ( .A(n17011), .ZN(n10165) );
  NAND2_X1 U11930 ( .A1(n10189), .A2(n10188), .ZN(n10187) );
  INV_X1 U11931 ( .A(n16996), .ZN(n10188) );
  OAI21_X1 U11932 ( .B1(n17010), .B2(n16995), .A(n17007), .ZN(n10189) );
  INV_X1 U11933 ( .A(n10666), .ZN(n9978) );
  NAND2_X1 U11934 ( .A1(n13371), .A2(n10524), .ZN(n16511) );
  AND2_X1 U11935 ( .A1(n13105), .A2(n13104), .ZN(n13366) );
  OAI21_X1 U11936 ( .B1(n17098), .B2(n10387), .A(n10392), .ZN(n10608) );
  INV_X1 U11937 ( .A(n10390), .ZN(n10387) );
  OR2_X1 U11938 ( .A1(n10392), .A2(n13355), .ZN(n10386) );
  NAND2_X1 U11939 ( .A1(n10390), .A2(n13354), .ZN(n10389) );
  AND2_X1 U11940 ( .A1(n17364), .A2(n9911), .ZN(n17137) );
  NAND2_X1 U11941 ( .A1(n17364), .A2(n9776), .ZN(n17143) );
  NAND2_X1 U11942 ( .A1(n17179), .A2(n12695), .ZN(n12704) );
  AND2_X1 U11943 ( .A1(n17475), .A2(n13169), .ZN(n17453) );
  NAND2_X1 U11944 ( .A1(n12625), .A2(n13090), .ZN(n10579) );
  AND2_X1 U11945 ( .A1(n12673), .A2(n10529), .ZN(n10528) );
  NAND2_X1 U11946 ( .A1(n9791), .A2(n10241), .ZN(n10240) );
  NAND2_X1 U11947 ( .A1(n10530), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10529) );
  INV_X1 U11948 ( .A(n9791), .ZN(n10242) );
  NAND2_X1 U11949 ( .A1(n10238), .A2(n10550), .ZN(n10235) );
  NAND2_X1 U11950 ( .A1(n12800), .A2(n12799), .ZN(n12804) );
  NAND2_X1 U11951 ( .A1(n12805), .A2(n14439), .ZN(n14336) );
  NAND2_X1 U11952 ( .A1(n10212), .A2(n10211), .ZN(n12420) );
  NAND2_X1 U11953 ( .A1(n10210), .A2(n10208), .ZN(n10317) );
  AND2_X1 U11954 ( .A1(n13164), .A2(n21088), .ZN(n12796) );
  NOR2_X1 U11955 ( .A1(n17539), .A2(n13829), .ZN(n14849) );
  AND3_X1 U11956 ( .A1(n10226), .A2(n14435), .A3(n14281), .ZN(n10224) );
  INV_X1 U11957 ( .A(n14856), .ZN(n14275) );
  NAND2_X2 U11958 ( .A1(n13254), .A2(n13253), .ZN(n20350) );
  NAND2_X1 U11959 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13253) );
  NAND2_X1 U11960 ( .A1(n13252), .A2(n17596), .ZN(n13254) );
  NOR2_X2 U11961 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n21042) );
  OAI21_X2 U11962 ( .B1(n18136), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n14858), 
        .ZN(n20896) );
  NAND2_X1 U11963 ( .A1(n12438), .A2(n20895), .ZN(n20903) );
  OR2_X1 U11964 ( .A1(n18269), .A2(n20183), .ZN(n10456) );
  NAND2_X1 U11965 ( .A1(n18596), .A2(P3_EBX_REG_29__SCAN_IN), .ZN(n10455) );
  NOR2_X1 U11966 ( .A1(n18313), .A2(n10450), .ZN(n18300) );
  NOR2_X1 U11967 ( .A1(n18330), .A2(n10450), .ZN(n18321) );
  AND3_X1 U11968 ( .A1(n14128), .A2(n14127), .A3(n14126), .ZN(n14206) );
  AND4_X1 U11969 ( .A1(n14121), .A2(n14120), .A3(n14119), .A4(n14118), .ZN(
        n14127) );
  AND4_X1 U11970 ( .A1(n14117), .A2(n14116), .A3(n14115), .A4(n14114), .ZN(
        n14128) );
  AND4_X1 U11971 ( .A1(n13921), .A2(n13920), .A3(n13919), .A4(n13918), .ZN(
        n13926) );
  AND4_X1 U11972 ( .A1(n13634), .A2(n13633), .A3(n13632), .A4(n13631), .ZN(
        n13650) );
  AND4_X1 U11973 ( .A1(n12041), .A2(n12040), .A3(n12039), .A4(n12038), .ZN(
        n12042) );
  AND4_X1 U11974 ( .A1(n12029), .A2(n12028), .A3(n12027), .A4(n12026), .ZN(
        n12045) );
  NAND2_X1 U11975 ( .A1(n9794), .A2(n19132), .ZN(n19070) );
  CLKBUF_X1 U11976 ( .A(n11877), .Z(n11878) );
  AND4_X1 U11977 ( .A1(n12064), .A2(n12063), .A3(n12062), .A4(n12061), .ZN(
        n12065) );
  AND4_X1 U11978 ( .A1(n12057), .A2(n12056), .A3(n12055), .A4(n12054), .ZN(
        n12067) );
  NOR2_X1 U11979 ( .A1(n12060), .A2(n12059), .ZN(n12066) );
  NAND2_X1 U11980 ( .A1(n17759), .A2(n19196), .ZN(n19132) );
  NOR2_X1 U11981 ( .A1(n12072), .A2(n12071), .ZN(n12073) );
  OR2_X1 U11982 ( .A1(n13876), .A2(n12070), .ZN(n12072) );
  NAND2_X1 U11983 ( .A1(n9827), .A2(n19198), .ZN(n17844) );
  AND4_X1 U11984 ( .A1(n14161), .A2(n14160), .A3(n14159), .A4(n14158), .ZN(
        n14162) );
  NAND2_X1 U11985 ( .A1(n19279), .A2(n14184), .ZN(n19264) );
  INV_X1 U11986 ( .A(n19273), .ZN(n10431) );
  AND2_X1 U11987 ( .A1(n13698), .A2(n12105), .ZN(n20062) );
  OR2_X1 U11988 ( .A1(n13697), .A2(n12104), .ZN(n12105) );
  INV_X1 U11989 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21528) );
  INV_X1 U11990 ( .A(n15654), .ZN(n21168) );
  AND2_X1 U11991 ( .A1(n11672), .A2(n11657), .ZN(n21209) );
  INV_X1 U11992 ( .A(n18057), .ZN(n18052) );
  XNOR2_X1 U11993 ( .A(n11863), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16010) );
  NAND2_X1 U11994 ( .A1(n10087), .A2(n16042), .ZN(n16021) );
  OR2_X1 U11995 ( .A1(n11839), .A2(n16029), .ZN(n10087) );
  NAND2_X1 U11996 ( .A1(n16240), .A2(n10088), .ZN(n16108) );
  NAND2_X1 U11997 ( .A1(n10092), .A2(n10089), .ZN(n10088) );
  NOR2_X1 U11998 ( .A1(n10097), .A2(n10090), .ZN(n10089) );
  AND2_X1 U11999 ( .A1(n16096), .A2(n16234), .ZN(n10092) );
  OR2_X1 U12000 ( .A1(n11824), .A2(n11802), .ZN(n21293) );
  INV_X1 U12001 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21561) );
  INV_X1 U12002 ( .A(n11716), .ZN(n10980) );
  INV_X1 U12003 ( .A(n10978), .ZN(n10979) );
  AOI21_X1 U12004 ( .B1(n16434), .B2(n16980), .A(n10160), .ZN(n16426) );
  AOI21_X1 U12005 ( .B1(n16859), .B2(n20330), .A(n10157), .ZN(n10156) );
  NAND2_X1 U12006 ( .A1(n16436), .A2(n10158), .ZN(n10157) );
  AOI21_X1 U12007 ( .B1(n20262), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n16435), .ZN(n10158) );
  AND2_X1 U12008 ( .A1(n13325), .A2(n13324), .ZN(n20330) );
  NAND2_X1 U12009 ( .A1(n20350), .A2(n20326), .ZN(n16740) );
  NAND2_X1 U12010 ( .A1(n13132), .A2(n13181), .ZN(n16853) );
  NAND2_X1 U12011 ( .A1(n20417), .A2(n10104), .ZN(n13736) );
  OAI21_X1 U12012 ( .B1(n13205), .B2(n13207), .A(n13206), .ZN(n16984) );
  NAND2_X1 U12013 ( .A1(n16992), .A2(n18108), .ZN(n10286) );
  AOI21_X1 U12014 ( .B1(n17260), .B2(n18107), .A(n16993), .ZN(n10459) );
  NAND2_X1 U12015 ( .A1(n20274), .A2(n18107), .ZN(n10435) );
  INV_X1 U12016 ( .A(n17073), .ZN(n10434) );
  NAND2_X1 U12017 ( .A1(n10397), .A2(n13351), .ZN(n17087) );
  INV_X1 U12018 ( .A(n18102), .ZN(n17244) );
  XNOR2_X1 U12019 ( .A(n13219), .B(n13218), .ZN(n15352) );
  NAND2_X1 U12020 ( .A1(n13240), .A2(n13237), .ZN(n10106) );
  NAND2_X1 U12021 ( .A1(n10413), .A2(n10415), .ZN(n13240) );
  AND2_X1 U12022 ( .A1(n16971), .A2(n18118), .ZN(n13191) );
  OR2_X1 U12023 ( .A1(n13219), .A2(n13179), .ZN(n16970) );
  NOR2_X1 U12024 ( .A1(n10381), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10377) );
  NAND2_X1 U12025 ( .A1(n17011), .A2(n17266), .ZN(n10343) );
  NAND2_X1 U12026 ( .A1(n17021), .A2(n10338), .ZN(n10001) );
  OAI211_X1 U12027 ( .C1(n17364), .C2(n17035), .A(n10120), .B(n10119), .ZN(
        n17313) );
  OR2_X1 U12028 ( .A1(n13362), .A2(n17035), .ZN(n10120) );
  AOI21_X1 U12029 ( .B1(n10604), .B2(n10606), .A(n10603), .ZN(n10602) );
  NAND2_X1 U12030 ( .A1(n13363), .A2(n17036), .ZN(n17056) );
  NAND2_X1 U12031 ( .A1(n10404), .A2(n13370), .ZN(n13363) );
  OAI21_X1 U12032 ( .B1(n17364), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n10054), .ZN(n10057) );
  NOR2_X1 U12033 ( .A1(n17500), .A2(n10055), .ZN(n10054) );
  NOR2_X1 U12034 ( .A1(n9770), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10055) );
  XNOR2_X1 U12035 ( .A(n10232), .B(n17068), .ZN(n17350) );
  NAND2_X1 U12036 ( .A1(n10233), .A2(n17075), .ZN(n10232) );
  NAND2_X1 U12037 ( .A1(n17078), .A2(n17076), .ZN(n10233) );
  NOR2_X1 U12038 ( .A1(n18129), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10253) );
  NAND2_X1 U12039 ( .A1(n10027), .A2(n10030), .ZN(n17377) );
  NAND2_X1 U12040 ( .A1(n17364), .A2(n10032), .ZN(n10027) );
  INV_X1 U12041 ( .A(n17371), .ZN(n10251) );
  OAI21_X1 U12042 ( .B1(n17364), .B2(n10031), .A(n10028), .ZN(n10033) );
  AOI21_X1 U12043 ( .B1(n10030), .B2(n10029), .A(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10028) );
  INV_X1 U12044 ( .A(n10032), .ZN(n10029) );
  NAND2_X1 U12045 ( .A1(n17364), .A2(n9908), .ZN(n10043) );
  AND2_X1 U12046 ( .A1(n13164), .A2(n13138), .ZN(n17505) );
  INV_X1 U12047 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21083) );
  INV_X1 U12048 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21054) );
  NAND2_X1 U12049 ( .A1(n14854), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n18136) );
  NOR2_X1 U12050 ( .A1(n20061), .A2(n18976), .ZN(n20233) );
  NAND2_X1 U12051 ( .A1(n20233), .A2(n18917), .ZN(n20231) );
  XNOR2_X1 U12052 ( .A(n11895), .B(n17802), .ZN(n11896) );
  NOR2_X1 U12053 ( .A1(n18266), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n12117) );
  NOR2_X1 U12054 ( .A1(n21986), .A2(n18589), .ZN(n18481) );
  INV_X1 U12055 ( .A(n18481), .ZN(n18593) );
  NOR2_X2 U12056 ( .A1(n20231), .A2(n20097), .ZN(n18578) );
  NOR2_X1 U12057 ( .A1(n10477), .A2(n17649), .ZN(n18706) );
  NOR2_X1 U12058 ( .A1(n18781), .A2(n18784), .ZN(n13850) );
  AND4_X1 U12059 ( .A1(n11959), .A2(n11958), .A3(n11957), .A4(n11956), .ZN(
        n11960) );
  AND4_X1 U12060 ( .A1(n11954), .A2(n11953), .A3(n11952), .A4(n11951), .ZN(
        n11961) );
  AND4_X1 U12061 ( .A1(n11950), .A2(n11949), .A3(n11948), .A4(n11947), .ZN(
        n11962) );
  AND2_X1 U12062 ( .A1(n18880), .A2(n10274), .ZN(n18857) );
  NOR2_X1 U12063 ( .A1(n19023), .A2(n17735), .ZN(n18880) );
  INV_X1 U12064 ( .A(n18872), .ZN(n18878) );
  INV_X1 U12065 ( .A(n18864), .ZN(n18877) );
  NAND2_X1 U12066 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n9896), .ZN(n10270) );
  INV_X1 U12067 ( .A(n18911), .ZN(n18883) );
  AND2_X1 U12068 ( .A1(n13878), .A2(n20212), .ZN(n13881) );
  AND2_X1 U12069 ( .A1(n13881), .A2(n13964), .ZN(n18911) );
  OR2_X1 U12070 ( .A1(n19026), .A2(n19196), .ZN(n10005) );
  INV_X1 U12071 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18914) );
  INV_X1 U12072 ( .A(n19362), .ZN(n10004) );
  OR2_X1 U12073 ( .A1(n19598), .A2(n19566), .ZN(n19564) );
  INV_X1 U12074 ( .A(n19564), .ZN(n19602) );
  OAI22_X1 U12075 ( .A1(n14853), .A2(n12472), .B1(n12438), .B2(n12491), .ZN(
        n12474) );
  OAI22_X1 U12076 ( .A1(n14853), .A2(n12439), .B1(n12438), .B2(n12458), .ZN(
        n12442) );
  INV_X1 U12077 ( .A(n14704), .ZN(n10219) );
  OAI211_X1 U12078 ( .C1(n10921), .C2(n10045), .A(n10077), .B(n11504), .ZN(
        n11514) );
  NAND2_X1 U12079 ( .A1(n10078), .A2(n14561), .ZN(n10077) );
  AOI21_X1 U12080 ( .B1(n15157), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A(
        n10066), .ZN(n15198) );
  AND2_X1 U12081 ( .A1(n9717), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10066) );
  AOI22_X1 U12082 ( .A1(n9727), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(n9717), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15202) );
  INV_X1 U12083 ( .A(n13344), .ZN(n10597) );
  OAI22_X1 U12084 ( .A1(n20551), .A2(n12334), .B1(n12970), .B2(n9934), .ZN(
        n12335) );
  AOI21_X1 U12085 ( .B1(n12207), .B2(n12590), .A(n12594), .ZN(n10199) );
  NAND2_X1 U12086 ( .A1(n12219), .A2(n12579), .ZN(n10200) );
  AOI22_X1 U12087 ( .A1(n9727), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9736), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12124) );
  AOI21_X1 U12088 ( .B1(n12900), .B2(n12600), .A(n10206), .ZN(n12603) );
  NOR2_X1 U12089 ( .A1(n14331), .A2(n12600), .ZN(n12210) );
  CLKBUF_X2 U12090 ( .A(n10892), .Z(n11435) );
  OR2_X1 U12091 ( .A1(n11021), .A2(n11020), .ZN(n11750) );
  OR2_X1 U12092 ( .A1(n11009), .A2(n11008), .ZN(n11740) );
  NAND2_X1 U12093 ( .A1(n10180), .A2(n9935), .ZN(n11031) );
  INV_X1 U12094 ( .A(n11030), .ZN(n9935) );
  OR2_X1 U12095 ( .A1(n10931), .A2(n10930), .ZN(n11700) );
  NOR2_X1 U12096 ( .A1(n10852), .A2(n10851), .ZN(n11711) );
  AOI21_X1 U12097 ( .B1(n9732), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A(n10409), .ZN(n15303) );
  AND2_X1 U12098 ( .A1(n9717), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10409) );
  AOI21_X1 U12099 ( .B1(n15158), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A(
        n10068), .ZN(n15267) );
  AND2_X1 U12100 ( .A1(n9717), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10068) );
  NAND2_X1 U12101 ( .A1(n9717), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n15257) );
  NAND2_X1 U12102 ( .A1(n9717), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n15244) );
  NAND2_X1 U12103 ( .A1(n9717), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n15238) );
  NAND2_X1 U12104 ( .A1(n9717), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n15224) );
  NAND2_X1 U12105 ( .A1(n9717), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n15218) );
  NAND2_X1 U12106 ( .A1(n9717), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n15164) );
  NAND2_X1 U12107 ( .A1(n9717), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n15156) );
  AOI22_X1 U12108 ( .A1(n9719), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9721), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12135) );
  INV_X1 U12109 ( .A(n13353), .ZN(n10394) );
  NOR2_X1 U12110 ( .A1(n10185), .A2(n10596), .ZN(n10384) );
  AND2_X1 U12111 ( .A1(n12471), .A2(n9884), .ZN(n10366) );
  NOR2_X1 U12112 ( .A1(n10337), .A2(n10368), .ZN(n10367) );
  INV_X1 U12113 ( .A(n12503), .ZN(n10368) );
  NAND2_X1 U12114 ( .A1(n12318), .A2(n15209), .ZN(n10401) );
  AND2_X1 U12115 ( .A1(n16421), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10076) );
  OAI21_X1 U12116 ( .B1(n12227), .B2(n14087), .A(n9790), .ZN(n10074) );
  INV_X1 U12117 ( .A(n12898), .ZN(n12215) );
  NAND2_X1 U12118 ( .A1(n12603), .A2(n12606), .ZN(n13146) );
  INV_X1 U12119 ( .A(n15275), .ZN(n15251) );
  NAND2_X1 U12120 ( .A1(n12898), .A2(n14331), .ZN(n12202) );
  INV_X1 U12121 ( .A(n12275), .ZN(n10122) );
  NAND2_X1 U12122 ( .A1(n15157), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n10026) );
  NAND2_X1 U12123 ( .A1(n15157), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n9998) );
  NAND2_X1 U12124 ( .A1(n9721), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n10129) );
  NAND3_X1 U12125 ( .A1(n12141), .A2(n12142), .A3(n10132), .ZN(n10131) );
  NAND2_X1 U12126 ( .A1(n10134), .A2(n12143), .ZN(n10133) );
  AOI22_X1 U12127 ( .A1(n9720), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(n9721), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12165) );
  NAND2_X1 U12128 ( .A1(n13147), .A2(n10124), .ZN(n12607) );
  AND2_X1 U12129 ( .A1(n10125), .A2(n12606), .ZN(n10124) );
  NAND2_X1 U12130 ( .A1(n12548), .A2(n12547), .ZN(n12559) );
  XNOR2_X1 U12131 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12558) );
  INV_X1 U12132 ( .A(n12549), .ZN(n12552) );
  AND2_X1 U12133 ( .A1(n13787), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11914) );
  AND2_X1 U12134 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11907) );
  NOR2_X1 U12135 ( .A1(n14170), .A2(n14206), .ZN(n14168) );
  AND4_X1 U12136 ( .A1(n11971), .A2(n11970), .A3(n11969), .A4(n11968), .ZN(
        n11984) );
  AND4_X1 U12137 ( .A1(n12012), .A2(n12011), .A3(n12010), .A4(n12009), .ZN(
        n12024) );
  NAND2_X1 U12138 ( .A1(n10657), .A2(n10622), .ZN(n10621) );
  INV_X1 U12139 ( .A(n15550), .ZN(n10622) );
  NOR2_X1 U12140 ( .A1(n15808), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10421) );
  INV_X1 U12141 ( .A(n15494), .ZN(n10547) );
  NOR2_X1 U12142 ( .A1(n10549), .A2(n15507), .ZN(n10548) );
  INV_X1 U12143 ( .A(n15527), .ZN(n10549) );
  INV_X1 U12144 ( .A(n10358), .ZN(n9966) );
  INV_X1 U12145 ( .A(n16003), .ZN(n10361) );
  OAI21_X1 U12146 ( .B1(n18044), .B2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10360) );
  NAND2_X1 U12147 ( .A1(n14507), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10177) );
  INV_X1 U12148 ( .A(n10179), .ZN(n10178) );
  OR2_X1 U12149 ( .A1(n11799), .A2(n21733), .ZN(n10921) );
  INV_X1 U12150 ( .A(n10921), .ZN(n10906) );
  OR2_X1 U12151 ( .A1(n10869), .A2(n10868), .ZN(n11717) );
  NOR2_X1 U12152 ( .A1(n10912), .A2(n10911), .ZN(n10913) );
  AND2_X2 U12153 ( .A1(n10706), .A2(n13805), .ZN(n10892) );
  OR2_X1 U12154 ( .A1(n11548), .A2(n11547), .ZN(n11551) );
  AOI21_X1 U12155 ( .B1(n10082), .B2(n10083), .A(n9817), .ZN(n10080) );
  NAND2_X1 U12156 ( .A1(n11524), .A2(n10082), .ZN(n10081) );
  INV_X1 U12157 ( .A(n11564), .ZN(n11554) );
  AOI22_X1 U12158 ( .A1(n11544), .A2(n11543), .B1(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n21733), .ZN(n11545) );
  NOR2_X1 U12159 ( .A1(n11542), .A2(n11541), .ZN(n11543) );
  AND2_X1 U12160 ( .A1(n11805), .A2(n14591), .ZN(n10558) );
  AOI22_X1 U12161 ( .A1(n9719), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n9730), .ZN(n12184) );
  NOR2_X1 U12162 ( .A1(n16972), .A2(n10488), .ZN(n10487) );
  AND2_X1 U12163 ( .A1(n12632), .A2(n12730), .ZN(n10513) );
  AND2_X1 U12164 ( .A1(n10509), .A2(n12628), .ZN(n10507) );
  AND2_X1 U12165 ( .A1(n16646), .A2(n10510), .ZN(n10509) );
  MUX2_X1 U12166 ( .A(P2_EBX_REG_3__SCAN_IN), .B(n12623), .S(n9987), .Z(n12657) );
  NAND2_X1 U12167 ( .A1(n9725), .A2(n16707), .ZN(n12621) );
  NOR2_X1 U12168 ( .A1(n10521), .A2(n10520), .ZN(n10519) );
  INV_X1 U12169 ( .A(n16570), .ZN(n10520) );
  NAND2_X1 U12170 ( .A1(n12844), .A2(n10522), .ZN(n10521) );
  INV_X1 U12171 ( .A(n16585), .ZN(n10522) );
  NAND2_X1 U12172 ( .A1(n9720), .A2(n12129), .ZN(n15181) );
  NAND2_X1 U12173 ( .A1(n9717), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n15283) );
  NAND2_X1 U12174 ( .A1(n9717), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n15289) );
  INV_X1 U12175 ( .A(n10653), .ZN(n10652) );
  OR2_X1 U12176 ( .A1(n10654), .A2(n16804), .ZN(n10653) );
  NAND2_X1 U12177 ( .A1(n10655), .A2(n16808), .ZN(n10654) );
  INV_X1 U12178 ( .A(n16811), .ZN(n10655) );
  AND2_X1 U12179 ( .A1(n12987), .A2(n10584), .ZN(n10583) );
  INV_X1 U12180 ( .A(n14603), .ZN(n10584) );
  INV_X1 U12181 ( .A(n14624), .ZN(n10578) );
  AOI22_X1 U12182 ( .A1(n9720), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9721), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12154) );
  INV_X1 U12183 ( .A(n12150), .ZN(n12151) );
  AOI22_X1 U12184 ( .A1(n12311), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9723), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12150) );
  NOR2_X1 U12185 ( .A1(n13301), .A2(n17030), .ZN(n13300) );
  NOR2_X1 U12186 ( .A1(n13292), .A2(n17049), .ZN(n10489) );
  INV_X1 U12187 ( .A(n16822), .ZN(n12844) );
  NAND2_X1 U12188 ( .A1(n13277), .A2(n10499), .ZN(n13282) );
  NAND2_X1 U12189 ( .A1(n13277), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13280) );
  AND2_X1 U12190 ( .A1(n14884), .A2(n12829), .ZN(n10518) );
  INV_X1 U12191 ( .A(n16627), .ZN(n12829) );
  AND2_X1 U12192 ( .A1(n13178), .A2(n13207), .ZN(n10526) );
  INV_X1 U12193 ( .A(n12542), .ZN(n12543) );
  INV_X1 U12194 ( .A(n13170), .ZN(n10283) );
  AND2_X1 U12195 ( .A1(n10039), .A2(n10038), .ZN(n10037) );
  INV_X1 U12196 ( .A(n16467), .ZN(n10038) );
  NAND2_X1 U12197 ( .A1(n12776), .A2(n10531), .ZN(n10064) );
  NOR2_X1 U12198 ( .A1(n16445), .A2(n12627), .ZN(n13201) );
  NOR2_X1 U12199 ( .A1(n17267), .A2(n17266), .ZN(n10554) );
  NAND2_X1 U12200 ( .A1(n9977), .A2(n17037), .ZN(n9976) );
  NAND2_X1 U12201 ( .A1(n17040), .A2(n17038), .ZN(n10373) );
  INV_X1 U12202 ( .A(n16499), .ZN(n10523) );
  AND2_X1 U12203 ( .A1(n13356), .A2(n9831), .ZN(n10069) );
  NOR2_X1 U12204 ( .A1(n16509), .A2(n10525), .ZN(n10524) );
  INV_X1 U12205 ( .A(n13373), .ZN(n10525) );
  INV_X1 U12206 ( .A(n13366), .ZN(n10587) );
  NOR2_X1 U12207 ( .A1(n17088), .A2(n10396), .ZN(n10395) );
  INV_X1 U12208 ( .A(n13351), .ZN(n10396) );
  NOR2_X1 U12209 ( .A1(n13345), .A2(n10422), .ZN(n10599) );
  NOR2_X1 U12210 ( .A1(n17388), .A2(n17456), .ZN(n10398) );
  XNOR2_X1 U12211 ( .A(n10403), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10611) );
  NOR2_X1 U12212 ( .A1(n12542), .A2(n12627), .ZN(n10403) );
  NAND2_X1 U12213 ( .A1(n17221), .A2(n17225), .ZN(n10023) );
  NAND2_X1 U12214 ( .A1(n12514), .A2(n12506), .ZN(n12508) );
  AND2_X1 U12215 ( .A1(n10515), .A2(n14499), .ZN(n10514) );
  INV_X1 U12216 ( .A(n20337), .ZN(n10530) );
  INV_X1 U12217 ( .A(n16695), .ZN(n10241) );
  OAI21_X1 U12218 ( .B1(n12690), .B2(n12676), .A(n10239), .ZN(n10238) );
  INV_X1 U12219 ( .A(n9863), .ZN(n10244) );
  OAI21_X1 U12220 ( .B1(n12690), .B2(n9863), .A(n10237), .ZN(n10236) );
  NAND2_X1 U12221 ( .A1(n12690), .A2(n12677), .ZN(n10237) );
  NAND2_X1 U12222 ( .A1(n13974), .A2(n13973), .ZN(n13976) );
  INV_X1 U12223 ( .A(n14727), .ZN(n14687) );
  OR2_X1 U12224 ( .A1(n15251), .A2(n17573), .ZN(n14001) );
  NAND2_X1 U12225 ( .A1(n10203), .A2(n10202), .ZN(n12575) );
  NAND2_X1 U12226 ( .A1(n14742), .A2(n17596), .ZN(n10202) );
  NAND2_X1 U12227 ( .A1(n12573), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10203) );
  AND2_X1 U12228 ( .A1(n12211), .A2(n12905), .ZN(n10163) );
  NAND2_X1 U12229 ( .A1(n12200), .A2(n12129), .ZN(n9943) );
  NAND2_X1 U12230 ( .A1(n12199), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9942) );
  INV_X1 U12231 ( .A(n19028), .ZN(n10448) );
  INV_X1 U12232 ( .A(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17641) );
  NAND2_X1 U12233 ( .A1(n14019), .A2(n11915), .ZN(n11972) );
  AND2_X1 U12234 ( .A1(n14054), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11915) );
  NOR2_X1 U12235 ( .A1(n13965), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10432) );
  AND2_X1 U12236 ( .A1(n11914), .A2(n14019), .ZN(n14099) );
  AND2_X1 U12237 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11908) );
  CLKBUF_X3 U12238 ( .A(n14099), .Z(n18760) );
  AND4_X1 U12239 ( .A1(n14132), .A2(n14131), .A3(n14130), .A4(n14129), .ZN(
        n14146) );
  AND4_X1 U12240 ( .A1(n13917), .A2(n13916), .A3(n13915), .A4(n13914), .ZN(
        n13927) );
  INV_X1 U12241 ( .A(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n18753) );
  NAND2_X1 U12242 ( .A1(n18235), .A2(n13673), .ZN(n13777) );
  NAND2_X1 U12244 ( .A1(n10439), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10438) );
  INV_X1 U12245 ( .A(n10440), .ZN(n10439) );
  OR2_X1 U12246 ( .A1(n10441), .A2(n19054), .ZN(n10440) );
  NAND2_X1 U12247 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10441) );
  NAND2_X1 U12248 ( .A1(n17844), .A2(n9812), .ZN(n10014) );
  AND2_X1 U12249 ( .A1(n19213), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11891) );
  NOR2_X1 U12250 ( .A1(n14207), .A2(n14206), .ZN(n14209) );
  AND4_X1 U12251 ( .A1(n12053), .A2(n12052), .A3(n12051), .A4(n12050), .ZN(
        n12068) );
  NAND2_X1 U12252 ( .A1(n19070), .A2(n10329), .ZN(n17765) );
  NAND2_X1 U12253 ( .A1(n10327), .A2(n10324), .ZN(n10329) );
  NAND2_X1 U12254 ( .A1(n10328), .A2(n17762), .ZN(n10327) );
  AND2_X1 U12255 ( .A1(n19073), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10316) );
  NAND2_X1 U12256 ( .A1(n17756), .A2(n17844), .ZN(n17761) );
  OR2_X1 U12257 ( .A1(n14218), .A2(n17755), .ZN(n14219) );
  AND4_X1 U12258 ( .A1(n14150), .A2(n14149), .A3(n14148), .A4(n14147), .ZN(
        n14165) );
  NAND2_X1 U12259 ( .A1(n19276), .A2(n14217), .ZN(n14223) );
  NAND2_X1 U12260 ( .A1(n14200), .A2(n10424), .ZN(n10320) );
  AND2_X1 U12261 ( .A1(n12089), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13681) );
  NOR2_X1 U12262 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14028) );
  NAND2_X1 U12263 ( .A1(n19650), .A2(n12079), .ZN(n13771) );
  AOI21_X1 U12264 ( .B1(n19615), .B2(n20116), .A(n20095), .ZN(n19625) );
  NAND2_X1 U12265 ( .A1(n13569), .A2(n10559), .ZN(n13571) );
  AND2_X1 U12266 ( .A1(n10796), .A2(n11805), .ZN(n10560) );
  AND2_X1 U12267 ( .A1(n11556), .A2(n11558), .ZN(n13575) );
  OR2_X1 U12268 ( .A1(n21200), .A2(n11673), .ZN(n21203) );
  INV_X1 U12269 ( .A(n13562), .ZN(n15651) );
  AND2_X1 U12270 ( .A1(n11611), .A2(n11610), .ZN(n15616) );
  NOR2_X1 U12271 ( .A1(n14875), .A2(n10543), .ZN(n15617) );
  AND2_X1 U12272 ( .A1(n11592), .A2(n11591), .ZN(n14839) );
  AND2_X1 U12273 ( .A1(n11654), .A2(n9734), .ZN(n14008) );
  INV_X1 U12274 ( .A(n15020), .ZN(n14547) );
  NOR2_X1 U12275 ( .A1(n11451), .A2(n15805), .ZN(n11452) );
  OR2_X1 U12276 ( .A1(n15800), .A2(n11455), .ZN(n11475) );
  AOI21_X1 U12277 ( .B1(n15807), .B2(n11278), .A(n11450), .ZN(n15392) );
  NAND2_X1 U12278 ( .A1(n11431), .A2(n11430), .ZN(n15407) );
  OR2_X1 U12279 ( .A1(n15831), .A2(n11455), .ZN(n11408) );
  NAND2_X1 U12280 ( .A1(n15442), .A2(n10634), .ZN(n15406) );
  OR2_X1 U12281 ( .A1(n11370), .A2(n11369), .ZN(n11389) );
  AOI21_X1 U12282 ( .B1(n15852), .B2(n11161), .A(n11368), .ZN(n15443) );
  OR2_X1 U12283 ( .A1(n15854), .A2(n11455), .ZN(n11351) );
  AND2_X1 U12284 ( .A1(n11320), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11321) );
  NAND2_X1 U12285 ( .A1(n11321), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11370) );
  NAND2_X1 U12286 ( .A1(n11317), .A2(n11316), .ZN(n15470) );
  AND2_X1 U12287 ( .A1(n11280), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11281) );
  INV_X1 U12288 ( .A(n11279), .ZN(n11280) );
  OR2_X1 U12289 ( .A1(n15874), .A2(n11455), .ZN(n11299) );
  AND2_X1 U12290 ( .A1(n11242), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11243) );
  NAND2_X1 U12291 ( .A1(n11262), .A2(n11261), .ZN(n15505) );
  OR2_X1 U12292 ( .A1(n15892), .A2(n11455), .ZN(n11262) );
  NAND2_X1 U12293 ( .A1(n11240), .A2(n11239), .ZN(n15504) );
  NAND2_X1 U12294 ( .A1(n11207), .A2(n11206), .ZN(n11241) );
  AND2_X1 U12295 ( .A1(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11206) );
  INV_X1 U12296 ( .A(n11205), .ZN(n11207) );
  INV_X1 U12297 ( .A(n14879), .ZN(n10620) );
  OR2_X1 U12298 ( .A1(n11177), .A2(n11135), .ZN(n11200) );
  NAND2_X1 U12299 ( .A1(n11101), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11177) );
  OR2_X1 U12300 ( .A1(n11093), .A2(n21130), .ZN(n11100) );
  AND2_X1 U12301 ( .A1(n11098), .A2(n11097), .ZN(n14880) );
  NAND2_X1 U12302 ( .A1(n11077), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11093) );
  AND3_X1 U12303 ( .A1(n11066), .A2(n11065), .A3(n11064), .ZN(n14819) );
  AND3_X1 U12304 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A3(n11046), .ZN(n11077) );
  CLKBUF_X1 U12305 ( .A(n14513), .Z(n14601) );
  NAND2_X1 U12306 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10960) );
  NOR2_X1 U12307 ( .A1(n10960), .A2(n21202), .ZN(n10961) );
  NAND2_X1 U12308 ( .A1(n15416), .A2(n9763), .ZN(n15378) );
  NAND2_X1 U12309 ( .A1(n15979), .A2(n16050), .ZN(n10182) );
  NAND2_X1 U12310 ( .A1(n15416), .A2(n10538), .ZN(n15405) );
  OAI21_X1 U12311 ( .B1(n15898), .B2(n10300), .A(n10299), .ZN(n10301) );
  INV_X1 U12312 ( .A(n10566), .ZN(n10300) );
  NOR2_X1 U12313 ( .A1(n15857), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15835) );
  NOR2_X1 U12314 ( .A1(n16252), .A2(n11830), .ZN(n10097) );
  NAND2_X1 U12315 ( .A1(n15526), .A2(n9868), .ZN(n15496) );
  NAND2_X1 U12316 ( .A1(n15526), .A2(n10548), .ZN(n15508) );
  NAND2_X1 U12317 ( .A1(n10094), .A2(n10091), .ZN(n16125) );
  INV_X1 U12318 ( .A(n10097), .ZN(n10094) );
  NOR2_X1 U12319 ( .A1(n10090), .A2(n10093), .ZN(n10091) );
  AND2_X1 U12320 ( .A1(n11627), .A2(n11626), .ZN(n15539) );
  AND2_X1 U12321 ( .A1(n11623), .A2(n11622), .ZN(n15551) );
  NOR2_X2 U12322 ( .A1(n15571), .A2(n15551), .ZN(n15553) );
  XNOR2_X1 U12323 ( .A(n15993), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15920) );
  NAND2_X1 U12324 ( .A1(n10293), .A2(n10292), .ZN(n15917) );
  INV_X1 U12325 ( .A(n15931), .ZN(n10294) );
  NAND2_X1 U12326 ( .A1(n10541), .A2(n15599), .ZN(n10540) );
  INV_X1 U12327 ( .A(n10543), .ZN(n10541) );
  NOR2_X1 U12328 ( .A1(n15959), .A2(n11766), .ZN(n15941) );
  NAND2_X1 U12329 ( .A1(n10542), .A2(n10674), .ZN(n15633) );
  INV_X1 U12330 ( .A(n14875), .ZN(n10542) );
  NOR2_X1 U12331 ( .A1(n15993), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10173) );
  INV_X1 U12332 ( .A(n10172), .ZN(n10174) );
  AND2_X1 U12333 ( .A1(n11760), .A2(n9876), .ZN(n10563) );
  NOR2_X1 U12334 ( .A1(n14521), .A2(n10536), .ZN(n14841) );
  NAND2_X1 U12335 ( .A1(n14072), .A2(n14071), .ZN(n10555) );
  NAND2_X1 U12336 ( .A1(n10533), .A2(n14452), .ZN(n10532) );
  INV_X1 U12337 ( .A(n14074), .ZN(n10533) );
  NAND2_X1 U12338 ( .A1(n18087), .A2(n21733), .ZN(n11686) );
  OR2_X1 U12339 ( .A1(n11824), .A2(n11818), .ZN(n14013) );
  OAI211_X1 U12340 ( .C1(n11541), .C2(n10903), .A(n10902), .B(n10901), .ZN(
        n10986) );
  CLKBUF_X1 U12341 ( .A(n14392), .Z(n21305) );
  NAND2_X1 U12342 ( .A1(n10952), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11682) );
  INV_X1 U12343 ( .A(n10838), .ZN(n10348) );
  NAND2_X1 U12344 ( .A1(n10858), .A2(n10838), .ZN(n10347) );
  OR3_X1 U12345 ( .A1(n13799), .A2(n13798), .A3(n13797), .ZN(n17997) );
  NAND2_X1 U12346 ( .A1(n21305), .A2(n21304), .ZN(n21413) );
  OR2_X1 U12347 ( .A1(n9707), .A2(n16317), .ZN(n21454) );
  INV_X1 U12348 ( .A(n10765), .ZN(n10768) );
  INV_X1 U12349 ( .A(n10766), .ZN(n10767) );
  NAND2_X1 U12350 ( .A1(n9707), .A2(n14752), .ZN(n21369) );
  NOR2_X1 U12351 ( .A1(n15020), .A2(n18057), .ZN(n14582) );
  INV_X1 U12352 ( .A(n14584), .ZN(n14576) );
  AND2_X1 U12353 ( .A1(n15370), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n18034) );
  OR2_X1 U12354 ( .A1(n17992), .A2(n18039), .ZN(n18025) );
  INV_X1 U12355 ( .A(n14854), .ZN(n14731) );
  NAND2_X1 U12356 ( .A1(n12571), .A2(n12570), .ZN(n12597) );
  NAND2_X1 U12357 ( .A1(n16430), .A2(n16736), .ZN(n10495) );
  NOR2_X1 U12358 ( .A1(n13295), .A2(n10490), .ZN(n10161) );
  NAND2_X1 U12359 ( .A1(n17043), .A2(n10491), .ZN(n10490) );
  INV_X1 U12360 ( .A(n17053), .ZN(n10491) );
  NOR2_X1 U12361 ( .A1(n16544), .A2(n17053), .ZN(n16517) );
  AND2_X1 U12362 ( .A1(n20350), .A2(n13295), .ZN(n16544) );
  AND2_X1 U12363 ( .A1(n13102), .A2(n13101), .ZN(n16533) );
  NOR2_X1 U12364 ( .A1(n16559), .A2(n10150), .ZN(n20266) );
  NOR2_X1 U12365 ( .A1(n20283), .A2(n13286), .ZN(n16577) );
  AND2_X1 U12366 ( .A1(n13277), .A2(n9751), .ZN(n13285) );
  AND2_X1 U12367 ( .A1(n12730), .A2(n16606), .ZN(n10061) );
  NOR2_X1 U12368 ( .A1(n16635), .A2(n16633), .ZN(n16619) );
  NOR2_X1 U12369 ( .A1(n12696), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12728) );
  NAND2_X1 U12370 ( .A1(n20310), .A2(n13270), .ZN(n20313) );
  AND2_X1 U12371 ( .A1(n16655), .A2(n17200), .ZN(n20310) );
  NOR2_X1 U12372 ( .A1(n12675), .A2(n12674), .ZN(n12688) );
  INV_X1 U12373 ( .A(n20354), .ZN(n10151) );
  NOR2_X1 U12374 ( .A1(n16722), .A2(n16715), .ZN(n16697) );
  OR2_X1 U12375 ( .A1(n14732), .A2(n18142), .ZN(n13461) );
  NOR2_X1 U12376 ( .A1(n14646), .A2(n10521), .ZN(n16586) );
  AOI21_X1 U12377 ( .B1(n9731), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A(
        n10067), .ZN(n15318) );
  AND2_X1 U12378 ( .A1(n9717), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10067) );
  AOI21_X1 U12379 ( .B1(n12310), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n10065), .ZN(n15330) );
  NAND2_X1 U12380 ( .A1(n16451), .A2(n10580), .ZN(n13132) );
  AND2_X1 U12381 ( .A1(n9764), .A2(n13180), .ZN(n10580) );
  NAND2_X1 U12382 ( .A1(n10645), .A2(n10642), .ZN(n16747) );
  NAND2_X1 U12383 ( .A1(n15296), .A2(n10647), .ZN(n10645) );
  NOR2_X1 U12384 ( .A1(n16748), .A2(n10648), .ZN(n10647) );
  AND2_X1 U12385 ( .A1(n13123), .A2(n13122), .ZN(n13210) );
  NAND2_X1 U12386 ( .A1(n16451), .A2(n9761), .ZN(n16439) );
  XNOR2_X1 U12387 ( .A(n15235), .B(n15232), .ZN(n16770) );
  NAND2_X1 U12388 ( .A1(n16770), .A2(n16769), .ZN(n16768) );
  NAND2_X1 U12389 ( .A1(n15063), .A2(n9746), .ZN(n16797) );
  INV_X1 U12390 ( .A(n16532), .ZN(n16929) );
  OR2_X1 U12391 ( .A1(n16816), .A2(n10654), .ZN(n16807) );
  INV_X1 U12392 ( .A(n16571), .ZN(n10588) );
  NAND2_X1 U12393 ( .A1(n15063), .A2(n15062), .ZN(n16816) );
  AND2_X1 U12394 ( .A1(n13094), .A2(n13093), .ZN(n16591) );
  NAND2_X1 U12395 ( .A1(n14619), .A2(n10589), .ZN(n16589) );
  AND2_X1 U12396 ( .A1(n14619), .A2(n14807), .ZN(n14806) );
  AND3_X1 U12397 ( .A1(n13056), .A2(n13055), .A3(n13054), .ZN(n14620) );
  AND3_X1 U12398 ( .A1(n13038), .A2(n13037), .A3(n13036), .ZN(n14639) );
  AND3_X1 U12399 ( .A1(n12986), .A2(n12985), .A3(n12984), .ZN(n14631) );
  OR2_X1 U12400 ( .A1(n16938), .A2(n14427), .ZN(n16946) );
  NAND2_X1 U12401 ( .A1(n12203), .A2(n10363), .ZN(n14422) );
  AND2_X1 U12402 ( .A1(n10206), .A2(n14866), .ZN(n10363) );
  INV_X1 U12403 ( .A(n10406), .ZN(n14421) );
  NAND2_X1 U12404 ( .A1(n12897), .A2(n12896), .ZN(n14418) );
  AOI22_X1 U12405 ( .A1(n12899), .A2(n12895), .B1(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n13145), .ZN(n12896) );
  OAI211_X1 U12406 ( .C1(n12942), .C2(n12904), .A(n12903), .B(n12916), .ZN(
        n14419) );
  INV_X1 U12407 ( .A(n13479), .ZN(n13550) );
  NAND2_X1 U12408 ( .A1(n10486), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10481) );
  NAND2_X1 U12409 ( .A1(n13312), .A2(n10483), .ZN(n10482) );
  OR2_X1 U12410 ( .A1(n13312), .A2(n13233), .ZN(n10484) );
  NAND2_X1 U12411 ( .A1(n10489), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13301) );
  INV_X1 U12412 ( .A(n10489), .ZN(n13298) );
  AND2_X1 U12413 ( .A1(n9751), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10498) );
  NOR2_X1 U12414 ( .A1(n17097), .A2(n10246), .ZN(n10245) );
  INV_X1 U12415 ( .A(n10248), .ZN(n10246) );
  NAND2_X1 U12416 ( .A1(n10036), .A2(n12844), .ZN(n16824) );
  INV_X1 U12417 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17172) );
  AND2_X1 U12418 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n13230) );
  INV_X1 U12419 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20340) );
  NOR2_X1 U12420 ( .A1(n9739), .A2(n13160), .ZN(n10167) );
  OR2_X1 U12421 ( .A1(n17278), .A2(n13172), .ZN(n13402) );
  INV_X1 U12422 ( .A(n12784), .ZN(n10417) );
  INV_X1 U12423 ( .A(n13188), .ZN(n10416) );
  NAND2_X1 U12424 ( .A1(n10110), .A2(n10108), .ZN(n10413) );
  NOR2_X1 U12425 ( .A1(n10418), .A2(n10109), .ZN(n10108) );
  INV_X1 U12426 ( .A(n10111), .ZN(n10109) );
  NAND2_X1 U12427 ( .A1(n16451), .A2(n16452), .ZN(n16438) );
  NOR2_X1 U12428 ( .A1(n17481), .A2(n9894), .ZN(n13161) );
  INV_X1 U12429 ( .A(n13159), .ZN(n10195) );
  AND2_X1 U12430 ( .A1(n13371), .A2(n9798), .ZN(n16498) );
  INV_X1 U12431 ( .A(n10609), .ZN(n10604) );
  INV_X1 U12432 ( .A(n10606), .ZN(n10605) );
  OR2_X1 U12433 ( .A1(n20264), .A2(n12760), .ZN(n17066) );
  AND2_X1 U12434 ( .A1(n18126), .A2(n17365), .ZN(n10032) );
  AND2_X1 U12435 ( .A1(n10042), .A2(n14834), .ZN(n10041) );
  NAND2_X1 U12436 ( .A1(n17364), .A2(n17381), .ZN(n17118) );
  NAND2_X1 U12437 ( .A1(n9972), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12540) );
  INV_X1 U12438 ( .A(n17206), .ZN(n9972) );
  INV_X1 U12439 ( .A(n10611), .ZN(n17193) );
  CLKBUF_X1 U12440 ( .A(n17204), .Z(n17205) );
  NOR2_X1 U12441 ( .A1(n17517), .A2(n13158), .ZN(n13162) );
  NAND2_X1 U12442 ( .A1(n17219), .A2(n17220), .ZN(n12684) );
  NAND2_X1 U12443 ( .A1(n9984), .A2(n12425), .ZN(n12513) );
  NAND2_X1 U12444 ( .A1(n9945), .A2(n12262), .ZN(n9944) );
  AND2_X1 U12445 ( .A1(n10205), .A2(n10204), .ZN(n17524) );
  AOI21_X1 U12446 ( .B1(n17361), .B2(n13157), .A(n13156), .ZN(n10204) );
  INV_X1 U12447 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13584) );
  AND2_X1 U12448 ( .A1(n12931), .A2(n12930), .ZN(n16689) );
  NAND2_X1 U12449 ( .A1(n10125), .A2(n14866), .ZN(n13153) );
  INV_X1 U12450 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n21861) );
  AND2_X1 U12451 ( .A1(n21058), .A2(n21072), .ZN(n21043) );
  INV_X1 U12452 ( .A(n21043), .ZN(n20752) );
  INV_X1 U12453 ( .A(n21062), .ZN(n20835) );
  NOR2_X2 U12454 ( .A1(n15337), .A2(n14862), .ZN(n20453) );
  NOR2_X2 U12455 ( .A1(n15338), .A2(n14862), .ZN(n20454) );
  NAND2_X1 U12456 ( .A1(n9719), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n10139) );
  INV_X1 U12457 ( .A(n20896), .ZN(n20623) );
  NOR2_X1 U12458 ( .A1(n20713), .A2(n20712), .ZN(n20894) );
  OAI21_X1 U12459 ( .B1(n12582), .B2(n12580), .A(n12597), .ZN(n14732) );
  AND2_X1 U12460 ( .A1(n19628), .A2(n18973), .ZN(n13673) );
  NOR2_X1 U12461 ( .A1(n14038), .A2(n12087), .ZN(n20061) );
  AND2_X1 U12462 ( .A1(n10445), .A2(n9888), .ZN(n18272) );
  NAND2_X1 U12463 ( .A1(n10450), .A2(n10448), .ZN(n10446) );
  NAND2_X1 U12464 ( .A1(n10448), .A2(n19040), .ZN(n10447) );
  NOR2_X1 U12465 ( .A1(n18292), .A2(n18293), .ZN(n18291) );
  NOR2_X1 U12466 ( .A1(n19058), .A2(n18300), .ZN(n18299) );
  NAND2_X1 U12468 ( .A1(n18349), .A2(n21897), .ZN(n18343) );
  NOR2_X1 U12469 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n18365), .ZN(n18349) );
  NAND2_X1 U12470 ( .A1(n18392), .A2(n18386), .ZN(n18381) );
  NOR2_X1 U12471 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n18414), .ZN(n18392) );
  NOR2_X1 U12472 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n18460), .ZN(n18445) );
  NOR2_X1 U12474 ( .A1(n10461), .A2(n21845), .ZN(n10460) );
  INV_X1 U12475 ( .A(n10462), .ZN(n10461) );
  NOR2_X1 U12476 ( .A1(n21874), .A2(n10463), .ZN(n10462) );
  INV_X1 U12477 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n10463) );
  NOR2_X1 U12478 ( .A1(n22097), .A2(n18541), .ZN(n10480) );
  AND4_X1 U12479 ( .A1(n11946), .A2(n11945), .A3(n11944), .A4(n11943), .ZN(
        n11963) );
  INV_X1 U12480 ( .A(n10668), .ZN(n10469) );
  NAND2_X1 U12481 ( .A1(n9821), .A2(n9741), .ZN(n10470) );
  NOR2_X1 U12482 ( .A1(n18925), .A2(n10265), .ZN(n10264) );
  NOR2_X1 U12483 ( .A1(n18862), .A2(n10275), .ZN(n10274) );
  NAND2_X1 U12484 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(P3_EAX_REG_16__SCAN_IN), 
        .ZN(n10275) );
  INV_X1 U12485 ( .A(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17678) );
  AND2_X1 U12486 ( .A1(n13840), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13784) );
  NOR2_X1 U12487 ( .A1(n18953), .A2(n18901), .ZN(n17711) );
  OR2_X1 U12488 ( .A1(n10270), .A2(n13885), .ZN(n10269) );
  AND2_X1 U12489 ( .A1(n13840), .A2(n13965), .ZN(n14466) );
  AND4_X1 U12490 ( .A1(n13951), .A2(n13950), .A3(n13949), .A4(n13948), .ZN(
        n13960) );
  AND4_X1 U12491 ( .A1(n13903), .A2(n13902), .A3(n13901), .A4(n13900), .ZN(
        n13904) );
  AND4_X1 U12492 ( .A1(n13895), .A2(n13894), .A3(n13893), .A4(n13892), .ZN(
        n13906) );
  AND3_X1 U12493 ( .A1(n19646), .A2(n19642), .A3(n18606), .ZN(n13874) );
  AOI21_X1 U12494 ( .B1(n13777), .B2(n20098), .A(n20215), .ZN(n18915) );
  INV_X1 U12495 ( .A(n18971), .ZN(n18918) );
  CLKBUF_X1 U12496 ( .A(n11892), .Z(n11893) );
  CLKBUF_X1 U12497 ( .A(n11870), .Z(n11871) );
  AND2_X1 U12498 ( .A1(n17767), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n19024) );
  NAND2_X1 U12499 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n19178) );
  CLKBUF_X1 U12500 ( .A(n11889), .Z(n11890) );
  INV_X1 U12501 ( .A(n19313), .ZN(n19306) );
  AND2_X1 U12502 ( .A1(n17767), .A2(n9899), .ZN(n17770) );
  NOR2_X1 U12503 ( .A1(n17903), .A2(n19034), .ZN(n10430) );
  OAI21_X1 U12504 ( .B1(n10333), .B2(n10332), .A(n10330), .ZN(n17808) );
  NOR2_X1 U12505 ( .A1(n10332), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10331) );
  OR2_X1 U12506 ( .A1(n17768), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10332) );
  NAND2_X1 U12507 ( .A1(n17767), .A2(n9893), .ZN(n19027) );
  NAND2_X1 U12508 ( .A1(n10012), .A2(n19034), .ZN(n19026) );
  NAND2_X1 U12509 ( .A1(n10315), .A2(n10313), .ZN(n19355) );
  NOR2_X1 U12510 ( .A1(n9767), .A2(n10314), .ZN(n10313) );
  INV_X1 U12511 ( .A(n17901), .ZN(n10314) );
  AND2_X1 U12512 ( .A1(n9859), .A2(n10018), .ZN(n19045) );
  AOI21_X1 U12513 ( .B1(n17765), .B2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n10019), .ZN(n10018) );
  AND2_X1 U12514 ( .A1(n10323), .A2(n19050), .ZN(n10019) );
  NAND2_X1 U12515 ( .A1(n10315), .A2(n10316), .ZN(n19384) );
  NOR2_X1 U12516 ( .A1(n17760), .A2(n10427), .ZN(n10426) );
  AND2_X1 U12517 ( .A1(n10323), .A2(n10428), .ZN(n10427) );
  NAND2_X1 U12518 ( .A1(n17761), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10429) );
  NAND2_X1 U12519 ( .A1(n10017), .A2(n17761), .ZN(n19175) );
  INV_X1 U12520 ( .A(n17760), .ZN(n10017) );
  INV_X1 U12521 ( .A(n19408), .ZN(n19513) );
  NAND2_X1 U12522 ( .A1(n14225), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17856) );
  INV_X1 U12523 ( .A(n14225), .ZN(n10020) );
  AOI21_X1 U12524 ( .B1(n14400), .B2(n10303), .A(n9804), .ZN(n10302) );
  NAND2_X1 U12525 ( .A1(n14187), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14402) );
  INV_X1 U12526 ( .A(n14182), .ZN(n10304) );
  NAND2_X1 U12527 ( .A1(n10013), .A2(n14194), .ZN(n14201) );
  NAND2_X1 U12528 ( .A1(n19331), .A2(n14178), .ZN(n19316) );
  NAND2_X1 U12529 ( .A1(n13705), .A2(n13704), .ZN(n20064) );
  AND2_X1 U12530 ( .A1(n20062), .A2(n13684), .ZN(n20063) );
  AND3_X1 U12531 ( .A1(n13698), .A2(n13697), .A3(n13696), .ZN(n20059) );
  NAND2_X1 U12532 ( .A1(n10259), .A2(n10258), .ZN(n13677) );
  NOR2_X1 U12533 ( .A1(n13689), .A2(n10262), .ZN(n10258) );
  INV_X1 U12534 ( .A(n12085), .ZN(n10259) );
  NOR2_X2 U12535 ( .A1(n14031), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14026) );
  NAND2_X1 U12536 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13775) );
  NOR2_X1 U12537 ( .A1(n10261), .A2(n13677), .ZN(n14038) );
  NOR2_X1 U12538 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19625), .ZN(n19862) );
  INV_X1 U12539 ( .A(n19862), .ZN(n19912) );
  OR3_X1 U12540 ( .A1(n17992), .A2(n13564), .A3(n21099), .ZN(n15373) );
  AND2_X1 U12541 ( .A1(n11672), .A2(n11670), .ZN(n21210) );
  NAND2_X1 U12542 ( .A1(n11672), .A2(n11671), .ZN(n21205) );
  INV_X1 U12543 ( .A(n21217), .ZN(n21146) );
  NAND2_X2 U12544 ( .A1(n14068), .A2(n14067), .ZN(n15709) );
  OR2_X1 U12545 ( .A1(n14063), .A2(n21099), .ZN(n14068) );
  NAND2_X1 U12546 ( .A1(n15786), .A2(n14595), .ZN(n15768) );
  INV_X1 U12547 ( .A(n15776), .ZN(n15770) );
  OR2_X1 U12548 ( .A1(n14596), .A2(n14547), .ZN(n15776) );
  INV_X1 U12549 ( .A(n13423), .ZN(n15786) );
  AND2_X1 U12550 ( .A1(n15768), .A2(n14596), .ZN(n15788) );
  NOR2_X1 U12551 ( .A1(n18095), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n21234) );
  INV_X1 U12552 ( .A(n21256), .ZN(n21235) );
  INV_X1 U12553 ( .A(n21821), .ZN(n21254) );
  OAI21_X1 U12554 ( .B1(n15391), .B2(n15392), .A(n15380), .ZN(n15816) );
  INV_X1 U12555 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n21130) );
  INV_X1 U12556 ( .A(n18056), .ZN(n15997) );
  INV_X1 U12557 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18062) );
  INV_X1 U12558 ( .A(n18061), .ZN(n18048) );
  XNOR2_X1 U12559 ( .A(n10423), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11855) );
  NAND2_X1 U12560 ( .A1(n10149), .A2(n10148), .ZN(n10423) );
  NAND2_X1 U12561 ( .A1(n11860), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10148) );
  NOR2_X1 U12562 ( .A1(n16021), .A2(n10084), .ZN(n16012) );
  NAND2_X1 U12563 ( .A1(n10085), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10084) );
  NAND2_X1 U12564 ( .A1(n16257), .A2(n11838), .ZN(n10085) );
  AND2_X1 U12565 ( .A1(n9745), .A2(n10145), .ZN(n15795) );
  OR3_X1 U12566 ( .A1(n16079), .A2(n16050), .A3(n16049), .ZN(n16030) );
  NAND2_X1 U12567 ( .A1(n11837), .A2(n10086), .ZN(n16042) );
  NAND2_X1 U12568 ( .A1(n16061), .A2(n9909), .ZN(n10086) );
  NOR2_X1 U12569 ( .A1(n10096), .A2(n9820), .ZN(n10095) );
  INV_X1 U12570 ( .A(n11832), .ZN(n10096) );
  NAND2_X1 U12571 ( .A1(n10181), .A2(n15845), .ZN(n15846) );
  INV_X1 U12572 ( .A(n15857), .ZN(n10181) );
  OAI21_X1 U12573 ( .B1(n15898), .B2(n9901), .A(n15909), .ZN(n15861) );
  NAND2_X1 U12574 ( .A1(n10569), .A2(n15993), .ZN(n15862) );
  AND2_X1 U12575 ( .A1(n16092), .A2(n16091), .ZN(n16123) );
  AND2_X1 U12576 ( .A1(n16186), .A2(n21912), .ZN(n14247) );
  INV_X1 U12577 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21306) );
  INV_X1 U12578 ( .A(n10047), .ZN(n21304) );
  CLKBUF_X1 U12579 ( .A(n14349), .Z(n21310) );
  INV_X1 U12580 ( .A(n17992), .ZN(n13816) );
  NOR2_X1 U12581 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n18087) );
  INV_X1 U12582 ( .A(n21404), .ZN(n21372) );
  INV_X1 U12583 ( .A(n21362), .ZN(n21365) );
  OAI21_X1 U12584 ( .B1(n21378), .B2(n21382), .A(n21377), .ZN(n21407) );
  OAI221_X1 U12585 ( .B1(n10670), .B2(n11673), .C1(n10670), .C2(n21458), .A(
        n21457), .ZN(n21476) );
  OR2_X1 U12586 ( .A1(n21455), .A2(n21532), .ZN(n21510) );
  INV_X1 U12587 ( .A(n21501), .ZN(n21506) );
  INV_X1 U12588 ( .A(n21510), .ZN(n21498) );
  OAI211_X1 U12589 ( .C1(n21679), .C2(n16282), .A(n14545), .B(n21677), .ZN(
        n14581) );
  OAI21_X1 U12590 ( .B1(n16322), .B2(n21518), .A(n21568), .ZN(n21521) );
  INV_X1 U12591 ( .A(n21611), .ZN(n21633) );
  INV_X1 U12592 ( .A(n21653), .ZN(n21624) );
  INV_X1 U12593 ( .A(n21649), .ZN(n16370) );
  INV_X1 U12594 ( .A(n21714), .ZN(n21598) );
  INV_X1 U12595 ( .A(n21723), .ZN(n21602) );
  OAI211_X1 U12596 ( .C1(n14758), .C2(n21654), .A(n21566), .B(n21457), .ZN(
        n21656) );
  INV_X1 U12597 ( .A(n21639), .ZN(n21670) );
  INV_X1 U12598 ( .A(n21576), .ZN(n21684) );
  INV_X1 U12599 ( .A(n16382), .ZN(n21685) );
  AND2_X1 U12600 ( .A1(n14553), .A2(n14576), .ZN(n21696) );
  INV_X1 U12601 ( .A(n16391), .ZN(n21697) );
  INV_X1 U12602 ( .A(n21644), .ZN(n21702) );
  INV_X1 U12603 ( .A(n21731), .ZN(n21717) );
  AND2_X1 U12604 ( .A1(n10799), .A2(n14576), .ZN(n21714) );
  INV_X1 U12605 ( .A(n16405), .ZN(n21715) );
  INV_X1 U12606 ( .A(n21720), .ZN(n21727) );
  OR2_X1 U12607 ( .A1(n21673), .A2(n21410), .ZN(n21731) );
  INV_X1 U12608 ( .A(n16410), .ZN(n21724) );
  INV_X1 U12609 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n20965) );
  OAI21_X1 U12610 ( .B1(n15343), .B2(n20341), .A(n13339), .ZN(n13340) );
  AOI21_X1 U12611 ( .B1(n13338), .B2(n16736), .A(n13337), .ZN(n13339) );
  INV_X1 U12612 ( .A(n20339), .ZN(n20262) );
  NAND2_X1 U12613 ( .A1(n16423), .A2(n13330), .ZN(n20292) );
  OR2_X1 U12614 ( .A1(n16423), .A2(n13327), .ZN(n20336) );
  INV_X1 U12615 ( .A(n20351), .ZN(n20326) );
  NAND2_X1 U12616 ( .A1(n10153), .A2(n10152), .ZN(n20349) );
  NAND2_X1 U12617 ( .A1(n10160), .A2(n20326), .ZN(n16742) );
  MUX2_X1 U12618 ( .A(n13584), .B(n16741), .S(n17596), .Z(n16739) );
  OR2_X1 U12619 ( .A1(n13002), .A2(n13001), .ZN(n14887) );
  OR2_X1 U12620 ( .A1(n12963), .A2(n12962), .ZN(n14815) );
  INV_X1 U12621 ( .A(n21072), .ZN(n21045) );
  NAND2_X1 U12622 ( .A1(n15296), .A2(n16753), .ZN(n10646) );
  INV_X1 U12623 ( .A(n10637), .ZN(n16762) );
  OR2_X1 U12624 ( .A1(n15339), .A2(n15337), .ZN(n16921) );
  OR2_X1 U12625 ( .A1(n15339), .A2(n15338), .ZN(n16941) );
  INV_X1 U12626 ( .A(n16941), .ZN(n20361) );
  INV_X1 U12627 ( .A(n16921), .ZN(n20362) );
  INV_X1 U12628 ( .A(n16946), .ZN(n20360) );
  NAND2_X1 U12629 ( .A1(n14333), .A2(n14332), .ZN(n14437) );
  AND2_X1 U12630 ( .A1(n20389), .A2(n16934), .ZN(n16963) );
  OR2_X1 U12631 ( .A1(n16938), .A2(n14426), .ZN(n20389) );
  INV_X1 U12632 ( .A(n16934), .ZN(n20385) );
  AND2_X1 U12633 ( .A1(n13628), .A2(n14733), .ZN(n20417) );
  INV_X2 U12634 ( .A(n13711), .ZN(n20425) );
  INV_X1 U12635 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18113) );
  NAND2_X1 U12636 ( .A1(n20239), .A2(n13227), .ZN(n18112) );
  NAND2_X1 U12637 ( .A1(n10411), .A2(n10410), .ZN(n13246) );
  AND2_X1 U12638 ( .A1(n10339), .A2(n10164), .ZN(n13216) );
  NOR2_X1 U12639 ( .A1(n10166), .A2(n10338), .ZN(n10164) );
  NAND2_X1 U12640 ( .A1(n10167), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10166) );
  NAND2_X1 U12641 ( .A1(n10187), .A2(n10186), .ZN(n16999) );
  NAND2_X1 U12642 ( .A1(n16996), .A2(n17007), .ZN(n10186) );
  NAND2_X1 U12643 ( .A1(n13161), .A2(n10338), .ZN(n17291) );
  NOR2_X1 U12644 ( .A1(n17036), .A2(n17035), .ZN(n17034) );
  OAI211_X1 U12645 ( .C1(n17364), .C2(n13361), .A(n10279), .B(n10278), .ZN(
        n17337) );
  OR2_X1 U12646 ( .A1(n9772), .A2(n13361), .ZN(n10279) );
  NAND2_X1 U12647 ( .A1(n10608), .A2(n10606), .ZN(n17060) );
  AND2_X1 U12648 ( .A1(n21906), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10256) );
  NAND2_X1 U12649 ( .A1(n12704), .A2(n12703), .ZN(n17166) );
  NAND2_X1 U12650 ( .A1(n17364), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17449) );
  AND2_X1 U12651 ( .A1(n17492), .A2(n17493), .ZN(n17475) );
  CLKBUF_X1 U12652 ( .A(n17487), .Z(n17488) );
  OR2_X1 U12653 ( .A1(n16688), .A2(n9747), .ZN(n10576) );
  NAND2_X1 U12654 ( .A1(n17524), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n17517) );
  NAND2_X1 U12655 ( .A1(n14439), .A2(n10040), .ZN(n14441) );
  INV_X1 U12656 ( .A(n12804), .ZN(n10040) );
  CLKBUF_X1 U12657 ( .A(n17234), .Z(n17235) );
  NAND2_X1 U12658 ( .A1(n10385), .A2(n17249), .ZN(n17531) );
  INV_X1 U12659 ( .A(n14849), .ZN(n21079) );
  INV_X1 U12660 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21065) );
  OR2_X1 U12661 ( .A1(n21058), .A2(n21072), .ZN(n21062) );
  NAND2_X1 U12662 ( .A1(n10641), .A2(n14282), .ZN(n14285) );
  INV_X1 U12663 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18043) );
  NAND2_X1 U12664 ( .A1(n13822), .A2(n14275), .ZN(n13826) );
  AOI21_X1 U12665 ( .B1(n14743), .B2(n20237), .A(n13618), .ZN(n17555) );
  INV_X1 U12666 ( .A(n20599), .ZN(n20606) );
  OAI21_X1 U12667 ( .B1(n20655), .B2(n21041), .A(n20654), .ZN(n20674) );
  NAND2_X1 U12668 ( .A1(n10371), .A2(n20834), .ZN(n10370) );
  OAI21_X1 U12669 ( .B1(n20783), .B2(n20751), .A(n20750), .ZN(n20774) );
  NOR2_X1 U12670 ( .A1(n20753), .A2(n21062), .ZN(n20829) );
  AOI21_X1 U12671 ( .B1(n20900), .B2(n14865), .A(n14864), .ZN(n20823) );
  INV_X1 U12672 ( .A(n20829), .ZN(n20867) );
  INV_X1 U12673 ( .A(n20587), .ZN(n20907) );
  INV_X1 U12674 ( .A(n20590), .ZN(n20914) );
  INV_X1 U12675 ( .A(n20469), .ZN(n20911) );
  INV_X1 U12676 ( .A(n20474), .ZN(n20921) );
  INV_X1 U12677 ( .A(n20595), .ZN(n20928) );
  INV_X1 U12678 ( .A(n20855), .ZN(n20934) );
  INV_X1 U12679 ( .A(n20479), .ZN(n20935) );
  INV_X1 U12680 ( .A(n20602), .ZN(n20941) );
  INV_X1 U12681 ( .A(n20672), .ZN(n20947) );
  INV_X1 U12682 ( .A(n20611), .ZN(n21835) );
  AND2_X1 U12683 ( .A1(n20903), .A2(n20902), .ZN(n20952) );
  INV_X1 U12684 ( .A(n18142), .ZN(n20237) );
  INV_X1 U12685 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20900) );
  NOR2_X1 U12686 ( .A1(n14750), .A2(n14749), .ZN(n18135) );
  NAND2_X1 U12687 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20965), .ZN(n21095) );
  NOR2_X1 U12688 ( .A1(n13673), .A2(n13672), .ZN(n20226) );
  AND2_X1 U12689 ( .A1(n12049), .A2(n12048), .ZN(n18975) );
  NAND2_X1 U12690 ( .A1(n20212), .A2(n20062), .ZN(n18976) );
  NOR2_X1 U12692 ( .A1(n18265), .A2(n10454), .ZN(n10453) );
  NAND2_X1 U12693 ( .A1(n10456), .A2(n10455), .ZN(n10454) );
  NOR2_X1 U12694 ( .A1(n18568), .A2(n12109), .ZN(n18283) );
  NAND2_X1 U12695 ( .A1(n10451), .A2(n19124), .ZN(n10449) );
  NOR2_X1 U12698 ( .A1(n18359), .A2(n10450), .ZN(n18352) );
  NOR2_X1 U12699 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n18381), .ZN(n18372) );
  NOR2_X1 U12700 ( .A1(n18370), .A2(n10450), .ZN(n18360) );
  NOR2_X1 U12701 ( .A1(n18378), .A2(n10450), .ZN(n18371) );
  NOR2_X1 U12703 ( .A1(n18379), .A2(n18380), .ZN(n18378) );
  NAND2_X1 U12704 ( .A1(n18406), .A2(n10444), .ZN(n18379) );
  NAND2_X1 U12705 ( .A1(n11894), .A2(n18396), .ZN(n10444) );
  NOR2_X1 U12707 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n18472), .ZN(n18471) );
  NAND2_X1 U12708 ( .A1(n18471), .A2(n18461), .ZN(n18460) );
  NOR2_X1 U12709 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n18540), .ZN(n18521) );
  NAND2_X1 U12710 ( .A1(n18550), .A2(n18541), .ZN(n18540) );
  INV_X1 U12712 ( .A(n18552), .ZN(n18589) );
  INV_X1 U12713 ( .A(n18575), .ZN(n18579) );
  OR2_X1 U12714 ( .A1(n20231), .A2(n12112), .ZN(n18522) );
  INV_X1 U12715 ( .A(n18578), .ZN(n18568) );
  OAI211_X1 U12716 ( .C1(n20109), .C2(n20102), .A(n18561), .B(n20229), .ZN(
        n18552) );
  NOR2_X1 U12717 ( .A1(n18610), .A2(n18609), .ZN(n18660) );
  NAND2_X1 U12718 ( .A1(n18808), .A2(n18670), .ZN(n18674) );
  NOR2_X1 U12719 ( .A1(n18709), .A2(n21897), .ZN(n17606) );
  NOR2_X1 U12720 ( .A1(n19654), .A2(n10476), .ZN(n10474) );
  NAND2_X1 U12721 ( .A1(n17686), .A2(n10475), .ZN(n17649) );
  INV_X1 U12722 ( .A(n17688), .ZN(n17686) );
  AND2_X1 U12723 ( .A1(n17686), .A2(P3_EBX_REG_18__SCAN_IN), .ZN(n17684) );
  AND2_X1 U12724 ( .A1(n14473), .A2(n10464), .ZN(n18727) );
  AND2_X1 U12725 ( .A1(n9771), .A2(P3_EBX_REG_16__SCAN_IN), .ZN(n10464) );
  NOR2_X1 U12726 ( .A1(n18423), .A2(n18438), .ZN(n10465) );
  NAND2_X1 U12727 ( .A1(n14473), .A2(n9771), .ZN(n18710) );
  NOR2_X1 U12728 ( .A1(n14472), .A2(n14471), .ZN(n14473) );
  NAND2_X1 U12729 ( .A1(n14473), .A2(P3_EBX_REG_13__SCAN_IN), .ZN(n14790) );
  NOR2_X1 U12730 ( .A1(n18747), .A2(n18751), .ZN(n14095) );
  AND2_X1 U12731 ( .A1(n9768), .A2(P3_EBX_REG_7__SCAN_IN), .ZN(n10478) );
  NAND2_X1 U12732 ( .A1(n10479), .A2(n10480), .ZN(n18792) );
  NAND2_X1 U12733 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n18799), .ZN(n18795) );
  INV_X1 U12734 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n22097) );
  NOR2_X1 U12735 ( .A1(n18795), .A2(n22097), .ZN(n18798) );
  AND2_X1 U12736 ( .A1(n18805), .A2(P3_EBX_REG_2__SCAN_IN), .ZN(n18799) );
  INV_X1 U12737 ( .A(n10466), .ZN(n18805) );
  AOI22_X1 U12738 ( .A1(n13848), .A2(n10468), .B1(n10668), .B2(n10467), .ZN(
        n10466) );
  NOR2_X1 U12739 ( .A1(n10471), .A2(n10469), .ZN(n10468) );
  INV_X1 U12740 ( .A(n10470), .ZN(n10467) );
  INV_X2 U12741 ( .A(n18812), .ZN(n18808) );
  OAI21_X1 U12742 ( .B1(n10473), .B2(n10471), .A(n10470), .ZN(n18814) );
  AND2_X1 U12743 ( .A1(n18814), .A2(n19654), .ZN(n18812) );
  NOR2_X1 U12744 ( .A1(n18993), .A2(n18831), .ZN(n18824) );
  INV_X1 U12745 ( .A(n18838), .ZN(n18832) );
  NAND2_X1 U12746 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n18832), .ZN(n18831) );
  INV_X1 U12747 ( .A(n18851), .ZN(n18847) );
  NAND2_X1 U12748 ( .A1(n18847), .A2(P3_EAX_REG_25__SCAN_IN), .ZN(n18846) );
  AND2_X1 U12749 ( .A1(n18880), .A2(n10271), .ZN(n18852) );
  NOR2_X1 U12750 ( .A1(n19654), .A2(n10273), .ZN(n10271) );
  AND2_X1 U12751 ( .A1(n18817), .A2(n17728), .ZN(n17727) );
  NAND2_X1 U12752 ( .A1(n18880), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n18879) );
  AND2_X1 U12753 ( .A1(n17711), .A2(n18606), .ZN(n18896) );
  OR2_X1 U12754 ( .A1(n13882), .A2(n10267), .ZN(n18901) );
  NAND2_X1 U12755 ( .A1(n10268), .A2(P3_EAX_REG_8__SCAN_IN), .ZN(n10267) );
  INV_X1 U12756 ( .A(n10269), .ZN(n10268) );
  NOR2_X1 U12757 ( .A1(n13882), .A2(n10269), .ZN(n18903) );
  INV_X1 U12758 ( .A(n18913), .ZN(n18900) );
  INV_X1 U12759 ( .A(n17942), .ZN(n17778) );
  AND2_X1 U12760 ( .A1(n13929), .A2(P3_EAX_REG_2__SCAN_IN), .ZN(n13930) );
  NOR2_X1 U12761 ( .A1(n13882), .A2(n18969), .ZN(n13908) );
  AND4_X1 U12762 ( .A1(n13646), .A2(n13645), .A3(n13644), .A4(n13643), .ZN(
        n13647) );
  AND4_X1 U12763 ( .A1(n13638), .A2(n13637), .A3(n13636), .A4(n13635), .ZN(
        n13649) );
  INV_X1 U12764 ( .A(n19022), .ZN(n19012) );
  OR2_X1 U12765 ( .A1(n20098), .A2(n18976), .ZN(n19022) );
  OAI21_X1 U12766 ( .B1(n19024), .B2(n19196), .A(n19026), .ZN(n17944) );
  INV_X1 U12767 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n19031) );
  NAND2_X1 U12768 ( .A1(n19132), .A2(n17764), .ZN(n19072) );
  INV_X1 U12769 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n19122) );
  OAI21_X1 U12770 ( .B1(n10312), .B2(n10311), .A(n10309), .ZN(n17926) );
  AND2_X1 U12771 ( .A1(n10310), .A2(n17920), .ZN(n10309) );
  OR2_X1 U12772 ( .A1(n17921), .A2(n19504), .ZN(n10310) );
  OAI21_X1 U12773 ( .B1(n17926), .B2(n10306), .A(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n10305) );
  NAND2_X1 U12774 ( .A1(n10308), .A2(n10307), .ZN(n10306) );
  NAND2_X1 U12775 ( .A1(n19497), .A2(n17939), .ZN(n10308) );
  INV_X1 U12776 ( .A(n17927), .ZN(n10307) );
  NOR2_X1 U12777 ( .A1(n19189), .A2(n9767), .ZN(n19059) );
  NAND2_X1 U12778 ( .A1(n19420), .A2(n19079), .ZN(n19395) );
  OR2_X1 U12779 ( .A1(n10261), .A2(n13871), .ZN(n13671) );
  NAND2_X1 U12780 ( .A1(n19198), .A2(n17856), .ZN(n17878) );
  NAND2_X1 U12781 ( .A1(n14214), .A2(n14213), .ZN(n19274) );
  INV_X1 U12782 ( .A(n20064), .ZN(n19587) );
  INV_X1 U12783 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20088) );
  INV_X1 U12784 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14032) );
  INV_X2 U12785 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13787) );
  NOR2_X1 U12786 ( .A1(n19627), .A2(n13781), .ZN(n14055) );
  INV_X1 U12787 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n21986) );
  INV_X1 U12789 ( .A(U212), .ZN(n18193) );
  OAI21_X1 U12790 ( .B1(n11797), .B2(n21143), .A(n11678), .ZN(n11679) );
  OAI21_X1 U12791 ( .B1(n16010), .B2(n21105), .A(n10362), .ZN(P1_U2969) );
  NAND2_X1 U12792 ( .A1(n16108), .A2(n11832), .ZN(n16082) );
  OAI21_X1 U12793 ( .B1(n10497), .B2(n20351), .A(n10492), .ZN(P2_U2826) );
  XNOR2_X1 U12794 ( .A(n16426), .B(n16975), .ZN(n10497) );
  AND2_X1 U12795 ( .A1(n10159), .A2(n10156), .ZN(n10155) );
  MUX2_X1 U12796 ( .A(n15352), .B(n15347), .S(n9713), .Z(n15348) );
  NAND2_X1 U12797 ( .A1(n10683), .A2(n15358), .ZN(n10105) );
  NAND2_X1 U12798 ( .A1(n16978), .A2(n18107), .ZN(n9916) );
  INV_X1 U12799 ( .A(n16970), .ZN(n16978) );
  NAND2_X1 U12800 ( .A1(n10285), .A2(n10284), .ZN(n16994) );
  NAND2_X1 U12801 ( .A1(n10286), .A2(n10459), .ZN(n10285) );
  NAND2_X1 U12802 ( .A1(n10288), .A2(n9808), .ZN(n10284) );
  INV_X1 U12803 ( .A(n17025), .ZN(n9999) );
  OR2_X1 U12804 ( .A1(n17299), .A2(n17252), .ZN(n10002) );
  NAND2_X1 U12805 ( .A1(n17297), .A2(n18108), .ZN(n10000) );
  NAND2_X1 U12806 ( .A1(n10435), .A2(n10434), .ZN(n10433) );
  NAND2_X1 U12807 ( .A1(n9793), .A2(n18105), .ZN(n9985) );
  INV_X1 U12808 ( .A(n9981), .ZN(n9980) );
  OAI21_X1 U12809 ( .B1(n17411), .B2(n17252), .A(n17141), .ZN(n9981) );
  OAI21_X1 U12810 ( .B1(n9782), .B2(n17500), .A(n10192), .ZN(P2_U3016) );
  OAI21_X1 U12811 ( .B1(n15352), .B2(n17518), .A(n9822), .ZN(n10193) );
  OR2_X1 U12812 ( .A1(n16970), .A2(n17518), .ZN(n10658) );
  NAND2_X1 U12813 ( .A1(n16986), .A2(n18126), .ZN(n10407) );
  OAI211_X1 U12814 ( .C1(n17261), .C2(n17500), .A(n17262), .B(n10318), .ZN(
        P2_U3019) );
  NAND2_X1 U12815 ( .A1(n10287), .A2(n16992), .ZN(n17261) );
  INV_X1 U12816 ( .A(n17285), .ZN(n10340) );
  NAND2_X1 U12817 ( .A1(n17286), .A2(n18126), .ZN(n10342) );
  NAND2_X1 U12818 ( .A1(n17313), .A2(n18126), .ZN(n17322) );
  OAI211_X1 U12819 ( .C1(n17056), .C2(n17500), .A(n13376), .B(n13377), .ZN(
        P2_U3025) );
  AOI21_X1 U12820 ( .B1(n17072), .B2(n10056), .A(n17348), .ZN(n17349) );
  INV_X1 U12821 ( .A(n10057), .ZN(n10056) );
  NAND2_X1 U12822 ( .A1(n9793), .A2(n18118), .ZN(n9986) );
  NAND2_X1 U12823 ( .A1(n10251), .A2(n18118), .ZN(n10250) );
  AOI21_X1 U12824 ( .B1(n17377), .B2(n10256), .A(n10255), .ZN(n10254) );
  NAND2_X1 U12825 ( .A1(n10615), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10614) );
  INV_X1 U12826 ( .A(n9983), .ZN(n9982) );
  NAND2_X1 U12827 ( .A1(n10073), .A2(n10071), .ZN(P2_U3035) );
  INV_X1 U12828 ( .A(n10072), .ZN(n10071) );
  NOR4_X1 U12829 ( .A1(n12117), .A2(n13380), .A3(n12116), .A4(n12115), .ZN(
        n12118) );
  NAND2_X1 U12830 ( .A1(n11896), .A2(n18598), .ZN(n12119) );
  OAI21_X1 U12831 ( .B1(n18260), .B2(n10457), .A(n10452), .ZN(P3_U2642) );
  INV_X1 U12832 ( .A(n10458), .ZN(n10457) );
  AND2_X1 U12833 ( .A1(n18268), .A2(n10453), .ZN(n10452) );
  AOI21_X1 U12834 ( .B1(n18262), .B2(n18261), .A(n18584), .ZN(n10458) );
  NAND2_X1 U12835 ( .A1(n18880), .A2(n10272), .ZN(n18856) );
  OR2_X1 U12836 ( .A1(n13882), .A2(n10270), .ZN(n18908) );
  AOI21_X1 U12837 ( .B1(n19602), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n9902), .ZN(n9918) );
  NAND2_X1 U12838 ( .A1(n10004), .A2(n19530), .ZN(n10003) );
  NAND2_X1 U12839 ( .A1(n19361), .A2(n19598), .ZN(n9917) );
  AND3_X1 U12841 ( .A1(n10359), .A2(n10358), .A3(n18050), .ZN(n9738) );
  NAND2_X1 U12842 ( .A1(n9774), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9739) );
  OR2_X1 U12843 ( .A1(n20217), .A2(n18243), .ZN(n9740) );
  OAI21_X1 U12844 ( .B1(n11699), .B2(n11820), .A(n11698), .ZN(n11707) );
  OAI21_X1 U12845 ( .B1(n10385), .B2(n10337), .A(n16695), .ZN(n17231) );
  NAND2_X1 U12846 ( .A1(n10628), .A2(n10629), .ZN(n15479) );
  NAND2_X1 U12847 ( .A1(n10620), .A2(n10657), .ZN(n15549) );
  AND2_X1 U12848 ( .A1(n16535), .A2(n16537), .ZN(n13371) );
  NAND2_X1 U12849 ( .A1(n14821), .A2(n14884), .ZN(n14883) );
  NAND2_X1 U12850 ( .A1(n15416), .A2(n15417), .ZN(n15402) );
  NAND2_X1 U12851 ( .A1(n14027), .A2(n11917), .ZN(n11974) );
  INV_X1 U12852 ( .A(n11974), .ZN(n18717) );
  AND2_X2 U12853 ( .A1(n10700), .A2(n13805), .ZN(n10938) );
  AND2_X1 U12854 ( .A1(n18917), .A2(n20212), .ZN(n9741) );
  AND2_X1 U12855 ( .A1(n12685), .A2(n10366), .ZN(n9742) );
  AND2_X1 U12856 ( .A1(n16532), .A2(n9869), .ZN(n13365) );
  AND2_X1 U12857 ( .A1(n12988), .A2(n10583), .ZN(n9743) );
  OR2_X1 U12858 ( .A1(n10420), .A2(n10419), .ZN(n9744) );
  INV_X1 U12859 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13229) );
  NOR2_X1 U12860 ( .A1(n17481), .A2(n13168), .ZN(n17457) );
  INV_X1 U12861 ( .A(n17457), .ZN(n10034) );
  NAND2_X1 U12862 ( .A1(n11775), .A2(n15909), .ZN(n9745) );
  AND2_X1 U12863 ( .A1(n9879), .A2(n15062), .ZN(n9746) );
  INV_X1 U12864 ( .A(n10561), .ZN(n15991) );
  OR2_X1 U12865 ( .A1(n16959), .A2(n16962), .ZN(n9747) );
  OR3_X1 U12866 ( .A1(n16434), .A2(n16433), .A3(n16740), .ZN(n9748) );
  INV_X1 U12867 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n19165) );
  AND4_X1 U12868 ( .A1(n10069), .A2(n12743), .A3(n13354), .A4(n13350), .ZN(
        n9749) );
  AND2_X1 U12869 ( .A1(n15909), .A2(n9901), .ZN(n9750) );
  INV_X1 U12870 ( .A(n17919), .ZN(n10312) );
  AND2_X1 U12871 ( .A1(n10499), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n9751) );
  AND2_X1 U12872 ( .A1(n10364), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n9752) );
  NAND2_X1 U12873 ( .A1(n10628), .A2(n10626), .ZN(n10631) );
  OR2_X1 U12874 ( .A1(n11553), .A2(n11554), .ZN(n9753) );
  INV_X1 U12875 ( .A(n10185), .ZN(n12695) );
  AND2_X1 U12876 ( .A1(n10382), .A2(n13204), .ZN(n9754) );
  NAND2_X1 U12877 ( .A1(n10116), .A2(n10115), .ZN(n9755) );
  NAND2_X1 U12878 ( .A1(n10339), .A2(n9910), .ZN(n17000) );
  NAND2_X1 U12879 ( .A1(n13570), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10920) );
  INV_X1 U12880 ( .A(n10920), .ZN(n10078) );
  INV_X1 U12881 ( .A(n12219), .ZN(n10104) );
  AND2_X1 U12882 ( .A1(n17026), .A2(n9976), .ZN(n9756) );
  AND2_X1 U12883 ( .A1(n10969), .A2(n9858), .ZN(n9757) );
  INV_X1 U12884 ( .A(n19196), .ZN(n10323) );
  NOR2_X1 U12885 ( .A1(n14521), .A2(n15350), .ZN(n9758) );
  NAND2_X1 U12886 ( .A1(n10364), .A2(n9880), .ZN(n9759) );
  NAND2_X1 U12887 ( .A1(n10951), .A2(n10950), .ZN(n9760) );
  AND2_X1 U12888 ( .A1(n9897), .A2(n16452), .ZN(n9761) );
  INV_X1 U12889 ( .A(n11829), .ZN(n10090) );
  AND2_X1 U12890 ( .A1(n10538), .A2(n10537), .ZN(n9762) );
  AND2_X1 U12891 ( .A1(n9762), .A2(n15379), .ZN(n9763) );
  AND2_X1 U12892 ( .A1(n9761), .A2(n10581), .ZN(n9764) );
  AND2_X1 U12893 ( .A1(n12636), .A2(n12638), .ZN(n9765) );
  AND2_X1 U12894 ( .A1(n10401), .A2(n12934), .ZN(n9766) );
  INV_X2 U12895 ( .A(n14466), .ZN(n13862) );
  NAND2_X1 U12896 ( .A1(n10316), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9767) );
  INV_X1 U12897 ( .A(n14200), .ZN(n10322) );
  AND2_X1 U12898 ( .A1(n10480), .A2(P3_EBX_REG_6__SCAN_IN), .ZN(n9768) );
  AND2_X1 U12899 ( .A1(n10474), .A2(P3_EBX_REG_20__SCAN_IN), .ZN(n9769) );
  AND2_X1 U12900 ( .A1(n17327), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9770) );
  AND2_X1 U12901 ( .A1(n10465), .A2(P3_EBX_REG_15__SCAN_IN), .ZN(n9771) );
  AND2_X1 U12902 ( .A1(n17327), .A2(n10405), .ZN(n9772) );
  AND2_X1 U12903 ( .A1(n13362), .A2(n17035), .ZN(n9773) );
  AND2_X1 U12904 ( .A1(n10554), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9774) );
  AND2_X1 U12905 ( .A1(n10460), .A2(P3_EBX_REG_25__SCAN_IN), .ZN(n9775) );
  AND2_X1 U12906 ( .A1(n10398), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9776) );
  AND2_X1 U12907 ( .A1(n10405), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9777) );
  AND2_X2 U12908 ( .A1(n15153), .A2(n14684), .ZN(n12350) );
  NAND2_X1 U12909 ( .A1(n16373), .A2(n10859), .ZN(n14754) );
  INV_X1 U12910 ( .A(n14238), .ZN(n11577) );
  NAND2_X1 U12911 ( .A1(n15898), .A2(n15897), .ZN(n15870) );
  AND2_X1 U12912 ( .A1(n10564), .A2(n9876), .ZN(n15999) );
  INV_X1 U12913 ( .A(n17607), .ZN(n17630) );
  NAND2_X1 U12914 ( .A1(n14028), .A2(n10432), .ZN(n17607) );
  AND2_X1 U12915 ( .A1(n17606), .A2(n10462), .ZN(n9779) );
  AND2_X1 U12916 ( .A1(n15416), .A2(n9762), .ZN(n9780) );
  NAND2_X1 U12917 ( .A1(n14019), .A2(n11907), .ZN(n9781) );
  INV_X1 U12918 ( .A(n10205), .ZN(n18129) );
  NAND2_X1 U12919 ( .A1(n13984), .A2(n17361), .ZN(n10205) );
  NOR2_X1 U12920 ( .A1(n16441), .A2(n16442), .ZN(n13205) );
  AND2_X1 U12921 ( .A1(n17854), .A2(n11891), .ZN(n11883) );
  XOR2_X1 U12922 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n13215), .Z(
        n9782) );
  AND2_X1 U12923 ( .A1(n10700), .A2(n10699), .ZN(n10756) );
  NAND2_X1 U12924 ( .A1(n14708), .A2(n15153), .ZN(n9783) );
  AND2_X1 U12925 ( .A1(n10801), .A2(n10817), .ZN(n11684) );
  NOR2_X1 U12926 ( .A1(n15504), .A2(n15505), .ZN(n15492) );
  NOR2_X1 U12927 ( .A1(n14879), .A2(n10621), .ZN(n15537) );
  NAND2_X1 U12928 ( .A1(n10504), .A2(n10505), .ZN(n12686) );
  NAND2_X1 U12929 ( .A1(n16532), .A2(n13103), .ZN(n13364) );
  NAND2_X1 U12930 ( .A1(n13371), .A2(n13373), .ZN(n13372) );
  OR2_X1 U12931 ( .A1(n10034), .A2(n10196), .ZN(n9785) );
  AND2_X1 U12932 ( .A1(n11240), .A2(n10052), .ZN(n9786) );
  OR2_X1 U12933 ( .A1(n10295), .A2(n10294), .ZN(n10290) );
  NAND2_X1 U12934 ( .A1(n10224), .A2(n10640), .ZN(n14333) );
  AND4_X1 U12935 ( .A1(n12203), .A2(n10206), .A3(n12211), .A4(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n9787) );
  AND2_X1 U12936 ( .A1(n10240), .A2(n10528), .ZN(n9788) );
  AND2_X1 U12937 ( .A1(n10583), .A2(n14642), .ZN(n9789) );
  AND2_X1 U12938 ( .A1(n13274), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13273) );
  NOR2_X1 U12939 ( .A1(n16552), .A2(n16802), .ZN(n16535) );
  AND3_X1 U12940 ( .A1(n9971), .A2(n12221), .A3(n9970), .ZN(n9790) );
  AND2_X1 U12941 ( .A1(n12671), .A2(n10243), .ZN(n9791) );
  AND3_X1 U12942 ( .A1(n14784), .A2(n14785), .A3(n10624), .ZN(n9792) );
  XOR2_X1 U12943 ( .A(n17078), .B(n17077), .Z(n9793) );
  NAND2_X1 U12944 ( .A1(n10508), .A2(n10509), .ZN(n12722) );
  AND2_X1 U12945 ( .A1(n17764), .A2(n19078), .ZN(n9794) );
  INV_X1 U12946 ( .A(n10074), .ZN(n12242) );
  INV_X1 U12947 ( .A(n13239), .ZN(n10412) );
  INV_X1 U12948 ( .A(n12290), .ZN(n10617) );
  INV_X1 U12949 ( .A(n9967), .ZN(n10958) );
  AND2_X1 U12950 ( .A1(n16953), .A2(n14807), .ZN(n9795) );
  AND3_X1 U12951 ( .A1(n12543), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        n10337), .ZN(n9796) );
  AND2_X1 U12952 ( .A1(n10415), .A2(n10412), .ZN(n9797) );
  NAND2_X1 U12953 ( .A1(n10354), .A2(n11737), .ZN(n18049) );
  NAND2_X1 U12954 ( .A1(n12541), .A2(n12540), .ZN(n17192) );
  AND2_X1 U12955 ( .A1(n10524), .A2(n10523), .ZN(n9798) );
  AND3_X1 U12956 ( .A1(n10153), .A2(n10152), .A3(n10151), .ZN(n9799) );
  AND2_X1 U12957 ( .A1(n15920), .A2(n15930), .ZN(n9800) );
  AND2_X1 U12958 ( .A1(n9760), .A2(n11030), .ZN(n9801) );
  INV_X1 U12959 ( .A(n12905), .ZN(n10206) );
  NAND2_X1 U12960 ( .A1(n10555), .A2(n11733), .ZN(n14503) );
  INV_X1 U12961 ( .A(n15993), .ZN(n15909) );
  INV_X1 U12962 ( .A(n12685), .ZN(n12515) );
  NAND2_X1 U12963 ( .A1(n12504), .A2(n12503), .ZN(n12685) );
  AND2_X1 U12964 ( .A1(n13822), .A2(n12266), .ZN(n9802) );
  AND2_X1 U12965 ( .A1(n12731), .A2(n12730), .ZN(n9803) );
  NAND2_X1 U12966 ( .A1(n16532), .A2(n10586), .ZN(n16495) );
  NAND2_X1 U12967 ( .A1(n10359), .A2(n10358), .ZN(n10562) );
  AND2_X1 U12968 ( .A1(n19265), .A2(n19264), .ZN(n9804) );
  AND2_X1 U12969 ( .A1(n10513), .A2(n12633), .ZN(n9805) );
  AND2_X1 U12970 ( .A1(n12207), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9806) );
  INV_X1 U12971 ( .A(n12694), .ZN(n10503) );
  INV_X1 U12972 ( .A(n14591), .ZN(n14069) );
  INV_X1 U12973 ( .A(n14561), .ZN(n10045) );
  NOR2_X1 U12974 ( .A1(n15366), .A2(n15365), .ZN(n9807) );
  AND2_X1 U12975 ( .A1(n10459), .A2(n17256), .ZN(n9808) );
  AND2_X1 U12976 ( .A1(n12901), .A2(n20433), .ZN(n9809) );
  NAND2_X1 U12977 ( .A1(n19476), .A2(n19188), .ZN(n19189) );
  INV_X1 U12978 ( .A(n19189), .ZN(n10315) );
  AND2_X1 U12979 ( .A1(n15979), .A2(n16176), .ZN(n9810) );
  NOR2_X1 U12980 ( .A1(n17362), .A2(n10616), .ZN(n9811) );
  AND2_X1 U12981 ( .A1(n17756), .A2(n19073), .ZN(n9812) );
  AND2_X1 U12982 ( .A1(n10035), .A2(n10033), .ZN(n9813) );
  OR2_X1 U12983 ( .A1(n17079), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9814) );
  NAND2_X1 U12984 ( .A1(n10163), .A2(n9939), .ZN(n9815) );
  INV_X1 U12985 ( .A(n12291), .ZN(n9992) );
  AND2_X1 U12986 ( .A1(n11541), .A2(n11561), .ZN(n9816) );
  AND2_X1 U12987 ( .A1(n11534), .A2(n11561), .ZN(n9817) );
  NAND2_X1 U12988 ( .A1(n12574), .A2(n10104), .ZN(n9818) );
  AND2_X1 U12989 ( .A1(n12504), .A2(n10367), .ZN(n9819) );
  INV_X1 U12990 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13965) );
  NOR2_X1 U12991 ( .A1(n16203), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9820) );
  AND3_X1 U12992 ( .A1(n13874), .A2(n13849), .A3(n19638), .ZN(n9821) );
  OR3_X1 U12993 ( .A1(n16514), .A2(n12627), .A3(n17035), .ZN(n17037) );
  INV_X1 U12994 ( .A(n17037), .ZN(n10113) );
  INV_X1 U12995 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n22046) );
  AND2_X1 U12996 ( .A1(n10044), .A2(n13176), .ZN(n9822) );
  OR2_X1 U12997 ( .A1(n14392), .A2(n11082), .ZN(n9823) );
  NAND2_X2 U12998 ( .A1(n9951), .A2(n9950), .ZN(n14331) );
  AND2_X1 U12999 ( .A1(n12145), .A2(n10129), .ZN(n9824) );
  AND4_X1 U13000 ( .A1(n12317), .A2(n12316), .A3(n12315), .A4(n12314), .ZN(
        n9825) );
  INV_X1 U13001 ( .A(n10031), .ZN(n10030) );
  NOR2_X1 U13002 ( .A1(n10034), .A2(n17366), .ZN(n10031) );
  OR2_X1 U13003 ( .A1(n15909), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9826) );
  AND2_X1 U13004 ( .A1(n17856), .A2(n10323), .ZN(n9827) );
  INV_X1 U13005 ( .A(n10596), .ZN(n10595) );
  OR2_X1 U13006 ( .A1(n13347), .A2(n10597), .ZN(n10596) );
  NAND3_X1 U13007 ( .A1(n13357), .A2(n12765), .A3(n17076), .ZN(n9828) );
  AND2_X1 U13008 ( .A1(n20059), .A2(n18973), .ZN(n9829) );
  AND2_X1 U13009 ( .A1(n14839), .A2(n14840), .ZN(n9830) );
  NAND2_X1 U13010 ( .A1(n10049), .A2(n11099), .ZN(n14879) );
  NAND2_X1 U13011 ( .A1(n13822), .A2(n12271), .ZN(n12280) );
  INV_X1 U13012 ( .A(n12280), .ZN(n9990) );
  AND3_X1 U13013 ( .A1(n13353), .A2(n17121), .A3(n10070), .ZN(n9831) );
  AND2_X1 U13014 ( .A1(n10591), .A2(n9938), .ZN(n9832) );
  AND2_X1 U13015 ( .A1(n11539), .A2(n11538), .ZN(n9833) );
  AND2_X1 U13016 ( .A1(n17606), .A2(n9775), .ZN(n18672) );
  NAND2_X1 U13017 ( .A1(n12213), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12219) );
  NAND2_X1 U13018 ( .A1(n16535), .A2(n10039), .ZN(n16466) );
  AND2_X1 U13019 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12299) );
  AND2_X1 U13020 ( .A1(n10014), .A2(n17763), .ZN(n9834) );
  INV_X1 U13021 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n19053) );
  AND2_X1 U13022 ( .A1(n10566), .A2(n10421), .ZN(n9835) );
  INV_X1 U13023 ( .A(n15470), .ZN(n11318) );
  NAND2_X1 U13024 ( .A1(n19045), .A2(n22049), .ZN(n9836) );
  AND2_X1 U13025 ( .A1(n16451), .A2(n9764), .ZN(n9837) );
  AND2_X1 U13026 ( .A1(n16996), .A2(n17026), .ZN(n9838) );
  AND3_X1 U13027 ( .A1(n15280), .A2(n16752), .A3(n10651), .ZN(n9839) );
  AND2_X1 U13028 ( .A1(n13824), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12312) );
  AND2_X1 U13029 ( .A1(n9701), .A2(n18108), .ZN(n9840) );
  AND2_X1 U13030 ( .A1(n9701), .A2(n18126), .ZN(n9841) );
  AND2_X1 U13031 ( .A1(n10552), .A2(n13170), .ZN(n9842) );
  AND2_X1 U13032 ( .A1(n9941), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9843) );
  AND2_X1 U13033 ( .A1(n9721), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n9844)
         );
  AND2_X1 U13034 ( .A1(n16977), .A2(n16976), .ZN(n9845) );
  AND2_X1 U13035 ( .A1(n10758), .A2(n10757), .ZN(n9846) );
  NAND2_X1 U13036 ( .A1(n11509), .A2(n11784), .ZN(n11553) );
  AND2_X1 U13037 ( .A1(n10225), .A2(n14278), .ZN(n9847) );
  AND2_X1 U13038 ( .A1(n9721), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n9848) );
  AND2_X1 U13039 ( .A1(n9798), .A2(n16482), .ZN(n9849) );
  NOR2_X1 U13040 ( .A1(n18291), .A2(n10450), .ZN(n9850) );
  AND2_X1 U13041 ( .A1(n10505), .A2(n10503), .ZN(n9851) );
  NOR2_X1 U13042 ( .A1(n10536), .A2(n10535), .ZN(n9852) );
  OR2_X1 U13043 ( .A1(n16437), .A2(n16980), .ZN(n9853) );
  NAND2_X1 U13044 ( .A1(n11552), .A2(n11564), .ZN(n9854) );
  INV_X1 U13045 ( .A(n12703), .ZN(n10422) );
  AND2_X1 U13046 ( .A1(n14281), .A2(n14435), .ZN(n9855) );
  AND2_X1 U13047 ( .A1(n10589), .A2(n10588), .ZN(n9856) );
  AND2_X1 U13048 ( .A1(n9789), .A2(n10582), .ZN(n9857) );
  AND2_X1 U13049 ( .A1(n9801), .A2(n11042), .ZN(n9858) );
  NAND2_X1 U13050 ( .A1(n19070), .A2(n19196), .ZN(n9859) );
  INV_X1 U13051 ( .A(n13204), .ZN(n10381) );
  AND2_X1 U13052 ( .A1(n9826), .A2(n11763), .ZN(n9860) );
  NAND2_X1 U13053 ( .A1(n10906), .A2(n11717), .ZN(n9861) );
  AND2_X1 U13054 ( .A1(n10646), .A2(n10649), .ZN(n9862) );
  AND2_X1 U13055 ( .A1(n11351), .A2(n11350), .ZN(n15457) );
  INV_X1 U13056 ( .A(n18050), .ZN(n10357) );
  INV_X1 U13057 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14352) );
  NAND2_X1 U13058 ( .A1(n10661), .A2(n16768), .ZN(n15256) );
  AND3_X1 U13059 ( .A1(n12937), .A2(n12936), .A3(n12935), .ZN(n16959) );
  INV_X1 U13060 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12088) );
  AND2_X1 U13061 ( .A1(n13831), .A2(n20237), .ZN(n16835) );
  INV_X1 U13062 ( .A(n12920), .ZN(n13106) );
  AND2_X1 U13063 ( .A1(n12796), .A2(n13145), .ZN(n18118) );
  NOR2_X1 U13064 ( .A1(n11875), .A2(n19053), .ZN(n17782) );
  INV_X1 U13065 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20834) );
  OR2_X1 U13066 ( .A1(n10337), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9863) );
  NOR2_X1 U13067 ( .A1(n16816), .A2(n16811), .ZN(n16806) );
  AND2_X1 U13068 ( .A1(n15063), .A2(n10227), .ZN(n9864) );
  NAND2_X1 U13069 ( .A1(n15526), .A2(n15527), .ZN(n15506) );
  NAND2_X1 U13070 ( .A1(n10036), .A2(n10519), .ZN(n16551) );
  NOR2_X1 U13071 ( .A1(n16816), .A2(n10653), .ZN(n16796) );
  NAND2_X1 U13072 ( .A1(n13289), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13292) );
  AND2_X1 U13073 ( .A1(n17606), .A2(n10460), .ZN(n9865) );
  NAND2_X1 U13074 ( .A1(n12796), .A2(n15209), .ZN(n17500) );
  INV_X1 U13075 ( .A(n17500), .ZN(n18126) );
  AND2_X1 U13076 ( .A1(n17606), .A2(P3_EBX_REG_22__SCAN_IN), .ZN(n9866) );
  AND2_X1 U13077 ( .A1(n18847), .A2(n10264), .ZN(n9867) );
  NOR2_X1 U13078 ( .A1(n14534), .A2(n14811), .ZN(n14812) );
  AND2_X1 U13079 ( .A1(n14812), .A2(n14822), .ZN(n14821) );
  INV_X1 U13080 ( .A(n12627), .ZN(n10337) );
  INV_X1 U13081 ( .A(n19505), .ZN(n19530) );
  NAND2_X1 U13082 ( .A1(n14619), .A2(n9795), .ZN(n16588) );
  NAND2_X1 U13083 ( .A1(n14812), .A2(n10041), .ZN(n14647) );
  NAND2_X1 U13084 ( .A1(n12988), .A2(n9789), .ZN(n14638) );
  AND2_X1 U13085 ( .A1(n10548), .A2(n10547), .ZN(n9868) );
  XNOR2_X1 U13086 ( .A(n11736), .B(n18080), .ZN(n18055) );
  NAND2_X1 U13087 ( .A1(n10576), .A2(n10579), .ZN(n14623) );
  AND2_X1 U13088 ( .A1(n14812), .A2(n10042), .ZN(n14833) );
  NAND2_X1 U13089 ( .A1(n14821), .A2(n10518), .ZN(n16613) );
  INV_X1 U13090 ( .A(n17057), .ZN(n10603) );
  OR2_X1 U13091 ( .A1(n16688), .A2(n16959), .ZN(n16958) );
  NAND2_X1 U13092 ( .A1(n12988), .A2(n12987), .ZN(n14602) );
  AND2_X1 U13093 ( .A1(n9957), .A2(n13142), .ZN(n13135) );
  AND2_X1 U13094 ( .A1(n13103), .A2(n10587), .ZN(n9869) );
  AND2_X1 U13095 ( .A1(n20057), .A2(n19598), .ZN(n19610) );
  INV_X1 U13096 ( .A(n19610), .ZN(n10311) );
  NAND2_X1 U13097 ( .A1(n13676), .A2(n13675), .ZN(n13687) );
  AND2_X1 U13098 ( .A1(n11826), .A2(n11825), .ZN(n16234) );
  AND2_X1 U13099 ( .A1(n14473), .A2(n10465), .ZN(n9870) );
  AND2_X1 U13100 ( .A1(n17686), .A2(n10474), .ZN(n9871) );
  AND2_X1 U13101 ( .A1(n12631), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n9872) );
  AND2_X1 U13103 ( .A1(n17500), .A2(n17361), .ZN(n9873) );
  NOR2_X1 U13104 ( .A1(n18352), .A2(n19124), .ZN(n9874) );
  AND2_X1 U13105 ( .A1(n10227), .A2(n16788), .ZN(n9875) );
  INV_X1 U13106 ( .A(n21305), .ZN(n10046) );
  INV_X2 U13107 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n17596) );
  OR2_X1 U13108 ( .A1(n12418), .A2(n12417), .ZN(n12934) );
  OR2_X1 U13109 ( .A1(n12664), .A2(n12657), .ZN(n10060) );
  INV_X1 U13110 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20085) );
  INV_X1 U13111 ( .A(n12318), .ZN(n10400) );
  NAND2_X1 U13112 ( .A1(n11745), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9876) );
  NOR2_X1 U13113 ( .A1(n12502), .A2(n12501), .ZN(n12943) );
  AND2_X1 U13114 ( .A1(n16774), .A2(n15213), .ZN(n9877) );
  NAND2_X1 U13115 ( .A1(n20062), .A2(n20218), .ZN(n9878) );
  AND2_X1 U13116 ( .A1(n10652), .A2(n15116), .ZN(n9879) );
  AND3_X1 U13117 ( .A1(n12203), .A2(n10206), .A3(n12211), .ZN(n9880) );
  AND2_X1 U13118 ( .A1(n15796), .A2(n16014), .ZN(n9881) );
  AND2_X1 U13119 ( .A1(n10429), .A2(n10426), .ZN(n9882) );
  AND3_X1 U13120 ( .A1(n12805), .A2(n14439), .A3(n10515), .ZN(n9883) );
  AND2_X1 U13121 ( .A1(n12470), .A2(n12627), .ZN(n9884) );
  AND2_X1 U13122 ( .A1(n10519), .A2(n12854), .ZN(n9885) );
  AND2_X1 U13123 ( .A1(n12393), .A2(n9766), .ZN(n9886) );
  OR2_X1 U13124 ( .A1(n11875), .A2(n10441), .ZN(n9887) );
  AND2_X1 U13125 ( .A1(n10446), .A2(n10451), .ZN(n9888) );
  AND2_X1 U13126 ( .A1(n9765), .A2(n10511), .ZN(n9889) );
  INV_X1 U13127 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10011) );
  INV_X1 U13128 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n12089) );
  INV_X1 U13129 ( .A(n18795), .ZN(n10479) );
  INV_X1 U13130 ( .A(n17218), .ZN(n18108) );
  NOR2_X1 U13131 ( .A1(n11875), .A2(n10440), .ZN(n11873) );
  AND2_X1 U13132 ( .A1(n10479), .A2(n9768), .ZN(n9891) );
  NOR2_X1 U13133 ( .A1(n14075), .A2(n14074), .ZN(n9892) );
  INV_X1 U13134 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10144) );
  NOR2_X1 U13135 ( .A1(n13687), .A2(n13771), .ZN(n13848) );
  INV_X1 U13136 ( .A(n13848), .ZN(n10473) );
  INV_X1 U13137 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n21733) );
  INV_X1 U13138 ( .A(n19073), .ZN(n10016) );
  INV_X1 U13139 ( .A(n17084), .ZN(n10150) );
  AND2_X1 U13140 ( .A1(n10323), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9893) );
  INV_X1 U13141 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14685) );
  OR3_X1 U13142 ( .A1(n10196), .A2(n13168), .A3(n10195), .ZN(n9894) );
  OR2_X1 U13143 ( .A1(n20211), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n9895) );
  AND2_X1 U13144 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(P3_EAX_REG_3__SCAN_IN), 
        .ZN(n9896) );
  NAND2_X1 U13145 ( .A1(n13121), .A2(n13120), .ZN(n9897) );
  NAND2_X1 U13146 ( .A1(n13110), .A2(n13109), .ZN(n9898) );
  AND2_X1 U13147 ( .A1(n10323), .A2(n10430), .ZN(n9899) );
  INV_X1 U13148 ( .A(n10486), .ZN(n10485) );
  NAND2_X1 U13149 ( .A1(n10487), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10486) );
  AND2_X1 U13150 ( .A1(n10526), .A2(n13218), .ZN(n9900) );
  INV_X1 U13151 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17573) );
  INV_X1 U13152 ( .A(n20187), .ZN(n20225) );
  INV_X1 U13153 ( .A(n16715), .ZN(n10154) );
  AND3_X1 U13154 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18534) );
  AND3_X1 U13155 ( .A1(n17854), .A2(n9737), .A3(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n19139) );
  INV_X1 U13156 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n10511) );
  NAND4_X1 U13157 ( .A1(n16107), .A2(n16141), .A3(n11772), .A4(n11771), .ZN(
        n9901) );
  AND2_X1 U13158 ( .A1(n19556), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n9902) );
  INV_X1 U13159 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10488) );
  NOR2_X1 U13160 ( .A1(n17328), .A2(n17340), .ZN(n10405) );
  AND2_X1 U13161 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n9774), .ZN(
        n9903) );
  AND2_X1 U13162 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n9904) );
  INV_X1 U13163 ( .A(n10273), .ZN(n10272) );
  NAND2_X1 U13164 ( .A1(n10274), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n10273) );
  INV_X1 U13165 ( .A(n10476), .ZN(n10475) );
  NAND2_X1 U13166 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(P3_EBX_REG_19__SCAN_IN), 
        .ZN(n10476) );
  AND2_X1 U13167 ( .A1(n17327), .A2(n9777), .ZN(n9905) );
  AND2_X1 U13168 ( .A1(n10264), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n9906) );
  AND2_X1 U13169 ( .A1(n9772), .A2(n13361), .ZN(n9907) );
  INV_X1 U13170 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10428) );
  INV_X1 U13171 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n10424) );
  INV_X1 U13172 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n10477) );
  INV_X1 U13173 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10510) );
  INV_X1 U13174 ( .A(n16050), .ZN(n10297) );
  INV_X1 U13175 ( .A(n16029), .ZN(n10147) );
  NAND2_X1 U13176 ( .A1(n17854), .A2(n9737), .ZN(n19164) );
  INV_X1 U13177 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n18554) );
  INV_X1 U13178 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n10266) );
  INV_X1 U13179 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n10265) );
  AND2_X1 U13180 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n9908) );
  AND2_X1 U13181 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n9909) );
  AND2_X1 U13182 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n9910) );
  INV_X1 U13183 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10500) );
  AND2_X1 U13184 ( .A1(n9776), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n9911) );
  INV_X1 U13185 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10338) );
  NOR2_X2 U13186 ( .A1(n15020), .A2(n18057), .ZN(n9912) );
  AND2_X2 U13187 ( .A1(n13435), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n15020)
         );
  NAND2_X1 U13188 ( .A1(n14395), .A2(n11683), .ZN(n18057) );
  OAI21_X1 U13189 ( .B1(n17411), .B2(n17534), .A(n17409), .ZN(n9983) );
  OR2_X1 U13190 ( .A1(n17287), .A2(n17534), .ZN(n10341) );
  OAI21_X1 U13191 ( .B1(n17436), .B2(n17534), .A(n17435), .ZN(n10072) );
  OR2_X1 U13192 ( .A1(n17263), .A2(n17534), .ZN(n10318) );
  OAI21_X1 U13193 ( .B1(n17378), .B2(n17534), .A(n10613), .ZN(n10612) );
  OR2_X1 U13194 ( .A1(n19912), .A2(n19911), .ZN(n19863) );
  AOI22_X2 U13195 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n9698), .B1(DATAI_25_), 
        .B2(n9912), .ZN(n21689) );
  AOI22_X2 U13196 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n9698), .B1(DATAI_21_), 
        .B2(n9912), .ZN(n21597) );
  AOI22_X2 U13197 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n9698), .B1(DATAI_18_), 
        .B2(n9912), .ZN(n21695) );
  AOI22_X2 U13198 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n9698), .B1(DATAI_24_), 
        .B2(n9912), .ZN(n21643) );
  NOR3_X2 U13199 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20110), .A3(
        n19839), .ZN(n19810) );
  INV_X1 U13200 ( .A(n9699), .ZN(n14658) );
  NOR2_X4 U13201 ( .A1(n21751), .A2(n21815), .ZN(n21789) );
  AOI22_X2 U13202 ( .A1(DATAI_22_), .A2(n9912), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n9698), .ZN(n21631) );
  AOI211_X1 U13203 ( .C1(n17376), .C2(n9701), .A(n17218), .B(n17101), .ZN(
        n17102) );
  XNOR2_X2 U13204 ( .A(n10169), .B(n10277), .ZN(n12682) );
  NAND2_X2 U13205 ( .A1(n10280), .A2(n10551), .ZN(n17093) );
  NAND4_X1 U13206 ( .A1(n12004), .A2(n12003), .A3(n12002), .A4(n12001), .ZN(
        n13674) );
  AOI21_X1 U13207 ( .B1(n9720), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A(n9914), .ZN(n12198) );
  OAI21_X2 U13208 ( .B1(n19347), .B2(n19082), .A(n19863), .ZN(n19212) );
  INV_X2 U13209 ( .A(n17966), .ZN(n19526) );
  NAND2_X2 U13210 ( .A1(n18244), .A2(n9895), .ZN(n19313) );
  INV_X2 U13212 ( .A(n18777), .ZN(n14968) );
  NAND4_X1 U13213 ( .A1(n9825), .A2(n12308), .A3(n12309), .A4(n12307), .ZN(
        n12929) );
  NAND2_X1 U13214 ( .A1(n10229), .A2(n9843), .ZN(n10118) );
  NOR2_X2 U13215 ( .A1(n10058), .A2(n12664), .ZN(n10504) );
  INV_X1 U13216 ( .A(n13237), .ZN(n10419) );
  AOI21_X1 U13217 ( .B1(n13409), .B2(n18105), .A(n13247), .ZN(n13248) );
  NAND3_X1 U13218 ( .A1(n12147), .A2(n12149), .A3(n12148), .ZN(n12152) );
  NAND2_X1 U13219 ( .A1(n16971), .A2(n18105), .ZN(n16977) );
  OAI22_X1 U13220 ( .A1(n12301), .A2(n12433), .B1(n20614), .B2(n12289), .ZN(
        n12294) );
  NAND2_X1 U13221 ( .A1(n10414), .A2(n10677), .ZN(n13190) );
  OAI211_X1 U13222 ( .C1(n17218), .C2(n16979), .A(n9845), .B(n9916), .ZN(
        P2_U2985) );
  NOR2_X1 U13223 ( .A1(n19264), .A2(n19265), .ZN(n19263) );
  NAND2_X1 U13224 ( .A1(n19332), .A2(n19333), .ZN(n19331) );
  NAND3_X1 U13225 ( .A1(n10003), .A2(n9918), .A3(n9917), .ZN(P3_U2835) );
  NAND2_X1 U13226 ( .A1(n14185), .A2(n10302), .ZN(n14187) );
  INV_X1 U13227 ( .A(n14400), .ZN(n14186) );
  OAI21_X1 U13228 ( .B1(n20551), .B2(n12285), .A(n10121), .ZN(n12286) );
  BUF_X4 U13229 ( .A(n17093), .Z(n17364) );
  AND3_X2 U13230 ( .A1(n13148), .A2(n20433), .A3(n12905), .ZN(n9920) );
  AND2_X1 U13231 ( .A1(n9920), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n9938) );
  NAND2_X1 U13232 ( .A1(n9919), .A2(n10591), .ZN(n9928) );
  AND2_X1 U13233 ( .A1(n14870), .A2(n9920), .ZN(n9919) );
  NAND2_X1 U13234 ( .A1(n12209), .A2(n9920), .ZN(n12585) );
  NAND3_X1 U13235 ( .A1(n9963), .A2(n11760), .A3(n11762), .ZN(n9923) );
  NAND3_X1 U13236 ( .A1(n9923), .A2(n9921), .A3(n9965), .ZN(n9924) );
  INV_X1 U13237 ( .A(n10359), .ZN(n9922) );
  NAND3_X1 U13238 ( .A1(n10172), .A2(n9860), .A3(n15906), .ZN(n10141) );
  NAND3_X1 U13239 ( .A1(n9738), .A2(n10557), .A3(n18055), .ZN(n9925) );
  NAND2_X2 U13240 ( .A1(n10175), .A2(n11735), .ZN(n10557) );
  AND2_X1 U13241 ( .A1(n12212), .A2(n12174), .ZN(n9929) );
  NAND2_X1 U13242 ( .A1(n10792), .A2(n11719), .ZN(n9930) );
  NAND2_X1 U13243 ( .A1(n9930), .A2(n9933), .ZN(n9931) );
  INV_X1 U13244 ( .A(n10806), .ZN(n11556) );
  NAND3_X1 U13245 ( .A1(n10770), .A2(n9932), .A3(n9931), .ZN(n10806) );
  NAND3_X1 U13246 ( .A1(n11799), .A2(n14591), .A3(n10821), .ZN(n9933) );
  INV_X1 U13247 ( .A(n9934), .ZN(n20685) );
  NAND2_X1 U13248 ( .A1(n9934), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n10371) );
  OAI22_X1 U13249 ( .A1(n20614), .A2(n12435), .B1(n9934), .B2(n13040), .ZN(
        n12436) );
  OAI22_X1 U13250 ( .A1(n20494), .A2(n12292), .B1(n13007), .B2(n9934), .ZN(
        n12293) );
  OR2_X1 U13251 ( .A1(n9937), .A2(n14753), .ZN(n14371) );
  NAND2_X1 U13252 ( .A1(n10840), .A2(n9937), .ZN(n13801) );
  XNOR2_X1 U13253 ( .A(n9937), .B(n14540), .ZN(n14349) );
  OAI211_X2 U13254 ( .C1(n10829), .C2(n10348), .A(n10347), .B(n10836), .ZN(
        n9937) );
  NAND2_X1 U13255 ( .A1(n9940), .A2(n14866), .ZN(n12208) );
  AND2_X1 U13256 ( .A1(n12212), .A2(n9940), .ZN(n9939) );
  AND2_X2 U13257 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14684) );
  NAND2_X2 U13258 ( .A1(n9943), .A2(n9942), .ZN(n12213) );
  INV_X1 U13259 ( .A(n12800), .ZN(n9945) );
  NAND3_X1 U13260 ( .A1(n9956), .A2(n12262), .A3(n12263), .ZN(n9946) );
  XNOR2_X2 U13261 ( .A(n12253), .B(n12252), .ZN(n12263) );
  NAND2_X2 U13262 ( .A1(n12244), .A2(n12243), .ZN(n9956) );
  NAND2_X1 U13263 ( .A1(n9954), .A2(n12129), .ZN(n9948) );
  NAND2_X1 U13264 ( .A1(n9952), .A2(n12129), .ZN(n9950) );
  NAND4_X1 U13265 ( .A1(n12126), .A2(n12128), .A3(n12127), .A4(n12125), .ZN(
        n9952) );
  NAND4_X1 U13266 ( .A1(n12124), .A2(n12121), .A3(n12122), .A4(n12123), .ZN(
        n9953) );
  NAND4_X1 U13267 ( .A1(n12164), .A2(n12165), .A3(n12166), .A4(n12167), .ZN(
        n9954) );
  NAND4_X1 U13268 ( .A1(n12163), .A2(n12162), .A3(n12160), .A4(n12161), .ZN(
        n9955) );
  XNOR2_X1 U13269 ( .A(n9956), .B(n12263), .ZN(n12274) );
  NAND3_X2 U13270 ( .A1(n9957), .A2(n14420), .A3(n13142), .ZN(n12223) );
  INV_X2 U13271 ( .A(n12227), .ZN(n13223) );
  NAND2_X2 U13272 ( .A1(n10053), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12227) );
  OR2_X1 U13273 ( .A1(n12227), .A2(n17526), .ZN(n9958) );
  INV_X1 U13274 ( .A(n9961), .ZN(n9960) );
  XNOR2_X2 U13275 ( .A(n9961), .B(n12242), .ZN(n12265) );
  NAND2_X1 U13276 ( .A1(n9962), .A2(n9990), .ZN(n20832) );
  NAND2_X1 U13277 ( .A1(n10231), .A2(n9962), .ZN(n10230) );
  AND2_X4 U13278 ( .A1(n10170), .A2(n13805), .ZN(n10871) );
  AND2_X2 U13279 ( .A1(n14352), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10170) );
  INV_X1 U13280 ( .A(n9876), .ZN(n9964) );
  NOR2_X1 U13281 ( .A1(n10355), .A2(n9964), .ZN(n9963) );
  NAND2_X1 U13282 ( .A1(n9966), .A2(n11762), .ZN(n9965) );
  AND4_X2 U13283 ( .A1(n9967), .A2(n10968), .A3(n10969), .A4(n9801), .ZN(
        n10353) );
  NAND3_X1 U13284 ( .A1(n9757), .A2(n9702), .A3(n9967), .ZN(n11748) );
  NAND2_X2 U13285 ( .A1(n9969), .A2(n9968), .ZN(n9967) );
  NAND2_X1 U13286 ( .A1(n14349), .A2(n21733), .ZN(n9969) );
  NAND2_X2 U13287 ( .A1(n9787), .A2(n10364), .ZN(n12248) );
  NAND2_X2 U13288 ( .A1(n12611), .A2(n12220), .ZN(n12879) );
  INV_X1 U13289 ( .A(n12540), .ZN(n10610) );
  AOI21_X1 U13290 ( .B1(n9994), .B2(n9840), .A(n17116), .ZN(n17117) );
  NAND2_X1 U13291 ( .A1(n9994), .A2(n9841), .ZN(n9993) );
  INV_X1 U13292 ( .A(n10554), .ZN(n9973) );
  NAND2_X2 U13293 ( .A1(n10339), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17011) );
  NAND2_X2 U13294 ( .A1(n10281), .A2(n10282), .ZN(n10339) );
  NOR2_X2 U13295 ( .A1(n17113), .A2(n17376), .ZN(n17101) );
  OAI21_X1 U13296 ( .B1(n17040), .B2(n10113), .A(n9756), .ZN(n9979) );
  INV_X1 U13297 ( .A(n17038), .ZN(n9977) );
  NAND2_X1 U13298 ( .A1(n10373), .A2(n17037), .ZN(n17027) );
  NAND2_X1 U13299 ( .A1(n17020), .A2(n10338), .ZN(n10190) );
  NAND2_X1 U13300 ( .A1(n17142), .A2(n9980), .ZN(P2_U3001) );
  NAND2_X1 U13301 ( .A1(n17410), .A2(n9982), .ZN(P2_U3033) );
  NAND4_X1 U13302 ( .A1(n9984), .A2(n12505), .A3(n12425), .A4(n17223), .ZN(
        n10215) );
  NAND3_X1 U13303 ( .A1(n17223), .A2(n12425), .A3(n9984), .ZN(n17221) );
  NAND2_X1 U13304 ( .A1(n17086), .A2(n9985), .ZN(P2_U2996) );
  NAND2_X1 U13305 ( .A1(n17360), .A2(n9986), .ZN(P2_U3028) );
  NAND2_X1 U13306 ( .A1(n12421), .A2(n10277), .ZN(n12423) );
  NAND3_X1 U13307 ( .A1(n10207), .A2(n10209), .A3(n12403), .ZN(n12422) );
  NOR2_X1 U13308 ( .A1(n12901), .A2(n12898), .ZN(n12893) );
  NAND2_X1 U13309 ( .A1(n12513), .A2(n9988), .ZN(n10216) );
  AND2_X2 U13310 ( .A1(n12275), .A2(n14287), .ZN(n9991) );
  OAI211_X1 U13311 ( .C1(n17387), .C2(n17534), .A(n9995), .B(n9993), .ZN(
        P2_U3031) );
  NOR2_X1 U13312 ( .A1(n17386), .A2(n17385), .ZN(n9995) );
  NOR2_X1 U13313 ( .A1(n9844), .A2(n9996), .ZN(n10140) );
  NAND3_X1 U13314 ( .A1(n9998), .A2(n12129), .A3(n9997), .ZN(n9996) );
  NAND3_X1 U13315 ( .A1(n10002), .A2(n10000), .A3(n9999), .ZN(P2_U2990) );
  NAND3_X1 U13316 ( .A1(n10006), .A2(n19027), .A3(n10005), .ZN(n19362) );
  NAND3_X1 U13317 ( .A1(n19025), .A2(n19026), .A3(n19196), .ZN(n10006) );
  NAND3_X1 U13318 ( .A1(n14213), .A2(n10431), .A3(n14214), .ZN(n19276) );
  NAND2_X1 U13319 ( .A1(n19302), .A2(n14205), .ZN(n19288) );
  NAND2_X1 U13320 ( .A1(n19302), .A2(n10008), .ZN(n14213) );
  OAI21_X1 U13321 ( .B1(n19326), .B2(n19325), .A(n10013), .ZN(n19327) );
  NAND2_X1 U13322 ( .A1(n19326), .A2(n19325), .ZN(n10013) );
  OAI21_X1 U13323 ( .B1(n19198), .B2(n19197), .A(n19196), .ZN(n19222) );
  NAND2_X1 U13324 ( .A1(n17204), .A2(n10552), .ZN(n10280) );
  NAND2_X1 U13325 ( .A1(n17487), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10021) );
  NAND3_X1 U13326 ( .A1(n10216), .A2(n10215), .A3(n12512), .ZN(n17487) );
  NAND2_X1 U13327 ( .A1(n10026), .A2(n10025), .ZN(n10024) );
  NAND2_X1 U13328 ( .A1(n10614), .A2(n9813), .ZN(P2_U3030) );
  INV_X1 U13329 ( .A(n10612), .ZN(n10035) );
  NAND2_X1 U13330 ( .A1(n10036), .A2(n9885), .ZN(n16552) );
  NOR2_X1 U13331 ( .A1(n14287), .A2(n17573), .ZN(n10218) );
  NOR2_X2 U13332 ( .A1(n21270), .A2(n10045), .ZN(n21260) );
  NAND2_X1 U13333 ( .A1(n10047), .A2(n11174), .ZN(n10977) );
  NAND2_X1 U13334 ( .A1(n10047), .A2(n11784), .ZN(n11715) );
  NAND2_X1 U13335 ( .A1(n10046), .A2(n21304), .ZN(n21529) );
  NAND2_X1 U13336 ( .A1(n10047), .A2(n9967), .ZN(n21673) );
  MUX2_X1 U13337 ( .A(n21672), .B(n14613), .S(n21304), .Z(n14386) );
  NAND2_X1 U13338 ( .A1(n10049), .A2(n10048), .ZN(n15528) );
  NAND4_X1 U13339 ( .A1(n12223), .A2(n12218), .A3(n13621), .A4(n14748), .ZN(
        n10053) );
  NAND2_X1 U13340 ( .A1(n9851), .A2(n10504), .ZN(n12629) );
  INV_X1 U13341 ( .A(n10060), .ZN(n12655) );
  INV_X1 U13342 ( .A(n10504), .ZN(n12675) );
  NAND2_X1 U13343 ( .A1(n12731), .A2(n10061), .ZN(n12740) );
  NAND2_X1 U13344 ( .A1(n12740), .A2(n9872), .ZN(n10063) );
  INV_X1 U13345 ( .A(n10062), .ZN(n12717) );
  NAND2_X1 U13346 ( .A1(n10063), .A2(n10062), .ZN(n20278) );
  NAND2_X1 U13347 ( .A1(n12731), .A2(n10513), .ZN(n10062) );
  NAND2_X1 U13348 ( .A1(n17424), .A2(n18126), .ZN(n10073) );
  NAND4_X1 U13349 ( .A1(n12450), .A2(n12447), .A3(n12449), .A4(n12448), .ZN(
        n12471) );
  NAND2_X1 U13350 ( .A1(n10081), .A2(n10080), .ZN(n11539) );
  INV_X1 U13351 ( .A(n16234), .ZN(n10093) );
  NAND2_X1 U13352 ( .A1(n10095), .A2(n16108), .ZN(n16068) );
  NAND2_X1 U13353 ( .A1(n16137), .A2(n16234), .ZN(n16240) );
  NAND4_X1 U13354 ( .A1(n10099), .A2(n10100), .A3(n10102), .A4(n10098), .ZN(
        n11782) );
  NAND3_X1 U13355 ( .A1(n10099), .A2(n10100), .A3(n10102), .ZN(n17992) );
  AND2_X1 U13356 ( .A1(n11545), .A2(n9854), .ZN(n10103) );
  INV_X1 U13357 ( .A(n10373), .ZN(n10107) );
  NAND2_X1 U13358 ( .A1(n10107), .A2(n10372), .ZN(n10110) );
  NAND2_X1 U13359 ( .A1(n10110), .A2(n10111), .ZN(n16997) );
  NAND2_X1 U13360 ( .A1(n10114), .A2(n13145), .ZN(n10346) );
  NOR2_X1 U13361 ( .A1(n10114), .A2(n10400), .ZN(n10335) );
  NAND4_X1 U13362 ( .A1(n12295), .A2(n12297), .A3(n12296), .A4(n12298), .ZN(
        n10114) );
  INV_X1 U13363 ( .A(n12611), .ZN(n10116) );
  NAND3_X1 U13364 ( .A1(n10118), .A2(n12238), .A3(n10117), .ZN(n12245) );
  NAND3_X1 U13365 ( .A1(n10116), .A2(n10104), .A3(n10115), .ZN(n12238) );
  NAND2_X1 U13366 ( .A1(n10229), .A2(n9941), .ZN(n12231) );
  NAND2_X1 U13367 ( .A1(n12230), .A2(n9806), .ZN(n10117) );
  NAND2_X1 U13368 ( .A1(n17364), .A2(n13362), .ZN(n17036) );
  NAND2_X1 U13369 ( .A1(n17364), .A2(n9773), .ZN(n10119) );
  NAND2_X2 U13370 ( .A1(n10123), .A2(n10122), .ZN(n12288) );
  NAND3_X1 U13371 ( .A1(n10123), .A2(n10122), .A3(n9802), .ZN(n20646) );
  OR2_X2 U13372 ( .A1(n12291), .A2(n12288), .ZN(n20551) );
  NAND2_X1 U13373 ( .A1(n10127), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10126) );
  NAND4_X1 U13374 ( .A1(n9824), .A2(n12146), .A3(n12144), .A4(n10128), .ZN(
        n10127) );
  NAND2_X1 U13375 ( .A1(n9720), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n10128) );
  NAND2_X1 U13376 ( .A1(n9721), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n10132) );
  NAND2_X1 U13377 ( .A1(n9719), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n10134) );
  NAND2_X2 U13378 ( .A1(n10138), .A2(n10135), .ZN(n20433) );
  NAND4_X1 U13379 ( .A1(n10137), .A2(n12169), .A3(n12170), .A4(n10136), .ZN(
        n10135) );
  NAND4_X1 U13380 ( .A1(n10140), .A2(n12172), .A3(n12171), .A4(n10139), .ZN(
        n10138) );
  NAND2_X2 U13381 ( .A1(n10143), .A2(n10141), .ZN(n15898) );
  NAND3_X1 U13382 ( .A1(n9745), .A2(n10145), .A3(n15796), .ZN(n11862) );
  NAND3_X1 U13383 ( .A1(n9745), .A2(n10145), .A3(n9881), .ZN(n10149) );
  NAND3_X1 U13384 ( .A1(n11738), .A2(n11748), .A3(n11784), .ZN(n11744) );
  NAND3_X1 U13385 ( .A1(n9748), .A2(n10155), .A3(n9853), .ZN(P2_U2827) );
  NOR2_X2 U13386 ( .A1(n16501), .A2(n17028), .ZN(n16487) );
  NOR2_X2 U13387 ( .A1(n10161), .A2(n10160), .ZN(n16501) );
  NAND4_X1 U13388 ( .A1(n11799), .A2(n10821), .A3(n14591), .A4(n10162), .ZN(
        n10802) );
  NAND2_X1 U13389 ( .A1(n17204), .A2(n9842), .ZN(n10281) );
  NAND2_X1 U13390 ( .A1(n9992), .A2(n10168), .ZN(n12433) );
  AND2_X4 U13391 ( .A1(n10707), .A2(n10170), .ZN(n10876) );
  NAND2_X1 U13392 ( .A1(n9835), .A2(n10171), .ZN(n11773) );
  NAND2_X1 U13393 ( .A1(n10172), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15981) );
  NAND2_X1 U13394 ( .A1(n10174), .A2(n10173), .ZN(n15982) );
  NAND2_X1 U13395 ( .A1(n10935), .A2(n9967), .ZN(n10959) );
  NAND2_X1 U13396 ( .A1(n10180), .A2(n10178), .ZN(n11699) );
  AOI21_X1 U13397 ( .B1(n10935), .B2(n9967), .A(n9760), .ZN(n10179) );
  AND2_X2 U13398 ( .A1(n15857), .A2(n10182), .ZN(n15812) );
  NAND3_X1 U13399 ( .A1(n9749), .A2(n17490), .A3(n17489), .ZN(n10184) );
  OAI21_X1 U13400 ( .B1(n17020), .B2(n10338), .A(n17018), .ZN(n10191) );
  AOI21_X2 U13401 ( .B1(n15357), .B2(n18118), .A(n10193), .ZN(n10192) );
  NAND3_X1 U13402 ( .A1(n10317), .A2(n12401), .A3(n12420), .ZN(n17248) );
  NAND3_X1 U13403 ( .A1(n10208), .A2(n10212), .A3(n12401), .ZN(n10207) );
  NAND3_X1 U13404 ( .A1(n10210), .A2(n12401), .A3(n10211), .ZN(n10209) );
  NAND2_X1 U13405 ( .A1(n17105), .A2(n10213), .ZN(P2_U2998) );
  NAND2_X1 U13406 ( .A1(n10214), .A2(n18105), .ZN(n10213) );
  INV_X1 U13407 ( .A(n17378), .ZN(n10214) );
  OAI21_X1 U13408 ( .B1(n20646), .B2(n12363), .A(n10220), .ZN(n12322) );
  INV_X1 U13409 ( .A(n10222), .ZN(n15278) );
  INV_X1 U13410 ( .A(n13998), .ZN(n10223) );
  NAND2_X1 U13411 ( .A1(n10223), .A2(n14282), .ZN(n10226) );
  NAND2_X1 U13412 ( .A1(n14279), .A2(n14278), .ZN(n14334) );
  NAND2_X1 U13413 ( .A1(n14279), .A2(n9847), .ZN(n14281) );
  NAND2_X1 U13414 ( .A1(n13144), .A2(n12228), .ZN(n10229) );
  OAI21_X1 U13415 ( .B1(n20460), .B2(n13006), .A(n10230), .ZN(n12282) );
  OAI22_X1 U13416 ( .A1(n20614), .A2(n12329), .B1(n12328), .B2(n20832), .ZN(
        n12330) );
  NAND2_X1 U13417 ( .A1(n10236), .A2(n10277), .ZN(n10234) );
  NAND2_X1 U13418 ( .A1(n12690), .A2(n10244), .ZN(n10239) );
  NAND3_X1 U13419 ( .A1(n10254), .A2(n10252), .A3(n10250), .ZN(P2_U3029) );
  NAND2_X1 U13420 ( .A1(n10260), .A2(n10257), .ZN(n13875) );
  OR2_X1 U13421 ( .A1(n12085), .A2(n13689), .ZN(n10263) );
  INV_X1 U13422 ( .A(n10263), .ZN(n13670) );
  INV_X1 U13423 ( .A(n10261), .ZN(n14033) );
  INV_X1 U13424 ( .A(n12086), .ZN(n10262) );
  NAND2_X1 U13425 ( .A1(n18847), .A2(n9906), .ZN(n18838) );
  NAND2_X1 U13426 ( .A1(n10277), .A2(n9819), .ZN(n10276) );
  NAND2_X1 U13427 ( .A1(n17364), .A2(n9772), .ZN(n17072) );
  NAND2_X1 U13428 ( .A1(n17364), .A2(n9907), .ZN(n10278) );
  NAND2_X1 U13429 ( .A1(n17364), .A2(n17327), .ZN(n17094) );
  INV_X1 U13430 ( .A(n12513), .ZN(n17222) );
  INV_X1 U13431 ( .A(n17001), .ZN(n10288) );
  OR2_X1 U13432 ( .A1(n17001), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10287) );
  OAI21_X1 U13433 ( .B1(n11855), .B2(n21105), .A(n10565), .ZN(P1_U2968) );
  NAND3_X1 U13434 ( .A1(n10293), .A2(n9800), .A3(n10292), .ZN(n10291) );
  INV_X1 U13435 ( .A(n10295), .ZN(n15928) );
  NAND2_X1 U13436 ( .A1(n11767), .A2(n15939), .ZN(n10295) );
  NAND2_X2 U13437 ( .A1(n14402), .A2(n14403), .ZN(n19188) );
  NAND3_X1 U13438 ( .A1(n17930), .A2(n17931), .A3(n10305), .ZN(n17933) );
  NOR2_X2 U13439 ( .A1(n19189), .A2(n17843), .ZN(n19405) );
  NAND2_X1 U13440 ( .A1(n10317), .A2(n12420), .ZN(n10385) );
  NAND2_X1 U13441 ( .A1(n14201), .A2(n10322), .ZN(n14202) );
  NOR2_X1 U13442 ( .A1(n14200), .A2(n10424), .ZN(n10321) );
  XNOR2_X1 U13443 ( .A(n14201), .B(n14200), .ZN(n19318) );
  NAND2_X1 U13444 ( .A1(n17759), .A2(n10325), .ZN(n10324) );
  INV_X1 U13445 ( .A(n19100), .ZN(n10328) );
  NAND2_X1 U13446 ( .A1(n19132), .A2(n19100), .ZN(n19160) );
  NAND2_X1 U13447 ( .A1(n19045), .A2(n10331), .ZN(n10330) );
  NAND2_X4 U13448 ( .A1(n11916), .A2(n14019), .ZN(n18715) );
  INV_X1 U13449 ( .A(n10335), .ZN(n10334) );
  INV_X1 U13450 ( .A(n12262), .ZN(n10336) );
  NAND3_X1 U13451 ( .A1(n10342), .A2(n10341), .A3(n10340), .ZN(P2_U3021) );
  NAND2_X1 U13452 ( .A1(n10345), .A2(n12211), .ZN(n10344) );
  INV_X2 U13453 ( .A(n13148), .ZN(n12211) );
  NAND3_X1 U13454 ( .A1(n12206), .A2(n9715), .A3(n12215), .ZN(n10345) );
  NAND2_X1 U13455 ( .A1(n10353), .A2(n10350), .ZN(n10349) );
  NAND2_X1 U13456 ( .A1(n11754), .A2(n11784), .ZN(n11759) );
  AND2_X1 U13457 ( .A1(n10352), .A2(n11042), .ZN(n10350) );
  INV_X1 U13458 ( .A(n11045), .ZN(n10352) );
  NAND2_X1 U13459 ( .A1(n10557), .A2(n18055), .ZN(n10354) );
  NOR2_X1 U13460 ( .A1(n10357), .A2(n11737), .ZN(n10355) );
  INV_X1 U13461 ( .A(n18055), .ZN(n10356) );
  INV_X1 U13462 ( .A(n18044), .ZN(n16000) );
  NAND2_X1 U13463 ( .A1(n10361), .A2(n10360), .ZN(n10359) );
  INV_X1 U13464 ( .A(n16989), .ZN(n10375) );
  NAND3_X1 U13465 ( .A1(n10379), .A2(n10376), .A3(n10374), .ZN(n16988) );
  NAND4_X1 U13466 ( .A1(n10379), .A2(n10376), .A3(n18118), .A4(n10374), .ZN(
        n10380) );
  NAND2_X1 U13467 ( .A1(n9754), .A2(n10375), .ZN(n10374) );
  NAND2_X1 U13468 ( .A1(n13200), .A2(n13201), .ZN(n10382) );
  INV_X1 U13469 ( .A(n10382), .ZN(n10378) );
  NAND3_X1 U13470 ( .A1(n16989), .A2(n10381), .A3(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10379) );
  NAND3_X1 U13471 ( .A1(n10407), .A2(n13214), .A3(n10380), .ZN(P2_U3018) );
  NAND2_X1 U13472 ( .A1(n10384), .A2(n17179), .ZN(n10383) );
  OAI21_X1 U13473 ( .B1(n17098), .B2(n10389), .A(n10386), .ZN(n10388) );
  NAND4_X1 U13474 ( .A1(n12340), .A2(n12337), .A3(n12339), .A4(n12338), .ZN(
        n10402) );
  NAND2_X1 U13475 ( .A1(n17364), .A2(n9905), .ZN(n10404) );
  NAND2_X2 U13476 ( .A1(n10406), .A2(n12589), .ZN(n13142) );
  NAND2_X2 U13477 ( .A1(n12213), .A2(n9735), .ZN(n12589) );
  AND2_X4 U13478 ( .A1(n10408), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14708) );
  NAND2_X1 U13479 ( .A1(n16997), .A2(n9797), .ZN(n10411) );
  NAND2_X1 U13480 ( .A1(n16997), .A2(n12784), .ZN(n10414) );
  AOI21_X1 U13481 ( .B1(n9797), .B2(n10418), .A(n9744), .ZN(n10410) );
  AOI21_X2 U13482 ( .B1(n10677), .B2(n10417), .A(n10416), .ZN(n10415) );
  INV_X1 U13483 ( .A(n10677), .ZN(n10418) );
  NAND2_X1 U13484 ( .A1(n11773), .A2(n15909), .ZN(n15827) );
  NAND2_X1 U13485 ( .A1(n10425), .A2(n14202), .ZN(n19304) );
  NAND2_X1 U13486 ( .A1(n19318), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10425) );
  XNOR2_X1 U13487 ( .A(n14223), .B(n14221), .ZN(n19268) );
  NAND3_X1 U13488 ( .A1(n12201), .A2(n12202), .A3(n14866), .ZN(n12606) );
  NAND2_X1 U13489 ( .A1(n13146), .A2(n13148), .ZN(n12205) );
  AND2_X1 U13490 ( .A1(n17072), .A2(n18108), .ZN(n10436) );
  INV_X1 U13491 ( .A(n10437), .ZN(n11870) );
  INV_X1 U13493 ( .A(n18545), .ZN(n10443) );
  NAND2_X1 U13494 ( .A1(n10443), .A2(n10442), .ZN(n11889) );
  AND2_X1 U13495 ( .A1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10442) );
  NAND2_X1 U13496 ( .A1(n10445), .A2(n10446), .ZN(n18280) );
  OAI21_X1 U13497 ( .B1(n18359), .B2(n10450), .A(n10449), .ZN(n18342) );
  NAND4_X2 U13498 ( .A1(n17854), .A2(n9737), .A3(n10673), .A4(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11882) );
  NAND3_X1 U13499 ( .A1(n12611), .A2(n12220), .A3(P2_REIP_REG_3__SCAN_IN), 
        .ZN(n12258) );
  NAND2_X2 U13500 ( .A1(n11897), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n18755) );
  NAND2_X1 U13501 ( .A1(n17686), .A2(n9769), .ZN(n18709) );
  NAND2_X1 U13502 ( .A1(n10479), .A2(n10478), .ZN(n18781) );
  NAND3_X1 U13503 ( .A1(n10484), .A2(n10482), .A3(n10481), .ZN(n13252) );
  NOR2_X2 U13504 ( .A1(n13290), .A2(n17071), .ZN(n13289) );
  NOR2_X1 U13505 ( .A1(n16970), .A2(n20345), .ZN(n10496) );
  NAND2_X1 U13506 ( .A1(n13277), .A2(n10498), .ZN(n13284) );
  NOR2_X2 U13507 ( .A1(n13262), .A2(n20340), .ZN(n13264) );
  INV_X1 U13508 ( .A(n12620), .ZN(n12592) );
  NAND2_X1 U13509 ( .A1(n12620), .A2(n9987), .ZN(n10501) );
  NAND2_X1 U13511 ( .A1(n10508), .A2(n10507), .ZN(n12719) );
  NAND2_X1 U13512 ( .A1(n12637), .A2(n9765), .ZN(n12647) );
  NAND2_X1 U13513 ( .A1(n12637), .A2(n12636), .ZN(n12653) );
  AND2_X2 U13514 ( .A1(n12637), .A2(n9889), .ZN(n12643) );
  NAND3_X1 U13515 ( .A1(n12650), .A2(n16996), .A3(n12775), .ZN(n12776) );
  NAND3_X1 U13516 ( .A1(n12805), .A2(n14439), .A3(n10514), .ZN(n14498) );
  INV_X1 U13517 ( .A(n14498), .ZN(n12818) );
  AND2_X1 U13518 ( .A1(n13205), .A2(n10526), .ZN(n13219) );
  AND2_X1 U13519 ( .A1(n13205), .A2(n13207), .ZN(n13177) );
  NAND2_X1 U13520 ( .A1(n13205), .A2(n9900), .ZN(n10527) );
  INV_X1 U13521 ( .A(n13198), .ZN(n10531) );
  NAND2_X1 U13522 ( .A1(n12208), .A2(n12174), .ZN(n12175) );
  INV_X1 U13523 ( .A(n14521), .ZN(n10534) );
  NAND2_X1 U13524 ( .A1(n10534), .A2(n9852), .ZN(n14876) );
  NOR2_X2 U13525 ( .A1(n14875), .A2(n10540), .ZN(n15601) );
  NAND2_X1 U13526 ( .A1(n17205), .A2(n12539), .ZN(n12541) );
  INV_X1 U13527 ( .A(n12539), .ZN(n10553) );
  XNOR2_X1 U13528 ( .A(n11732), .B(n11827), .ZN(n14072) );
  NAND2_X1 U13529 ( .A1(n11731), .A2(n11730), .ZN(n11732) );
  XNOR2_X1 U13530 ( .A(n10557), .B(n10356), .ZN(n18083) );
  AND2_X2 U13531 ( .A1(n10558), .A2(n10796), .ZN(n11555) );
  NAND2_X1 U13532 ( .A1(n10560), .A2(n9724), .ZN(n10559) );
  NAND2_X1 U13533 ( .A1(n18049), .A2(n18050), .ZN(n10564) );
  AOI21_X1 U13534 ( .B1(n10564), .B2(n10563), .A(n10562), .ZN(n10561) );
  NAND2_X1 U13535 ( .A1(n15898), .A2(n10572), .ZN(n10569) );
  NAND3_X1 U13536 ( .A1(n16373), .A2(n10859), .A3(n21733), .ZN(n10574) );
  NAND2_X1 U13537 ( .A1(n16688), .A2(n10579), .ZN(n10575) );
  NAND2_X1 U13538 ( .A1(n10575), .A2(n10577), .ZN(n12948) );
  AND2_X2 U13539 ( .A1(n16532), .A2(n10585), .ZN(n16483) );
  AND2_X1 U13540 ( .A1(n13349), .A2(n17109), .ZN(n10600) );
  OAI21_X1 U13541 ( .B1(n17078), .B2(n10605), .A(n10602), .ZN(n13359) );
  AND2_X1 U13542 ( .A1(n17363), .A2(n17380), .ZN(n10616) );
  OAI21_X2 U13543 ( .B1(n13801), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n10856), 
        .ZN(n10969) );
  NAND4_X1 U13544 ( .A1(n10760), .A2(n10686), .A3(n9846), .A4(n10759), .ZN(
        n10769) );
  NAND3_X1 U13545 ( .A1(n14784), .A2(n10623), .A3(n14785), .ZN(n14845) );
  NAND2_X1 U13546 ( .A1(n14784), .A2(n14785), .ZN(n14788) );
  INV_X1 U13547 ( .A(n14819), .ZN(n10624) );
  INV_X1 U13548 ( .A(n10631), .ZN(n15469) );
  AND2_X1 U13549 ( .A1(n15442), .A2(n10635), .ZN(n15418) );
  NAND2_X1 U13550 ( .A1(n15442), .A2(n15443), .ZN(n15431) );
  NAND2_X1 U13551 ( .A1(n12201), .A2(n12202), .ZN(n12604) );
  NAND2_X1 U13552 ( .A1(n14284), .A2(n14282), .ZN(n10640) );
  NAND3_X1 U13553 ( .A1(n15280), .A2(n16752), .A3(n10650), .ZN(n10649) );
  NAND3_X1 U13554 ( .A1(n15280), .A2(n16752), .A3(n10643), .ZN(n10642) );
  NAND2_X1 U13555 ( .A1(n15280), .A2(n16752), .ZN(n16758) );
  INV_X1 U13556 ( .A(n16757), .ZN(n10651) );
  INV_X1 U13557 ( .A(n16979), .ZN(n13194) );
  OR2_X1 U13558 ( .A1(n16938), .A2(n12905), .ZN(n16934) );
  NAND2_X1 U13559 ( .A1(n13231), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13271) );
  INV_X1 U13560 ( .A(n13267), .ZN(n13231) );
  NAND2_X1 U13561 ( .A1(n12818), .A2(n12817), .ZN(n14534) );
  OAI21_X1 U13562 ( .B1(n13193), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n13215), .ZN(n16979) );
  NOR2_X1 U13563 ( .A1(n18271), .A2(n10450), .ZN(n18262) );
  AND2_X1 U13564 ( .A1(n15063), .A2(n14433), .ZN(n14654) );
  NOR2_X4 U13565 ( .A1(n14591), .A2(n10952), .ZN(n10992) );
  NAND2_X1 U13566 ( .A1(n11569), .A2(n11781), .ZN(n14350) );
  NAND2_X1 U13567 ( .A1(n10803), .A2(n14561), .ZN(n11806) );
  INV_X1 U13568 ( .A(n14561), .ZN(n11661) );
  XNOR2_X1 U13569 ( .A(n10813), .B(n10833), .ZN(n10857) );
  AND2_X2 U13571 ( .A1(n15157), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12451) );
  AOI22_X1 U13572 ( .A1(n15157), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9730), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12130) );
  OAI211_X1 U13573 ( .C1(n12248), .C2(n16707), .A(n12250), .B(n12249), .ZN(
        n12251) );
  INV_X1 U13574 ( .A(n21105), .ZN(n11864) );
  NOR2_X1 U13575 ( .A1(n14342), .A2(n14056), .ZN(n10656) );
  AND4_X1 U13576 ( .A1(n11185), .A2(n15569), .A3(n15568), .A4(n15598), .ZN(
        n10657) );
  INV_X1 U13577 ( .A(n11455), .ZN(n11278) );
  NOR2_X1 U13578 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11161) );
  NAND2_X1 U13579 ( .A1(n13422), .A2(n13421), .ZN(n15781) );
  OR3_X1 U13580 ( .A1(n16012), .A2(n11839), .A3(n13815), .ZN(n10659) );
  NOR2_X1 U13581 ( .A1(n11658), .A2(n13570), .ZN(n10660) );
  NAND2_X2 U13582 ( .A1(n15786), .A2(n14594), .ZN(n15790) );
  AND2_X1 U13583 ( .A1(n11808), .A2(n15651), .ZN(n10663) );
  AND2_X1 U13584 ( .A1(n12217), .A2(n12905), .ZN(n10665) );
  NOR3_X1 U13585 ( .A1(n16500), .A2(n12627), .A3(n12772), .ZN(n10666) );
  AND2_X1 U13586 ( .A1(n15979), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10667) );
  AND2_X1 U13587 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n10668) );
  INV_X1 U13588 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n15370) );
  INV_X1 U13589 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10830) );
  INV_X1 U13590 ( .A(n12341), .ZN(n12523) );
  NAND2_X1 U13591 ( .A1(n18112), .A2(n13457), .ZN(n17242) );
  INV_X1 U13592 ( .A(n17242), .ZN(n18107) );
  INV_X1 U13593 ( .A(n15338), .ZN(n15337) );
  NAND2_X2 U13594 ( .A1(n13455), .A2(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n15338)
         );
  NOR2_X1 U13595 ( .A1(n21453), .A2(n21480), .ZN(n10670) );
  INV_X1 U13596 ( .A(n17252), .ZN(n18105) );
  AND2_X1 U13597 ( .A1(n12130), .A2(n12129), .ZN(n10671) );
  AND2_X1 U13598 ( .A1(n15253), .A2(n15274), .ZN(n10672) );
  NOR2_X1 U13599 ( .A1(n19214), .A2(n19306), .ZN(n19123) );
  INV_X1 U13600 ( .A(n19123), .ZN(n19082) );
  INV_X1 U13601 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n20107) );
  AND2_X1 U13602 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10673) );
  AND2_X1 U13603 ( .A1(n15630), .A2(n15629), .ZN(n10674) );
  AND2_X1 U13604 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10675) );
  XNOR2_X1 U13605 ( .A(n13397), .B(n13396), .ZN(n15361) );
  AND4_X1 U13606 ( .A1(n12345), .A2(n12344), .A3(n12343), .A4(n12342), .ZN(
        n10676) );
  INV_X1 U13607 ( .A(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n19819) );
  INV_X1 U13608 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n13232) );
  INV_X1 U13609 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20307) );
  AND2_X1 U13610 ( .A1(n12792), .A2(n13203), .ZN(n10677) );
  OR2_X1 U13611 ( .A1(n13201), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10678) );
  AND2_X1 U13612 ( .A1(n16992), .A2(n13197), .ZN(n10679) );
  OR3_X1 U13613 ( .A1(n13392), .A2(n13391), .A3(n13390), .ZN(P3_U2640) );
  NAND2_X2 U13614 ( .A1(n12159), .A2(n12158), .ZN(n12905) );
  AND2_X1 U13615 ( .A1(n18102), .A2(n13252), .ZN(n10681) );
  INV_X1 U13616 ( .A(n11972), .ZN(n14112) );
  OR2_X1 U13617 ( .A1(n15352), .A2(n17242), .ZN(n10683) );
  INV_X1 U13618 ( .A(n17530), .ZN(n14288) );
  AND4_X1 U13619 ( .A1(n10774), .A2(n10773), .A3(n10772), .A4(n10771), .ZN(
        n10685) );
  AND4_X1 U13620 ( .A1(n10764), .A2(n10763), .A3(n10762), .A4(n10761), .ZN(
        n10686) );
  AND4_X1 U13621 ( .A1(n10735), .A2(n10734), .A3(n10733), .A4(n10732), .ZN(
        n10687) );
  AND4_X1 U13622 ( .A1(n10779), .A2(n10778), .A3(n10777), .A4(n10776), .ZN(
        n10688) );
  NOR2_X2 U13623 ( .A1(n21673), .A2(n21532), .ZN(n10689) );
  INV_X1 U13624 ( .A(n12589), .ZN(n12207) );
  NAND2_X1 U13625 ( .A1(n12215), .A2(n9715), .ZN(n12201) );
  OAI21_X1 U13626 ( .B1(n11022), .B2(n11541), .A(n11041), .ZN(n11023) );
  INV_X1 U13627 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11533) );
  INV_X1 U13628 ( .A(n11023), .ZN(n11024) );
  AOI22_X1 U13629 ( .A1(n10780), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10775), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10760) );
  NAND2_X1 U13630 ( .A1(n12559), .A2(n12558), .ZN(n12561) );
  INV_X1 U13631 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12506) );
  INV_X1 U13632 ( .A(n11507), .ZN(n11518) );
  BUF_X1 U13633 ( .A(n10780), .Z(n11462) );
  OR2_X1 U13634 ( .A1(n10949), .A2(n10948), .ZN(n11696) );
  NAND2_X1 U13635 ( .A1(n10811), .A2(n10810), .ZN(n10813) );
  AOI22_X1 U13636 ( .A1(n10845), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10943), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10743) );
  INV_X1 U13637 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n12628) );
  OR2_X1 U13638 ( .A1(n12879), .A2(n20981), .ZN(n12250) );
  AOI22_X1 U13639 ( .A1(n9736), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(n9726), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12128) );
  AND2_X1 U13640 ( .A1(n11546), .A2(n11549), .ZN(n11562) );
  NOR2_X1 U13641 ( .A1(n10995), .A2(n10694), .ZN(n10974) );
  NAND2_X1 U13642 ( .A1(n11781), .A2(n14577), .ZN(n11719) );
  AOI22_X1 U13643 ( .A1(n9727), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n9736), .ZN(n12147) );
  AND2_X1 U13644 ( .A1(n12183), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12187) );
  AND4_X1 U13645 ( .A1(n12534), .A2(n12533), .A3(n12532), .A4(n12531), .ZN(
        n12535) );
  OR2_X1 U13646 ( .A1(n13582), .A2(n12378), .ZN(n12398) );
  INV_X1 U13647 ( .A(n16689), .ZN(n12932) );
  INV_X1 U13648 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n22096) );
  AOI22_X1 U13649 ( .A1(n9727), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_10__2__SCAN_IN), .B2(n9736), .ZN(n12169) );
  NAND2_X1 U13650 ( .A1(n21083), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12549) );
  NOR2_X1 U13651 ( .A1(n19646), .A2(n13690), .ZN(n13680) );
  INV_X1 U13652 ( .A(n15420), .ZN(n11409) );
  INV_X1 U13653 ( .A(n11319), .ZN(n11320) );
  INV_X1 U13654 ( .A(n11241), .ZN(n11242) );
  NOR2_X1 U13655 ( .A1(n11100), .A2(n15985), .ZN(n11101) );
  NAND2_X1 U13656 ( .A1(n11053), .A2(n11052), .ZN(n14785) );
  AND2_X1 U13657 ( .A1(n11584), .A2(n11583), .ZN(n14452) );
  AND2_X1 U13658 ( .A1(n11551), .A2(n11550), .ZN(n11564) );
  INV_X1 U13659 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n12638) );
  INV_X1 U13660 ( .A(n16554), .ZN(n12854) );
  INV_X1 U13661 ( .A(n14648), .ZN(n12839) );
  AND2_X1 U13662 ( .A1(n13100), .A2(n13099), .ZN(n16927) );
  INV_X1 U13663 ( .A(n14620), .ZN(n13057) );
  NAND2_X1 U13664 ( .A1(n12929), .A2(n15209), .ZN(n12318) );
  AND2_X1 U13665 ( .A1(n13674), .A2(n19654), .ZN(n13675) );
  INV_X1 U13666 ( .A(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n18688) );
  AND4_X1 U13667 ( .A1(n11932), .A2(n11931), .A3(n11930), .A4(n11929), .ZN(
        n11941) );
  INV_X1 U13668 ( .A(n14567), .ZN(n10803) );
  INV_X1 U13669 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n21202) );
  AND2_X1 U13670 ( .A1(n11605), .A2(n11604), .ZN(n15630) );
  NAND2_X1 U13671 ( .A1(n11452), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11501) );
  OR2_X1 U13672 ( .A1(n15821), .A2(n11455), .ZN(n11431) );
  INV_X1 U13673 ( .A(n15529), .ZN(n11239) );
  INV_X1 U13674 ( .A(n11682), .ZN(n11497) );
  NAND2_X1 U13675 ( .A1(n9823), .A2(n10967), .ZN(n14448) );
  INV_X1 U13676 ( .A(n16203), .ZN(n16198) );
  NAND2_X1 U13677 ( .A1(n10919), .A2(n10918), .ZN(n14540) );
  INV_X1 U13678 ( .A(n16533), .ZN(n13103) );
  INV_X1 U13679 ( .A(n16740), .ZN(n16706) );
  OR2_X1 U13680 ( .A1(n15252), .A2(n15254), .ZN(n15274) );
  INV_X1 U13681 ( .A(n16474), .ZN(n16477) );
  AND2_X1 U13682 ( .A1(n13096), .A2(n13095), .ZN(n16571) );
  INV_X1 U13683 ( .A(n14627), .ZN(n12967) );
  OR2_X1 U13684 ( .A1(n12268), .A2(n12267), .ZN(n12269) );
  AND2_X1 U13685 ( .A1(n13112), .A2(n13111), .ZN(n16484) );
  AND2_X1 U13686 ( .A1(n17075), .A2(n17067), .ZN(n13354) );
  INV_X1 U13687 ( .A(n12627), .ZN(n12946) );
  NAND2_X1 U13688 ( .A1(n13823), .A2(n20834), .ZN(n14277) );
  NAND2_X1 U13689 ( .A1(n20226), .A2(n13848), .ZN(n19560) );
  AND4_X1 U13690 ( .A1(n14125), .A2(n14124), .A3(n14123), .A4(n14122), .ZN(
        n14126) );
  AND4_X1 U13691 ( .A1(n12021), .A2(n12020), .A3(n12019), .A4(n12018), .ZN(
        n12022) );
  OR2_X1 U13692 ( .A1(n17985), .A2(n17690), .ZN(n12053) );
  INV_X1 U13693 ( .A(n19498), .ZN(n19450) );
  INV_X1 U13694 ( .A(n13775), .ZN(n14027) );
  OR2_X1 U13695 ( .A1(n17985), .A2(n14799), .ZN(n11945) );
  INV_X1 U13696 ( .A(n21210), .ZN(n21126) );
  AND2_X1 U13697 ( .A1(n11635), .A2(n11634), .ZN(n15494) );
  INV_X1 U13698 ( .A(n11161), .ZN(n11455) );
  NAND2_X1 U13699 ( .A1(n11040), .A2(n11039), .ZN(n14600) );
  OR2_X1 U13700 ( .A1(n11410), .A2(n15408), .ZN(n11451) );
  NAND2_X1 U13701 ( .A1(n11243), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11279) );
  INV_X1 U13702 ( .A(n10992), .ZN(n11492) );
  INV_X1 U13703 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n15985) );
  NAND2_X1 U13704 ( .A1(n14384), .A2(n11174), .ZN(n10985) );
  AND2_X1 U13705 ( .A1(n11642), .A2(n11641), .ZN(n15444) );
  NOR2_X1 U13706 ( .A1(n16252), .A2(n14247), .ZN(n16207) );
  AND2_X1 U13707 ( .A1(n21415), .A2(n21442), .ZN(n21420) );
  OR2_X1 U13708 ( .A1(n21455), .A2(n21369), .ZN(n16313) );
  INV_X1 U13709 ( .A(n21696), .ZN(n21585) );
  INV_X1 U13710 ( .A(n21375), .ZN(n21568) );
  OR2_X1 U13711 ( .A1(n21673), .A2(n21454), .ZN(n21647) );
  INV_X1 U13712 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21665) );
  AOI221_X1 U13713 ( .B1(n21823), .B2(n21800), .C1(n14378), .C2(n21800), .A(
        P1_STATE2_REG_0__SCAN_IN), .ZN(n16321) );
  INV_X1 U13714 ( .A(n21679), .ZN(n21667) );
  INV_X1 U13715 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n20277) );
  AND3_X1 U13716 ( .A1(n20260), .A2(n20351), .A3(n18130), .ZN(n13330) );
  INV_X1 U13717 ( .A(n15208), .ZN(n16775) );
  AND3_X1 U13718 ( .A1(n12941), .A2(n12940), .A3(n12939), .ZN(n16962) );
  OAI21_X1 U13719 ( .B1(n14731), .B2(n14687), .A(n13611), .ZN(n14425) );
  NOR2_X1 U13720 ( .A1(n10681), .A2(n13235), .ZN(n13236) );
  AND2_X2 U13721 ( .A1(n12270), .A2(n12269), .ZN(n13822) );
  NOR2_X1 U13722 ( .A1(n21047), .A2(n20712), .ZN(n20651) );
  OR2_X1 U13723 ( .A1(n20619), .A2(n20752), .ZN(n20498) );
  AND2_X1 U13724 ( .A1(n20646), .A2(n20645), .ZN(n20653) );
  INV_X1 U13725 ( .A(n20714), .ZN(n20721) );
  NAND3_X1 U13726 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n21042), .A3(n20896), 
        .ZN(n14862) );
  NAND2_X1 U13727 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20896), .ZN(n20450) );
  INV_X1 U13728 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n14742) );
  OR3_X1 U13729 ( .A1(n13695), .A2(n13694), .A3(n13693), .ZN(n13696) );
  NOR2_X1 U13730 ( .A1(n13387), .A2(n13386), .ZN(n13388) );
  NOR2_X1 U13732 ( .A1(n18341), .A2(n10450), .ZN(n18331) );
  NOR2_X1 U13733 ( .A1(n20162), .A2(n18385), .ZN(n18358) );
  AND4_X1 U13734 ( .A1(n11912), .A2(n11911), .A3(n11910), .A4(n11909), .ZN(
        n11922) );
  AND4_X1 U13735 ( .A1(n14142), .A2(n14141), .A3(n14140), .A4(n14139), .ZN(
        n14143) );
  AND4_X1 U13736 ( .A1(n13957), .A2(n13956), .A3(n13955), .A4(n13954), .ZN(
        n13958) );
  AND4_X1 U13737 ( .A1(n12033), .A2(n12032), .A3(n12031), .A4(n12030), .ZN(
        n12044) );
  AND4_X1 U13738 ( .A1(n14154), .A2(n14153), .A3(n14152), .A4(n14151), .ZN(
        n14164) );
  AND2_X1 U13739 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n19450), .ZN(
        n19476) );
  INV_X1 U13740 ( .A(n19702), .ZN(n19703) );
  OR2_X1 U13741 ( .A1(n13792), .A2(n13570), .ZN(n13564) );
  OR2_X1 U13742 ( .A1(n21200), .A2(n15370), .ZN(n15033) );
  XNOR2_X1 U13743 ( .A(n11503), .B(n11674), .ZN(n15035) );
  AND2_X1 U13744 ( .A1(n21820), .A2(n11568), .ZN(n21200) );
  INV_X1 U13745 ( .A(n15704), .ZN(n15697) );
  NOR2_X1 U13746 ( .A1(n15776), .A2(n18147), .ZN(n13438) );
  NAND2_X1 U13747 ( .A1(n13798), .A2(n13800), .ZN(n13422) );
  INV_X1 U13748 ( .A(n14330), .ZN(n21270) );
  INV_X1 U13749 ( .A(n14658), .ZN(n21275) );
  NOR2_X1 U13750 ( .A1(n11034), .A2(n18062), .ZN(n11046) );
  INV_X1 U13751 ( .A(n13800), .ZN(n21099) );
  AND2_X1 U13752 ( .A1(n10659), .A2(n11851), .ZN(n11852) );
  INV_X1 U13753 ( .A(n18077), .ZN(n16221) );
  INV_X1 U13754 ( .A(n21291), .ZN(n18072) );
  INV_X1 U13755 ( .A(n21294), .ZN(n21286) );
  INV_X1 U13756 ( .A(n21293), .ZN(n21282) );
  NAND2_X1 U13757 ( .A1(n13816), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21800) );
  OAI22_X1 U13758 ( .A1(n21316), .A2(n21315), .B1(n21571), .B2(n21450), .ZN(
        n21339) );
  OAI211_X1 U13759 ( .C1(n21316), .C2(n21314), .A(n21313), .B(n21568), .ZN(
        n21340) );
  OAI22_X1 U13760 ( .A1(n21382), .A2(n21381), .B1(n21571), .B2(n21380), .ZN(
        n21406) );
  OAI21_X1 U13761 ( .B1(n21421), .B2(n21418), .A(n21417), .ZN(n21446) );
  INV_X1 U13762 ( .A(n21471), .ZN(n21475) );
  OR2_X1 U13763 ( .A1(n9707), .A2(n14752), .ZN(n21532) );
  INV_X1 U13764 ( .A(n16313), .ZN(n14588) );
  INV_X1 U13765 ( .A(n16323), .ZN(n21520) );
  OAI22_X1 U13766 ( .A1(n21573), .A2(n21572), .B1(n21571), .B2(n21570), .ZN(
        n21605) );
  OR2_X1 U13767 ( .A1(n14614), .A2(n21416), .ZN(n21635) );
  INV_X1 U13768 ( .A(n21529), .ZN(n21534) );
  INV_X1 U13769 ( .A(n21581), .ZN(n21690) );
  INV_X1 U13770 ( .A(n21593), .ZN(n21708) );
  AND2_X1 U13771 ( .A1(n14591), .A2(n14576), .ZN(n21723) );
  INV_X1 U13772 ( .A(n18092), .ZN(n21822) );
  INV_X1 U13773 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n21097) );
  OAI21_X1 U13774 ( .B1(n15367), .B2(n16740), .A(n9807), .ZN(n15368) );
  INV_X1 U13775 ( .A(n16483), .ZN(n16496) );
  INV_X1 U13776 ( .A(n20336), .ZN(n16736) );
  INV_X1 U13777 ( .A(n20292), .ZN(n20344) );
  INV_X1 U13778 ( .A(n20345), .ZN(n20329) );
  OR2_X1 U13779 ( .A1(n13072), .A2(n13071), .ZN(n15057) );
  OR2_X1 U13780 ( .A1(n13020), .A2(n13019), .ZN(n16837) );
  INV_X1 U13781 ( .A(n16840), .ZN(n16830) );
  OR2_X1 U13782 ( .A1(n15089), .A2(n15088), .ZN(n16808) );
  INV_X1 U13783 ( .A(n20389), .ZN(n20373) );
  OR2_X1 U13784 ( .A1(n16938), .A2(n14429), .ZN(n15339) );
  AND2_X1 U13785 ( .A1(n18112), .A2(n13588), .ZN(n18102) );
  INV_X1 U13786 ( .A(n13139), .ZN(n20343) );
  INV_X1 U13787 ( .A(n18112), .ZN(n17214) );
  INV_X1 U13788 ( .A(n13350), .ZN(n17097) );
  INV_X1 U13789 ( .A(n17518), .ZN(n18120) );
  OAI21_X1 U13790 ( .B1(n17561), .B2(n17564), .A(n17560), .ZN(n20455) );
  INV_X1 U13791 ( .A(n20498), .ZN(n21833) );
  OAI21_X1 U13792 ( .B1(n20555), .B2(n20554), .A(n20553), .ZN(n20571) );
  OAI21_X1 U13793 ( .B1(n20584), .B2(n20583), .A(n20582), .ZN(n20607) );
  OR3_X1 U13794 ( .A1(n20624), .A2(n20623), .A3(n20622), .ZN(n20641) );
  INV_X1 U13795 ( .A(n20650), .ZN(n20893) );
  AND2_X1 U13796 ( .A1(n20787), .A2(n20785), .ZN(n20806) );
  NOR2_X2 U13797 ( .A1(n20722), .A2(n20752), .ZN(n20824) );
  AND2_X1 U13798 ( .A1(n20838), .A2(n20833), .ZN(n20863) );
  OAI21_X1 U13799 ( .B1(n17581), .B2(n17584), .A(n17580), .ZN(n20887) );
  INV_X1 U13800 ( .A(n20725), .ZN(n20905) );
  AND2_X1 U13801 ( .A1(READY12_REG_SCAN_IN), .A2(READY21_REG_SCAN_IN), .ZN(
        n20959) );
  AND2_X1 U13802 ( .A1(n14052), .A2(n20107), .ZN(n20230) );
  NAND2_X1 U13803 ( .A1(n13389), .A2(n13388), .ZN(n13390) );
  NAND2_X1 U13804 ( .A1(n18332), .A2(n21874), .ZN(n18326) );
  NAND2_X1 U13805 ( .A1(n18372), .A2(n18368), .ZN(n18365) );
  NAND2_X1 U13806 ( .A1(n18521), .A2(n18513), .ZN(n18512) );
  NOR2_X1 U13807 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n18574), .ZN(n18550) );
  INV_X1 U13808 ( .A(n18522), .ZN(n18596) );
  INV_X1 U13809 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n18802) );
  INV_X1 U13810 ( .A(n18861), .ZN(n17728) );
  NAND2_X1 U13811 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n18896), .ZN(n18895) );
  NAND2_X2 U13812 ( .A1(n13881), .A2(n19654), .ZN(n18902) );
  AND2_X1 U13813 ( .A1(n19348), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n19236) );
  NAND2_X1 U13814 ( .A1(n17798), .A2(n17797), .ZN(n17873) );
  INV_X1 U13815 ( .A(n19204), .ZN(n19254) );
  NAND2_X1 U13816 ( .A1(n19183), .A2(n19082), .ZN(n19344) );
  NAND4_X1 U13817 ( .A1(n14165), .A2(n14164), .A3(n14163), .A4(n14162), .ZN(
        n17942) );
  NAND2_X1 U13818 ( .A1(n19598), .A2(n19587), .ZN(n19605) );
  INV_X1 U13819 ( .A(n17856), .ZN(n19209) );
  INV_X1 U13820 ( .A(n19603), .ZN(n19566) );
  AND2_X1 U13821 ( .A1(n13702), .A2(n20212), .ZN(n19598) );
  NOR2_X1 U13822 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n21986), .ZN(
        n20095) );
  CLKBUF_X1 U13823 ( .A(n19676), .Z(n19744) );
  INV_X1 U13824 ( .A(n19880), .ZN(n19882) );
  INV_X1 U13825 ( .A(n20018), .ZN(n19946) );
  INV_X1 U13826 ( .A(n20006), .ZN(n19969) );
  INV_X2 U13827 ( .A(n19863), .ZN(n20002) );
  INV_X1 U13828 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n22024) );
  NOR2_X1 U13829 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13456), .ZN(n18218)
         );
  INV_X1 U13830 ( .A(n11679), .ZN(n11680) );
  INV_X1 U13831 ( .A(n21209), .ZN(n21143) );
  OR2_X1 U13832 ( .A1(n15035), .A2(n15033), .ZN(n15654) );
  AND2_X1 U13833 ( .A1(n15654), .A2(n15653), .ZN(n21215) );
  INV_X1 U13834 ( .A(n15976), .ZN(n15794) );
  INV_X1 U13835 ( .A(n21220), .ZN(n14599) );
  INV_X1 U13836 ( .A(n21231), .ZN(n21237) );
  OR3_X1 U13837 ( .A1(n18025), .A2(n13751), .A3(n21099), .ZN(n21256) );
  NOR2_X1 U13838 ( .A1(n15373), .A2(n14251), .ZN(n14330) );
  NAND2_X1 U13839 ( .A1(n18061), .A2(n13746), .ZN(n18056) );
  NAND2_X1 U13840 ( .A1(n21105), .A2(n11687), .ZN(n18061) );
  AND2_X1 U13841 ( .A1(n11853), .A2(n11852), .ZN(n11854) );
  OR3_X1 U13842 ( .A1(n21290), .A2(n21278), .A3(n18080), .ZN(n18077) );
  OR2_X2 U13843 ( .A1(n11824), .A2(n11796), .ZN(n21294) );
  INV_X1 U13844 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n21303) );
  OR2_X1 U13845 ( .A1(n21413), .A2(n21454), .ZN(n21362) );
  OR2_X1 U13846 ( .A1(n21413), .A2(n21532), .ZN(n21404) );
  OR2_X1 U13847 ( .A1(n21413), .A2(n21369), .ZN(n21443) );
  OR2_X1 U13848 ( .A1(n21413), .A2(n21410), .ZN(n21471) );
  OR2_X1 U13849 ( .A1(n21455), .A2(n21454), .ZN(n21501) );
  AOI22_X1 U13850 ( .A1(n16286), .A2(n16284), .B1(n16281), .B2(n21379), .ZN(
        n16316) );
  OR2_X1 U13851 ( .A1(n21455), .A2(n21410), .ZN(n16323) );
  NAND2_X1 U13852 ( .A1(n21534), .A2(n16318), .ZN(n21559) );
  NAND2_X1 U13853 ( .A1(n21534), .A2(n21533), .ZN(n21609) );
  NAND2_X1 U13854 ( .A1(n21534), .A2(n14606), .ZN(n21627) );
  NAND2_X1 U13855 ( .A1(n21534), .A2(n14607), .ZN(n21653) );
  AOI21_X1 U13856 ( .B1(n16375), .B2(n16376), .A(n21416), .ZN(n16417) );
  OR2_X1 U13857 ( .A1(n21673), .A2(n21369), .ZN(n21720) );
  NAND2_X1 U13858 ( .A1(n21749), .A2(n21815), .ZN(n21736) );
  NAND2_X1 U13859 ( .A1(n13249), .A2(n14736), .ZN(n16423) );
  INV_X1 U13860 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n20712) );
  AOI21_X1 U13861 ( .B1(n15361), .B2(n20330), .A(n15368), .ZN(n15369) );
  INV_X1 U13862 ( .A(n20330), .ZN(n20341) );
  INV_X1 U13863 ( .A(n17163), .ZN(n17429) );
  NAND2_X1 U13864 ( .A1(n20292), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20339) );
  OR2_X1 U13865 ( .A1(n16423), .A2(n13250), .ZN(n20345) );
  INV_X1 U13866 ( .A(n17320), .ZN(n16791) );
  NAND2_X1 U13867 ( .A1(n16835), .A2(n12905), .ZN(n16840) );
  INV_X1 U13868 ( .A(n16938), .ZN(n16965) );
  AND2_X1 U13869 ( .A1(n16946), .A2(n15339), .ZN(n20393) );
  OR2_X1 U13870 ( .A1(n20417), .A2(n20426), .ZN(n13711) );
  OR2_X1 U13871 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14857), .ZN(n20419) );
  INV_X1 U13872 ( .A(n20417), .ZN(n20428) );
  NAND2_X1 U13873 ( .A1(n13468), .A2(n16419), .ZN(n13625) );
  OR2_X1 U13874 ( .A1(n21087), .A2(n13217), .ZN(n17218) );
  OR2_X1 U13875 ( .A1(n20239), .A2(n15209), .ZN(n17252) );
  NOR2_X1 U13876 ( .A1(n13192), .A2(n13191), .ZN(n13196) );
  INV_X1 U13877 ( .A(n18118), .ZN(n17534) );
  NAND2_X1 U13878 ( .A1(n20714), .A2(n20656), .ZN(n20518) );
  NOR2_X1 U13879 ( .A1(n20523), .A2(n20522), .ZN(n21841) );
  INV_X1 U13880 ( .A(n21836), .ZN(n20575) );
  NAND2_X1 U13881 ( .A1(n20543), .A2(n20835), .ZN(n20599) );
  INV_X1 U13882 ( .A(n20669), .ZN(n20677) );
  AOI21_X1 U13883 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n20710), .A(n20709), 
        .ZN(n20748) );
  INV_X1 U13884 ( .A(n20755), .ZN(n20778) );
  INV_X1 U13885 ( .A(n20779), .ZN(n20810) );
  AOI21_X1 U13886 ( .B1(n14861), .B2(n14860), .A(n14859), .ZN(n20828) );
  AOI22_X1 U13887 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20454), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n20453), .ZN(n20855) );
  AOI211_X2 U13888 ( .C1(n17585), .C2(n17584), .A(n20623), .B(n17583), .ZN(
        n20891) );
  NOR2_X1 U13889 ( .A1(n20898), .A2(n20897), .ZN(n20957) );
  INV_X1 U13890 ( .A(n21040), .ZN(n20958) );
  NAND2_X1 U13891 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18914), .ZN(n20109) );
  INV_X1 U13892 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18807) );
  OR2_X1 U13893 ( .A1(n18902), .A2(n19650), .ZN(n18864) );
  AND2_X1 U13894 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17727), .ZN(n17721) );
  INV_X1 U13895 ( .A(n18902), .ZN(n18907) );
  NOR2_X1 U13896 ( .A1(n18949), .A2(n18895), .ZN(n17746) );
  INV_X1 U13897 ( .A(n14215), .ZN(n17755) );
  OR2_X1 U13898 ( .A1(n18902), .A2(n13964), .ZN(n18913) );
  NAND2_X1 U13899 ( .A1(n18916), .A2(n18915), .ZN(n18971) );
  OR2_X1 U13900 ( .A1(n19342), .A2(n17778), .ZN(n19204) );
  AND2_X1 U13901 ( .A1(n19093), .A2(n19092), .ZN(n19186) );
  INV_X1 U13902 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n19524) );
  INV_X1 U13903 ( .A(n19344), .ZN(n19309) );
  OR2_X1 U13904 ( .A1(n18244), .A2(n18973), .ZN(n19334) );
  OR2_X1 U13905 ( .A1(n19605), .A2(n17778), .ZN(n19505) );
  INV_X1 U13906 ( .A(n19556), .ZN(n19603) );
  INV_X1 U13907 ( .A(n19598), .ZN(n19575) );
  INV_X1 U13908 ( .A(n19723), .ZN(n19718) );
  INV_X1 U13909 ( .A(n19789), .ZN(n19776) );
  INV_X1 U13910 ( .A(n19811), .ZN(n19807) );
  INV_X1 U13911 ( .A(n19835), .ZN(n19833) );
  INV_X1 U13912 ( .A(n20048), .ZN(n20036) );
  INV_X1 U13913 ( .A(n20220), .ZN(n20116) );
  INV_X1 U13914 ( .A(n20197), .ZN(n20117) );
  INV_X1 U13915 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n20137) );
  INV_X1 U13916 ( .A(n18191), .ZN(n18195) );
  NAND2_X1 U13917 ( .A1(n13343), .A2(n13342), .ZN(P2_U2825) );
  NAND2_X1 U13918 ( .A1(n10780), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10693) );
  NAND2_X1 U13919 ( .A1(n10845), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10692) );
  NAND2_X1 U13920 ( .A1(n10775), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n10691) );
  NAND2_X1 U13921 ( .A1(n10846), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n10690) );
  NAND2_X1 U13922 ( .A1(n10871), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10698) );
  INV_X1 U13923 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10694) );
  NAND2_X1 U13924 ( .A1(n10892), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10697) );
  NAND2_X1 U13925 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n10696) );
  NAND2_X1 U13926 ( .A1(n10938), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n10695) );
  AND2_X2 U13927 ( .A1(n10705), .A2(n14351), .ZN(n10727) );
  NAND2_X1 U13928 ( .A1(n10727), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n10704) );
  AND2_X2 U13929 ( .A1(n10706), .A2(n10699), .ZN(n10741) );
  NAND2_X1 U13930 ( .A1(n10741), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n10703) );
  NAND2_X1 U13931 ( .A1(n10943), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n10702) );
  NAND2_X1 U13932 ( .A1(n10756), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10701) );
  NAND2_X1 U13933 ( .A1(n11111), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n10711) );
  NAND2_X1 U13934 ( .A1(n10889), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n10710) );
  NAND2_X1 U13935 ( .A1(n10884), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10709) );
  AND2_X4 U13936 ( .A1(n10707), .A2(n14351), .ZN(n10937) );
  NAND2_X1 U13937 ( .A1(n10937), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10708) );
  AOI22_X1 U13938 ( .A1(n11111), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10871), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10719) );
  AOI22_X1 U13939 ( .A1(n10775), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10938), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10718) );
  AOI22_X1 U13940 ( .A1(n10756), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10943), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10717) );
  NAND4_X1 U13941 ( .A1(n10720), .A2(n10719), .A3(n10718), .A4(n10717), .ZN(
        n10726) );
  AOI22_X1 U13942 ( .A1(n10892), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10846), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10724) );
  AOI22_X1 U13943 ( .A1(n10884), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10876), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10723) );
  AOI22_X1 U13944 ( .A1(n10727), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10741), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10722) );
  AOI22_X1 U13945 ( .A1(n10889), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10937), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10721) );
  NAND4_X1 U13946 ( .A1(n10724), .A2(n10723), .A3(n10722), .A4(n10721), .ZN(
        n10725) );
  INV_X2 U13947 ( .A(n10799), .ZN(n10821) );
  AOI22_X1 U13948 ( .A1(n10780), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10775), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10731) );
  AOI22_X1 U13949 ( .A1(n10741), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10756), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10730) );
  AOI22_X1 U13950 ( .A1(n10727), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10943), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10729) );
  AOI22_X1 U13951 ( .A1(n10845), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10846), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10728) );
  AOI22_X1 U13952 ( .A1(n11111), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10889), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10735) );
  AOI22_X1 U13953 ( .A1(n10884), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10937), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10734) );
  AOI22_X1 U13954 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10871), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10733) );
  AOI22_X1 U13955 ( .A1(n10892), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10938), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10732) );
  AOI22_X1 U13956 ( .A1(n10780), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10727), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10740) );
  AOI22_X1 U13957 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10739) );
  AOI22_X1 U13958 ( .A1(n11111), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10889), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10738) );
  AOI22_X1 U13959 ( .A1(n10884), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10871), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10737) );
  NAND4_X1 U13960 ( .A1(n10740), .A2(n10739), .A3(n10738), .A4(n10737), .ZN(
        n10766) );
  AOI22_X1 U13961 ( .A1(n10937), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10938), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10745) );
  AOI22_X1 U13962 ( .A1(n10741), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10756), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10744) );
  AOI22_X1 U13963 ( .A1(n10775), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10846), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10742) );
  NAND4_X1 U13964 ( .A1(n10745), .A2(n10744), .A3(n10743), .A4(n10742), .ZN(
        n10765) );
  AOI22_X1 U13965 ( .A1(n10780), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10775), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10749) );
  AOI22_X1 U13966 ( .A1(n10741), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10756), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10748) );
  AOI22_X1 U13967 ( .A1(n10727), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10943), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10747) );
  AOI22_X1 U13968 ( .A1(n10845), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10846), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10746) );
  NAND4_X1 U13969 ( .A1(n10749), .A2(n10748), .A3(n10747), .A4(n10746), .ZN(
        n10755) );
  AOI22_X1 U13970 ( .A1(n11111), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10889), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10753) );
  AOI22_X1 U13971 ( .A1(n10884), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10937), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10752) );
  AOI22_X1 U13972 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10871), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10751) );
  AOI22_X1 U13973 ( .A1(n10892), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10938), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10750) );
  NAND4_X1 U13974 ( .A1(n10753), .A2(n10752), .A3(n10751), .A4(n10750), .ZN(
        n10754) );
  AOI22_X1 U13975 ( .A1(n10741), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10756), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10759) );
  AOI22_X1 U13976 ( .A1(n10727), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10943), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10758) );
  AOI22_X1 U13977 ( .A1(n10845), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10846), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10757) );
  AOI22_X1 U13978 ( .A1(n11111), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10889), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10764) );
  AOI22_X1 U13979 ( .A1(n10884), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10937), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10763) );
  AOI22_X1 U13980 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10871), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10762) );
  AOI22_X1 U13981 ( .A1(n10892), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10938), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10761) );
  NAND2_X2 U13982 ( .A1(n10768), .A2(n10767), .ZN(n14577) );
  AOI22_X1 U13983 ( .A1(n11111), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10889), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10774) );
  AOI22_X1 U13984 ( .A1(n10884), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10937), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10773) );
  AOI22_X1 U13985 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10871), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10772) );
  AOI22_X1 U13986 ( .A1(n10892), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10938), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10771) );
  AOI22_X1 U13987 ( .A1(n10780), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10775), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10779) );
  AOI22_X1 U13988 ( .A1(n10741), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10756), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10778) );
  AOI22_X1 U13989 ( .A1(n10727), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10943), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10777) );
  AOI22_X1 U13990 ( .A1(n10845), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10846), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10776) );
  AOI22_X1 U13991 ( .A1(n11111), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10889), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10784) );
  AOI22_X1 U13992 ( .A1(n10884), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10780), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10783) );
  AOI22_X1 U13993 ( .A1(n10845), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10846), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10782) );
  AOI22_X1 U13994 ( .A1(n10727), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10756), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10781) );
  NAND4_X1 U13995 ( .A1(n10784), .A2(n10783), .A3(n10782), .A4(n10781), .ZN(
        n10791) );
  AOI22_X1 U13996 ( .A1(n10741), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10943), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10789) );
  AOI22_X1 U13997 ( .A1(n10775), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10938), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10788) );
  AOI22_X1 U13998 ( .A1(n10937), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10871), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10786) );
  AOI22_X1 U13999 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10785) );
  AND2_X1 U14000 ( .A1(n10786), .A2(n10785), .ZN(n10787) );
  NAND3_X1 U14001 ( .A1(n10789), .A2(n10788), .A3(n10787), .ZN(n10790) );
  OR2_X4 U14002 ( .A1(n10791), .A2(n10790), .ZN(n14561) );
  NAND2_X1 U14003 ( .A1(n11556), .A2(n10663), .ZN(n11792) );
  INV_X1 U14004 ( .A(n14553), .ZN(n11569) );
  INV_X1 U14005 ( .A(n14350), .ZN(n10794) );
  NAND2_X1 U14006 ( .A1(n10792), .A2(n13420), .ZN(n11800) );
  XNOR2_X1 U14007 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n11658) );
  NAND2_X1 U14008 ( .A1(n11555), .A2(n10660), .ZN(n10797) );
  AND2_X4 U14009 ( .A1(n14561), .A2(n9724), .ZN(n14238) );
  NAND2_X1 U14010 ( .A1(n11555), .A2(n14238), .ZN(n11794) );
  NAND4_X1 U14011 ( .A1(n11792), .A2(n11800), .A3(n10797), .A4(n11794), .ZN(
        n10798) );
  NAND2_X1 U14012 ( .A1(n10798), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10812) );
  NAND2_X1 U14013 ( .A1(n10816), .A2(n10799), .ZN(n10800) );
  AND2_X1 U14014 ( .A1(n10800), .A2(n14591), .ZN(n10817) );
  NAND2_X1 U14015 ( .A1(n11684), .A2(n10795), .ZN(n11786) );
  NAND2_X1 U14016 ( .A1(n11786), .A2(n16270), .ZN(n10827) );
  NAND2_X1 U14017 ( .A1(n11661), .A2(n9724), .ZN(n21825) );
  NAND2_X1 U14018 ( .A1(n11808), .A2(n15028), .ZN(n10805) );
  NAND2_X1 U14019 ( .A1(n14557), .A2(n9724), .ZN(n11807) );
  OAI211_X1 U14020 ( .C1(n21825), .C2(n10795), .A(n10805), .B(n10804), .ZN(
        n10820) );
  NOR2_X1 U14021 ( .A1(n10820), .A2(n10794), .ZN(n10807) );
  NAND2_X1 U14022 ( .A1(n10806), .A2(n13570), .ZN(n10825) );
  NAND3_X1 U14023 ( .A1(n10827), .A2(n10807), .A3(n10825), .ZN(n11819) );
  NAND2_X1 U14024 ( .A1(n11819), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10808) );
  NAND2_X1 U14025 ( .A1(n10834), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10811) );
  NAND2_X1 U14026 ( .A1(n21665), .A2(n21561), .ZN(n21453) );
  NAND2_X1 U14027 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n10914) );
  NAND2_X1 U14028 ( .A1(n21453), .A2(n10914), .ZN(n16324) );
  OR2_X1 U14029 ( .A1(n18034), .A2(n21665), .ZN(n10831) );
  OAI21_X1 U14030 ( .B1(n11686), .B2(n16324), .A(n10831), .ZN(n10809) );
  INV_X1 U14031 ( .A(n10809), .ZN(n10810) );
  INV_X1 U14032 ( .A(n10857), .ZN(n10829) );
  NAND2_X1 U14033 ( .A1(n10834), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10815) );
  MUX2_X1 U14034 ( .A(n18034), .B(n11686), .S(n21561), .Z(n10814) );
  AND2_X1 U14035 ( .A1(n13562), .A2(n11654), .ZN(n15374) );
  OAI21_X1 U14036 ( .B1(n10816), .B2(n10799), .A(n14553), .ZN(n10819) );
  INV_X1 U14037 ( .A(n10817), .ZN(n10818) );
  AOI22_X1 U14038 ( .A1(n15374), .A2(n10819), .B1(n10818), .B2(n11798), .ZN(
        n10824) );
  INV_X1 U14039 ( .A(n10820), .ZN(n10823) );
  INV_X1 U14040 ( .A(n18087), .ZN(n21802) );
  NOR2_X1 U14041 ( .A1(n21802), .A2(n21733), .ZN(n10822) );
  NAND2_X1 U14042 ( .A1(n10794), .A2(n10821), .ZN(n11816) );
  OAI211_X1 U14043 ( .C1(n10827), .C2(n11661), .A(n10826), .B(n10825), .ZN(
        n10990) );
  NAND2_X1 U14044 ( .A1(n10831), .A2(n10830), .ZN(n10832) );
  NAND2_X1 U14045 ( .A1(n10833), .A2(n10832), .ZN(n10838) );
  NOR2_X1 U14046 ( .A1(n18034), .A2(n21306), .ZN(n10835) );
  INV_X1 U14047 ( .A(n11686), .ZN(n10917) );
  XNOR2_X1 U14048 ( .A(n10914), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n14759) );
  NAND2_X1 U14049 ( .A1(n10917), .A2(n14759), .ZN(n10837) );
  NAND2_X1 U14050 ( .A1(n10839), .A2(n10837), .ZN(n10836) );
  NAND4_X1 U14051 ( .A1(n10859), .A2(n10839), .A3(n10838), .A4(n10837), .ZN(
        n10840) );
  INV_X1 U14052 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10853) );
  AOI22_X1 U14053 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11393), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10844) );
  AOI22_X1 U14054 ( .A1(n10936), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10870), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10843) );
  AOI22_X1 U14055 ( .A1(n10890), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10871), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10842) );
  AOI22_X1 U14056 ( .A1(n11435), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11324), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10841) );
  NAND4_X1 U14057 ( .A1(n10844), .A2(n10843), .A3(n10842), .A4(n10841), .ZN(
        n10852) );
  AOI22_X1 U14058 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11269), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10850) );
  AOI22_X1 U14059 ( .A1(n10741), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10849) );
  AOI22_X1 U14060 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10848) );
  INV_X1 U14061 ( .A(n10846), .ZN(n10877) );
  AOI22_X1 U14062 ( .A1(n11335), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10847) );
  NAND4_X1 U14063 ( .A1(n10850), .A2(n10849), .A3(n10848), .A4(n10847), .ZN(
        n10851) );
  OAI22_X1 U14064 ( .A1(n11541), .A2(n10853), .B1(n11711), .B2(n10920), .ZN(
        n10855) );
  NOR2_X1 U14065 ( .A1(n11711), .A2(n10921), .ZN(n10854) );
  XNOR2_X1 U14066 ( .A(n10855), .B(n10854), .ZN(n10856) );
  AOI22_X1 U14067 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10870), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10863) );
  AOI22_X1 U14068 ( .A1(n11435), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11462), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10862) );
  AOI22_X1 U14069 ( .A1(n10845), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11413), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10861) );
  AOI22_X1 U14070 ( .A1(n10741), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10860) );
  NAND4_X1 U14071 ( .A1(n10863), .A2(n10862), .A3(n10861), .A4(n10860), .ZN(
        n10869) );
  AOI22_X1 U14072 ( .A1(n10936), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11393), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10867) );
  AOI22_X1 U14073 ( .A1(n10890), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10871), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10866) );
  AOI22_X1 U14074 ( .A1(n11269), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10938), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10865) );
  AOI22_X1 U14075 ( .A1(n10891), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10864) );
  NAND4_X1 U14076 ( .A1(n10867), .A2(n10866), .A3(n10865), .A4(n10864), .ZN(
        n10868) );
  BUF_X1 U14077 ( .A(n10889), .Z(n11393) );
  BUF_X1 U14078 ( .A(n10937), .Z(n10870) );
  AOI22_X1 U14079 ( .A1(n11393), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10870), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10875) );
  AOI22_X1 U14080 ( .A1(n10727), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11412), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10874) );
  AOI22_X1 U14081 ( .A1(n11435), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10871), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10873) );
  AOI22_X1 U14082 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10938), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10872) );
  NAND4_X1 U14083 ( .A1(n10875), .A2(n10874), .A3(n10873), .A4(n10872), .ZN(
        n10883) );
  AOI22_X1 U14084 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10936), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10881) );
  BUF_X1 U14085 ( .A(n10876), .Z(n10890) );
  AOI22_X1 U14086 ( .A1(n10890), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11269), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10880) );
  AOI22_X1 U14087 ( .A1(n10845), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10879) );
  AOI22_X1 U14088 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10878) );
  NAND4_X1 U14089 ( .A1(n10881), .A2(n10880), .A3(n10879), .A4(n10878), .ZN(
        n10882) );
  AOI22_X1 U14090 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10870), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10888) );
  AOI22_X1 U14091 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11335), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10887) );
  AOI22_X1 U14092 ( .A1(n10936), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10871), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10886) );
  AOI22_X1 U14093 ( .A1(n11269), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10938), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10885) );
  NAND4_X1 U14094 ( .A1(n10888), .A2(n10887), .A3(n10886), .A4(n10885), .ZN(
        n10899) );
  AOI22_X1 U14095 ( .A1(n11393), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10890), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10897) );
  BUF_X1 U14096 ( .A(n10943), .Z(n10891) );
  AOI22_X1 U14097 ( .A1(n10727), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10896) );
  AOI22_X1 U14098 ( .A1(n10741), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10895) );
  AOI22_X1 U14099 ( .A1(n11435), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10894) );
  NAND4_X1 U14100 ( .A1(n10897), .A2(n10896), .A3(n10895), .A4(n10894), .ZN(
        n10898) );
  XNOR2_X1 U14101 ( .A(n11755), .B(n11724), .ZN(n10900) );
  INV_X1 U14102 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10903) );
  AOI21_X1 U14103 ( .B1(n13570), .B2(n11724), .A(n21733), .ZN(n10902) );
  NAND2_X1 U14104 ( .A1(n10795), .A2(n11755), .ZN(n10901) );
  NAND2_X1 U14105 ( .A1(n10987), .A2(n10986), .ZN(n10905) );
  NAND2_X1 U14106 ( .A1(n10906), .A2(n11755), .ZN(n10904) );
  INV_X1 U14107 ( .A(n11755), .ZN(n11746) );
  NAND2_X1 U14108 ( .A1(n10906), .A2(n11746), .ZN(n10909) );
  NAND2_X1 U14109 ( .A1(n11509), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10908) );
  NAND2_X1 U14110 ( .A1(n10078), .A2(n11717), .ZN(n10907) );
  INV_X1 U14111 ( .A(n10910), .ZN(n10911) );
  NAND2_X1 U14112 ( .A1(n10834), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10919) );
  OAI21_X1 U14113 ( .B1(n10914), .B2(n21306), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10916) );
  INV_X1 U14114 ( .A(n10914), .ZN(n21661) );
  NAND2_X1 U14115 ( .A1(n11533), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n21480) );
  INV_X1 U14116 ( .A(n21480), .ZN(n10915) );
  NAND2_X1 U14117 ( .A1(n21661), .A2(n10915), .ZN(n14585) );
  NAND2_X1 U14118 ( .A1(n10916), .A2(n14585), .ZN(n21312) );
  INV_X1 U14119 ( .A(n18034), .ZN(n18028) );
  AOI22_X1 U14120 ( .A1(n10917), .A2(n21312), .B1(n18028), .B2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10918) );
  INV_X1 U14121 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10933) );
  AOI22_X1 U14122 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11393), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10925) );
  AOI22_X1 U14123 ( .A1(n10936), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10870), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10924) );
  AOI22_X1 U14124 ( .A1(n10890), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11434), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10923) );
  AOI22_X1 U14125 ( .A1(n11435), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11324), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10922) );
  NAND4_X1 U14126 ( .A1(n10925), .A2(n10924), .A3(n10923), .A4(n10922), .ZN(
        n10931) );
  INV_X1 U14127 ( .A(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n22117) );
  AOI22_X1 U14128 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11269), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10929) );
  AOI22_X1 U14129 ( .A1(n10741), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10928) );
  AOI22_X1 U14130 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10927) );
  AOI22_X1 U14131 ( .A1(n11335), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10926) );
  NAND4_X1 U14132 ( .A1(n10929), .A2(n10928), .A3(n10927), .A4(n10926), .ZN(
        n10930) );
  NAND2_X1 U14133 ( .A1(n11552), .A2(n11700), .ZN(n10932) );
  OAI21_X1 U14134 ( .B1(n10933), .B2(n11541), .A(n10932), .ZN(n10934) );
  AOI22_X1 U14135 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11393), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10942) );
  AOI22_X1 U14136 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n10936), .B1(
        n10870), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10941) );
  AOI22_X1 U14137 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10890), .B1(
        n11434), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10940) );
  AOI22_X1 U14138 ( .A1(n11435), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11324), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10939) );
  NAND4_X1 U14139 ( .A1(n10942), .A2(n10941), .A3(n10940), .A4(n10939), .ZN(
        n10949) );
  AOI22_X1 U14140 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n11462), .B1(
        n11269), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10947) );
  AOI22_X1 U14141 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11412), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10946) );
  AOI22_X1 U14142 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n11413), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10945) );
  AOI22_X1 U14143 ( .A1(n11335), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10944) );
  NAND4_X1 U14144 ( .A1(n10947), .A2(n10946), .A3(n10945), .A4(n10944), .ZN(
        n10948) );
  NAND2_X1 U14145 ( .A1(n11552), .A2(n11696), .ZN(n10951) );
  NAND2_X1 U14146 ( .A1(n11509), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10950) );
  NAND2_X1 U14147 ( .A1(n10961), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11034) );
  OAI21_X1 U14148 ( .B1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n10961), .A(
        n11034), .ZN(n21194) );
  NAND2_X1 U14149 ( .A1(n10792), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10995) );
  INV_X1 U14150 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18089) );
  OAI21_X1 U14151 ( .B1(n21528), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n10952), .ZN(n10954) );
  NAND2_X1 U14152 ( .A1(n10992), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n10953) );
  OAI211_X1 U14153 ( .C1(n10995), .C2(n18089), .A(n10954), .B(n10953), .ZN(
        n10955) );
  OAI21_X1 U14154 ( .B1(n11455), .B2(n21194), .A(n10955), .ZN(n10956) );
  NAND2_X1 U14155 ( .A1(n10957), .A2(n10958), .ZN(n14391) );
  NAND2_X1 U14156 ( .A1(n10959), .A2(n14391), .ZN(n14392) );
  INV_X1 U14157 ( .A(n10960), .ZN(n10963) );
  INV_X1 U14158 ( .A(n10961), .ZN(n10962) );
  OAI21_X1 U14159 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n10963), .A(
        n10962), .ZN(n21216) );
  AOI22_X1 U14160 ( .A1(n11497), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n11278), .B2(n21216), .ZN(n10965) );
  NAND2_X1 U14161 ( .A1(n10992), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n10964) );
  OAI211_X1 U14162 ( .C1(n10995), .C2(n14352), .A(n10965), .B(n10964), .ZN(
        n10966) );
  INV_X1 U14163 ( .A(n10966), .ZN(n10967) );
  NAND2_X1 U14164 ( .A1(n14512), .A2(n14448), .ZN(n10999) );
  INV_X1 U14165 ( .A(n9702), .ZN(n10970) );
  XNOR2_X1 U14166 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n15662) );
  NAND2_X1 U14167 ( .A1(n15662), .A2(n11278), .ZN(n10971) );
  NAND2_X1 U14168 ( .A1(n10971), .A2(n11682), .ZN(n10972) );
  AOI21_X1 U14169 ( .B1(n10992), .B2(P1_EAX_REG_2__SCAN_IN), .A(n10972), .ZN(
        n10973) );
  INV_X1 U14170 ( .A(n10973), .ZN(n10975) );
  NOR2_X1 U14171 ( .A1(n10975), .A2(n10974), .ZN(n10976) );
  NAND2_X1 U14172 ( .A1(n10977), .A2(n10976), .ZN(n14341) );
  NAND2_X1 U14173 ( .A1(n10992), .A2(P1_EAX_REG_1__SCAN_IN), .ZN(n10982) );
  NAND2_X1 U14174 ( .A1(n10952), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10981) );
  OAI211_X1 U14175 ( .C1(n10995), .C2(n10830), .A(n10982), .B(n10981), .ZN(
        n10983) );
  INV_X1 U14176 ( .A(n10983), .ZN(n10984) );
  NAND2_X1 U14177 ( .A1(n10985), .A2(n10984), .ZN(n14058) );
  NAND2_X1 U14178 ( .A1(n14752), .A2(n10821), .ZN(n10988) );
  NAND2_X1 U14179 ( .A1(n10988), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13738) );
  INV_X1 U14180 ( .A(n10990), .ZN(n10991) );
  XNOR2_X1 U14181 ( .A(n10989), .B(n10991), .ZN(n14542) );
  NAND2_X1 U14182 ( .A1(n10952), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10994) );
  NAND2_X1 U14183 ( .A1(n10992), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n10993) );
  OAI211_X1 U14184 ( .C1(n10995), .C2(n10144), .A(n10994), .B(n10993), .ZN(
        n10996) );
  AOI21_X1 U14185 ( .B1(n14542), .B2(n11174), .A(n10996), .ZN(n13739) );
  OR2_X1 U14186 ( .A1(n13738), .A2(n13739), .ZN(n13740) );
  NAND2_X1 U14187 ( .A1(n13739), .A2(n11278), .ZN(n10997) );
  NAND2_X1 U14188 ( .A1(n13740), .A2(n10997), .ZN(n14057) );
  NAND2_X1 U14189 ( .A1(n14058), .A2(n14057), .ZN(n14056) );
  INV_X1 U14190 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n15658) );
  OR2_X1 U14191 ( .A1(n11682), .A2(n15658), .ZN(n14340) );
  NAND2_X1 U14192 ( .A1(n14056), .A2(n14340), .ZN(n10998) );
  NAND2_X1 U14193 ( .A1(n14341), .A2(n10998), .ZN(n14447) );
  AOI22_X1 U14194 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11393), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11003) );
  AOI22_X1 U14195 ( .A1(n10936), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10870), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11002) );
  AOI22_X1 U14196 ( .A1(n10890), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11434), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11001) );
  INV_X1 U14197 ( .A(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n21894) );
  AOI22_X1 U14198 ( .A1(n11435), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11324), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11000) );
  NAND4_X1 U14199 ( .A1(n11003), .A2(n11002), .A3(n11001), .A4(n11000), .ZN(
        n11009) );
  AOI22_X1 U14200 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11269), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11007) );
  AOI22_X1 U14201 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11006) );
  AOI22_X1 U14202 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11005) );
  AOI22_X1 U14203 ( .A1(n11335), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11004) );
  NAND4_X1 U14204 ( .A1(n11007), .A2(n11006), .A3(n11005), .A4(n11004), .ZN(
        n11008) );
  NAND2_X1 U14205 ( .A1(n11552), .A2(n11740), .ZN(n11011) );
  NAND2_X1 U14206 ( .A1(n11509), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11010) );
  INV_X1 U14207 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11022) );
  AOI22_X1 U14208 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11393), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11015) );
  AOI22_X1 U14209 ( .A1(n10936), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10870), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11014) );
  AOI22_X1 U14210 ( .A1(n10890), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11434), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11013) );
  AOI22_X1 U14211 ( .A1(n11435), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11324), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11012) );
  NAND4_X1 U14212 ( .A1(n11015), .A2(n11014), .A3(n11013), .A4(n11012), .ZN(
        n11021) );
  AOI22_X1 U14213 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11269), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11019) );
  AOI22_X1 U14214 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11018) );
  AOI22_X1 U14215 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11017) );
  AOI22_X1 U14216 ( .A1(n11335), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11016) );
  NAND4_X1 U14217 ( .A1(n11019), .A2(n11018), .A3(n11017), .A4(n11016), .ZN(
        n11020) );
  NAND2_X1 U14218 ( .A1(n11552), .A2(n11750), .ZN(n11041) );
  NAND2_X1 U14219 ( .A1(n11738), .A2(n11174), .ZN(n11029) );
  INV_X1 U14220 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11026) );
  XNOR2_X1 U14221 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B(n11046), .ZN(
        n21172) );
  NAND2_X1 U14222 ( .A1(n21172), .A2(n11278), .ZN(n11025) );
  OAI21_X1 U14223 ( .B1(n11026), .B2(n11682), .A(n11025), .ZN(n11027) );
  AOI21_X1 U14224 ( .B1(n10992), .B2(P1_EAX_REG_6__SCAN_IN), .A(n11027), .ZN(
        n11028) );
  NAND2_X1 U14225 ( .A1(n11029), .A2(n11028), .ZN(n14827) );
  NAND2_X1 U14226 ( .A1(n11032), .A2(n11031), .ZN(n11694) );
  INV_X1 U14227 ( .A(n11694), .ZN(n11033) );
  NAND2_X1 U14228 ( .A1(n11033), .A2(n11174), .ZN(n11040) );
  INV_X1 U14229 ( .A(n11034), .ZN(n11036) );
  INV_X1 U14230 ( .A(n11046), .ZN(n11035) );
  OAI21_X1 U14231 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n11036), .A(
        n11035), .ZN(n21182) );
  NAND2_X1 U14232 ( .A1(n21182), .A2(n11278), .ZN(n11037) );
  OAI21_X1 U14233 ( .B1(n18062), .B2(n11682), .A(n11037), .ZN(n11038) );
  AOI21_X1 U14234 ( .B1(n10992), .B2(P1_EAX_REG_5__SCAN_IN), .A(n11038), .ZN(
        n11039) );
  INV_X1 U14235 ( .A(n11041), .ZN(n11042) );
  INV_X1 U14236 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11044) );
  NAND2_X1 U14237 ( .A1(n11552), .A2(n11755), .ZN(n11043) );
  OAI21_X1 U14238 ( .B1(n11044), .B2(n11541), .A(n11043), .ZN(n11045) );
  NAND2_X1 U14239 ( .A1(n11754), .A2(n11174), .ZN(n11053) );
  INV_X1 U14240 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n21154) );
  INV_X1 U14241 ( .A(n11077), .ZN(n11049) );
  NAND2_X1 U14242 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n11046), .ZN(
        n11047) );
  NAND2_X1 U14243 ( .A1(n21154), .A2(n11047), .ZN(n11048) );
  NAND2_X1 U14244 ( .A1(n11049), .A2(n11048), .ZN(n21162) );
  NAND2_X1 U14245 ( .A1(n21162), .A2(n11161), .ZN(n11050) );
  OAI21_X1 U14246 ( .B1(n21154), .B2(n11682), .A(n11050), .ZN(n11051) );
  AOI21_X1 U14247 ( .B1(n10992), .B2(P1_EAX_REG_7__SCAN_IN), .A(n11051), .ZN(
        n11052) );
  AOI22_X1 U14248 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10936), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11057) );
  AOI22_X1 U14249 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11434), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11056) );
  AOI22_X1 U14250 ( .A1(n11335), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11412), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11055) );
  AOI22_X1 U14251 ( .A1(n10780), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11269), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11054) );
  NAND4_X1 U14252 ( .A1(n11057), .A2(n11056), .A3(n11055), .A4(n11054), .ZN(
        n11063) );
  AOI22_X1 U14253 ( .A1(n11393), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10937), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11061) );
  AOI22_X1 U14254 ( .A1(n11435), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11324), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11060) );
  AOI22_X1 U14255 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11059) );
  AOI22_X1 U14256 ( .A1(n10943), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11058) );
  NAND4_X1 U14257 ( .A1(n11061), .A2(n11060), .A3(n11059), .A4(n11058), .ZN(
        n11062) );
  OAI21_X1 U14258 ( .B1(n11063), .B2(n11062), .A(n11174), .ZN(n11066) );
  XNOR2_X1 U14259 ( .A(n11077), .B(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n21145) );
  AOI22_X1 U14260 ( .A1(n21145), .A2(n11161), .B1(n11497), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11065) );
  NAND2_X1 U14261 ( .A1(n10992), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11064) );
  AOI22_X1 U14262 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10889), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11070) );
  AOI22_X1 U14263 ( .A1(n10936), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10937), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11069) );
  AOI22_X1 U14264 ( .A1(n11335), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11434), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11068) );
  AOI22_X1 U14265 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11067) );
  NAND4_X1 U14266 ( .A1(n11070), .A2(n11069), .A3(n11068), .A4(n11067), .ZN(
        n11076) );
  AOI22_X1 U14267 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11435), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11074) );
  AOI22_X1 U14268 ( .A1(n11269), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11324), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11073) );
  AOI22_X1 U14269 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11072) );
  AOI22_X1 U14270 ( .A1(n10780), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10846), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11071) );
  NAND4_X1 U14271 ( .A1(n11074), .A2(n11073), .A3(n11072), .A4(n11071), .ZN(
        n11075) );
  NOR2_X1 U14272 ( .A1(n11076), .A2(n11075), .ZN(n11081) );
  XOR2_X1 U14273 ( .A(n21130), .B(n11093), .Z(n21134) );
  INV_X1 U14274 ( .A(n21134), .ZN(n11078) );
  AOI22_X1 U14275 ( .A1(n11497), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(
        n11278), .B2(n11078), .ZN(n11080) );
  NAND2_X1 U14276 ( .A1(n10992), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11079) );
  OAI211_X1 U14277 ( .C1(n11082), .C2(n11081), .A(n11080), .B(n11079), .ZN(
        n14846) );
  AOI22_X1 U14278 ( .A1(n10889), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10890), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11086) );
  AOI22_X1 U14279 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11412), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11085) );
  AOI22_X1 U14280 ( .A1(n11435), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11269), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11084) );
  AOI22_X1 U14281 ( .A1(n10780), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11083) );
  NAND4_X1 U14282 ( .A1(n11086), .A2(n11085), .A3(n11084), .A4(n11083), .ZN(
        n11092) );
  AOI22_X1 U14283 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10937), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11090) );
  AOI22_X1 U14284 ( .A1(n10936), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11434), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11089) );
  AOI22_X1 U14285 ( .A1(n11335), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11324), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11088) );
  AOI22_X1 U14286 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10943), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11087) );
  NAND4_X1 U14287 ( .A1(n11090), .A2(n11089), .A3(n11088), .A4(n11087), .ZN(
        n11091) );
  OR2_X1 U14288 ( .A1(n11092), .A2(n11091), .ZN(n11095) );
  XNOR2_X1 U14289 ( .A(n11100), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15987) );
  NOR2_X1 U14290 ( .A1(n15987), .A2(n11455), .ZN(n11094) );
  AOI21_X1 U14291 ( .B1(n11174), .B2(n11095), .A(n11094), .ZN(n11098) );
  NOR2_X1 U14292 ( .A1(n11682), .A2(n15985), .ZN(n11096) );
  AOI21_X1 U14293 ( .B1(n10992), .B2(P1_EAX_REG_10__SCAN_IN), .A(n11096), .ZN(
        n11097) );
  INV_X1 U14294 ( .A(n14880), .ZN(n11099) );
  NAND2_X1 U14295 ( .A1(n10992), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n11106) );
  INV_X1 U14296 ( .A(n11101), .ZN(n11103) );
  INV_X1 U14297 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11102) );
  NAND2_X1 U14298 ( .A1(n11103), .A2(n11102), .ZN(n11104) );
  NAND2_X1 U14299 ( .A1(n11177), .A2(n11104), .ZN(n15974) );
  AOI22_X1 U14300 ( .A1(n15974), .A2(n11278), .B1(n11497), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11105) );
  NAND2_X1 U14301 ( .A1(n11106), .A2(n11105), .ZN(n15565) );
  AOI22_X1 U14302 ( .A1(n10936), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10870), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11110) );
  AOI22_X1 U14303 ( .A1(n11435), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11434), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11109) );
  AOI22_X1 U14304 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11324), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11108) );
  AOI22_X1 U14305 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11107) );
  NAND4_X1 U14306 ( .A1(n11110), .A2(n11109), .A3(n11108), .A4(n11107), .ZN(
        n11117) );
  AOI22_X1 U14307 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11393), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11115) );
  AOI22_X1 U14308 ( .A1(n10890), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11269), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11114) );
  AOI22_X1 U14309 ( .A1(n11335), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11113) );
  AOI22_X1 U14310 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11112) );
  NAND4_X1 U14311 ( .A1(n11115), .A2(n11114), .A3(n11113), .A4(n11112), .ZN(
        n11116) );
  OR2_X1 U14312 ( .A1(n11117), .A2(n11116), .ZN(n11118) );
  AND2_X1 U14313 ( .A1(n11174), .A2(n11118), .ZN(n15595) );
  OR2_X1 U14314 ( .A1(n15565), .A2(n15595), .ZN(n11134) );
  AOI22_X1 U14315 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11269), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11122) );
  AOI22_X1 U14316 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n11435), .B1(
        n11324), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11121) );
  AOI22_X1 U14317 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n11412), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11120) );
  AOI22_X1 U14318 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n11335), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11119) );
  NAND4_X1 U14319 ( .A1(n11122), .A2(n11121), .A3(n11120), .A4(n11119), .ZN(
        n11128) );
  AOI22_X1 U14320 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11393), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11126) );
  AOI22_X1 U14321 ( .A1(n10936), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10870), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11125) );
  AOI22_X1 U14322 ( .A1(n10890), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11434), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11124) );
  AOI22_X1 U14323 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11123) );
  NAND4_X1 U14324 ( .A1(n11126), .A2(n11125), .A3(n11124), .A4(n11123), .ZN(
        n11127) );
  OAI21_X1 U14325 ( .B1(n11128), .B2(n11127), .A(n11174), .ZN(n11133) );
  NAND2_X1 U14326 ( .A1(n10992), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n11132) );
  INV_X1 U14327 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11129) );
  XNOR2_X1 U14328 ( .A(n11177), .B(n11129), .ZN(n15963) );
  NAND2_X1 U14329 ( .A1(n15963), .A2(n11278), .ZN(n11131) );
  NAND2_X1 U14330 ( .A1(n11497), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11130) );
  NAND4_X1 U14331 ( .A1(n11133), .A2(n11132), .A3(n11131), .A4(n11130), .ZN(
        n15596) );
  AND2_X1 U14332 ( .A1(n11134), .A2(n15596), .ZN(n11185) );
  INV_X1 U14333 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n21228) );
  NAND2_X1 U14334 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11135) );
  INV_X1 U14335 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11160) );
  NOR2_X1 U14336 ( .A1(n11200), .A2(n11160), .ZN(n11136) );
  XNOR2_X1 U14337 ( .A(n11136), .B(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15934) );
  NAND2_X1 U14338 ( .A1(n15934), .A2(n11278), .ZN(n11149) );
  AOI22_X1 U14339 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11393), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11140) );
  AOI22_X1 U14340 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11335), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11139) );
  AOI22_X1 U14341 ( .A1(n10936), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11434), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11138) );
  AOI22_X1 U14342 ( .A1(n11269), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11324), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11137) );
  NAND4_X1 U14343 ( .A1(n11140), .A2(n11139), .A3(n11138), .A4(n11137), .ZN(
        n11146) );
  AOI22_X1 U14344 ( .A1(n10870), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10890), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11144) );
  AOI22_X1 U14345 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11143) );
  AOI22_X1 U14346 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11142) );
  AOI22_X1 U14347 ( .A1(n11435), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11141) );
  NAND4_X1 U14348 ( .A1(n11144), .A2(n11143), .A3(n11142), .A4(n11141), .ZN(
        n11145) );
  OR2_X1 U14349 ( .A1(n11146), .A2(n11145), .ZN(n11147) );
  AOI22_X1 U14350 ( .A1(n11174), .A2(n11147), .B1(n11497), .B2(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11148) );
  OAI211_X1 U14351 ( .C1(n11492), .C2(n21228), .A(n11149), .B(n11148), .ZN(
        n15569) );
  AOI22_X1 U14352 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10890), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11153) );
  AOI22_X1 U14353 ( .A1(n11435), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11462), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11152) );
  AOI22_X1 U14354 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11412), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11151) );
  AOI22_X1 U14355 ( .A1(n11335), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11150) );
  NAND4_X1 U14356 ( .A1(n11153), .A2(n11152), .A3(n11151), .A4(n11150), .ZN(
        n11159) );
  AOI22_X1 U14357 ( .A1(n11393), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10870), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11157) );
  AOI22_X1 U14358 ( .A1(n10936), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11434), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11156) );
  AOI22_X1 U14359 ( .A1(n11269), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11324), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11155) );
  AOI22_X1 U14360 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10943), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11154) );
  NAND4_X1 U14361 ( .A1(n11157), .A2(n11156), .A3(n11155), .A4(n11154), .ZN(
        n11158) );
  OAI21_X1 U14362 ( .B1(n11159), .B2(n11158), .A(n11174), .ZN(n11165) );
  XNOR2_X1 U14363 ( .A(n11200), .B(n11160), .ZN(n15946) );
  NAND2_X1 U14364 ( .A1(n15946), .A2(n11161), .ZN(n11164) );
  NAND2_X1 U14365 ( .A1(n10992), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n11163) );
  NAND2_X1 U14366 ( .A1(n11497), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11162) );
  NAND4_X1 U14367 ( .A1(n11165), .A2(n11164), .A3(n11163), .A4(n11162), .ZN(
        n15568) );
  AOI22_X1 U14368 ( .A1(n10936), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10870), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11169) );
  AOI22_X1 U14369 ( .A1(n11335), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11412), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11168) );
  AOI22_X1 U14370 ( .A1(n11434), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11324), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11167) );
  AOI22_X1 U14371 ( .A1(n11269), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11166) );
  NAND4_X1 U14372 ( .A1(n11169), .A2(n11168), .A3(n11167), .A4(n11166), .ZN(
        n11176) );
  AOI22_X1 U14373 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11393), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11173) );
  AOI22_X1 U14374 ( .A1(n10890), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11435), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11172) );
  AOI22_X1 U14375 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11171) );
  AOI22_X1 U14376 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11170) );
  NAND4_X1 U14377 ( .A1(n11173), .A2(n11172), .A3(n11171), .A4(n11170), .ZN(
        n11175) );
  OAI21_X1 U14378 ( .B1(n11176), .B2(n11175), .A(n11174), .ZN(n11184) );
  INV_X1 U14379 ( .A(n11177), .ZN(n11178) );
  NAND2_X1 U14380 ( .A1(n11178), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11180) );
  INV_X1 U14381 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11179) );
  XNOR2_X1 U14382 ( .A(n11180), .B(n11179), .ZN(n15950) );
  NAND2_X1 U14383 ( .A1(n15950), .A2(n11161), .ZN(n11183) );
  NAND2_X1 U14384 ( .A1(n10992), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n11182) );
  NAND2_X1 U14385 ( .A1(n11497), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11181) );
  NAND4_X1 U14386 ( .A1(n11184), .A2(n11183), .A3(n11182), .A4(n11181), .ZN(
        n15598) );
  INV_X1 U14387 ( .A(n16270), .ZN(n11186) );
  AOI22_X1 U14388 ( .A1(n11393), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10870), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11190) );
  AOI22_X1 U14389 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11412), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11189) );
  AOI22_X1 U14390 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11434), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11188) );
  AOI22_X1 U14391 ( .A1(n11335), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11324), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11187) );
  NAND4_X1 U14392 ( .A1(n11190), .A2(n11189), .A3(n11188), .A4(n11187), .ZN(
        n11196) );
  AOI22_X1 U14393 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10936), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11194) );
  AOI22_X1 U14394 ( .A1(n11435), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11269), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11193) );
  AOI22_X1 U14395 ( .A1(n10780), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11192) );
  AOI22_X1 U14396 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11191) );
  NAND4_X1 U14397 ( .A1(n11194), .A2(n11193), .A3(n11192), .A4(n11191), .ZN(
        n11195) );
  NOR2_X1 U14398 ( .A1(n11196), .A2(n11195), .ZN(n11199) );
  INV_X1 U14399 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15923) );
  AOI21_X1 U14400 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15923), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11197) );
  AOI21_X1 U14401 ( .B1(n10992), .B2(P1_EAX_REG_16__SCAN_IN), .A(n11197), .ZN(
        n11198) );
  OAI21_X1 U14402 ( .B1(n11472), .B2(n11199), .A(n11198), .ZN(n11204) );
  XNOR2_X1 U14403 ( .A(n11205), .B(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15921) );
  NAND2_X1 U14404 ( .A1(n15921), .A2(n11278), .ZN(n11203) );
  NAND2_X1 U14405 ( .A1(n11204), .A2(n11203), .ZN(n15550) );
  INV_X1 U14406 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n22100) );
  OAI21_X1 U14407 ( .B1(n11205), .B2(n15923), .A(n22100), .ZN(n11208) );
  AND2_X1 U14408 ( .A1(n11208), .A2(n11241), .ZN(n15912) );
  AOI22_X1 U14409 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10937), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11212) );
  AOI22_X1 U14410 ( .A1(n11335), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11412), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11211) );
  AOI22_X1 U14411 ( .A1(n10780), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11269), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11210) );
  AOI22_X1 U14412 ( .A1(n10936), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11324), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11209) );
  NAND4_X1 U14413 ( .A1(n11212), .A2(n11211), .A3(n11210), .A4(n11209), .ZN(
        n11218) );
  AOI22_X1 U14414 ( .A1(n10890), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11435), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11216) );
  AOI22_X1 U14415 ( .A1(n11393), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11434), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11215) );
  AOI22_X1 U14416 ( .A1(n10943), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11214) );
  AOI22_X1 U14417 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11213) );
  NAND4_X1 U14418 ( .A1(n11216), .A2(n11215), .A3(n11214), .A4(n11213), .ZN(
        n11217) );
  OR2_X1 U14419 ( .A1(n11218), .A2(n11217), .ZN(n11219) );
  NAND2_X1 U14420 ( .A1(n11494), .A2(n11219), .ZN(n11222) );
  NOR2_X1 U14421 ( .A1(n11682), .A2(n22100), .ZN(n11220) );
  AOI21_X1 U14422 ( .B1(n10992), .B2(P1_EAX_REG_17__SCAN_IN), .A(n11220), .ZN(
        n11221) );
  OAI211_X1 U14423 ( .C1(n15912), .C2(n11455), .A(n11222), .B(n11221), .ZN(
        n15538) );
  INV_X1 U14424 ( .A(n15528), .ZN(n11240) );
  AOI22_X1 U14425 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11412), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11226) );
  AOI22_X1 U14426 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11413), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11225) );
  AOI22_X1 U14427 ( .A1(n10870), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11269), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11224) );
  AOI22_X1 U14428 ( .A1(n11434), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10943), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11223) );
  NAND4_X1 U14429 ( .A1(n11226), .A2(n11225), .A3(n11224), .A4(n11223), .ZN(
        n11234) );
  AOI22_X1 U14430 ( .A1(n10889), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11435), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11232) );
  NAND2_X1 U14431 ( .A1(n10936), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n11228) );
  NAND2_X1 U14432 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n11227) );
  AND3_X1 U14433 ( .A1(n11228), .A2(n11455), .A3(n11227), .ZN(n11231) );
  AOI22_X1 U14434 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10846), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11230) );
  AOI22_X1 U14435 ( .A1(n11335), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11324), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11229) );
  NAND4_X1 U14436 ( .A1(n11232), .A2(n11231), .A3(n11230), .A4(n11229), .ZN(
        n11233) );
  NAND2_X1 U14437 ( .A1(n11472), .A2(n11455), .ZN(n11311) );
  OAI21_X1 U14438 ( .B1(n11234), .B2(n11233), .A(n11311), .ZN(n11236) );
  AOI22_X1 U14439 ( .A1(n10992), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n10952), .ZN(n11235) );
  NAND2_X1 U14440 ( .A1(n11236), .A2(n11235), .ZN(n11238) );
  XNOR2_X1 U14441 ( .A(n11241), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15901) );
  NAND2_X1 U14442 ( .A1(n15901), .A2(n11161), .ZN(n11237) );
  NAND2_X1 U14443 ( .A1(n11238), .A2(n11237), .ZN(n15529) );
  INV_X1 U14444 ( .A(n11243), .ZN(n11245) );
  INV_X1 U14445 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n11244) );
  NAND2_X1 U14446 ( .A1(n11245), .A2(n11244), .ZN(n11246) );
  NAND2_X1 U14447 ( .A1(n11279), .A2(n11246), .ZN(n15892) );
  AOI22_X1 U14448 ( .A1(n10936), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11434), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11250) );
  AOI22_X1 U14449 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11335), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11249) );
  AOI22_X1 U14450 ( .A1(n10890), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11269), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11248) );
  AOI22_X1 U14451 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11247) );
  NAND4_X1 U14452 ( .A1(n11250), .A2(n11249), .A3(n11248), .A4(n11247), .ZN(
        n11256) );
  AOI22_X1 U14453 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11393), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11254) );
  AOI22_X1 U14454 ( .A1(n10870), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11435), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11253) );
  AOI22_X1 U14455 ( .A1(n11324), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11252) );
  AOI22_X1 U14456 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11251) );
  NAND4_X1 U14457 ( .A1(n11254), .A2(n11253), .A3(n11252), .A4(n11251), .ZN(
        n11255) );
  NOR2_X1 U14458 ( .A1(n11256), .A2(n11255), .ZN(n11260) );
  NAND2_X1 U14459 ( .A1(n10952), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11257) );
  NAND2_X1 U14460 ( .A1(n11455), .A2(n11257), .ZN(n11258) );
  AOI21_X1 U14461 ( .B1(n10992), .B2(P1_EAX_REG_19__SCAN_IN), .A(n11258), .ZN(
        n11259) );
  OAI21_X1 U14462 ( .B1(n11472), .B2(n11260), .A(n11259), .ZN(n11261) );
  XNOR2_X1 U14463 ( .A(n11279), .B(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15884) );
  AOI22_X1 U14464 ( .A1(n10992), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n10952), .ZN(n11277) );
  AOI22_X1 U14465 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11435), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11266) );
  AOI22_X1 U14466 ( .A1(n10936), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11413), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11265) );
  AOI22_X1 U14467 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n11335), .B1(
        n11434), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11264) );
  AOI22_X1 U14468 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n11462), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11263) );
  NAND4_X1 U14469 ( .A1(n11266), .A2(n11265), .A3(n11264), .A4(n11263), .ZN(
        n11275) );
  NAND2_X1 U14470 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11268) );
  NAND2_X1 U14471 ( .A1(n10870), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11267) );
  AND3_X1 U14472 ( .A1(n11268), .A2(n11267), .A3(n11455), .ZN(n11273) );
  AOI22_X1 U14473 ( .A1(n11393), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11324), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11272) );
  AOI22_X1 U14474 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n11269), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11271) );
  AOI22_X1 U14475 ( .A1(n10890), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11270) );
  NAND4_X1 U14476 ( .A1(n11273), .A2(n11272), .A3(n11271), .A4(n11270), .ZN(
        n11274) );
  OAI21_X1 U14477 ( .B1(n11275), .B2(n11274), .A(n11311), .ZN(n11276) );
  AOI22_X1 U14478 ( .A1(n15884), .A2(n11278), .B1(n11277), .B2(n11276), .ZN(
        n15493) );
  INV_X1 U14479 ( .A(n11281), .ZN(n11282) );
  INV_X1 U14480 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15483) );
  NAND2_X1 U14481 ( .A1(n11282), .A2(n15483), .ZN(n11283) );
  NAND2_X1 U14482 ( .A1(n11319), .A2(n11283), .ZN(n15874) );
  AOI22_X1 U14483 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11393), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11287) );
  AOI22_X1 U14484 ( .A1(n10936), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10890), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11286) );
  AOI22_X1 U14485 ( .A1(n10780), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11324), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11285) );
  AOI22_X1 U14486 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11284) );
  NAND4_X1 U14487 ( .A1(n11287), .A2(n11286), .A3(n11285), .A4(n11284), .ZN(
        n11293) );
  AOI22_X1 U14488 ( .A1(n10937), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11434), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11291) );
  AOI22_X1 U14489 ( .A1(n11435), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11269), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11290) );
  AOI22_X1 U14490 ( .A1(n11335), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11289) );
  AOI22_X1 U14491 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10943), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11288) );
  NAND4_X1 U14492 ( .A1(n11291), .A2(n11290), .A3(n11289), .A4(n11288), .ZN(
        n11292) );
  NOR2_X1 U14493 ( .A1(n11293), .A2(n11292), .ZN(n11297) );
  NAND2_X1 U14494 ( .A1(n10952), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11294) );
  NAND2_X1 U14495 ( .A1(n11455), .A2(n11294), .ZN(n11295) );
  AOI21_X1 U14496 ( .B1(n10992), .B2(P1_EAX_REG_21__SCAN_IN), .A(n11295), .ZN(
        n11296) );
  OAI21_X1 U14497 ( .B1(n11472), .B2(n11297), .A(n11296), .ZN(n11298) );
  NAND2_X1 U14498 ( .A1(n11299), .A2(n11298), .ZN(n15480) );
  XNOR2_X1 U14499 ( .A(n11319), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15867) );
  NAND2_X1 U14500 ( .A1(n15867), .A2(n11161), .ZN(n11317) );
  AOI22_X1 U14501 ( .A1(n10936), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11462), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11303) );
  AOI22_X1 U14502 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11269), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11302) );
  AOI22_X1 U14503 ( .A1(n11335), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11434), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11301) );
  AOI22_X1 U14504 ( .A1(n10889), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11324), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11300) );
  NAND4_X1 U14505 ( .A1(n11303), .A2(n11302), .A3(n11301), .A4(n11300), .ZN(
        n11313) );
  AOI22_X1 U14506 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11435), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11310) );
  NAND2_X1 U14507 ( .A1(n10937), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11306) );
  NAND2_X1 U14508 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11305) );
  AND3_X1 U14509 ( .A1(n11306), .A2(n11455), .A3(n11305), .ZN(n11309) );
  AOI22_X1 U14510 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11308) );
  AOI22_X1 U14511 ( .A1(n10741), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10846), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11307) );
  NAND4_X1 U14512 ( .A1(n11310), .A2(n11309), .A3(n11308), .A4(n11307), .ZN(
        n11312) );
  OAI21_X1 U14513 ( .B1(n11313), .B2(n11312), .A(n11311), .ZN(n11315) );
  AOI22_X1 U14514 ( .A1(n10992), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n10952), .ZN(n11314) );
  NAND2_X1 U14515 ( .A1(n11315), .A2(n11314), .ZN(n11316) );
  INV_X1 U14516 ( .A(n11321), .ZN(n11322) );
  INV_X1 U14517 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15459) );
  NAND2_X1 U14518 ( .A1(n11322), .A2(n15459), .ZN(n11323) );
  NAND2_X1 U14519 ( .A1(n11370), .A2(n11323), .ZN(n15854) );
  AOI22_X1 U14520 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11393), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11328) );
  AOI22_X1 U14521 ( .A1(n10936), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10870), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11327) );
  AOI22_X1 U14522 ( .A1(n10890), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11434), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11326) );
  AOI22_X1 U14523 ( .A1(n11435), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11324), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11325) );
  NAND4_X1 U14524 ( .A1(n11328), .A2(n11327), .A3(n11326), .A4(n11325), .ZN(
        n11334) );
  AOI22_X1 U14525 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11269), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11332) );
  AOI22_X1 U14526 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11331) );
  AOI22_X1 U14527 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11330) );
  AOI22_X1 U14528 ( .A1(n11335), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11329) );
  NAND4_X1 U14529 ( .A1(n11332), .A2(n11331), .A3(n11330), .A4(n11329), .ZN(
        n11333) );
  NOR2_X1 U14530 ( .A1(n11334), .A2(n11333), .ZN(n11352) );
  AOI22_X1 U14531 ( .A1(n11393), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10870), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11339) );
  AOI22_X1 U14532 ( .A1(n10890), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11435), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11338) );
  AOI22_X1 U14533 ( .A1(n11335), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11269), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11337) );
  AOI22_X1 U14534 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11336) );
  NAND4_X1 U14535 ( .A1(n11339), .A2(n11338), .A3(n11337), .A4(n11336), .ZN(
        n11345) );
  AOI22_X1 U14536 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10936), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11343) );
  AOI22_X1 U14537 ( .A1(n11434), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11324), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11342) );
  AOI22_X1 U14538 ( .A1(n10727), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11341) );
  AOI22_X1 U14539 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11340) );
  NAND4_X1 U14540 ( .A1(n11343), .A2(n11342), .A3(n11341), .A4(n11340), .ZN(
        n11344) );
  NOR2_X1 U14541 ( .A1(n11345), .A2(n11344), .ZN(n11353) );
  XNOR2_X1 U14542 ( .A(n11352), .B(n11353), .ZN(n11349) );
  NAND2_X1 U14543 ( .A1(n10952), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11346) );
  NAND2_X1 U14544 ( .A1(n11455), .A2(n11346), .ZN(n11347) );
  AOI21_X1 U14545 ( .B1(n10992), .B2(P1_EAX_REG_23__SCAN_IN), .A(n11347), .ZN(
        n11348) );
  OAI21_X1 U14546 ( .B1(n11472), .B2(n11349), .A(n11348), .ZN(n11350) );
  XNOR2_X1 U14547 ( .A(n11370), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15852) );
  NOR2_X1 U14548 ( .A1(n11353), .A2(n11352), .ZN(n11383) );
  AOI22_X1 U14549 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11393), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11357) );
  AOI22_X1 U14550 ( .A1(n10936), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10870), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11356) );
  INV_X1 U14551 ( .A(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n21848) );
  AOI22_X1 U14552 ( .A1(n10890), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11434), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11355) );
  AOI22_X1 U14553 ( .A1(n11435), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11324), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11354) );
  NAND4_X1 U14554 ( .A1(n11357), .A2(n11356), .A3(n11355), .A4(n11354), .ZN(
        n11363) );
  AOI22_X1 U14555 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11269), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11361) );
  AOI22_X1 U14556 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11360) );
  AOI22_X1 U14557 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11359) );
  AOI22_X1 U14558 ( .A1(n11335), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11358) );
  NAND4_X1 U14559 ( .A1(n11361), .A2(n11360), .A3(n11359), .A4(n11358), .ZN(
        n11362) );
  OR2_X1 U14560 ( .A1(n11363), .A2(n11362), .ZN(n11382) );
  INV_X1 U14561 ( .A(n11382), .ZN(n11364) );
  XNOR2_X1 U14562 ( .A(n11383), .B(n11364), .ZN(n11367) );
  INV_X1 U14563 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n15734) );
  NAND2_X1 U14564 ( .A1(n10952), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11365) );
  OAI211_X1 U14565 ( .C1(n11492), .C2(n15734), .A(n11455), .B(n11365), .ZN(
        n11366) );
  AOI21_X1 U14566 ( .B1(n11367), .B2(n11494), .A(n11366), .ZN(n11368) );
  INV_X1 U14567 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15848) );
  INV_X1 U14568 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15434) );
  OAI21_X1 U14569 ( .B1(n11370), .B2(n15848), .A(n15434), .ZN(n11371) );
  NAND2_X1 U14570 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11369) );
  NAND2_X1 U14571 ( .A1(n11371), .A2(n11389), .ZN(n15841) );
  AOI22_X1 U14572 ( .A1(n10936), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10890), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11375) );
  AOI22_X1 U14573 ( .A1(n11393), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10870), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11374) );
  AOI22_X1 U14574 ( .A1(n11335), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11373) );
  AOI22_X1 U14575 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11372) );
  NAND4_X1 U14576 ( .A1(n11375), .A2(n11374), .A3(n11373), .A4(n11372), .ZN(
        n11381) );
  AOI22_X1 U14577 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11434), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11379) );
  AOI22_X1 U14578 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11269), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11378) );
  AOI22_X1 U14579 ( .A1(n11435), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11324), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11377) );
  AOI22_X1 U14580 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11376) );
  NAND4_X1 U14581 ( .A1(n11379), .A2(n11378), .A3(n11377), .A4(n11376), .ZN(
        n11380) );
  NOR2_X1 U14582 ( .A1(n11381), .A2(n11380), .ZN(n11392) );
  NAND2_X1 U14583 ( .A1(n11383), .A2(n11382), .ZN(n11391) );
  XNOR2_X1 U14584 ( .A(n11392), .B(n11391), .ZN(n11384) );
  NOR2_X1 U14585 ( .A1(n11384), .A2(n11472), .ZN(n11387) );
  INV_X1 U14586 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n15728) );
  NAND2_X1 U14587 ( .A1(n10952), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11385) );
  OAI211_X1 U14588 ( .C1(n11492), .C2(n15728), .A(n11455), .B(n11385), .ZN(
        n11386) );
  OAI22_X1 U14589 ( .A1(n15841), .A2(n11455), .B1(n11387), .B2(n11386), .ZN(
        n15433) );
  INV_X1 U14590 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n22033) );
  NAND2_X1 U14591 ( .A1(n11389), .A2(n22033), .ZN(n11390) );
  NAND2_X1 U14592 ( .A1(n11410), .A2(n11390), .ZN(n15831) );
  NOR2_X1 U14593 ( .A1(n11392), .A2(n11391), .ZN(n11425) );
  AOI22_X1 U14594 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11393), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11397) );
  AOI22_X1 U14595 ( .A1(n10936), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10870), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11396) );
  AOI22_X1 U14596 ( .A1(n10890), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10871), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11395) );
  AOI22_X1 U14597 ( .A1(n11435), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11324), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11394) );
  NAND4_X1 U14598 ( .A1(n11397), .A2(n11396), .A3(n11395), .A4(n11394), .ZN(
        n11403) );
  AOI22_X1 U14599 ( .A1(n10780), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11269), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11401) );
  AOI22_X1 U14600 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11400) );
  AOI22_X1 U14601 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11399) );
  AOI22_X1 U14602 ( .A1(n11335), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10893), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11398) );
  NAND4_X1 U14603 ( .A1(n11401), .A2(n11400), .A3(n11399), .A4(n11398), .ZN(
        n11402) );
  OR2_X1 U14604 ( .A1(n11403), .A2(n11402), .ZN(n11424) );
  XNOR2_X1 U14605 ( .A(n11425), .B(n11424), .ZN(n11406) );
  AOI21_X1 U14606 ( .B1(n22033), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11404) );
  AOI21_X1 U14607 ( .B1(n10992), .B2(P1_EAX_REG_26__SCAN_IN), .A(n11404), .ZN(
        n11405) );
  OAI21_X1 U14608 ( .B1(n11406), .B2(n11472), .A(n11405), .ZN(n11407) );
  NAND2_X1 U14609 ( .A1(n11408), .A2(n11407), .ZN(n15420) );
  INV_X1 U14610 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15408) );
  NAND2_X1 U14611 ( .A1(n11410), .A2(n15408), .ZN(n11411) );
  NAND2_X1 U14612 ( .A1(n11451), .A2(n11411), .ZN(n15821) );
  AOI22_X1 U14613 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n10889), .B1(
        n10870), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11417) );
  AOI22_X1 U14614 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n11413), .B1(
        n11412), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11416) );
  AOI22_X1 U14615 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n11335), .B1(
        n11269), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11415) );
  AOI22_X1 U14616 ( .A1(n11435), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11324), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11414) );
  NAND4_X1 U14617 ( .A1(n11417), .A2(n11416), .A3(n11415), .A4(n11414), .ZN(
        n11423) );
  AOI22_X1 U14618 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10936), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11421) );
  AOI22_X1 U14619 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n10890), .B1(
        n11434), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11420) );
  AOI22_X1 U14620 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10846), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11419) );
  AOI22_X1 U14621 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n11478), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11418) );
  NAND4_X1 U14622 ( .A1(n11421), .A2(n11420), .A3(n11419), .A4(n11418), .ZN(
        n11422) );
  NOR2_X1 U14623 ( .A1(n11423), .A2(n11422), .ZN(n11433) );
  NAND2_X1 U14624 ( .A1(n11425), .A2(n11424), .ZN(n11432) );
  XNOR2_X1 U14625 ( .A(n11433), .B(n11432), .ZN(n11429) );
  NAND2_X1 U14626 ( .A1(n10952), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11426) );
  NAND2_X1 U14627 ( .A1(n11455), .A2(n11426), .ZN(n11427) );
  AOI21_X1 U14628 ( .B1(n10992), .B2(P1_EAX_REG_27__SCAN_IN), .A(n11427), .ZN(
        n11428) );
  OAI21_X1 U14629 ( .B1(n11429), .B2(n11472), .A(n11428), .ZN(n11430) );
  XNOR2_X1 U14630 ( .A(n11451), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15807) );
  NOR2_X1 U14631 ( .A1(n11433), .A2(n11432), .ZN(n11457) );
  AOI22_X1 U14632 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10889), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11439) );
  AOI22_X1 U14633 ( .A1(n10936), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10937), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11438) );
  AOI22_X1 U14634 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11434), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11437) );
  INV_X1 U14635 ( .A(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n22081) );
  AOI22_X1 U14636 ( .A1(n11435), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11324), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11436) );
  NAND4_X1 U14637 ( .A1(n11439), .A2(n11438), .A3(n11437), .A4(n11436), .ZN(
        n11445) );
  AOI22_X1 U14638 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11269), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11443) );
  AOI22_X1 U14639 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11442) );
  AOI22_X1 U14640 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10943), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11441) );
  AOI22_X1 U14641 ( .A1(n11335), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10846), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11440) );
  NAND4_X1 U14642 ( .A1(n11443), .A2(n11442), .A3(n11441), .A4(n11440), .ZN(
        n11444) );
  OR2_X1 U14643 ( .A1(n11445), .A2(n11444), .ZN(n11456) );
  INV_X1 U14644 ( .A(n11456), .ZN(n11446) );
  XNOR2_X1 U14645 ( .A(n11457), .B(n11446), .ZN(n11449) );
  INV_X1 U14646 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n15715) );
  NAND2_X1 U14647 ( .A1(n10952), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11447) );
  OAI211_X1 U14648 ( .C1(n11492), .C2(n15715), .A(n11455), .B(n11447), .ZN(
        n11448) );
  AOI21_X1 U14649 ( .B1(n11449), .B2(n11494), .A(n11448), .ZN(n11450) );
  INV_X1 U14650 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15805) );
  INV_X1 U14651 ( .A(n11452), .ZN(n11453) );
  INV_X1 U14652 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n11469) );
  NAND2_X1 U14653 ( .A1(n11453), .A2(n11469), .ZN(n11454) );
  NAND2_X1 U14654 ( .A1(n11501), .A2(n11454), .ZN(n15800) );
  NAND2_X1 U14655 ( .A1(n11457), .A2(n11456), .ZN(n11476) );
  AOI22_X1 U14656 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10889), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11461) );
  AOI22_X1 U14657 ( .A1(n10936), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10871), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11460) );
  AOI22_X1 U14658 ( .A1(n10876), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11435), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11459) );
  AOI22_X1 U14659 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11269), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11458) );
  NAND4_X1 U14660 ( .A1(n11461), .A2(n11460), .A3(n11459), .A4(n11458), .ZN(
        n11468) );
  AOI22_X1 U14661 ( .A1(n10870), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11324), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11466) );
  AOI22_X1 U14662 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11465) );
  AOI22_X1 U14663 ( .A1(n11335), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10891), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11464) );
  AOI22_X1 U14664 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10846), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11463) );
  NAND4_X1 U14665 ( .A1(n11466), .A2(n11465), .A3(n11464), .A4(n11463), .ZN(
        n11467) );
  NOR2_X1 U14666 ( .A1(n11468), .A2(n11467), .ZN(n11477) );
  XNOR2_X1 U14667 ( .A(n11476), .B(n11477), .ZN(n11473) );
  AOI21_X1 U14668 ( .B1(n11469), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11470) );
  AOI21_X1 U14669 ( .B1(n10992), .B2(P1_EAX_REG_29__SCAN_IN), .A(n11470), .ZN(
        n11471) );
  OAI21_X1 U14670 ( .B1(n11473), .B2(n11472), .A(n11471), .ZN(n11474) );
  NAND2_X1 U14671 ( .A1(n11475), .A2(n11474), .ZN(n15382) );
  XNOR2_X1 U14672 ( .A(n11501), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15036) );
  NOR2_X1 U14673 ( .A1(n11477), .A2(n11476), .ZN(n11490) );
  AOI22_X1 U14674 ( .A1(n10889), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10871), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11482) );
  AOI22_X1 U14675 ( .A1(n10727), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11481) );
  AOI22_X1 U14676 ( .A1(n11335), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10943), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11480) );
  AOI22_X1 U14677 ( .A1(n10780), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10846), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11479) );
  NAND4_X1 U14678 ( .A1(n11482), .A2(n11481), .A3(n11480), .A4(n11479), .ZN(
        n11488) );
  AOI22_X1 U14679 ( .A1(n11304), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10937), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11486) );
  AOI22_X1 U14680 ( .A1(n10936), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10876), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11485) );
  AOI22_X1 U14681 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11269), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11484) );
  AOI22_X1 U14682 ( .A1(n11435), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11324), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11483) );
  NAND4_X1 U14683 ( .A1(n11486), .A2(n11485), .A3(n11484), .A4(n11483), .ZN(
        n11487) );
  NOR2_X1 U14684 ( .A1(n11488), .A2(n11487), .ZN(n11489) );
  XNOR2_X1 U14685 ( .A(n11490), .B(n11489), .ZN(n11495) );
  INV_X1 U14686 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n15023) );
  OAI21_X1 U14687 ( .B1(n21528), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n10952), .ZN(n11491) );
  OAI21_X1 U14688 ( .B1(n11492), .B2(n15023), .A(n11491), .ZN(n11493) );
  AOI21_X1 U14689 ( .B1(n11495), .B2(n11494), .A(n11493), .ZN(n11496) );
  AOI21_X1 U14690 ( .B1(n15036), .B2(n11161), .A(n11496), .ZN(n11856) );
  NAND2_X1 U14691 ( .A1(n15381), .A2(n11856), .ZN(n11500) );
  AOI22_X1 U14692 ( .A1(n10992), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n11497), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11498) );
  INV_X1 U14693 ( .A(n11498), .ZN(n11499) );
  INV_X1 U14694 ( .A(n11501), .ZN(n11502) );
  NAND2_X1 U14695 ( .A1(n11502), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11503) );
  INV_X1 U14696 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11674) );
  NAND2_X1 U14697 ( .A1(n10816), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11504) );
  INV_X1 U14698 ( .A(n11514), .ZN(n11505) );
  NAND2_X1 U14699 ( .A1(n11505), .A2(n14561), .ZN(n11540) );
  XNOR2_X1 U14700 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11519) );
  NAND2_X1 U14701 ( .A1(n21561), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11507) );
  XNOR2_X1 U14702 ( .A(n11519), .B(n11518), .ZN(n11559) );
  INV_X1 U14703 ( .A(n11559), .ZN(n11517) );
  NAND2_X1 U14704 ( .A1(n10816), .A2(n9724), .ZN(n11506) );
  NAND2_X1 U14705 ( .A1(n11506), .A2(n11661), .ZN(n11525) );
  OAI21_X1 U14706 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21561), .A(
        n11507), .ZN(n11508) );
  INV_X1 U14707 ( .A(n11508), .ZN(n11510) );
  OAI211_X1 U14708 ( .C1(n11557), .C2(n13570), .A(n11525), .B(n11510), .ZN(
        n11513) );
  NAND2_X1 U14709 ( .A1(n11552), .A2(n11510), .ZN(n11511) );
  NAND2_X1 U14710 ( .A1(n11553), .A2(n11511), .ZN(n11512) );
  OAI211_X1 U14711 ( .C1(n11514), .C2(n11517), .A(n11513), .B(n11512), .ZN(
        n11516) );
  NAND2_X1 U14712 ( .A1(n11514), .A2(n11517), .ZN(n11515) );
  OAI211_X1 U14713 ( .C1(n11540), .C2(n11517), .A(n11516), .B(n11515), .ZN(
        n11524) );
  NAND2_X1 U14714 ( .A1(n11519), .A2(n11518), .ZN(n11521) );
  NAND2_X1 U14715 ( .A1(n21665), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11520) );
  NAND2_X1 U14716 ( .A1(n11521), .A2(n11520), .ZN(n11530) );
  XNOR2_X1 U14717 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11529) );
  XNOR2_X1 U14718 ( .A(n11530), .B(n11529), .ZN(n11560) );
  INV_X1 U14719 ( .A(n11560), .ZN(n11526) );
  NAND2_X1 U14720 ( .A1(n11552), .A2(n11526), .ZN(n11522) );
  OAI211_X1 U14721 ( .C1(n11526), .C2(n11541), .A(n11522), .B(n11525), .ZN(
        n11523) );
  INV_X1 U14722 ( .A(n11525), .ZN(n11527) );
  NAND3_X1 U14723 ( .A1(n11527), .A2(n11526), .A3(n11552), .ZN(n11528) );
  NAND2_X1 U14724 ( .A1(n11530), .A2(n11529), .ZN(n11532) );
  NAND2_X1 U14725 ( .A1(n21306), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11531) );
  MUX2_X1 U14726 ( .A(n11533), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n11536) );
  XNOR2_X1 U14727 ( .A(n11537), .B(n11536), .ZN(n11561) );
  INV_X1 U14728 ( .A(n11553), .ZN(n11534) );
  NOR2_X1 U14729 ( .A1(n14352), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11535) );
  NAND2_X1 U14730 ( .A1(n11541), .A2(n11562), .ZN(n11538) );
  INV_X1 U14731 ( .A(n11540), .ZN(n11544) );
  INV_X1 U14732 ( .A(n11562), .ZN(n11542) );
  INV_X1 U14733 ( .A(n11546), .ZN(n11548) );
  NOR2_X1 U14734 ( .A1(n18089), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n11547) );
  INV_X1 U14735 ( .A(n11549), .ZN(n11550) );
  NOR2_X1 U14736 ( .A1(n11557), .A2(n9724), .ZN(n11558) );
  NOR4_X1 U14737 ( .A1(n11562), .A2(n11561), .A3(n11560), .A4(n11559), .ZN(
        n11563) );
  NOR2_X1 U14738 ( .A1(n11564), .A2(n11563), .ZN(n13573) );
  NAND2_X1 U14739 ( .A1(n13563), .A2(n13800), .ZN(n15371) );
  NOR2_X1 U14740 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n21823) );
  NAND2_X1 U14741 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21823), .ZN(n18030) );
  NAND2_X1 U14742 ( .A1(n11161), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n11565) );
  MUX2_X1 U14743 ( .A(n18030), .B(n11565), .S(n21733), .Z(n11566) );
  INV_X1 U14744 ( .A(n11566), .ZN(n11567) );
  OR2_X2 U14745 ( .A1(n11686), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21291) );
  NOR2_X1 U14746 ( .A1(n11567), .A2(n18072), .ZN(n11568) );
  NAND2_X1 U14747 ( .A1(n13425), .A2(n21168), .ZN(n11681) );
  INV_X1 U14748 ( .A(n14008), .ZN(n11811) );
  INV_X1 U14749 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16014) );
  NOR2_X1 U14750 ( .A1(n14238), .A2(n16014), .ZN(n11570) );
  AOI21_X1 U14751 ( .B1(n11811), .B2(P1_EBX_REG_30__SCAN_IN), .A(n11570), .ZN(
        n15030) );
  NAND2_X2 U14752 ( .A1(n9703), .A2(n14238), .ZN(n11576) );
  INV_X1 U14753 ( .A(n11581), .ZN(n11650) );
  NAND2_X1 U14754 ( .A1(n9714), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11571) );
  AND2_X1 U14755 ( .A1(n11607), .A2(n11571), .ZN(n11572) );
  NAND2_X1 U14756 ( .A1(n9734), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n11574) );
  OAI21_X1 U14757 ( .B1(n9703), .B2(P1_EBX_REG_0__SCAN_IN), .A(n11574), .ZN(
        n14009) );
  XNOR2_X1 U14758 ( .A(n11575), .B(n14009), .ZN(n14239) );
  NAND2_X1 U14759 ( .A1(n14239), .A2(n14238), .ZN(n14237) );
  NAND2_X1 U14760 ( .A1(n14237), .A2(n11575), .ZN(n14075) );
  MUX2_X1 U14761 ( .A(n11576), .B(n9734), .S(P1_EBX_REG_2__SCAN_IN), .Z(n11580) );
  NAND2_X1 U14762 ( .A1(n11577), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11578) );
  AND2_X1 U14763 ( .A1(n11607), .A2(n11578), .ZN(n11579) );
  AND2_X1 U14764 ( .A1(n11580), .A2(n11579), .ZN(n14074) );
  INV_X1 U14765 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n21204) );
  NAND2_X1 U14766 ( .A1(n11624), .A2(n21204), .ZN(n11584) );
  INV_X1 U14767 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21300) );
  NAND2_X1 U14768 ( .A1(n14238), .A2(n21204), .ZN(n11582) );
  OAI211_X1 U14769 ( .C1(n9703), .C2(n21300), .A(n11582), .B(n9734), .ZN(
        n11583) );
  INV_X1 U14770 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n14509) );
  NAND2_X1 U14771 ( .A1(n9734), .A2(n14509), .ZN(n11586) );
  INV_X1 U14772 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n21192) );
  NAND2_X1 U14773 ( .A1(n14238), .A2(n21192), .ZN(n11585) );
  NAND3_X1 U14774 ( .A1(n11586), .A2(n11654), .A3(n11585), .ZN(n11587) );
  OAI21_X1 U14775 ( .B1(n11576), .B2(P1_EBX_REG_4__SCAN_IN), .A(n11587), .ZN(
        n14522) );
  INV_X1 U14776 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18080) );
  NAND2_X1 U14777 ( .A1(n18080), .A2(n14008), .ZN(n11589) );
  MUX2_X1 U14778 ( .A(n11649), .B(n11654), .S(P1_EBX_REG_5__SCAN_IN), .Z(
        n11588) );
  NAND2_X1 U14779 ( .A1(n11589), .A2(n11588), .ZN(n15350) );
  INV_X1 U14780 ( .A(n15350), .ZN(n11590) );
  MUX2_X1 U14781 ( .A(n11649), .B(n11654), .S(P1_EBX_REG_7__SCAN_IN), .Z(
        n11592) );
  INV_X1 U14782 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18069) );
  NAND2_X1 U14783 ( .A1(n14008), .A2(n18069), .ZN(n11591) );
  MUX2_X1 U14784 ( .A(n11576), .B(n9734), .S(P1_EBX_REG_6__SCAN_IN), .Z(n11595) );
  NAND2_X1 U14785 ( .A1(n11577), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11593) );
  AND2_X1 U14786 ( .A1(n11607), .A2(n11593), .ZN(n11594) );
  NAND2_X1 U14787 ( .A1(n11595), .A2(n11594), .ZN(n14840) );
  MUX2_X1 U14788 ( .A(n11576), .B(n9734), .S(P1_EBX_REG_8__SCAN_IN), .Z(n11598) );
  NAND2_X1 U14789 ( .A1(n11577), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11596) );
  AND2_X1 U14790 ( .A1(n11607), .A2(n11596), .ZN(n11597) );
  NAND2_X1 U14791 ( .A1(n11598), .A2(n11597), .ZN(n15705) );
  INV_X1 U14792 ( .A(n14876), .ZN(n11602) );
  MUX2_X1 U14793 ( .A(n11649), .B(n11654), .S(P1_EBX_REG_9__SCAN_IN), .Z(
        n11600) );
  INV_X1 U14794 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15992) );
  NAND2_X1 U14795 ( .A1(n14008), .A2(n15992), .ZN(n11599) );
  NAND2_X1 U14796 ( .A1(n11600), .A2(n11599), .ZN(n14877) );
  INV_X1 U14797 ( .A(n14877), .ZN(n11601) );
  INV_X1 U14798 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15703) );
  NAND2_X1 U14799 ( .A1(n11624), .A2(n15703), .ZN(n11605) );
  INV_X1 U14800 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16206) );
  NAND2_X1 U14801 ( .A1(n14238), .A2(n15703), .ZN(n11603) );
  OAI211_X1 U14802 ( .C1(n9703), .C2(n16206), .A(n11603), .B(n9734), .ZN(
        n11604) );
  MUX2_X1 U14803 ( .A(n11576), .B(n9734), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n11609) );
  NAND2_X1 U14804 ( .A1(n11577), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11606) );
  AND2_X1 U14805 ( .A1(n11607), .A2(n11606), .ZN(n11608) );
  NAND2_X1 U14806 ( .A1(n11609), .A2(n11608), .ZN(n15629) );
  MUX2_X1 U14807 ( .A(n11576), .B(n9734), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n11611) );
  NAND2_X1 U14808 ( .A1(n11577), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11610) );
  INV_X1 U14809 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n15699) );
  NAND2_X1 U14810 ( .A1(n11624), .A2(n15699), .ZN(n11614) );
  INV_X1 U14811 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11840) );
  NAND2_X1 U14812 ( .A1(n14238), .A2(n15699), .ZN(n11612) );
  OAI211_X1 U14813 ( .C1(n9703), .C2(n11840), .A(n11612), .B(n9734), .ZN(
        n11613) );
  MUX2_X1 U14814 ( .A(n11576), .B(n9734), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n11616) );
  NAND2_X1 U14815 ( .A1(n11577), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11615) );
  NAND2_X1 U14816 ( .A1(n11616), .A2(n11615), .ZN(n15581) );
  NAND2_X1 U14817 ( .A1(n15601), .A2(n15581), .ZN(n15570) );
  MUX2_X1 U14818 ( .A(n11649), .B(n11654), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n11618) );
  INV_X1 U14819 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n22124) );
  NAND2_X1 U14820 ( .A1(n14008), .A2(n22124), .ZN(n11617) );
  NAND2_X1 U14821 ( .A1(n11618), .A2(n11617), .ZN(n15573) );
  OR2_X2 U14822 ( .A1(n15570), .A2(n15573), .ZN(n15571) );
  INV_X1 U14823 ( .A(n11576), .ZN(n11651) );
  INV_X1 U14824 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n11619) );
  NAND2_X1 U14825 ( .A1(n11651), .A2(n11619), .ZN(n11623) );
  INV_X1 U14826 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16162) );
  NAND2_X1 U14827 ( .A1(n9734), .A2(n16162), .ZN(n11621) );
  NAND2_X1 U14828 ( .A1(n14238), .A2(n11619), .ZN(n11620) );
  NAND3_X1 U14829 ( .A1(n11621), .A2(n11654), .A3(n11620), .ZN(n11622) );
  INV_X1 U14830 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n15694) );
  NAND2_X1 U14831 ( .A1(n11624), .A2(n15694), .ZN(n11627) );
  INV_X1 U14832 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16147) );
  NAND2_X1 U14833 ( .A1(n14238), .A2(n15694), .ZN(n11625) );
  OAI211_X1 U14834 ( .C1(n9703), .C2(n16147), .A(n11625), .B(n9734), .ZN(
        n11626) );
  AND2_X2 U14835 ( .A1(n15553), .A2(n15539), .ZN(n15526) );
  MUX2_X1 U14836 ( .A(n11576), .B(n9734), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n11629) );
  NAND2_X1 U14837 ( .A1(n11577), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11628) );
  NAND2_X1 U14838 ( .A1(n11629), .A2(n11628), .ZN(n15527) );
  INV_X1 U14839 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11771) );
  INV_X1 U14840 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n22099) );
  NAND2_X1 U14841 ( .A1(n14238), .A2(n22099), .ZN(n11630) );
  OAI211_X1 U14842 ( .C1(n9703), .C2(n11771), .A(n11630), .B(n9734), .ZN(
        n11631) );
  OAI21_X1 U14843 ( .B1(n11649), .B2(P1_EBX_REG_19__SCAN_IN), .A(n11631), .ZN(
        n15507) );
  INV_X1 U14844 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n15691) );
  NAND2_X1 U14845 ( .A1(n11651), .A2(n15691), .ZN(n11635) );
  INV_X1 U14846 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11772) );
  NAND2_X1 U14847 ( .A1(n9734), .A2(n11772), .ZN(n11633) );
  NAND2_X1 U14848 ( .A1(n14238), .A2(n15691), .ZN(n11632) );
  NAND3_X1 U14849 ( .A1(n11633), .A2(n11654), .A3(n11632), .ZN(n11634) );
  MUX2_X1 U14850 ( .A(n11649), .B(n11654), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n11637) );
  INV_X1 U14851 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16107) );
  NAND2_X1 U14852 ( .A1(n14008), .A2(n16107), .ZN(n11636) );
  NAND2_X1 U14853 ( .A1(n11637), .A2(n11636), .ZN(n15482) );
  MUX2_X1 U14854 ( .A(n11576), .B(n9734), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n11639) );
  NAND2_X1 U14855 ( .A1(n11577), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11638) );
  NAND2_X1 U14856 ( .A1(n11639), .A2(n11638), .ZN(n15467) );
  NAND2_X1 U14857 ( .A1(n15481), .A2(n15467), .ZN(n15453) );
  MUX2_X1 U14858 ( .A(n11649), .B(n11654), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n11640) );
  OAI21_X1 U14859 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n11811), .A(
        n11640), .ZN(n15454) );
  MUX2_X1 U14860 ( .A(n11576), .B(n9734), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n11642) );
  NAND2_X1 U14861 ( .A1(n11577), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11641) );
  MUX2_X1 U14862 ( .A(n11649), .B(n11654), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n11644) );
  INV_X1 U14863 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16060) );
  NAND2_X1 U14864 ( .A1(n14008), .A2(n16060), .ZN(n11643) );
  AND2_X1 U14865 ( .A1(n11644), .A2(n11643), .ZN(n15430) );
  MUX2_X1 U14866 ( .A(n11576), .B(n9734), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n11646) );
  NAND2_X1 U14867 ( .A1(n11577), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11645) );
  NAND2_X1 U14868 ( .A1(n11646), .A2(n11645), .ZN(n15417) );
  INV_X1 U14869 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16041) );
  INV_X1 U14870 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n15684) );
  NAND2_X1 U14871 ( .A1(n14238), .A2(n15684), .ZN(n11647) );
  OAI211_X1 U14872 ( .C1(n9703), .C2(n16041), .A(n11647), .B(n9734), .ZN(
        n11648) );
  OAI21_X1 U14873 ( .B1(n11649), .B2(P1_EBX_REG_27__SCAN_IN), .A(n11648), .ZN(
        n15403) );
  MUX2_X1 U14874 ( .A(n11651), .B(n11650), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n11652) );
  AOI21_X1 U14875 ( .B1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n11577), .A(
        n11652), .ZN(n15399) );
  INV_X1 U14876 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11838) );
  NOR2_X1 U14877 ( .A1(n11577), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n11653) );
  AOI21_X1 U14878 ( .B1(n14008), .B2(n11838), .A(n11653), .ZN(n15027) );
  MUX2_X1 U14879 ( .A(n15027), .B(n11653), .S(n9703), .Z(n15379) );
  AOI22_X1 U14881 ( .A1(n11811), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n11577), .ZN(n11655) );
  NOR2_X1 U14882 ( .A1(n21820), .A2(n13570), .ZN(n11672) );
  NAND2_X1 U14883 ( .A1(n14561), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n11668) );
  NAND2_X1 U14884 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n18092) );
  AND2_X1 U14885 ( .A1(n18092), .A2(n21528), .ZN(n18022) );
  NOR2_X1 U14886 ( .A1(n11668), .A2(n18022), .ZN(n11657) );
  AND2_X1 U14887 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(P1_REIP_REG_29__SCAN_IN), 
        .ZN(n11666) );
  INV_X1 U14888 ( .A(n11658), .ZN(n11660) );
  INV_X1 U14889 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n11659) );
  NAND2_X1 U14890 ( .A1(n11660), .A2(n11659), .ZN(n18039) );
  NAND2_X1 U14891 ( .A1(n11661), .A2(n18039), .ZN(n11777) );
  AND2_X1 U14892 ( .A1(n11777), .A2(n18022), .ZN(n11670) );
  OR2_X1 U14893 ( .A1(n21210), .A2(n21200), .ZN(n15628) );
  INV_X1 U14894 ( .A(n15628), .ZN(n15675) );
  AOI21_X1 U14895 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(P1_REIP_REG_28__SCAN_IN), 
        .A(n15675), .ZN(n11665) );
  INV_X1 U14896 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n15829) );
  INV_X1 U14897 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n21775) );
  INV_X1 U14898 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n21138) );
  NAND4_X1 U14899 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n21125)
         );
  NAND4_X1 U14900 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(P1_REIP_REG_7__SCAN_IN), 
        .A3(P1_REIP_REG_6__SCAN_IN), .A4(P1_REIP_REG_5__SCAN_IN), .ZN(n21124)
         );
  NOR3_X1 U14901 ( .A1(n21138), .A2(n21125), .A3(n21124), .ZN(n15644) );
  NAND2_X1 U14902 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n15644), .ZN(n15645) );
  INV_X1 U14903 ( .A(n15645), .ZN(n11662) );
  AND2_X1 U14904 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n11662), .ZN(n15613) );
  AND2_X1 U14905 ( .A1(n15613), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n15515) );
  INV_X1 U14906 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n21770) );
  NAND2_X1 U14907 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(P1_REIP_REG_14__SCAN_IN), 
        .ZN(n15555) );
  NAND2_X1 U14908 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n15558) );
  NOR3_X1 U14909 ( .A1(n21770), .A2(n15555), .A3(n15558), .ZN(n15520) );
  NAND2_X1 U14910 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n15520), .ZN(n15512) );
  INV_X1 U14911 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n15890) );
  NOR2_X1 U14912 ( .A1(n15512), .A2(n15890), .ZN(n11663) );
  NAND2_X1 U14913 ( .A1(n15515), .A2(n11663), .ZN(n15497) );
  NOR2_X1 U14914 ( .A1(n21775), .A2(n15497), .ZN(n15472) );
  AND3_X1 U14915 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .A3(n15472), .ZN(n15460) );
  AND2_X1 U14916 ( .A1(n15460), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n15435) );
  AND2_X1 U14917 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n11664) );
  NAND2_X1 U14918 ( .A1(n15435), .A2(n11664), .ZN(n15421) );
  NOR2_X1 U14919 ( .A1(n15829), .A2(n15421), .ZN(n15410) );
  INV_X1 U14920 ( .A(n21200), .ZN(n21123) );
  OAI21_X1 U14921 ( .B1(n21126), .B2(n15410), .A(n21123), .ZN(n15425) );
  NOR2_X1 U14922 ( .A1(n11665), .A2(n15425), .ZN(n15395) );
  OAI21_X1 U14923 ( .B1(n11666), .B2(n15675), .A(n15395), .ZN(n15031) );
  AND3_X1 U14924 ( .A1(n21210), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n15410), 
        .ZN(n15394) );
  NAND2_X1 U14925 ( .A1(n15394), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n15383) );
  INV_X1 U14926 ( .A(n11666), .ZN(n11667) );
  NOR3_X1 U14927 ( .A1(n15383), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n11667), 
        .ZN(n11677) );
  INV_X1 U14928 ( .A(n11668), .ZN(n11669) );
  NOR2_X1 U14929 ( .A1(n11670), .A2(n11669), .ZN(n11671) );
  INV_X1 U14930 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n11675) );
  INV_X1 U14931 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n11673) );
  OAI22_X1 U14932 ( .A1(n21205), .A2(n11675), .B1(n11674), .B2(n21203), .ZN(
        n11676) );
  AOI211_X1 U14933 ( .C1(n15031), .C2(P1_REIP_REG_31__SCAN_IN), .A(n11677), 
        .B(n11676), .ZN(n11678) );
  NAND2_X1 U14934 ( .A1(n11681), .A2(n11680), .ZN(P1_U2809) );
  NOR2_X1 U14935 ( .A1(n11682), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n14395) );
  AND2_X1 U14936 ( .A1(n21733), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n11683) );
  NAND2_X1 U14937 ( .A1(n16270), .A2(n13570), .ZN(n11685) );
  NAND2_X1 U14938 ( .A1(n13414), .A2(n11808), .ZN(n18011) );
  NOR2_X2 U14939 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21679) );
  NAND2_X1 U14940 ( .A1(n11686), .A2(n21667), .ZN(n21818) );
  NAND2_X1 U14941 ( .A1(n21818), .A2(n21733), .ZN(n11687) );
  NAND2_X1 U14942 ( .A1(n21733), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n18021) );
  NAND2_X1 U14943 ( .A1(n21528), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n11688) );
  NAND2_X1 U14944 ( .A1(n18021), .A2(n11688), .ZN(n13746) );
  NAND2_X1 U14945 ( .A1(n18072), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n11849) );
  NAND2_X1 U14946 ( .A1(n18048), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11689) );
  OAI211_X1 U14947 ( .C1(n15035), .C2(n18056), .A(n11849), .B(n11689), .ZN(
        n11690) );
  INV_X1 U14948 ( .A(n11784), .ZN(n11820) );
  NAND2_X1 U14949 ( .A1(n11717), .A2(n11724), .ZN(n11710) );
  NAND2_X1 U14950 ( .A1(n11710), .A2(n11711), .ZN(n11709) );
  NAND2_X1 U14951 ( .A1(n11709), .A2(n11700), .ZN(n11695) );
  INV_X1 U14952 ( .A(n11696), .ZN(n11691) );
  OR2_X1 U14953 ( .A1(n11695), .A2(n11691), .ZN(n11739) );
  XNOR2_X1 U14954 ( .A(n11739), .B(n11740), .ZN(n11692) );
  NAND2_X1 U14955 ( .A1(n11692), .A2(n11798), .ZN(n11693) );
  INV_X1 U14956 ( .A(n11695), .ZN(n11697) );
  OAI211_X1 U14957 ( .C1(n11697), .C2(n11696), .A(n11798), .B(n11739), .ZN(
        n11698) );
  INV_X1 U14958 ( .A(n11700), .ZN(n11701) );
  XNOR2_X1 U14959 ( .A(n11709), .B(n11701), .ZN(n11702) );
  NAND2_X1 U14960 ( .A1(n11702), .A2(n11798), .ZN(n11703) );
  AND2_X2 U14961 ( .A1(n11704), .A2(n11703), .ZN(n11705) );
  INV_X2 U14962 ( .A(n11705), .ZN(n14507) );
  NAND2_X1 U14963 ( .A1(n11705), .A2(n21300), .ZN(n11706) );
  OAI21_X1 U14964 ( .B1(n11707), .B2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n11706), .ZN(n11708) );
  INV_X1 U14965 ( .A(n11708), .ZN(n11734) );
  OAI21_X1 U14966 ( .B1(n11711), .B2(n11710), .A(n11709), .ZN(n11713) );
  NAND2_X1 U14967 ( .A1(n13570), .A2(n14553), .ZN(n11723) );
  INV_X1 U14968 ( .A(n11723), .ZN(n11712) );
  AOI21_X1 U14969 ( .B1(n11713), .B2(n11798), .A(n11712), .ZN(n11714) );
  NAND2_X1 U14970 ( .A1(n11715), .A2(n11714), .ZN(n14071) );
  NAND2_X1 U14971 ( .A1(n14561), .A2(n11716), .ZN(n11722) );
  INV_X1 U14972 ( .A(n11724), .ZN(n11718) );
  XNOR2_X1 U14973 ( .A(n11718), .B(n11717), .ZN(n11720) );
  AOI21_X1 U14974 ( .B1(n11720), .B2(n11798), .A(n11719), .ZN(n11721) );
  NAND2_X1 U14975 ( .A1(n16317), .A2(n11784), .ZN(n11727) );
  OAI21_X1 U14976 ( .B1(n21825), .B2(n11724), .A(n11723), .ZN(n11725) );
  INV_X1 U14977 ( .A(n11725), .ZN(n11726) );
  NAND2_X1 U14978 ( .A1(n11727), .A2(n11726), .ZN(n13743) );
  NAND2_X1 U14979 ( .A1(n13743), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11728) );
  XNOR2_X1 U14980 ( .A(n11729), .B(n11728), .ZN(n14059) );
  NAND2_X1 U14981 ( .A1(n14059), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11731) );
  INV_X1 U14982 ( .A(n11728), .ZN(n13744) );
  NAND2_X1 U14983 ( .A1(n11729), .A2(n13744), .ZN(n11730) );
  INV_X1 U14984 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11827) );
  NAND2_X1 U14985 ( .A1(n11732), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11733) );
  NAND2_X1 U14986 ( .A1(n11734), .A2(n14503), .ZN(n11735) );
  NAND2_X1 U14987 ( .A1(n11736), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11737) );
  INV_X1 U14988 ( .A(n11739), .ZN(n11741) );
  NAND2_X1 U14989 ( .A1(n11741), .A2(n11740), .ZN(n11749) );
  XNOR2_X1 U14990 ( .A(n11749), .B(n11750), .ZN(n11742) );
  NAND2_X1 U14991 ( .A1(n11742), .A2(n11798), .ZN(n11743) );
  NAND2_X1 U14992 ( .A1(n11744), .A2(n11743), .ZN(n11745) );
  NOR2_X1 U14993 ( .A1(n11820), .A2(n11746), .ZN(n11747) );
  INV_X1 U14994 ( .A(n11749), .ZN(n11751) );
  NAND2_X1 U14995 ( .A1(n11751), .A2(n11750), .ZN(n11756) );
  NAND2_X1 U14996 ( .A1(n11798), .A2(n11755), .ZN(n11752) );
  OR2_X1 U14997 ( .A1(n11756), .A2(n11752), .ZN(n11753) );
  XNOR2_X1 U14998 ( .A(n11756), .B(n11755), .ZN(n11757) );
  NAND2_X1 U14999 ( .A1(n11757), .A2(n11798), .ZN(n11758) );
  NOR2_X1 U15000 ( .A1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11761) );
  OR2_X1 U15001 ( .A1(n15979), .A2(n15992), .ZN(n11762) );
  NAND2_X1 U15002 ( .A1(n15979), .A2(n15992), .ZN(n11763) );
  NAND2_X1 U15003 ( .A1(n15979), .A2(n11840), .ZN(n11764) );
  NAND2_X1 U15004 ( .A1(n15939), .A2(n11764), .ZN(n15959) );
  INV_X1 U15005 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16214) );
  NAND2_X1 U15006 ( .A1(n15979), .A2(n16214), .ZN(n15957) );
  NAND2_X1 U15007 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11765) );
  NAND2_X1 U15008 ( .A1(n15979), .A2(n11765), .ZN(n15955) );
  NAND2_X1 U15009 ( .A1(n15957), .A2(n15955), .ZN(n11766) );
  INV_X1 U15010 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16176) );
  OR2_X1 U15011 ( .A1(n15979), .A2(n16176), .ZN(n11767) );
  NAND2_X1 U15012 ( .A1(n15979), .A2(n22124), .ZN(n15930) );
  NOR2_X1 U15013 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15953) );
  NAND2_X1 U15014 ( .A1(n15953), .A2(n16214), .ZN(n15904) );
  NAND2_X1 U15015 ( .A1(n16162), .A2(n16147), .ZN(n11768) );
  NOR2_X1 U15016 ( .A1(n15904), .A2(n11768), .ZN(n11769) );
  NOR2_X1 U15017 ( .A1(n15993), .A2(n11769), .ZN(n11770) );
  XNOR2_X1 U15018 ( .A(n15993), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15897) );
  AND2_X1 U15019 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16096) );
  NAND2_X1 U15020 ( .A1(n16096), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16093) );
  INV_X1 U15021 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16141) );
  INV_X1 U15022 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16069) );
  NAND2_X1 U15023 ( .A1(n16060), .A2(n16069), .ZN(n15808) );
  AND2_X1 U15024 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16048) );
  NAND2_X1 U15025 ( .A1(n16048), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16050) );
  AND2_X1 U15026 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16029) );
  INV_X1 U15027 ( .A(n11773), .ZN(n11774) );
  NOR2_X1 U15028 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16028) );
  INV_X1 U15029 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16049) );
  NAND3_X1 U15030 ( .A1(n11774), .A2(n16028), .A3(n16049), .ZN(n11775) );
  NOR2_X1 U15031 ( .A1(n15993), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15796) );
  AND2_X1 U15032 ( .A1(n13573), .A2(n18092), .ZN(n13417) );
  NAND2_X1 U15033 ( .A1(n14561), .A2(n18039), .ZN(n11776) );
  NAND2_X1 U15034 ( .A1(n13417), .A2(n11776), .ZN(n11783) );
  AND2_X1 U15035 ( .A1(n11777), .A2(n18092), .ZN(n11779) );
  INV_X1 U15036 ( .A(n10792), .ZN(n14593) );
  NAND2_X1 U15037 ( .A1(n14593), .A2(n9724), .ZN(n11778) );
  AOI21_X1 U15038 ( .B1(n11555), .B2(n11779), .A(n11778), .ZN(n11780) );
  MUX2_X1 U15039 ( .A(n11783), .B(n11782), .S(n11781), .Z(n11790) );
  INV_X1 U15040 ( .A(n13575), .ZN(n11788) );
  INV_X1 U15041 ( .A(n13414), .ZN(n11787) );
  AND2_X1 U15042 ( .A1(n11784), .A2(n10821), .ZN(n11789) );
  NOR2_X1 U15043 ( .A1(n11789), .A2(n13570), .ZN(n11785) );
  AND2_X1 U15044 ( .A1(n11786), .A2(n11785), .ZN(n11804) );
  AOI21_X1 U15045 ( .B1(n11788), .B2(n11787), .A(n11804), .ZN(n13796) );
  NAND2_X1 U15046 ( .A1(n17992), .A2(n11789), .ZN(n13794) );
  NAND3_X1 U15047 ( .A1(n11790), .A2(n13796), .A3(n13794), .ZN(n11791) );
  INV_X1 U15048 ( .A(n11792), .ZN(n18086) );
  OR2_X1 U15049 ( .A1(n11808), .A2(n15651), .ZN(n11793) );
  NAND2_X1 U15050 ( .A1(n13414), .A2(n11793), .ZN(n13569) );
  OAI211_X1 U15051 ( .C1(n10795), .C2(n11800), .A(n13569), .B(n11794), .ZN(
        n11795) );
  NOR2_X1 U15052 ( .A1(n18086), .A2(n11795), .ZN(n11796) );
  INV_X1 U15053 ( .A(n11797), .ZN(n11803) );
  NAND2_X1 U15054 ( .A1(n11555), .A2(n11798), .ZN(n18024) );
  OAI21_X1 U15055 ( .B1(n11800), .B2(n11799), .A(n18024), .ZN(n11801) );
  INV_X1 U15056 ( .A(n11801), .ZN(n11802) );
  NAND2_X1 U15057 ( .A1(n11803), .A2(n21282), .ZN(n11853) );
  INV_X1 U15058 ( .A(n11804), .ZN(n11815) );
  INV_X1 U15059 ( .A(n11805), .ZN(n11810) );
  OAI21_X1 U15060 ( .B1(n11808), .B2(n11806), .A(n11807), .ZN(n11809) );
  AOI21_X1 U15061 ( .B1(n11811), .B2(n11810), .A(n11809), .ZN(n11814) );
  INV_X1 U15062 ( .A(n11684), .ZN(n11812) );
  NAND2_X1 U15063 ( .A1(n11812), .A2(n9703), .ZN(n11813) );
  NAND4_X1 U15064 ( .A1(n11815), .A2(n11814), .A3(n10825), .A4(n11813), .ZN(
        n13802) );
  INV_X1 U15065 ( .A(n11816), .ZN(n11817) );
  NOR2_X1 U15066 ( .A1(n13802), .A2(n11817), .ZN(n11818) );
  NAND2_X1 U15067 ( .A1(n13575), .A2(n14561), .ZN(n17995) );
  OR2_X1 U15068 ( .A1(n11819), .A2(n11820), .ZN(n13807) );
  NAND2_X1 U15069 ( .A1(n16252), .A2(n16203), .ZN(n16257) );
  NAND2_X1 U15070 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16259) );
  INV_X1 U15071 ( .A(n16259), .ZN(n16237) );
  AND2_X1 U15072 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16237), .ZN(
        n16229) );
  NAND2_X1 U15073 ( .A1(n16229), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16222) );
  NAND2_X1 U15074 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11821) );
  NOR2_X1 U15075 ( .A1(n16222), .A2(n11821), .ZN(n16215) );
  NAND2_X1 U15076 ( .A1(n16215), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11828) );
  NAND2_X1 U15077 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21278) );
  INV_X1 U15078 ( .A(n21278), .ZN(n16251) );
  NAND3_X1 U15079 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n16251), .ZN(n16255) );
  OR2_X1 U15080 ( .A1(n18080), .A2(n16255), .ZN(n16200) );
  OR2_X1 U15081 ( .A1(n11828), .A2(n16200), .ZN(n16185) );
  NAND3_X1 U15082 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16148) );
  INV_X1 U15083 ( .A(n16148), .ZN(n11822) );
  AND2_X1 U15084 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n11822), .ZN(
        n16138) );
  NAND2_X1 U15085 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16138), .ZN(
        n11844) );
  NOR2_X1 U15086 ( .A1(n11840), .A2(n11844), .ZN(n16091) );
  INV_X1 U15087 ( .A(n16091), .ZN(n11823) );
  NOR2_X1 U15088 ( .A1(n16185), .A2(n11823), .ZN(n11830) );
  INV_X1 U15089 ( .A(n14013), .ZN(n16086) );
  INV_X1 U15090 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21912) );
  NAND2_X1 U15091 ( .A1(n16086), .A2(n21912), .ZN(n11826) );
  NAND2_X1 U15092 ( .A1(n11824), .A2(n21291), .ZN(n11825) );
  INV_X1 U15093 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14243) );
  OAI21_X1 U15094 ( .B1(n21912), .B2(n14243), .A(n11827), .ZN(n16212) );
  NAND3_X1 U15095 ( .A1(n16251), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        n16212), .ZN(n16236) );
  NOR2_X1 U15096 ( .A1(n11828), .A2(n16236), .ZN(n16134) );
  NAND2_X1 U15097 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n16134), .ZN(
        n11842) );
  OAI21_X1 U15098 ( .B1(n11844), .B2(n11842), .A(n16198), .ZN(n11829) );
  INV_X1 U15099 ( .A(n16096), .ZN(n16114) );
  INV_X1 U15100 ( .A(n16257), .ZN(n16137) );
  NAND2_X1 U15101 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11831) );
  NAND2_X1 U15102 ( .A1(n16257), .A2(n11831), .ZN(n11832) );
  INV_X1 U15103 ( .A(n16186), .ZN(n16089) );
  NAND2_X1 U15104 ( .A1(n16089), .A2(n16050), .ZN(n11835) );
  INV_X1 U15105 ( .A(n16048), .ZN(n11833) );
  NAND2_X1 U15106 ( .A1(n16086), .A2(n11833), .ZN(n11834) );
  OAI211_X1 U15107 ( .C1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n16203), .A(
        n11835), .B(n11834), .ZN(n11836) );
  NOR2_X1 U15108 ( .A1(n16068), .A2(n11836), .ZN(n16061) );
  INV_X1 U15109 ( .A(n11837), .ZN(n11839) );
  INV_X1 U15110 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13815) );
  NOR2_X1 U15111 ( .A1(n16185), .A2(n11840), .ZN(n11841) );
  NAND2_X1 U15112 ( .A1(n16207), .A2(n11841), .ZN(n16066) );
  INV_X1 U15113 ( .A(n11842), .ZN(n16177) );
  NAND2_X1 U15114 ( .A1(n16198), .A2(n16177), .ZN(n11843) );
  NAND2_X1 U15115 ( .A1(n16066), .A2(n11843), .ZN(n16161) );
  INV_X1 U15116 ( .A(n11844), .ZN(n11845) );
  NAND2_X1 U15117 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n11845), .ZN(
        n11846) );
  NOR2_X1 U15118 ( .A1(n16093), .A2(n11846), .ZN(n11847) );
  NAND2_X1 U15119 ( .A1(n16161), .A2(n11847), .ZN(n16079) );
  INV_X1 U15120 ( .A(n16030), .ZN(n16038) );
  NAND3_X1 U15121 ( .A1(n16038), .A2(n16029), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16013) );
  NOR3_X1 U15122 ( .A1(n16013), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n16014), .ZN(n11848) );
  INV_X1 U15123 ( .A(n11849), .ZN(n11850) );
  NOR2_X1 U15124 ( .A1(n11848), .A2(n11850), .ZN(n11851) );
  OAI21_X1 U15125 ( .B1(n11855), .B2(n21294), .A(n11854), .ZN(P1_U3000) );
  INV_X1 U15126 ( .A(n15043), .ZN(n15019) );
  NAND2_X1 U15127 ( .A1(n15019), .A2(n18052), .ZN(n11866) );
  INV_X1 U15128 ( .A(n15036), .ZN(n11858) );
  NAND2_X1 U15129 ( .A1(n18072), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n16011) );
  NAND2_X1 U15130 ( .A1(n18048), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11857) );
  OAI211_X1 U15131 ( .C1(n11858), .C2(n18056), .A(n16011), .B(n11857), .ZN(
        n11859) );
  INV_X1 U15132 ( .A(n11859), .ZN(n11865) );
  INV_X1 U15133 ( .A(n11860), .ZN(n11861) );
  NAND2_X1 U15134 ( .A1(n11862), .A2(n11861), .ZN(n11863) );
  NAND2_X1 U15135 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17880) );
  INV_X1 U15136 ( .A(n17880), .ZN(n11867) );
  AND2_X2 U15137 ( .A1(n17879), .A2(n18426), .ZN(n17854) );
  NAND2_X1 U15138 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18427) );
  INV_X1 U15140 ( .A(n19178), .ZN(n11868) );
  NOR2_X2 U15141 ( .A1(n11882), .A2(n19122), .ZN(n11877) );
  NAND2_X1 U15142 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n19054) );
  CLKBUF_X1 U15143 ( .A(n11869), .Z(n11872) );
  NAND2_X1 U15144 ( .A1(n11869), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11886) );
  CLKBUF_X1 U15145 ( .A(n11886), .Z(n17785) );
  OAI21_X1 U15146 ( .B1(n11872), .B2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n17785), .ZN(n17829) );
  INV_X1 U15147 ( .A(n17829), .ZN(n18273) );
  AOI21_X1 U15148 ( .B1(n11871), .B2(n19031), .A(n11872), .ZN(n19028) );
  OAI21_X1 U15149 ( .B1(n11873), .B2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n11871), .ZN(n19040) );
  INV_X1 U15150 ( .A(n19040), .ZN(n18293) );
  INV_X1 U15151 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n19056) );
  INV_X1 U15152 ( .A(n9887), .ZN(n11876) );
  NAND2_X1 U15153 ( .A1(n11876), .A2(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11874) );
  AOI21_X1 U15154 ( .B1(n19056), .B2(n11874), .A(n11873), .ZN(n19058) );
  INV_X1 U15155 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n19068) );
  AOI22_X1 U15156 ( .A1(n11876), .A2(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        n19068), .B2(n9887), .ZN(n19076) );
  INV_X1 U15157 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n19347) );
  NOR2_X1 U15158 ( .A1(n19347), .A2(n11875), .ZN(n11879) );
  INV_X1 U15159 ( .A(n11879), .ZN(n19051) );
  AOI21_X1 U15160 ( .B1(n19053), .B2(n19051), .A(n11876), .ZN(n19083) );
  INV_X1 U15161 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n19096) );
  NAND3_X1 U15162 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n11878), .A3(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11880) );
  AOI21_X1 U15163 ( .B1(n19096), .B2(n11880), .A(n11879), .ZN(n19099) );
  INV_X1 U15164 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n21843) );
  NAND2_X1 U15165 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n11878), .ZN(
        n11881) );
  XOR2_X1 U15166 ( .A(n21843), .B(n11881), .Z(n19115) );
  NOR2_X1 U15167 ( .A1(n19347), .A2(n11882), .ZN(n11884) );
  INV_X1 U15168 ( .A(n11884), .ZN(n19094) );
  AOI22_X1 U15169 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n11878), .B1(
        n19122), .B2(n19094), .ZN(n19124) );
  INV_X1 U15170 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n19143) );
  INV_X1 U15171 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n19154) );
  NAND2_X1 U15172 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n11883), .ZN(
        n18428) );
  INV_X1 U15173 ( .A(n18428), .ZN(n17840) );
  NAND3_X1 U15174 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A3(n17840), .ZN(n18396) );
  INV_X1 U15175 ( .A(n18396), .ZN(n11888) );
  NAND2_X1 U15176 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n11888), .ZN(
        n19141) );
  OR2_X1 U15177 ( .A1(n19154), .A2(n19141), .ZN(n11885) );
  AOI21_X1 U15178 ( .B1(n19143), .B2(n11885), .A(n11884), .ZN(n19146) );
  XOR2_X1 U15179 ( .A(n19154), .B(n19141), .Z(n19157) );
  OAI21_X1 U15180 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n11888), .A(
        n19141), .ZN(n19173) );
  INV_X1 U15181 ( .A(n19173), .ZN(n18380) );
  INV_X1 U15182 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n18263) );
  NOR2_X2 U15183 ( .A1(n11886), .A2(n18263), .ZN(n11892) );
  NAND2_X1 U15184 ( .A1(n11892), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11887) );
  NOR2_X1 U15185 ( .A1(n19347), .A2(n11890), .ZN(n18535) );
  NAND2_X1 U15186 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18535), .ZN(
        n18519) );
  NOR2_X1 U15187 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18519), .ZN(
        n18527) );
  NAND3_X1 U15188 ( .A1(n18426), .A2(n11891), .A3(n18527), .ZN(n18398) );
  NOR2_X1 U15190 ( .A1(n18320), .A2(n10450), .ZN(n18314) );
  AOI21_X1 U15193 ( .B1(n18263), .B2(n17785), .A(n11893), .ZN(n18261) );
  NOR2_X1 U15194 ( .A1(n18260), .A2(n10450), .ZN(n13378) );
  INV_X1 U15195 ( .A(n13378), .ZN(n11895) );
  INV_X1 U15196 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n17800) );
  XNOR2_X1 U15197 ( .A(n11893), .B(n17800), .ZN(n17802) );
  INV_X1 U15198 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n13932) );
  INV_X1 U15199 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n20216) );
  NAND3_X1 U15200 ( .A1(n13932), .A2(n20107), .A3(n20216), .ZN(n20115) );
  NOR2_X1 U15201 ( .A1(n18914), .A2(n20115), .ZN(n18598) );
  NAND2_X1 U15202 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n20218) );
  NAND2_X1 U15203 ( .A1(n9712), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11902) );
  AND2_X4 U15204 ( .A1(n11898), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14457) );
  NAND2_X1 U15205 ( .A1(n14457), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11901) );
  NAND2_X1 U15206 ( .A1(n9705), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11900) );
  NAND2_X1 U15207 ( .A1(n18652), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11899) );
  INV_X2 U15208 ( .A(n13862), .ZN(n14951) );
  NAND2_X1 U15209 ( .A1(n14951), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11906) );
  INV_X2 U15210 ( .A(n13784), .ZN(n18777) );
  NAND2_X1 U15211 ( .A1(n14968), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11905) );
  INV_X1 U15212 ( .A(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n18693) );
  OR2_X1 U15213 ( .A1(n18775), .A2(n18693), .ZN(n11904) );
  INV_X1 U15214 ( .A(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n18696) );
  OR2_X1 U15215 ( .A1(n18773), .A2(n18696), .ZN(n11903) );
  NAND2_X1 U15216 ( .A1(n18760), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11912) );
  NAND2_X1 U15217 ( .A1(n17630), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11911) );
  INV_X2 U15218 ( .A(n9781), .ZN(n18616) );
  NAND2_X1 U15219 ( .A1(n18616), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11910) );
  AND2_X2 U15220 ( .A1(n14028), .A2(n11908), .ZN(n12013) );
  NAND2_X1 U15221 ( .A1(n12013), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11909) );
  INV_X1 U15222 ( .A(n14031), .ZN(n11913) );
  INV_X2 U15223 ( .A(n11955), .ZN(n13659) );
  INV_X1 U15224 ( .A(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14906) );
  OAI22_X1 U15225 ( .A1(n11955), .A2(n14906), .B1(n11972), .B2(n18688), .ZN(
        n11920) );
  NOR2_X1 U15226 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11916) );
  INV_X1 U15227 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18794) );
  INV_X2 U15228 ( .A(n18717), .ZN(n18764) );
  INV_X1 U15229 ( .A(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11918) );
  OAI22_X1 U15230 ( .A1(n18715), .A2(n18794), .B1(n18764), .B2(n11918), .ZN(
        n11919) );
  NOR2_X1 U15231 ( .A1(n11920), .A2(n11919), .ZN(n11921) );
  NAND2_X1 U15232 ( .A1(n9712), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11928) );
  NAND2_X1 U15233 ( .A1(n14457), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n11927) );
  NAND2_X1 U15234 ( .A1(n9706), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11926) );
  NAND2_X1 U15235 ( .A1(n18652), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n11925) );
  NAND2_X1 U15236 ( .A1(n14951), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n11932) );
  NAND2_X1 U15237 ( .A1(n18646), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n11931) );
  INV_X1 U15238 ( .A(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17670) );
  OR2_X1 U15239 ( .A1(n18775), .A2(n17670), .ZN(n11930) );
  INV_X1 U15240 ( .A(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17671) );
  OR2_X1 U15241 ( .A1(n18773), .A2(n17671), .ZN(n11929) );
  INV_X1 U15242 ( .A(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n18729) );
  INV_X1 U15243 ( .A(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n18735) );
  OAI22_X1 U15244 ( .A1(n11955), .A2(n18729), .B1(n17695), .B2(n18735), .ZN(
        n11934) );
  OAI22_X1 U15245 ( .A1(n18715), .A2(n18807), .B1(n18764), .B2(n17678), .ZN(
        n11933) );
  NOR2_X1 U15246 ( .A1(n11934), .A2(n11933), .ZN(n11940) );
  NAND2_X1 U15247 ( .A1(n18760), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n11938) );
  NAND2_X1 U15248 ( .A1(n17630), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n11937) );
  NAND2_X1 U15249 ( .A1(n18616), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n11936) );
  NAND2_X1 U15250 ( .A1(n12013), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n11935) );
  NAND2_X1 U15251 ( .A1(n9712), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11946) );
  INV_X1 U15252 ( .A(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14799) );
  NAND2_X1 U15253 ( .A1(n9706), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11944) );
  NAND2_X1 U15254 ( .A1(n18652), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11943) );
  NAND2_X1 U15255 ( .A1(n14951), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11950) );
  NAND2_X1 U15256 ( .A1(n14968), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11949) );
  INV_X1 U15257 ( .A(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n18614) );
  OR2_X1 U15258 ( .A1(n18775), .A2(n18614), .ZN(n11948) );
  INV_X1 U15259 ( .A(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14930) );
  OR2_X1 U15260 ( .A1(n18773), .A2(n14930), .ZN(n11947) );
  NAND2_X1 U15261 ( .A1(n14896), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11954) );
  NAND2_X1 U15262 ( .A1(n17630), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11953) );
  NAND2_X1 U15263 ( .A1(n18616), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11952) );
  NAND2_X1 U15264 ( .A1(n12013), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11951) );
  NAND2_X1 U15265 ( .A1(n13659), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11959) );
  NAND2_X1 U15266 ( .A1(n10682), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11958) );
  NAND2_X1 U15267 ( .A1(n14112), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11957) );
  NAND2_X1 U15268 ( .A1(n18717), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11956) );
  NAND3_X1 U15269 ( .A1(n19646), .A2(n19634), .A3(n19654), .ZN(n12071) );
  INV_X1 U15270 ( .A(n12071), .ZN(n12049) );
  NAND2_X1 U15271 ( .A1(n9712), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11967) );
  NAND2_X1 U15272 ( .A1(n14457), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11966) );
  NAND2_X1 U15273 ( .A1(n9705), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11965) );
  NAND2_X1 U15274 ( .A1(n18652), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11964) );
  NAND2_X1 U15275 ( .A1(n14951), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11971) );
  NAND2_X1 U15276 ( .A1(n14968), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11970) );
  INV_X1 U15277 ( .A(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17624) );
  OR2_X1 U15278 ( .A1(n18775), .A2(n17624), .ZN(n11969) );
  INV_X1 U15279 ( .A(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17627) );
  OR2_X1 U15280 ( .A1(n18773), .A2(n17627), .ZN(n11968) );
  INV_X1 U15281 ( .A(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11973) );
  INV_X1 U15282 ( .A(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14291) );
  OAI22_X1 U15283 ( .A1(n18763), .A2(n11973), .B1(n17695), .B2(n14291), .ZN(
        n11977) );
  INV_X1 U15284 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11975) );
  OAI22_X1 U15285 ( .A1(n18715), .A2(n11975), .B1(n11974), .B2(n17641), .ZN(
        n11976) );
  NOR2_X1 U15286 ( .A1(n11977), .A2(n11976), .ZN(n11983) );
  NAND2_X1 U15287 ( .A1(n14896), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11981) );
  NAND2_X1 U15288 ( .A1(n17630), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11980) );
  NAND2_X1 U15290 ( .A1(n17631), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11979) );
  NAND2_X1 U15291 ( .A1(n12013), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11978) );
  NAND2_X1 U15292 ( .A1(n9712), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11989) );
  NAND2_X1 U15293 ( .A1(n14457), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n11988) );
  NAND2_X1 U15294 ( .A1(n9705), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11987) );
  NAND2_X1 U15295 ( .A1(n18652), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n11986) );
  NAND2_X1 U15296 ( .A1(n14951), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n11993) );
  NAND2_X1 U15297 ( .A1(n14968), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11992) );
  INV_X1 U15298 ( .A(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17653) );
  OR2_X1 U15299 ( .A1(n18775), .A2(n17653), .ZN(n11991) );
  INV_X1 U15300 ( .A(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17655) );
  OR2_X1 U15301 ( .A1(n18773), .A2(n17655), .ZN(n11990) );
  INV_X1 U15302 ( .A(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14991) );
  INV_X1 U15303 ( .A(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13897) );
  OAI22_X1 U15304 ( .A1(n11955), .A2(n14991), .B1(n14983), .B2(n13897), .ZN(
        n11996) );
  INV_X1 U15305 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11994) );
  INV_X2 U15306 ( .A(n18717), .ZN(n17698) );
  INV_X1 U15307 ( .A(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14979) );
  OAI22_X1 U15308 ( .A1(n18715), .A2(n11994), .B1(n17698), .B2(n14979), .ZN(
        n11995) );
  NOR2_X1 U15309 ( .A1(n11996), .A2(n11995), .ZN(n12002) );
  NAND2_X1 U15310 ( .A1(n14896), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n12000) );
  NAND2_X1 U15311 ( .A1(n17630), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n11999) );
  NAND2_X1 U15312 ( .A1(n17631), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n11998) );
  INV_X2 U15313 ( .A(n17608), .ZN(n18692) );
  NAND2_X1 U15314 ( .A1(n18692), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11997) );
  NAND2_X1 U15315 ( .A1(n19642), .A2(n13674), .ZN(n12047) );
  NAND2_X1 U15316 ( .A1(n18624), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n12008) );
  NAND2_X1 U15317 ( .A1(n13784), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n12007) );
  NAND2_X1 U15318 ( .A1(n18742), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n12006) );
  INV_X1 U15319 ( .A(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n18637) );
  OR2_X1 U15320 ( .A1(n18775), .A2(n18637), .ZN(n12005) );
  NAND2_X1 U15321 ( .A1(n9712), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n12012) );
  NAND2_X1 U15322 ( .A1(n14457), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n12011) );
  NAND2_X1 U15323 ( .A1(n9706), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n12010) );
  NAND2_X1 U15324 ( .A1(n18652), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n12009) );
  NAND2_X1 U15325 ( .A1(n18760), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n12017) );
  NAND2_X1 U15326 ( .A1(n17630), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n12016) );
  NAND2_X1 U15327 ( .A1(n17631), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n12015) );
  NAND2_X1 U15328 ( .A1(n12013), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n12014) );
  NAND2_X1 U15329 ( .A1(n13659), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n12021) );
  NAND2_X1 U15330 ( .A1(n10682), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12020) );
  NAND2_X1 U15331 ( .A1(n14112), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n12019) );
  NAND2_X1 U15332 ( .A1(n18717), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n12018) );
  NAND2_X1 U15333 ( .A1(n14457), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12029) );
  NAND2_X1 U15334 ( .A1(n9712), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12028) );
  NAND2_X1 U15335 ( .A1(n9705), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12027) );
  NAND2_X1 U15336 ( .A1(n18652), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12026) );
  NAND2_X1 U15337 ( .A1(n14968), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12033) );
  NAND2_X1 U15338 ( .A1(n14951), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12032) );
  INV_X1 U15339 ( .A(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14916) );
  OR2_X1 U15340 ( .A1(n18775), .A2(n14916), .ZN(n12031) );
  INV_X1 U15341 ( .A(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n18714) );
  OR2_X1 U15342 ( .A1(n18773), .A2(n18714), .ZN(n12030) );
  OAI22_X1 U15343 ( .A1(n18613), .A2(n18753), .B1(n17695), .B2(n19819), .ZN(
        n12037) );
  INV_X1 U15344 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12035) );
  INV_X1 U15345 ( .A(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n18756) );
  NAND2_X1 U15346 ( .A1(n18616), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12034) );
  OAI21_X1 U15347 ( .B1(n12035), .B2(n18715), .A(n12034), .ZN(n12036) );
  NOR2_X1 U15348 ( .A1(n12037), .A2(n12036), .ZN(n12043) );
  NAND2_X1 U15349 ( .A1(n14896), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12041) );
  NAND2_X1 U15350 ( .A1(n18692), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12040) );
  NAND2_X1 U15351 ( .A1(n18717), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12039) );
  NAND2_X1 U15352 ( .A1(n17630), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12038) );
  NAND2_X1 U15353 ( .A1(n19650), .A2(n18917), .ZN(n12046) );
  NOR2_X1 U15354 ( .A1(n12047), .A2(n12046), .ZN(n12048) );
  INV_X1 U15355 ( .A(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17690) );
  NAND2_X1 U15356 ( .A1(n9705), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12052) );
  NAND2_X1 U15357 ( .A1(n9712), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n12051) );
  NAND2_X1 U15358 ( .A1(n18652), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12050) );
  NAND2_X1 U15359 ( .A1(n14968), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12057) );
  NAND2_X1 U15360 ( .A1(n14951), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12056) );
  INV_X1 U15361 ( .A(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17694) );
  OR2_X1 U15362 ( .A1(n18775), .A2(n17694), .ZN(n12055) );
  INV_X1 U15363 ( .A(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17699) );
  OR2_X1 U15364 ( .A1(n18773), .A2(n17699), .ZN(n12054) );
  INV_X1 U15365 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18809) );
  OAI22_X1 U15366 ( .A1(n9781), .A2(n14943), .B1(n18715), .B2(n18809), .ZN(
        n12060) );
  INV_X1 U15367 ( .A(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12058) );
  OAI22_X1 U15368 ( .A1(n17695), .A2(n17689), .B1(n17698), .B2(n12058), .ZN(
        n12059) );
  NAND2_X1 U15369 ( .A1(n13659), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12064) );
  NAND2_X1 U15370 ( .A1(n14896), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12063) );
  INV_X2 U15371 ( .A(n17608), .ZN(n17693) );
  NAND2_X1 U15372 ( .A1(n17693), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12062) );
  NAND2_X1 U15373 ( .A1(n17630), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12061) );
  NAND4_X1 U15374 ( .A1(n19638), .A2(n19628), .A3(n19642), .A4(n19654), .ZN(
        n12069) );
  AND2_X2 U15375 ( .A1(n12086), .A2(n13690), .ZN(n18235) );
  NAND2_X1 U15376 ( .A1(n19628), .A2(n20217), .ZN(n13876) );
  NAND2_X1 U15377 ( .A1(n19638), .A2(n13685), .ZN(n12070) );
  NOR2_X1 U15378 ( .A1(n19646), .A2(n13685), .ZN(n13964) );
  INV_X1 U15379 ( .A(n13964), .ZN(n12075) );
  NOR2_X1 U15380 ( .A1(n19628), .A2(n18973), .ZN(n13672) );
  INV_X1 U15381 ( .A(n13672), .ZN(n12074) );
  NOR2_X1 U15382 ( .A1(n12075), .A2(n12074), .ZN(n13688) );
  INV_X1 U15383 ( .A(n13688), .ZN(n12077) );
  AOI21_X1 U15384 ( .B1(n12077), .B2(n13676), .A(n19638), .ZN(n12085) );
  OAI211_X1 U15385 ( .C1(n13680), .C2(n19650), .A(n19628), .B(n13771), .ZN(
        n12084) );
  AOI21_X1 U15386 ( .B1(n18917), .B2(n19638), .A(n18606), .ZN(n12083) );
  INV_X1 U15387 ( .A(n13691), .ZN(n12078) );
  NAND2_X1 U15388 ( .A1(n12078), .A2(n12079), .ZN(n12082) );
  OAI21_X1 U15389 ( .B1(n19646), .B2(n12079), .A(n19634), .ZN(n12080) );
  OAI21_X1 U15390 ( .B1(n12080), .B2(n13673), .A(n13691), .ZN(n12081) );
  NAND4_X1 U15391 ( .A1(n12084), .A2(n12083), .A3(n12082), .A4(n12081), .ZN(
        n13689) );
  MUX2_X1 U15392 ( .A(n12088), .B(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n13692) );
  NAND2_X1 U15393 ( .A1(n13692), .A2(n13681), .ZN(n12103) );
  NAND2_X1 U15394 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n12088), .ZN(
        n12090) );
  NAND2_X1 U15395 ( .A1(n12103), .A2(n12090), .ZN(n12101) );
  MUX2_X1 U15396 ( .A(n20085), .B(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n12100) );
  NAND2_X1 U15397 ( .A1(n12101), .A2(n12100), .ZN(n12092) );
  NAND2_X1 U15398 ( .A1(n20085), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12091) );
  NAND2_X1 U15399 ( .A1(n12092), .A2(n12091), .ZN(n12093) );
  NAND2_X1 U15400 ( .A1(n12093), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12097) );
  OAI22_X1 U15401 ( .A1(n12093), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n20088), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n12095) );
  AOI21_X1 U15402 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n12097), .A(
        n12095), .ZN(n12094) );
  AOI21_X1 U15403 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20088), .A(
        n12094), .ZN(n13698) );
  NAND2_X1 U15404 ( .A1(n12095), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12099) );
  NOR2_X1 U15405 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20088), .ZN(
        n12096) );
  NAND2_X1 U15406 ( .A1(n12097), .A2(n12096), .ZN(n12098) );
  NAND2_X1 U15407 ( .A1(n12099), .A2(n12098), .ZN(n13694) );
  XNOR2_X1 U15408 ( .A(n12101), .B(n12100), .ZN(n12102) );
  OAI21_X1 U15409 ( .B1(n13681), .B2(n13692), .A(n12103), .ZN(n12104) );
  NAND2_X1 U15410 ( .A1(n18973), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n12111) );
  AOI211_X4 U15411 ( .C1(n20216), .C2(n20218), .A(n20231), .B(n12111), .ZN(
        n18575) );
  NAND2_X1 U15412 ( .A1(n18580), .A2(n18802), .ZN(n18574) );
  INV_X1 U15413 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n18541) );
  INV_X1 U15414 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n18513) );
  INV_X1 U15415 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n18480) );
  NAND2_X1 U15416 ( .A1(n18491), .A2(n18480), .ZN(n18472) );
  INV_X1 U15417 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n18461) );
  INV_X1 U15418 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n18438) );
  NAND2_X1 U15419 ( .A1(n18445), .A2(n18438), .ZN(n18437) );
  INV_X1 U15420 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n18415) );
  NAND2_X1 U15421 ( .A1(n18419), .A2(n18415), .ZN(n18414) );
  INV_X1 U15422 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n18386) );
  INV_X1 U15423 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n18368) );
  INV_X1 U15424 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n21897) );
  INV_X1 U15425 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n21874) );
  INV_X1 U15426 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n18306) );
  NAND2_X1 U15427 ( .A1(n18312), .A2(n18306), .ZN(n18305) );
  INV_X1 U15428 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n18669) );
  NAND2_X1 U15429 ( .A1(n18290), .A2(n18669), .ZN(n18284) );
  INV_X1 U15430 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n18661) );
  NAND2_X1 U15431 ( .A1(n18270), .A2(n18661), .ZN(n12113) );
  NAND2_X1 U15432 ( .A1(n18575), .A2(n12113), .ZN(n18266) );
  INV_X1 U15433 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n20131) );
  NOR2_X2 U15434 ( .A1(n22024), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n20187) );
  INV_X1 U15435 ( .A(n20225), .ZN(n20208) );
  NAND2_X2 U15436 ( .A1(n20208), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n20189) );
  NOR2_X1 U15437 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n20118) );
  INV_X1 U15438 ( .A(n20118), .ZN(n12106) );
  NAND3_X1 U15439 ( .A1(n20131), .A2(n20189), .A3(n12106), .ZN(n20215) );
  NAND2_X1 U15440 ( .A1(n20215), .A2(n20217), .ZN(n12108) );
  INV_X1 U15441 ( .A(n20218), .ZN(n20121) );
  NOR2_X1 U15442 ( .A1(P3_STATEBS16_REG_SCAN_IN), .A2(n20121), .ZN(n12107) );
  NAND2_X1 U15443 ( .A1(n12108), .A2(n12107), .ZN(n20097) );
  INV_X1 U15444 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n20176) );
  INV_X1 U15445 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n20173) );
  INV_X1 U15446 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n20162) );
  INV_X1 U15447 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n20159) );
  INV_X1 U15448 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n20155) );
  INV_X1 U15449 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n20151) );
  NAND2_X1 U15450 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n18567) );
  NOR2_X1 U15451 ( .A1(n20137), .A2(n18567), .ZN(n18553) );
  NAND3_X1 U15452 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(P3_REIP_REG_4__SCAN_IN), 
        .A3(n18553), .ZN(n18514) );
  NAND3_X1 U15453 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(P3_REIP_REG_7__SCAN_IN), 
        .A3(P3_REIP_REG_6__SCAN_IN), .ZN(n18465) );
  NAND2_X1 U15454 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_9__SCAN_IN), 
        .ZN(n18477) );
  NOR4_X1 U15455 ( .A1(n20151), .A2(n18514), .A3(n18465), .A4(n18477), .ZN(
        n18448) );
  NAND2_X1 U15456 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n18448), .ZN(n18435) );
  NOR2_X1 U15457 ( .A1(n20155), .A2(n18435), .ZN(n18420) );
  NAND2_X1 U15458 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n18420), .ZN(n18421) );
  NOR2_X1 U15459 ( .A1(n20159), .A2(n18421), .ZN(n18395) );
  NAND2_X1 U15460 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n18395), .ZN(n18385) );
  NAND4_X1 U15461 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n18358), .A3(
        P3_REIP_REG_19__SCAN_IN), .A4(P3_REIP_REG_18__SCAN_IN), .ZN(n18329) );
  NAND2_X1 U15462 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .ZN(n18337) );
  NOR3_X1 U15463 ( .A1(n20173), .A2(n18329), .A3(n18337), .ZN(n18311) );
  NAND2_X1 U15464 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n18311), .ZN(n18301) );
  NOR2_X1 U15465 ( .A1(n20176), .A2(n18301), .ZN(n18289) );
  NAND2_X1 U15466 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n18289), .ZN(n12109) );
  NAND4_X1 U15467 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n18283), .ZN(n13383) );
  NOR2_X1 U15468 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n13383), .ZN(n13380) );
  NAND3_X1 U15469 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n12110) );
  NOR2_X1 U15470 ( .A1(n21986), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n20110) );
  INV_X1 U15471 ( .A(n20110), .ZN(n20102) );
  NOR2_X1 U15472 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n14052) );
  AND2_X2 U15473 ( .A1(n20230), .A2(n13932), .ZN(n19556) );
  NOR2_X1 U15474 ( .A1(n19556), .A2(n18598), .ZN(n18561) );
  INV_X1 U15475 ( .A(n20233), .ZN(n20229) );
  AND2_X1 U15476 ( .A1(n18578), .A2(n12109), .ZN(n18288) );
  NOR2_X1 U15477 ( .A1(n18589), .A2(n18288), .ZN(n18287) );
  INV_X1 U15478 ( .A(n18287), .ZN(n18296) );
  AOI21_X1 U15479 ( .B1(n18578), .B2(n12110), .A(n18296), .ZN(n18269) );
  INV_X1 U15480 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n22051) );
  OAI22_X1 U15481 ( .A1(n18269), .A2(n22051), .B1(n17800), .B2(n18593), .ZN(
        n12116) );
  NAND2_X1 U15482 ( .A1(n20097), .A2(n12111), .ZN(n12112) );
  NOR2_X1 U15483 ( .A1(n18579), .A2(n12113), .ZN(n13379) );
  OAI21_X1 U15484 ( .B1(n18596), .B2(n13379), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n12114) );
  INV_X1 U15485 ( .A(n12114), .ZN(n12115) );
  NAND2_X1 U15486 ( .A1(n12119), .A2(n12118), .ZN(P3_U2641) );
  INV_X1 U15487 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12273) );
  AOI22_X1 U15488 ( .A1(n9719), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9721), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12123) );
  AND2_X4 U15489 ( .A1(n12313), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12311) );
  INV_X2 U15490 ( .A(n15259), .ZN(n12190) );
  AOI22_X1 U15491 ( .A1(n12311), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n15323), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12122) );
  AOI22_X1 U15492 ( .A1(n15157), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9730), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12121) );
  AOI22_X1 U15493 ( .A1(n9732), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(n9729), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12127) );
  AOI22_X1 U15494 ( .A1(n9720), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(n9721), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12126) );
  AOI22_X1 U15495 ( .A1(n12311), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9723), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12125) );
  AOI22_X1 U15496 ( .A1(n12311), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n15323), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12133) );
  AOI22_X1 U15497 ( .A1(n9720), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(n9721), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12132) );
  AOI22_X1 U15498 ( .A1(n9728), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(n9727), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12131) );
  NAND4_X1 U15499 ( .A1(n12132), .A2(n12133), .A3(n10671), .A4(n12131), .ZN(
        n12140) );
  AOI22_X1 U15500 ( .A1(n9732), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(n9729), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12136) );
  AOI22_X1 U15501 ( .A1(n12311), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9723), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12134) );
  AOI22_X1 U15502 ( .A1(n9728), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9727), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12137) );
  NAND2_X1 U15503 ( .A1(n12138), .A2(n12137), .ZN(n12139) );
  AOI22_X1 U15504 ( .A1(n9728), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(n9727), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12143) );
  AOI22_X1 U15505 ( .A1(n15157), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9730), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12142) );
  AOI22_X1 U15506 ( .A1(n12311), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12190), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12141) );
  AOI22_X1 U15507 ( .A1(n9727), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_10__3__SCAN_IN), .B2(n9728), .ZN(n12146) );
  AOI22_X1 U15508 ( .A1(n9732), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(n9730), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12145) );
  AOI22_X1 U15509 ( .A1(n12311), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12190), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12144) );
  NAND2_X1 U15510 ( .A1(n12900), .A2(n13148), .ZN(n12217) );
  AOI22_X1 U15511 ( .A1(n9719), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(n9721), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12149) );
  AOI22_X1 U15512 ( .A1(n9732), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(n9730), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12148) );
  AOI22_X1 U15513 ( .A1(n9728), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9727), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12156) );
  AOI22_X1 U15514 ( .A1(n9731), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(n9730), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12155) );
  AOI22_X1 U15515 ( .A1(n12311), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9723), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12153) );
  NAND4_X1 U15516 ( .A1(n12156), .A2(n12155), .A3(n12154), .A4(n12153), .ZN(
        n12157) );
  NAND2_X1 U15517 ( .A1(n12157), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12158) );
  AOI22_X1 U15518 ( .A1(n9732), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(n9720), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12163) );
  AOI22_X1 U15519 ( .A1(n12311), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9723), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12162) );
  AOI22_X1 U15520 ( .A1(n9736), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9726), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12161) );
  AOI22_X1 U15521 ( .A1(n9730), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9721), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12160) );
  AOI22_X1 U15522 ( .A1(n9731), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(n9730), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12166) );
  AOI22_X1 U15523 ( .A1(n12311), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9723), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12164) );
  INV_X1 U15524 ( .A(n12210), .ZN(n12168) );
  NAND2_X1 U15525 ( .A1(n12168), .A2(n12202), .ZN(n12173) );
  AOI22_X1 U15526 ( .A1(n12311), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n15323), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12170) );
  AOI22_X1 U15527 ( .A1(n9736), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(n9727), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12172) );
  AOI22_X1 U15528 ( .A1(n12311), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12190), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12171) );
  NAND2_X1 U15529 ( .A1(n12173), .A2(n20433), .ZN(n12176) );
  AOI22_X1 U15530 ( .A1(n9728), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(n9727), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12181) );
  AOI22_X1 U15531 ( .A1(n9732), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(n9729), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12180) );
  AOI22_X1 U15532 ( .A1(n9719), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(n9721), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12179) );
  AOI22_X1 U15533 ( .A1(n12311), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12190), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12178) );
  AND4_X1 U15534 ( .A1(n12181), .A2(n12180), .A3(n12179), .A4(n12178), .ZN(
        n12182) );
  NAND2_X1 U15535 ( .A1(n12182), .A2(n12129), .ZN(n12189) );
  AOI22_X1 U15536 ( .A1(n15157), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9721), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12183) );
  AOI22_X1 U15537 ( .A1(n9736), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9727), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12186) );
  AOI22_X1 U15538 ( .A1(n12311), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12190), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12185) );
  NAND4_X1 U15539 ( .A1(n12187), .A2(n12186), .A3(n12185), .A4(n12184), .ZN(
        n12188) );
  AOI22_X1 U15540 ( .A1(n9728), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(n9727), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12194) );
  AOI22_X1 U15541 ( .A1(n9732), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(n9730), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12193) );
  AOI22_X1 U15542 ( .A1(n9720), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(n9721), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12192) );
  AOI22_X1 U15543 ( .A1(n12311), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12190), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12191) );
  NAND4_X1 U15544 ( .A1(n12194), .A2(n12193), .A3(n12192), .A4(n12191), .ZN(
        n12200) );
  AOI22_X1 U15545 ( .A1(n12311), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n15323), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12197) );
  AOI22_X1 U15546 ( .A1(n9728), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9727), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12196) );
  AOI22_X1 U15547 ( .A1(n9729), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9721), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12195) );
  NAND4_X1 U15548 ( .A1(n12198), .A2(n12197), .A3(n12196), .A4(n12195), .ZN(
        n12199) );
  NOR2_X2 U15549 ( .A1(n12898), .A2(n9715), .ZN(n12203) );
  INV_X1 U15550 ( .A(n12208), .ZN(n12209) );
  NAND2_X1 U15551 ( .A1(n12245), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12214) );
  NOR2_X1 U15552 ( .A1(n12213), .A2(n12600), .ZN(n12212) );
  AND2_X1 U15553 ( .A1(n12905), .A2(n14331), .ZN(n14428) );
  AND2_X1 U15554 ( .A1(n12600), .A2(n12905), .ZN(n12216) );
  INV_X1 U15555 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n20979) );
  NAND2_X1 U15556 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12221) );
  AND3_X1 U15557 ( .A1(n14420), .A2(n12207), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n12222) );
  OAI22_X1 U15558 ( .A1(n12245), .A2(n12222), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n12809), .ZN(n12226) );
  INV_X1 U15559 ( .A(n12223), .ZN(n12224) );
  AOI22_X1 U15560 ( .A1(n12224), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n16421), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n12225) );
  NAND2_X1 U15561 ( .A1(n12226), .A2(n12225), .ZN(n12268) );
  BUF_X4 U15562 ( .A(n12227), .Z(n12890) );
  INV_X1 U15563 ( .A(n12228), .ZN(n12229) );
  NAND2_X1 U15564 ( .A1(n12230), .A2(n12229), .ZN(n13143) );
  NAND2_X1 U15565 ( .A1(n13143), .A2(n12231), .ZN(n12232) );
  NAND2_X1 U15566 ( .A1(n12232), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12241) );
  NAND2_X1 U15567 ( .A1(n12809), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n12239) );
  INV_X1 U15568 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n12235) );
  INV_X1 U15569 ( .A(n16421), .ZN(n14746) );
  NAND2_X1 U15570 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12233) );
  AND2_X1 U15571 ( .A1(n14746), .A2(n12233), .ZN(n12234) );
  INV_X1 U15572 ( .A(n12236), .ZN(n12237) );
  OAI211_X2 U15573 ( .C1(n12890), .C2(n13584), .A(n12241), .B(n12240), .ZN(
        n12267) );
  NAND2_X1 U15574 ( .A1(n12268), .A2(n12267), .ZN(n12264) );
  NAND2_X1 U15575 ( .A1(n12265), .A2(n12264), .ZN(n12244) );
  NAND2_X1 U15576 ( .A1(n12254), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12247) );
  AOI21_X1 U15577 ( .B1(n17596), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n12246) );
  INV_X1 U15578 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n16707) );
  INV_X1 U15579 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n20981) );
  NAND2_X1 U15580 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12249) );
  AOI21_X2 U15581 ( .B1(n13223), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n12251), .ZN(n12252) );
  NAND2_X1 U15582 ( .A1(n12254), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12256) );
  NAND2_X1 U15583 ( .A1(n16421), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12255) );
  NAND2_X1 U15584 ( .A1(n12256), .A2(n12255), .ZN(n12261) );
  INV_X1 U15585 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n12259) );
  NAND2_X1 U15586 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12257) );
  OAI211_X1 U15587 ( .C1(n12248), .C2(n12259), .A(n12258), .B(n12257), .ZN(
        n12260) );
  BUF_X1 U15588 ( .A(n12264), .Z(n12270) );
  BUF_X1 U15589 ( .A(n12265), .Z(n12266) );
  XNOR2_X2 U15590 ( .A(n12266), .B(n12270), .ZN(n16718) );
  INV_X1 U15591 ( .A(n13822), .ZN(n13833) );
  NAND2_X1 U15592 ( .A1(n16718), .A2(n13833), .ZN(n12290) );
  INV_X1 U15593 ( .A(n12266), .ZN(n12271) );
  INV_X1 U15594 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12272) );
  OAI22_X1 U15595 ( .A1(n12273), .A2(n20757), .B1(n12429), .B2(n12272), .ZN(
        n12278) );
  INV_X1 U15596 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12276) );
  INV_X1 U15597 ( .A(n12274), .ZN(n12275) );
  OR2_X4 U15598 ( .A1(n12288), .A2(n12280), .ZN(n20580) );
  NOR2_X1 U15599 ( .A1(n12278), .A2(n12277), .ZN(n12298) );
  INV_X1 U15600 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15092) );
  INV_X1 U15601 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12279) );
  OAI22_X1 U15602 ( .A1(n15092), .A2(n20526), .B1(n12426), .B2(n12279), .ZN(
        n12283) );
  INV_X1 U15603 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13006) );
  INV_X1 U15604 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12281) );
  NOR2_X1 U15605 ( .A1(n12283), .A2(n12282), .ZN(n12297) );
  INV_X1 U15606 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12284) );
  OAI22_X1 U15607 ( .A1(n12284), .A2(n14853), .B1(n12438), .B2(n20931), .ZN(
        n12287) );
  INV_X1 U15608 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12285) );
  INV_X1 U15609 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12302) );
  NOR2_X1 U15610 ( .A1(n12287), .A2(n12286), .ZN(n12296) );
  INV_X1 U15611 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12301) );
  OR2_X2 U15612 ( .A1(n12288), .A2(n12290), .ZN(n20614) );
  INV_X1 U15613 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12289) );
  INV_X1 U15614 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12292) );
  INV_X1 U15615 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13007) );
  NOR2_X1 U15616 ( .A1(n12294), .A2(n12293), .ZN(n12295) );
  AOI22_X1 U15617 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n15148), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12309) );
  INV_X1 U15618 ( .A(n12299), .ZN(n12300) );
  OAI22_X1 U15619 ( .A1(n15145), .A2(n12302), .B1(n15143), .B2(n12301), .ZN(
        n12306) );
  NAND2_X1 U15620 ( .A1(n15172), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n12304) );
  NAND2_X1 U15621 ( .A1(n12350), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n12303) );
  OAI211_X1 U15622 ( .C1(n13078), .C2(n20931), .A(n12304), .B(n12303), .ZN(
        n12305) );
  NOR2_X1 U15623 ( .A1(n12306), .A2(n12305), .ZN(n12308) );
  AND2_X2 U15624 ( .A1(n9728), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12362) );
  AND2_X2 U15625 ( .A1(n9721), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12412) );
  AOI22_X1 U15626 ( .A1(n12362), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12412), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12307) );
  INV_X1 U15627 ( .A(n12310), .ZN(n14698) );
  NAND2_X1 U15628 ( .A1(n9730), .A2(n12129), .ZN(n15179) );
  INV_X2 U15629 ( .A(n15179), .ZN(n15125) );
  AOI22_X1 U15630 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n15125), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12317) );
  AND2_X2 U15631 ( .A1(n12311), .A2(n12129), .ZN(n12341) );
  AND2_X2 U15632 ( .A1(n15323), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12525) );
  AOI22_X1 U15633 ( .A1(n12341), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12525), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12316) );
  AND2_X2 U15634 ( .A1(n15153), .A2(n12313), .ZN(n15171) );
  AOI22_X1 U15635 ( .A1(n12371), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n15171), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12315) );
  AND2_X2 U15636 ( .A1(n12311), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12524) );
  NAND2_X1 U15637 ( .A1(n12524), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n12314) );
  INV_X1 U15638 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12363) );
  INV_X1 U15639 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12320) );
  INV_X1 U15640 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12319) );
  OAI22_X1 U15641 ( .A1(n12320), .A2(n20580), .B1(n20757), .B2(n12319), .ZN(
        n12321) );
  NOR2_X1 U15642 ( .A1(n12322), .A2(n12321), .ZN(n12340) );
  INV_X1 U15643 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n15066) );
  INV_X1 U15644 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n20917) );
  OAI22_X1 U15645 ( .A1(n15066), .A2(n20526), .B1(n12438), .B2(n20917), .ZN(
        n12326) );
  INV_X1 U15646 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12324) );
  INV_X1 U15647 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12323) );
  OAI22_X1 U15648 ( .A1(n12324), .A2(n12429), .B1(n12426), .B2(n12323), .ZN(
        n12325) );
  NOR2_X1 U15649 ( .A1(n12326), .A2(n12325), .ZN(n12339) );
  INV_X1 U15650 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12969) );
  INV_X1 U15651 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12327) );
  OAI22_X1 U15652 ( .A1(n12969), .A2(n20460), .B1(n14853), .B2(n12327), .ZN(
        n12331) );
  INV_X1 U15653 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12329) );
  INV_X1 U15654 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12328) );
  NOR2_X1 U15655 ( .A1(n12331), .A2(n12330), .ZN(n12338) );
  INV_X1 U15656 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12333) );
  INV_X1 U15657 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12332) );
  OAI22_X1 U15658 ( .A1(n12333), .A2(n20494), .B1(n17579), .B2(n12332), .ZN(
        n12336) );
  INV_X1 U15659 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12334) );
  INV_X1 U15660 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12970) );
  NOR2_X1 U15661 ( .A1(n12336), .A2(n12335), .ZN(n12337) );
  AOI22_X1 U15662 ( .A1(n12371), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n15171), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12345) );
  NAND2_X1 U15663 ( .A1(n12524), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12344) );
  NAND2_X1 U15664 ( .A1(n12341), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12343) );
  NAND2_X1 U15665 ( .A1(n12525), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12342) );
  NAND2_X1 U15666 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12349) );
  NAND2_X1 U15667 ( .A1(n12362), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12348) );
  NAND2_X1 U15668 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12347) );
  NAND2_X1 U15669 ( .A1(n12412), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12346) );
  NAND4_X1 U15670 ( .A1(n12349), .A2(n12348), .A3(n12347), .A4(n12346), .ZN(
        n12356) );
  INV_X2 U15671 ( .A(n9783), .ZN(n15172) );
  AOI22_X1 U15672 ( .A1(n15172), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12350), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12354) );
  NAND2_X1 U15673 ( .A1(n15176), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12353) );
  NAND2_X1 U15674 ( .A1(n15177), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12352) );
  NAND2_X1 U15675 ( .A1(n15173), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12351) );
  NAND4_X1 U15676 ( .A1(n12354), .A2(n12353), .A3(n12352), .A4(n12351), .ZN(
        n12355) );
  NOR2_X1 U15677 ( .A1(n12356), .A2(n12355), .ZN(n12361) );
  INV_X1 U15678 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12358) );
  INV_X1 U15679 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12357) );
  OAI22_X1 U15680 ( .A1(n15181), .A2(n12358), .B1(n15179), .B2(n12357), .ZN(
        n12359) );
  INV_X1 U15681 ( .A(n12904), .ZN(n12587) );
  NAND2_X1 U15682 ( .A1(n12587), .A2(n15209), .ZN(n13582) );
  AOI22_X1 U15683 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n12362), .B1(
        n12379), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12370) );
  AOI22_X1 U15684 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n15148), .B1(
        n12451), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12369) );
  OAI22_X1 U15685 ( .A1(n12363), .A2(n15145), .B1(n15143), .B2(n17573), .ZN(
        n12367) );
  NAND2_X1 U15686 ( .A1(n15171), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12365) );
  NAND2_X1 U15687 ( .A1(n15172), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n12364) );
  OAI211_X1 U15688 ( .C1(n13078), .C2(n20917), .A(n12365), .B(n12364), .ZN(
        n12366) );
  NOR2_X1 U15689 ( .A1(n12367), .A2(n12366), .ZN(n12368) );
  NAND3_X1 U15690 ( .A1(n12370), .A2(n12369), .A3(n12368), .ZN(n12377) );
  AOI22_X1 U15691 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12341), .B1(
        n12524), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12375) );
  AOI22_X1 U15692 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n12412), .B1(
        n15125), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12374) );
  AOI22_X1 U15693 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12371), .B1(
        n12350), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12373) );
  NAND2_X1 U15694 ( .A1(n12525), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12372) );
  NAND4_X1 U15695 ( .A1(n12375), .A2(n12374), .A3(n12373), .A4(n12372), .ZN(
        n12376) );
  INV_X1 U15696 ( .A(n12909), .ZN(n12378) );
  AOI22_X1 U15697 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n12379), .B1(
        n15148), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12386) );
  INV_X1 U15698 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12991) );
  NAND2_X1 U15699 ( .A1(n15172), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n12381) );
  NAND2_X1 U15700 ( .A1(n12350), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n12380) );
  OAI211_X1 U15701 ( .C1(n15143), .C2(n12991), .A(n12381), .B(n12380), .ZN(
        n12382) );
  INV_X1 U15702 ( .A(n12382), .ZN(n12385) );
  AOI22_X1 U15703 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n15177), .B1(
        n15173), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12384) );
  AOI22_X1 U15704 ( .A1(n12362), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12412), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12383) );
  NAND4_X1 U15705 ( .A1(n12386), .A2(n12385), .A3(n12384), .A4(n12383), .ZN(
        n12392) );
  AOI22_X1 U15706 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n15125), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12390) );
  AOI22_X1 U15707 ( .A1(n12524), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12525), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12389) );
  AOI22_X1 U15708 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n12371), .B1(
        n15171), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12388) );
  NAND2_X1 U15709 ( .A1(n12341), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n12387) );
  NAND4_X1 U15710 ( .A1(n12390), .A2(n12389), .A3(n12388), .A4(n12387), .ZN(
        n12391) );
  INV_X1 U15711 ( .A(n12591), .ZN(n12397) );
  NAND2_X1 U15712 ( .A1(n12398), .A2(n12397), .ZN(n12393) );
  NAND2_X1 U15713 ( .A1(n13582), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12394) );
  XNOR2_X1 U15714 ( .A(n12904), .B(n12909), .ZN(n12395) );
  XNOR2_X1 U15715 ( .A(n12394), .B(n12395), .ZN(n13604) );
  NAND2_X1 U15716 ( .A1(n13604), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13603) );
  INV_X1 U15717 ( .A(n12394), .ZN(n13583) );
  NAND2_X1 U15718 ( .A1(n13583), .A2(n12395), .ZN(n12396) );
  NAND2_X1 U15719 ( .A1(n13603), .A2(n12396), .ZN(n12399) );
  INV_X1 U15720 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21972) );
  XNOR2_X1 U15721 ( .A(n12399), .B(n21972), .ZN(n13595) );
  XNOR2_X1 U15722 ( .A(n12398), .B(n12397), .ZN(n13594) );
  NAND2_X1 U15723 ( .A1(n13595), .A2(n13594), .ZN(n13972) );
  NAND2_X1 U15724 ( .A1(n12399), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12400) );
  NAND2_X1 U15725 ( .A1(n13972), .A2(n12400), .ZN(n12402) );
  XNOR2_X1 U15726 ( .A(n12402), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n17249) );
  INV_X1 U15727 ( .A(n17249), .ZN(n12401) );
  NAND2_X1 U15728 ( .A1(n12402), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12403) );
  AOI22_X1 U15729 ( .A1(n12362), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12379), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12411) );
  AOI22_X1 U15730 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n15148), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12410) );
  INV_X1 U15731 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12406) );
  NAND2_X1 U15732 ( .A1(n15171), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12405) );
  NAND2_X1 U15733 ( .A1(n15172), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n12404) );
  OAI211_X1 U15734 ( .C1(n13078), .C2(n12406), .A(n12405), .B(n12404), .ZN(
        n12407) );
  INV_X1 U15735 ( .A(n12407), .ZN(n12409) );
  AOI22_X1 U15736 ( .A1(n15177), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n15176), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12408) );
  NAND4_X1 U15737 ( .A1(n12411), .A2(n12410), .A3(n12409), .A4(n12408), .ZN(
        n12418) );
  AOI22_X1 U15738 ( .A1(n12524), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12341), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12416) );
  AOI22_X1 U15739 ( .A1(n15125), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12412), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12415) );
  AOI22_X1 U15740 ( .A1(n12371), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12350), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12414) );
  NAND2_X1 U15741 ( .A1(n12525), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n12413) );
  NAND4_X1 U15742 ( .A1(n12416), .A2(n12415), .A3(n12414), .A4(n12413), .ZN(
        n12417) );
  INV_X1 U15743 ( .A(n12934), .ZN(n12419) );
  NAND2_X1 U15744 ( .A1(n12420), .A2(n12419), .ZN(n12421) );
  INV_X1 U15745 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n22037) );
  INV_X1 U15746 ( .A(n12422), .ZN(n12424) );
  NAND2_X1 U15747 ( .A1(n12424), .A2(n12423), .ZN(n12425) );
  INV_X1 U15748 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12428) );
  INV_X1 U15749 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12427) );
  OAI22_X1 U15750 ( .A1(n12428), .A2(n20551), .B1(n12426), .B2(n12427), .ZN(
        n12432) );
  INV_X1 U15751 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15119) );
  INV_X1 U15752 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12430) );
  OAI22_X1 U15753 ( .A1(n15119), .A2(n20526), .B1(n12429), .B2(n12430), .ZN(
        n12431) );
  NOR2_X1 U15754 ( .A1(n12432), .A2(n12431), .ZN(n12450) );
  INV_X1 U15755 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14494) );
  INV_X1 U15756 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12434) );
  OAI22_X1 U15757 ( .A1(n14494), .A2(n12433), .B1(n20580), .B2(n12434), .ZN(
        n12437) );
  INV_X1 U15758 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12435) );
  INV_X1 U15759 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13040) );
  NOR2_X1 U15760 ( .A1(n12437), .A2(n12436), .ZN(n12449) );
  INV_X1 U15761 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12439) );
  INV_X1 U15762 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12458) );
  INV_X1 U15763 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12455) );
  INV_X1 U15764 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12440) );
  OAI22_X1 U15765 ( .A1(n12455), .A2(n20646), .B1(n20832), .B2(n12440), .ZN(
        n12441) );
  NOR2_X1 U15766 ( .A1(n12442), .A2(n12441), .ZN(n12448) );
  INV_X1 U15767 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13039) );
  INV_X1 U15768 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12452) );
  OAI22_X1 U15769 ( .A1(n13039), .A2(n20460), .B1(n20757), .B2(n12452), .ZN(
        n12446) );
  INV_X1 U15770 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12444) );
  INV_X1 U15771 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12443) );
  OAI22_X1 U15772 ( .A1(n12444), .A2(n20494), .B1(n17579), .B2(n12443), .ZN(
        n12445) );
  NOR2_X1 U15773 ( .A1(n12446), .A2(n12445), .ZN(n12447) );
  INV_X1 U15774 ( .A(n12451), .ZN(n12453) );
  OAI22_X1 U15775 ( .A1(n12435), .A2(n15181), .B1(n12453), .B2(n12452), .ZN(
        n12454) );
  INV_X1 U15776 ( .A(n12454), .ZN(n12463) );
  AOI22_X1 U15777 ( .A1(n12362), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12379), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12462) );
  OAI22_X1 U15778 ( .A1(n15145), .A2(n12455), .B1(n15143), .B2(n14494), .ZN(
        n12460) );
  NAND2_X1 U15779 ( .A1(n15171), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n12457) );
  NAND2_X1 U15780 ( .A1(n15172), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n12456) );
  OAI211_X1 U15781 ( .C1(n13078), .C2(n12458), .A(n12457), .B(n12456), .ZN(
        n12459) );
  NOR2_X1 U15782 ( .A1(n12460), .A2(n12459), .ZN(n12461) );
  NAND3_X1 U15783 ( .A1(n12463), .A2(n12462), .A3(n12461), .ZN(n12469) );
  AOI22_X1 U15784 ( .A1(n12524), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12341), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12467) );
  AOI22_X1 U15785 ( .A1(n15125), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12412), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12466) );
  AOI22_X1 U15786 ( .A1(n12371), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12350), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12465) );
  NAND2_X1 U15787 ( .A1(n12525), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n12464) );
  NAND4_X1 U15788 ( .A1(n12467), .A2(n12466), .A3(n12465), .A4(n12464), .ZN(
        n12468) );
  NAND2_X1 U15789 ( .A1(n12624), .A2(n15209), .ZN(n12470) );
  INV_X1 U15790 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12472) );
  INV_X1 U15791 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12491) );
  INV_X1 U15792 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n15141) );
  INV_X1 U15793 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12488) );
  OAI22_X1 U15794 ( .A1(n15141), .A2(n20551), .B1(n20646), .B2(n12488), .ZN(
        n12473) );
  NOR2_X1 U15795 ( .A1(n12474), .A2(n12473), .ZN(n12487) );
  INV_X1 U15796 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n15139) );
  INV_X1 U15797 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n15135) );
  OAI22_X1 U15798 ( .A1(n15139), .A2(n20526), .B1(n12426), .B2(n15135), .ZN(
        n12477) );
  INV_X1 U15799 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13061) );
  INV_X1 U15800 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12475) );
  OAI22_X1 U15801 ( .A1(n13061), .A2(n20460), .B1(n20832), .B2(n12475), .ZN(
        n12476) );
  NOR2_X1 U15802 ( .A1(n12477), .A2(n12476), .ZN(n12486) );
  INV_X1 U15803 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n15132) );
  INV_X1 U15804 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n15144) );
  OAI22_X1 U15805 ( .A1(n15132), .A2(n20757), .B1(n12429), .B2(n15144), .ZN(
        n12480) );
  INV_X1 U15806 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12478) );
  OAI22_X1 U15807 ( .A1(n12478), .A2(n20580), .B1(n17579), .B2(n20884), .ZN(
        n12479) );
  NOR2_X1 U15808 ( .A1(n12480), .A2(n12479), .ZN(n12485) );
  INV_X1 U15809 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n20449) );
  INV_X1 U15810 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12481) );
  OAI22_X1 U15811 ( .A1(n20449), .A2(n12433), .B1(n20614), .B2(n12481), .ZN(
        n12483) );
  INV_X1 U15812 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n15142) );
  INV_X1 U15813 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13058) );
  NOR2_X1 U15814 ( .A1(n12483), .A2(n12482), .ZN(n12484) );
  NAND4_X1 U15815 ( .A1(n12487), .A2(n12486), .A3(n12485), .A4(n12484), .ZN(
        n12504) );
  AOI22_X1 U15816 ( .A1(n12362), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12379), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12496) );
  OAI22_X1 U15817 ( .A1(n15145), .A2(n12488), .B1(n15143), .B2(n20449), .ZN(
        n12493) );
  NAND2_X1 U15818 ( .A1(n15171), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n12490) );
  NAND2_X1 U15819 ( .A1(n15172), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n12489) );
  OAI211_X1 U15820 ( .C1(n13078), .C2(n12491), .A(n12490), .B(n12489), .ZN(
        n12492) );
  NOR2_X1 U15821 ( .A1(n12493), .A2(n12492), .ZN(n12495) );
  AOI22_X1 U15822 ( .A1(n15148), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n15125), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12494) );
  NAND3_X1 U15823 ( .A1(n12496), .A2(n12495), .A3(n12494), .ZN(n12502) );
  AOI22_X1 U15824 ( .A1(n12524), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12341), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12500) );
  AOI22_X1 U15825 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12412), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12499) );
  AOI22_X1 U15826 ( .A1(n12371), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12350), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12498) );
  NAND2_X1 U15827 ( .A1(n12525), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n12497) );
  NAND4_X1 U15828 ( .A1(n12500), .A2(n12499), .A3(n12498), .A4(n12497), .ZN(
        n12501) );
  NAND2_X1 U15829 ( .A1(n12943), .A2(n15209), .ZN(n12503) );
  INV_X1 U15830 ( .A(n12514), .ZN(n12505) );
  INV_X1 U15831 ( .A(n12682), .ZN(n12507) );
  NAND2_X1 U15832 ( .A1(n12508), .A2(n12507), .ZN(n12511) );
  NAND2_X1 U15833 ( .A1(n12685), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12509) );
  NAND2_X1 U15834 ( .A1(n12682), .A2(n12509), .ZN(n12510) );
  NAND2_X1 U15835 ( .A1(n12511), .A2(n12510), .ZN(n12512) );
  NAND2_X1 U15836 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n12519) );
  NAND2_X1 U15837 ( .A1(n12362), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n12518) );
  NAND2_X1 U15838 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n12517) );
  NAND2_X1 U15839 ( .A1(n12412), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n12516) );
  AOI22_X1 U15840 ( .A1(n15148), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n15125), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12537) );
  INV_X1 U15841 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12522) );
  NAND2_X1 U15842 ( .A1(n15171), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n12521) );
  NAND2_X1 U15843 ( .A1(n12371), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n12520) );
  OAI211_X1 U15844 ( .C1(n12523), .C2(n12522), .A(n12521), .B(n12520), .ZN(
        n12530) );
  INV_X1 U15845 ( .A(n12524), .ZN(n12528) );
  INV_X1 U15846 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12527) );
  INV_X1 U15847 ( .A(n12525), .ZN(n15136) );
  INV_X1 U15848 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12526) );
  OAI22_X1 U15849 ( .A1(n12528), .A2(n12527), .B1(n15136), .B2(n12526), .ZN(
        n12529) );
  NOR2_X1 U15850 ( .A1(n12530), .A2(n12529), .ZN(n12536) );
  AOI22_X1 U15851 ( .A1(n15172), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12350), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12534) );
  NAND2_X1 U15852 ( .A1(n15173), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n12533) );
  NAND2_X1 U15853 ( .A1(n15176), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12532) );
  NAND2_X1 U15854 ( .A1(n15177), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n12531) );
  AND4_X2 U15855 ( .A1(n12538), .A2(n12537), .A3(n12536), .A4(n12535), .ZN(
        n12627) );
  INV_X1 U15856 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17474) );
  NAND2_X1 U15857 ( .A1(n17206), .A2(n17474), .ZN(n12539) );
  NAND4_X1 U15858 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A4(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12544) );
  NAND2_X1 U15859 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17388) );
  NOR2_X1 U15860 ( .A1(n12544), .A2(n17388), .ZN(n17381) );
  AND3_X1 U15861 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17325) );
  NAND2_X1 U15862 ( .A1(n17381), .A2(n17325), .ZN(n13360) );
  NAND3_X1 U15863 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12545) );
  OR2_X1 U15864 ( .A1(n13360), .A2(n12545), .ZN(n13368) );
  AND2_X1 U15865 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n13159) );
  NAND2_X1 U15866 ( .A1(n13159), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12546) );
  NOR2_X1 U15867 ( .A1(n13368), .A2(n12546), .ZN(n13170) );
  INV_X1 U15868 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17266) );
  INV_X1 U15869 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17267) );
  INV_X1 U15870 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n13197) );
  MUX2_X1 U15871 ( .A(n22046), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n12588) );
  NAND2_X1 U15872 ( .A1(n12588), .A2(n12552), .ZN(n12548) );
  NAND2_X1 U15873 ( .A1(n22046), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12547) );
  XNOR2_X1 U15874 ( .A(n12559), .B(n12558), .ZN(n12579) );
  INV_X1 U15875 ( .A(n12579), .ZN(n12590) );
  OAI21_X1 U15876 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21083), .A(
        n12549), .ZN(n12581) );
  INV_X1 U15877 ( .A(n12581), .ZN(n12586) );
  NAND2_X1 U15878 ( .A1(n12588), .A2(n12586), .ZN(n12550) );
  NAND2_X1 U15879 ( .A1(n12207), .A2(n12550), .ZN(n12556) );
  XNOR2_X1 U15880 ( .A(n12588), .B(n12552), .ZN(n12580) );
  INV_X1 U15881 ( .A(n12580), .ZN(n12554) );
  OAI21_X1 U15882 ( .B1(n12581), .B2(n12580), .A(n12579), .ZN(n12553) );
  OAI211_X1 U15883 ( .C1(n12551), .C2(n12554), .A(n9941), .B(n12553), .ZN(
        n12555) );
  AND2_X1 U15884 ( .A1(n12556), .A2(n12555), .ZN(n12557) );
  NAND2_X1 U15885 ( .A1(n21065), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12560) );
  NAND3_X1 U15886 ( .A1(n12569), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A3(
        n14742), .ZN(n12567) );
  INV_X1 U15887 ( .A(n12563), .ZN(n12564) );
  XNOR2_X1 U15888 ( .A(n12565), .B(n12564), .ZN(n12566) );
  NAND2_X1 U15889 ( .A1(n12567), .A2(n12566), .ZN(n12594) );
  NAND2_X1 U15890 ( .A1(n18043), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12568) );
  NAND2_X1 U15891 ( .A1(n12569), .A2(n12568), .ZN(n12571) );
  NAND2_X1 U15892 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n14742), .ZN(
        n12570) );
  NOR2_X1 U15893 ( .A1(n12572), .A2(n12574), .ZN(n12573) );
  OAI211_X1 U15894 ( .C1(n12575), .C2(n14870), .A(n13627), .B(n12600), .ZN(
        n12618) );
  INV_X1 U15895 ( .A(n13627), .ZN(n12576) );
  NAND2_X2 U15896 ( .A1(n20976), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n21030) );
  NOR2_X1 U15897 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n20236) );
  INV_X1 U15898 ( .A(n20236), .ZN(n20970) );
  NAND3_X1 U15899 ( .A1(n20965), .A2(n21030), .A3(n20970), .ZN(n20964) );
  NOR2_X1 U15900 ( .A1(n20964), .A2(n20959), .ZN(n13609) );
  NAND3_X1 U15901 ( .A1(n12576), .A2(n13609), .A3(n12174), .ZN(n12617) );
  OR2_X1 U15902 ( .A1(n12577), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13619) );
  INV_X1 U15903 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n12578) );
  OAI21_X1 U15904 ( .B1(n12379), .B2(n13619), .A(n12578), .ZN(n21076) );
  OR2_X1 U15905 ( .A1(n12594), .A2(n12579), .ZN(n12582) );
  NOR2_X1 U15906 ( .A1(n12582), .A2(n12581), .ZN(n12583) );
  NOR2_X1 U15907 ( .A1(n14732), .A2(n12583), .ZN(n12584) );
  MUX2_X1 U15908 ( .A(n21076), .B(n12584), .S(n17538), .Z(n18134) );
  NAND2_X1 U15909 ( .A1(n18134), .A2(n13145), .ZN(n21089) );
  NOR2_X1 U15910 ( .A1(n21089), .A2(n12585), .ZN(n12615) );
  NOR2_X1 U15911 ( .A1(n12585), .A2(n9941), .ZN(n21088) );
  INV_X1 U15912 ( .A(n21088), .ZN(n14738) );
  MUX2_X1 U15913 ( .A(n12587), .B(n12586), .S(n12589), .Z(n12659) );
  NAND2_X1 U15914 ( .A1(n12659), .A2(n12588), .ZN(n12593) );
  MUX2_X1 U15915 ( .A(n12591), .B(n12590), .S(n12589), .Z(n12620) );
  NAND2_X1 U15916 ( .A1(n12593), .A2(n12592), .ZN(n12596) );
  INV_X1 U15917 ( .A(n12594), .ZN(n12595) );
  NAND2_X1 U15918 ( .A1(n12596), .A2(n12595), .ZN(n12599) );
  AND2_X1 U15919 ( .A1(n12597), .A2(n15209), .ZN(n12598) );
  NAND2_X1 U15920 ( .A1(n12599), .A2(n12598), .ZN(n21087) );
  NOR2_X1 U15921 ( .A1(n14732), .A2(n20959), .ZN(n13610) );
  INV_X1 U15922 ( .A(n20964), .ZN(n14733) );
  NAND3_X1 U15923 ( .A1(n13610), .A2(n12611), .A3(n14733), .ZN(n12610) );
  NAND2_X1 U15924 ( .A1(n15209), .A2(n12600), .ZN(n12601) );
  NAND2_X1 U15925 ( .A1(n12601), .A2(n9941), .ZN(n12602) );
  NAND3_X1 U15926 ( .A1(n12603), .A2(n20433), .A3(n12602), .ZN(n12608) );
  NAND2_X1 U15927 ( .A1(n12604), .A2(n12905), .ZN(n12605) );
  NAND2_X1 U15928 ( .A1(n12605), .A2(n16419), .ZN(n13147) );
  AOI21_X1 U15929 ( .B1(n9815), .B2(n12608), .A(n12607), .ZN(n12609) );
  AND2_X1 U15930 ( .A1(n12610), .A2(n12609), .ZN(n13613) );
  MUX2_X1 U15931 ( .A(n12611), .B(n12174), .S(n12551), .Z(n12612) );
  NAND2_X1 U15932 ( .A1(n12612), .A2(n13610), .ZN(n12613) );
  OAI211_X1 U15933 ( .C1(n14738), .C2(n21087), .A(n13613), .B(n12613), .ZN(
        n12614) );
  NOR2_X1 U15934 ( .A1(n12615), .A2(n12614), .ZN(n12616) );
  NAND3_X1 U15935 ( .A1(n12618), .A2(n12617), .A3(n12616), .ZN(n12619) );
  NAND3_X1 U15936 ( .A1(n17538), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n18142) );
  NOR2_X1 U15937 ( .A1(P2_EBX_REG_0__SCAN_IN), .A2(P2_EBX_REG_1__SCAN_IN), 
        .ZN(n12622) );
  MUX2_X1 U15938 ( .A(n12622), .B(n12909), .S(n9987), .Z(n12666) );
  INV_X1 U15939 ( .A(n12929), .ZN(n12623) );
  INV_X1 U15940 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n20334) );
  MUX2_X1 U15941 ( .A(n20334), .B(n12934), .S(n9987), .Z(n12656) );
  MUX2_X1 U15942 ( .A(P2_EBX_REG_5__SCAN_IN), .B(n12624), .S(n9987), .Z(n12674) );
  INV_X1 U15943 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n12626) );
  INV_X1 U15944 ( .A(n12943), .ZN(n12625) );
  MUX2_X1 U15945 ( .A(n12626), .B(n12625), .S(n9987), .Z(n12687) );
  MUX2_X1 U15946 ( .A(P2_EBX_REG_7__SCAN_IN), .B(n12627), .S(n9987), .Z(n12694) );
  INV_X1 U15947 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n21858) );
  NOR2_X1 U15948 ( .A1(n9987), .A2(n21858), .ZN(n12692) );
  INV_X1 U15949 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n16646) );
  NAND2_X1 U15950 ( .A1(n12631), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12630) );
  NAND2_X1 U15951 ( .A1(n12631), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n12730) );
  OAI21_X1 U15952 ( .B1(P2_EBX_REG_15__SCAN_IN), .B2(P2_EBX_REG_14__SCAN_IN), 
        .A(n12631), .ZN(n12632) );
  OAI21_X1 U15953 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(P2_EBX_REG_16__SCAN_IN), 
        .A(n12631), .ZN(n12633) );
  OAI21_X1 U15954 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(P2_EBX_REG_18__SCAN_IN), 
        .A(n12631), .ZN(n12634) );
  NOR2_X2 U15955 ( .A1(n12745), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12706) );
  INV_X1 U15956 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n12635) );
  NAND2_X1 U15957 ( .A1(n12706), .A2(n12635), .ZN(n12768) );
  NAND2_X1 U15958 ( .A1(n12768), .A2(n12726), .ZN(n12708) );
  NAND2_X1 U15959 ( .A1(n12631), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12766) );
  NAND2_X1 U15960 ( .A1(n12708), .A2(n12766), .ZN(n12770) );
  INV_X1 U15961 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n12868) );
  NOR2_X1 U15962 ( .A1(n9987), .A2(n12868), .ZN(n12651) );
  INV_X1 U15963 ( .A(n12651), .ZN(n12636) );
  INV_X1 U15964 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n16767) );
  NAND2_X1 U15965 ( .A1(n12643), .A2(n16767), .ZN(n12781) );
  NAND2_X1 U15966 ( .A1(n12781), .A2(n12726), .ZN(n13242) );
  NAND2_X1 U15967 ( .A1(n12631), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12779) );
  NAND2_X1 U15968 ( .A1(n13242), .A2(n12779), .ZN(n12783) );
  INV_X1 U15969 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n16432) );
  NOR2_X1 U15970 ( .A1(n9987), .A2(n16432), .ZN(n12777) );
  INV_X1 U15971 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n22023) );
  NOR2_X1 U15972 ( .A1(n9987), .A2(n22023), .ZN(n12793) );
  NOR2_X2 U15973 ( .A1(n9778), .A2(n12793), .ZN(n13241) );
  AND2_X1 U15974 ( .A1(n12631), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12639) );
  XNOR2_X1 U15975 ( .A(n13241), .B(n12639), .ZN(n13338) );
  AOI21_X1 U15976 ( .B1(n13338), .B2(n10337), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13239) );
  NAND3_X1 U15977 ( .A1(n13338), .A2(n12946), .A3(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13238) );
  NAND2_X1 U15978 ( .A1(n10412), .A2(n13238), .ZN(n12795) );
  NAND2_X1 U15979 ( .A1(n12631), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n12640) );
  OAI211_X1 U15980 ( .C1(n12643), .C2(n12640), .A(n12726), .B(n12781), .ZN(
        n12785) );
  OR2_X1 U15981 ( .A1(n12785), .A2(n12627), .ZN(n12641) );
  NAND3_X1 U15982 ( .A1(n12647), .A2(n12631), .A3(P2_EBX_REG_25__SCAN_IN), 
        .ZN(n12642) );
  NAND2_X1 U15983 ( .A1(n12642), .A2(n12726), .ZN(n12644) );
  OR2_X1 U15984 ( .A1(n12644), .A2(n12643), .ZN(n12787) );
  AND2_X1 U15985 ( .A1(n12631), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12646) );
  INV_X1 U15986 ( .A(n12726), .ZN(n12645) );
  AOI21_X1 U15987 ( .B1(n12653), .B2(n12646), .A(n12645), .ZN(n12648) );
  NAND2_X1 U15988 ( .A1(n12648), .A2(n12647), .ZN(n16485) );
  NAND2_X1 U15989 ( .A1(n17018), .A2(n10338), .ZN(n12649) );
  AND2_X1 U15990 ( .A1(n17008), .A2(n12649), .ZN(n12650) );
  NAND2_X1 U15991 ( .A1(n12770), .A2(n12651), .ZN(n12652) );
  NAND2_X1 U15992 ( .A1(n12653), .A2(n12652), .ZN(n16500) );
  OR2_X1 U15993 ( .A1(n16500), .A2(n12627), .ZN(n12654) );
  XNOR2_X1 U15994 ( .A(n12654), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17026) );
  XNOR2_X1 U15995 ( .A(n12655), .B(n12656), .ZN(n20337) );
  NAND2_X1 U15996 ( .A1(n12664), .A2(n12657), .ZN(n12658) );
  NAND2_X1 U15997 ( .A1(n10060), .A2(n12658), .ZN(n16695) );
  MUX2_X1 U15998 ( .A(n12659), .B(P2_EBX_REG_0__SCAN_IN), .S(n12631), .Z(
        n16735) );
  NAND2_X1 U15999 ( .A1(n16735), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13586) );
  INV_X1 U16000 ( .A(n13586), .ZN(n12661) );
  AND3_X1 U16001 ( .A1(n12631), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n12660) );
  NOR2_X1 U16002 ( .A1(n12666), .A2(n12660), .ZN(n12662) );
  NAND2_X1 U16003 ( .A1(n12661), .A2(n12662), .ZN(n13601) );
  INV_X1 U16004 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14087) );
  NAND2_X1 U16005 ( .A1(n13601), .A2(n14087), .ZN(n12663) );
  INV_X1 U16006 ( .A(n12662), .ZN(n16724) );
  NAND2_X1 U16007 ( .A1(n13586), .A2(n16724), .ZN(n13600) );
  AND2_X1 U16008 ( .A1(n12663), .A2(n13600), .ZN(n13592) );
  OAI21_X1 U16009 ( .B1(n12666), .B2(n12665), .A(n12664), .ZN(n16711) );
  XNOR2_X1 U16010 ( .A(n16711), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13591) );
  NAND2_X1 U16011 ( .A1(n13592), .A2(n13591), .ZN(n12669) );
  INV_X1 U16012 ( .A(n16711), .ZN(n12667) );
  NAND2_X1 U16013 ( .A1(n12667), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12668) );
  NAND2_X1 U16014 ( .A1(n12669), .A2(n12668), .ZN(n17240) );
  NAND2_X1 U16015 ( .A1(n20337), .A2(n22037), .ZN(n12672) );
  OAI21_X1 U16016 ( .B1(n17240), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n12672), .ZN(n12670) );
  INV_X1 U16017 ( .A(n12670), .ZN(n12671) );
  NAND3_X1 U16018 ( .A1(n17240), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n12672), .ZN(n12673) );
  XNOR2_X1 U16019 ( .A(n12675), .B(n12674), .ZN(n20322) );
  AND2_X1 U16020 ( .A1(n20322), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12677) );
  INV_X1 U16021 ( .A(n12677), .ZN(n12676) );
  OAI21_X1 U16022 ( .B1(n12627), .B2(n12506), .A(n20322), .ZN(n12678) );
  OAI21_X1 U16023 ( .B1(n20322), .B2(n12506), .A(n12678), .ZN(n12679) );
  INV_X1 U16024 ( .A(n20322), .ZN(n12681) );
  AOI21_X1 U16025 ( .B1(n20322), .B2(n10337), .A(n12506), .ZN(n12680) );
  OAI21_X1 U16026 ( .B1(n12682), .B2(n12681), .A(n12680), .ZN(n12683) );
  OR2_X1 U16027 ( .A1(n12688), .A2(n12687), .ZN(n12689) );
  AND2_X1 U16028 ( .A1(n12686), .A2(n12689), .ZN(n16682) );
  INV_X1 U16029 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17494) );
  NAND2_X1 U16030 ( .A1(n12629), .A2(n12692), .ZN(n12693) );
  NAND2_X1 U16031 ( .A1(n12696), .A2(n12693), .ZN(n16652) );
  NOR2_X1 U16032 ( .A1(n16652), .A2(n12627), .ZN(n12700) );
  NAND2_X1 U16033 ( .A1(n12700), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17195) );
  XNOR2_X1 U16034 ( .A(n12686), .B(n10503), .ZN(n16665) );
  NAND2_X1 U16035 ( .A1(n16665), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17209) );
  AND2_X1 U16036 ( .A1(n17195), .A2(n17209), .ZN(n17180) );
  NAND2_X1 U16037 ( .A1(n12631), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12697) );
  MUX2_X1 U16038 ( .A(n12631), .B(n12697), .S(n12696), .Z(n12699) );
  INV_X1 U16039 ( .A(n12728), .ZN(n12698) );
  NAND2_X1 U16040 ( .A1(n12699), .A2(n12698), .ZN(n20308) );
  INV_X1 U16041 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17456) );
  OAI21_X1 U16042 ( .B1(n20308), .B2(n12627), .A(n17456), .ZN(n17184) );
  INV_X1 U16043 ( .A(n12700), .ZN(n12701) );
  INV_X1 U16044 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17469) );
  NAND2_X1 U16045 ( .A1(n12701), .A2(n17469), .ZN(n17194) );
  INV_X1 U16046 ( .A(n16665), .ZN(n12702) );
  NAND2_X1 U16047 ( .A1(n12702), .A2(n17474), .ZN(n17208) );
  AND2_X1 U16048 ( .A1(n17194), .A2(n17208), .ZN(n17181) );
  AND2_X1 U16049 ( .A1(n17184), .A2(n17181), .ZN(n12703) );
  NAND2_X1 U16050 ( .A1(n12631), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n12705) );
  NOR2_X1 U16051 ( .A1(n12706), .A2(n12705), .ZN(n12707) );
  OR2_X1 U16052 ( .A1(n12708), .A2(n12707), .ZN(n16529) );
  INV_X1 U16053 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n13370) );
  NAND2_X1 U16054 ( .A1(n12747), .A2(n13370), .ZN(n13356) );
  NAND2_X1 U16055 ( .A1(n12631), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12709) );
  MUX2_X1 U16056 ( .A(n12709), .B(n12631), .S(n12734), .Z(n12710) );
  INV_X1 U16057 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n16557) );
  NAND2_X1 U16058 ( .A1(n12734), .A2(n16557), .ZN(n12712) );
  AND2_X1 U16059 ( .A1(n12710), .A2(n12712), .ZN(n16564) );
  NAND2_X1 U16060 ( .A1(n16564), .A2(n12946), .ZN(n12763) );
  INV_X1 U16061 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17328) );
  NAND2_X1 U16062 ( .A1(n12763), .A2(n17328), .ZN(n17075) );
  AND2_X1 U16063 ( .A1(n12631), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n12711) );
  NAND2_X1 U16064 ( .A1(n12712), .A2(n12711), .ZN(n12713) );
  NAND2_X1 U16065 ( .A1(n12713), .A2(n12745), .ZN(n20264) );
  OR2_X1 U16066 ( .A1(n20264), .A2(n12627), .ZN(n12714) );
  INV_X1 U16067 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17340) );
  NAND2_X1 U16068 ( .A1(n12714), .A2(n17340), .ZN(n17067) );
  NAND2_X1 U16069 ( .A1(n12631), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n12715) );
  INV_X1 U16070 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n12847) );
  NAND2_X1 U16071 ( .A1(n12717), .A2(n12847), .ZN(n12735) );
  OAI211_X1 U16072 ( .C1(n12717), .C2(n12715), .A(n12726), .B(n12735), .ZN(
        n16592) );
  OR2_X1 U16073 ( .A1(n16592), .A2(n12627), .ZN(n12716) );
  XNOR2_X1 U16074 ( .A(n12716), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13350) );
  INV_X1 U16075 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n16606) );
  OR2_X1 U16076 ( .A1(n20278), .A2(n12627), .ZN(n12718) );
  INV_X1 U16077 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17380) );
  NAND2_X1 U16078 ( .A1(n12718), .A2(n17380), .ZN(n17110) );
  AND3_X1 U16079 ( .A1(n12719), .A2(n12631), .A3(P2_EBX_REG_12__SCAN_IN), .ZN(
        n12720) );
  NOR2_X1 U16080 ( .A1(n12731), .A2(n12720), .ZN(n16616) );
  NAND2_X1 U16081 ( .A1(n16616), .A2(n12946), .ZN(n12721) );
  INV_X1 U16082 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17418) );
  NAND2_X1 U16083 ( .A1(n12721), .A2(n17418), .ZN(n17145) );
  AND3_X1 U16084 ( .A1(n12722), .A2(n12631), .A3(P2_EBX_REG_11__SCAN_IN), .ZN(
        n12723) );
  NOR2_X1 U16085 ( .A1(n12724), .A2(n12723), .ZN(n16629) );
  NAND2_X1 U16086 ( .A1(n16629), .A2(n12946), .ZN(n12725) );
  INV_X1 U16087 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17431) );
  NAND2_X1 U16088 ( .A1(n12725), .A2(n17431), .ZN(n17154) );
  AND2_X1 U16089 ( .A1(n17145), .A2(n17154), .ZN(n13346) );
  NAND2_X1 U16090 ( .A1(n12631), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n12727) );
  OAI211_X1 U16091 ( .C1(n12728), .C2(n12727), .A(n12726), .B(n12722), .ZN(
        n16643) );
  OR2_X1 U16092 ( .A1(n16643), .A2(n12627), .ZN(n12729) );
  INV_X1 U16093 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17432) );
  NAND2_X1 U16094 ( .A1(n12729), .A2(n17432), .ZN(n17168) );
  NOR2_X1 U16095 ( .A1(n12731), .A2(n12730), .ZN(n12732) );
  NOR2_X1 U16096 ( .A1(n9803), .A2(n12732), .ZN(n12750) );
  NAND2_X1 U16097 ( .A1(n12750), .A2(n12946), .ZN(n12733) );
  INV_X1 U16098 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17402) );
  NAND2_X1 U16099 ( .A1(n12733), .A2(n17402), .ZN(n17132) );
  AND4_X1 U16100 ( .A1(n17110), .A2(n13346), .A3(n17168), .A4(n17132), .ZN(
        n12743) );
  INV_X1 U16101 ( .A(n12734), .ZN(n12737) );
  NAND3_X1 U16102 ( .A1(n12735), .A2(n12631), .A3(P2_EBX_REG_17__SCAN_IN), 
        .ZN(n12736) );
  NAND2_X1 U16103 ( .A1(n12737), .A2(n12736), .ZN(n16574) );
  OR2_X1 U16104 ( .A1(n16574), .A2(n12627), .ZN(n12738) );
  INV_X1 U16105 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21906) );
  NAND2_X1 U16106 ( .A1(n12738), .A2(n21906), .ZN(n13353) );
  NAND2_X1 U16107 ( .A1(n12631), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n12739) );
  MUX2_X1 U16108 ( .A(n12739), .B(n12631), .S(n9803), .Z(n12741) );
  AND2_X1 U16109 ( .A1(n12741), .A2(n12740), .ZN(n16604) );
  NAND2_X1 U16110 ( .A1(n16604), .A2(n12946), .ZN(n12761) );
  INV_X1 U16111 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12742) );
  NAND2_X1 U16112 ( .A1(n12761), .A2(n12742), .ZN(n17121) );
  NAND2_X1 U16113 ( .A1(n12631), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12744) );
  XNOR2_X1 U16114 ( .A(n12745), .B(n12744), .ZN(n16548) );
  NAND2_X1 U16115 ( .A1(n16548), .A2(n12946), .ZN(n12746) );
  INV_X1 U16116 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n13361) );
  NAND2_X1 U16117 ( .A1(n12746), .A2(n13361), .ZN(n17058) );
  INV_X1 U16118 ( .A(n12747), .ZN(n12748) );
  NAND2_X1 U16119 ( .A1(n12748), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13357) );
  NAND2_X1 U16120 ( .A1(n10337), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12749) );
  OR2_X1 U16121 ( .A1(n16574), .A2(n12749), .ZN(n13352) );
  INV_X1 U16122 ( .A(n12750), .ZN(n20293) );
  NAND2_X1 U16123 ( .A1(n10337), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12751) );
  OR2_X1 U16124 ( .A1(n20293), .A2(n12751), .ZN(n17131) );
  INV_X1 U16125 ( .A(n20308), .ZN(n12753) );
  AND2_X1 U16126 ( .A1(n10337), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12752) );
  NAND2_X1 U16127 ( .A1(n12753), .A2(n12752), .ZN(n17183) );
  NAND2_X1 U16128 ( .A1(n10337), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12754) );
  OR2_X1 U16129 ( .A1(n16643), .A2(n12754), .ZN(n17167) );
  AND2_X1 U16130 ( .A1(n17183), .A2(n17167), .ZN(n13344) );
  AND2_X1 U16131 ( .A1(n10337), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12755) );
  NAND2_X1 U16132 ( .A1(n16616), .A2(n12755), .ZN(n17144) );
  NAND3_X1 U16133 ( .A1(n16629), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        n10337), .ZN(n17155) );
  AND4_X1 U16134 ( .A1(n17131), .A2(n13344), .A3(n17144), .A4(n17155), .ZN(
        n12758) );
  NAND2_X1 U16135 ( .A1(n10337), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12756) );
  OR2_X1 U16136 ( .A1(n16592), .A2(n12756), .ZN(n13351) );
  NAND2_X1 U16137 ( .A1(n10337), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12757) );
  OR2_X1 U16138 ( .A1(n20278), .A2(n12757), .ZN(n17109) );
  AND4_X1 U16139 ( .A1(n13352), .A2(n12758), .A3(n13351), .A4(n17109), .ZN(
        n12762) );
  AND2_X1 U16140 ( .A1(n10337), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12759) );
  NAND2_X1 U16141 ( .A1(n16548), .A2(n12759), .ZN(n17057) );
  NAND2_X1 U16142 ( .A1(n10337), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12760) );
  INV_X1 U16143 ( .A(n12761), .ZN(n13348) );
  NAND2_X1 U16144 ( .A1(n13348), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17123) );
  AND4_X1 U16145 ( .A1(n12762), .A2(n17057), .A3(n17066), .A4(n17123), .ZN(
        n12765) );
  INV_X1 U16146 ( .A(n12763), .ZN(n12764) );
  NAND2_X1 U16147 ( .A1(n12764), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17076) );
  INV_X1 U16148 ( .A(n12766), .ZN(n12767) );
  NAND2_X1 U16149 ( .A1(n12768), .A2(n12767), .ZN(n12769) );
  NAND2_X1 U16150 ( .A1(n12770), .A2(n12769), .ZN(n16514) );
  OR2_X1 U16151 ( .A1(n16514), .A2(n12627), .ZN(n12771) );
  INV_X1 U16152 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17035) );
  NAND2_X1 U16153 ( .A1(n12771), .A2(n17035), .ZN(n17038) );
  INV_X1 U16154 ( .A(n17018), .ZN(n12773) );
  INV_X1 U16155 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12772) );
  AOI21_X1 U16156 ( .B1(n12773), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n10666), .ZN(n12774) );
  INV_X1 U16157 ( .A(n12774), .ZN(n12775) );
  INV_X1 U16158 ( .A(n12777), .ZN(n12778) );
  XNOR2_X1 U16159 ( .A(n12783), .B(n12778), .ZN(n16431) );
  NAND2_X1 U16160 ( .A1(n16431), .A2(n12946), .ZN(n12791) );
  NAND2_X1 U16161 ( .A1(n12791), .A2(n13197), .ZN(n13202) );
  INV_X1 U16162 ( .A(n12779), .ZN(n12780) );
  NAND2_X1 U16163 ( .A1(n12781), .A2(n12780), .ZN(n12782) );
  NAND2_X1 U16164 ( .A1(n12783), .A2(n12782), .ZN(n16445) );
  INV_X1 U16165 ( .A(n12791), .ZN(n12790) );
  NAND2_X1 U16166 ( .A1(n12946), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12786) );
  OR2_X1 U16167 ( .A1(n12785), .A2(n12786), .ZN(n12789) );
  INV_X1 U16168 ( .A(n12787), .ZN(n16480) );
  AND2_X1 U16169 ( .A1(n12946), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12788) );
  NAND2_X1 U16170 ( .A1(n16480), .A2(n12788), .ZN(n17007) );
  NAND2_X1 U16171 ( .A1(n12789), .A2(n17007), .ZN(n13198) );
  AOI21_X1 U16172 ( .B1(n12790), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n13198), .ZN(n12792) );
  INV_X1 U16173 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13160) );
  OAI21_X1 U16174 ( .B1(n12794), .B2(n12627), .A(n13160), .ZN(n13188) );
  INV_X1 U16175 ( .A(n12794), .ZN(n16430) );
  NAND3_X1 U16176 ( .A1(n16430), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n10337), .ZN(n13237) );
  INV_X1 U16177 ( .A(n12798), .ZN(n12799) );
  NAND2_X1 U16178 ( .A1(n13220), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n12802) );
  NAND2_X1 U16179 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n12801) );
  OAI211_X1 U16180 ( .C1(n12857), .C2(n20334), .A(n12802), .B(n12801), .ZN(
        n12803) );
  AOI21_X1 U16181 ( .B1(n12812), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n12803), .ZN(n14440) );
  INV_X1 U16182 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n22065) );
  NAND2_X1 U16183 ( .A1(n13220), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n12807) );
  NAND2_X1 U16184 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12806) );
  OAI211_X1 U16185 ( .C1(n12857), .C2(n22065), .A(n12807), .B(n12806), .ZN(
        n12808) );
  AOI21_X1 U16186 ( .B1(n12812), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n12808), .ZN(n14337) );
  AOI22_X1 U16187 ( .A1(n13220), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12811) );
  NAND2_X1 U16188 ( .A1(n12809), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n12810) );
  OAI211_X1 U16189 ( .C1(n12890), .C2(n17494), .A(n12811), .B(n12810), .ZN(
        n14499) );
  INV_X1 U16190 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n12815) );
  INV_X1 U16191 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n20990) );
  OR2_X1 U16192 ( .A1(n12879), .A2(n20990), .ZN(n12814) );
  NAND2_X1 U16193 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12813) );
  OAI211_X1 U16194 ( .C1(n12248), .C2(n12815), .A(n12814), .B(n12813), .ZN(
        n12816) );
  AOI21_X1 U16195 ( .B1(n12812), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n12816), .ZN(n14535) );
  INV_X1 U16196 ( .A(n14535), .ZN(n12817) );
  NAND2_X1 U16197 ( .A1(n13220), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n12820) );
  NAND2_X1 U16198 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12819) );
  OAI211_X1 U16199 ( .C1(n12857), .C2(n21858), .A(n12820), .B(n12819), .ZN(
        n12821) );
  AOI21_X1 U16200 ( .B1(n13223), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n12821), .ZN(n14811) );
  AOI22_X1 U16201 ( .A1(n13220), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12823) );
  NAND2_X1 U16202 ( .A1(n12809), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12822) );
  OAI211_X1 U16203 ( .C1(n12890), .C2(n17456), .A(n12823), .B(n12822), .ZN(
        n14822) );
  NAND2_X1 U16204 ( .A1(n12812), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12825) );
  AOI22_X1 U16205 ( .A1(n13220), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n12824) );
  OAI211_X1 U16206 ( .C1(n12248), .C2(n16646), .A(n12825), .B(n12824), .ZN(
        n14884) );
  NAND2_X1 U16207 ( .A1(n13220), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n12827) );
  NAND2_X1 U16208 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12826) );
  OAI211_X1 U16209 ( .C1(n12857), .C2(n12628), .A(n12827), .B(n12826), .ZN(
        n12828) );
  AOI21_X1 U16210 ( .B1(n12812), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n12828), .ZN(n16627) );
  INV_X1 U16211 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n12832) );
  NAND2_X1 U16212 ( .A1(n13220), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n12831) );
  NAND2_X1 U16213 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12830) );
  OAI211_X1 U16214 ( .C1(n12857), .C2(n12832), .A(n12831), .B(n12830), .ZN(
        n12833) );
  AOI21_X1 U16215 ( .B1(n12812), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n12833), .ZN(n16614) );
  AOI22_X1 U16216 ( .A1(n13220), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n12835) );
  NAND2_X1 U16217 ( .A1(n12809), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n12834) );
  OAI211_X1 U16218 ( .C1(n12890), .C2(n17402), .A(n12835), .B(n12834), .ZN(
        n14834) );
  NAND2_X1 U16219 ( .A1(n13220), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n12837) );
  NAND2_X1 U16220 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12836) );
  OAI211_X1 U16221 ( .C1(n12857), .C2(n16606), .A(n12837), .B(n12836), .ZN(
        n12838) );
  AOI21_X1 U16222 ( .B1(n12812), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n12838), .ZN(n14648) );
  NAND2_X1 U16223 ( .A1(n12840), .A2(n12839), .ZN(n14646) );
  INV_X1 U16224 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n22063) );
  INV_X1 U16225 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n21003) );
  OR2_X1 U16226 ( .A1(n12879), .A2(n21003), .ZN(n12842) );
  NAND2_X1 U16227 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12841) );
  OAI211_X1 U16228 ( .C1(n12857), .C2(n22063), .A(n12842), .B(n12841), .ZN(
        n12843) );
  AOI21_X1 U16229 ( .B1(n13223), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n12843), .ZN(n16822) );
  INV_X1 U16230 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n21005) );
  OR2_X1 U16231 ( .A1(n12879), .A2(n21005), .ZN(n12846) );
  NAND2_X1 U16232 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n12845) );
  OAI211_X1 U16233 ( .C1(n12857), .C2(n12847), .A(n12846), .B(n12845), .ZN(
        n12848) );
  AOI21_X1 U16234 ( .B1(n13223), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n12848), .ZN(n16585) );
  AOI22_X1 U16235 ( .A1(n13220), .A2(P2_REIP_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n12850) );
  NAND2_X1 U16236 ( .A1(n12809), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n12849) );
  OAI211_X1 U16237 ( .C1(n12890), .C2(n21906), .A(n12850), .B(n12849), .ZN(
        n16570) );
  NAND2_X1 U16238 ( .A1(n13220), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n12852) );
  NAND2_X1 U16239 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n12851) );
  OAI211_X1 U16240 ( .C1(n12857), .C2(n16557), .A(n12852), .B(n12851), .ZN(
        n12853) );
  AOI21_X1 U16241 ( .B1(n12812), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n12853), .ZN(n16554) );
  INV_X1 U16242 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n21989) );
  INV_X1 U16243 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n21010) );
  OR2_X1 U16244 ( .A1(n12879), .A2(n21010), .ZN(n12856) );
  NAND2_X1 U16245 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n12855) );
  OAI211_X1 U16246 ( .C1(n12857), .C2(n21989), .A(n12856), .B(n12855), .ZN(
        n12858) );
  AOI21_X1 U16247 ( .B1(n12812), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n12858), .ZN(n16802) );
  AOI22_X1 U16248 ( .A1(n13220), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n12860) );
  NAND2_X1 U16249 ( .A1(n12809), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12859) );
  OAI211_X1 U16250 ( .C1(n12890), .C2(n13361), .A(n12860), .B(n12859), .ZN(
        n16537) );
  AOI22_X1 U16251 ( .A1(n13220), .A2(P2_REIP_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n12862) );
  NAND2_X1 U16252 ( .A1(n12809), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n12861) );
  OAI211_X1 U16253 ( .C1(n12890), .C2(n13370), .A(n12862), .B(n12861), .ZN(
        n13373) );
  INV_X1 U16254 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n16515) );
  INV_X1 U16255 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n21015) );
  OR2_X1 U16256 ( .A1(n12879), .A2(n21015), .ZN(n12864) );
  NAND2_X1 U16257 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12863) );
  OAI211_X1 U16258 ( .C1(n12857), .C2(n16515), .A(n12864), .B(n12863), .ZN(
        n12865) );
  AOI21_X1 U16259 ( .B1(n12812), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n12865), .ZN(n16509) );
  INV_X1 U16260 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n21017) );
  OR2_X1 U16261 ( .A1(n12879), .A2(n21017), .ZN(n12867) );
  NAND2_X1 U16262 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n12866) );
  OAI211_X1 U16263 ( .C1(n12857), .C2(n12868), .A(n12867), .B(n12866), .ZN(
        n12869) );
  AOI21_X1 U16264 ( .B1(n13223), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n12869), .ZN(n16499) );
  AOI22_X1 U16265 ( .A1(n13220), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n12871) );
  NAND2_X1 U16266 ( .A1(n12809), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12870) );
  OAI211_X1 U16267 ( .C1(n12890), .C2(n10338), .A(n12871), .B(n12870), .ZN(
        n16482) );
  INV_X1 U16268 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n21021) );
  OR2_X1 U16269 ( .A1(n12879), .A2(n21021), .ZN(n12873) );
  NAND2_X1 U16270 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n12872) );
  OAI211_X1 U16271 ( .C1(n12857), .C2(n10511), .A(n12873), .B(n12872), .ZN(
        n12874) );
  AOI21_X1 U16272 ( .B1(n12812), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n12874), .ZN(n16467) );
  INV_X1 U16273 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n21023) );
  OR2_X1 U16274 ( .A1(n12879), .A2(n21023), .ZN(n12876) );
  NAND2_X1 U16275 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12875) );
  OAI211_X1 U16276 ( .C1(n12857), .C2(n16767), .A(n12876), .B(n12875), .ZN(
        n12877) );
  AOI21_X1 U16277 ( .B1(n12812), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n12877), .ZN(n16455) );
  INV_X1 U16278 ( .A(n16455), .ZN(n12878) );
  INV_X1 U16279 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n12882) );
  INV_X1 U16280 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n21967) );
  OR2_X1 U16281 ( .A1(n12879), .A2(n21967), .ZN(n12881) );
  NAND2_X1 U16282 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12880) );
  OAI211_X1 U16283 ( .C1(n12857), .C2(n12882), .A(n12881), .B(n12880), .ZN(
        n12883) );
  AOI21_X1 U16284 ( .B1(n12812), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n12883), .ZN(n16442) );
  AOI22_X1 U16285 ( .A1(n13220), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n12885) );
  NAND2_X1 U16286 ( .A1(n12809), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n12884) );
  OAI211_X1 U16287 ( .C1(n12890), .C2(n13197), .A(n12885), .B(n12884), .ZN(
        n13207) );
  NAND2_X1 U16288 ( .A1(n12812), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12887) );
  AOI22_X1 U16289 ( .A1(n13220), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n12886) );
  OAI211_X1 U16290 ( .C1(n22023), .C2(n12857), .A(n12887), .B(n12886), .ZN(
        n13178) );
  INV_X1 U16291 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13401) );
  AOI22_X1 U16292 ( .A1(n13220), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n12889) );
  NAND2_X1 U16293 ( .A1(n12809), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12888) );
  OAI211_X1 U16294 ( .C1(n12890), .C2(n13401), .A(n12889), .B(n12888), .ZN(
        n13218) );
  NAND2_X1 U16295 ( .A1(n14713), .A2(n15209), .ZN(n12891) );
  NAND2_X1 U16296 ( .A1(n12891), .A2(n12223), .ZN(n12892) );
  NAND2_X1 U16297 ( .A1(n12920), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n12897) );
  INV_X1 U16298 ( .A(n12908), .ZN(n12899) );
  INV_X1 U16299 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n12894) );
  NAND2_X1 U16300 ( .A1(n20834), .A2(n12894), .ZN(n12895) );
  NAND3_X1 U16301 ( .A1(n12551), .A2(n9987), .A3(n20834), .ZN(n12942) );
  AND2_X1 U16302 ( .A1(n21083), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n21080) );
  INV_X1 U16303 ( .A(n21080), .ZN(n20839) );
  NAND2_X1 U16304 ( .A1(n12899), .A2(n20839), .ZN(n12903) );
  INV_X1 U16305 ( .A(n14426), .ZN(n12902) );
  NAND2_X1 U16306 ( .A1(n12901), .A2(n20834), .ZN(n12927) );
  NAND2_X1 U16307 ( .A1(n12902), .A2(n12919), .ZN(n12916) );
  NAND2_X1 U16308 ( .A1(n14418), .A2(n14419), .ZN(n12914) );
  NOR2_X1 U16309 ( .A1(n12905), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12918) );
  AOI22_X1 U16310 ( .A1(n12918), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n12919), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12907) );
  NAND2_X1 U16311 ( .A1(n12920), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n12906) );
  NAND2_X1 U16312 ( .A1(n12907), .A2(n12906), .ZN(n12912) );
  XNOR2_X1 U16313 ( .A(n12914), .B(n12912), .ZN(n14083) );
  AOI22_X1 U16314 ( .A1(n14426), .A2(n12908), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12911) );
  INV_X2 U16315 ( .A(n12942), .ZN(n13090) );
  NAND2_X1 U16316 ( .A1(n13090), .A2(n12909), .ZN(n12910) );
  AND2_X1 U16317 ( .A1(n12911), .A2(n12910), .ZN(n14082) );
  NAND2_X1 U16318 ( .A1(n14083), .A2(n14082), .ZN(n14085) );
  INV_X1 U16319 ( .A(n12912), .ZN(n12913) );
  NAND2_X1 U16320 ( .A1(n12914), .A2(n12913), .ZN(n12915) );
  NAND2_X1 U16321 ( .A1(n14085), .A2(n12915), .ZN(n12925) );
  NAND2_X1 U16322 ( .A1(n13090), .A2(n12591), .ZN(n12917) );
  OAI211_X1 U16323 ( .C1(n20834), .C2(n21065), .A(n12917), .B(n12916), .ZN(
        n12923) );
  XNOR2_X1 U16324 ( .A(n12925), .B(n12923), .ZN(n13974) );
  AOI22_X1 U16325 ( .A1(n13127), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n13126), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12922) );
  NAND2_X1 U16326 ( .A1(n13114), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n12921) );
  AND2_X1 U16327 ( .A1(n12922), .A2(n12921), .ZN(n13973) );
  INV_X1 U16328 ( .A(n12923), .ZN(n12924) );
  NAND2_X1 U16329 ( .A1(n12925), .A2(n12924), .ZN(n12926) );
  NAND2_X1 U16330 ( .A1(n13976), .A2(n12926), .ZN(n16690) );
  INV_X1 U16331 ( .A(n16690), .ZN(n12933) );
  INV_X2 U16332 ( .A(n13106), .ZN(n13114) );
  INV_X1 U16333 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n17526) );
  OAI22_X1 U16334 ( .A1(n12927), .A2(n17526), .B1(n21054), .B2(n20834), .ZN(
        n12928) );
  AOI21_X1 U16335 ( .B1(P2_REIP_REG_3__SCAN_IN), .B2(n13114), .A(n12928), .ZN(
        n12931) );
  AOI22_X1 U16336 ( .A1(n13090), .A2(n12929), .B1(n13127), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n12930) );
  NAND2_X1 U16337 ( .A1(n12933), .A2(n12932), .ZN(n16688) );
  AOI22_X1 U16338 ( .A1(n13127), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n13126), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12937) );
  NAND2_X1 U16339 ( .A1(n13114), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n12936) );
  NAND2_X1 U16340 ( .A1(n13090), .A2(n12934), .ZN(n12935) );
  AOI22_X1 U16341 ( .A1(n13127), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n13126), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12941) );
  NAND2_X1 U16342 ( .A1(n13114), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n12940) );
  NAND2_X1 U16343 ( .A1(n13090), .A2(n12938), .ZN(n12939) );
  AOI22_X1 U16344 ( .A1(n13127), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n13126), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12945) );
  NAND2_X1 U16345 ( .A1(n13114), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n12944) );
  NAND2_X1 U16346 ( .A1(n12945), .A2(n12944), .ZN(n14624) );
  NAND2_X1 U16347 ( .A1(n13090), .A2(n12946), .ZN(n12947) );
  NAND2_X1 U16348 ( .A1(n12948), .A2(n12947), .ZN(n14635) );
  AOI22_X1 U16349 ( .A1(n13127), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n13126), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n12950) );
  NAND2_X1 U16350 ( .A1(n13114), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n12949) );
  NAND2_X1 U16351 ( .A1(n12950), .A2(n12949), .ZN(n14634) );
  NAND2_X1 U16352 ( .A1(n14635), .A2(n14634), .ZN(n14626) );
  INV_X1 U16353 ( .A(n14626), .ZN(n12968) );
  AOI22_X1 U16354 ( .A1(n13127), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n13126), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12966) );
  NAND2_X1 U16355 ( .A1(n13114), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n12965) );
  AOI22_X1 U16356 ( .A1(n12362), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12379), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12957) );
  AOI22_X1 U16357 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n15148), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12956) );
  INV_X1 U16358 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17566) );
  NAND2_X1 U16359 ( .A1(n15171), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12952) );
  NAND2_X1 U16360 ( .A1(n15172), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12951) );
  OAI211_X1 U16361 ( .C1(n13078), .C2(n17566), .A(n12952), .B(n12951), .ZN(
        n12953) );
  INV_X1 U16362 ( .A(n12953), .ZN(n12955) );
  AOI22_X1 U16363 ( .A1(n15177), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n15176), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12954) );
  NAND4_X1 U16364 ( .A1(n12957), .A2(n12956), .A3(n12955), .A4(n12954), .ZN(
        n12963) );
  AOI22_X1 U16365 ( .A1(n12524), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12341), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12961) );
  AOI22_X1 U16366 ( .A1(n15125), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12412), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12960) );
  AOI22_X1 U16367 ( .A1(n12371), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12350), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12959) );
  NAND2_X1 U16368 ( .A1(n12525), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12958) );
  NAND4_X1 U16369 ( .A1(n12961), .A2(n12960), .A3(n12959), .A4(n12958), .ZN(
        n12962) );
  NAND2_X1 U16370 ( .A1(n13090), .A2(n14815), .ZN(n12964) );
  NAND2_X1 U16371 ( .A1(n12968), .A2(n12967), .ZN(n14625) );
  AOI22_X1 U16372 ( .A1(n13127), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n13126), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12986) );
  NAND2_X1 U16373 ( .A1(n13114), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n12985) );
  AOI22_X1 U16374 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n12362), .B1(
        n12379), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12977) );
  AOI22_X1 U16375 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n15148), .B1(
        n12451), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12976) );
  OAI22_X1 U16376 ( .A1(n12970), .A2(n15145), .B1(n15143), .B2(n12969), .ZN(
        n12974) );
  NAND2_X1 U16377 ( .A1(n15171), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n12972) );
  NAND2_X1 U16378 ( .A1(n15172), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n12971) );
  OAI211_X1 U16379 ( .C1(n13078), .C2(n17573), .A(n12972), .B(n12971), .ZN(
        n12973) );
  NOR2_X1 U16380 ( .A1(n12974), .A2(n12973), .ZN(n12975) );
  NAND3_X1 U16381 ( .A1(n12977), .A2(n12976), .A3(n12975), .ZN(n12983) );
  AOI22_X1 U16382 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n12341), .B1(
        n12524), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12981) );
  AOI22_X1 U16383 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n12412), .B1(
        n15125), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12980) );
  AOI22_X1 U16384 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12371), .B1(
        n12350), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12979) );
  NAND2_X1 U16385 ( .A1(n12525), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12978) );
  NAND4_X1 U16386 ( .A1(n12981), .A2(n12980), .A3(n12979), .A4(n12978), .ZN(
        n12982) );
  NAND2_X1 U16387 ( .A1(n13090), .A2(n14820), .ZN(n12984) );
  AOI22_X1 U16388 ( .A1(n13127), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n13126), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n13005) );
  NAND2_X1 U16389 ( .A1(n13114), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n13004) );
  AOI22_X1 U16390 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12379), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12996) );
  NAND2_X1 U16391 ( .A1(n15172), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n12990) );
  NAND2_X1 U16392 ( .A1(n12350), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n12989) );
  OAI211_X1 U16393 ( .C1(n13078), .C2(n12991), .A(n12990), .B(n12989), .ZN(
        n12992) );
  INV_X1 U16394 ( .A(n12992), .ZN(n12995) );
  AOI22_X1 U16395 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n15177), .B1(
        n15176), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12994) );
  AOI22_X1 U16396 ( .A1(n12362), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n15125), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12993) );
  NAND4_X1 U16397 ( .A1(n12996), .A2(n12995), .A3(n12994), .A4(n12993), .ZN(
        n13002) );
  AOI22_X1 U16398 ( .A1(n12524), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12341), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13000) );
  AOI22_X1 U16399 ( .A1(n15148), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12412), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12999) );
  AOI22_X1 U16400 ( .A1(n12371), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n15171), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12998) );
  NAND2_X1 U16401 ( .A1(n12525), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n12997) );
  NAND4_X1 U16402 ( .A1(n13000), .A2(n12999), .A3(n12998), .A4(n12997), .ZN(
        n13001) );
  NAND2_X1 U16403 ( .A1(n13090), .A2(n14887), .ZN(n13003) );
  INV_X1 U16404 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n17159) );
  AOI22_X1 U16405 ( .A1(n13127), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n13126), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n13022) );
  AOI22_X1 U16406 ( .A1(n12362), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12379), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13014) );
  AOI22_X1 U16407 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n15148), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13013) );
  OAI22_X1 U16408 ( .A1(n15145), .A2(n13007), .B1(n15143), .B2(n13006), .ZN(
        n13011) );
  NAND2_X1 U16409 ( .A1(n15171), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n13009) );
  NAND2_X1 U16410 ( .A1(n15172), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n13008) );
  OAI211_X1 U16411 ( .C1(n13078), .C2(n12301), .A(n13009), .B(n13008), .ZN(
        n13010) );
  NOR2_X1 U16412 ( .A1(n13011), .A2(n13010), .ZN(n13012) );
  NAND3_X1 U16413 ( .A1(n13014), .A2(n13013), .A3(n13012), .ZN(n13020) );
  AOI22_X1 U16414 ( .A1(n12524), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12341), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13018) );
  AOI22_X1 U16415 ( .A1(n15125), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12412), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13017) );
  AOI22_X1 U16416 ( .A1(n12371), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12350), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13016) );
  NAND2_X1 U16417 ( .A1(n12525), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n13015) );
  NAND4_X1 U16418 ( .A1(n13018), .A2(n13017), .A3(n13016), .A4(n13015), .ZN(
        n13019) );
  NAND2_X1 U16419 ( .A1(n13090), .A2(n16837), .ZN(n13021) );
  OAI211_X1 U16420 ( .C1(n13106), .C2(n17159), .A(n13022), .B(n13021), .ZN(
        n14642) );
  AOI22_X1 U16421 ( .A1(n13127), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n13126), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n13038) );
  NAND2_X1 U16422 ( .A1(n13114), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n13037) );
  AOI22_X1 U16423 ( .A1(n12362), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12451), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13029) );
  NAND2_X1 U16424 ( .A1(n15172), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n13024) );
  NAND2_X1 U16425 ( .A1(n12350), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n13023) );
  OAI211_X1 U16426 ( .C1(n13078), .C2(n20442), .A(n13024), .B(n13023), .ZN(
        n13025) );
  INV_X1 U16427 ( .A(n13025), .ZN(n13028) );
  AOI22_X1 U16428 ( .A1(n15177), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n15176), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13027) );
  AOI22_X1 U16429 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n15125), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13026) );
  NAND4_X1 U16430 ( .A1(n13029), .A2(n13028), .A3(n13027), .A4(n13026), .ZN(
        n13035) );
  AOI22_X1 U16431 ( .A1(n12524), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12341), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13033) );
  AOI22_X1 U16432 ( .A1(n15148), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12412), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13032) );
  AOI22_X1 U16433 ( .A1(n12371), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n15171), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13031) );
  NAND2_X1 U16434 ( .A1(n12525), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n13030) );
  NAND4_X1 U16435 ( .A1(n13033), .A2(n13032), .A3(n13031), .A4(n13030), .ZN(
        n13034) );
  OR2_X1 U16436 ( .A1(n13035), .A2(n13034), .ZN(n16831) );
  NAND2_X1 U16437 ( .A1(n13090), .A2(n16831), .ZN(n13036) );
  AOI22_X1 U16438 ( .A1(n13127), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n13126), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n13056) );
  NAND2_X1 U16439 ( .A1(n13114), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n13055) );
  AOI22_X1 U16440 ( .A1(n12362), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12379), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13047) );
  AOI22_X1 U16441 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15148), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13046) );
  OAI22_X1 U16442 ( .A1(n15145), .A2(n13040), .B1(n15143), .B2(n13039), .ZN(
        n13044) );
  NAND2_X1 U16443 ( .A1(n15171), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n13042) );
  NAND2_X1 U16444 ( .A1(n15172), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n13041) );
  OAI211_X1 U16445 ( .C1(n13078), .C2(n14494), .A(n13042), .B(n13041), .ZN(
        n13043) );
  NOR2_X1 U16446 ( .A1(n13044), .A2(n13043), .ZN(n13045) );
  NAND3_X1 U16447 ( .A1(n13047), .A2(n13046), .A3(n13045), .ZN(n13053) );
  AOI22_X1 U16448 ( .A1(n12524), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12341), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13051) );
  AOI22_X1 U16449 ( .A1(n15125), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12412), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13050) );
  AOI22_X1 U16450 ( .A1(n12371), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12350), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13049) );
  NAND2_X1 U16451 ( .A1(n12525), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n13048) );
  NAND4_X1 U16452 ( .A1(n13051), .A2(n13050), .A3(n13049), .A4(n13048), .ZN(
        n13052) );
  NAND2_X1 U16453 ( .A1(n13090), .A2(n15056), .ZN(n13054) );
  AND2_X2 U16454 ( .A1(n14617), .A2(n13057), .ZN(n14619) );
  INV_X1 U16455 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n17125) );
  AOI22_X1 U16456 ( .A1(n13127), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n13126), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n13074) );
  AOI22_X1 U16457 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n15148), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13066) );
  OAI22_X1 U16458 ( .A1(n15145), .A2(n13058), .B1(n13078), .B2(n20449), .ZN(
        n13063) );
  NAND2_X1 U16459 ( .A1(n15172), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n13060) );
  NAND2_X1 U16460 ( .A1(n12350), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n13059) );
  OAI211_X1 U16461 ( .C1(n15143), .C2(n13061), .A(n13060), .B(n13059), .ZN(
        n13062) );
  NOR2_X1 U16462 ( .A1(n13063), .A2(n13062), .ZN(n13065) );
  AOI22_X1 U16463 ( .A1(n12362), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12412), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13064) );
  NAND3_X1 U16464 ( .A1(n13066), .A2(n13065), .A3(n13064), .ZN(n13072) );
  AOI22_X1 U16465 ( .A1(n12524), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12341), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13070) );
  AOI22_X1 U16466 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n15125), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13069) );
  AOI22_X1 U16467 ( .A1(n12371), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n15171), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13068) );
  NAND2_X1 U16468 ( .A1(n12525), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n13067) );
  NAND4_X1 U16469 ( .A1(n13070), .A2(n13069), .A3(n13068), .A4(n13067), .ZN(
        n13071) );
  NAND2_X1 U16470 ( .A1(n13090), .A2(n15057), .ZN(n13073) );
  OAI211_X1 U16471 ( .C1(n13106), .C2(n17125), .A(n13074), .B(n13073), .ZN(
        n14807) );
  AOI22_X1 U16472 ( .A1(n13127), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n13126), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n13092) );
  AOI22_X1 U16473 ( .A1(n12362), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12379), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13083) );
  AOI22_X1 U16474 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n15148), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13082) );
  INV_X1 U16475 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15180) );
  INV_X1 U16476 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13075) );
  OAI22_X1 U16477 ( .A1(n15145), .A2(n15180), .B1(n15143), .B2(n13075), .ZN(
        n13080) );
  INV_X1 U16478 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n20458) );
  NAND2_X1 U16479 ( .A1(n15171), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n13077) );
  NAND2_X1 U16480 ( .A1(n15172), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n13076) );
  OAI211_X1 U16481 ( .C1(n13078), .C2(n20458), .A(n13077), .B(n13076), .ZN(
        n13079) );
  NOR2_X1 U16482 ( .A1(n13080), .A2(n13079), .ZN(n13081) );
  NAND3_X1 U16483 ( .A1(n13083), .A2(n13082), .A3(n13081), .ZN(n13089) );
  AOI22_X1 U16484 ( .A1(n12524), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12341), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13087) );
  AOI22_X1 U16485 ( .A1(n15125), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12412), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13086) );
  AOI22_X1 U16486 ( .A1(n12371), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12350), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13085) );
  NAND2_X1 U16487 ( .A1(n12525), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n13084) );
  NAND4_X1 U16488 ( .A1(n13087), .A2(n13086), .A3(n13085), .A4(n13084), .ZN(
        n13088) );
  OR2_X1 U16489 ( .A1(n13089), .A2(n13088), .ZN(n16815) );
  NAND2_X1 U16490 ( .A1(n13090), .A2(n16815), .ZN(n13091) );
  OAI211_X1 U16491 ( .C1(n13106), .C2(n21003), .A(n13092), .B(n13091), .ZN(
        n16953) );
  AOI22_X1 U16492 ( .A1(n13127), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n13126), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n13094) );
  NAND2_X1 U16493 ( .A1(n13114), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n13093) );
  AOI22_X1 U16494 ( .A1(n13127), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n13126), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n13096) );
  NAND2_X1 U16495 ( .A1(n13114), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n13095) );
  AOI22_X1 U16496 ( .A1(n13127), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n13126), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n13098) );
  NAND2_X1 U16497 ( .A1(n13114), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n13097) );
  NAND2_X1 U16498 ( .A1(n13098), .A2(n13097), .ZN(n16566) );
  NAND2_X1 U16499 ( .A1(n16573), .A2(n16566), .ZN(n16565) );
  AOI22_X1 U16500 ( .A1(n13127), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n13126), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n13100) );
  NAND2_X1 U16501 ( .A1(n13114), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n13099) );
  NOR2_X4 U16502 ( .A1(n16565), .A2(n16927), .ZN(n16532) );
  AOI22_X1 U16503 ( .A1(n13127), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n13126), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n13102) );
  NAND2_X1 U16504 ( .A1(n13114), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n13101) );
  AOI22_X1 U16505 ( .A1(n13127), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n13126), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n13105) );
  NAND2_X1 U16506 ( .A1(n13114), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n13104) );
  AOI22_X1 U16507 ( .A1(n13127), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n13126), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n13108) );
  NAND2_X1 U16508 ( .A1(n13114), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n13107) );
  NAND2_X1 U16509 ( .A1(n13108), .A2(n13107), .ZN(n16512) );
  AOI22_X1 U16510 ( .A1(n13127), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n13126), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n13110) );
  NAND2_X1 U16511 ( .A1(n12920), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n13109) );
  AOI22_X1 U16512 ( .A1(n13127), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n13126), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n13112) );
  NAND2_X1 U16513 ( .A1(n13114), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n13111) );
  INV_X1 U16514 ( .A(n16484), .ZN(n13113) );
  NAND2_X1 U16515 ( .A1(n16483), .A2(n13113), .ZN(n16474) );
  AOI22_X1 U16516 ( .A1(n13127), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n13126), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n13116) );
  NAND2_X1 U16517 ( .A1(n13114), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n13115) );
  NAND2_X1 U16518 ( .A1(n13116), .A2(n13115), .ZN(n16476) );
  INV_X1 U16519 ( .A(n16476), .ZN(n13117) );
  NOR2_X2 U16520 ( .A1(n16474), .A2(n13117), .ZN(n16451) );
  AOI22_X1 U16521 ( .A1(n13127), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n13126), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13119) );
  NAND2_X1 U16522 ( .A1(n13114), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n13118) );
  NAND2_X1 U16523 ( .A1(n13119), .A2(n13118), .ZN(n16452) );
  AOI22_X1 U16524 ( .A1(n13127), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n13126), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13121) );
  NAND2_X1 U16525 ( .A1(n12920), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n13120) );
  AOI22_X1 U16526 ( .A1(n13127), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n13126), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n13123) );
  NAND2_X1 U16527 ( .A1(n12920), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n13122) );
  AOI22_X1 U16528 ( .A1(n13127), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n13126), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13125) );
  NAND2_X1 U16529 ( .A1(n12920), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n13124) );
  NAND2_X1 U16530 ( .A1(n13125), .A2(n13124), .ZN(n13180) );
  INV_X1 U16531 ( .A(n13132), .ZN(n13131) );
  AOI22_X1 U16532 ( .A1(n13127), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n13126), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13129) );
  NAND2_X1 U16533 ( .A1(n12920), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n13128) );
  AND2_X1 U16534 ( .A1(n13129), .A2(n13128), .ZN(n13133) );
  INV_X1 U16535 ( .A(n13133), .ZN(n13130) );
  NAND2_X1 U16536 ( .A1(n13131), .A2(n13130), .ZN(n13397) );
  NAND2_X1 U16537 ( .A1(n13132), .A2(n13133), .ZN(n13134) );
  NAND2_X2 U16538 ( .A1(n13397), .A2(n13134), .ZN(n15343) );
  NAND2_X1 U16539 ( .A1(n9755), .A2(n13135), .ZN(n14730) );
  NAND2_X1 U16540 ( .A1(n14736), .A2(n13145), .ZN(n13137) );
  NAND2_X1 U16541 ( .A1(n14730), .A2(n13137), .ZN(n13138) );
  NAND2_X1 U16542 ( .A1(n21042), .A2(n16421), .ZN(n13139) );
  NAND2_X1 U16543 ( .A1(n20343), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n15354) );
  NAND2_X1 U16544 ( .A1(n15209), .A2(n20433), .ZN(n13140) );
  NOR2_X1 U16545 ( .A1(n13140), .A2(n12631), .ZN(n13141) );
  AND2_X1 U16546 ( .A1(n13135), .A2(n13141), .ZN(n14727) );
  NAND2_X1 U16547 ( .A1(n13164), .A2(n14727), .ZN(n17361) );
  NAND2_X1 U16548 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14091) );
  INV_X1 U16549 ( .A(n14091), .ZN(n13986) );
  NAND2_X1 U16550 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13986), .ZN(
        n13157) );
  NAND2_X1 U16551 ( .A1(n21972), .A2(n14091), .ZN(n13163) );
  INV_X1 U16552 ( .A(n13163), .ZN(n13156) );
  NAND2_X1 U16553 ( .A1(n13143), .A2(n13142), .ZN(n13154) );
  MUX2_X1 U16554 ( .A(n13144), .B(n20433), .S(n14870), .Z(n13151) );
  NAND2_X1 U16555 ( .A1(n13146), .A2(n13145), .ZN(n14706) );
  NAND2_X1 U16556 ( .A1(n14706), .A2(n13147), .ZN(n13149) );
  NAND2_X1 U16557 ( .A1(n13149), .A2(n13148), .ZN(n13150) );
  NAND2_X1 U16558 ( .A1(n13151), .A2(n13150), .ZN(n13152) );
  AOI21_X1 U16559 ( .B1(n13154), .B2(n13153), .A(n13152), .ZN(n14711) );
  NAND2_X1 U16560 ( .A1(n14711), .A2(n9759), .ZN(n13155) );
  NAND2_X1 U16561 ( .A1(n13164), .A2(n13155), .ZN(n13984) );
  NOR2_X1 U16562 ( .A1(n22037), .A2(n12506), .ZN(n17508) );
  INV_X1 U16563 ( .A(n17508), .ZN(n13158) );
  NAND2_X1 U16564 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13162), .ZN(
        n17481) );
  NAND2_X1 U16565 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n13168) );
  NOR2_X1 U16566 ( .A1(n13368), .A2(n13370), .ZN(n13362) );
  NAND2_X1 U16567 ( .A1(n13161), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17278) );
  NAND2_X1 U16568 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13172) );
  NAND2_X1 U16569 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13182) );
  NOR2_X1 U16570 ( .A1(n13182), .A2(n13160), .ZN(n13174) );
  INV_X1 U16571 ( .A(n13174), .ZN(n13400) );
  NOR2_X1 U16572 ( .A1(n13402), .A2(n13400), .ZN(n13175) );
  NAND2_X1 U16573 ( .A1(n13162), .A2(n17494), .ZN(n17492) );
  OR2_X1 U16574 ( .A1(n17361), .A2(n13163), .ZN(n13980) );
  OAI211_X1 U16575 ( .C1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .C2(n13984), .A(
        n13980), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13166) );
  INV_X1 U16576 ( .A(n13164), .ZN(n13165) );
  INV_X1 U16577 ( .A(n20343), .ZN(n20260) );
  NAND2_X1 U16578 ( .A1(n13165), .A2(n20260), .ZN(n18115) );
  OAI21_X1 U16579 ( .B1(n13984), .B2(n13986), .A(n18115), .ZN(n13985) );
  NOR2_X1 U16580 ( .A1(n13166), .A2(n13985), .ZN(n17525) );
  NAND2_X1 U16581 ( .A1(n17525), .A2(n17508), .ZN(n13167) );
  NAND2_X1 U16582 ( .A1(n18129), .A2(n18115), .ZN(n17502) );
  NAND2_X1 U16583 ( .A1(n13167), .A2(n17502), .ZN(n17493) );
  NAND2_X1 U16584 ( .A1(n10205), .A2(n13168), .ZN(n13169) );
  NAND2_X1 U16585 ( .A1(n17453), .A2(n13170), .ZN(n17290) );
  NAND2_X1 U16586 ( .A1(n17290), .A2(n17502), .ZN(n13171) );
  NAND2_X1 U16587 ( .A1(n17291), .A2(n13171), .ZN(n17282) );
  INV_X1 U16588 ( .A(n13172), .ZN(n17265) );
  NOR2_X1 U16589 ( .A1(n18129), .A2(n17265), .ZN(n13173) );
  NOR2_X1 U16590 ( .A1(n17282), .A2(n13173), .ZN(n17257) );
  OAI211_X1 U16591 ( .C1(n18129), .C2(n13174), .A(n17257), .B(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13405) );
  OAI21_X1 U16592 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n13175), .A(
        n13405), .ZN(n13176) );
  NOR2_X1 U16593 ( .A1(n13177), .A2(n13178), .ZN(n13179) );
  OR2_X1 U16594 ( .A1(n9837), .A2(n13180), .ZN(n13181) );
  INV_X1 U16595 ( .A(n13402), .ZN(n13184) );
  NOR2_X1 U16596 ( .A1(n13182), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13183) );
  INV_X1 U16597 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n21028) );
  NOR2_X1 U16598 ( .A1(n13139), .A2(n21028), .ZN(n16974) );
  AOI21_X1 U16599 ( .B1(n13184), .B2(n13183), .A(n16974), .ZN(n13187) );
  INV_X1 U16600 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17256) );
  NAND2_X1 U16601 ( .A1(n13184), .A2(n17256), .ZN(n17255) );
  NAND2_X1 U16602 ( .A1(n17257), .A2(n17255), .ZN(n13209) );
  NAND2_X1 U16603 ( .A1(n13197), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13185) );
  NOR2_X1 U16604 ( .A1(n13402), .A2(n13185), .ZN(n13208) );
  OAI21_X1 U16605 ( .B1(n13209), .B2(n13208), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13186) );
  OAI211_X1 U16606 ( .C1(n16853), .C2(n18123), .A(n13187), .B(n13186), .ZN(
        n13192) );
  NAND2_X1 U16607 ( .A1(n13237), .A2(n13188), .ZN(n13189) );
  XNOR2_X1 U16608 ( .A(n13190), .B(n13189), .ZN(n16971) );
  NAND2_X1 U16609 ( .A1(n13194), .A2(n18126), .ZN(n13195) );
  NAND3_X1 U16610 ( .A1(n10658), .A2(n13196), .A3(n13195), .ZN(P2_U3017) );
  XNOR2_X1 U16611 ( .A(n13199), .B(n13201), .ZN(n16989) );
  INV_X1 U16612 ( .A(n13199), .ZN(n13200) );
  NAND2_X1 U16613 ( .A1(n13203), .A2(n13202), .ZN(n13204) );
  INV_X1 U16614 ( .A(n13177), .ZN(n13206) );
  INV_X1 U16615 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n21026) );
  NOR2_X1 U16616 ( .A1(n13139), .A2(n21026), .ZN(n16982) );
  AOI211_X1 U16617 ( .C1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n13209), .A(
        n16982), .B(n13208), .ZN(n13212) );
  XOR2_X1 U16618 ( .A(n13210), .B(n16439), .Z(n16859) );
  NAND2_X1 U16619 ( .A1(n16859), .A2(n17505), .ZN(n13211) );
  OAI211_X1 U16620 ( .C1(n16984), .C2(n17518), .A(n13212), .B(n13211), .ZN(
        n13213) );
  INV_X1 U16621 ( .A(n13213), .ZN(n13214) );
  XNOR2_X1 U16622 ( .A(n13216), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13413) );
  AND2_X1 U16623 ( .A1(n21088), .A2(n20237), .ZN(n13225) );
  INV_X1 U16624 ( .A(n13225), .ZN(n13217) );
  INV_X1 U16625 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n13332) );
  AOI22_X1 U16626 ( .A1(n13220), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n13221) );
  OAI21_X1 U16627 ( .B1(n12857), .B2(n13332), .A(n13221), .ZN(n13222) );
  AOI21_X1 U16628 ( .B1(n13223), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n13222), .ZN(n13224) );
  NAND2_X1 U16629 ( .A1(n21089), .A2(n21087), .ZN(n13226) );
  NAND2_X1 U16630 ( .A1(n13226), .A2(n13225), .ZN(n20239) );
  NOR2_X1 U16631 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17545) );
  OR2_X1 U16632 ( .A1(n21042), .A2(n17545), .ZN(n21055) );
  NAND2_X1 U16633 ( .A1(n21055), .A2(n17596), .ZN(n13227) );
  AND2_X1 U16634 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n13457) );
  AND2_X1 U16635 ( .A1(n20712), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13256) );
  INV_X1 U16636 ( .A(n13256), .ZN(n13228) );
  NAND2_X1 U16637 ( .A1(n17596), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n14856) );
  NAND2_X1 U16638 ( .A1(n13228), .A2(n14856), .ZN(n13588) );
  NAND2_X1 U16639 ( .A1(n13260), .A2(n13230), .ZN(n13267) );
  NOR2_X2 U16640 ( .A1(n13271), .A2(n17172), .ZN(n13274) );
  AND2_X2 U16641 ( .A1(n13273), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13277) );
  INV_X1 U16642 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n13279) );
  NOR2_X2 U16643 ( .A1(n13284), .A2(n13232), .ZN(n13257) );
  NAND2_X1 U16644 ( .A1(n13257), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13290) );
  INV_X1 U16645 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17071) );
  INV_X1 U16646 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17049) );
  INV_X1 U16647 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n13297) );
  INV_X1 U16648 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17030) );
  NAND2_X1 U16649 ( .A1(n13300), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13303) );
  INV_X1 U16650 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17012) );
  OR2_X2 U16651 ( .A1(n13303), .A2(n17012), .ZN(n13310) );
  INV_X1 U16652 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n13309) );
  NOR2_X2 U16653 ( .A1(n13310), .A2(n13309), .ZN(n13308) );
  AND2_X2 U16654 ( .A1(n13308), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13312) );
  INV_X1 U16655 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16972) );
  INV_X1 U16656 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n13336) );
  INV_X1 U16657 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13233) );
  INV_X1 U16658 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n13395) );
  NOR2_X1 U16659 ( .A1(n13139), .A2(n13395), .ZN(n13404) );
  AOI21_X1 U16660 ( .B1(n17214), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n13404), .ZN(n13234) );
  INV_X1 U16661 ( .A(n13234), .ZN(n13235) );
  OAI21_X1 U16662 ( .B1(n15359), .B2(n17242), .A(n13236), .ZN(n13247) );
  INV_X1 U16663 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n15347) );
  NAND2_X1 U16664 ( .A1(n13241), .A2(n15347), .ZN(n13243) );
  MUX2_X1 U16665 ( .A(n13243), .B(n13242), .S(n9987), .Z(n15362) );
  NOR2_X1 U16666 ( .A1(n15362), .A2(n12627), .ZN(n13244) );
  XNOR2_X1 U16667 ( .A(n13244), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13245) );
  XNOR2_X1 U16668 ( .A(n13246), .B(n13245), .ZN(n13409) );
  OAI21_X1 U16669 ( .B1(n13413), .B2(n17218), .A(n13248), .ZN(P2_U2983) );
  INV_X1 U16670 ( .A(n15352), .ZN(n13251) );
  INV_X1 U16671 ( .A(n13461), .ZN(n13249) );
  NOR2_X1 U16672 ( .A1(n20959), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n13326) );
  NAND2_X1 U16673 ( .A1(n12207), .A2(n13326), .ZN(n13250) );
  NAND2_X1 U16674 ( .A1(n13251), .A2(n20329), .ZN(n13343) );
  NOR2_X1 U16675 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13255) );
  NAND2_X1 U16676 ( .A1(n13256), .A2(n13255), .ZN(n20351) );
  INV_X1 U16677 ( .A(n13257), .ZN(n13288) );
  INV_X1 U16678 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n13258) );
  NAND2_X1 U16679 ( .A1(n13288), .A2(n13258), .ZN(n13259) );
  NAND2_X1 U16680 ( .A1(n13290), .A2(n13259), .ZN(n17084) );
  XNOR2_X1 U16681 ( .A(n13260), .B(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17212) );
  AOI21_X1 U16682 ( .B1(n18113), .B2(n13263), .A(n13260), .ZN(n18101) );
  AOI21_X1 U16683 ( .B1(n20340), .B2(n13262), .A(n13264), .ZN(n20354) );
  INV_X1 U16684 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16741) );
  MUX2_X1 U16685 ( .A(n14087), .B(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .S(n17596), .Z(n16719) );
  NAND2_X1 U16686 ( .A1(n16739), .A2(n16719), .ZN(n16722) );
  AOI21_X1 U16687 ( .B1(n21861), .B2(n13229), .A(n13261), .ZN(n16715) );
  OAI21_X1 U16688 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n13261), .A(
        n13262), .ZN(n17243) );
  OAI21_X1 U16689 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n13264), .A(
        n13263), .ZN(n20324) );
  NOR2_X1 U16690 ( .A1(n18101), .A2(n16681), .ZN(n16667) );
  AND2_X1 U16691 ( .A1(n17212), .A2(n16667), .ZN(n16655) );
  NAND2_X1 U16692 ( .A1(n13260), .A2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13266) );
  INV_X1 U16693 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n13265) );
  NAND2_X1 U16694 ( .A1(n13266), .A2(n13265), .ZN(n13268) );
  NAND2_X1 U16695 ( .A1(n13268), .A2(n13267), .ZN(n17200) );
  NAND2_X1 U16696 ( .A1(n13267), .A2(n20307), .ZN(n13269) );
  AND2_X1 U16697 ( .A1(n13271), .A2(n13269), .ZN(n20311) );
  INV_X1 U16698 ( .A(n20311), .ZN(n13270) );
  AND2_X1 U16699 ( .A1(n13271), .A2(n17172), .ZN(n13272) );
  NOR2_X1 U16700 ( .A1(n13274), .A2(n13272), .ZN(n17174) );
  NOR2_X1 U16701 ( .A1(n13274), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13275) );
  OR2_X1 U16702 ( .A1(n13273), .A2(n13275), .ZN(n17161) );
  INV_X1 U16703 ( .A(n17161), .ZN(n16633) );
  NOR2_X1 U16704 ( .A1(n13273), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13276) );
  OR2_X1 U16705 ( .A1(n13277), .A2(n13276), .ZN(n17150) );
  AND2_X1 U16706 ( .A1(n16619), .A2(n17150), .ZN(n20296) );
  OR2_X1 U16707 ( .A1(n13277), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13278) );
  NAND2_X1 U16708 ( .A1(n13280), .A2(n13278), .ZN(n20297) );
  AND2_X1 U16709 ( .A1(n20296), .A2(n20297), .ZN(n20299) );
  NAND2_X1 U16710 ( .A1(n13280), .A2(n13279), .ZN(n13281) );
  NAND2_X1 U16711 ( .A1(n13282), .A2(n13281), .ZN(n17126) );
  NAND2_X1 U16712 ( .A1(n20299), .A2(n17126), .ZN(n20280) );
  AND2_X1 U16713 ( .A1(n13282), .A2(n20277), .ZN(n13283) );
  NOR2_X1 U16714 ( .A1(n13285), .A2(n13283), .ZN(n20281) );
  OR2_X1 U16715 ( .A1(n20280), .A2(n20281), .ZN(n20283) );
  OAI21_X1 U16716 ( .B1(n13285), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n13284), .ZN(n17100) );
  INV_X1 U16717 ( .A(n17100), .ZN(n13286) );
  NAND2_X1 U16718 ( .A1(n13232), .A2(n13284), .ZN(n13287) );
  NAND2_X1 U16719 ( .A1(n13288), .A2(n13287), .ZN(n17090) );
  INV_X1 U16720 ( .A(n13289), .ZN(n13293) );
  NAND2_X1 U16721 ( .A1(n13290), .A2(n17071), .ZN(n13291) );
  NAND2_X1 U16722 ( .A1(n13293), .A2(n13291), .ZN(n17069) );
  AND2_X1 U16723 ( .A1(n20266), .A2(n17069), .ZN(n20269) );
  INV_X1 U16724 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n16539) );
  NAND2_X1 U16725 ( .A1(n13293), .A2(n16539), .ZN(n13294) );
  NAND2_X1 U16726 ( .A1(n13292), .A2(n13294), .ZN(n17062) );
  NAND2_X1 U16727 ( .A1(n20269), .A2(n17062), .ZN(n13295) );
  NAND2_X1 U16728 ( .A1(n13292), .A2(n17049), .ZN(n13296) );
  AND2_X1 U16729 ( .A1(n13298), .A2(n13296), .ZN(n17053) );
  NAND2_X1 U16730 ( .A1(n13298), .A2(n13297), .ZN(n13299) );
  NAND2_X1 U16731 ( .A1(n13301), .A2(n13299), .ZN(n17043) );
  INV_X1 U16732 ( .A(n13300), .ZN(n13305) );
  NAND2_X1 U16733 ( .A1(n13301), .A2(n17030), .ZN(n13302) );
  AND2_X1 U16734 ( .A1(n13305), .A2(n13302), .ZN(n17028) );
  INV_X1 U16735 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n13304) );
  NAND2_X1 U16736 ( .A1(n13305), .A2(n13304), .ZN(n13306) );
  NAND2_X1 U16737 ( .A1(n13303), .A2(n13306), .ZN(n17022) );
  AOI21_X1 U16738 ( .B1(n16487), .B2(n17022), .A(n10160), .ZN(n16470) );
  NAND2_X1 U16739 ( .A1(n13303), .A2(n17012), .ZN(n13307) );
  AND2_X1 U16740 ( .A1(n13310), .A2(n13307), .ZN(n17014) );
  NOR2_X2 U16741 ( .A1(n16470), .A2(n17014), .ZN(n16457) );
  INV_X1 U16742 ( .A(n13308), .ZN(n13313) );
  NAND2_X1 U16743 ( .A1(n13310), .A2(n13309), .ZN(n13311) );
  NAND2_X1 U16744 ( .A1(n13313), .A2(n13311), .ZN(n17004) );
  AOI21_X2 U16745 ( .B1(n16457), .B2(n17004), .A(n10160), .ZN(n16443) );
  INV_X1 U16746 ( .A(n13312), .ZN(n13315) );
  INV_X1 U16747 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n22083) );
  NAND2_X1 U16748 ( .A1(n13313), .A2(n22083), .ZN(n13314) );
  NAND2_X1 U16749 ( .A1(n13315), .A2(n10488), .ZN(n13316) );
  NAND2_X1 U16750 ( .A1(n13317), .A2(n13316), .ZN(n16980) );
  NAND2_X1 U16751 ( .A1(n13317), .A2(n16972), .ZN(n13318) );
  AND2_X1 U16752 ( .A1(n13319), .A2(n13318), .ZN(n16975) );
  NOR2_X1 U16753 ( .A1(n16426), .A2(n16975), .ZN(n13320) );
  XNOR2_X1 U16754 ( .A(n13319), .B(n13336), .ZN(n15355) );
  OAI21_X1 U16755 ( .B1(n13320), .B2(n15355), .A(n20326), .ZN(n13322) );
  OAI21_X2 U16756 ( .B1(n13320), .B2(n10160), .A(n15355), .ZN(n15367) );
  INV_X1 U16757 ( .A(n15367), .ZN(n13321) );
  AOI21_X1 U16758 ( .B1(n16742), .B2(n13322), .A(n13321), .ZN(n13341) );
  INV_X1 U16759 ( .A(n16423), .ZN(n13325) );
  NAND2_X1 U16760 ( .A1(n14733), .A2(n13326), .ZN(n14747) );
  INV_X1 U16761 ( .A(n14747), .ZN(n13323) );
  AND2_X1 U16762 ( .A1(n13323), .A2(n16419), .ZN(n13324) );
  INV_X1 U16763 ( .A(n13326), .ZN(n13331) );
  NAND3_X1 U16764 ( .A1(n12207), .A2(P2_EBX_REG_31__SCAN_IN), .A3(n13331), 
        .ZN(n13327) );
  NOR2_X1 U16765 ( .A1(n20834), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20647) );
  INV_X1 U16766 ( .A(n20647), .ZN(n13328) );
  NOR2_X1 U16767 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n13328), .ZN(n13329) );
  NAND2_X1 U16768 ( .A1(n13329), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n18130) );
  AND3_X1 U16769 ( .A1(n14870), .A2(n13332), .A3(n13331), .ZN(n13333) );
  AOI21_X1 U16770 ( .B1(n14747), .B2(n16419), .A(n13333), .ZN(n13334) );
  OR2_X2 U16771 ( .A1(n16423), .A2(n13334), .ZN(n20335) );
  INV_X1 U16772 ( .A(n20335), .ZN(n20295) );
  AOI22_X1 U16773 ( .A1(P2_EBX_REG_30__SCAN_IN), .A2(n20295), .B1(n20344), 
        .B2(P2_REIP_REG_30__SCAN_IN), .ZN(n13335) );
  OAI21_X1 U16774 ( .B1(n13336), .B2(n20339), .A(n13335), .ZN(n13337) );
  INV_X1 U16775 ( .A(n17168), .ZN(n13345) );
  NAND2_X1 U16776 ( .A1(n17144), .A2(n17155), .ZN(n13347) );
  INV_X1 U16777 ( .A(n17121), .ZN(n17107) );
  OAI21_X1 U16778 ( .B1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(n13348), .ZN(n13349) );
  NAND2_X1 U16779 ( .A1(n13353), .A2(n13352), .ZN(n17088) );
  INV_X1 U16780 ( .A(n13354), .ZN(n13355) );
  NAND2_X1 U16781 ( .A1(n13357), .A2(n13356), .ZN(n13358) );
  XNOR2_X1 U16782 ( .A(n13359), .B(n13358), .ZN(n17047) );
  NAND2_X1 U16783 ( .A1(n17047), .A2(n18118), .ZN(n13377) );
  INV_X1 U16784 ( .A(n13360), .ZN(n17327) );
  AOI21_X1 U16785 ( .B1(n13366), .B2(n13364), .A(n13365), .ZN(n16909) );
  NAND2_X1 U16786 ( .A1(n10205), .A2(n13368), .ZN(n13367) );
  AND2_X1 U16787 ( .A1(n17453), .A2(n13367), .ZN(n17302) );
  NAND2_X1 U16788 ( .A1(n20343), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n17048) );
  INV_X1 U16789 ( .A(n13368), .ZN(n13369) );
  NAND3_X1 U16790 ( .A1(n17457), .A2(n13369), .A3(n13370), .ZN(n17301) );
  OAI211_X1 U16791 ( .C1(n17302), .C2(n13370), .A(n17048), .B(n17301), .ZN(
        n13375) );
  OAI21_X1 U16792 ( .B1(n13371), .B2(n13373), .A(n13372), .ZN(n17050) );
  NOR2_X1 U16793 ( .A1(n17050), .A2(n17518), .ZN(n13374) );
  AOI211_X1 U16794 ( .C1(n17505), .C2(n16909), .A(n13375), .B(n13374), .ZN(
        n13376) );
  NAND2_X1 U16795 ( .A1(n10451), .A2(n18598), .ZN(n18525) );
  NOR3_X1 U16796 ( .A1(n17802), .A2(n13378), .A3(n18525), .ZN(n13392) );
  INV_X1 U16797 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n18610) );
  AND2_X1 U16798 ( .A1(n13379), .A2(n18610), .ZN(n13391) );
  INV_X1 U16799 ( .A(n13380), .ZN(n13381) );
  INV_X1 U16800 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n20186) );
  AOI21_X1 U16801 ( .B1(n18269), .B2(n13381), .A(n20186), .ZN(n13382) );
  INV_X1 U16802 ( .A(n13382), .ZN(n13389) );
  NOR3_X1 U16803 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n22051), .A3(n13383), 
        .ZN(n13384) );
  AOI21_X1 U16804 ( .B1(n18596), .B2(P3_EBX_REG_31__SCAN_IN), .A(n13384), .ZN(
        n13385) );
  INV_X1 U16805 ( .A(n13385), .ZN(n13387) );
  INV_X1 U16806 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n17787) );
  NOR2_X1 U16807 ( .A1(n18593), .A2(n17787), .ZN(n13386) );
  NAND2_X1 U16808 ( .A1(n13126), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13394) );
  NAND2_X1 U16809 ( .A1(n13127), .A2(P2_EAX_REG_31__SCAN_IN), .ZN(n13393) );
  OAI211_X1 U16810 ( .C1(n13106), .C2(n13395), .A(n13394), .B(n13393), .ZN(
        n13396) );
  NAND2_X1 U16811 ( .A1(n15361), .A2(n17505), .ZN(n13408) );
  INV_X1 U16812 ( .A(n17282), .ZN(n13399) );
  INV_X1 U16813 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13398) );
  AOI21_X1 U16814 ( .B1(n13399), .B2(n18129), .A(n13398), .ZN(n13406) );
  NOR4_X1 U16815 ( .A1(n13402), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n13401), .A4(n13400), .ZN(n13403) );
  AOI211_X1 U16816 ( .C1(n13406), .C2(n13405), .A(n13404), .B(n13403), .ZN(
        n13407) );
  OAI211_X1 U16817 ( .C1(n15359), .C2(n17518), .A(n13408), .B(n13407), .ZN(
        n13411) );
  NOR2_X1 U16818 ( .A1(n13411), .A2(n13410), .ZN(n13412) );
  OAI21_X1 U16819 ( .B1(n13413), .B2(n17500), .A(n13412), .ZN(P2_U3015) );
  NAND2_X1 U16820 ( .A1(n13414), .A2(n15651), .ZN(n13806) );
  OR2_X1 U16821 ( .A1(n11794), .A2(n21822), .ZN(n13415) );
  NAND2_X1 U16822 ( .A1(n18086), .A2(n13417), .ZN(n13418) );
  AND4_X1 U16823 ( .A1(n14069), .A2(n10795), .A3(n13800), .A4(n10799), .ZN(
        n14065) );
  NAND2_X1 U16824 ( .A1(n13420), .A2(n14065), .ZN(n13421) );
  AND2_X1 U16825 ( .A1(n15786), .A2(n14069), .ZN(n13424) );
  NAND2_X1 U16826 ( .A1(n13425), .A2(n13424), .ZN(n13441) );
  NAND2_X1 U16827 ( .A1(n15781), .A2(n10792), .ZN(n14596) );
  NOR4_X1 U16828 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(
        P1_ADDRESS_REG_15__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_13__SCAN_IN), .ZN(n13429) );
  NOR4_X1 U16829 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_20__SCAN_IN), .A3(P1_ADDRESS_REG_19__SCAN_IN), .A4(
        P1_ADDRESS_REG_18__SCAN_IN), .ZN(n13428) );
  NOR4_X1 U16830 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(
        P1_ADDRESS_REG_6__SCAN_IN), .A3(P1_ADDRESS_REG_5__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13427) );
  NOR4_X1 U16831 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(
        P1_ADDRESS_REG_11__SCAN_IN), .A3(P1_ADDRESS_REG_10__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n13426) );
  AND4_X1 U16832 ( .A1(n13429), .A2(n13428), .A3(n13427), .A4(n13426), .ZN(
        n13434) );
  NOR4_X1 U16833 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_4__SCAN_IN), .ZN(n13432) );
  NOR4_X1 U16834 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n13431) );
  NOR4_X1 U16835 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n13430) );
  INV_X1 U16836 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n21754) );
  AND4_X1 U16837 ( .A1(n13432), .A2(n13431), .A3(n13430), .A4(n21754), .ZN(
        n13433) );
  NAND2_X1 U16838 ( .A1(n13434), .A2(n13433), .ZN(n13435) );
  AOI22_X1 U16839 ( .A1(n13436), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n13423), .ZN(n13437) );
  INV_X1 U16840 ( .A(n13437), .ZN(n13439) );
  INV_X1 U16841 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n18147) );
  NOR2_X1 U16842 ( .A1(n13439), .A2(n13438), .ZN(n13440) );
  NAND2_X1 U16843 ( .A1(n13441), .A2(n13440), .ZN(P1_U2873) );
  NOR2_X1 U16844 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13443) );
  NOR4_X1 U16845 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13442) );
  NAND4_X1 U16846 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13443), .A4(n13442), .ZN(n13456) );
  INV_X1 U16847 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21816) );
  NOR3_X1 U16848 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n21816), .ZN(n13445) );
  NOR4_X1 U16849 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13444) );
  NAND4_X1 U16850 ( .A1(n15020), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13445), .A4(
        n13444), .ZN(U214) );
  NOR4_X1 U16851 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n13449) );
  NOR4_X1 U16852 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n13448) );
  NOR4_X1 U16853 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n13447) );
  NOR4_X1 U16854 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_7__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n13446) );
  AND4_X1 U16855 ( .A1(n13449), .A2(n13448), .A3(n13447), .A4(n13446), .ZN(
        n13454) );
  NOR4_X1 U16856 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_1__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n13452) );
  NOR4_X1 U16857 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n13451) );
  NOR4_X1 U16858 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n13450) );
  INV_X1 U16859 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20978) );
  AND4_X1 U16860 ( .A1(n13452), .A2(n13451), .A3(n13450), .A4(n20978), .ZN(
        n13453) );
  NAND2_X1 U16861 ( .A1(n13454), .A2(n13453), .ZN(n13455) );
  NOR2_X1 U16862 ( .A1(n15338), .A2(n13456), .ZN(n18146) );
  NAND2_X1 U16863 ( .A1(n18146), .A2(U214), .ZN(U212) );
  INV_X1 U16864 ( .A(n20959), .ZN(n17597) );
  NAND2_X1 U16865 ( .A1(n17597), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13458) );
  INV_X1 U16866 ( .A(n13457), .ZN(n21044) );
  MUX2_X1 U16867 ( .A(n13458), .B(n21044), .S(n17596), .Z(n13460) );
  NAND2_X1 U16868 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n14857) );
  INV_X1 U16869 ( .A(n14857), .ZN(n13459) );
  NAND2_X1 U16870 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13459), .ZN(n18041) );
  INV_X1 U16871 ( .A(n18041), .ZN(n18133) );
  AOI21_X1 U16872 ( .B1(n13460), .B2(n20900), .A(n18133), .ZN(P2_U3178) );
  NOR2_X1 U16873 ( .A1(n13461), .A2(n13621), .ZN(n20348) );
  INV_X1 U16874 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n13463) );
  NOR2_X1 U16875 ( .A1(n13461), .A2(n10116), .ZN(n13468) );
  NAND2_X1 U16876 ( .A1(n13468), .A2(n14870), .ZN(n13469) );
  AND2_X1 U16877 ( .A1(n21042), .A2(n17538), .ZN(n13464) );
  INV_X1 U16878 ( .A(n13464), .ZN(n13462) );
  OAI211_X1 U16879 ( .C1(n20348), .C2(n13463), .A(n13469), .B(n13462), .ZN(
        P2_U2814) );
  INV_X1 U16880 ( .A(n13142), .ZN(n13466) );
  OAI21_X1 U16881 ( .B1(n13464), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n16423), 
        .ZN(n13465) );
  OAI21_X1 U16882 ( .B1(n13466), .B2(n16423), .A(n13465), .ZN(P2_U3612) );
  INV_X1 U16883 ( .A(n17545), .ZN(n17553) );
  NOR2_X1 U16884 ( .A1(n17553), .A2(n17596), .ZN(n17595) );
  AOI22_X1 U16885 ( .A1(n16423), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n17595), 
        .B2(n20900), .ZN(n13467) );
  INV_X1 U16886 ( .A(n13467), .ZN(P2_U2816) );
  INV_X1 U16887 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n20398) );
  OR2_X1 U16888 ( .A1(n13469), .A2(n20959), .ZN(n13472) );
  OR2_X1 U16889 ( .A1(n13472), .A2(n15209), .ZN(n13479) );
  INV_X1 U16890 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n14327) );
  OR2_X1 U16891 ( .A1(n15338), .A2(n14327), .ZN(n13471) );
  NAND2_X1 U16892 ( .A1(n15338), .A2(BUF2_REG_15__SCAN_IN), .ZN(n13470) );
  AND2_X1 U16893 ( .A1(n13471), .A2(n13470), .ZN(n16955) );
  NAND2_X1 U16894 ( .A1(n13472), .A2(n13625), .ZN(n20432) );
  INV_X1 U16895 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13473) );
  OAI222_X1 U16896 ( .A1(n13625), .A2(n20398), .B1(n13479), .B2(n16955), .C1(
        n20432), .C2(n13473), .ZN(P2_U2982) );
  INV_X1 U16897 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n20407) );
  INV_X1 U16898 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n18180) );
  OR2_X1 U16899 ( .A1(n15338), .A2(n18180), .ZN(n13475) );
  NAND2_X1 U16900 ( .A1(n15338), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13474) );
  NAND2_X1 U16901 ( .A1(n13475), .A2(n13474), .ZN(n16869) );
  INV_X1 U16902 ( .A(n16869), .ZN(n13476) );
  NOR2_X1 U16903 ( .A1(n13479), .A2(n13476), .ZN(n20429) );
  INV_X1 U16904 ( .A(n20429), .ZN(n13478) );
  NAND2_X1 U16905 ( .A1(n13533), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13477) );
  OAI211_X1 U16906 ( .C1(n20407), .C2(n13625), .A(n13478), .B(n13477), .ZN(
        P2_U2977) );
  INV_X2 U16907 ( .A(n13625), .ZN(n20430) );
  AOI22_X1 U16908 ( .A1(n13533), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_5__SCAN_IN), .B2(n20430), .ZN(n13483) );
  INV_X1 U16909 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n14574) );
  OR2_X1 U16910 ( .A1(n15338), .A2(n14574), .ZN(n13481) );
  NAND2_X1 U16911 ( .A1(n15338), .A2(BUF2_REG_5__SCAN_IN), .ZN(n13480) );
  AND2_X1 U16912 ( .A1(n13481), .A2(n13480), .ZN(n20443) );
  INV_X1 U16913 ( .A(n20443), .ZN(n13482) );
  NAND2_X1 U16914 ( .A1(n13550), .A2(n13482), .ZN(n13542) );
  NAND2_X1 U16915 ( .A1(n13483), .A2(n13542), .ZN(P2_U2972) );
  AOI22_X1 U16916 ( .A1(n13533), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_13__SCAN_IN), .B2(n20430), .ZN(n13486) );
  INV_X1 U16917 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n14670) );
  OR2_X1 U16918 ( .A1(n15338), .A2(n14670), .ZN(n13485) );
  NAND2_X1 U16919 ( .A1(n15338), .A2(BUF2_REG_13__SCAN_IN), .ZN(n13484) );
  NAND2_X1 U16920 ( .A1(n13485), .A2(n13484), .ZN(n16846) );
  NAND2_X1 U16921 ( .A1(n13550), .A2(n16846), .ZN(n13546) );
  NAND2_X1 U16922 ( .A1(n13486), .A2(n13546), .ZN(P2_U2980) );
  AOI22_X1 U16923 ( .A1(n13533), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(
        P2_EAX_REG_17__SCAN_IN), .B2(n20430), .ZN(n13491) );
  INV_X1 U16924 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n13487) );
  OR2_X1 U16925 ( .A1(n15338), .A2(n13487), .ZN(n13489) );
  NAND2_X1 U16926 ( .A1(n15338), .A2(BUF2_REG_1__SCAN_IN), .ZN(n13488) );
  AND2_X1 U16927 ( .A1(n13489), .A2(n13488), .ZN(n20394) );
  INV_X1 U16928 ( .A(n20394), .ZN(n13490) );
  NAND2_X1 U16929 ( .A1(n13550), .A2(n13490), .ZN(n13495) );
  NAND2_X1 U16930 ( .A1(n13491), .A2(n13495), .ZN(P2_U2953) );
  AOI22_X1 U16931 ( .A1(n13533), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_12__SCAN_IN), .B2(n20430), .ZN(n13494) );
  INV_X1 U16932 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n14271) );
  OR2_X1 U16933 ( .A1(n15338), .A2(n14271), .ZN(n13493) );
  NAND2_X1 U16934 ( .A1(n15338), .A2(BUF2_REG_12__SCAN_IN), .ZN(n13492) );
  NAND2_X1 U16935 ( .A1(n13493), .A2(n13492), .ZN(n16854) );
  NAND2_X1 U16936 ( .A1(n13550), .A2(n16854), .ZN(n13540) );
  NAND2_X1 U16937 ( .A1(n13494), .A2(n13540), .ZN(P2_U2979) );
  AOI22_X1 U16938 ( .A1(n13533), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(
        P2_EAX_REG_1__SCAN_IN), .B2(n20430), .ZN(n13496) );
  NAND2_X1 U16939 ( .A1(n13496), .A2(n13495), .ZN(P2_U2968) );
  AOI22_X1 U16940 ( .A1(n13533), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_4__SCAN_IN), .B2(n20430), .ZN(n13499) );
  INV_X1 U16941 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n14259) );
  OR2_X1 U16942 ( .A1(n15338), .A2(n14259), .ZN(n13498) );
  NAND2_X1 U16943 ( .A1(n15338), .A2(BUF2_REG_4__SCAN_IN), .ZN(n13497) );
  AND2_X1 U16944 ( .A1(n13498), .A2(n13497), .ZN(n20377) );
  INV_X1 U16945 ( .A(n20377), .ZN(n16918) );
  NAND2_X1 U16946 ( .A1(n13550), .A2(n16918), .ZN(n13534) );
  NAND2_X1 U16947 ( .A1(n13499), .A2(n13534), .ZN(P2_U2971) );
  AOI22_X1 U16948 ( .A1(n13533), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_6__SCAN_IN), .B2(n20430), .ZN(n13503) );
  INV_X1 U16949 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n13500) );
  OR2_X1 U16950 ( .A1(n15338), .A2(n13500), .ZN(n13502) );
  NAND2_X1 U16951 ( .A1(n15338), .A2(BUF2_REG_6__SCAN_IN), .ZN(n13501) );
  NAND2_X1 U16952 ( .A1(n13502), .A2(n13501), .ZN(n16901) );
  NAND2_X1 U16953 ( .A1(n13550), .A2(n16901), .ZN(n13554) );
  NAND2_X1 U16954 ( .A1(n13503), .A2(n13554), .ZN(P2_U2973) );
  AOI22_X1 U16955 ( .A1(n13533), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(
        P2_EAX_REG_7__SCAN_IN), .B2(n20430), .ZN(n13507) );
  INV_X1 U16956 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n13504) );
  OR2_X1 U16957 ( .A1(n15338), .A2(n13504), .ZN(n13506) );
  NAND2_X1 U16958 ( .A1(n15338), .A2(BUF2_REG_7__SCAN_IN), .ZN(n13505) );
  NAND2_X1 U16959 ( .A1(n13506), .A2(n13505), .ZN(n16893) );
  NAND2_X1 U16960 ( .A1(n13550), .A2(n16893), .ZN(n13544) );
  NAND2_X1 U16961 ( .A1(n13507), .A2(n13544), .ZN(P2_U2974) );
  AOI22_X1 U16962 ( .A1(n13533), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_9__SCAN_IN), .B2(n20430), .ZN(n13510) );
  INV_X1 U16963 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n14319) );
  OR2_X1 U16964 ( .A1(n15338), .A2(n14319), .ZN(n13509) );
  NAND2_X1 U16965 ( .A1(n15338), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13508) );
  NAND2_X1 U16966 ( .A1(n13509), .A2(n13508), .ZN(n16877) );
  NAND2_X1 U16967 ( .A1(n13550), .A2(n16877), .ZN(n13552) );
  NAND2_X1 U16968 ( .A1(n13510), .A2(n13552), .ZN(P2_U2976) );
  AOI22_X1 U16969 ( .A1(n13533), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_2__SCAN_IN), .B2(n20430), .ZN(n13514) );
  INV_X1 U16970 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n13511) );
  OR2_X1 U16971 ( .A1(n15338), .A2(n13511), .ZN(n13513) );
  NAND2_X1 U16972 ( .A1(n15338), .A2(BUF2_REG_2__SCAN_IN), .ZN(n13512) );
  NAND2_X1 U16973 ( .A1(n13513), .A2(n13512), .ZN(n20434) );
  NAND2_X1 U16974 ( .A1(n13550), .A2(n20434), .ZN(n13538) );
  NAND2_X1 U16975 ( .A1(n13514), .A2(n13538), .ZN(P2_U2969) );
  AOI22_X1 U16976 ( .A1(n13533), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_3__SCAN_IN), .B2(n20430), .ZN(n13519) );
  INV_X1 U16977 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n13515) );
  OR2_X1 U16978 ( .A1(n15338), .A2(n13515), .ZN(n13517) );
  NAND2_X1 U16979 ( .A1(n15338), .A2(BUF2_REG_3__SCAN_IN), .ZN(n13516) );
  AND2_X1 U16980 ( .A1(n13517), .A2(n13516), .ZN(n20437) );
  INV_X1 U16981 ( .A(n20437), .ZN(n13518) );
  NAND2_X1 U16982 ( .A1(n13550), .A2(n13518), .ZN(n13536) );
  NAND2_X1 U16983 ( .A1(n13519), .A2(n13536), .ZN(P2_U2970) );
  AOI22_X1 U16984 ( .A1(n13533), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_11__SCAN_IN), .B2(n20430), .ZN(n13523) );
  INV_X1 U16985 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n13520) );
  OR2_X1 U16986 ( .A1(n15338), .A2(n13520), .ZN(n13522) );
  NAND2_X1 U16987 ( .A1(n15338), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13521) );
  NAND2_X1 U16988 ( .A1(n13522), .A2(n13521), .ZN(n16863) );
  NAND2_X1 U16989 ( .A1(n13550), .A2(n16863), .ZN(n13558) );
  NAND2_X1 U16990 ( .A1(n13523), .A2(n13558), .ZN(P2_U2978) );
  AOI22_X1 U16991 ( .A1(n13533), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n20430), 
        .B2(P2_EAX_REG_0__SCAN_IN), .ZN(n13527) );
  INV_X1 U16992 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n13524) );
  OR2_X1 U16993 ( .A1(n15338), .A2(n13524), .ZN(n13526) );
  NAND2_X1 U16994 ( .A1(n15338), .A2(BUF2_REG_0__SCAN_IN), .ZN(n13525) );
  NAND2_X1 U16995 ( .A1(n13526), .A2(n13525), .ZN(n20359) );
  NAND2_X1 U16996 ( .A1(n13550), .A2(n20359), .ZN(n13561) );
  NAND2_X1 U16997 ( .A1(n13527), .A2(n13561), .ZN(P2_U2967) );
  INV_X1 U16998 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13730) );
  INV_X1 U16999 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n15021) );
  OR2_X1 U17000 ( .A1(n15338), .A2(n15021), .ZN(n13529) );
  NAND2_X1 U17001 ( .A1(n15338), .A2(BUF2_REG_14__SCAN_IN), .ZN(n13528) );
  NAND2_X1 U17002 ( .A1(n13529), .A2(n13528), .ZN(n15340) );
  NAND2_X1 U17003 ( .A1(n13550), .A2(n15340), .ZN(n13532) );
  NAND2_X1 U17004 ( .A1(n13533), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13530) );
  OAI211_X1 U17005 ( .C1(n13730), .C2(n13625), .A(n13532), .B(n13530), .ZN(
        P2_U2966) );
  INV_X1 U17006 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n20400) );
  NAND2_X1 U17007 ( .A1(n13533), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n13531) );
  OAI211_X1 U17008 ( .C1(n20400), .C2(n13625), .A(n13532), .B(n13531), .ZN(
        P2_U2981) );
  AOI22_X1 U17009 ( .A1(n13533), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n20430), .ZN(n13535) );
  NAND2_X1 U17010 ( .A1(n13535), .A2(n13534), .ZN(P2_U2956) );
  AOI22_X1 U17011 ( .A1(n13533), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_19__SCAN_IN), .B2(n20430), .ZN(n13537) );
  NAND2_X1 U17012 ( .A1(n13537), .A2(n13536), .ZN(P2_U2955) );
  AOI22_X1 U17013 ( .A1(n13533), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_18__SCAN_IN), .B2(n20430), .ZN(n13539) );
  NAND2_X1 U17014 ( .A1(n13539), .A2(n13538), .ZN(P2_U2954) );
  AOI22_X1 U17015 ( .A1(n13533), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_28__SCAN_IN), .B2(n20430), .ZN(n13541) );
  NAND2_X1 U17016 ( .A1(n13541), .A2(n13540), .ZN(P2_U2964) );
  AOI22_X1 U17017 ( .A1(n13533), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_21__SCAN_IN), .B2(n20430), .ZN(n13543) );
  NAND2_X1 U17018 ( .A1(n13543), .A2(n13542), .ZN(P2_U2957) );
  AOI22_X1 U17019 ( .A1(n13533), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(
        P2_EAX_REG_23__SCAN_IN), .B2(n20430), .ZN(n13545) );
  NAND2_X1 U17020 ( .A1(n13545), .A2(n13544), .ZN(P2_U2959) );
  AOI22_X1 U17021 ( .A1(n13533), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n20430), .ZN(n13547) );
  NAND2_X1 U17022 ( .A1(n13547), .A2(n13546), .ZN(P2_U2965) );
  AOI22_X1 U17023 ( .A1(n13533), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_24__SCAN_IN), .B2(n20430), .ZN(n13551) );
  INV_X1 U17024 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n14309) );
  OR2_X1 U17025 ( .A1(n15338), .A2(n14309), .ZN(n13549) );
  NAND2_X1 U17026 ( .A1(n15338), .A2(BUF2_REG_8__SCAN_IN), .ZN(n13548) );
  NAND2_X1 U17027 ( .A1(n13549), .A2(n13548), .ZN(n16885) );
  NAND2_X1 U17028 ( .A1(n13550), .A2(n16885), .ZN(n13556) );
  NAND2_X1 U17029 ( .A1(n13551), .A2(n13556), .ZN(P2_U2960) );
  AOI22_X1 U17030 ( .A1(n13533), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_25__SCAN_IN), .B2(n20430), .ZN(n13553) );
  NAND2_X1 U17031 ( .A1(n13553), .A2(n13552), .ZN(P2_U2961) );
  AOI22_X1 U17032 ( .A1(n13533), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n20430), .ZN(n13555) );
  NAND2_X1 U17033 ( .A1(n13555), .A2(n13554), .ZN(P2_U2958) );
  AOI22_X1 U17034 ( .A1(n13533), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_8__SCAN_IN), .B2(n20430), .ZN(n13557) );
  NAND2_X1 U17035 ( .A1(n13557), .A2(n13556), .ZN(P2_U2975) );
  AOI22_X1 U17036 ( .A1(n13533), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n20430), .ZN(n13559) );
  NAND2_X1 U17037 ( .A1(n13559), .A2(n13558), .ZN(P2_U2963) );
  INV_X1 U17038 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n22094) );
  NAND2_X1 U17039 ( .A1(n13533), .A2(P2_UWORD_REG_0__SCAN_IN), .ZN(n13560) );
  OAI211_X1 U17040 ( .C1(n22094), .C2(n13625), .A(n13561), .B(n13560), .ZN(
        P2_U2952) );
  INV_X1 U17041 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13581) );
  NAND2_X1 U17042 ( .A1(n17992), .A2(n13562), .ZN(n13567) );
  INV_X1 U17043 ( .A(n13563), .ZN(n13565) );
  NAND2_X1 U17044 ( .A1(n13565), .A2(n13564), .ZN(n13566) );
  NAND2_X1 U17045 ( .A1(n13567), .A2(n13566), .ZN(n21100) );
  NAND2_X1 U17046 ( .A1(n21825), .A2(n11806), .ZN(n13568) );
  AOI21_X1 U17047 ( .B1(n13568), .B2(n18039), .A(n21822), .ZN(n21824) );
  OR2_X1 U17048 ( .A1(n21100), .A2(n21824), .ZN(n18013) );
  AND2_X1 U17049 ( .A1(n18013), .A2(n13800), .ZN(n21107) );
  INV_X1 U17050 ( .A(n13807), .ZN(n13572) );
  MUX2_X1 U17051 ( .A(n13572), .B(n13571), .S(n17992), .Z(n13577) );
  INV_X1 U17052 ( .A(n13573), .ZN(n13574) );
  AND2_X1 U17053 ( .A1(n13575), .A2(n13574), .ZN(n13576) );
  OR2_X1 U17054 ( .A1(n13577), .A2(n13576), .ZN(n13578) );
  NAND2_X1 U17055 ( .A1(n13578), .A2(n14591), .ZN(n18012) );
  INV_X1 U17056 ( .A(n18012), .ZN(n13579) );
  NAND2_X1 U17057 ( .A1(n13579), .A2(n21107), .ZN(n13580) );
  OAI21_X1 U17058 ( .B1(n13581), .B2(n21107), .A(n13580), .ZN(P1_U3484) );
  INV_X1 U17059 ( .A(n13582), .ZN(n13585) );
  AOI21_X1 U17060 ( .B1(n13585), .B2(n13584), .A(n13583), .ZN(n18125) );
  NOR2_X1 U17061 ( .A1(n20260), .A2(n12235), .ZN(n18119) );
  OAI21_X1 U17062 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n16735), .A(
        n13586), .ZN(n18114) );
  NOR2_X1 U17063 ( .A1(n17252), .A2(n18114), .ZN(n13587) );
  AOI211_X1 U17064 ( .C1(n18125), .C2(n18108), .A(n18119), .B(n13587), .ZN(
        n13590) );
  OAI21_X1 U17065 ( .B1(n17214), .B2(n13588), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13589) );
  OAI211_X1 U17066 ( .C1(n13833), .C2(n17242), .A(n13590), .B(n13589), .ZN(
        P2_U3014) );
  INV_X1 U17067 ( .A(n13591), .ZN(n13593) );
  XNOR2_X1 U17068 ( .A(n13593), .B(n13592), .ZN(n13978) );
  NOR2_X1 U17069 ( .A1(n20260), .A2(n20981), .ZN(n13977) );
  AOI21_X1 U17070 ( .B1(n17214), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n13977), .ZN(n13597) );
  OR2_X1 U17071 ( .A1(n13595), .A2(n13594), .ZN(n13971) );
  NAND3_X1 U17072 ( .A1(n13971), .A2(n13972), .A3(n18108), .ZN(n13596) );
  OAI211_X1 U17073 ( .C1(n17244), .C2(n10154), .A(n13597), .B(n13596), .ZN(
        n13598) );
  AOI21_X1 U17074 ( .B1(n18105), .B2(n13978), .A(n13598), .ZN(n13599) );
  OAI21_X1 U17075 ( .B1(n12275), .B2(n17242), .A(n13599), .ZN(P2_U3012) );
  NAND2_X1 U17076 ( .A1(n13601), .A2(n13600), .ZN(n13602) );
  XNOR2_X1 U17077 ( .A(n13602), .B(n14087), .ZN(n14088) );
  OAI21_X1 U17078 ( .B1(n13604), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n13603), .ZN(n14094) );
  OR2_X1 U17079 ( .A1(n13139), .A2(n20979), .ZN(n14086) );
  OAI21_X1 U17080 ( .B1(n17218), .B2(n14094), .A(n14086), .ZN(n13606) );
  NOR2_X1 U17081 ( .A1(n17244), .A2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13605) );
  AOI211_X1 U17082 ( .C1(n17214), .C2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13606), .B(n13605), .ZN(n13608) );
  NAND2_X1 U17083 ( .A1(n16718), .A2(n18107), .ZN(n13607) );
  OAI211_X1 U17084 ( .C1(n14088), .C2(n17252), .A(n13608), .B(n13607), .ZN(
        P2_U3013) );
  INV_X1 U17085 ( .A(n13621), .ZN(n13624) );
  NAND2_X1 U17086 ( .A1(n13624), .A2(n13609), .ZN(n13616) );
  NAND3_X1 U17087 ( .A1(n13610), .A2(n13142), .A3(n14736), .ZN(n13611) );
  INV_X1 U17088 ( .A(n14425), .ZN(n13615) );
  INV_X1 U17089 ( .A(n14730), .ZN(n13612) );
  NAND2_X1 U17090 ( .A1(n14731), .A2(n13612), .ZN(n13830) );
  AND2_X1 U17091 ( .A1(n13830), .A2(n13613), .ZN(n13614) );
  OAI211_X1 U17092 ( .C1(n13627), .C2(n13616), .A(n13615), .B(n13614), .ZN(
        n14743) );
  NAND2_X1 U17093 ( .A1(n17596), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13617) );
  OAI21_X1 U17094 ( .B1(n18041), .B2(n12578), .A(n13617), .ZN(n13618) );
  INV_X1 U17095 ( .A(n17555), .ZN(n13623) );
  NAND2_X1 U17096 ( .A1(n15209), .A2(n13619), .ZN(n13620) );
  OR2_X1 U17097 ( .A1(n13621), .A2(n13620), .ZN(n14737) );
  OR3_X1 U17098 ( .A1(n17555), .A2(n14737), .A3(n17553), .ZN(n13622) );
  OAI21_X1 U17099 ( .B1(n13623), .B2(n14742), .A(n13622), .ZN(P2_U3595) );
  NAND2_X1 U17100 ( .A1(n13624), .A2(n20237), .ZN(n13626) );
  OAI21_X1 U17101 ( .B1(n13627), .B2(n13626), .A(n13625), .ZN(n13628) );
  INV_X2 U17102 ( .A(n20419), .ZN(n20426) );
  INV_X1 U17103 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n13630) );
  INV_X1 U17104 ( .A(n13736), .ZN(n20395) );
  AOI22_X1 U17105 ( .A1(n20395), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n20426), 
        .B2(P2_UWORD_REG_1__SCAN_IN), .ZN(n13629) );
  OAI21_X1 U17106 ( .B1(n13711), .B2(n13630), .A(n13629), .ZN(P2_U2934) );
  NAND2_X1 U17107 ( .A1(n14457), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n13634) );
  NAND2_X1 U17108 ( .A1(n9712), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n13633) );
  NAND2_X1 U17109 ( .A1(n9705), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n13632) );
  NAND2_X1 U17110 ( .A1(n18652), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n13631) );
  NAND2_X1 U17111 ( .A1(n18624), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n13638) );
  NAND2_X1 U17112 ( .A1(n14968), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13637) );
  INV_X1 U17113 ( .A(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14945) );
  OR2_X1 U17114 ( .A1(n18773), .A2(n14945), .ZN(n13636) );
  OR2_X1 U17115 ( .A1(n18775), .A2(n14943), .ZN(n13635) );
  INV_X2 U17116 ( .A(n13659), .ZN(n18763) );
  NAND2_X1 U17117 ( .A1(n14896), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n13639) );
  OAI21_X1 U17118 ( .B1(n17689), .B2(n18763), .A(n13639), .ZN(n13641) );
  INV_X1 U17119 ( .A(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17697) );
  INV_X1 U17120 ( .A(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14952) );
  OAI22_X1 U17121 ( .A1(n17695), .A2(n17697), .B1(n11974), .B2(n14952), .ZN(
        n13640) );
  NOR2_X1 U17122 ( .A1(n13641), .A2(n13640), .ZN(n13648) );
  NAND2_X1 U17123 ( .A1(n17693), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n13646) );
  NAND2_X1 U17124 ( .A1(n17631), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n13645) );
  NAND2_X1 U17125 ( .A1(n17630), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n13644) );
  INV_X1 U17126 ( .A(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13642) );
  OR2_X1 U17127 ( .A1(n18715), .A2(n13642), .ZN(n13643) );
  NAND4_X2 U17128 ( .A1(n13650), .A2(n13649), .A3(n13648), .A4(n13647), .ZN(
        n14188) );
  XNOR2_X1 U17129 ( .A(n14188), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13703) );
  NAND2_X1 U17130 ( .A1(n9712), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n13654) );
  NAND2_X1 U17131 ( .A1(n14457), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n13653) );
  NAND2_X1 U17132 ( .A1(n9705), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n13652) );
  NAND2_X1 U17133 ( .A1(n18652), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n13651) );
  AND4_X1 U17134 ( .A1(n13654), .A2(n13653), .A3(n13652), .A4(n13651), .ZN(
        n13669) );
  NAND2_X1 U17135 ( .A1(n18624), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n13658) );
  NAND2_X1 U17136 ( .A1(n14968), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13657) );
  OR2_X1 U17137 ( .A1(n18775), .A2(n18756), .ZN(n13656) );
  INV_X1 U17138 ( .A(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n18752) );
  OR2_X1 U17139 ( .A1(n18773), .A2(n18752), .ZN(n13655) );
  AND4_X1 U17140 ( .A1(n13658), .A2(n13657), .A3(n13656), .A4(n13655), .ZN(
        n13668) );
  INV_X2 U17141 ( .A(n14112), .ZN(n14983) );
  INV_X1 U17142 ( .A(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18762) );
  OAI22_X1 U17143 ( .A1(n18613), .A2(n19819), .B1(n14983), .B2(n18762), .ZN(
        n13661) );
  INV_X1 U17144 ( .A(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n18776) );
  OAI22_X1 U17145 ( .A1(n18715), .A2(n18776), .B1(n18764), .B2(n18753), .ZN(
        n13660) );
  NOR2_X1 U17146 ( .A1(n13661), .A2(n13660), .ZN(n13667) );
  NAND2_X1 U17147 ( .A1(n14896), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n13665) );
  NAND2_X1 U17148 ( .A1(n17630), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n13664) );
  NAND2_X1 U17149 ( .A1(n17631), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n13663) );
  NAND2_X1 U17150 ( .A1(n17693), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n13662) );
  AND4_X1 U17151 ( .A1(n13665), .A2(n13664), .A3(n13663), .A4(n13662), .ZN(
        n13666) );
  NAND4_X1 U17152 ( .A1(n13669), .A2(n13668), .A3(n13667), .A4(n13666), .ZN(
        n14174) );
  OR2_X1 U17153 ( .A1(n14174), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13936) );
  XNOR2_X1 U17154 ( .A(n13703), .B(n13936), .ZN(n19339) );
  OR2_X1 U17155 ( .A1(n13690), .A2(n13674), .ZN(n13871) );
  INV_X1 U17156 ( .A(n13871), .ZN(n13773) );
  NOR2_X4 U17157 ( .A1(n19526), .A2(n20058), .ZN(n19438) );
  NOR2_X4 U17158 ( .A1(n19477), .A2(n18973), .ZN(n20057) );
  XNOR2_X1 U17159 ( .A(n13690), .B(n18973), .ZN(n13678) );
  AOI21_X1 U17160 ( .B1(n20215), .B2(n13678), .A(n20121), .ZN(n18241) );
  INV_X1 U17161 ( .A(n18241), .ZN(n13679) );
  NOR2_X1 U17162 ( .A1(n13680), .A2(n13679), .ZN(n13686) );
  INV_X1 U17163 ( .A(n13681), .ZN(n13683) );
  NAND2_X1 U17164 ( .A1(n13965), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n13682) );
  NAND2_X1 U17165 ( .A1(n13683), .A2(n13682), .ZN(n13693) );
  OR2_X1 U17166 ( .A1(n13697), .A2(n13693), .ZN(n13684) );
  AND3_X1 U17167 ( .A1(n19634), .A2(n13685), .A3(n18973), .ZN(n13849) );
  AOI22_X1 U17168 ( .A1(n20062), .A2(n13686), .B1(n20063), .B2(n13849), .ZN(
        n13701) );
  INV_X1 U17169 ( .A(n18235), .ZN(n18242) );
  INV_X1 U17170 ( .A(n13687), .ZN(n13705) );
  AOI211_X1 U17171 ( .C1(n18242), .C2(n13687), .A(n13689), .B(n13688), .ZN(
        n13780) );
  OAI21_X1 U17172 ( .B1(n13691), .B2(n13690), .A(n19642), .ZN(n13699) );
  INV_X1 U17173 ( .A(n13692), .ZN(n13695) );
  NAND2_X1 U17174 ( .A1(n13699), .A2(n20059), .ZN(n13700) );
  NAND3_X1 U17175 ( .A1(n13701), .A2(n13780), .A3(n13700), .ZN(n13702) );
  AND2_X1 U17176 ( .A1(n14174), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13935) );
  NAND2_X1 U17177 ( .A1(n13703), .A2(n13935), .ZN(n14192) );
  OAI21_X1 U17178 ( .B1(n13703), .B2(n13935), .A(n14192), .ZN(n19341) );
  AND3_X1 U17179 ( .A1(n13849), .A2(n19642), .A3(n18917), .ZN(n13704) );
  AND2_X1 U17180 ( .A1(n19477), .A2(n19598), .ZN(n19497) );
  INV_X1 U17181 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19590) );
  OAI211_X1 U17182 ( .C1(n19604), .C2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n19497), .B(n19590), .ZN(n13707) );
  AND2_X1 U17183 ( .A1(n19566), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n19338) );
  INV_X1 U17184 ( .A(n19338), .ZN(n13706) );
  OAI211_X1 U17185 ( .C1(n19341), .C2(n19605), .A(n13707), .B(n13706), .ZN(
        n13709) );
  INV_X1 U17186 ( .A(n19438), .ZN(n19427) );
  INV_X1 U17187 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19606) );
  NAND3_X1 U17188 ( .A1(n19598), .A2(n19427), .A3(n19606), .ZN(n19611) );
  AOI21_X1 U17189 ( .B1(n19564), .B2(n19611), .A(n19590), .ZN(n13708) );
  AOI211_X1 U17190 ( .C1(n19339), .C2(n19610), .A(n13709), .B(n13708), .ZN(
        n13710) );
  INV_X1 U17191 ( .A(n13710), .ZN(P3_U2861) );
  INV_X1 U17192 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13713) );
  AOI22_X1 U17193 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n20425), .B1(n20426), 
        .B2(P2_UWORD_REG_6__SCAN_IN), .ZN(n13712) );
  OAI21_X1 U17194 ( .B1(n13713), .B2(n13736), .A(n13712), .ZN(P2_U2929) );
  INV_X1 U17195 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n13715) );
  AOI22_X1 U17196 ( .A1(n20426), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n20425), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13714) );
  OAI21_X1 U17197 ( .B1(n13715), .B2(n13736), .A(n13714), .ZN(P2_U2932) );
  INV_X1 U17198 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13717) );
  AOI22_X1 U17199 ( .A1(n20426), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n20425), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13716) );
  OAI21_X1 U17200 ( .B1(n13717), .B2(n13736), .A(n13716), .ZN(P2_U2931) );
  INV_X1 U17201 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n13719) );
  AOI22_X1 U17202 ( .A1(n20426), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n20425), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13718) );
  OAI21_X1 U17203 ( .B1(n13719), .B2(n13736), .A(n13718), .ZN(P2_U2930) );
  INV_X1 U17204 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13721) );
  AOI22_X1 U17205 ( .A1(n20426), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n20425), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13720) );
  OAI21_X1 U17206 ( .B1(n13721), .B2(n13736), .A(n13720), .ZN(P2_U2927) );
  INV_X1 U17207 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n13723) );
  AOI22_X1 U17208 ( .A1(n20426), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n20425), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13722) );
  OAI21_X1 U17209 ( .B1(n13723), .B2(n13736), .A(n13722), .ZN(P2_U2926) );
  INV_X1 U17210 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n13725) );
  AOI22_X1 U17211 ( .A1(n20426), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n20425), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13724) );
  OAI21_X1 U17212 ( .B1(n13725), .B2(n13736), .A(n13724), .ZN(P2_U2924) );
  INV_X1 U17213 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13727) );
  AOI22_X1 U17214 ( .A1(n20426), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n20425), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13726) );
  OAI21_X1 U17215 ( .B1(n13727), .B2(n13736), .A(n13726), .ZN(P2_U2933) );
  AOI22_X1 U17216 ( .A1(n20426), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n20425), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13728) );
  OAI21_X1 U17217 ( .B1(n22094), .B2(n13736), .A(n13728), .ZN(P2_U2935) );
  AOI22_X1 U17218 ( .A1(n20426), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n20425), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n13729) );
  OAI21_X1 U17219 ( .B1(n13730), .B2(n13736), .A(n13729), .ZN(P2_U2921) );
  INV_X1 U17220 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n13732) );
  AOI22_X1 U17221 ( .A1(n20426), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n20425), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13731) );
  OAI21_X1 U17222 ( .B1(n13732), .B2(n13736), .A(n13731), .ZN(P2_U2928) );
  INV_X1 U17223 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n13734) );
  AOI22_X1 U17224 ( .A1(n20426), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n20425), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13733) );
  OAI21_X1 U17225 ( .B1(n13734), .B2(n13736), .A(n13733), .ZN(P2_U2923) );
  INV_X1 U17226 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n13737) );
  AOI22_X1 U17227 ( .A1(n20426), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n20425), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13735) );
  OAI21_X1 U17228 ( .B1(n13737), .B2(n13736), .A(n13735), .ZN(P2_U2922) );
  INV_X1 U17229 ( .A(n13738), .ZN(n13742) );
  INV_X1 U17230 ( .A(n13739), .ZN(n13741) );
  OAI21_X1 U17231 ( .B1(n13742), .B2(n13741), .A(n13740), .ZN(n15681) );
  INV_X1 U17232 ( .A(n13743), .ZN(n13745) );
  AOI21_X1 U17233 ( .B1(n13745), .B2(n21912), .A(n13744), .ZN(n14007) );
  INV_X1 U17234 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n21812) );
  NOR2_X1 U17235 ( .A1(n21291), .A2(n21812), .ZN(n14011) );
  INV_X1 U17236 ( .A(n13746), .ZN(n13748) );
  INV_X1 U17237 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13747) );
  AOI21_X1 U17238 ( .B1(n18061), .B2(n13748), .A(n13747), .ZN(n13749) );
  AOI211_X1 U17239 ( .C1(n14007), .C2(n11864), .A(n14011), .B(n13749), .ZN(
        n13750) );
  OAI21_X1 U17240 ( .B1(n18057), .B2(n15681), .A(n13750), .ZN(P1_U2999) );
  INV_X1 U17241 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13753) );
  AND2_X1 U17242 ( .A1(n17995), .A2(n18024), .ZN(n13751) );
  NAND2_X1 U17243 ( .A1(n21235), .A2(n9724), .ZN(n13789) );
  NAND2_X1 U17244 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n18095) );
  INV_X1 U17245 ( .A(n21234), .ZN(n21821) );
  NOR2_X4 U17246 ( .A1(n21235), .A2(n21254), .ZN(n21231) );
  AOI22_X1 U17247 ( .A1(n21234), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n21231), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13752) );
  OAI21_X1 U17248 ( .B1(n13753), .B2(n13789), .A(n13752), .ZN(P1_U2918) );
  AOI22_X1 U17249 ( .A1(n21254), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n21231), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13754) );
  OAI21_X1 U17250 ( .B1(n15734), .B2(n13789), .A(n13754), .ZN(P1_U2912) );
  INV_X1 U17251 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13756) );
  AOI22_X1 U17252 ( .A1(n21234), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n21231), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13755) );
  OAI21_X1 U17253 ( .B1(n13756), .B2(n13789), .A(n13755), .ZN(P1_U2916) );
  INV_X1 U17254 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13758) );
  AOI22_X1 U17255 ( .A1(n21234), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n21231), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13757) );
  OAI21_X1 U17256 ( .B1(n13758), .B2(n13789), .A(n13757), .ZN(P1_U2915) );
  INV_X1 U17257 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13760) );
  AOI22_X1 U17258 ( .A1(n21234), .A2(P1_UWORD_REG_0__SCAN_IN), .B1(n21231), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13759) );
  OAI21_X1 U17259 ( .B1(n13760), .B2(n13789), .A(n13759), .ZN(P1_U2920) );
  INV_X1 U17260 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13762) );
  AOI22_X1 U17261 ( .A1(n21234), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n21231), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13761) );
  OAI21_X1 U17262 ( .B1(n13762), .B2(n13789), .A(n13761), .ZN(P1_U2913) );
  INV_X1 U17263 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13764) );
  AOI22_X1 U17264 ( .A1(n21234), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n21231), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13763) );
  OAI21_X1 U17265 ( .B1(n13764), .B2(n13789), .A(n13763), .ZN(P1_U2917) );
  INV_X1 U17266 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n14326) );
  AOI22_X1 U17267 ( .A1(n21234), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n21231), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13765) );
  OAI21_X1 U17268 ( .B1(n14326), .B2(n13789), .A(n13765), .ZN(P1_U2909) );
  AOI22_X1 U17269 ( .A1(n21254), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n21231), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13766) );
  OAI21_X1 U17270 ( .B1(n15728), .B2(n13789), .A(n13766), .ZN(P1_U2911) );
  INV_X1 U17271 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13768) );
  AOI22_X1 U17272 ( .A1(n21234), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n21231), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13767) );
  OAI21_X1 U17273 ( .B1(n13768), .B2(n13789), .A(n13767), .ZN(P1_U2914) );
  INV_X1 U17274 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n14316) );
  AOI22_X1 U17275 ( .A1(n21254), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n21231), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13769) );
  OAI21_X1 U17276 ( .B1(n14316), .B2(n13789), .A(n13769), .ZN(P1_U2910) );
  INV_X1 U17277 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n15710) );
  AOI22_X1 U17278 ( .A1(n21254), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n21231), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13770) );
  OAI21_X1 U17279 ( .B1(n15710), .B2(n13789), .A(n13770), .ZN(P1_U2907) );
  INV_X1 U17280 ( .A(n13771), .ZN(n13772) );
  AOI21_X1 U17281 ( .B1(n13773), .B2(n13772), .A(n10263), .ZN(n14029) );
  INV_X1 U17282 ( .A(n14029), .ZN(n13774) );
  AOI21_X1 U17283 ( .B1(n19604), .B2(n13775), .A(n13774), .ZN(n13776) );
  NOR2_X1 U17284 ( .A1(n13775), .A2(n13965), .ZN(n14040) );
  NAND2_X1 U17285 ( .A1(n14031), .A2(n14054), .ZN(n14039) );
  OAI21_X1 U17286 ( .B1(n13776), .B2(n14040), .A(n14039), .ZN(n20070) );
  NOR2_X1 U17287 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n21986), .ZN(n19627) );
  INV_X1 U17288 ( .A(n20062), .ZN(n18240) );
  NOR2_X1 U17289 ( .A1(n20121), .A2(n18240), .ZN(n13778) );
  NAND2_X1 U17290 ( .A1(n18975), .A2(n20217), .ZN(n20098) );
  AOI22_X1 U17291 ( .A1(n20059), .A2(n13848), .B1(n13778), .B2(n18915), .ZN(
        n13779) );
  NAND3_X1 U17292 ( .A1(n13780), .A2(n13779), .A3(n13875), .ZN(n20073) );
  INV_X1 U17293 ( .A(n20073), .ZN(n20082) );
  INV_X1 U17294 ( .A(n20212), .ZN(n20105) );
  INV_X1 U17295 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n19616) );
  NAND3_X1 U17296 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n20198)
         );
  OAI22_X1 U17297 ( .A1(n20082), .A2(n20105), .B1(n19616), .B2(n20198), .ZN(
        n13781) );
  AOI21_X1 U17298 ( .B1(n14052), .B2(n20070), .A(n14055), .ZN(n13788) );
  NOR2_X1 U17299 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19604), .ZN(
        n14021) );
  INV_X1 U17300 ( .A(n14021), .ZN(n13782) );
  AOI22_X1 U17301 ( .A1(n20058), .A2(n14039), .B1(n14027), .B2(n13782), .ZN(
        n13783) );
  NOR2_X1 U17302 ( .A1(n13783), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n20071) );
  INV_X1 U17303 ( .A(n14040), .ZN(n13785) );
  INV_X2 U17304 ( .A(n18777), .ZN(n18646) );
  AOI21_X1 U17305 ( .B1(n13787), .B2(n13785), .A(n18646), .ZN(n18566) );
  AOI22_X1 U17306 ( .A1(n20071), .A2(n14052), .B1(n20095), .B2(n18566), .ZN(
        n13786) );
  OAI22_X1 U17307 ( .A1(n13788), .A2(n13787), .B1(n14055), .B2(n13786), .ZN(
        P3_U3285) );
  INV_X1 U17308 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n13791) );
  INV_X1 U17309 ( .A(n13789), .ZN(n21225) );
  AOI22_X1 U17310 ( .A1(n21225), .A2(P1_EAX_REG_28__SCAN_IN), .B1(n21254), 
        .B2(P1_UWORD_REG_12__SCAN_IN), .ZN(n13790) );
  OAI21_X1 U17311 ( .B1(n21237), .B2(n13791), .A(n13790), .ZN(P1_U2908) );
  NAND2_X1 U17312 ( .A1(n17995), .A2(n13792), .ZN(n13793) );
  NAND2_X1 U17313 ( .A1(n13793), .A2(n18092), .ZN(n13795) );
  OAI21_X1 U17314 ( .B1(n18025), .B2(n13795), .A(n14063), .ZN(n13799) );
  OAI21_X1 U17315 ( .B1(n14557), .B2(n11806), .A(n13796), .ZN(n13797) );
  NOR2_X1 U17316 ( .A1(n21733), .A2(n18095), .ZN(n14348) );
  AOI22_X1 U17317 ( .A1(n13800), .A2(n17997), .B1(P1_FLUSH_REG_SCAN_IN), .B2(
        n14348), .ZN(n18091) );
  OAI21_X1 U17318 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n11673), .A(n18091), 
        .ZN(n18088) );
  INV_X1 U17319 ( .A(n18088), .ZN(n21804) );
  INV_X1 U17320 ( .A(n13802), .ZN(n13804) );
  NOR2_X1 U17321 ( .A1(n13420), .A2(n11555), .ZN(n13803) );
  NAND3_X1 U17322 ( .A1(n13804), .A2(n13803), .A3(n9700), .ZN(n16273) );
  INV_X1 U17323 ( .A(n16273), .ZN(n15015) );
  OR2_X1 U17324 ( .A1(n13801), .A2(n15015), .ZN(n13814) );
  XNOR2_X1 U17325 ( .A(n13805), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13817) );
  OR2_X1 U17326 ( .A1(n14350), .A2(n13817), .ZN(n13811) );
  NAND2_X1 U17327 ( .A1(n13807), .A2(n13806), .ZN(n14356) );
  NAND2_X1 U17328 ( .A1(n14356), .A2(n13817), .ZN(n13810) );
  INV_X1 U17329 ( .A(n17995), .ZN(n15014) );
  XNOR2_X1 U17330 ( .A(n10694), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13808) );
  NAND2_X1 U17331 ( .A1(n15014), .A2(n13808), .ZN(n13809) );
  OAI211_X1 U17332 ( .C1(n16273), .C2(n13811), .A(n13810), .B(n13809), .ZN(
        n13812) );
  INV_X1 U17333 ( .A(n13812), .ZN(n13813) );
  NAND2_X1 U17334 ( .A1(n13814), .A2(n13813), .ZN(n14366) );
  NOR2_X1 U17335 ( .A1(n15370), .A2(n21912), .ZN(n16275) );
  OAI22_X1 U17336 ( .A1(n13815), .A2(n14243), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16274) );
  INV_X1 U17337 ( .A(n16274), .ZN(n13819) );
  INV_X1 U17338 ( .A(n21800), .ZN(n16277) );
  INV_X1 U17339 ( .A(n13817), .ZN(n13818) );
  AOI222_X1 U17340 ( .A1(n14366), .A2(n18087), .B1(n16275), .B2(n13819), .C1(
        n16277), .C2(n13818), .ZN(n13821) );
  NAND2_X1 U17341 ( .A1(n21804), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13820) );
  OAI21_X1 U17342 ( .B1(n21804), .B2(n13821), .A(n13820), .ZN(P1_U3472) );
  NAND2_X1 U17343 ( .A1(n14331), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13823) );
  AOI22_X1 U17344 ( .A1(n14277), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n21042), .B2(n21083), .ZN(n13825) );
  NOR2_X1 U17345 ( .A1(n17596), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13827) );
  OAI211_X1 U17346 ( .C1(n15209), .C2(n17566), .A(n9715), .B(n13827), .ZN(
        n13828) );
  INV_X1 U17347 ( .A(n13828), .ZN(n13829) );
  NAND2_X1 U17348 ( .A1(n13830), .A2(n9759), .ZN(n13831) );
  INV_X1 U17349 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n13832) );
  MUX2_X1 U17350 ( .A(n13833), .B(n13832), .S(n9713), .Z(n13834) );
  OAI21_X1 U17351 ( .B1(n21079), .B2(n16840), .A(n13834), .ZN(P2_U2887) );
  NAND2_X1 U17352 ( .A1(n14277), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13836) );
  NAND2_X1 U17353 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20521) );
  NAND2_X1 U17354 ( .A1(n22046), .A2(n21083), .ZN(n20678) );
  NAND2_X1 U17355 ( .A1(n20521), .A2(n20678), .ZN(n20618) );
  INV_X1 U17356 ( .A(n20618), .ZN(n20613) );
  NAND2_X1 U17357 ( .A1(n20613), .A2(n21042), .ZN(n20751) );
  NAND2_X1 U17358 ( .A1(n13836), .A2(n20751), .ZN(n13837) );
  INV_X1 U17359 ( .A(n16718), .ZN(n14712) );
  NOR2_X1 U17360 ( .A1(n14712), .A2(n9713), .ZN(n13838) );
  AOI21_X1 U17361 ( .B1(P2_EBX_REG_1__SCAN_IN), .B2(n9713), .A(n13838), .ZN(
        n13839) );
  OAI21_X1 U17362 ( .B1(n21045), .B2(n16840), .A(n13839), .ZN(P2_U2886) );
  INV_X1 U17363 ( .A(n14038), .ZN(n13841) );
  NOR2_X1 U17364 ( .A1(n13840), .A2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n19614) );
  NOR2_X1 U17365 ( .A1(n13841), .A2(n19614), .ZN(n20065) );
  NAND2_X1 U17366 ( .A1(n20065), .A2(n14052), .ZN(n13842) );
  INV_X1 U17367 ( .A(n14055), .ZN(n14049) );
  INV_X1 U17368 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n20069) );
  OAI22_X1 U17369 ( .A1(n14055), .A2(n13842), .B1(n14049), .B2(n20069), .ZN(
        P3_U3284) );
  NAND2_X1 U17370 ( .A1(n18552), .A2(n18568), .ZN(n13846) );
  NAND2_X1 U17371 ( .A1(n20233), .A2(n19628), .ZN(n18565) );
  INV_X1 U17372 ( .A(n14052), .ZN(n13967) );
  NAND3_X1 U17373 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n13967), .A3(
        n18552), .ZN(n13843) );
  OAI21_X1 U17374 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18565), .A(
        n13843), .ZN(n13845) );
  INV_X1 U17375 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n18815) );
  AOI21_X1 U17376 ( .B1(n18522), .B2(n18579), .A(n18815), .ZN(n13844) );
  AOI211_X1 U17377 ( .C1(n13846), .C2(P3_REIP_REG_0__SCAN_IN), .A(n13845), .B(
        n13844), .ZN(n13847) );
  INV_X1 U17378 ( .A(n13847), .ZN(P3_U2671) );
  INV_X1 U17379 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n18788) );
  INV_X1 U17380 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n18784) );
  NAND2_X1 U17381 ( .A1(n13850), .A2(P3_EBX_REG_9__SCAN_IN), .ZN(n18747) );
  NAND2_X1 U17382 ( .A1(n18747), .A2(n18808), .ZN(n18750) );
  NOR2_X1 U17383 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n13850), .ZN(n13870) );
  AOI22_X1 U17384 ( .A1(n9712), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n14457), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13861) );
  INV_X1 U17385 ( .A(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17696) );
  OAI22_X1 U17386 ( .A1(n18763), .A2(n17697), .B1(n14983), .B2(n17696), .ZN(
        n13853) );
  INV_X1 U17387 ( .A(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13851) );
  OAI22_X1 U17388 ( .A1(n18715), .A2(n13851), .B1(n17698), .B2(n17689), .ZN(
        n13852) );
  NOR2_X1 U17389 ( .A1(n13853), .A2(n13852), .ZN(n13860) );
  AOI22_X1 U17390 ( .A1(n9705), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n18652), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13859) );
  NAND2_X1 U17391 ( .A1(n18760), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n13857) );
  NAND2_X1 U17392 ( .A1(n17630), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n13856) );
  NAND2_X1 U17393 ( .A1(n18616), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n13855) );
  NAND2_X1 U17394 ( .A1(n17693), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n13854) );
  AND4_X1 U17395 ( .A1(n13857), .A2(n13856), .A3(n13855), .A4(n13854), .ZN(
        n13858) );
  NAND4_X1 U17396 ( .A1(n13861), .A2(n13860), .A3(n13859), .A4(n13858), .ZN(
        n13869) );
  NAND2_X1 U17397 ( .A1(n14951), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13867) );
  NAND2_X1 U17398 ( .A1(n14968), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n13866) );
  OR2_X1 U17399 ( .A1(n18775), .A2(n17690), .ZN(n13865) );
  INV_X1 U17400 ( .A(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13863) );
  OR2_X1 U17401 ( .A1(n18773), .A2(n13863), .ZN(n13864) );
  NAND4_X1 U17402 ( .A1(n13867), .A2(n13866), .A3(n13865), .A4(n13864), .ZN(
        n13868) );
  NOR2_X1 U17403 ( .A1(n13869), .A2(n13868), .ZN(n13887) );
  OAI22_X1 U17404 ( .A1(n18750), .A2(n13870), .B1(n13887), .B2(n18808), .ZN(
        P3_U2694) );
  NOR2_X1 U17405 ( .A1(n13871), .A2(n19650), .ZN(n13873) );
  AOI21_X1 U17406 ( .B1(n13874), .B2(n13873), .A(n13872), .ZN(n13877) );
  OAI21_X1 U17407 ( .B1(n13877), .B2(n13876), .A(n13875), .ZN(n13878) );
  NAND2_X1 U17408 ( .A1(n13881), .A2(n18606), .ZN(n18863) );
  INV_X1 U17409 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n18972) );
  OAI22_X1 U17410 ( .A1(n18863), .A2(P3_EAX_REG_0__SCAN_IN), .B1(n13881), .B2(
        n18972), .ZN(n13879) );
  AOI21_X1 U17411 ( .B1(n18911), .B2(n14174), .A(n13879), .ZN(n13880) );
  OAI21_X1 U17412 ( .B1(n18913), .B2(n19624), .A(n13880), .ZN(P3_U2735) );
  INV_X1 U17413 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n21987) );
  INV_X1 U17414 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n18969) );
  AOI211_X1 U17415 ( .C1(n13882), .C2(n18969), .A(n13908), .B(n18907), .ZN(
        n13883) );
  AOI21_X1 U17416 ( .B1(n18911), .B2(n14188), .A(n13883), .ZN(n13884) );
  OAI21_X1 U17417 ( .B1(n21987), .B2(n18913), .A(n13884), .ZN(P3_U2734) );
  INV_X1 U17418 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n19007) );
  NAND4_X1 U17419 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .A3(P3_EAX_REG_7__SCAN_IN), .A4(P3_EAX_REG_6__SCAN_IN), .ZN(n13885) );
  AND2_X1 U17420 ( .A1(n18903), .A2(n18606), .ZN(n17750) );
  AOI22_X1 U17421 ( .A1(n17750), .A2(P3_EAX_REG_8__SCAN_IN), .B1(
        P3_EAX_REG_9__SCAN_IN), .B2(n18902), .ZN(n13886) );
  INV_X1 U17422 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n18953) );
  OAI222_X1 U17423 ( .A1(n18913), .A2(n19007), .B1(n18883), .B2(n13887), .C1(
        n13886), .C2(n18896), .ZN(P3_U2726) );
  INV_X1 U17424 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n19637) );
  NAND2_X1 U17425 ( .A1(n9712), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n13891) );
  NAND2_X1 U17426 ( .A1(n14457), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n13890) );
  NAND2_X1 U17427 ( .A1(n9706), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n13889) );
  NAND2_X1 U17428 ( .A1(n18652), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n13888) );
  NAND2_X1 U17429 ( .A1(n18624), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n13895) );
  NAND2_X1 U17430 ( .A1(n18646), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13894) );
  INV_X1 U17431 ( .A(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14982) );
  OR2_X1 U17432 ( .A1(n18775), .A2(n14982), .ZN(n13893) );
  INV_X1 U17433 ( .A(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14984) );
  OR2_X1 U17434 ( .A1(n18773), .A2(n14984), .ZN(n13892) );
  INV_X1 U17435 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13896) );
  OAI22_X1 U17436 ( .A1(n18613), .A2(n13897), .B1(n14983), .B2(n13896), .ZN(
        n13899) );
  INV_X1 U17437 ( .A(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14978) );
  OAI22_X1 U17438 ( .A1(n18715), .A2(n14978), .B1(n18764), .B2(n14991), .ZN(
        n13898) );
  NOR2_X1 U17439 ( .A1(n13899), .A2(n13898), .ZN(n13905) );
  NAND2_X1 U17440 ( .A1(n14896), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n13903) );
  NAND2_X1 U17441 ( .A1(n18759), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n13902) );
  NAND2_X1 U17442 ( .A1(n17631), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n13901) );
  NAND2_X1 U17443 ( .A1(n17693), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n13900) );
  NAND4_X1 U17444 ( .A1(n13907), .A2(n13906), .A3(n13905), .A4(n13904), .ZN(
        n14195) );
  INV_X1 U17445 ( .A(n14195), .ZN(n14197) );
  INV_X1 U17446 ( .A(n13908), .ZN(n13909) );
  NOR2_X1 U17447 ( .A1(n19654), .A2(n13909), .ZN(n13929) );
  NAND2_X1 U17448 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n13930), .ZN(n13962) );
  INV_X1 U17449 ( .A(n13962), .ZN(n13911) );
  AOI21_X1 U17450 ( .B1(n18902), .B2(P3_EAX_REG_3__SCAN_IN), .A(n13930), .ZN(
        n13910) );
  OAI222_X1 U17451 ( .A1(n18913), .A2(n19637), .B1(n18883), .B2(n14197), .C1(
        n13911), .C2(n13910), .ZN(P3_U2732) );
  AOI22_X1 U17452 ( .A1(n13659), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18616), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13913) );
  INV_X2 U17453 ( .A(n17607), .ZN(n18759) );
  AOI22_X1 U17454 ( .A1(n18759), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n18692), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13912) );
  AND2_X1 U17455 ( .A1(n13913), .A2(n13912), .ZN(n13928) );
  NAND2_X1 U17456 ( .A1(n14457), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n13917) );
  NAND2_X1 U17457 ( .A1(n9706), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n13916) );
  NAND2_X1 U17458 ( .A1(n9712), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n13915) );
  NAND2_X1 U17459 ( .A1(n18652), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n13914) );
  NAND2_X1 U17460 ( .A1(n18646), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n13921) );
  NAND2_X1 U17461 ( .A1(n18624), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n13920) );
  INV_X1 U17462 ( .A(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n18730) );
  OR2_X1 U17463 ( .A1(n18775), .A2(n18730), .ZN(n13919) );
  INV_X1 U17464 ( .A(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n18728) );
  OR2_X1 U17465 ( .A1(n18773), .A2(n18728), .ZN(n13918) );
  INV_X1 U17466 ( .A(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18734) );
  NAND2_X1 U17467 ( .A1(n14896), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n13922) );
  OAI21_X1 U17468 ( .B1(n18734), .B2(n17695), .A(n13922), .ZN(n13924) );
  INV_X1 U17469 ( .A(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17680) );
  OAI22_X1 U17470 ( .A1(n18715), .A2(n17680), .B1(n18764), .B2(n18729), .ZN(
        n13923) );
  NOR2_X1 U17471 ( .A1(n13924), .A2(n13923), .ZN(n13925) );
  NAND4_X1 U17472 ( .A1(n13928), .A2(n13927), .A3(n13926), .A4(n13925), .ZN(
        n14189) );
  INV_X1 U17473 ( .A(n14189), .ZN(n14111) );
  INV_X1 U17474 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n19633) );
  AOI21_X1 U17475 ( .B1(n18902), .B2(P3_EAX_REG_2__SCAN_IN), .A(n13929), .ZN(
        n13931) );
  OAI222_X1 U17476 ( .A1(n18883), .A2(n14111), .B1(n18913), .B2(n19633), .C1(
        n13931), .C2(n13930), .ZN(P3_U2733) );
  NAND2_X1 U17477 ( .A1(n13932), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19214) );
  NAND2_X1 U17478 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n19615) );
  NAND2_X1 U17479 ( .A1(n21986), .A2(n19615), .ZN(n20211) );
  NAND2_X1 U17480 ( .A1(n20057), .A2(n20059), .ZN(n13934) );
  NAND2_X1 U17481 ( .A1(n20063), .A2(n19587), .ZN(n13933) );
  NAND3_X1 U17482 ( .A1(n18914), .A2(n19214), .A3(n19313), .ZN(n13942) );
  OR2_X2 U17483 ( .A1(n18244), .A2(n20217), .ZN(n19342) );
  INV_X1 U17484 ( .A(n13935), .ZN(n13937) );
  AND2_X1 U17485 ( .A1(n13937), .A2(n13936), .ZN(n13939) );
  INV_X1 U17486 ( .A(n13939), .ZN(n19609) );
  NOR2_X1 U17487 ( .A1(n19342), .A2(n19609), .ZN(n13941) );
  INV_X1 U17488 ( .A(n19556), .ZN(n19613) );
  INV_X1 U17489 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n13938) );
  OAI22_X1 U17490 ( .A1(n19334), .A2(n13939), .B1(n19613), .B2(n13938), .ZN(
        n13940) );
  AOI211_X1 U17491 ( .C1(n13942), .C2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n13941), .B(n13940), .ZN(n13943) );
  INV_X1 U17492 ( .A(n13943), .ZN(P3_U2830) );
  NAND2_X1 U17493 ( .A1(n9712), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n13947) );
  NAND2_X1 U17494 ( .A1(n14457), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n13946) );
  NAND2_X1 U17495 ( .A1(n9705), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n13945) );
  NAND2_X1 U17496 ( .A1(n18652), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n13944) );
  NAND2_X1 U17497 ( .A1(n18624), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n13951) );
  NAND2_X1 U17498 ( .A1(n18646), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n13950) );
  INV_X1 U17499 ( .A(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14892) );
  OR2_X1 U17500 ( .A1(n18775), .A2(n14892), .ZN(n13949) );
  INV_X1 U17501 ( .A(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14893) );
  OR2_X1 U17502 ( .A1(n18773), .A2(n14893), .ZN(n13948) );
  INV_X1 U17503 ( .A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n18695) );
  OAI22_X1 U17504 ( .A1(n18613), .A2(n18688), .B1(n14983), .B2(n18695), .ZN(
        n13953) );
  INV_X1 U17505 ( .A(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14467) );
  OAI22_X1 U17506 ( .A1(n18715), .A2(n14467), .B1(n18764), .B2(n14906), .ZN(
        n13952) );
  NOR2_X1 U17507 ( .A1(n13953), .A2(n13952), .ZN(n13959) );
  NAND2_X1 U17508 ( .A1(n14896), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n13957) );
  NAND2_X1 U17509 ( .A1(n18759), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n13956) );
  NAND2_X1 U17510 ( .A1(n17631), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n13955) );
  NAND2_X1 U17511 ( .A1(n17693), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n13954) );
  NAND4_X1 U17512 ( .A1(n13961), .A2(n13960), .A3(n13959), .A4(n13958), .ZN(
        n14208) );
  INV_X1 U17513 ( .A(n14208), .ZN(n14210) );
  INV_X1 U17514 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n19645) );
  INV_X1 U17515 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n18963) );
  NOR2_X1 U17516 ( .A1(n18963), .A2(n13962), .ZN(n18906) );
  AOI21_X1 U17517 ( .B1(n18902), .B2(P3_EAX_REG_5__SCAN_IN), .A(n18906), .ZN(
        n13963) );
  NAND2_X1 U17518 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n18906), .ZN(n17749) );
  INV_X1 U17519 ( .A(n17749), .ZN(n17752) );
  OAI222_X1 U17520 ( .A1(n18883), .A2(n14210), .B1(n18913), .B2(n19645), .C1(
        n13963), .C2(n17752), .ZN(P3_U2730) );
  NAND2_X1 U17521 ( .A1(n20095), .A2(n13965), .ZN(n13970) );
  NOR2_X1 U17522 ( .A1(n19526), .A2(n13964), .ZN(n14022) );
  MUX2_X1 U17523 ( .A(n19410), .B(n14022), .S(n13965), .Z(n20076) );
  NAND2_X1 U17524 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n19606), .ZN(n13966) );
  OAI211_X1 U17525 ( .C1(n20076), .C2(n13967), .A(n14049), .B(n13966), .ZN(
        n13968) );
  OAI21_X1 U17526 ( .B1(n14049), .B2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n13968), .ZN(n13969) );
  OAI21_X1 U17527 ( .B1(n14055), .B2(n13970), .A(n13969), .ZN(P3_U3290) );
  NAND3_X1 U17528 ( .A1(n18126), .A2(n13972), .A3(n13971), .ZN(n13982) );
  OR2_X1 U17529 ( .A1(n13974), .A2(n13973), .ZN(n13975) );
  NAND2_X1 U17530 ( .A1(n13976), .A2(n13975), .ZN(n14530) );
  AOI21_X1 U17531 ( .B1(n17505), .B2(n14530), .A(n13977), .ZN(n13981) );
  NAND2_X1 U17532 ( .A1(n18118), .A2(n13978), .ZN(n13979) );
  NAND4_X1 U17533 ( .A1(n13982), .A2(n13981), .A3(n13980), .A4(n13979), .ZN(
        n13983) );
  AOI21_X1 U17534 ( .B1(n14704), .B2(n18120), .A(n13983), .ZN(n13991) );
  INV_X1 U17535 ( .A(n13984), .ZN(n17363) );
  NAND2_X1 U17536 ( .A1(n17363), .A2(n13986), .ZN(n13989) );
  INV_X1 U17537 ( .A(n17361), .ZN(n13987) );
  AOI21_X1 U17538 ( .B1(n13987), .B2(n13986), .A(n13985), .ZN(n13988) );
  MUX2_X1 U17539 ( .A(n13989), .B(n13988), .S(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n13990) );
  NAND2_X1 U17540 ( .A1(n13991), .A2(n13990), .ZN(P2_U3044) );
  NAND2_X1 U17541 ( .A1(n14704), .A2(n14275), .ZN(n13995) );
  NAND2_X1 U17542 ( .A1(n20521), .A2(n21065), .ZN(n13993) );
  NAND2_X1 U17543 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20892) );
  INV_X1 U17544 ( .A(n20892), .ZN(n13992) );
  NAND2_X1 U17545 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13992), .ZN(
        n17558) );
  AND2_X1 U17546 ( .A1(n13993), .A2(n17558), .ZN(n14850) );
  AOI22_X1 U17547 ( .A1(n14277), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n21042), .B2(n14850), .ZN(n13994) );
  NAND2_X1 U17548 ( .A1(n14000), .A2(n13999), .ZN(n14004) );
  INV_X1 U17549 ( .A(n17539), .ZN(n14002) );
  NAND2_X1 U17550 ( .A1(n14002), .A2(n14001), .ZN(n14003) );
  XNOR2_X2 U17551 ( .A(n14283), .B(n14284), .ZN(n21058) );
  INV_X1 U17552 ( .A(n21058), .ZN(n16705) );
  MUX2_X1 U17553 ( .A(P2_EBX_REG_2__SCAN_IN), .B(n14704), .S(n16835), .Z(
        n14005) );
  AOI21_X1 U17554 ( .B1(n16705), .B2(n16830), .A(n14005), .ZN(n14006) );
  INV_X1 U17555 ( .A(n14006), .ZN(P2_U2885) );
  INV_X1 U17556 ( .A(n14007), .ZN(n14018) );
  NAND2_X1 U17557 ( .A1(n14008), .A2(n21912), .ZN(n14010) );
  NAND2_X1 U17558 ( .A1(n14010), .A2(n14009), .ZN(n15674) );
  INV_X1 U17559 ( .A(n15674), .ZN(n14012) );
  AOI21_X1 U17560 ( .B1(n21282), .B2(n14012), .A(n14011), .ZN(n14017) );
  AOI21_X1 U17561 ( .B1(n16198), .B2(n21912), .A(n10093), .ZN(n14244) );
  INV_X1 U17562 ( .A(n14244), .ZN(n14015) );
  NAND3_X1 U17563 ( .A1(n16203), .A2(n14013), .A3(n21912), .ZN(n14014) );
  OAI21_X1 U17564 ( .B1(n16089), .B2(n14015), .A(n14014), .ZN(n14016) );
  OAI211_X1 U17565 ( .C1(n14018), .C2(n21294), .A(n14017), .B(n14016), .ZN(
        P1_U3031) );
  INV_X1 U17566 ( .A(n14019), .ZN(n14020) );
  NAND2_X1 U17567 ( .A1(n14020), .A2(n14031), .ZN(n17605) );
  OAI22_X1 U17568 ( .A1(n14022), .A2(n17605), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n14021), .ZN(n20077) );
  INV_X1 U17569 ( .A(n20095), .ZN(n14050) );
  NOR2_X1 U17570 ( .A1(n18914), .A2(n19606), .ZN(n14047) );
  INV_X1 U17571 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n17775) );
  OAI22_X1 U17572 ( .A1(n17775), .A2(n19590), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14045) );
  NAND2_X1 U17573 ( .A1(n14047), .A2(n14045), .ZN(n14023) );
  OAI211_X1 U17574 ( .C1(n14050), .C2(n17605), .A(n14049), .B(n14023), .ZN(
        n14024) );
  AOI21_X1 U17575 ( .B1(n20077), .B2(n14052), .A(n14024), .ZN(n14025) );
  AOI21_X1 U17576 ( .B1(n14055), .B2(n14032), .A(n14025), .ZN(P3_U3289) );
  INV_X1 U17577 ( .A(n14026), .ZN(n14044) );
  NOR2_X1 U17578 ( .A1(n14028), .A2(n14027), .ZN(n14037) );
  OAI21_X1 U17579 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n14033), .A(
        n14029), .ZN(n14030) );
  AND2_X1 U17580 ( .A1(n14031), .A2(n14030), .ZN(n14035) );
  NOR2_X1 U17581 ( .A1(n14033), .A2(n14032), .ZN(n14034) );
  MUX2_X1 U17582 ( .A(n14035), .B(n14034), .S(n14054), .Z(n14036) );
  AOI21_X1 U17583 ( .B1(n14038), .B2(n14037), .A(n14036), .ZN(n14043) );
  INV_X1 U17584 ( .A(n14039), .ZN(n14041) );
  OR2_X1 U17585 ( .A1(n14041), .A2(n14040), .ZN(n18582) );
  NAND2_X1 U17586 ( .A1(n20058), .A2(n18582), .ZN(n14042) );
  OAI211_X1 U17587 ( .C1(n17966), .C2(n14044), .A(n14043), .B(n14042), .ZN(
        n20074) );
  INV_X1 U17588 ( .A(n14045), .ZN(n14046) );
  NAND2_X1 U17589 ( .A1(n14047), .A2(n14046), .ZN(n14048) );
  OAI211_X1 U17590 ( .C1(n14050), .C2(n18582), .A(n14049), .B(n14048), .ZN(
        n14051) );
  AOI21_X1 U17591 ( .B1(n20074), .B2(n14052), .A(n14051), .ZN(n14053) );
  AOI21_X1 U17592 ( .B1(n14055), .B2(n14054), .A(n14053), .ZN(P3_U3288) );
  OAI21_X1 U17593 ( .B1(n14058), .B2(n14057), .A(n14056), .ZN(n15673) );
  XOR2_X1 U17594 ( .A(n14059), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n14242) );
  NAND2_X1 U17595 ( .A1(n14242), .A2(n11864), .ZN(n14062) );
  INV_X1 U17596 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n21806) );
  NOR2_X1 U17597 ( .A1(n21291), .A2(n21806), .ZN(n14246) );
  NOR2_X1 U17598 ( .A1(n18056), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14060) );
  AOI211_X1 U17599 ( .C1(n18048), .C2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n14246), .B(n14060), .ZN(n14061) );
  OAI211_X1 U17600 ( .C1(n18057), .C2(n15673), .A(n14062), .B(n14061), .ZN(
        P1_U2998) );
  INV_X1 U17601 ( .A(n14064), .ZN(n14066) );
  NAND3_X1 U17602 ( .A1(n14066), .A2(n14238), .A3(n14065), .ZN(n14067) );
  INV_X1 U17603 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n14070) );
  OAI222_X1 U17604 ( .A1(n15681), .A2(n15702), .B1(n15709), .B2(n14070), .C1(
        n15674), .C2(n15704), .ZN(P1_U2872) );
  XNOR2_X1 U17605 ( .A(n14072), .B(n14071), .ZN(n14347) );
  NOR2_X1 U17606 ( .A1(n16203), .A2(n21912), .ZN(n14073) );
  MUX2_X1 U17607 ( .A(n16207), .B(n14073), .S(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n14080) );
  AND2_X1 U17608 ( .A1(n14075), .A2(n14074), .ZN(n14076) );
  OR2_X1 U17609 ( .A1(n14076), .A2(n9892), .ZN(n15655) );
  OAI21_X1 U17610 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n16252), .A(
        n16234), .ZN(n14077) );
  NOR2_X1 U17611 ( .A1(n16203), .A2(n16212), .ZN(n21280) );
  AOI21_X1 U17612 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n14077), .A(
        n21280), .ZN(n14078) );
  NAND2_X1 U17613 ( .A1(n18072), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n14344) );
  OAI211_X1 U17614 ( .C1(n21293), .C2(n15655), .A(n14078), .B(n14344), .ZN(
        n14079) );
  AOI21_X1 U17615 ( .B1(n14080), .B2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n14079), .ZN(n14081) );
  OAI21_X1 U17616 ( .B1(n14347), .B2(n21294), .A(n14081), .ZN(P1_U3029) );
  OR2_X1 U17617 ( .A1(n14083), .A2(n14082), .ZN(n14084) );
  AND2_X1 U17618 ( .A1(n14085), .A2(n14084), .ZN(n14525) );
  INV_X1 U17619 ( .A(n14525), .ZN(n21067) );
  OAI21_X1 U17620 ( .B1(n18115), .B2(n14087), .A(n14086), .ZN(n14090) );
  OAI22_X1 U17621 ( .A1(n17534), .A2(n14088), .B1(n14712), .B2(n17518), .ZN(
        n14089) );
  AOI211_X1 U17622 ( .C1(n17505), .C2(n21067), .A(n14090), .B(n14089), .ZN(
        n14093) );
  OAI211_X1 U17623 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n10205), .B(n14091), .ZN(n14092) );
  OAI211_X1 U17624 ( .C1(n17500), .C2(n14094), .A(n14093), .B(n14092), .ZN(
        P2_U3045) );
  INV_X1 U17625 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n18751) );
  NAND2_X1 U17626 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n14095), .ZN(n14472) );
  OAI21_X1 U17627 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n14095), .A(n14472), .ZN(
        n14110) );
  INV_X1 U17628 ( .A(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14096) );
  OAI22_X1 U17629 ( .A1(n9704), .A2(n14984), .B1(n17985), .B2(n14096), .ZN(
        n14098) );
  INV_X1 U17630 ( .A(n18652), .ZN(n18754) );
  OAI22_X1 U17631 ( .A1(n18755), .A2(n14982), .B1(n18754), .B2(n14991), .ZN(
        n14097) );
  NOR2_X1 U17632 ( .A1(n14098), .A2(n14097), .ZN(n14105) );
  AOI22_X1 U17633 ( .A1(n18759), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17693), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14104) );
  AOI22_X1 U17634 ( .A1(n18760), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17631), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14103) );
  INV_X1 U17635 ( .A(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17654) );
  OAI22_X1 U17636 ( .A1(n13896), .A2(n18613), .B1(n17695), .B2(n17654), .ZN(
        n14101) );
  INV_X1 U17637 ( .A(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14992) );
  OAI22_X1 U17638 ( .A1(n18715), .A2(n14992), .B1(n17698), .B2(n13897), .ZN(
        n14100) );
  NOR2_X1 U17639 ( .A1(n14101), .A2(n14100), .ZN(n14102) );
  AND4_X1 U17640 ( .A1(n14105), .A2(n14104), .A3(n14103), .A4(n14102), .ZN(
        n14108) );
  INV_X1 U17641 ( .A(n18775), .ZN(n18743) );
  AOI22_X1 U17642 ( .A1(n18743), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n18742), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14107) );
  AOI22_X1 U17643 ( .A1(n14951), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13784), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14106) );
  NAND3_X1 U17644 ( .A1(n14108), .A2(n14107), .A3(n14106), .ZN(n17744) );
  NAND2_X1 U17645 ( .A1(n18812), .A2(n17744), .ZN(n14109) );
  OAI21_X1 U17646 ( .B1(n14110), .B2(n18812), .A(n14109), .ZN(P3_U2692) );
  NAND2_X1 U17647 ( .A1(n14188), .A2(n14174), .ZN(n14173) );
  NAND2_X1 U17648 ( .A1(n14173), .A2(n14111), .ZN(n14171) );
  NAND2_X1 U17649 ( .A1(n14171), .A2(n14195), .ZN(n14170) );
  AOI22_X1 U17650 ( .A1(n14112), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n18760), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14117) );
  INV_X1 U17651 ( .A(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14996) );
  OAI22_X1 U17652 ( .A1(n18613), .A2(n14291), .B1(n18715), .B2(n14996), .ZN(
        n14113) );
  INV_X1 U17653 ( .A(n14113), .ZN(n14116) );
  AOI22_X1 U17654 ( .A1(n17631), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18717), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14115) );
  INV_X1 U17655 ( .A(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17625) );
  AOI22_X1 U17656 ( .A1(n18759), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n18692), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14114) );
  NAND2_X1 U17657 ( .A1(n18646), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n14121) );
  NAND2_X1 U17658 ( .A1(n18624), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n14120) );
  INV_X1 U17659 ( .A(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15000) );
  OR2_X1 U17660 ( .A1(n18773), .A2(n15000), .ZN(n14119) );
  INV_X1 U17661 ( .A(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14999) );
  OR2_X1 U17662 ( .A1(n18775), .A2(n14999), .ZN(n14118) );
  NAND2_X1 U17663 ( .A1(n14457), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n14125) );
  NAND2_X1 U17664 ( .A1(n9712), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n14124) );
  NAND2_X1 U17665 ( .A1(n9706), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n14123) );
  NAND2_X1 U17666 ( .A1(n18652), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n14122) );
  NAND2_X1 U17667 ( .A1(n14168), .A2(n14208), .ZN(n14167) );
  NAND2_X1 U17668 ( .A1(n9712), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n14132) );
  NAND2_X1 U17669 ( .A1(n14457), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n14131) );
  NAND2_X1 U17670 ( .A1(n9706), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n14130) );
  NAND2_X1 U17671 ( .A1(n18652), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n14129) );
  NAND2_X1 U17672 ( .A1(n18624), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n14136) );
  NAND2_X1 U17673 ( .A1(n18646), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n14135) );
  INV_X1 U17674 ( .A(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n18636) );
  OR2_X1 U17675 ( .A1(n18775), .A2(n18636), .ZN(n14134) );
  INV_X1 U17676 ( .A(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n18640) );
  OR2_X1 U17677 ( .A1(n18773), .A2(n18640), .ZN(n14133) );
  INV_X1 U17678 ( .A(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17615) );
  INV_X1 U17679 ( .A(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14479) );
  OAI22_X1 U17680 ( .A1(n18763), .A2(n17615), .B1(n14983), .B2(n14479), .ZN(
        n14138) );
  INV_X1 U17681 ( .A(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14487) );
  INV_X1 U17682 ( .A(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n18647) );
  OAI22_X1 U17683 ( .A1(n18715), .A2(n14487), .B1(n18764), .B2(n18647), .ZN(
        n14137) );
  NOR2_X1 U17684 ( .A1(n14138), .A2(n14137), .ZN(n14144) );
  NAND2_X1 U17685 ( .A1(n14896), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n14142) );
  NAND2_X1 U17686 ( .A1(n18759), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n14141) );
  INV_X1 U17687 ( .A(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17616) );
  NAND2_X1 U17688 ( .A1(n17631), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n14140) );
  NAND2_X1 U17689 ( .A1(n17693), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n14139) );
  NAND4_X1 U17690 ( .A1(n14146), .A2(n14145), .A3(n14144), .A4(n14143), .ZN(
        n14215) );
  NOR2_X1 U17691 ( .A1(n14167), .A2(n17755), .ZN(n14166) );
  NAND2_X1 U17692 ( .A1(n9712), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n14150) );
  NAND2_X1 U17693 ( .A1(n14457), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n14149) );
  NAND2_X1 U17694 ( .A1(n9705), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n14148) );
  NAND2_X1 U17695 ( .A1(n18652), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n14147) );
  NAND2_X1 U17696 ( .A1(n18624), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n14154) );
  NAND2_X1 U17697 ( .A1(n18646), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n14153) );
  INV_X1 U17698 ( .A(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n18612) );
  OR2_X1 U17699 ( .A1(n18775), .A2(n18612), .ZN(n14152) );
  INV_X1 U17700 ( .A(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n18618) );
  OR2_X1 U17701 ( .A1(n18773), .A2(n18618), .ZN(n14151) );
  INV_X1 U17702 ( .A(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14926) );
  INV_X1 U17703 ( .A(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14929) );
  OAI22_X1 U17704 ( .A1(n18763), .A2(n14926), .B1(n14983), .B2(n14929), .ZN(
        n14157) );
  INV_X1 U17705 ( .A(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14155) );
  INV_X1 U17706 ( .A(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n18626) );
  OAI22_X1 U17707 ( .A1(n18715), .A2(n14155), .B1(n18764), .B2(n18626), .ZN(
        n14156) );
  NOR2_X1 U17708 ( .A1(n14157), .A2(n14156), .ZN(n14163) );
  NAND2_X1 U17709 ( .A1(n18760), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n14161) );
  NAND2_X1 U17710 ( .A1(n17630), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n14160) );
  NAND2_X1 U17711 ( .A1(n17631), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n14159) );
  NAND2_X1 U17712 ( .A1(n17693), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n14158) );
  AND2_X1 U17713 ( .A1(n14166), .A2(n17942), .ZN(n14401) );
  XNOR2_X1 U17714 ( .A(n14166), .B(n17778), .ZN(n19265) );
  XNOR2_X1 U17715 ( .A(n14167), .B(n14215), .ZN(n14182) );
  XNOR2_X1 U17716 ( .A(n14168), .B(n14210), .ZN(n14169) );
  NAND2_X1 U17717 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n14169), .ZN(
        n14181) );
  XOR2_X1 U17718 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n14169), .Z(
        n19291) );
  INV_X1 U17719 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19569) );
  INV_X1 U17720 ( .A(n14206), .ZN(n18910) );
  XNOR2_X1 U17721 ( .A(n14170), .B(n18910), .ZN(n19298) );
  XNOR2_X1 U17722 ( .A(n14171), .B(n14197), .ZN(n14172) );
  NAND2_X1 U17723 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n14172), .ZN(
        n14179) );
  XOR2_X1 U17724 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n14172), .Z(
        n19317) );
  XNOR2_X1 U17725 ( .A(n14173), .B(n14189), .ZN(n14177) );
  INV_X1 U17726 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19592) );
  OR2_X1 U17727 ( .A1(n14177), .A2(n19592), .ZN(n14178) );
  INV_X1 U17728 ( .A(n14188), .ZN(n14190) );
  AOI21_X1 U17729 ( .B1(n14188), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14175) );
  MUX2_X1 U17730 ( .A(n14175), .B(n14188), .S(n14174), .Z(n14176) );
  AOI21_X1 U17731 ( .B1(n14190), .B2(n19590), .A(n14176), .ZN(n19333) );
  XNOR2_X1 U17732 ( .A(n14177), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n19332) );
  NAND2_X1 U17733 ( .A1(n19317), .A2(n19316), .ZN(n19315) );
  NAND2_X1 U17734 ( .A1(n14179), .A2(n19315), .ZN(n19299) );
  NAND2_X1 U17735 ( .A1(n19298), .A2(n19299), .ZN(n19297) );
  NOR2_X1 U17736 ( .A1(n19298), .A2(n19299), .ZN(n14180) );
  NAND2_X1 U17737 ( .A1(n19291), .A2(n19290), .ZN(n19289) );
  NAND2_X1 U17738 ( .A1(n14182), .A2(n14183), .ZN(n14184) );
  INV_X1 U17739 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n22078) );
  NOR2_X2 U17740 ( .A1(n19263), .A2(n22078), .ZN(n14400) );
  NAND2_X1 U17741 ( .A1(n14401), .A2(n14186), .ZN(n14185) );
  OAI21_X1 U17742 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n14187), .A(
        n14402), .ZN(n17889) );
  OR2_X1 U17743 ( .A1(n19605), .A2(n17942), .ZN(n19504) );
  OAI21_X1 U17744 ( .B1(n14189), .B2(n14188), .A(n14198), .ZN(n14193) );
  XNOR2_X1 U17745 ( .A(n14193), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n19326) );
  NAND2_X1 U17746 ( .A1(n14190), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14191) );
  NAND2_X1 U17747 ( .A1(n14192), .A2(n14191), .ZN(n19325) );
  OR2_X1 U17748 ( .A1(n14193), .A2(n19592), .ZN(n14194) );
  INV_X1 U17749 ( .A(n14198), .ZN(n14196) );
  NAND2_X1 U17750 ( .A1(n14198), .A2(n14197), .ZN(n14199) );
  NAND2_X1 U17751 ( .A1(n14207), .A2(n14199), .ZN(n14200) );
  XNOR2_X1 U17752 ( .A(n14207), .B(n14206), .ZN(n14203) );
  XNOR2_X1 U17753 ( .A(n14203), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19303) );
  INV_X1 U17754 ( .A(n14203), .ZN(n14204) );
  NAND2_X1 U17755 ( .A1(n14204), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n14205) );
  INV_X1 U17756 ( .A(n14209), .ZN(n14211) );
  NAND2_X1 U17757 ( .A1(n14211), .A2(n14210), .ZN(n14212) );
  NAND2_X1 U17758 ( .A1(n14218), .A2(n14212), .ZN(n19286) );
  XNOR2_X1 U17759 ( .A(n14218), .B(n14215), .ZN(n14216) );
  XNOR2_X1 U17760 ( .A(n14216), .B(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n19273) );
  NAND2_X1 U17761 ( .A1(n14216), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14217) );
  NAND2_X1 U17762 ( .A1(n14219), .A2(n17778), .ZN(n14220) );
  NAND2_X1 U17763 ( .A1(n19196), .A2(n14220), .ZN(n14221) );
  NAND2_X1 U17764 ( .A1(n19268), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n19267) );
  INV_X1 U17765 ( .A(n14221), .ZN(n14222) );
  NAND2_X1 U17766 ( .A1(n14223), .A2(n14222), .ZN(n14224) );
  INV_X1 U17767 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n19546) );
  NAND3_X1 U17768 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19448) );
  INV_X1 U17769 ( .A(n19448), .ZN(n14226) );
  OAI21_X1 U17770 ( .B1(n19606), .B2(n19590), .A(n19592), .ZN(n19584) );
  NOR2_X1 U17771 ( .A1(n19592), .A2(n19590), .ZN(n19562) );
  OAI21_X1 U17772 ( .B1(n17966), .B2(n19606), .A(n19410), .ZN(n19593) );
  AOI22_X1 U17773 ( .A1(n20058), .A2(n19584), .B1(n19562), .B2(n19593), .ZN(
        n19576) );
  NOR2_X1 U17774 ( .A1(n19576), .A2(n19575), .ZN(n19570) );
  NAND2_X1 U17775 ( .A1(n14226), .A2(n19570), .ZN(n19547) );
  NOR3_X1 U17776 ( .A1(n22078), .A2(n19546), .A3(n19547), .ZN(n14405) );
  INV_X1 U17777 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n14410) );
  NAND2_X1 U17778 ( .A1(n14226), .A2(n19584), .ZN(n14413) );
  INV_X1 U17779 ( .A(n14413), .ZN(n14228) );
  NAND2_X1 U17780 ( .A1(n14226), .A2(n19562), .ZN(n14411) );
  NOR2_X1 U17781 ( .A1(n17966), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n19591) );
  NOR2_X1 U17782 ( .A1(n19526), .A2(n19604), .ZN(n19561) );
  INV_X1 U17783 ( .A(n19561), .ZN(n19589) );
  OAI21_X1 U17784 ( .B1(n14411), .B2(n19591), .A(n19589), .ZN(n14227) );
  OAI21_X1 U17785 ( .B1(n19560), .B2(n14228), .A(n14227), .ZN(n19544) );
  AOI211_X1 U17786 ( .C1(n19477), .C2(n19546), .A(n22078), .B(n19544), .ZN(
        n14229) );
  INV_X1 U17787 ( .A(n14229), .ZN(n19535) );
  AOI21_X1 U17788 ( .B1(n19497), .B2(n19535), .A(n19602), .ZN(n14230) );
  NAND2_X1 U17789 ( .A1(n19556), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n17881) );
  OAI21_X1 U17790 ( .B1(n14230), .B2(n14410), .A(n17881), .ZN(n14231) );
  AOI21_X1 U17791 ( .B1(n14405), .B2(n14410), .A(n14231), .ZN(n14234) );
  NAND2_X1 U17792 ( .A1(n17878), .A2(n19196), .ZN(n14232) );
  NAND2_X1 U17793 ( .A1(n17844), .A2(n14232), .ZN(n17886) );
  NAND2_X1 U17794 ( .A1(n17886), .A2(n19530), .ZN(n14233) );
  OAI211_X1 U17795 ( .C1(n19504), .C2(n17878), .A(n14234), .B(n14233), .ZN(
        n14235) );
  INV_X1 U17796 ( .A(n14235), .ZN(n14236) );
  OAI21_X1 U17797 ( .B1(n17889), .B2(n10311), .A(n14236), .ZN(P3_U2854) );
  OAI21_X1 U17798 ( .B1(n14239), .B2(n14238), .A(n14237), .ZN(n15671) );
  INV_X1 U17799 ( .A(n15671), .ZN(n14241) );
  INV_X1 U17800 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n14240) );
  OAI222_X1 U17801 ( .A1(n15673), .A2(n15702), .B1(n15704), .B2(n14241), .C1(
        n15709), .C2(n14240), .ZN(P1_U2871) );
  INV_X1 U17802 ( .A(n14242), .ZN(n14250) );
  NOR2_X1 U17803 ( .A1(n14244), .A2(n14243), .ZN(n14245) );
  AOI211_X1 U17804 ( .C1(n21282), .C2(n15671), .A(n14246), .B(n14245), .ZN(
        n14249) );
  OR3_X1 U17805 ( .A1(n16137), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n14247), .ZN(n14248) );
  OAI211_X1 U17806 ( .C1(n14250), .C2(n21294), .A(n14249), .B(n14248), .ZN(
        P1_U3030) );
  AND2_X1 U17807 ( .A1(n21825), .A2(n21822), .ZN(n14251) );
  INV_X1 U17808 ( .A(n14330), .ZN(n21274) );
  AOI22_X1 U17809 ( .A1(n9699), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n21274), .ZN(n14255) );
  NAND2_X1 U17810 ( .A1(n14547), .A2(DATAI_3_), .ZN(n14253) );
  NAND2_X1 U17811 ( .A1(n15020), .A2(BUF1_REG_3__SCAN_IN), .ZN(n14252) );
  AND2_X1 U17812 ( .A1(n14253), .A2(n14252), .ZN(n15757) );
  INV_X1 U17813 ( .A(n15757), .ZN(n14254) );
  NAND2_X1 U17814 ( .A1(n21260), .A2(n14254), .ZN(n14661) );
  NAND2_X1 U17815 ( .A1(n14255), .A2(n14661), .ZN(P1_U2940) );
  AOI22_X1 U17816 ( .A1(n9699), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n21274), .ZN(n14258) );
  INV_X1 U17817 ( .A(DATAI_2_), .ZN(n14257) );
  NAND2_X1 U17818 ( .A1(n15020), .A2(BUF1_REG_2__SCAN_IN), .ZN(n14256) );
  OAI21_X1 U17819 ( .B1(n15020), .B2(n14257), .A(n14256), .ZN(n15762) );
  NAND2_X1 U17820 ( .A1(n21260), .A2(n15762), .ZN(n14663) );
  NAND2_X1 U17821 ( .A1(n14258), .A2(n14663), .ZN(P1_U2939) );
  AOI22_X1 U17822 ( .A1(n9699), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n21274), .ZN(n14262) );
  INV_X1 U17823 ( .A(DATAI_4_), .ZN(n14260) );
  MUX2_X1 U17824 ( .A(n14260), .B(n14259), .S(n15020), .Z(n15753) );
  INV_X1 U17825 ( .A(n15753), .ZN(n14261) );
  NAND2_X1 U17826 ( .A1(n21260), .A2(n14261), .ZN(n14678) );
  NAND2_X1 U17827 ( .A1(n14262), .A2(n14678), .ZN(P1_U2941) );
  AOI22_X1 U17828 ( .A1(n9699), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n21274), .ZN(n14266) );
  NAND2_X1 U17829 ( .A1(n14547), .A2(DATAI_1_), .ZN(n14264) );
  NAND2_X1 U17830 ( .A1(n15020), .A2(BUF1_REG_1__SCAN_IN), .ZN(n14263) );
  AND2_X1 U17831 ( .A1(n14264), .A2(n14263), .ZN(n15767) );
  INV_X1 U17832 ( .A(n15767), .ZN(n14265) );
  NAND2_X1 U17833 ( .A1(n21260), .A2(n14265), .ZN(n14659) );
  NAND2_X1 U17834 ( .A1(n14266), .A2(n14659), .ZN(P1_U2938) );
  AOI22_X1 U17835 ( .A1(n9699), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n21274), .ZN(n14270) );
  NAND2_X1 U17836 ( .A1(n14547), .A2(DATAI_7_), .ZN(n14268) );
  NAND2_X1 U17837 ( .A1(n15020), .A2(BUF1_REG_7__SCAN_IN), .ZN(n14267) );
  AND2_X1 U17838 ( .A1(n14268), .A2(n14267), .ZN(n15739) );
  INV_X1 U17839 ( .A(n15739), .ZN(n14269) );
  NAND2_X1 U17840 ( .A1(n21260), .A2(n14269), .ZN(n14682) );
  NAND2_X1 U17841 ( .A1(n14270), .A2(n14682), .ZN(P1_U2959) );
  INV_X1 U17842 ( .A(P1_UWORD_REG_12__SCAN_IN), .ZN(n22052) );
  INV_X1 U17843 ( .A(DATAI_12_), .ZN(n14272) );
  MUX2_X1 U17844 ( .A(n14272), .B(n14271), .S(n15020), .Z(n15789) );
  INV_X1 U17845 ( .A(n15789), .ZN(n14273) );
  NAND2_X1 U17846 ( .A1(n21260), .A2(n14273), .ZN(n21268) );
  NAND2_X1 U17847 ( .A1(n9699), .A2(P1_EAX_REG_28__SCAN_IN), .ZN(n14274) );
  OAI211_X1 U17848 ( .C1(n14330), .C2(n22052), .A(n21268), .B(n14274), .ZN(
        P1_U2949) );
  NAND2_X1 U17849 ( .A1(n17530), .A2(n14275), .ZN(n14279) );
  INV_X1 U17850 ( .A(n20521), .ZN(n20780) );
  NAND2_X1 U17851 ( .A1(n21054), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20617) );
  INV_X1 U17852 ( .A(n20617), .ZN(n20612) );
  NAND2_X1 U17853 ( .A1(n20780), .A2(n20612), .ZN(n20649) );
  NAND2_X1 U17854 ( .A1(n17558), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14276) );
  NAND2_X1 U17855 ( .A1(n20649), .A2(n14276), .ZN(n20545) );
  AOI22_X1 U17856 ( .A1(n14277), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n21042), .B2(n20545), .ZN(n14278) );
  NAND2_X1 U17857 ( .A1(n14334), .A2(n14280), .ZN(n14435) );
  AND2_X4 U17858 ( .A1(n14333), .A2(n14286), .ZN(n21047) );
  MUX2_X1 U17859 ( .A(n12259), .B(n14288), .S(n16835), .Z(n14289) );
  OAI21_X1 U17860 ( .B1(n20713), .B2(n16840), .A(n14289), .ZN(P2_U2884) );
  INV_X1 U17861 ( .A(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17626) );
  OAI22_X1 U17862 ( .A1(n18613), .A2(n17626), .B1(n14983), .B2(n17625), .ZN(
        n14290) );
  INV_X1 U17863 ( .A(n14290), .ZN(n14297) );
  AOI22_X1 U17864 ( .A1(n18760), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17631), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14296) );
  AOI22_X1 U17865 ( .A1(n18759), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12013), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14295) );
  INV_X1 U17866 ( .A(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14292) );
  OAI22_X1 U17867 ( .A1(n18715), .A2(n14292), .B1(n17698), .B2(n14291), .ZN(
        n14293) );
  INV_X1 U17868 ( .A(n14293), .ZN(n14294) );
  AND4_X1 U17869 ( .A1(n14297), .A2(n14296), .A3(n14295), .A4(n14294), .ZN(
        n14305) );
  AOI22_X1 U17870 ( .A1(n18743), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18742), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14304) );
  AOI22_X1 U17871 ( .A1(n14951), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n14968), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14303) );
  NAND2_X1 U17872 ( .A1(n9712), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n14301) );
  NAND2_X1 U17873 ( .A1(n14457), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n14300) );
  NAND2_X1 U17874 ( .A1(n9706), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n14299) );
  NAND2_X1 U17875 ( .A1(n18652), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n14298) );
  AND4_X1 U17876 ( .A1(n14301), .A2(n14300), .A3(n14299), .A4(n14298), .ZN(
        n14302) );
  AND4_X1 U17877 ( .A1(n14305), .A2(n14304), .A3(n14303), .A4(n14302), .ZN(
        n17743) );
  NOR2_X1 U17878 ( .A1(n14472), .A2(n19654), .ZN(n14491) );
  INV_X1 U17879 ( .A(n14491), .ZN(n14306) );
  NAND3_X1 U17880 ( .A1(n14306), .A2(P3_EBX_REG_12__SCAN_IN), .A3(n18808), 
        .ZN(n14308) );
  INV_X1 U17881 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n14471) );
  NAND2_X1 U17882 ( .A1(n14491), .A2(n14471), .ZN(n14307) );
  OAI211_X1 U17883 ( .C1(n17743), .C2(n18808), .A(n14308), .B(n14307), .ZN(
        P3_U2691) );
  NAND2_X1 U17884 ( .A1(n21270), .A2(P1_UWORD_REG_8__SCAN_IN), .ZN(n14312) );
  INV_X1 U17885 ( .A(DATAI_8_), .ZN(n14310) );
  MUX2_X1 U17886 ( .A(n14310), .B(n14309), .S(n15020), .Z(n15735) );
  INV_X1 U17887 ( .A(n15735), .ZN(n14311) );
  NAND2_X1 U17888 ( .A1(n21260), .A2(n14311), .ZN(n14317) );
  OAI211_X1 U17889 ( .C1(n14658), .C2(n15734), .A(n14312), .B(n14317), .ZN(
        P1_U2945) );
  NAND2_X1 U17890 ( .A1(n21274), .A2(P1_UWORD_REG_10__SCAN_IN), .ZN(n14315) );
  INV_X1 U17891 ( .A(DATAI_10_), .ZN(n14313) );
  MUX2_X1 U17892 ( .A(n14313), .B(n18180), .S(n15020), .Z(n15723) );
  INV_X1 U17893 ( .A(n15723), .ZN(n14314) );
  NAND2_X1 U17894 ( .A1(n21260), .A2(n14314), .ZN(n21264) );
  OAI211_X1 U17895 ( .C1(n14658), .C2(n14316), .A(n14315), .B(n21264), .ZN(
        P1_U2947) );
  INV_X1 U17896 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n21241) );
  NAND2_X1 U17897 ( .A1(n21274), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n14318) );
  OAI211_X1 U17898 ( .C1(n14658), .C2(n21241), .A(n14318), .B(n14317), .ZN(
        P1_U2960) );
  NAND2_X1 U17899 ( .A1(n21274), .A2(P1_UWORD_REG_9__SCAN_IN), .ZN(n14322) );
  INV_X1 U17900 ( .A(DATAI_9_), .ZN(n14320) );
  MUX2_X1 U17901 ( .A(n14320), .B(n14319), .S(n15020), .Z(n15729) );
  INV_X1 U17902 ( .A(n15729), .ZN(n14321) );
  NAND2_X1 U17903 ( .A1(n21260), .A2(n14321), .ZN(n21262) );
  OAI211_X1 U17904 ( .C1(n14658), .C2(n15728), .A(n14322), .B(n21262), .ZN(
        P1_U2946) );
  NAND2_X1 U17905 ( .A1(n21274), .A2(P1_UWORD_REG_11__SCAN_IN), .ZN(n14325) );
  INV_X1 U17906 ( .A(DATAI_11_), .ZN(n14324) );
  NAND2_X1 U17907 ( .A1(n15020), .A2(BUF1_REG_11__SCAN_IN), .ZN(n14323) );
  OAI21_X1 U17908 ( .B1(n15020), .B2(n14324), .A(n14323), .ZN(n15791) );
  NAND2_X1 U17909 ( .A1(n21260), .A2(n15791), .ZN(n21266) );
  OAI211_X1 U17910 ( .C1(n14658), .C2(n14326), .A(n14325), .B(n21266), .ZN(
        P1_U2948) );
  INV_X1 U17911 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n21229) );
  INV_X1 U17912 ( .A(n21260), .ZN(n14329) );
  INV_X1 U17913 ( .A(DATAI_15_), .ZN(n14328) );
  MUX2_X1 U17914 ( .A(n14328), .B(n14327), .S(n15020), .Z(n15780) );
  OAI222_X1 U17915 ( .A1(n14658), .A2(n21228), .B1(n14330), .B2(n21229), .C1(
        n14329), .C2(n15780), .ZN(P1_U2967) );
  NAND2_X1 U17916 ( .A1(n14331), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n14332) );
  AND2_X1 U17917 ( .A1(n14334), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n14335) );
  AND2_X1 U17918 ( .A1(n15275), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n14433) );
  XNOR2_X1 U17919 ( .A(n14654), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14339) );
  AOI21_X1 U17920 ( .B1(n14337), .B2(n14336), .A(n9883), .ZN(n20328) );
  INV_X1 U17921 ( .A(n20328), .ZN(n17507) );
  MUX2_X1 U17922 ( .A(n22065), .B(n17507), .S(n16835), .Z(n14338) );
  OAI21_X1 U17923 ( .B1(n14339), .B2(n16840), .A(n14338), .ZN(P2_U2882) );
  NAND2_X1 U17924 ( .A1(n14341), .A2(n14340), .ZN(n14342) );
  AOI21_X1 U17925 ( .B1(n14056), .B2(n14342), .A(n10656), .ZN(n14445) );
  NAND2_X1 U17926 ( .A1(n18048), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14343) );
  OAI211_X1 U17927 ( .C1(n18056), .C2(n15662), .A(n14344), .B(n14343), .ZN(
        n14345) );
  AOI21_X1 U17928 ( .B1(n14445), .B2(n18052), .A(n14345), .ZN(n14346) );
  OAI21_X1 U17929 ( .B1(n21105), .B2(n14347), .A(n14346), .ZN(P1_U2997) );
  INV_X1 U17930 ( .A(n14348), .ZN(n18099) );
  NAND2_X1 U17931 ( .A1(n21310), .A2(n16273), .ZN(n14365) );
  INV_X1 U17932 ( .A(n10700), .ZN(n14353) );
  OAI211_X1 U17933 ( .C1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C2(n13805), .A(
        n10877), .B(n14353), .ZN(n21801) );
  OR2_X1 U17934 ( .A1(n14350), .A2(n21801), .ZN(n14362) );
  INV_X1 U17935 ( .A(n14351), .ZN(n14355) );
  MUX2_X1 U17936 ( .A(n14353), .B(n14352), .S(n13805), .Z(n14354) );
  NAND3_X1 U17937 ( .A1(n14356), .A2(n14355), .A3(n14354), .ZN(n14361) );
  NAND2_X1 U17938 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14358) );
  INV_X1 U17939 ( .A(n14358), .ZN(n14357) );
  MUX2_X1 U17940 ( .A(n14358), .B(n14357), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n14359) );
  OR2_X1 U17941 ( .A1(n17995), .A2(n14359), .ZN(n14360) );
  OAI211_X1 U17942 ( .C1(n16273), .C2(n14362), .A(n14361), .B(n14360), .ZN(
        n14363) );
  INV_X1 U17943 ( .A(n14363), .ZN(n14364) );
  NAND2_X1 U17944 ( .A1(n14365), .A2(n14364), .ZN(n21799) );
  MUX2_X1 U17945 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n21799), .S(
        n17997), .Z(n18006) );
  NAND2_X1 U17946 ( .A1(n18006), .A2(n15370), .ZN(n14369) );
  NOR2_X1 U17947 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n15370), .ZN(n14373) );
  NAND2_X1 U17948 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n14373), .ZN(
        n14368) );
  MUX2_X1 U17949 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14366), .S(
        n17997), .Z(n18005) );
  AOI22_X1 U17950 ( .A1(n14373), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n18005), .B2(n15370), .ZN(n14367) );
  AOI21_X1 U17951 ( .B1(n14369), .B2(n14368), .A(n14367), .ZN(n18018) );
  INV_X1 U17952 ( .A(n10699), .ZN(n14370) );
  AND2_X1 U17953 ( .A1(n18018), .A2(n14370), .ZN(n14377) );
  INV_X1 U17954 ( .A(n14540), .ZN(n14753) );
  XNOR2_X1 U17955 ( .A(n14371), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n21183) );
  NAND2_X1 U17956 ( .A1(n21183), .A2(n18086), .ZN(n14372) );
  MUX2_X1 U17957 ( .A(n18089), .B(n14372), .S(n17997), .Z(n14375) );
  NAND2_X1 U17958 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n14373), .ZN(
        n14374) );
  OAI21_X1 U17959 ( .B1(n14375), .B2(P1_STATE2_REG_1__SCAN_IN), .A(n14374), 
        .ZN(n18016) );
  NOR3_X1 U17960 ( .A1(n14377), .A2(n18016), .A3(P1_FLUSH_REG_SCAN_IN), .ZN(
        n14376) );
  INV_X1 U17961 ( .A(n18095), .ZN(n14378) );
  OAI21_X1 U17962 ( .B1(n18099), .B2(n14376), .A(n14757), .ZN(n21302) );
  INV_X1 U17963 ( .A(n14377), .ZN(n14380) );
  INV_X1 U17964 ( .A(n18016), .ZN(n14379) );
  NAND3_X1 U17965 ( .A1(n14380), .A2(n14379), .A3(n14378), .ZN(n18031) );
  INV_X1 U17966 ( .A(n18031), .ZN(n14382) );
  INV_X1 U17967 ( .A(n14542), .ZN(n15676) );
  NAND2_X1 U17968 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n11673), .ZN(n14394) );
  INV_X1 U17969 ( .A(n14394), .ZN(n16268) );
  OAI22_X1 U17970 ( .A1(n14752), .A2(n21667), .B1(n15676), .B2(n16268), .ZN(
        n14381) );
  OAI21_X1 U17971 ( .B1(n14382), .B2(n14381), .A(n21302), .ZN(n14383) );
  OAI21_X1 U17972 ( .B1(n21302), .B2(n21561), .A(n14383), .ZN(P1_U3478) );
  NOR2_X1 U17973 ( .A1(n13801), .A2(n16268), .ZN(n14387) );
  INV_X1 U17974 ( .A(n9707), .ZN(n14385) );
  NOR3_X1 U17975 ( .A1(n14385), .A2(n21528), .A3(n21667), .ZN(n14613) );
  AOI21_X1 U17976 ( .B1(n9707), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n21667), 
        .ZN(n21672) );
  OAI21_X1 U17977 ( .B1(n14387), .B2(n14386), .A(n21302), .ZN(n14388) );
  OAI21_X1 U17978 ( .B1(n21302), .B2(n21306), .A(n14388), .ZN(P1_U3476) );
  INV_X1 U17979 ( .A(n21302), .ZN(n14399) );
  NOR2_X1 U17980 ( .A1(n9702), .A2(n14389), .ZN(n14390) );
  MUX2_X1 U17981 ( .A(n21673), .B(n21455), .S(n9707), .Z(n14393) );
  NAND2_X1 U17982 ( .A1(n14393), .A2(n21529), .ZN(n14396) );
  NOR2_X1 U17983 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n21667), .ZN(n21484) );
  AOI222_X1 U17984 ( .A1(n14396), .A2(n14395), .B1(n10046), .B2(n21484), .C1(
        n21310), .C2(n14394), .ZN(n14398) );
  NAND2_X1 U17985 ( .A1(n14399), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14397) );
  OAI21_X1 U17986 ( .B1(n14399), .B2(n14398), .A(n14397), .ZN(P1_U3475) );
  NAND2_X1 U17987 ( .A1(n14401), .A2(n14400), .ZN(n14403) );
  INV_X1 U17988 ( .A(n19504), .ZN(n14404) );
  AOI222_X1 U17989 ( .A1(n19188), .A2(n19610), .B1(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n14405), .C1(n19209), .C2(
        n14404), .ZN(n19519) );
  OR2_X1 U17990 ( .A1(n19198), .A2(n10323), .ZN(n17977) );
  INV_X1 U17991 ( .A(n17977), .ZN(n17975) );
  NOR2_X1 U17992 ( .A1(n17856), .A2(n19196), .ZN(n19200) );
  NOR2_X1 U17993 ( .A1(n17975), .A2(n19200), .ZN(n14406) );
  INV_X1 U17994 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17974) );
  XOR2_X1 U17995 ( .A(n14406), .B(n17974), .Z(n17875) );
  INV_X1 U17996 ( .A(n17875), .ZN(n14408) );
  INV_X1 U17997 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n14407) );
  OAI22_X1 U17998 ( .A1(n19505), .A2(n14408), .B1(n19613), .B2(n14407), .ZN(
        n14409) );
  INV_X1 U17999 ( .A(n14409), .ZN(n14417) );
  NOR3_X1 U18000 ( .A1(n22078), .A2(n19546), .A3(n14410), .ZN(n19449) );
  INV_X1 U18001 ( .A(n19449), .ZN(n14412) );
  NOR2_X1 U18002 ( .A1(n14412), .A2(n14411), .ZN(n19495) );
  INV_X1 U18003 ( .A(n19591), .ZN(n19452) );
  OAI21_X1 U18004 ( .B1(n19495), .B2(n19561), .A(n19452), .ZN(n14415) );
  INV_X1 U18005 ( .A(n19188), .ZN(n17857) );
  NOR2_X1 U18006 ( .A1(n14413), .A2(n14412), .ZN(n17890) );
  NOR2_X1 U18007 ( .A1(n17890), .A2(n19560), .ZN(n19473) );
  OR2_X1 U18008 ( .A1(n20064), .A2(n17942), .ZN(n19401) );
  NOR2_X1 U18009 ( .A1(n19209), .A2(n19401), .ZN(n14414) );
  AOI211_X1 U18010 ( .C1(n17857), .C2(n20057), .A(n19473), .B(n14414), .ZN(
        n19512) );
  NAND2_X1 U18011 ( .A1(n19598), .A2(n19512), .ZN(n17962) );
  OAI211_X1 U18012 ( .C1(n14415), .C2(n17962), .A(n19603), .B(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n14416) );
  OAI211_X1 U18013 ( .C1(n19519), .C2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n14417), .B(n14416), .ZN(P3_U2853) );
  XNOR2_X1 U18014 ( .A(n14419), .B(n14418), .ZN(n18122) );
  XNOR2_X1 U18015 ( .A(n21079), .B(n18122), .ZN(n14432) );
  NAND2_X1 U18016 ( .A1(n14421), .A2(n14420), .ZN(n14423) );
  NOR2_X1 U18017 ( .A1(n14423), .A2(n14422), .ZN(n14424) );
  OAI21_X4 U18018 ( .B1(n14425), .B2(n14424), .A(n20237), .ZN(n16938) );
  INV_X1 U18019 ( .A(n18122), .ZN(n16734) );
  AOI22_X1 U18020 ( .A1(n20385), .A2(n16734), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n16938), .ZN(n14431) );
  NAND2_X1 U18021 ( .A1(n12631), .A2(n12905), .ZN(n14427) );
  INV_X1 U18022 ( .A(n14428), .ZN(n14429) );
  INV_X1 U18023 ( .A(n20393), .ZN(n14809) );
  NAND2_X1 U18024 ( .A1(n14809), .A2(n20359), .ZN(n14430) );
  OAI211_X1 U18025 ( .C1(n14432), .C2(n20389), .A(n14431), .B(n14430), .ZN(
        P2_U2919) );
  INV_X1 U18026 ( .A(n14433), .ZN(n14434) );
  NAND2_X1 U18027 ( .A1(n14435), .A2(n14434), .ZN(n14436) );
  NOR2_X1 U18028 ( .A1(n14437), .A2(n14436), .ZN(n14438) );
  NOR2_X1 U18029 ( .A1(n14654), .A2(n14438), .ZN(n20372) );
  INV_X1 U18030 ( .A(n20372), .ZN(n14444) );
  NAND2_X1 U18031 ( .A1(n14441), .A2(n14440), .ZN(n14442) );
  NAND2_X1 U18032 ( .A1(n14336), .A2(n14442), .ZN(n20346) );
  MUX2_X1 U18033 ( .A(n20346), .B(n20334), .S(n9713), .Z(n14443) );
  OAI21_X1 U18034 ( .B1(n14444), .B2(n16840), .A(n14443), .ZN(P2_U2883) );
  INV_X1 U18035 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n14446) );
  INV_X1 U18036 ( .A(n14445), .ZN(n15666) );
  OAI222_X1 U18037 ( .A1(n15655), .A2(n15704), .B1(n14446), .B2(n15709), .C1(
        n15666), .C2(n15702), .ZN(P1_U2870) );
  INV_X1 U18038 ( .A(n14447), .ZN(n14449) );
  OR2_X1 U18039 ( .A1(n14449), .A2(n14448), .ZN(n14450) );
  NAND2_X1 U18040 ( .A1(n14449), .A2(n14448), .ZN(n14514) );
  AND2_X1 U18041 ( .A1(n14450), .A2(n14514), .ZN(n21220) );
  NOR2_X1 U18042 ( .A1(n9892), .A2(n14452), .ZN(n14453) );
  OR2_X1 U18043 ( .A1(n14451), .A2(n14453), .ZN(n21292) );
  INV_X1 U18044 ( .A(n21292), .ZN(n21208) );
  INV_X1 U18045 ( .A(n15709), .ZN(n15696) );
  AOI22_X1 U18046 ( .A1(n15697), .A2(n21208), .B1(n15696), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n14454) );
  OAI21_X1 U18047 ( .B1(n14599), .B2(n15702), .A(n14454), .ZN(P1_U2869) );
  NOR2_X1 U18048 ( .A1(n9704), .A2(n14893), .ZN(n14456) );
  OAI22_X1 U18049 ( .A1(n18755), .A2(n14892), .B1(n18754), .B2(n14906), .ZN(
        n14455) );
  AOI211_X1 U18050 ( .C1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .C2(n14457), .A(
        n14456), .B(n14455), .ZN(n14464) );
  AOI22_X1 U18051 ( .A1(n18759), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17693), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14463) );
  AOI22_X1 U18052 ( .A1(n18760), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n18616), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14462) );
  INV_X1 U18053 ( .A(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n18694) );
  OAI22_X1 U18054 ( .A1(n18763), .A2(n18695), .B1(n14983), .B2(n18694), .ZN(
        n14460) );
  INV_X1 U18055 ( .A(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14458) );
  OAI22_X1 U18056 ( .A1(n18715), .A2(n14458), .B1(n17698), .B2(n18688), .ZN(
        n14459) );
  NOR2_X1 U18057 ( .A1(n14460), .A2(n14459), .ZN(n14461) );
  NAND4_X1 U18058 ( .A1(n14464), .A2(n14463), .A3(n14462), .A4(n14461), .ZN(
        n14470) );
  INV_X1 U18059 ( .A(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14465) );
  INV_X1 U18060 ( .A(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n18689) );
  OAI22_X1 U18061 ( .A1(n14465), .A2(n18775), .B1(n18773), .B2(n18689), .ZN(
        n14469) );
  OAI22_X1 U18062 ( .A1(n18794), .A2(n13862), .B1(n18777), .B2(n14467), .ZN(
        n14468) );
  OR3_X1 U18063 ( .A1(n14470), .A2(n14469), .A3(n14468), .ZN(n18890) );
  INV_X1 U18064 ( .A(n18890), .ZN(n14475) );
  OAI211_X1 U18065 ( .C1(P3_EBX_REG_13__SCAN_IN), .C2(n14473), .A(n18808), .B(
        n14790), .ZN(n14474) );
  OAI21_X1 U18066 ( .B1(n14475), .B2(n18808), .A(n14474), .ZN(P3_U2690) );
  INV_X1 U18067 ( .A(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14476) );
  OAI22_X1 U18068 ( .A1(n9704), .A2(n18640), .B1(n17985), .B2(n14476), .ZN(
        n14478) );
  OAI22_X1 U18069 ( .A1(n18755), .A2(n18636), .B1(n18754), .B2(n18647), .ZN(
        n14477) );
  NOR2_X1 U18070 ( .A1(n14478), .A2(n14477), .ZN(n14486) );
  INV_X1 U18071 ( .A(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n22118) );
  AOI22_X1 U18072 ( .A1(n18759), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12013), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14485) );
  AOI22_X1 U18073 ( .A1(n18760), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n18616), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14484) );
  INV_X1 U18074 ( .A(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n18639) );
  OAI22_X1 U18075 ( .A1(n18613), .A2(n14479), .B1(n17695), .B2(n18639), .ZN(
        n14482) );
  INV_X1 U18076 ( .A(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14480) );
  OAI22_X1 U18077 ( .A1(n18715), .A2(n14480), .B1(n17698), .B2(n17615), .ZN(
        n14481) );
  NOR2_X1 U18078 ( .A1(n14482), .A2(n14481), .ZN(n14483) );
  NAND4_X1 U18079 ( .A1(n14486), .A2(n14485), .A3(n14484), .A4(n14483), .ZN(
        n14490) );
  INV_X1 U18080 ( .A(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17614) );
  OAI22_X1 U18081 ( .A1(n18775), .A2(n17616), .B1(n18773), .B2(n17614), .ZN(
        n14489) );
  INV_X1 U18082 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18790) );
  OAI22_X1 U18083 ( .A1(n18790), .A2(n13862), .B1(n18777), .B2(n14487), .ZN(
        n14488) );
  NOR3_X1 U18084 ( .A1(n14490), .A2(n14489), .A3(n14488), .ZN(n17740) );
  INV_X1 U18085 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n18423) );
  NAND4_X1 U18086 ( .A1(n14491), .A2(P3_EBX_REG_13__SCAN_IN), .A3(n18423), 
        .A4(P3_EBX_REG_12__SCAN_IN), .ZN(n14493) );
  NAND3_X1 U18087 ( .A1(n18808), .A2(n14790), .A3(P3_EBX_REG_14__SCAN_IN), 
        .ZN(n14492) );
  OAI211_X1 U18088 ( .C1(n17740), .C2(n18808), .A(n14493), .B(n14492), .ZN(
        P3_U2689) );
  INV_X1 U18089 ( .A(n14654), .ZN(n14495) );
  NOR2_X1 U18090 ( .A1(n14495), .A2(n14494), .ZN(n14497) );
  NAND2_X1 U18091 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14650) );
  INV_X1 U18092 ( .A(n14650), .ZN(n14496) );
  NAND2_X1 U18093 ( .A1(n14654), .A2(n14496), .ZN(n14814) );
  OAI211_X1 U18094 ( .C1(n14497), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n16830), .B(n14814), .ZN(n14502) );
  OR2_X1 U18095 ( .A1(n9883), .A2(n14499), .ZN(n14500) );
  NAND2_X1 U18096 ( .A1(n14498), .A2(n14500), .ZN(n17496) );
  INV_X1 U18097 ( .A(n17496), .ZN(n18106) );
  NAND2_X1 U18098 ( .A1(n18106), .A2(n16835), .ZN(n14501) );
  OAI211_X1 U18099 ( .C1(n16835), .C2(n12626), .A(n14502), .B(n14501), .ZN(
        P2_U2881) );
  XNOR2_X1 U18100 ( .A(n14503), .B(n21300), .ZN(n14508) );
  XNOR2_X1 U18101 ( .A(n14508), .B(n14507), .ZN(n21295) );
  AOI22_X1 U18102 ( .A1(n18048), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n18072), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n14504) );
  OAI21_X1 U18103 ( .B1(n21216), .B2(n18056), .A(n14504), .ZN(n14505) );
  AOI21_X1 U18104 ( .B1(n21220), .B2(n18052), .A(n14505), .ZN(n14506) );
  OAI21_X1 U18105 ( .B1(n21295), .B2(n21105), .A(n14506), .ZN(P1_U2996) );
  AOI22_X1 U18106 ( .A1(n14508), .A2(n14507), .B1(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n14503), .ZN(n14511) );
  XNOR2_X1 U18107 ( .A(n11707), .B(n14509), .ZN(n14510) );
  XNOR2_X1 U18108 ( .A(n14511), .B(n14510), .ZN(n21287) );
  INV_X1 U18109 ( .A(n21287), .ZN(n14519) );
  INV_X1 U18110 ( .A(n14512), .ZN(n14515) );
  AOI21_X1 U18111 ( .B1(n14515), .B2(n14514), .A(n14601), .ZN(n14520) );
  NAND2_X1 U18112 ( .A1(n18072), .A2(P1_REIP_REG_4__SCAN_IN), .ZN(n21283) );
  NAND2_X1 U18113 ( .A1(n18048), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n14516) );
  OAI211_X1 U18114 ( .C1(n18056), .C2(n21194), .A(n21283), .B(n14516), .ZN(
        n14517) );
  AOI21_X1 U18115 ( .B1(n14520), .B2(n18052), .A(n14517), .ZN(n14518) );
  OAI21_X1 U18116 ( .B1(n14519), .B2(n21105), .A(n14518), .ZN(P1_U2995) );
  INV_X1 U18117 ( .A(n14520), .ZN(n21195) );
  OAI21_X1 U18118 ( .B1(n14451), .B2(n14522), .A(n14521), .ZN(n14523) );
  INV_X1 U18119 ( .A(n14523), .ZN(n21281) );
  AOI22_X1 U18120 ( .A1(n15697), .A2(n21281), .B1(n15696), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n14524) );
  OAI21_X1 U18121 ( .B1(n21195), .B2(n15702), .A(n14524), .ZN(P1_U2868) );
  XOR2_X1 U18122 ( .A(n14530), .B(n21058), .Z(n14529) );
  NAND2_X1 U18123 ( .A1(n21045), .A2(n14525), .ZN(n14526) );
  OAI21_X1 U18124 ( .B1(n21045), .B2(n14525), .A(n14526), .ZN(n20387) );
  NOR2_X1 U18125 ( .A1(n21079), .A2(n18122), .ZN(n20388) );
  NOR2_X1 U18126 ( .A1(n20387), .A2(n20388), .ZN(n20386) );
  INV_X1 U18127 ( .A(n14526), .ZN(n14527) );
  NOR2_X1 U18128 ( .A1(n20386), .A2(n14527), .ZN(n14528) );
  NOR2_X1 U18129 ( .A1(n14528), .A2(n14529), .ZN(n16957) );
  AOI21_X1 U18130 ( .B1(n14529), .B2(n14528), .A(n16957), .ZN(n14533) );
  INV_X1 U18131 ( .A(n14530), .ZN(n21056) );
  INV_X1 U18132 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n20423) );
  OAI22_X1 U18133 ( .A1(n21056), .A2(n16934), .B1(n16965), .B2(n20423), .ZN(
        n14531) );
  AOI21_X1 U18134 ( .B1(n14809), .B2(n20434), .A(n14531), .ZN(n14532) );
  OAI21_X1 U18135 ( .B1(n14533), .B2(n20389), .A(n14532), .ZN(P2_U2917) );
  XOR2_X1 U18136 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B(n14814), .Z(n14538)
         );
  NAND2_X1 U18137 ( .A1(n14498), .A2(n14535), .ZN(n14536) );
  NAND2_X1 U18138 ( .A1(n14534), .A2(n14536), .ZN(n17476) );
  MUX2_X1 U18139 ( .A(n17476), .B(n12815), .S(n9713), .Z(n14537) );
  OAI21_X1 U18140 ( .B1(n14538), .B2(n16840), .A(n14537), .ZN(P2_U2880) );
  NOR2_X1 U18141 ( .A1(n21665), .A2(n21480), .ZN(n16282) );
  INV_X1 U18142 ( .A(n21455), .ZN(n14539) );
  NOR2_X1 U18143 ( .A1(n14539), .A2(n21667), .ZN(n21485) );
  OR2_X1 U18144 ( .A1(n13801), .A2(n14540), .ZN(n21479) );
  NAND2_X1 U18145 ( .A1(n10829), .A2(n14542), .ZN(n21659) );
  OR2_X1 U18146 ( .A1(n21479), .A2(n21659), .ZN(n14543) );
  NAND2_X1 U18147 ( .A1(n14543), .A2(n14585), .ZN(n14546) );
  INV_X1 U18148 ( .A(n14546), .ZN(n14544) );
  OAI21_X1 U18149 ( .B1(n21485), .B2(n21672), .A(n14544), .ZN(n14545) );
  NAND2_X1 U18150 ( .A1(n14581), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n14552) );
  AOI22_X1 U18151 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n9698), .B1(DATAI_30_), 
        .B2(n14582), .ZN(n21721) );
  INV_X1 U18152 ( .A(n21721), .ZN(n21628) );
  AOI22_X1 U18153 ( .A1(n14546), .A2(n21679), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n16282), .ZN(n14586) );
  NAND2_X1 U18154 ( .A1(n14547), .A2(DATAI_6_), .ZN(n14549) );
  NAND2_X1 U18155 ( .A1(n15020), .A2(BUF1_REG_6__SCAN_IN), .ZN(n14548) );
  AND2_X1 U18156 ( .A1(n14549), .A2(n14548), .ZN(n15743) );
  OR2_X1 U18157 ( .A1(n15743), .A2(n14757), .ZN(n16405) );
  NAND2_X1 U18158 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n16321), .ZN(n14584) );
  OAI22_X1 U18159 ( .A1(n14586), .A2(n16405), .B1(n14585), .B2(n21598), .ZN(
        n14550) );
  AOI21_X1 U18160 ( .B1(n14588), .B2(n21628), .A(n14550), .ZN(n14551) );
  OAI211_X1 U18161 ( .C1(n21631), .C2(n16323), .A(n14552), .B(n14551), .ZN(
        P1_U3095) );
  AOI22_X2 U18162 ( .A1(DATAI_19_), .A2(n9912), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n9698), .ZN(n21701) );
  NAND2_X1 U18163 ( .A1(n14581), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n14556) );
  AOI22_X1 U18164 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n9698), .B1(DATAI_27_), 
        .B2(n14582), .ZN(n21586) );
  INV_X1 U18165 ( .A(n21586), .ZN(n21698) );
  OR2_X1 U18166 ( .A1(n15757), .A2(n14757), .ZN(n16391) );
  OAI22_X1 U18167 ( .A1(n14586), .A2(n16391), .B1(n14585), .B2(n21585), .ZN(
        n14554) );
  AOI21_X1 U18168 ( .B1(n14588), .B2(n21698), .A(n14554), .ZN(n14555) );
  OAI211_X1 U18169 ( .C1(n21701), .C2(n16323), .A(n14556), .B(n14555), .ZN(
        P1_U3092) );
  NAND2_X1 U18170 ( .A1(n14581), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n14560) );
  AOI22_X1 U18171 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n9698), .B1(DATAI_26_), 
        .B2(n14582), .ZN(n21618) );
  INV_X1 U18172 ( .A(n21618), .ZN(n21692) );
  AND2_X1 U18173 ( .A1(n15762), .A2(n16321), .ZN(n21691) );
  INV_X1 U18174 ( .A(n21691), .ZN(n16356) );
  NAND2_X1 U18175 ( .A1(n14557), .A2(n14576), .ZN(n21581) );
  OAI22_X1 U18176 ( .A1(n14586), .A2(n16356), .B1(n14585), .B2(n21581), .ZN(
        n14558) );
  AOI21_X1 U18177 ( .B1(n14588), .B2(n21692), .A(n14558), .ZN(n14559) );
  OAI211_X1 U18178 ( .C1(n21695), .C2(n16323), .A(n14560), .B(n14559), .ZN(
        P1_U3091) );
  AOI22_X1 U18179 ( .A1(DATAI_17_), .A2(n14582), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n9698), .ZN(n21577) );
  NAND2_X1 U18180 ( .A1(n14581), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n14564) );
  INV_X1 U18181 ( .A(n21689), .ZN(n16351) );
  OR2_X1 U18182 ( .A1(n15767), .A2(n14757), .ZN(n16382) );
  NAND2_X1 U18183 ( .A1(n14561), .A2(n14576), .ZN(n21576) );
  OAI22_X1 U18184 ( .A1(n14586), .A2(n16382), .B1(n14585), .B2(n21576), .ZN(
        n14562) );
  AOI21_X1 U18185 ( .B1(n14588), .B2(n16351), .A(n14562), .ZN(n14563) );
  OAI211_X1 U18186 ( .C1(n21577), .C2(n16323), .A(n14564), .B(n14563), .ZN(
        P1_U3090) );
  AOI22_X1 U18187 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n9698), .B1(DATAI_16_), 
        .B2(n14582), .ZN(n21683) );
  NAND2_X1 U18188 ( .A1(n14581), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n14570) );
  INV_X1 U18189 ( .A(n21643), .ZN(n21680) );
  INV_X1 U18190 ( .A(DATAI_0_), .ZN(n14566) );
  NAND2_X1 U18191 ( .A1(n15020), .A2(BUF1_REG_0__SCAN_IN), .ZN(n14565) );
  OAI21_X1 U18192 ( .B1(n15020), .B2(n14566), .A(n14565), .ZN(n15773) );
  AND2_X1 U18193 ( .A1(n15773), .A2(n16321), .ZN(n21671) );
  INV_X1 U18194 ( .A(n21671), .ZN(n16326) );
  NAND2_X1 U18195 ( .A1(n9724), .A2(n14576), .ZN(n21639) );
  OAI22_X1 U18196 ( .A1(n14586), .A2(n16326), .B1(n14585), .B2(n21639), .ZN(
        n14568) );
  AOI21_X1 U18197 ( .B1(n14588), .B2(n21680), .A(n14568), .ZN(n14569) );
  OAI211_X1 U18198 ( .C1(n21683), .C2(n16323), .A(n14570), .B(n14569), .ZN(
        P1_U3089) );
  AOI22_X2 U18199 ( .A1(DATAI_23_), .A2(n9912), .B1(BUF1_REG_23__SCAN_IN), 
        .B2(n9698), .ZN(n21732) );
  NAND2_X1 U18200 ( .A1(n14581), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n14573) );
  AOI22_X1 U18201 ( .A1(DATAI_31_), .A2(n14582), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n9698), .ZN(n21610) );
  INV_X1 U18202 ( .A(n21610), .ZN(n21726) );
  OR2_X1 U18203 ( .A1(n15739), .A2(n14757), .ZN(n16410) );
  OAI22_X1 U18204 ( .A1(n14586), .A2(n16410), .B1(n14585), .B2(n21602), .ZN(
        n14571) );
  AOI21_X1 U18205 ( .B1(n14588), .B2(n21726), .A(n14571), .ZN(n14572) );
  OAI211_X1 U18206 ( .C1(n21732), .C2(n16323), .A(n14573), .B(n14572), .ZN(
        P1_U3096) );
  NAND2_X1 U18207 ( .A1(n14581), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n14580) );
  AOI22_X1 U18208 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n9698), .B1(DATAI_29_), 
        .B2(n14582), .ZN(n21713) );
  INV_X1 U18209 ( .A(n21713), .ZN(n21546) );
  INV_X1 U18210 ( .A(DATAI_5_), .ZN(n14575) );
  MUX2_X1 U18211 ( .A(n14575), .B(n14574), .S(n15020), .Z(n15748) );
  NOR2_X2 U18212 ( .A1(n15748), .A2(n14757), .ZN(n21709) );
  INV_X1 U18213 ( .A(n21709), .ZN(n16363) );
  NAND2_X1 U18214 ( .A1(n14577), .A2(n14576), .ZN(n21593) );
  OAI22_X1 U18215 ( .A1(n14586), .A2(n16363), .B1(n14585), .B2(n21593), .ZN(
        n14578) );
  AOI21_X1 U18216 ( .B1(n14588), .B2(n21546), .A(n14578), .ZN(n14579) );
  OAI211_X1 U18217 ( .C1(n21597), .C2(n16323), .A(n14580), .B(n14579), .ZN(
        P1_U3094) );
  AOI22_X2 U18218 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n9698), .B1(DATAI_20_), 
        .B2(n9912), .ZN(n21646) );
  NAND2_X1 U18219 ( .A1(n14581), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n14590) );
  AOI22_X1 U18220 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n9698), .B1(DATAI_28_), 
        .B2(n14582), .ZN(n21707) );
  INV_X1 U18221 ( .A(n21707), .ZN(n21621) );
  NOR2_X2 U18222 ( .A1(n15753), .A2(n14757), .ZN(n21703) );
  INV_X1 U18223 ( .A(n21703), .ZN(n16303) );
  OR2_X1 U18224 ( .A1(n10795), .A2(n14584), .ZN(n21644) );
  OAI22_X1 U18225 ( .A1(n14586), .A2(n16303), .B1(n14585), .B2(n21644), .ZN(
        n14587) );
  AOI21_X1 U18226 ( .B1(n14588), .B2(n21621), .A(n14587), .ZN(n14589) );
  OAI211_X1 U18227 ( .C1(n21646), .C2(n16323), .A(n14590), .B(n14589), .ZN(
        P1_U3093) );
  AND2_X1 U18228 ( .A1(n10816), .A2(n14591), .ZN(n14595) );
  INV_X1 U18229 ( .A(n14595), .ZN(n14592) );
  AND2_X1 U18230 ( .A1(n14593), .A2(n14592), .ZN(n14594) );
  INV_X1 U18231 ( .A(n15773), .ZN(n14597) );
  INV_X1 U18232 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n21257) );
  OAI222_X1 U18233 ( .A1(n15681), .A2(n15790), .B1(n15788), .B2(n14597), .C1(
        n15781), .C2(n21257), .ZN(P1_U2904) );
  INV_X1 U18234 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n14598) );
  OAI222_X1 U18235 ( .A1(n14599), .A2(n15790), .B1(n15788), .B2(n15757), .C1(
        n14598), .C2(n15786), .ZN(P1_U2901) );
  INV_X1 U18236 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n21248) );
  OAI222_X1 U18237 ( .A1(n21195), .A2(n15790), .B1(n15753), .B2(n15788), .C1(
        n21248), .C2(n15786), .ZN(P1_U2900) );
  INV_X1 U18238 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n21253) );
  OAI222_X1 U18239 ( .A1(n15673), .A2(n15790), .B1(n15788), .B2(n15767), .C1(
        n15786), .C2(n21253), .ZN(P1_U2903) );
  NAND2_X1 U18240 ( .A1(n14600), .A2(n14601), .ZN(n14826) );
  OAI21_X1 U18241 ( .B1(n14601), .B2(n14600), .A(n14826), .ZN(n21178) );
  INV_X1 U18242 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n21246) );
  OAI222_X1 U18243 ( .A1(n21178), .A2(n15790), .B1(n15748), .B2(n15788), .C1(
        n15781), .C2(n21246), .ZN(P1_U2899) );
  AOI21_X1 U18244 ( .B1(n14603), .B2(n14602), .A(n9743), .ZN(n17441) );
  INV_X1 U18245 ( .A(n17441), .ZN(n14605) );
  AOI22_X1 U18246 ( .A1(n14809), .A2(n16869), .B1(P2_EAX_REG_10__SCAN_IN), 
        .B2(n16938), .ZN(n14604) );
  OAI21_X1 U18247 ( .B1(n14605), .B2(n16963), .A(n14604), .ZN(P2_U2909) );
  INV_X1 U18248 ( .A(n21369), .ZN(n14606) );
  INV_X1 U18249 ( .A(n21410), .ZN(n14607) );
  INV_X1 U18250 ( .A(n21683), .ZN(n21535) );
  INV_X1 U18251 ( .A(n21310), .ZN(n14608) );
  INV_X1 U18252 ( .A(n13801), .ZN(n21309) );
  INV_X1 U18253 ( .A(n21565), .ZN(n14609) );
  NOR2_X1 U18254 ( .A1(n11533), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n21560) );
  NAND2_X1 U18255 ( .A1(n21560), .A2(n21661), .ZN(n21612) );
  OAI21_X1 U18256 ( .B1(n14609), .B2(n21659), .A(n21612), .ZN(n14610) );
  AND2_X1 U18257 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21560), .ZN(
        n14612) );
  AOI22_X1 U18258 ( .A1(n14610), .A2(n21679), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14612), .ZN(n21611) );
  OAI22_X1 U18259 ( .A1(n21611), .A2(n16326), .B1(n21639), .B2(n21612), .ZN(
        n14611) );
  AOI21_X1 U18260 ( .B1(n21624), .B2(n21535), .A(n14611), .ZN(n14616) );
  AOI21_X1 U18261 ( .B1(n21534), .B2(n14613), .A(n14612), .ZN(n14614) );
  INV_X1 U18262 ( .A(n21677), .ZN(n21416) );
  NAND2_X1 U18263 ( .A1(n21635), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n14615) );
  OAI211_X1 U18264 ( .C1(n21643), .C2(n21627), .A(n14616), .B(n14615), .ZN(
        P1_U3121) );
  AOI21_X1 U18265 ( .B1(n14620), .B2(n14618), .A(n14619), .ZN(n20304) );
  INV_X1 U18266 ( .A(n20304), .ZN(n14622) );
  INV_X1 U18267 ( .A(n16846), .ZN(n14621) );
  INV_X1 U18268 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n20402) );
  OAI222_X1 U18269 ( .A1(n14622), .A2(n16963), .B1(n14621), .B2(n20393), .C1(
        n20402), .C2(n16965), .ZN(P2_U2906) );
  XNOR2_X1 U18270 ( .A(n14623), .B(n14624), .ZN(n17495) );
  INV_X1 U18271 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n20415) );
  INV_X1 U18272 ( .A(n16901), .ZN(n20446) );
  OAI222_X1 U18273 ( .A1(n17495), .A2(n16963), .B1(n20415), .B2(n16965), .C1(
        n20393), .C2(n20446), .ZN(P2_U2913) );
  NAND2_X1 U18274 ( .A1(n14626), .A2(n14627), .ZN(n14628) );
  NAND2_X1 U18275 ( .A1(n14625), .A2(n14628), .ZN(n17463) );
  INV_X1 U18276 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n20411) );
  INV_X1 U18277 ( .A(n16885), .ZN(n14629) );
  OAI222_X1 U18278 ( .A1(n17463), .A2(n16963), .B1(n16965), .B2(n20411), .C1(
        n20393), .C2(n14629), .ZN(P2_U2911) );
  INV_X1 U18279 ( .A(n14602), .ZN(n14630) );
  AOI21_X1 U18280 ( .B1(n14631), .B2(n14625), .A(n14630), .ZN(n20319) );
  INV_X1 U18281 ( .A(n20319), .ZN(n14633) );
  INV_X1 U18282 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n20409) );
  INV_X1 U18283 ( .A(n16877), .ZN(n14632) );
  OAI222_X1 U18284 ( .A1(n14633), .A2(n16963), .B1(n16965), .B2(n20409), .C1(
        n20393), .C2(n14632), .ZN(P2_U2910) );
  OR2_X1 U18285 ( .A1(n14635), .A2(n14634), .ZN(n14636) );
  AND2_X1 U18286 ( .A1(n14626), .A2(n14636), .ZN(n17479) );
  INV_X1 U18287 ( .A(n17479), .ZN(n14637) );
  INV_X1 U18288 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n20413) );
  INV_X1 U18289 ( .A(n16893), .ZN(n20452) );
  OAI222_X1 U18290 ( .A1(n14637), .A2(n16963), .B1(n20413), .B2(n16965), .C1(
        n20393), .C2(n20452), .ZN(P2_U2912) );
  NAND2_X1 U18291 ( .A1(n14638), .A2(n14639), .ZN(n14640) );
  NAND2_X1 U18292 ( .A1(n14618), .A2(n14640), .ZN(n17413) );
  INV_X1 U18293 ( .A(n16854), .ZN(n14641) );
  INV_X1 U18294 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n20404) );
  OAI222_X1 U18295 ( .A1(n17413), .A2(n16963), .B1(n14641), .B2(n20393), .C1(
        n20404), .C2(n16965), .ZN(P2_U2907) );
  OR2_X1 U18296 ( .A1(n9743), .A2(n14642), .ZN(n14643) );
  AND2_X1 U18297 ( .A1(n14638), .A2(n14643), .ZN(n17427) );
  INV_X1 U18298 ( .A(n17427), .ZN(n14645) );
  INV_X1 U18299 ( .A(n16863), .ZN(n14644) );
  INV_X1 U18300 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n21936) );
  OAI222_X1 U18301 ( .A1(n14645), .A2(n16963), .B1(n14644), .B2(n20393), .C1(
        n21936), .C2(n16965), .ZN(P2_U2908) );
  NAND2_X1 U18302 ( .A1(n14647), .A2(n14648), .ZN(n14649) );
  NAND2_X1 U18303 ( .A1(n14646), .A2(n14649), .ZN(n17395) );
  NOR2_X1 U18304 ( .A1(n14650), .A2(n20458), .ZN(n14651) );
  NAND4_X1 U18305 ( .A1(n16837), .A2(n14887), .A3(n16831), .A4(n14651), .ZN(
        n14653) );
  NAND2_X1 U18306 ( .A1(n14815), .A2(n14820), .ZN(n14652) );
  NOR2_X1 U18307 ( .A1(n14653), .A2(n14652), .ZN(n15061) );
  NAND2_X1 U18308 ( .A1(n14654), .A2(n15061), .ZN(n16829) );
  INV_X1 U18309 ( .A(n15056), .ZN(n14832) );
  NOR2_X1 U18310 ( .A1(n16829), .A2(n14832), .ZN(n14655) );
  NAND2_X1 U18311 ( .A1(n14655), .A2(n15057), .ZN(n16821) );
  OAI211_X1 U18312 ( .C1(n14655), .C2(n15057), .A(n16821), .B(n16830), .ZN(
        n14657) );
  NAND2_X1 U18313 ( .A1(n9713), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n14656) );
  OAI211_X1 U18314 ( .C1(n17395), .C2(n9713), .A(n14657), .B(n14656), .ZN(
        P2_U2873) );
  AOI22_X1 U18315 ( .A1(n21275), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n21274), .ZN(n14660) );
  NAND2_X1 U18316 ( .A1(n14660), .A2(n14659), .ZN(P1_U2953) );
  AOI22_X1 U18317 ( .A1(n21275), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n21274), .ZN(n14662) );
  NAND2_X1 U18318 ( .A1(n14662), .A2(n14661), .ZN(P1_U2955) );
  AOI22_X1 U18319 ( .A1(n21275), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n21274), .ZN(n14664) );
  NAND2_X1 U18320 ( .A1(n14664), .A2(n14663), .ZN(P1_U2954) );
  AOI22_X1 U18321 ( .A1(n21275), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n21274), .ZN(n14665) );
  NAND2_X1 U18322 ( .A1(n21260), .A2(n15773), .ZN(n14666) );
  NAND2_X1 U18323 ( .A1(n14665), .A2(n14666), .ZN(P1_U2937) );
  AOI22_X1 U18324 ( .A1(n21275), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n21274), .ZN(n14667) );
  NAND2_X1 U18325 ( .A1(n14667), .A2(n14666), .ZN(P1_U2952) );
  AOI22_X1 U18326 ( .A1(n21275), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n21274), .ZN(n14669) );
  INV_X1 U18327 ( .A(n15743), .ZN(n14668) );
  NAND2_X1 U18328 ( .A1(n21260), .A2(n14668), .ZN(n14680) );
  NAND2_X1 U18329 ( .A1(n14669), .A2(n14680), .ZN(P1_U2958) );
  AOI22_X1 U18330 ( .A1(n21275), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n21274), .ZN(n14673) );
  INV_X1 U18331 ( .A(DATAI_13_), .ZN(n14671) );
  MUX2_X1 U18332 ( .A(n14671), .B(n14670), .S(n15020), .Z(n15785) );
  INV_X1 U18333 ( .A(n15785), .ZN(n14672) );
  NAND2_X1 U18334 ( .A1(n21260), .A2(n14672), .ZN(n21272) );
  NAND2_X1 U18335 ( .A1(n14673), .A2(n21272), .ZN(P1_U2950) );
  AOI22_X1 U18336 ( .A1(n21275), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n21274), .ZN(n14675) );
  INV_X1 U18337 ( .A(n15748), .ZN(n14674) );
  NAND2_X1 U18338 ( .A1(n21260), .A2(n14674), .ZN(n14676) );
  NAND2_X1 U18339 ( .A1(n14675), .A2(n14676), .ZN(P1_U2942) );
  AOI22_X1 U18340 ( .A1(n21275), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n21274), .ZN(n14677) );
  NAND2_X1 U18341 ( .A1(n14677), .A2(n14676), .ZN(P1_U2957) );
  AOI22_X1 U18342 ( .A1(n21275), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n21274), .ZN(n14679) );
  NAND2_X1 U18343 ( .A1(n14679), .A2(n14678), .ZN(P1_U2956) );
  AOI22_X1 U18344 ( .A1(n21275), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n21274), .ZN(n14681) );
  NAND2_X1 U18345 ( .A1(n14681), .A2(n14680), .ZN(P1_U2943) );
  AOI22_X1 U18346 ( .A1(n21275), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n21274), .ZN(n14683) );
  NAND2_X1 U18347 ( .A1(n14683), .A2(n14682), .ZN(P1_U2944) );
  INV_X1 U18348 ( .A(n14711), .ZN(n14716) );
  INV_X1 U18349 ( .A(n14684), .ZN(n14688) );
  OAI21_X1 U18350 ( .B1(n14713), .B2(n14688), .A(n21964), .ZN(n14686) );
  NAND2_X1 U18351 ( .A1(n14713), .A2(n14685), .ZN(n14710) );
  AND2_X1 U18352 ( .A1(n14686), .A2(n14710), .ZN(n14690) );
  NAND2_X1 U18353 ( .A1(n14687), .A2(n14730), .ZN(n14700) );
  NAND2_X1 U18354 ( .A1(n14688), .A2(n21964), .ZN(n14697) );
  AOI22_X1 U18355 ( .A1(n14700), .A2(n14697), .B1(n12299), .B2(n14713), .ZN(
        n14689) );
  MUX2_X1 U18356 ( .A(n14690), .B(n14689), .S(n12129), .Z(n14692) );
  NAND2_X1 U18357 ( .A1(n12223), .A2(n9759), .ZN(n14701) );
  OAI211_X1 U18358 ( .C1(n12310), .C2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n14701), .B(n15143), .ZN(n14691) );
  NAND2_X1 U18359 ( .A1(n14692), .A2(n14691), .ZN(n14693) );
  AOI21_X1 U18360 ( .B1(n17530), .B2(n14716), .A(n14693), .ZN(n17554) );
  MUX2_X1 U18361 ( .A(n12129), .B(n17554), .S(n14743), .Z(n14726) );
  INV_X1 U18362 ( .A(n14710), .ZN(n14696) );
  INV_X1 U18363 ( .A(n14713), .ZN(n14694) );
  NOR2_X1 U18364 ( .A1(n14694), .A2(n14685), .ZN(n14695) );
  MUX2_X1 U18365 ( .A(n14696), .B(n14695), .S(n21964), .Z(n14703) );
  NAND2_X1 U18366 ( .A1(n14698), .A2(n14697), .ZN(n14699) );
  MUX2_X1 U18367 ( .A(n14701), .B(n14700), .S(n14699), .Z(n14702) );
  AOI211_X1 U18368 ( .C1(n14704), .C2(n14716), .A(n14703), .B(n14702), .ZN(
        n17549) );
  NAND2_X1 U18369 ( .A1(n17549), .A2(n14743), .ZN(n14705) );
  OAI21_X1 U18370 ( .B1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n14743), .A(
        n14705), .ZN(n14725) );
  INV_X1 U18371 ( .A(n13135), .ZN(n14707) );
  NAND2_X1 U18372 ( .A1(n14707), .A2(n14706), .ZN(n14714) );
  OAI21_X1 U18373 ( .B1(n12312), .B2(n14708), .A(n14714), .ZN(n14709) );
  OAI211_X1 U18374 ( .C1(n14712), .C2(n14711), .A(n14710), .B(n14709), .ZN(
        n17546) );
  INV_X1 U18375 ( .A(n17546), .ZN(n14717) );
  MUX2_X1 U18376 ( .A(n14714), .B(n14713), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n14715) );
  AOI21_X1 U18377 ( .B1(n13822), .B2(n14716), .A(n14715), .ZN(n17537) );
  OAI211_X1 U18378 ( .C1(n14717), .C2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n17537), .ZN(n14718) );
  OAI211_X1 U18379 ( .C1(n22046), .C2(n17546), .A(n14718), .B(n14743), .ZN(
        n14719) );
  NOR2_X1 U18380 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n14719), .ZN(
        n14723) );
  INV_X1 U18381 ( .A(n14726), .ZN(n14722) );
  AOI21_X1 U18382 ( .B1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n14719), .A(
        n14725), .ZN(n14720) );
  OR3_X1 U18383 ( .A1(n14723), .A2(n14722), .A3(n14720), .ZN(n14721) );
  AOI22_X1 U18384 ( .A1(n14723), .A2(n14722), .B1(n21054), .B2(n14721), .ZN(
        n14724) );
  OAI22_X1 U18385 ( .A1(n14726), .A2(n14725), .B1(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n14724), .ZN(n14745) );
  NAND2_X1 U18386 ( .A1(n14731), .A2(n14727), .ZN(n14729) );
  NAND2_X1 U18387 ( .A1(n14736), .A2(n14732), .ZN(n14728) );
  OAI211_X1 U18388 ( .C1(n14731), .C2(n14730), .A(n14729), .B(n14728), .ZN(
        n21086) );
  INV_X1 U18389 ( .A(n14732), .ZN(n14735) );
  OR2_X1 U18390 ( .A1(n13142), .A2(n14733), .ZN(n14734) );
  NAND2_X1 U18391 ( .A1(n14734), .A2(n17597), .ZN(n16418) );
  NAND3_X1 U18392 ( .A1(n14736), .A2(n14735), .A3(n16418), .ZN(n20238) );
  NOR2_X1 U18393 ( .A1(P2_FLUSH_REG_SCAN_IN), .A2(P2_MORE_REG_SCAN_IN), .ZN(
        n14739) );
  OAI211_X1 U18394 ( .C1(n20238), .C2(n14739), .A(n14738), .B(n14737), .ZN(
        n14740) );
  NOR2_X1 U18395 ( .A1(n21086), .A2(n14740), .ZN(n14741) );
  OAI21_X1 U18396 ( .B1(n14743), .B2(n14742), .A(n14741), .ZN(n14744) );
  NOR2_X1 U18397 ( .A1(n14745), .A2(n14744), .ZN(n18143) );
  INV_X1 U18398 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n17538) );
  AOI21_X1 U18399 ( .B1(n18143), .B2(n17538), .A(n17596), .ZN(n14750) );
  OAI211_X1 U18400 ( .C1(n14748), .C2(n14747), .A(P2_STATE2_REG_2__SCAN_IN), 
        .B(n14746), .ZN(n14749) );
  OAI21_X1 U18401 ( .B1(n18135), .B2(n17596), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n14751) );
  NAND2_X1 U18402 ( .A1(n14751), .A2(n18041), .ZN(P2_U3593) );
  OAI21_X1 U18403 ( .B1(n21727), .B2(n10689), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n14756) );
  OR2_X1 U18404 ( .A1(n13801), .A2(n14753), .ZN(n21660) );
  INV_X1 U18405 ( .A(n21660), .ZN(n14755) );
  NAND2_X1 U18406 ( .A1(n14755), .A2(n21564), .ZN(n14760) );
  AOI21_X1 U18407 ( .B1(n14756), .B2(n14760), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n14758) );
  NOR2_X1 U18408 ( .A1(n11533), .A2(n21306), .ZN(n21662) );
  INV_X1 U18409 ( .A(n21662), .ZN(n21664) );
  NOR3_X1 U18410 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21665), .A3(
        n21664), .ZN(n21654) );
  OAI21_X1 U18411 ( .B1(n11533), .B2(n16324), .A(P1_STATE2_REG_2__SCAN_IN), 
        .ZN(n21566) );
  OR2_X1 U18412 ( .A1(n14759), .A2(n10952), .ZN(n21571) );
  INV_X1 U18413 ( .A(n21571), .ZN(n16325) );
  NAND2_X1 U18414 ( .A1(n21656), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n14763) );
  NAND2_X1 U18415 ( .A1(n14759), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21451) );
  INV_X1 U18416 ( .A(n16324), .ZN(n21311) );
  NAND2_X1 U18417 ( .A1(n21311), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21570) );
  OAI22_X1 U18418 ( .A1(n14760), .A2(n21667), .B1(n21451), .B2(n21570), .ZN(
        n21655) );
  INV_X1 U18419 ( .A(n21655), .ZN(n14780) );
  INV_X1 U18420 ( .A(n21654), .ZN(n14779) );
  OAI22_X1 U18421 ( .A1(n14780), .A2(n16326), .B1(n21639), .B2(n14779), .ZN(
        n14761) );
  AOI21_X1 U18422 ( .B1(n10689), .B2(n21680), .A(n14761), .ZN(n14762) );
  OAI211_X1 U18423 ( .C1(n21683), .C2(n21720), .A(n14763), .B(n14762), .ZN(
        P1_U3145) );
  NAND2_X1 U18424 ( .A1(n21656), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n14766) );
  OAI22_X1 U18425 ( .A1(n14780), .A2(n16410), .B1(n21602), .B2(n14779), .ZN(
        n14764) );
  AOI21_X1 U18426 ( .B1(n10689), .B2(n21726), .A(n14764), .ZN(n14765) );
  OAI211_X1 U18427 ( .C1(n21732), .C2(n21720), .A(n14766), .B(n14765), .ZN(
        P1_U3152) );
  NAND2_X1 U18428 ( .A1(n21656), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n14769) );
  OAI22_X1 U18429 ( .A1(n14780), .A2(n16356), .B1(n21581), .B2(n14779), .ZN(
        n14767) );
  AOI21_X1 U18430 ( .B1(n10689), .B2(n21692), .A(n14767), .ZN(n14768) );
  OAI211_X1 U18431 ( .C1(n21695), .C2(n21720), .A(n14769), .B(n14768), .ZN(
        P1_U3147) );
  NAND2_X1 U18432 ( .A1(n21656), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n14772) );
  OAI22_X1 U18433 ( .A1(n14780), .A2(n16382), .B1(n21576), .B2(n14779), .ZN(
        n14770) );
  AOI21_X1 U18434 ( .B1(n10689), .B2(n16351), .A(n14770), .ZN(n14771) );
  OAI211_X1 U18435 ( .C1(n21577), .C2(n21720), .A(n14772), .B(n14771), .ZN(
        P1_U3146) );
  NAND2_X1 U18436 ( .A1(n21656), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n14775) );
  OAI22_X1 U18437 ( .A1(n14780), .A2(n16303), .B1(n14779), .B2(n21644), .ZN(
        n14773) );
  AOI21_X1 U18438 ( .B1(n10689), .B2(n21621), .A(n14773), .ZN(n14774) );
  OAI211_X1 U18439 ( .C1(n21646), .C2(n21720), .A(n14775), .B(n14774), .ZN(
        P1_U3149) );
  NAND2_X1 U18440 ( .A1(n21656), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n14778) );
  OAI22_X1 U18441 ( .A1(n14780), .A2(n16405), .B1(n21598), .B2(n14779), .ZN(
        n14776) );
  AOI21_X1 U18442 ( .B1(n10689), .B2(n21628), .A(n14776), .ZN(n14777) );
  OAI211_X1 U18443 ( .C1(n21631), .C2(n21720), .A(n14778), .B(n14777), .ZN(
        P1_U3151) );
  NAND2_X1 U18444 ( .A1(n21656), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n14783) );
  OAI22_X1 U18445 ( .A1(n14780), .A2(n16363), .B1(n21593), .B2(n14779), .ZN(
        n14781) );
  AOI21_X1 U18446 ( .B1(n10689), .B2(n21546), .A(n14781), .ZN(n14782) );
  OAI211_X1 U18447 ( .C1(n21597), .C2(n21720), .A(n14783), .B(n14782), .ZN(
        P1_U3150) );
  INV_X1 U18448 ( .A(n14784), .ZN(n14787) );
  INV_X1 U18449 ( .A(n14785), .ZN(n14786) );
  NAND2_X1 U18450 ( .A1(n14787), .A2(n14786), .ZN(n14789) );
  AND2_X1 U18451 ( .A1(n14789), .A2(n14788), .ZN(n21159) );
  INV_X1 U18452 ( .A(n21159), .ZN(n14843) );
  INV_X1 U18453 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n22079) );
  OAI222_X1 U18454 ( .A1(n14843), .A2(n15790), .B1(n15739), .B2(n15788), .C1(
        n15781), .C2(n22079), .ZN(P1_U2897) );
  OAI21_X1 U18455 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n9870), .A(n18710), .ZN(
        n14805) );
  AOI22_X1 U18456 ( .A1(n13659), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14896), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14795) );
  AOI22_X1 U18457 ( .A1(n10682), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n18616), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14794) );
  AOI22_X1 U18458 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18759), .B1(
        n18692), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14793) );
  INV_X1 U18459 ( .A(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n18617) );
  OAI22_X1 U18460 ( .A1(n17695), .A2(n18617), .B1(n17698), .B2(n14926), .ZN(
        n14791) );
  INV_X1 U18461 ( .A(n14791), .ZN(n14792) );
  NAND4_X1 U18462 ( .A1(n14795), .A2(n14794), .A3(n14793), .A4(n14792), .ZN(
        n14803) );
  AOI22_X1 U18463 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n9712), .B1(
        n14457), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14797) );
  AOI22_X1 U18464 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n9705), .B1(
        n18652), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14796) );
  NAND2_X1 U18465 ( .A1(n14797), .A2(n14796), .ZN(n14802) );
  INV_X1 U18466 ( .A(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14798) );
  OAI22_X1 U18467 ( .A1(n14799), .A2(n18775), .B1(n18773), .B2(n14798), .ZN(
        n14801) );
  INV_X1 U18468 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18785) );
  OAI22_X1 U18469 ( .A1(n18785), .A2(n13862), .B1(n18777), .B2(n14155), .ZN(
        n14800) );
  OR4_X1 U18470 ( .A1(n14803), .A2(n14802), .A3(n14801), .A4(n14800), .ZN(
        n18886) );
  NAND2_X1 U18471 ( .A1(n18812), .A2(n18886), .ZN(n14804) );
  OAI21_X1 U18472 ( .B1(n14805), .B2(n18812), .A(n14804), .ZN(P3_U2688) );
  NOR2_X1 U18473 ( .A1(n14619), .A2(n14807), .ZN(n14808) );
  OR2_X1 U18474 ( .A1(n14806), .A2(n14808), .ZN(n16602) );
  AOI22_X1 U18475 ( .A1(n14809), .A2(n15340), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n16938), .ZN(n14810) );
  OAI21_X1 U18476 ( .B1(n16602), .B2(n16963), .A(n14810), .ZN(P2_U2905) );
  AND2_X1 U18477 ( .A1(n14534), .A2(n14811), .ZN(n14813) );
  OR2_X1 U18478 ( .A1(n14813), .A2(n14812), .ZN(n17461) );
  NOR2_X1 U18479 ( .A1(n14814), .A2(n20458), .ZN(n14816) );
  NAND2_X1 U18480 ( .A1(n14816), .A2(n14815), .ZN(n14886) );
  OAI211_X1 U18481 ( .C1(n14816), .C2(n14815), .A(n14886), .B(n16830), .ZN(
        n14818) );
  NAND2_X1 U18482 ( .A1(n9713), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n14817) );
  OAI211_X1 U18483 ( .C1(n17461), .C2(n9713), .A(n14818), .B(n14817), .ZN(
        P2_U2879) );
  AOI21_X1 U18484 ( .B1(n14819), .B2(n14788), .A(n9792), .ZN(n21148) );
  INV_X1 U18485 ( .A(n21148), .ZN(n15707) );
  OAI222_X1 U18486 ( .A1(n15707), .A2(n15790), .B1(n15735), .B2(n15788), .C1(
        n21241), .C2(n15786), .ZN(P1_U2896) );
  INV_X1 U18487 ( .A(n14820), .ZN(n14885) );
  XNOR2_X1 U18488 ( .A(n14886), .B(n14885), .ZN(n14825) );
  NOR2_X1 U18489 ( .A1(n14812), .A2(n14822), .ZN(n14823) );
  OR2_X1 U18490 ( .A1(n14821), .A2(n14823), .ZN(n20316) );
  MUX2_X1 U18491 ( .A(n20316), .B(n10510), .S(n9713), .Z(n14824) );
  OAI21_X1 U18492 ( .B1(n14825), .B2(n16840), .A(n14824), .ZN(P2_U2878) );
  INV_X1 U18493 ( .A(n14826), .ZN(n14828) );
  NOR2_X1 U18494 ( .A1(n14828), .A2(n14827), .ZN(n14829) );
  NOR2_X1 U18495 ( .A1(n14784), .A2(n14829), .ZN(n21169) );
  INV_X1 U18496 ( .A(n21169), .ZN(n14831) );
  INV_X1 U18497 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n21244) );
  OAI222_X1 U18498 ( .A1(n14831), .A2(n15790), .B1(n15743), .B2(n15788), .C1(
        n15781), .C2(n21244), .ZN(P1_U2898) );
  XNOR2_X1 U18499 ( .A(n9758), .B(n14840), .ZN(n18071) );
  INV_X1 U18500 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n14830) );
  OAI222_X1 U18501 ( .A1(n14831), .A2(n15702), .B1(n15704), .B2(n18071), .C1(
        n15709), .C2(n14830), .ZN(P1_U2866) );
  XNOR2_X1 U18502 ( .A(n16829), .B(n14832), .ZN(n14838) );
  INV_X1 U18503 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n14836) );
  OR2_X1 U18504 ( .A1(n14833), .A2(n14834), .ZN(n14835) );
  AND2_X1 U18505 ( .A1(n14647), .A2(n14835), .ZN(n17140) );
  INV_X1 U18506 ( .A(n17140), .ZN(n20301) );
  MUX2_X1 U18507 ( .A(n14836), .B(n20301), .S(n16835), .Z(n14837) );
  OAI21_X1 U18508 ( .B1(n14838), .B2(n16840), .A(n14837), .ZN(P2_U2874) );
  AOI21_X1 U18509 ( .B1(n9758), .B2(n14840), .A(n14839), .ZN(n14842) );
  OR2_X1 U18510 ( .A1(n14842), .A2(n14841), .ZN(n18063) );
  INV_X1 U18511 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n14844) );
  OAI222_X1 U18512 ( .A1(n18063), .A2(n15704), .B1(n14844), .B2(n15709), .C1(
        n15702), .C2(n14843), .ZN(P1_U2865) );
  OR2_X1 U18513 ( .A1(n9792), .A2(n14846), .ZN(n14847) );
  NAND2_X1 U18514 ( .A1(n14845), .A2(n14847), .ZN(n21133) );
  INV_X1 U18515 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n14848) );
  OAI222_X1 U18516 ( .A1(n21133), .A2(n15790), .B1(n15729), .B2(n15788), .C1(
        n14848), .C2(n15786), .ZN(P1_U2895) );
  OAI21_X1 U18517 ( .B1(n20824), .B2(n20829), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n14861) );
  AND2_X1 U18518 ( .A1(n14850), .A2(n20618), .ZN(n20546) );
  NAND2_X1 U18519 ( .A1(n20545), .A2(n20546), .ZN(n14860) );
  NAND3_X1 U18520 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n22046), .ZN(n20836) );
  NOR2_X1 U18521 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20836), .ZN(
        n20822) );
  INV_X1 U18522 ( .A(n20822), .ZN(n14851) );
  AND2_X1 U18523 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n14851), .ZN(n14852) );
  NAND2_X1 U18524 ( .A1(n14853), .A2(n14852), .ZN(n14863) );
  NAND2_X1 U18525 ( .A1(n17596), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n14855) );
  NAND2_X1 U18526 ( .A1(n14856), .A2(n14855), .ZN(n18138) );
  NAND2_X1 U18527 ( .A1(n18138), .A2(n14857), .ZN(n14858) );
  OAI211_X1 U18528 ( .C1(n20822), .C2(n20834), .A(n14863), .B(n20896), .ZN(
        n14859) );
  INV_X1 U18529 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14869) );
  AOI22_X1 U18530 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20454), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n20453), .ZN(n20479) );
  AOI22_X1 U18531 ( .A1(n20829), .A2(n20935), .B1(n20824), .B2(n20934), .ZN(
        n14868) );
  NAND3_X1 U18532 ( .A1(n20545), .A2(n20834), .A3(n20546), .ZN(n14865) );
  INV_X1 U18533 ( .A(n14863), .ZN(n14864) );
  AND2_X1 U18534 ( .A1(n20896), .A2(n16918), .ZN(n20933) );
  NOR2_X2 U18535 ( .A1(n14866), .A2(n20450), .ZN(n20932) );
  AOI22_X1 U18536 ( .A1(n20823), .A2(n20933), .B1(n20822), .B2(n20932), .ZN(
        n14867) );
  OAI211_X1 U18537 ( .C1(n20828), .C2(n14869), .A(n14868), .B(n14867), .ZN(
        P2_U3148) );
  INV_X1 U18538 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14873) );
  AOI22_X1 U18539 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20454), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n20453), .ZN(n20587) );
  AOI22_X1 U18540 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n20453), .B1(
        BUF1_REG_24__SCAN_IN), .B2(n20454), .ZN(n20843) );
  INV_X1 U18541 ( .A(n20843), .ZN(n20906) );
  AOI22_X1 U18542 ( .A1(n20829), .A2(n20907), .B1(n20824), .B2(n20906), .ZN(
        n14872) );
  NAND2_X1 U18543 ( .A1(n20359), .A2(n20896), .ZN(n20725) );
  INV_X1 U18544 ( .A(n20450), .ZN(n17570) );
  AND2_X1 U18545 ( .A1(n14870), .A2(n17570), .ZN(n20904) );
  AOI22_X1 U18546 ( .A1(n20823), .A2(n20905), .B1(n20904), .B2(n20822), .ZN(
        n14871) );
  OAI211_X1 U18547 ( .C1(n20828), .C2(n14873), .A(n14872), .B(n14871), .ZN(
        P2_U3144) );
  INV_X1 U18548 ( .A(n15788), .ZN(n15792) );
  AOI22_X1 U18549 ( .A1(n15792), .A2(n15762), .B1(P1_EAX_REG_2__SCAN_IN), .B2(
        n13423), .ZN(n14874) );
  OAI21_X1 U18550 ( .B1(n15666), .B2(n15790), .A(n14874), .ZN(P1_U2902) );
  NAND2_X1 U18551 ( .A1(n14876), .A2(n14877), .ZN(n14878) );
  NAND2_X1 U18552 ( .A1(n14875), .A2(n14878), .ZN(n21127) );
  INV_X1 U18553 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n21985) );
  OAI222_X1 U18554 ( .A1(n21127), .A2(n15704), .B1(n15709), .B2(n21985), .C1(
        n15702), .C2(n21133), .ZN(P1_U2863) );
  NAND2_X1 U18555 ( .A1(n14845), .A2(n14880), .ZN(n14881) );
  NAND2_X1 U18556 ( .A1(n14879), .A2(n14881), .ZN(n15990) );
  XNOR2_X1 U18557 ( .A(n14875), .B(n15629), .ZN(n16233) );
  AOI22_X1 U18558 ( .A1(n16233), .A2(n15697), .B1(n15696), .B2(
        P1_EBX_REG_10__SCAN_IN), .ZN(n14882) );
  OAI21_X1 U18559 ( .B1(n15990), .B2(n15702), .A(n14882), .ZN(P1_U2862) );
  OAI21_X1 U18560 ( .B1(n14821), .B2(n14884), .A(n14883), .ZN(n17438) );
  NOR2_X1 U18561 ( .A1(n14886), .A2(n14885), .ZN(n14888) );
  NAND2_X1 U18562 ( .A1(n14888), .A2(n14887), .ZN(n16836) );
  OAI211_X1 U18563 ( .C1(n14888), .C2(n14887), .A(n16836), .B(n16830), .ZN(
        n14890) );
  NAND2_X1 U18564 ( .A1(n9713), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n14889) );
  OAI211_X1 U18565 ( .C1(n17438), .C2(n9713), .A(n14890), .B(n14889), .ZN(
        P2_U2877) );
  INV_X1 U18566 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n14891) );
  OAI222_X1 U18567 ( .A1(n15990), .A2(n15790), .B1(n15723), .B2(n15788), .C1(
        n14891), .C2(n15786), .ZN(P1_U2894) );
  AND2_X1 U18568 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n18604) );
  NAND2_X1 U18569 ( .A1(n18814), .A2(n18606), .ZN(n18816) );
  INV_X1 U18570 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n21981) );
  NAND2_X1 U18571 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n18727), .ZN(n17688) );
  NAND2_X1 U18572 ( .A1(n18672), .A2(P3_EBX_REG_26__SCAN_IN), .ZN(n18670) );
  OAI21_X1 U18573 ( .B1(n18604), .B2(n18816), .A(n18674), .ZN(n18664) );
  AOI22_X1 U18574 ( .A1(n9712), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14457), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14904) );
  OAI22_X1 U18575 ( .A1(n18613), .A2(n18693), .B1(n14983), .B2(n14892), .ZN(
        n14895) );
  OAI22_X1 U18576 ( .A1(n18715), .A2(n14893), .B1(n17698), .B2(n18694), .ZN(
        n14894) );
  NOR2_X1 U18577 ( .A1(n14895), .A2(n14894), .ZN(n14903) );
  AOI22_X1 U18578 ( .A1(n9706), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n18652), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14902) );
  NAND2_X1 U18579 ( .A1(n14896), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n14900) );
  NAND2_X1 U18580 ( .A1(n18759), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n14899) );
  NAND2_X1 U18581 ( .A1(n17631), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n14898) );
  NAND2_X1 U18582 ( .A1(n18692), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n14897) );
  AND4_X1 U18583 ( .A1(n14900), .A2(n14899), .A3(n14898), .A4(n14897), .ZN(
        n14901) );
  NAND4_X1 U18584 ( .A1(n14904), .A2(n14903), .A3(n14902), .A4(n14901), .ZN(
        n14912) );
  NAND2_X1 U18585 ( .A1(n18624), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n14910) );
  NAND2_X1 U18586 ( .A1(n14968), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n14909) );
  INV_X1 U18587 ( .A(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14905) );
  OR2_X1 U18588 ( .A1(n18775), .A2(n14905), .ZN(n14908) );
  OR2_X1 U18589 ( .A1(n18773), .A2(n14906), .ZN(n14907) );
  NAND4_X1 U18590 ( .A1(n14910), .A2(n14909), .A3(n14908), .A4(n14907), .ZN(
        n14911) );
  NOR2_X1 U18591 ( .A1(n14912), .A2(n14911), .ZN(n18635) );
  NOR2_X1 U18592 ( .A1(n17985), .A2(n18776), .ZN(n14915) );
  INV_X1 U18593 ( .A(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14913) );
  OAI22_X1 U18594 ( .A1(n18755), .A2(n14913), .B1(n18754), .B2(n18762), .ZN(
        n14914) );
  AOI211_X1 U18595 ( .C1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .C2(n9712), .A(
        n14915), .B(n14914), .ZN(n14922) );
  AOI22_X1 U18596 ( .A1(n18759), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n18692), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14921) );
  AOI22_X1 U18597 ( .A1(n18760), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18616), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14920) );
  OAI22_X1 U18598 ( .A1(n18613), .A2(n14916), .B1(n14983), .B2(n18756), .ZN(
        n14918) );
  INV_X1 U18599 ( .A(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n18761) );
  OAI22_X1 U18600 ( .A1(n18715), .A2(n18752), .B1(n17698), .B2(n18761), .ZN(
        n14917) );
  NOR2_X1 U18601 ( .A1(n14918), .A2(n14917), .ZN(n14919) );
  NAND4_X1 U18602 ( .A1(n14922), .A2(n14921), .A3(n14920), .A4(n14919), .ZN(
        n14925) );
  INV_X1 U18603 ( .A(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n21925) );
  OAI22_X1 U18604 ( .A1(n18775), .A2(n21925), .B1(n18773), .B2(n18753), .ZN(
        n14924) );
  INV_X1 U18605 ( .A(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18765) );
  OAI22_X1 U18606 ( .A1(n18714), .A2(n18777), .B1(n13862), .B2(n18765), .ZN(
        n14923) );
  NOR3_X1 U18607 ( .A1(n14925), .A2(n14924), .A3(n14923), .ZN(n18684) );
  NOR2_X1 U18608 ( .A1(n18754), .A2(n14926), .ZN(n14928) );
  OAI22_X1 U18609 ( .A1(n14798), .A2(n9704), .B1(n17985), .B2(n18785), .ZN(
        n14927) );
  AOI211_X1 U18610 ( .C1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .C2(n9706), .A(
        n14928), .B(n14927), .ZN(n14936) );
  AOI22_X1 U18611 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18692), .B1(
        n17630), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14935) );
  AOI22_X1 U18612 ( .A1(n18760), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n18616), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14934) );
  OAI22_X1 U18613 ( .A1(n18617), .A2(n18613), .B1(n14983), .B2(n18614), .ZN(
        n14932) );
  OAI22_X1 U18614 ( .A1(n18715), .A2(n14930), .B1(n17698), .B2(n14929), .ZN(
        n14931) );
  NOR2_X1 U18615 ( .A1(n14932), .A2(n14931), .ZN(n14933) );
  NAND4_X1 U18616 ( .A1(n14936), .A2(n14935), .A3(n14934), .A4(n14933), .ZN(
        n14942) );
  INV_X1 U18617 ( .A(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14938) );
  INV_X1 U18618 ( .A(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14937) );
  OAI22_X1 U18619 ( .A1(n18775), .A2(n14938), .B1(n18773), .B2(n14937), .ZN(
        n14941) );
  INV_X1 U18620 ( .A(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14939) );
  OAI22_X1 U18621 ( .A1(n14155), .A2(n13862), .B1(n18777), .B2(n14939), .ZN(
        n14940) );
  NOR3_X1 U18622 ( .A1(n14942), .A2(n14941), .A3(n14940), .ZN(n18685) );
  NOR2_X1 U18623 ( .A1(n18684), .A2(n18685), .ZN(n18683) );
  OAI22_X1 U18624 ( .A1(n18613), .A2(n17694), .B1(n14983), .B2(n14943), .ZN(
        n14944) );
  INV_X1 U18625 ( .A(n14944), .ZN(n14950) );
  AOI22_X1 U18626 ( .A1(n18760), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n18616), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14949) );
  AOI22_X1 U18627 ( .A1(n18759), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n18692), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14948) );
  OAI22_X1 U18628 ( .A1(n18715), .A2(n14945), .B1(n17698), .B2(n17696), .ZN(
        n14946) );
  INV_X1 U18629 ( .A(n14946), .ZN(n14947) );
  AND4_X1 U18630 ( .A1(n14950), .A2(n14949), .A3(n14948), .A4(n14947), .ZN(
        n14961) );
  NAND2_X1 U18631 ( .A1(n14951), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n14957) );
  NAND2_X1 U18632 ( .A1(n14968), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n14956) );
  OR2_X1 U18633 ( .A1(n18773), .A2(n14952), .ZN(n14955) );
  INV_X1 U18634 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14953) );
  OR2_X1 U18635 ( .A1(n18775), .A2(n14953), .ZN(n14954) );
  AND4_X1 U18636 ( .A1(n14957), .A2(n14956), .A3(n14955), .A4(n14954), .ZN(
        n14960) );
  AOI22_X1 U18637 ( .A1(n9712), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n14457), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14959) );
  AOI22_X1 U18638 ( .A1(n9705), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n18652), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14958) );
  NAND4_X1 U18639 ( .A1(n14961), .A2(n14960), .A3(n14959), .A4(n14958), .ZN(
        n18681) );
  AND2_X1 U18640 ( .A1(n18683), .A2(n18681), .ZN(n18679) );
  OAI22_X1 U18641 ( .A1(n18613), .A2(n17670), .B1(n14983), .B2(n18730), .ZN(
        n14962) );
  INV_X1 U18642 ( .A(n14962), .ZN(n14967) );
  AOI22_X1 U18643 ( .A1(n18760), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18616), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n14966) );
  AOI22_X1 U18644 ( .A1(n18759), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n18692), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14965) );
  INV_X1 U18645 ( .A(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n18733) );
  OAI22_X1 U18646 ( .A1(n18715), .A2(n18728), .B1(n17698), .B2(n18733), .ZN(
        n14963) );
  INV_X1 U18647 ( .A(n14963), .ZN(n14964) );
  AND4_X1 U18648 ( .A1(n14967), .A2(n14966), .A3(n14965), .A4(n14964), .ZN(
        n14977) );
  NAND2_X1 U18649 ( .A1(n18624), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n14973) );
  NAND2_X1 U18650 ( .A1(n14968), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n14972) );
  INV_X1 U18651 ( .A(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14969) );
  OR2_X1 U18652 ( .A1(n18775), .A2(n14969), .ZN(n14971) );
  OR2_X1 U18653 ( .A1(n18773), .A2(n18729), .ZN(n14970) );
  AND4_X1 U18654 ( .A1(n14973), .A2(n14972), .A3(n14971), .A4(n14970), .ZN(
        n14976) );
  AOI22_X1 U18655 ( .A1(n9712), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14457), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14975) );
  AOI22_X1 U18656 ( .A1(n9705), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n18652), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14974) );
  NAND4_X1 U18657 ( .A1(n14977), .A2(n14976), .A3(n14975), .A4(n14974), .ZN(
        n18677) );
  NAND2_X1 U18658 ( .A1(n18679), .A2(n18677), .ZN(n18676) );
  NOR2_X1 U18659 ( .A1(n18754), .A2(n13896), .ZN(n14981) );
  OAI22_X1 U18660 ( .A1(n9704), .A2(n14979), .B1(n17985), .B2(n14978), .ZN(
        n14980) );
  AOI211_X1 U18661 ( .C1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .C2(n9706), .A(
        n14981), .B(n14980), .ZN(n14990) );
  INV_X1 U18662 ( .A(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17650) );
  AOI22_X1 U18663 ( .A1(n18759), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18692), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14989) );
  AOI22_X1 U18664 ( .A1(n18760), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18616), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14988) );
  OAI22_X1 U18665 ( .A1(n18613), .A2(n17653), .B1(n14983), .B2(n14982), .ZN(
        n14986) );
  OAI22_X1 U18666 ( .A1(n18715), .A2(n14984), .B1(n17698), .B2(n17654), .ZN(
        n14985) );
  NOR2_X1 U18667 ( .A1(n14986), .A2(n14985), .ZN(n14987) );
  NAND4_X1 U18668 ( .A1(n14990), .A2(n14989), .A3(n14988), .A4(n14987), .ZN(
        n14995) );
  OAI22_X1 U18669 ( .A1(n18775), .A2(n14096), .B1(n18773), .B2(n14991), .ZN(
        n14994) );
  OAI22_X1 U18670 ( .A1(n13862), .A2(n14992), .B1(n18777), .B2(n17655), .ZN(
        n14993) );
  NOR3_X1 U18671 ( .A1(n14995), .A2(n14994), .A3(n14993), .ZN(n18671) );
  NOR2_X1 U18672 ( .A1(n18676), .A2(n18671), .ZN(n18837) );
  OAI22_X1 U18673 ( .A1(n9704), .A2(n17641), .B1(n17985), .B2(n14996), .ZN(
        n14998) );
  INV_X1 U18674 ( .A(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17640) );
  OAI22_X1 U18675 ( .A1(n18755), .A2(n17640), .B1(n18754), .B2(n17626), .ZN(
        n14997) );
  NOR2_X1 U18676 ( .A1(n14998), .A2(n14997), .ZN(n15006) );
  AOI22_X1 U18677 ( .A1(n18759), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n18692), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n15005) );
  AOI22_X1 U18678 ( .A1(n18760), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18616), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15004) );
  OAI22_X1 U18679 ( .A1(n18613), .A2(n17624), .B1(n11972), .B2(n14999), .ZN(
        n15002) );
  OAI22_X1 U18680 ( .A1(n18715), .A2(n15000), .B1(n17698), .B2(n17625), .ZN(
        n15001) );
  NOR2_X1 U18681 ( .A1(n15002), .A2(n15001), .ZN(n15003) );
  AND4_X1 U18682 ( .A1(n15006), .A2(n15005), .A3(n15004), .A4(n15003), .ZN(
        n15009) );
  AOI22_X1 U18683 ( .A1(n18743), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18742), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15008) );
  AOI22_X1 U18684 ( .A1(n14951), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n18646), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15007) );
  NAND3_X1 U18685 ( .A1(n15009), .A2(n15008), .A3(n15007), .ZN(n18836) );
  NAND2_X1 U18686 ( .A1(n18837), .A2(n18836), .ZN(n18835) );
  XOR2_X1 U18687 ( .A(n18635), .B(n18835), .Z(n18830) );
  AOI22_X1 U18688 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n18664), .B1(n18812), 
        .B2(n18830), .ZN(n15013) );
  INV_X1 U18689 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n15011) );
  INV_X1 U18690 ( .A(n18670), .ZN(n15010) );
  NAND3_X1 U18691 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n15011), .A3(n15010), 
        .ZN(n15012) );
  NAND2_X1 U18692 ( .A1(n15013), .A2(n15012), .ZN(P3_U2675) );
  AOI21_X1 U18693 ( .B1(n18087), .B2(n15014), .A(n21804), .ZN(n15018) );
  OAI22_X1 U18694 ( .A1(n15676), .A2(n15015), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n16270), .ZN(n17993) );
  OAI22_X1 U18695 ( .A1(n21800), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n15370), .ZN(n15016) );
  AOI21_X1 U18696 ( .B1(n18087), .B2(n17993), .A(n15016), .ZN(n15017) );
  OAI22_X1 U18697 ( .A1(n15018), .A2(n10144), .B1(n15017), .B2(n21804), .ZN(
        P1_U3474) );
  INV_X1 U18698 ( .A(DATAI_14_), .ZN(n15022) );
  MUX2_X1 U18699 ( .A(n15022), .B(n15021), .S(n15020), .Z(n21258) );
  OAI22_X1 U18700 ( .A1(n15768), .A2(n21258), .B1(n15023), .B2(n15781), .ZN(
        n15024) );
  AOI21_X1 U18701 ( .B1(BUF1_REG_30__SCAN_IN), .B2(n15770), .A(n15024), .ZN(
        n15026) );
  NAND2_X1 U18702 ( .A1(n13436), .A2(DATAI_30_), .ZN(n15025) );
  OAI211_X1 U18703 ( .C1(n15043), .C2(n15790), .A(n15026), .B(n15025), .ZN(
        P1_U2874) );
  AOI22_X1 U18704 ( .A1(n15378), .A2(n9703), .B1(n15027), .B2(n9780), .ZN(
        n15029) );
  XOR2_X1 U18705 ( .A(n15030), .B(n15029), .Z(n16017) );
  INV_X1 U18706 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n15042) );
  INV_X1 U18707 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n15798) );
  NOR2_X1 U18708 ( .A1(n15383), .A2(n15798), .ZN(n15032) );
  OAI21_X1 U18709 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(n15032), .A(n15031), 
        .ZN(n15038) );
  INV_X1 U18710 ( .A(n15033), .ZN(n15034) );
  AOI22_X1 U18711 ( .A1(n21146), .A2(n15036), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n21190), .ZN(n15037) );
  OAI211_X1 U18712 ( .C1(n21205), .C2(n15042), .A(n15038), .B(n15037), .ZN(
        n15039) );
  AOI21_X1 U18713 ( .B1(n16017), .B2(n21209), .A(n15039), .ZN(n15040) );
  OAI21_X1 U18714 ( .B1(n15043), .B2(n15654), .A(n15040), .ZN(P1_U2810) );
  INV_X1 U18715 ( .A(n16017), .ZN(n15041) );
  OAI222_X1 U18716 ( .A1(n15702), .A2(n15043), .B1(n15709), .B2(n15042), .C1(
        n15041), .C2(n15704), .ZN(P1_U2842) );
  AOI22_X1 U18717 ( .A1(n12362), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12379), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15049) );
  AOI22_X1 U18718 ( .A1(n15148), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12451), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15048) );
  AOI22_X1 U18719 ( .A1(n15172), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n15171), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15045) );
  NAND2_X1 U18720 ( .A1(n15173), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n15044) );
  AND2_X1 U18721 ( .A1(n15045), .A2(n15044), .ZN(n15047) );
  AOI22_X1 U18722 ( .A1(n15177), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n15176), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15046) );
  NAND4_X1 U18723 ( .A1(n15049), .A2(n15048), .A3(n15047), .A4(n15046), .ZN(
        n15055) );
  AOI22_X1 U18724 ( .A1(n12524), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12341), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15053) );
  AOI22_X1 U18725 ( .A1(n15125), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12412), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15052) );
  AOI22_X1 U18726 ( .A1(n12371), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12350), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15051) );
  NAND2_X1 U18727 ( .A1(n12525), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n15050) );
  NAND4_X1 U18728 ( .A1(n15053), .A2(n15052), .A3(n15051), .A4(n15050), .ZN(
        n15054) );
  OR2_X1 U18729 ( .A1(n15055), .A2(n15054), .ZN(n16817) );
  NAND3_X1 U18730 ( .A1(n16817), .A2(n15056), .A3(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15059) );
  NAND2_X1 U18731 ( .A1(n16815), .A2(n15057), .ZN(n15058) );
  NOR2_X1 U18732 ( .A1(n15059), .A2(n15058), .ZN(n15060) );
  AND3_X1 U18733 ( .A1(n15061), .A2(n15275), .A3(n15060), .ZN(n15062) );
  AOI22_X1 U18734 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n12362), .B1(
        n12379), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n15071) );
  AOI22_X1 U18735 ( .A1(n15148), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12451), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15070) );
  INV_X1 U18736 ( .A(n15171), .ZN(n15140) );
  NAND2_X1 U18737 ( .A1(n15173), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n15065) );
  NAND2_X1 U18738 ( .A1(n15172), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n15064) );
  OAI211_X1 U18739 ( .C1(n15140), .C2(n15066), .A(n15065), .B(n15064), .ZN(
        n15067) );
  INV_X1 U18740 ( .A(n15067), .ZN(n15069) );
  AOI22_X1 U18741 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n15177), .B1(
        n15176), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15068) );
  NAND4_X1 U18742 ( .A1(n15071), .A2(n15070), .A3(n15069), .A4(n15068), .ZN(
        n15077) );
  AOI22_X1 U18743 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12341), .B1(
        n12524), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15075) );
  AOI22_X1 U18744 ( .A1(n15125), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12412), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n15074) );
  AOI22_X1 U18745 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12371), .B1(
        n12350), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n15073) );
  NAND2_X1 U18746 ( .A1(n12525), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n15072) );
  NAND4_X1 U18747 ( .A1(n15075), .A2(n15074), .A3(n15073), .A4(n15072), .ZN(
        n15076) );
  NOR2_X1 U18748 ( .A1(n15077), .A2(n15076), .ZN(n16811) );
  AOI22_X1 U18749 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n12362), .B1(
        n12379), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15083) );
  AOI22_X1 U18750 ( .A1(n15148), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12451), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15082) );
  AOI22_X1 U18751 ( .A1(n15172), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n15171), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15079) );
  NAND2_X1 U18752 ( .A1(n15173), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n15078) );
  AND2_X1 U18753 ( .A1(n15079), .A2(n15078), .ZN(n15081) );
  AOI22_X1 U18754 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n15177), .B1(
        n15176), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15080) );
  NAND4_X1 U18755 ( .A1(n15083), .A2(n15082), .A3(n15081), .A4(n15080), .ZN(
        n15089) );
  AOI22_X1 U18756 ( .A1(n12524), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12341), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15087) );
  AOI22_X1 U18757 ( .A1(n15125), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12412), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15086) );
  AOI22_X1 U18758 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n12371), .B1(
        n12350), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15085) );
  NAND2_X1 U18759 ( .A1(n12525), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n15084) );
  NAND4_X1 U18760 ( .A1(n15087), .A2(n15086), .A3(n15085), .A4(n15084), .ZN(
        n15088) );
  AOI22_X1 U18761 ( .A1(n12362), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12379), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15097) );
  AOI22_X1 U18762 ( .A1(n15148), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12451), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15096) );
  NAND2_X1 U18763 ( .A1(n15173), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n15091) );
  NAND2_X1 U18764 ( .A1(n15172), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n15090) );
  OAI211_X1 U18765 ( .C1(n15140), .C2(n15092), .A(n15091), .B(n15090), .ZN(
        n15093) );
  INV_X1 U18766 ( .A(n15093), .ZN(n15095) );
  AOI22_X1 U18767 ( .A1(n15177), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n15176), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15094) );
  NAND4_X1 U18768 ( .A1(n15097), .A2(n15096), .A3(n15095), .A4(n15094), .ZN(
        n15103) );
  AOI22_X1 U18769 ( .A1(n12524), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12341), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15101) );
  AOI22_X1 U18770 ( .A1(n15125), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12412), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15100) );
  AOI22_X1 U18771 ( .A1(n12371), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12350), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15099) );
  NAND2_X1 U18772 ( .A1(n12525), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n15098) );
  NAND4_X1 U18773 ( .A1(n15101), .A2(n15100), .A3(n15099), .A4(n15098), .ZN(
        n15102) );
  NOR2_X1 U18774 ( .A1(n15103), .A2(n15102), .ZN(n16804) );
  AOI22_X1 U18775 ( .A1(n12362), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12379), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15109) );
  AOI22_X1 U18776 ( .A1(n15148), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12451), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15108) );
  AOI22_X1 U18777 ( .A1(n15172), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n15171), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15105) );
  NAND2_X1 U18778 ( .A1(n15173), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n15104) );
  AND2_X1 U18779 ( .A1(n15105), .A2(n15104), .ZN(n15107) );
  AOI22_X1 U18780 ( .A1(n15177), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n15176), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15106) );
  NAND4_X1 U18781 ( .A1(n15109), .A2(n15108), .A3(n15107), .A4(n15106), .ZN(
        n15115) );
  AOI22_X1 U18782 ( .A1(n12524), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12341), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15113) );
  AOI22_X1 U18783 ( .A1(n15125), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12412), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15112) );
  AOI22_X1 U18784 ( .A1(n12371), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12350), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15111) );
  NAND2_X1 U18785 ( .A1(n12525), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n15110) );
  NAND4_X1 U18786 ( .A1(n15113), .A2(n15112), .A3(n15111), .A4(n15110), .ZN(
        n15114) );
  NOR2_X1 U18787 ( .A1(n15115), .A2(n15114), .ZN(n16800) );
  INV_X1 U18788 ( .A(n16800), .ZN(n15116) );
  AOI22_X1 U18789 ( .A1(n12362), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12379), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15124) );
  AOI22_X1 U18790 ( .A1(n15148), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12451), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15123) );
  NAND2_X1 U18791 ( .A1(n15173), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n15118) );
  NAND2_X1 U18792 ( .A1(n15172), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n15117) );
  OAI211_X1 U18793 ( .C1(n15140), .C2(n15119), .A(n15118), .B(n15117), .ZN(
        n15120) );
  INV_X1 U18794 ( .A(n15120), .ZN(n15122) );
  AOI22_X1 U18795 ( .A1(n15177), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n15176), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15121) );
  NAND4_X1 U18796 ( .A1(n15124), .A2(n15123), .A3(n15122), .A4(n15121), .ZN(
        n15131) );
  AOI22_X1 U18797 ( .A1(n12524), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12341), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15129) );
  AOI22_X1 U18798 ( .A1(n15125), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12412), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15128) );
  AOI22_X1 U18799 ( .A1(n12371), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12350), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15127) );
  NAND2_X1 U18800 ( .A1(n12525), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n15126) );
  NAND4_X1 U18801 ( .A1(n15129), .A2(n15128), .A3(n15127), .A4(n15126), .ZN(
        n15130) );
  NOR2_X1 U18802 ( .A1(n15131), .A2(n15130), .ZN(n16792) );
  NOR2_X1 U18803 ( .A1(n15179), .A2(n15132), .ZN(n15138) );
  AOI22_X1 U18804 ( .A1(n12524), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12341), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n15134) );
  AOI22_X1 U18805 ( .A1(n12371), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12350), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n15133) );
  OAI211_X1 U18806 ( .C1(n15136), .C2(n15135), .A(n15134), .B(n15133), .ZN(
        n15137) );
  AOI211_X1 U18807 ( .C1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .C2(n12412), .A(
        n15138), .B(n15137), .ZN(n15152) );
  OAI22_X1 U18808 ( .A1(n9783), .A2(n15141), .B1(n15140), .B2(n15139), .ZN(
        n15147) );
  OAI22_X1 U18809 ( .A1(n15145), .A2(n15144), .B1(n15143), .B2(n15142), .ZN(
        n15146) );
  AOI211_X1 U18810 ( .C1(n15173), .C2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n15147), .B(n15146), .ZN(n15151) );
  AOI22_X1 U18811 ( .A1(n12362), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12379), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n15150) );
  AOI22_X1 U18812 ( .A1(n15148), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12451), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n15149) );
  NAND4_X1 U18813 ( .A1(n15152), .A2(n15151), .A3(n15150), .A4(n15149), .ZN(
        n16788) );
  INV_X1 U18814 ( .A(n16773), .ZN(n15215) );
  AND2_X1 U18815 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15154) );
  OR2_X1 U18816 ( .A1(n15154), .A2(n15153), .ZN(n15327) );
  NAND2_X1 U18817 ( .A1(n15326), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n15155) );
  AND3_X1 U18818 ( .A1(n15156), .A2(n15327), .A3(n15155), .ZN(n15162) );
  AOI22_X1 U18819 ( .A1(n15320), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n15323), .ZN(n15161) );
  AOI22_X1 U18820 ( .A1(n9732), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(n9727), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15160) );
  AOI22_X1 U18821 ( .A1(n9729), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n15158), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n15159) );
  NAND4_X1 U18822 ( .A1(n15162), .A2(n15161), .A3(n15160), .A4(n15159), .ZN(
        n15170) );
  INV_X1 U18823 ( .A(n15327), .ZN(n15305) );
  NAND2_X1 U18824 ( .A1(n15326), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n15163) );
  AND3_X1 U18825 ( .A1(n15164), .A2(n15305), .A3(n15163), .ZN(n15168) );
  AOI22_X1 U18826 ( .A1(n15320), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n15323), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15167) );
  AOI22_X1 U18827 ( .A1(n15157), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9727), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n15166) );
  AOI22_X1 U18828 ( .A1(n9730), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n15158), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15165) );
  NAND4_X1 U18829 ( .A1(n15168), .A2(n15167), .A3(n15166), .A4(n15165), .ZN(
        n15169) );
  AND2_X1 U18830 ( .A1(n15170), .A2(n15169), .ZN(n15212) );
  AOI22_X1 U18831 ( .A1(n12362), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12379), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n15186) );
  AOI22_X1 U18832 ( .A1(n15172), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n15171), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15175) );
  NAND2_X1 U18833 ( .A1(n15173), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n15174) );
  AND2_X1 U18834 ( .A1(n15175), .A2(n15174), .ZN(n15185) );
  AOI22_X1 U18835 ( .A1(n15177), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n15176), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15184) );
  INV_X1 U18836 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n15178) );
  OAI22_X1 U18837 ( .A1(n15181), .A2(n15180), .B1(n15179), .B2(n15178), .ZN(
        n15182) );
  INV_X1 U18838 ( .A(n15182), .ZN(n15183) );
  NAND4_X1 U18839 ( .A1(n15186), .A2(n15185), .A3(n15184), .A4(n15183), .ZN(
        n15192) );
  AOI22_X1 U18840 ( .A1(n12524), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12341), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15190) );
  AOI22_X1 U18841 ( .A1(n12451), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12412), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15189) );
  AOI22_X1 U18842 ( .A1(n12371), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12350), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15188) );
  NAND2_X1 U18843 ( .A1(n12525), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n15187) );
  NAND4_X1 U18844 ( .A1(n15190), .A2(n15189), .A3(n15188), .A4(n15187), .ZN(
        n15191) );
  OR2_X1 U18845 ( .A1(n15192), .A2(n15191), .ZN(n15210) );
  AOI22_X1 U18846 ( .A1(n9727), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12190), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15197) );
  NAND2_X1 U18847 ( .A1(n15326), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n15194) );
  NAND2_X1 U18848 ( .A1(n15158), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n15193) );
  AND3_X1 U18849 ( .A1(n15305), .A2(n15194), .A3(n15193), .ZN(n15196) );
  AOI22_X1 U18850 ( .A1(n15320), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9730), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n15195) );
  NAND4_X1 U18851 ( .A1(n15198), .A2(n15197), .A3(n15196), .A4(n15195), .ZN(
        n15206) );
  AOI22_X1 U18852 ( .A1(n15320), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12190), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15204) );
  NAND2_X1 U18853 ( .A1(n15326), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n15200) );
  NAND2_X1 U18854 ( .A1(n15158), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n15199) );
  AND3_X1 U18855 ( .A1(n15200), .A2(n15327), .A3(n15199), .ZN(n15203) );
  AOI22_X1 U18856 ( .A1(n15157), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9729), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15201) );
  NAND4_X1 U18857 ( .A1(n15204), .A2(n15203), .A3(n15202), .A4(n15201), .ZN(
        n15205) );
  AND2_X1 U18858 ( .A1(n15206), .A2(n15205), .ZN(n15208) );
  AND2_X1 U18859 ( .A1(n15210), .A2(n15208), .ZN(n15207) );
  NAND2_X1 U18860 ( .A1(n15207), .A2(n15212), .ZN(n15216) );
  OAI211_X1 U18861 ( .C1(n15212), .C2(n15207), .A(n15275), .B(n15216), .ZN(
        n16778) );
  NOR2_X1 U18862 ( .A1(n15209), .A2(n16775), .ZN(n15211) );
  XNOR2_X1 U18863 ( .A(n15211), .B(n15210), .ZN(n16776) );
  NOR2_X1 U18864 ( .A1(n16778), .A2(n16776), .ZN(n15214) );
  INV_X1 U18865 ( .A(n16776), .ZN(n16774) );
  NAND2_X1 U18866 ( .A1(n15209), .A2(n15212), .ZN(n16777) );
  NOR2_X1 U18867 ( .A1(n16777), .A2(n16775), .ZN(n15213) );
  INV_X1 U18868 ( .A(n15216), .ZN(n15231) );
  NAND2_X1 U18869 ( .A1(n15326), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n15217) );
  AND3_X1 U18870 ( .A1(n15218), .A2(n15327), .A3(n15217), .ZN(n15222) );
  AOI22_X1 U18871 ( .A1(n15320), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12190), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15221) );
  AOI22_X1 U18872 ( .A1(n9732), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(n9727), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15220) );
  AOI22_X1 U18873 ( .A1(n12310), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n15158), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15219) );
  NAND4_X1 U18874 ( .A1(n15222), .A2(n15221), .A3(n15220), .A4(n15219), .ZN(
        n15230) );
  NAND2_X1 U18875 ( .A1(n15326), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n15223) );
  AND3_X1 U18876 ( .A1(n15224), .A2(n15305), .A3(n15223), .ZN(n15228) );
  AOI22_X1 U18877 ( .A1(n15320), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n15323), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15227) );
  AOI22_X1 U18878 ( .A1(n9731), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9727), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15226) );
  AOI22_X1 U18879 ( .A1(n9730), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n15158), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15225) );
  NAND4_X1 U18880 ( .A1(n15228), .A2(n15227), .A3(n15226), .A4(n15225), .ZN(
        n15229) );
  AND2_X1 U18881 ( .A1(n15230), .A2(n15229), .ZN(n15233) );
  NAND2_X1 U18882 ( .A1(n15231), .A2(n15233), .ZN(n15252) );
  OAI211_X1 U18883 ( .C1(n15231), .C2(n15233), .A(n15275), .B(n15252), .ZN(
        n15236) );
  INV_X1 U18884 ( .A(n15236), .ZN(n15232) );
  INV_X1 U18885 ( .A(n15233), .ZN(n15234) );
  NOR2_X1 U18886 ( .A1(n13145), .A2(n15234), .ZN(n16769) );
  NAND2_X1 U18887 ( .A1(n15326), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n15237) );
  AND3_X1 U18888 ( .A1(n15238), .A2(n15327), .A3(n15237), .ZN(n15242) );
  AOI22_X1 U18889 ( .A1(n15320), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n15323), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15241) );
  AOI22_X1 U18890 ( .A1(n9732), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(n9727), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15240) );
  AOI22_X1 U18891 ( .A1(n12310), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n15158), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15239) );
  NAND4_X1 U18892 ( .A1(n15242), .A2(n15241), .A3(n15240), .A4(n15239), .ZN(
        n15250) );
  NAND2_X1 U18893 ( .A1(n15326), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n15243) );
  AND3_X1 U18894 ( .A1(n15244), .A2(n15305), .A3(n15243), .ZN(n15248) );
  AOI22_X1 U18895 ( .A1(n15320), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n15323), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15247) );
  AOI22_X1 U18896 ( .A1(n9732), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9727), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15246) );
  AOI22_X1 U18897 ( .A1(n12310), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n15158), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15245) );
  NAND4_X1 U18898 ( .A1(n15248), .A2(n15247), .A3(n15246), .A4(n15245), .ZN(
        n15249) );
  NAND2_X1 U18899 ( .A1(n15250), .A2(n15249), .ZN(n15254) );
  AOI21_X1 U18900 ( .B1(n15252), .B2(n15254), .A(n15251), .ZN(n15253) );
  INV_X1 U18901 ( .A(n15254), .ZN(n15255) );
  NAND2_X1 U18902 ( .A1(n15209), .A2(n15255), .ZN(n16763) );
  INV_X1 U18903 ( .A(n15274), .ZN(n15276) );
  INV_X1 U18904 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15258) );
  OAI211_X1 U18905 ( .C1(n15259), .C2(n15258), .A(n15257), .B(n15327), .ZN(
        n15260) );
  INV_X1 U18906 ( .A(n15260), .ZN(n15264) );
  AOI22_X1 U18907 ( .A1(n15320), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n15157), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15263) );
  AOI22_X1 U18908 ( .A1(n15326), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9727), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15262) );
  AOI22_X1 U18909 ( .A1(n12310), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n15158), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15261) );
  NAND4_X1 U18910 ( .A1(n15264), .A2(n15263), .A3(n15262), .A4(n15261), .ZN(
        n15272) );
  INV_X1 U18911 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n20879) );
  AOI22_X1 U18912 ( .A1(n15320), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9731), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n15270) );
  AOI22_X1 U18913 ( .A1(n9727), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12190), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15269) );
  NAND2_X1 U18914 ( .A1(n15326), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n15266) );
  NAND2_X1 U18915 ( .A1(n12310), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n15265) );
  AND3_X1 U18916 ( .A1(n15305), .A2(n15266), .A3(n15265), .ZN(n15268) );
  NAND4_X1 U18917 ( .A1(n15270), .A2(n15269), .A3(n15268), .A4(n15267), .ZN(
        n15271) );
  NAND2_X1 U18918 ( .A1(n15272), .A2(n15271), .ZN(n15273) );
  INV_X1 U18919 ( .A(n15273), .ZN(n15281) );
  OR2_X1 U18920 ( .A1(n15274), .A2(n15273), .ZN(n16751) );
  OAI211_X1 U18921 ( .C1(n15276), .C2(n15281), .A(n16751), .B(n15275), .ZN(
        n15279) );
  INV_X1 U18922 ( .A(n15279), .ZN(n15277) );
  NAND2_X1 U18923 ( .A1(n15278), .A2(n15279), .ZN(n15280) );
  NAND2_X1 U18924 ( .A1(n15209), .A2(n15281), .ZN(n16757) );
  INV_X1 U18925 ( .A(n16752), .ZN(n15296) );
  NAND2_X1 U18926 ( .A1(n15326), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n15282) );
  AND3_X1 U18927 ( .A1(n15283), .A2(n15327), .A3(n15282), .ZN(n15287) );
  AOI22_X1 U18928 ( .A1(n15320), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12190), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15286) );
  AOI22_X1 U18929 ( .A1(n15157), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9727), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15285) );
  AOI22_X1 U18930 ( .A1(n12310), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n15158), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15284) );
  NAND4_X1 U18931 ( .A1(n15287), .A2(n15286), .A3(n15285), .A4(n15284), .ZN(
        n15295) );
  NAND2_X1 U18932 ( .A1(n15326), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n15288) );
  AND3_X1 U18933 ( .A1(n15289), .A2(n15305), .A3(n15288), .ZN(n15293) );
  AOI22_X1 U18934 ( .A1(n15320), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n15323), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15292) );
  AOI22_X1 U18935 ( .A1(n9732), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9727), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15291) );
  AOI22_X1 U18936 ( .A1(n12310), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15158), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15290) );
  NAND4_X1 U18937 ( .A1(n15293), .A2(n15292), .A3(n15291), .A4(n15290), .ZN(
        n15294) );
  AND2_X1 U18938 ( .A1(n15295), .A2(n15294), .ZN(n16753) );
  NAND2_X1 U18939 ( .A1(n13145), .A2(n16753), .ZN(n15297) );
  NOR2_X1 U18940 ( .A1(n16751), .A2(n15297), .ZN(n15314) );
  AOI22_X1 U18941 ( .A1(n15320), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n15326), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n15302) );
  AOI22_X1 U18942 ( .A1(n12310), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9727), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n15301) );
  NAND2_X1 U18943 ( .A1(n15158), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n15299) );
  NAND2_X1 U18944 ( .A1(n12190), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n15298) );
  AND3_X1 U18945 ( .A1(n15299), .A2(n15298), .A3(n15327), .ZN(n15300) );
  NAND4_X1 U18946 ( .A1(n15303), .A2(n15302), .A3(n15301), .A4(n15300), .ZN(
        n15312) );
  NAND2_X1 U18947 ( .A1(n9717), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n15306) );
  NAND2_X1 U18948 ( .A1(n15326), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n15304) );
  AND3_X1 U18949 ( .A1(n15306), .A2(n15305), .A3(n15304), .ZN(n15310) );
  AOI22_X1 U18950 ( .A1(n15320), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12190), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n15309) );
  AOI22_X1 U18951 ( .A1(n12310), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9727), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n15308) );
  AOI22_X1 U18952 ( .A1(n9731), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n15158), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n15307) );
  NAND4_X1 U18953 ( .A1(n15310), .A2(n15309), .A3(n15308), .A4(n15307), .ZN(
        n15311) );
  AND2_X1 U18954 ( .A1(n15312), .A2(n15311), .ZN(n15313) );
  NAND2_X1 U18955 ( .A1(n15314), .A2(n15313), .ZN(n15315) );
  OAI21_X1 U18956 ( .B1(n15314), .B2(n15313), .A(n15315), .ZN(n16748) );
  INV_X1 U18957 ( .A(n15315), .ZN(n15316) );
  NOR2_X1 U18958 ( .A1(n16747), .A2(n15316), .ZN(n15336) );
  INV_X1 U18959 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15319) );
  AOI21_X1 U18960 ( .B1(n12190), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n15327), .ZN(n15317) );
  OAI211_X1 U18961 ( .C1(n9722), .C2(n15319), .A(n15318), .B(n15317), .ZN(
        n15334) );
  AOI22_X1 U18962 ( .A1(n15320), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n15326), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15322) );
  AOI22_X1 U18963 ( .A1(n12310), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9727), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n15321) );
  NAND2_X1 U18964 ( .A1(n15322), .A2(n15321), .ZN(n15333) );
  AOI22_X1 U18965 ( .A1(n15320), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n15157), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15325) );
  AOI22_X1 U18966 ( .A1(n9727), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12190), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15324) );
  NAND2_X1 U18967 ( .A1(n15325), .A2(n15324), .ZN(n15332) );
  NAND2_X1 U18968 ( .A1(n15326), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n15329) );
  NAND2_X1 U18969 ( .A1(n15158), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n15328) );
  NAND4_X1 U18970 ( .A1(n15330), .A2(n15329), .A3(n15328), .A4(n15327), .ZN(
        n15331) );
  OAI22_X1 U18971 ( .A1(n15334), .A2(n15333), .B1(n15332), .B2(n15331), .ZN(
        n15335) );
  XNOR2_X1 U18972 ( .A(n15336), .B(n15335), .ZN(n15349) );
  INV_X1 U18973 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n15342) );
  AOI22_X1 U18974 ( .A1(n20360), .A2(n15340), .B1(P2_EAX_REG_30__SCAN_IN), 
        .B2(n16938), .ZN(n15341) );
  OAI21_X1 U18975 ( .B1(n15342), .B2(n16941), .A(n15341), .ZN(n15345) );
  NOR2_X1 U18976 ( .A1(n15343), .A2(n16934), .ZN(n15344) );
  OAI21_X1 U18977 ( .B1(n15349), .B2(n20389), .A(n15346), .ZN(P2_U2889) );
  OAI21_X1 U18978 ( .B1(n15349), .B2(n16840), .A(n15348), .ZN(P2_U2857) );
  AOI21_X1 U18979 ( .B1(n15350), .B2(n14521), .A(n9758), .ZN(n21175) );
  AOI22_X1 U18980 ( .A1(n15697), .A2(n21175), .B1(n15696), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n15351) );
  OAI21_X1 U18981 ( .B1(n21178), .B2(n15702), .A(n15351), .ZN(P1_U2867) );
  NAND2_X1 U18982 ( .A1(n17214), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15353) );
  OAI211_X1 U18983 ( .C1(n17244), .C2(n15355), .A(n15354), .B(n15353), .ZN(
        n15356) );
  INV_X1 U18984 ( .A(n15356), .ZN(n15358) );
  OAI21_X1 U18985 ( .B1(n17218), .B2(n9782), .A(n10684), .ZN(P2_U2984) );
  NAND2_X1 U18986 ( .A1(n9713), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n15360) );
  OAI21_X1 U18987 ( .B1(n15359), .B2(n9713), .A(n15360), .ZN(P2_U2856) );
  NOR2_X1 U18988 ( .A1(n15362), .A2(n20336), .ZN(n15366) );
  NAND2_X1 U18989 ( .A1(n20262), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15364) );
  AOI22_X1 U18990 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n20295), .B1(n20344), 
        .B2(P2_REIP_REG_31__SCAN_IN), .ZN(n15363) );
  NAND2_X1 U18991 ( .A1(n15364), .A2(n15363), .ZN(n15365) );
  OAI21_X1 U18992 ( .B1(n15359), .B2(n20345), .A(n15369), .ZN(P2_U2824) );
  NAND2_X1 U18993 ( .A1(n15370), .A2(n21679), .ZN(n21102) );
  NAND2_X1 U18994 ( .A1(n15371), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n15372)
         );
  NAND3_X1 U18995 ( .A1(n15373), .A2(n21102), .A3(n15372), .ZN(P1_U2801) );
  INV_X1 U18996 ( .A(n15374), .ZN(n15377) );
  INV_X1 U18997 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n15375) );
  NAND2_X1 U18998 ( .A1(n21102), .A2(n15375), .ZN(n15376) );
  MUX2_X1 U18999 ( .A(n15377), .B(n15376), .S(n21820), .Z(P1_U3487) );
  OAI21_X1 U19000 ( .B1(n9780), .B2(n15379), .A(n15378), .ZN(n16022) );
  NAND2_X1 U19001 ( .A1(n15802), .A2(n21168), .ZN(n15390) );
  INV_X1 U19002 ( .A(n15395), .ZN(n15388) );
  NOR2_X1 U19003 ( .A1(n15383), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n15387) );
  INV_X1 U19004 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n15682) );
  INV_X1 U19005 ( .A(n15800), .ZN(n15384) );
  AOI22_X1 U19006 ( .A1(n21146), .A2(n15384), .B1(
        P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n21190), .ZN(n15385) );
  OAI21_X1 U19007 ( .B1(n21205), .B2(n15682), .A(n15385), .ZN(n15386) );
  AOI211_X1 U19008 ( .C1(n15388), .C2(P1_REIP_REG_29__SCAN_IN), .A(n15387), 
        .B(n15386), .ZN(n15389) );
  OAI211_X1 U19009 ( .C1(n16022), .C2(n21143), .A(n15390), .B(n15389), .ZN(
        P1_U2811) );
  INV_X1 U19010 ( .A(n15807), .ZN(n15393) );
  OAI22_X1 U19011 ( .A1(n9710), .A2(n15393), .B1(n15805), .B2(n21203), .ZN(
        n15398) );
  INV_X1 U19012 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n15804) );
  INV_X1 U19013 ( .A(n15394), .ZN(n15396) );
  AOI21_X1 U19014 ( .B1(n15804), .B2(n15396), .A(n15395), .ZN(n15397) );
  AOI211_X1 U19015 ( .C1(n21173), .C2(P1_EBX_REG_28__SCAN_IN), .A(n15398), .B(
        n15397), .ZN(n15401) );
  AOI21_X1 U19016 ( .B1(n15399), .B2(n15405), .A(n9780), .ZN(n15683) );
  NAND2_X1 U19017 ( .A1(n15683), .A2(n21209), .ZN(n15400) );
  OAI211_X1 U19018 ( .C1(n15816), .C2(n15654), .A(n15401), .B(n15400), .ZN(
        P1_U2812) );
  NAND2_X1 U19019 ( .A1(n15402), .A2(n15403), .ZN(n15404) );
  NAND2_X1 U19020 ( .A1(n15405), .A2(n15404), .ZN(n16037) );
  AOI21_X1 U19021 ( .B1(n15407), .B2(n15406), .A(n15391), .ZN(n15823) );
  NAND2_X1 U19022 ( .A1(n15823), .A2(n21168), .ZN(n15415) );
  OAI22_X1 U19023 ( .A1(n9710), .A2(n15821), .B1(n15408), .B2(n21203), .ZN(
        n15413) );
  INV_X1 U19024 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n15409) );
  NAND3_X1 U19025 ( .A1(n21210), .A2(n15410), .A3(n15409), .ZN(n15411) );
  OAI21_X1 U19026 ( .B1(n15684), .B2(n21205), .A(n15411), .ZN(n15412) );
  AOI211_X1 U19027 ( .C1(n15425), .C2(P1_REIP_REG_27__SCAN_IN), .A(n15413), 
        .B(n15412), .ZN(n15414) );
  OAI211_X1 U19028 ( .C1(n21143), .C2(n16037), .A(n15415), .B(n15414), .ZN(
        P1_U2813) );
  OAI21_X1 U19029 ( .B1(n15416), .B2(n15417), .A(n15402), .ZN(n16047) );
  INV_X1 U19030 ( .A(n15418), .ZN(n15432) );
  INV_X1 U19031 ( .A(n15406), .ZN(n15419) );
  AOI21_X1 U19032 ( .B1(n15420), .B2(n15432), .A(n15419), .ZN(n15833) );
  NAND2_X1 U19033 ( .A1(n15833), .A2(n21168), .ZN(n15427) );
  OAI21_X1 U19034 ( .B1(n21126), .B2(n15421), .A(n15829), .ZN(n15424) );
  INV_X1 U19035 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n15685) );
  NOR2_X1 U19036 ( .A1(n21205), .A2(n15685), .ZN(n15423) );
  OAI22_X1 U19037 ( .A1(n9710), .A2(n15831), .B1(n22033), .B2(n21203), .ZN(
        n15422) );
  AOI211_X1 U19038 ( .C1(n15425), .C2(n15424), .A(n15423), .B(n15422), .ZN(
        n15426) );
  OAI211_X1 U19039 ( .C1(n16047), .C2(n21143), .A(n15427), .B(n15426), .ZN(
        P1_U2814) );
  INV_X1 U19040 ( .A(n15416), .ZN(n15429) );
  OAI21_X1 U19041 ( .B1(n15430), .B2(n15428), .A(n15429), .ZN(n16057) );
  AOI21_X1 U19042 ( .B1(n15433), .B2(n15431), .A(n15418), .ZN(n15843) );
  NAND2_X1 U19043 ( .A1(n15843), .A2(n21168), .ZN(n15441) );
  OAI21_X1 U19044 ( .B1(n21126), .B2(n15435), .A(n21123), .ZN(n15445) );
  OAI22_X1 U19045 ( .A1(n9710), .A2(n15841), .B1(n15434), .B2(n21203), .ZN(
        n15439) );
  INV_X1 U19046 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n15686) );
  INV_X1 U19047 ( .A(n15435), .ZN(n15447) );
  OAI21_X1 U19048 ( .B1(n15447), .B2(P1_REIP_REG_25__SCAN_IN), .A(
        P1_REIP_REG_24__SCAN_IN), .ZN(n15436) );
  OAI211_X1 U19049 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(P1_REIP_REG_24__SCAN_IN), .A(n21210), .B(n15436), .ZN(n15437) );
  OAI21_X1 U19050 ( .B1(n15686), .B2(n21205), .A(n15437), .ZN(n15438) );
  AOI211_X1 U19051 ( .C1(n15445), .C2(P1_REIP_REG_25__SCAN_IN), .A(n15439), 
        .B(n15438), .ZN(n15440) );
  OAI211_X1 U19052 ( .C1(n16057), .C2(n21143), .A(n15441), .B(n15440), .ZN(
        P1_U2815) );
  OAI21_X1 U19053 ( .B1(n15442), .B2(n15443), .A(n15431), .ZN(n15849) );
  AOI21_X1 U19054 ( .B1(n15444), .B2(n10662), .A(n15428), .ZN(n16075) );
  INV_X1 U19055 ( .A(n15445), .ZN(n15462) );
  INV_X1 U19056 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n22018) );
  INV_X1 U19057 ( .A(n15852), .ZN(n15446) );
  OAI22_X1 U19058 ( .A1(n9710), .A2(n15446), .B1(n15848), .B2(n21203), .ZN(
        n15449) );
  NOR3_X1 U19059 ( .A1(n21126), .A2(P1_REIP_REG_24__SCAN_IN), .A3(n15447), 
        .ZN(n15448) );
  AOI211_X1 U19060 ( .C1(P1_EBX_REG_24__SCAN_IN), .C2(n21173), .A(n15449), .B(
        n15448), .ZN(n15450) );
  OAI21_X1 U19061 ( .B1(n15462), .B2(n22018), .A(n15450), .ZN(n15451) );
  AOI21_X1 U19062 ( .B1(n16075), .B2(n21209), .A(n15451), .ZN(n15452) );
  OAI21_X1 U19063 ( .B1(n15849), .B2(n15654), .A(n15452), .ZN(P1_U2816) );
  NAND2_X1 U19064 ( .A1(n15453), .A2(n15454), .ZN(n15455) );
  NAND2_X1 U19065 ( .A1(n10662), .A2(n15455), .ZN(n16085) );
  INV_X1 U19066 ( .A(n15442), .ZN(n15456) );
  OAI21_X1 U19067 ( .B1(n15457), .B2(n9786), .A(n15456), .ZN(n15860) );
  INV_X1 U19068 ( .A(n15860), .ZN(n15458) );
  NAND2_X1 U19069 ( .A1(n15458), .A2(n21168), .ZN(n15466) );
  OAI22_X1 U19070 ( .A1(n9710), .A2(n15854), .B1(n15459), .B2(n21203), .ZN(
        n15464) );
  AOI21_X1 U19071 ( .B1(n21210), .B2(n15460), .A(P1_REIP_REG_23__SCAN_IN), 
        .ZN(n15461) );
  NOR2_X1 U19072 ( .A1(n15462), .A2(n15461), .ZN(n15463) );
  AOI211_X1 U19073 ( .C1(P1_EBX_REG_23__SCAN_IN), .C2(n21173), .A(n15464), .B(
        n15463), .ZN(n15465) );
  OAI211_X1 U19074 ( .C1(n16085), .C2(n21143), .A(n15466), .B(n15465), .ZN(
        P1_U2817) );
  OR2_X1 U19075 ( .A1(n15481), .A2(n15467), .ZN(n15468) );
  NAND2_X1 U19076 ( .A1(n15453), .A2(n15468), .ZN(n16101) );
  AOI21_X1 U19077 ( .B1(n15470), .B2(n10631), .A(n9786), .ZN(n15864) );
  NAND2_X1 U19078 ( .A1(n15864), .A2(n21168), .ZN(n15478) );
  OAI21_X1 U19079 ( .B1(n21126), .B2(n15472), .A(n21123), .ZN(n15498) );
  INV_X1 U19080 ( .A(n15867), .ZN(n15471) );
  INV_X1 U19081 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15865) );
  OAI22_X1 U19082 ( .A1(n9710), .A2(n15471), .B1(n15865), .B2(n21203), .ZN(
        n15476) );
  INV_X1 U19083 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n15689) );
  INV_X1 U19084 ( .A(n15472), .ZN(n15484) );
  OAI21_X1 U19085 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(n15484), .A(
        P1_REIP_REG_21__SCAN_IN), .ZN(n15473) );
  OAI211_X1 U19086 ( .C1(P1_REIP_REG_21__SCAN_IN), .C2(P1_REIP_REG_22__SCAN_IN), .A(n21210), .B(n15473), .ZN(n15474) );
  OAI21_X1 U19087 ( .B1(n15689), .B2(n21205), .A(n15474), .ZN(n15475) );
  AOI211_X1 U19088 ( .C1(n15498), .C2(P1_REIP_REG_22__SCAN_IN), .A(n15476), 
        .B(n15475), .ZN(n15477) );
  OAI211_X1 U19089 ( .C1(n16101), .C2(n21143), .A(n15478), .B(n15477), .ZN(
        P1_U2818) );
  AOI21_X1 U19090 ( .B1(n15480), .B2(n15479), .A(n15469), .ZN(n15876) );
  INV_X1 U19091 ( .A(n15876), .ZN(n15752) );
  AOI21_X1 U19092 ( .B1(n15482), .B2(n15496), .A(n15481), .ZN(n16110) );
  INV_X1 U19093 ( .A(n15498), .ZN(n15489) );
  INV_X1 U19094 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n15488) );
  OAI22_X1 U19095 ( .A1(n9710), .A2(n15874), .B1(n15483), .B2(n21203), .ZN(
        n15486) );
  NOR3_X1 U19096 ( .A1(n21126), .A2(P1_REIP_REG_21__SCAN_IN), .A3(n15484), 
        .ZN(n15485) );
  AOI211_X1 U19097 ( .C1(P1_EBX_REG_21__SCAN_IN), .C2(n21173), .A(n15486), .B(
        n15485), .ZN(n15487) );
  OAI21_X1 U19098 ( .B1(n15489), .B2(n15488), .A(n15487), .ZN(n15490) );
  AOI21_X1 U19099 ( .B1(n16110), .B2(n21209), .A(n15490), .ZN(n15491) );
  OAI21_X1 U19100 ( .B1(n15752), .B2(n15654), .A(n15491), .ZN(P1_U2819) );
  OAI21_X1 U19101 ( .B1(n15492), .B2(n15493), .A(n15479), .ZN(n15881) );
  NAND2_X1 U19102 ( .A1(n15508), .A2(n15494), .ZN(n15495) );
  NAND2_X1 U19103 ( .A1(n15496), .A2(n15495), .ZN(n15692) );
  INV_X1 U19104 ( .A(n15692), .ZN(n16119) );
  NOR2_X1 U19105 ( .A1(n21126), .A2(n15497), .ZN(n15499) );
  OAI21_X1 U19106 ( .B1(n15499), .B2(P1_REIP_REG_20__SCAN_IN), .A(n15498), 
        .ZN(n15501) );
  AOI22_X1 U19107 ( .A1(n21146), .A2(n15884), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n21190), .ZN(n15500) );
  OAI211_X1 U19108 ( .C1(n15691), .C2(n21205), .A(n15501), .B(n15500), .ZN(
        n15502) );
  AOI21_X1 U19109 ( .B1(n16119), .B2(n21209), .A(n15502), .ZN(n15503) );
  OAI21_X1 U19110 ( .B1(n15881), .B2(n15654), .A(n15503), .ZN(P1_U2820) );
  AOI21_X1 U19111 ( .B1(n15505), .B2(n15504), .A(n15492), .ZN(n15894) );
  INV_X1 U19112 ( .A(n15506), .ZN(n15510) );
  INV_X1 U19113 ( .A(n15507), .ZN(n15509) );
  OAI21_X1 U19114 ( .B1(n15510), .B2(n15509), .A(n15508), .ZN(n16122) );
  INV_X1 U19115 ( .A(n21291), .ZN(n21189) );
  AOI21_X1 U19116 ( .B1(n21190), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n21189), .ZN(n15511) );
  OAI21_X1 U19117 ( .B1(n9710), .B2(n15892), .A(n15511), .ZN(n15514) );
  NAND2_X1 U19118 ( .A1(n21210), .A2(n15515), .ZN(n15603) );
  NOR3_X1 U19119 ( .A1(n15603), .A2(P1_REIP_REG_19__SCAN_IN), .A3(n15512), 
        .ZN(n15513) );
  AOI211_X1 U19120 ( .C1(P1_EBX_REG_19__SCAN_IN), .C2(n21173), .A(n15514), .B(
        n15513), .ZN(n15523) );
  INV_X1 U19121 ( .A(n15515), .ZN(n15516) );
  NAND2_X1 U19122 ( .A1(n21210), .A2(n15516), .ZN(n15517) );
  AND2_X1 U19123 ( .A1(n15517), .A2(n21123), .ZN(n15615) );
  INV_X1 U19124 ( .A(n15520), .ZN(n15518) );
  NAND2_X1 U19125 ( .A1(n15628), .A2(n15518), .ZN(n15519) );
  NAND2_X1 U19126 ( .A1(n15615), .A2(n15519), .ZN(n15541) );
  INV_X1 U19127 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n21771) );
  NAND2_X1 U19128 ( .A1(n21771), .A2(n15520), .ZN(n15521) );
  NOR2_X1 U19129 ( .A1(n15603), .A2(n15521), .ZN(n15534) );
  OAI21_X1 U19130 ( .B1(n15541), .B2(n15534), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n15522) );
  OAI211_X1 U19131 ( .C1(n16122), .C2(n21143), .A(n15523), .B(n15522), .ZN(
        n15524) );
  AOI21_X1 U19132 ( .B1(n15894), .B2(n21168), .A(n15524), .ZN(n15525) );
  INV_X1 U19133 ( .A(n15525), .ZN(P1_U2821) );
  OAI21_X1 U19134 ( .B1(n15526), .B2(n15527), .A(n15506), .ZN(n16132) );
  XNOR2_X1 U19135 ( .A(n15528), .B(n15529), .ZN(n15903) );
  INV_X1 U19136 ( .A(n15903), .ZN(n15530) );
  NAND2_X1 U19137 ( .A1(n15530), .A2(n21168), .ZN(n15536) );
  INV_X1 U19138 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n15693) );
  INV_X1 U19139 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15896) );
  OAI21_X1 U19140 ( .B1(n21203), .B2(n15896), .A(n21291), .ZN(n15531) );
  AOI21_X1 U19141 ( .B1(n21146), .B2(n15901), .A(n15531), .ZN(n15532) );
  OAI21_X1 U19142 ( .B1(n21205), .B2(n15693), .A(n15532), .ZN(n15533) );
  AOI211_X1 U19143 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(n15541), .A(n15534), 
        .B(n15533), .ZN(n15535) );
  OAI211_X1 U19144 ( .C1(n16132), .C2(n21143), .A(n15536), .B(n15535), .ZN(
        P1_U2822) );
  OAI21_X1 U19145 ( .B1(n15537), .B2(n15538), .A(n15528), .ZN(n15913) );
  NOR2_X1 U19146 ( .A1(n15553), .A2(n15539), .ZN(n15540) );
  OR2_X1 U19147 ( .A1(n15526), .A2(n15540), .ZN(n16150) );
  INV_X1 U19148 ( .A(n16150), .ZN(n15547) );
  INV_X1 U19149 ( .A(n15603), .ZN(n15586) );
  NAND3_X1 U19150 ( .A1(n15586), .A2(P1_REIP_REG_13__SCAN_IN), .A3(
        P1_REIP_REG_14__SCAN_IN), .ZN(n15575) );
  NOR2_X1 U19151 ( .A1(n15575), .A2(n15558), .ZN(n15542) );
  OAI21_X1 U19152 ( .B1(n15542), .B2(P1_REIP_REG_17__SCAN_IN), .A(n15541), 
        .ZN(n15545) );
  OAI21_X1 U19153 ( .B1(n21203), .B2(n22100), .A(n21291), .ZN(n15543) );
  AOI21_X1 U19154 ( .B1(n21146), .B2(n15912), .A(n15543), .ZN(n15544) );
  OAI211_X1 U19155 ( .C1(n15694), .C2(n21205), .A(n15545), .B(n15544), .ZN(
        n15546) );
  AOI21_X1 U19156 ( .B1(n15547), .B2(n21209), .A(n15546), .ZN(n15548) );
  OAI21_X1 U19157 ( .B1(n15913), .B2(n15654), .A(n15548), .ZN(P1_U2823) );
  AOI21_X1 U19158 ( .B1(n15550), .B2(n15549), .A(n15537), .ZN(n15925) );
  INV_X1 U19159 ( .A(n15925), .ZN(n15779) );
  AND2_X1 U19160 ( .A1(n15571), .A2(n15551), .ZN(n15552) );
  NOR2_X1 U19161 ( .A1(n15553), .A2(n15552), .ZN(n16165) );
  INV_X1 U19162 ( .A(n15615), .ZN(n15554) );
  AOI21_X1 U19163 ( .B1(n15555), .B2(n15628), .A(n15554), .ZN(n15588) );
  INV_X1 U19164 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n15562) );
  NAND2_X1 U19165 ( .A1(n21146), .A2(n15921), .ZN(n15556) );
  OAI211_X1 U19166 ( .C1(n21203), .C2(n15923), .A(n15556), .B(n21291), .ZN(
        n15557) );
  AOI21_X1 U19167 ( .B1(n21173), .B2(P1_EBX_REG_16__SCAN_IN), .A(n15557), .ZN(
        n15561) );
  INV_X1 U19168 ( .A(n15575), .ZN(n15559) );
  OAI211_X1 U19169 ( .C1(P1_REIP_REG_16__SCAN_IN), .C2(P1_REIP_REG_15__SCAN_IN), .A(n15559), .B(n15558), .ZN(n15560) );
  OAI211_X1 U19170 ( .C1(n15588), .C2(n15562), .A(n15561), .B(n15560), .ZN(
        n15563) );
  AOI21_X1 U19171 ( .B1(n21209), .B2(n16165), .A(n15563), .ZN(n15564) );
  OAI21_X1 U19172 ( .B1(n15779), .B2(n15654), .A(n15564), .ZN(P1_U2824) );
  INV_X1 U19173 ( .A(n15595), .ZN(n15625) );
  INV_X1 U19174 ( .A(n15565), .ZN(n15593) );
  INV_X1 U19175 ( .A(n15594), .ZN(n15566) );
  OAI21_X1 U19176 ( .B1(n15625), .B2(n14879), .A(n15566), .ZN(n15567) );
  NAND3_X1 U19177 ( .A1(n15567), .A2(n15598), .A3(n15596), .ZN(n15597) );
  INV_X1 U19178 ( .A(n15568), .ZN(n15584) );
  NOR2_X1 U19179 ( .A1(n15597), .A2(n15584), .ZN(n15583) );
  OAI21_X1 U19180 ( .B1(n15583), .B2(n15569), .A(n15549), .ZN(n15938) );
  INV_X1 U19181 ( .A(n15571), .ZN(n15572) );
  AOI21_X1 U19182 ( .B1(n15573), .B2(n15570), .A(n15572), .ZN(n16172) );
  INV_X1 U19183 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n21860) );
  AOI21_X1 U19184 ( .B1(n21190), .B2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n21189), .ZN(n15574) );
  OAI21_X1 U19185 ( .B1(n9710), .B2(n15934), .A(n15574), .ZN(n15577) );
  NOR2_X1 U19186 ( .A1(n15575), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n15576) );
  AOI211_X1 U19187 ( .C1(P1_EBX_REG_15__SCAN_IN), .C2(n21173), .A(n15577), .B(
        n15576), .ZN(n15578) );
  OAI21_X1 U19188 ( .B1(n15588), .B2(n21860), .A(n15578), .ZN(n15579) );
  AOI21_X1 U19189 ( .B1(n21209), .B2(n16172), .A(n15579), .ZN(n15580) );
  OAI21_X1 U19190 ( .B1(n15938), .B2(n15654), .A(n15580), .ZN(P1_U2825) );
  OR2_X1 U19191 ( .A1(n15601), .A2(n15581), .ZN(n15582) );
  NAND2_X1 U19192 ( .A1(n15570), .A2(n15582), .ZN(n16180) );
  AOI21_X1 U19193 ( .B1(n15584), .B2(n15597), .A(n15583), .ZN(n15948) );
  NAND2_X1 U19194 ( .A1(n15948), .A2(n21168), .ZN(n15592) );
  NAND2_X1 U19195 ( .A1(n21190), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15585) );
  OAI211_X1 U19196 ( .C1(n9710), .C2(n15946), .A(n21291), .B(n15585), .ZN(
        n15590) );
  AOI21_X1 U19197 ( .B1(n15586), .B2(P1_REIP_REG_13__SCAN_IN), .A(
        P1_REIP_REG_14__SCAN_IN), .ZN(n15587) );
  NOR2_X1 U19198 ( .A1(n15588), .A2(n15587), .ZN(n15589) );
  AOI211_X1 U19199 ( .C1(P1_EBX_REG_14__SCAN_IN), .C2(n21173), .A(n15590), .B(
        n15589), .ZN(n15591) );
  OAI211_X1 U19200 ( .C1(n16180), .C2(n21143), .A(n15592), .B(n15591), .ZN(
        P1_U2826) );
  AOI21_X1 U19201 ( .B1(n15593), .B2(n14879), .A(n15594), .ZN(n15626) );
  AOI21_X1 U19202 ( .B1(n15626), .B2(n15595), .A(n15594), .ZN(n15611) );
  INV_X1 U19203 ( .A(n15596), .ZN(n15610) );
  NOR2_X1 U19204 ( .A1(n15611), .A2(n15610), .ZN(n15609) );
  OAI21_X1 U19205 ( .B1(n15609), .B2(n15598), .A(n15597), .ZN(n15962) );
  NOR2_X1 U19206 ( .A1(n15617), .A2(n15599), .ZN(n15600) );
  OR2_X1 U19207 ( .A1(n15601), .A2(n15600), .ZN(n15700) );
  INV_X1 U19208 ( .A(n15700), .ZN(n16189) );
  INV_X1 U19209 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n22109) );
  AOI21_X1 U19210 ( .B1(n21190), .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n21189), .ZN(n15602) );
  OAI21_X1 U19211 ( .B1(n9710), .B2(n15950), .A(n15602), .ZN(n15605) );
  NOR2_X1 U19212 ( .A1(n15603), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n15604) );
  AOI211_X1 U19213 ( .C1(P1_EBX_REG_13__SCAN_IN), .C2(n21173), .A(n15605), .B(
        n15604), .ZN(n15606) );
  OAI21_X1 U19214 ( .B1(n15615), .B2(n22109), .A(n15606), .ZN(n15607) );
  AOI21_X1 U19215 ( .B1(n21209), .B2(n16189), .A(n15607), .ZN(n15608) );
  OAI21_X1 U19216 ( .B1(n15962), .B2(n15654), .A(n15608), .ZN(P1_U2827) );
  AOI21_X1 U19217 ( .B1(n15611), .B2(n15610), .A(n15609), .ZN(n15612) );
  INV_X1 U19218 ( .A(n15612), .ZN(n15970) );
  AOI21_X1 U19219 ( .B1(n21210), .B2(n15613), .A(P1_REIP_REG_12__SCAN_IN), 
        .ZN(n15614) );
  NOR2_X1 U19220 ( .A1(n15615), .A2(n15614), .ZN(n15623) );
  AND2_X1 U19221 ( .A1(n15633), .A2(n15616), .ZN(n15618) );
  OR2_X1 U19222 ( .A1(n15618), .A2(n15617), .ZN(n16197) );
  NOR2_X1 U19223 ( .A1(n16197), .A2(n21143), .ZN(n15622) );
  INV_X1 U19224 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n15701) );
  NOR2_X1 U19225 ( .A1(n21205), .A2(n15701), .ZN(n15621) );
  NAND2_X1 U19226 ( .A1(n21190), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15619) );
  OAI211_X1 U19227 ( .C1(n9710), .C2(n15963), .A(n21291), .B(n15619), .ZN(
        n15620) );
  NOR4_X1 U19228 ( .A1(n15623), .A2(n15622), .A3(n15621), .A4(n15620), .ZN(
        n15624) );
  OAI21_X1 U19229 ( .B1(n15970), .B2(n15654), .A(n15624), .ZN(P1_U2828) );
  XNOR2_X1 U19230 ( .A(n15626), .B(n15625), .ZN(n15976) );
  OR2_X1 U19231 ( .A1(n21200), .A2(n15645), .ZN(n15627) );
  NAND2_X1 U19232 ( .A1(n15628), .A2(n15627), .ZN(n15643) );
  INV_X1 U19233 ( .A(n15643), .ZN(n15640) );
  INV_X1 U19234 ( .A(n15629), .ZN(n15632) );
  INV_X1 U19235 ( .A(n15630), .ZN(n15631) );
  OAI21_X1 U19236 ( .B1(n14875), .B2(n15632), .A(n15631), .ZN(n15634) );
  NAND2_X1 U19237 ( .A1(n15634), .A2(n15633), .ZN(n16220) );
  AOI21_X1 U19238 ( .B1(n21190), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n21189), .ZN(n15635) );
  OAI21_X1 U19239 ( .B1(n9710), .B2(n15974), .A(n15635), .ZN(n15637) );
  NOR3_X1 U19240 ( .A1(n21126), .A2(P1_REIP_REG_11__SCAN_IN), .A3(n15645), 
        .ZN(n15636) );
  AOI211_X1 U19241 ( .C1(P1_EBX_REG_11__SCAN_IN), .C2(n21173), .A(n15637), .B(
        n15636), .ZN(n15638) );
  OAI21_X1 U19242 ( .B1(n21143), .B2(n16220), .A(n15638), .ZN(n15639) );
  AOI21_X1 U19243 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n15640), .A(n15639), 
        .ZN(n15641) );
  OAI21_X1 U19244 ( .B1(n15794), .B2(n15654), .A(n15641), .ZN(P1_U2829) );
  AOI22_X1 U19245 ( .A1(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n21190), .B1(
        n21209), .B2(n16233), .ZN(n15642) );
  OAI211_X1 U19246 ( .C1(n15643), .C2(n15984), .A(n15642), .B(n21291), .ZN(
        n15649) );
  AOI22_X1 U19247 ( .A1(n15987), .A2(n21146), .B1(n21173), .B2(
        P1_EBX_REG_10__SCAN_IN), .ZN(n15647) );
  NAND3_X1 U19248 ( .A1(n21210), .A2(n15645), .A3(n15644), .ZN(n15646) );
  NAND2_X1 U19249 ( .A1(n15647), .A2(n15646), .ZN(n15648) );
  NOR2_X1 U19250 ( .A1(n15649), .A2(n15648), .ZN(n15650) );
  OAI21_X1 U19251 ( .B1(n15654), .B2(n15990), .A(n15650), .ZN(P1_U2830) );
  INV_X1 U19252 ( .A(n21820), .ZN(n15652) );
  NAND2_X1 U19253 ( .A1(n15652), .A2(n15651), .ZN(n15653) );
  INV_X1 U19254 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n21201) );
  AND3_X1 U19255 ( .A1(n21210), .A2(n21201), .A3(P1_REIP_REG_1__SCAN_IN), .ZN(
        n15664) );
  INV_X1 U19256 ( .A(n15655), .ZN(n15656) );
  NAND2_X1 U19257 ( .A1(n21209), .A2(n15656), .ZN(n15661) );
  NOR2_X1 U19258 ( .A1(n21820), .A2(n11806), .ZN(n21207) );
  AOI21_X1 U19259 ( .B1(n21210), .B2(n21806), .A(n21200), .ZN(n15657) );
  OAI22_X1 U19260 ( .A1(n21203), .A2(n15658), .B1(n21201), .B2(n15657), .ZN(
        n15659) );
  AOI21_X1 U19261 ( .B1(n21309), .B2(n21207), .A(n15659), .ZN(n15660) );
  OAI211_X1 U19262 ( .C1(n9710), .C2(n15662), .A(n15661), .B(n15660), .ZN(
        n15663) );
  AOI211_X1 U19263 ( .C1(P1_EBX_REG_2__SCAN_IN), .C2(n21173), .A(n15664), .B(
        n15663), .ZN(n15665) );
  OAI21_X1 U19264 ( .B1(n15666), .B2(n21215), .A(n15665), .ZN(P1_U2838) );
  AOI22_X1 U19265 ( .A1(n21190), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n21200), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n15668) );
  NAND2_X1 U19266 ( .A1(n21207), .A2(n21564), .ZN(n15667) );
  OAI211_X1 U19267 ( .C1(n9710), .C2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n15668), .B(n15667), .ZN(n15670) );
  OAI22_X1 U19268 ( .A1(n21126), .A2(P1_REIP_REG_1__SCAN_IN), .B1(n14240), 
        .B2(n21205), .ZN(n15669) );
  AOI211_X1 U19269 ( .C1(n21209), .C2(n15671), .A(n15670), .B(n15669), .ZN(
        n15672) );
  OAI21_X1 U19270 ( .B1(n21215), .B2(n15673), .A(n15672), .ZN(P1_U2839) );
  OAI22_X1 U19271 ( .A1(n15675), .A2(n21812), .B1(n21143), .B2(n15674), .ZN(
        n15678) );
  INV_X1 U19272 ( .A(n21207), .ZN(n21184) );
  NOR2_X1 U19273 ( .A1(n21184), .A2(n15676), .ZN(n15677) );
  AOI211_X1 U19274 ( .C1(n21173), .C2(P1_EBX_REG_0__SCAN_IN), .A(n15678), .B(
        n15677), .ZN(n15680) );
  OAI21_X1 U19275 ( .B1(n21146), .B2(n21190), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15679) );
  OAI211_X1 U19276 ( .C1(n21215), .C2(n15681), .A(n15680), .B(n15679), .ZN(
        P1_U2840) );
  OAI22_X1 U19277 ( .A1(n11797), .A2(n15704), .B1(n11675), .B2(n15709), .ZN(
        P1_U2841) );
  INV_X1 U19278 ( .A(n15802), .ZN(n15714) );
  OAI222_X1 U19279 ( .A1(n15682), .A2(n15709), .B1(n15704), .B2(n16022), .C1(
        n15714), .C2(n15702), .ZN(P1_U2843) );
  INV_X1 U19280 ( .A(n15683), .ZN(n16036) );
  INV_X1 U19281 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n21984) );
  OAI222_X1 U19282 ( .A1(n16036), .A2(n15704), .B1(n21984), .B2(n15709), .C1(
        n15816), .C2(n15702), .ZN(P1_U2844) );
  INV_X1 U19283 ( .A(n15823), .ZN(n15722) );
  OAI222_X1 U19284 ( .A1(n15684), .A2(n15709), .B1(n15704), .B2(n16037), .C1(
        n15722), .C2(n15702), .ZN(P1_U2845) );
  INV_X1 U19285 ( .A(n15833), .ZN(n15727) );
  OAI222_X1 U19286 ( .A1(n16047), .A2(n15704), .B1(n15685), .B2(n15709), .C1(
        n15727), .C2(n15702), .ZN(P1_U2846) );
  INV_X1 U19287 ( .A(n15843), .ZN(n15733) );
  OAI222_X1 U19288 ( .A1(n16057), .A2(n15704), .B1(n15686), .B2(n15709), .C1(
        n15733), .C2(n15702), .ZN(P1_U2847) );
  AOI22_X1 U19289 ( .A1(n16075), .A2(n15697), .B1(n15696), .B2(
        P1_EBX_REG_24__SCAN_IN), .ZN(n15687) );
  OAI21_X1 U19290 ( .B1(n15849), .B2(n15702), .A(n15687), .ZN(P1_U2848) );
  INV_X1 U19291 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n15688) );
  OAI222_X1 U19292 ( .A1(n16085), .A2(n15704), .B1(n15688), .B2(n15709), .C1(
        n15860), .C2(n15702), .ZN(P1_U2849) );
  INV_X1 U19293 ( .A(n15864), .ZN(n15747) );
  OAI222_X1 U19294 ( .A1(n16101), .A2(n15704), .B1(n15689), .B2(n15709), .C1(
        n15747), .C2(n15702), .ZN(P1_U2850) );
  AOI22_X1 U19295 ( .A1(n16110), .A2(n15697), .B1(n15696), .B2(
        P1_EBX_REG_21__SCAN_IN), .ZN(n15690) );
  OAI21_X1 U19296 ( .B1(n15752), .B2(n15702), .A(n15690), .ZN(P1_U2851) );
  OAI222_X1 U19297 ( .A1(n15692), .A2(n15704), .B1(n15691), .B2(n15709), .C1(
        n15881), .C2(n15702), .ZN(P1_U2852) );
  INV_X1 U19298 ( .A(n15894), .ZN(n15761) );
  OAI222_X1 U19299 ( .A1(n16122), .A2(n15704), .B1(n22099), .B2(n15709), .C1(
        n15761), .C2(n15702), .ZN(P1_U2853) );
  OAI222_X1 U19300 ( .A1(n16132), .A2(n15704), .B1(n15693), .B2(n15709), .C1(
        n15702), .C2(n15903), .ZN(P1_U2854) );
  OAI222_X1 U19301 ( .A1(n16150), .A2(n15704), .B1(n15694), .B2(n15709), .C1(
        n15913), .C2(n15702), .ZN(P1_U2855) );
  AOI22_X1 U19302 ( .A1(n16165), .A2(n15697), .B1(n15696), .B2(
        P1_EBX_REG_16__SCAN_IN), .ZN(n15695) );
  OAI21_X1 U19303 ( .B1(n15779), .B2(n15702), .A(n15695), .ZN(P1_U2856) );
  AOI22_X1 U19304 ( .A1(n16172), .A2(n15697), .B1(n15696), .B2(
        P1_EBX_REG_15__SCAN_IN), .ZN(n15698) );
  OAI21_X1 U19305 ( .B1(n15938), .B2(n15702), .A(n15698), .ZN(P1_U2857) );
  INV_X1 U19306 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n22110) );
  INV_X1 U19307 ( .A(n15948), .ZN(n15783) );
  OAI222_X1 U19308 ( .A1(n16180), .A2(n15704), .B1(n22110), .B2(n15709), .C1(
        n15783), .C2(n15702), .ZN(P1_U2858) );
  OAI222_X1 U19309 ( .A1(n15700), .A2(n15704), .B1(n15699), .B2(n15709), .C1(
        n15962), .C2(n15702), .ZN(P1_U2859) );
  OAI222_X1 U19310 ( .A1(n16197), .A2(n15704), .B1(n15701), .B2(n15709), .C1(
        n15970), .C2(n15702), .ZN(P1_U2860) );
  OAI222_X1 U19311 ( .A1(n16220), .A2(n15704), .B1(n15703), .B2(n15709), .C1(
        n15794), .C2(n15702), .ZN(P1_U2861) );
  OR2_X1 U19312 ( .A1(n14841), .A2(n15705), .ZN(n15706) );
  NAND2_X1 U19313 ( .A1(n14876), .A2(n15706), .ZN(n21142) );
  INV_X1 U19314 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n15708) );
  OAI222_X1 U19315 ( .A1(n21142), .A2(n15704), .B1(n15709), .B2(n15708), .C1(
        n15702), .C2(n15707), .ZN(P1_U2864) );
  OAI22_X1 U19316 ( .A1(n15768), .A2(n15785), .B1(n15710), .B2(n15781), .ZN(
        n15711) );
  AOI21_X1 U19317 ( .B1(BUF1_REG_29__SCAN_IN), .B2(n15770), .A(n15711), .ZN(
        n15713) );
  NAND2_X1 U19318 ( .A1(n13436), .A2(DATAI_29_), .ZN(n15712) );
  OAI211_X1 U19319 ( .C1(n15714), .C2(n15790), .A(n15713), .B(n15712), .ZN(
        P1_U2875) );
  OAI22_X1 U19320 ( .A1(n15768), .A2(n15789), .B1(n15715), .B2(n15781), .ZN(
        n15716) );
  AOI21_X1 U19321 ( .B1(BUF1_REG_28__SCAN_IN), .B2(n15770), .A(n15716), .ZN(
        n15718) );
  NAND2_X1 U19322 ( .A1(n13436), .A2(DATAI_28_), .ZN(n15717) );
  OAI211_X1 U19323 ( .C1(n15816), .C2(n15790), .A(n15718), .B(n15717), .ZN(
        P1_U2876) );
  INV_X1 U19324 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n18153) );
  INV_X1 U19325 ( .A(n15768), .ZN(n15774) );
  AOI22_X1 U19326 ( .A1(n15774), .A2(n15791), .B1(P1_EAX_REG_27__SCAN_IN), 
        .B2(n13423), .ZN(n15719) );
  OAI21_X1 U19327 ( .B1(n18153), .B2(n15776), .A(n15719), .ZN(n15720) );
  AOI21_X1 U19328 ( .B1(n13436), .B2(DATAI_27_), .A(n15720), .ZN(n15721) );
  OAI21_X1 U19329 ( .B1(n15722), .B2(n15790), .A(n15721), .ZN(P1_U2877) );
  OAI22_X1 U19330 ( .A1(n15768), .A2(n15723), .B1(n14316), .B2(n15781), .ZN(
        n15724) );
  AOI21_X1 U19331 ( .B1(n15770), .B2(BUF1_REG_26__SCAN_IN), .A(n15724), .ZN(
        n15726) );
  NAND2_X1 U19332 ( .A1(n13436), .A2(DATAI_26_), .ZN(n15725) );
  OAI211_X1 U19333 ( .C1(n15727), .C2(n15790), .A(n15726), .B(n15725), .ZN(
        P1_U2878) );
  OAI22_X1 U19334 ( .A1(n15768), .A2(n15729), .B1(n15728), .B2(n15781), .ZN(
        n15730) );
  AOI21_X1 U19335 ( .B1(n15770), .B2(BUF1_REG_25__SCAN_IN), .A(n15730), .ZN(
        n15732) );
  NAND2_X1 U19336 ( .A1(n13436), .A2(DATAI_25_), .ZN(n15731) );
  OAI211_X1 U19337 ( .C1(n15733), .C2(n15790), .A(n15732), .B(n15731), .ZN(
        P1_U2879) );
  OAI22_X1 U19338 ( .A1(n15768), .A2(n15735), .B1(n15734), .B2(n15781), .ZN(
        n15736) );
  AOI21_X1 U19339 ( .B1(n15770), .B2(BUF1_REG_24__SCAN_IN), .A(n15736), .ZN(
        n15738) );
  NAND2_X1 U19340 ( .A1(n13436), .A2(DATAI_24_), .ZN(n15737) );
  OAI211_X1 U19341 ( .C1(n15849), .C2(n15790), .A(n15738), .B(n15737), .ZN(
        P1_U2880) );
  OAI22_X1 U19342 ( .A1(n15768), .A2(n15739), .B1(n13762), .B2(n15781), .ZN(
        n15740) );
  AOI21_X1 U19343 ( .B1(n15770), .B2(BUF1_REG_23__SCAN_IN), .A(n15740), .ZN(
        n15742) );
  NAND2_X1 U19344 ( .A1(n13436), .A2(DATAI_23_), .ZN(n15741) );
  OAI211_X1 U19345 ( .C1(n15860), .C2(n15790), .A(n15742), .B(n15741), .ZN(
        P1_U2881) );
  OAI22_X1 U19346 ( .A1(n15768), .A2(n15743), .B1(n13768), .B2(n15781), .ZN(
        n15744) );
  AOI21_X1 U19347 ( .B1(n15770), .B2(BUF1_REG_22__SCAN_IN), .A(n15744), .ZN(
        n15746) );
  NAND2_X1 U19348 ( .A1(n13436), .A2(DATAI_22_), .ZN(n15745) );
  OAI211_X1 U19349 ( .C1(n15747), .C2(n15790), .A(n15746), .B(n15745), .ZN(
        P1_U2882) );
  OAI22_X1 U19350 ( .A1(n15768), .A2(n15748), .B1(n13758), .B2(n15781), .ZN(
        n15749) );
  AOI21_X1 U19351 ( .B1(n15770), .B2(BUF1_REG_21__SCAN_IN), .A(n15749), .ZN(
        n15751) );
  NAND2_X1 U19352 ( .A1(n13436), .A2(DATAI_21_), .ZN(n15750) );
  OAI211_X1 U19353 ( .C1(n15752), .C2(n15790), .A(n15751), .B(n15750), .ZN(
        P1_U2883) );
  OAI22_X1 U19354 ( .A1(n15768), .A2(n15753), .B1(n13756), .B2(n15781), .ZN(
        n15754) );
  AOI21_X1 U19355 ( .B1(n15770), .B2(BUF1_REG_20__SCAN_IN), .A(n15754), .ZN(
        n15756) );
  NAND2_X1 U19356 ( .A1(n13436), .A2(DATAI_20_), .ZN(n15755) );
  OAI211_X1 U19357 ( .C1(n15881), .C2(n15790), .A(n15756), .B(n15755), .ZN(
        P1_U2884) );
  OAI22_X1 U19358 ( .A1(n15768), .A2(n15757), .B1(n13764), .B2(n15781), .ZN(
        n15758) );
  AOI21_X1 U19359 ( .B1(n15770), .B2(BUF1_REG_19__SCAN_IN), .A(n15758), .ZN(
        n15760) );
  NAND2_X1 U19360 ( .A1(n13436), .A2(DATAI_19_), .ZN(n15759) );
  OAI211_X1 U19361 ( .C1(n15761), .C2(n15790), .A(n15760), .B(n15759), .ZN(
        P1_U2885) );
  INV_X1 U19362 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n18168) );
  AOI22_X1 U19363 ( .A1(n15774), .A2(n15762), .B1(P1_EAX_REG_18__SCAN_IN), 
        .B2(n13423), .ZN(n15763) );
  OAI21_X1 U19364 ( .B1(n15776), .B2(n18168), .A(n15763), .ZN(n15764) );
  AOI21_X1 U19365 ( .B1(n13436), .B2(DATAI_18_), .A(n15764), .ZN(n15765) );
  OAI21_X1 U19366 ( .B1(n15903), .B2(n15790), .A(n15765), .ZN(P1_U2886) );
  INV_X1 U19367 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n15766) );
  OAI22_X1 U19368 ( .A1(n15768), .A2(n15767), .B1(n15766), .B2(n15781), .ZN(
        n15769) );
  AOI21_X1 U19369 ( .B1(n15770), .B2(BUF1_REG_17__SCAN_IN), .A(n15769), .ZN(
        n15772) );
  NAND2_X1 U19370 ( .A1(n13436), .A2(DATAI_17_), .ZN(n15771) );
  OAI211_X1 U19371 ( .C1(n15913), .C2(n15790), .A(n15772), .B(n15771), .ZN(
        P1_U2887) );
  AOI22_X1 U19372 ( .A1(n15774), .A2(n15773), .B1(P1_EAX_REG_16__SCAN_IN), 
        .B2(n13423), .ZN(n15775) );
  OAI21_X1 U19373 ( .B1(n15776), .B2(n18171), .A(n15775), .ZN(n15777) );
  AOI21_X1 U19374 ( .B1(n13436), .B2(DATAI_16_), .A(n15777), .ZN(n15778) );
  OAI21_X1 U19375 ( .B1(n15779), .B2(n15790), .A(n15778), .ZN(P1_U2888) );
  OAI222_X1 U19376 ( .A1(n15938), .A2(n15790), .B1(n15788), .B2(n15780), .C1(
        n21228), .C2(n15786), .ZN(P1_U2889) );
  INV_X1 U19377 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n15782) );
  OAI222_X1 U19378 ( .A1(n15783), .A2(n15790), .B1(n21258), .B2(n15788), .C1(
        n15782), .C2(n15781), .ZN(P1_U2890) );
  INV_X1 U19379 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n15784) );
  OAI222_X1 U19380 ( .A1(n15962), .A2(n15790), .B1(n15785), .B2(n15788), .C1(
        n15784), .C2(n15786), .ZN(P1_U2891) );
  INV_X1 U19381 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n15787) );
  OAI222_X1 U19382 ( .A1(n15970), .A2(n15790), .B1(n15789), .B2(n15788), .C1(
        n15787), .C2(n15786), .ZN(P1_U2892) );
  AOI22_X1 U19383 ( .A1(n15792), .A2(n15791), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n13423), .ZN(n15793) );
  OAI21_X1 U19384 ( .B1(n15794), .B2(n15790), .A(n15793), .ZN(P1_U2893) );
  NOR2_X1 U19385 ( .A1(n15796), .A2(n10667), .ZN(n15797) );
  XNOR2_X1 U19386 ( .A(n15795), .B(n15797), .ZN(n16026) );
  NOR2_X1 U19387 ( .A1(n21291), .A2(n15798), .ZN(n16020) );
  AOI21_X1 U19388 ( .B1(n18048), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n16020), .ZN(n15799) );
  OAI21_X1 U19389 ( .B1(n15800), .B2(n18056), .A(n15799), .ZN(n15801) );
  AOI21_X1 U19390 ( .B1(n15802), .B2(n18052), .A(n15801), .ZN(n15803) );
  OAI21_X1 U19391 ( .B1(n21105), .B2(n16026), .A(n15803), .ZN(P1_U2970) );
  NOR2_X1 U19392 ( .A1(n21291), .A2(n15804), .ZN(n16032) );
  NOR2_X1 U19393 ( .A1(n18061), .A2(n15805), .ZN(n15806) );
  AOI211_X1 U19394 ( .C1(n15997), .C2(n15807), .A(n16032), .B(n15806), .ZN(
        n15815) );
  NOR3_X1 U19395 ( .A1(n15808), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15811) );
  NAND2_X1 U19396 ( .A1(n15812), .A2(n16041), .ZN(n15810) );
  MUX2_X1 U19397 ( .A(n16041), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n15979), .Z(n15809) );
  OAI211_X1 U19398 ( .C1(n15812), .C2(n15811), .A(n15810), .B(n15809), .ZN(
        n15813) );
  XNOR2_X1 U19399 ( .A(n15813), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16027) );
  NAND2_X1 U19400 ( .A1(n16027), .A2(n11864), .ZN(n15814) );
  OAI211_X1 U19401 ( .C1(n15816), .C2(n18057), .A(n15815), .B(n15814), .ZN(
        P1_U2971) );
  MUX2_X1 U19402 ( .A(n15818), .B(n15817), .S(n15979), .Z(n15819) );
  XNOR2_X1 U19403 ( .A(n15819), .B(n16041), .ZN(n16046) );
  NAND2_X1 U19404 ( .A1(n18072), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n16040) );
  NAND2_X1 U19405 ( .A1(n18048), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15820) );
  OAI211_X1 U19406 ( .C1(n18056), .C2(n15821), .A(n16040), .B(n15820), .ZN(
        n15822) );
  AOI21_X1 U19407 ( .B1(n15823), .B2(n18052), .A(n15822), .ZN(n15824) );
  OAI21_X1 U19408 ( .B1(n21105), .B2(n16046), .A(n15824), .ZN(P1_U2972) );
  NAND2_X1 U19409 ( .A1(n15857), .A2(n10297), .ZN(n15825) );
  NAND2_X1 U19410 ( .A1(n15825), .A2(n15993), .ZN(n15826) );
  NAND2_X1 U19411 ( .A1(n15827), .A2(n15826), .ZN(n15828) );
  XNOR2_X1 U19412 ( .A(n15828), .B(n16049), .ZN(n16056) );
  NOR2_X1 U19413 ( .A1(n21291), .A2(n15829), .ZN(n16052) );
  AOI21_X1 U19414 ( .B1(n18048), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n16052), .ZN(n15830) );
  OAI21_X1 U19415 ( .B1(n15831), .B2(n18056), .A(n15830), .ZN(n15832) );
  AOI21_X1 U19416 ( .B1(n15833), .B2(n18052), .A(n15832), .ZN(n15834) );
  OAI21_X1 U19417 ( .B1(n21105), .B2(n16056), .A(n15834), .ZN(P1_U2973) );
  MUX2_X1 U19418 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n15835), .S(
        n15909), .Z(n15838) );
  NAND2_X1 U19419 ( .A1(n15836), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15845) );
  NAND2_X1 U19420 ( .A1(n15845), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15837) );
  NAND2_X1 U19421 ( .A1(n15838), .A2(n15837), .ZN(n15839) );
  XNOR2_X1 U19422 ( .A(n15839), .B(n16060), .ZN(n16065) );
  NAND2_X1 U19423 ( .A1(n18072), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n16059) );
  NAND2_X1 U19424 ( .A1(n18048), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15840) );
  OAI211_X1 U19425 ( .C1(n18056), .C2(n15841), .A(n16059), .B(n15840), .ZN(
        n15842) );
  AOI21_X1 U19426 ( .B1(n15843), .B2(n18052), .A(n15842), .ZN(n15844) );
  OAI21_X1 U19427 ( .B1(n21105), .B2(n16065), .A(n15844), .ZN(P1_U2974) );
  MUX2_X1 U19428 ( .A(n15846), .B(n15845), .S(n15979), .Z(n15847) );
  XNOR2_X1 U19429 ( .A(n15847), .B(n16069), .ZN(n16077) );
  NAND2_X1 U19430 ( .A1(n18072), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n16072) );
  OAI21_X1 U19431 ( .B1(n18061), .B2(n15848), .A(n16072), .ZN(n15851) );
  NOR2_X1 U19432 ( .A1(n15849), .A2(n18057), .ZN(n15850) );
  AOI211_X1 U19433 ( .C1(n15997), .C2(n15852), .A(n15851), .B(n15850), .ZN(
        n15853) );
  OAI21_X1 U19434 ( .B1(n21105), .B2(n16077), .A(n15853), .ZN(P1_U2975) );
  INV_X1 U19435 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n21779) );
  NOR2_X1 U19436 ( .A1(n21291), .A2(n21779), .ZN(n16081) );
  NOR2_X1 U19437 ( .A1(n18056), .A2(n15854), .ZN(n15855) );
  AOI211_X1 U19438 ( .C1(n18048), .C2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16081), .B(n15855), .ZN(n15859) );
  XNOR2_X1 U19439 ( .A(n15909), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15856) );
  XNOR2_X1 U19440 ( .A(n15857), .B(n15856), .ZN(n16078) );
  NAND2_X1 U19441 ( .A1(n16078), .A2(n11864), .ZN(n15858) );
  OAI211_X1 U19442 ( .C1(n15860), .C2(n18057), .A(n15859), .B(n15858), .ZN(
        P1_U2976) );
  NAND2_X1 U19443 ( .A1(n15862), .A2(n15861), .ZN(n15863) );
  XOR2_X1 U19444 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n15863), .Z(
        n16104) );
  NAND2_X1 U19445 ( .A1(n15864), .A2(n18052), .ZN(n15869) );
  INV_X1 U19446 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21971) );
  NOR2_X1 U19447 ( .A1(n21291), .A2(n21971), .ZN(n16094) );
  NOR2_X1 U19448 ( .A1(n18061), .A2(n15865), .ZN(n15866) );
  AOI211_X1 U19449 ( .C1(n15997), .C2(n15867), .A(n16094), .B(n15866), .ZN(
        n15868) );
  OAI211_X1 U19450 ( .C1(n16104), .C2(n21105), .A(n15869), .B(n15868), .ZN(
        P1_U2977) );
  NOR2_X1 U19451 ( .A1(n15993), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15878) );
  OAI21_X1 U19452 ( .B1(n15979), .B2(n16141), .A(n15870), .ZN(n15889) );
  OAI22_X1 U19453 ( .A1(n15889), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n15909), .B2(n15870), .ZN(n15871) );
  OAI21_X1 U19454 ( .B1(n16096), .B2(n15878), .A(n15871), .ZN(n15872) );
  XNOR2_X1 U19455 ( .A(n15872), .B(n16107), .ZN(n16112) );
  NAND2_X1 U19456 ( .A1(n18072), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n16106) );
  NAND2_X1 U19457 ( .A1(n18048), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15873) );
  OAI211_X1 U19458 ( .C1(n18056), .C2(n15874), .A(n16106), .B(n15873), .ZN(
        n15875) );
  AOI21_X1 U19459 ( .B1(n15876), .B2(n18052), .A(n15875), .ZN(n15877) );
  OAI21_X1 U19460 ( .B1(n21105), .B2(n16112), .A(n15877), .ZN(P1_U2978) );
  INV_X1 U19461 ( .A(n15878), .ZN(n15887) );
  NAND2_X1 U19462 ( .A1(n15993), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15886) );
  OAI22_X1 U19463 ( .A1(n15889), .A2(n15887), .B1(n15870), .B2(n15886), .ZN(
        n15879) );
  XNOR2_X1 U19464 ( .A(n15879), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16121) );
  INV_X1 U19465 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15880) );
  NAND2_X1 U19466 ( .A1(n18072), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n16115) );
  OAI21_X1 U19467 ( .B1(n18061), .B2(n15880), .A(n16115), .ZN(n15883) );
  NOR2_X1 U19468 ( .A1(n15881), .A2(n18057), .ZN(n15882) );
  AOI211_X1 U19469 ( .C1(n15997), .C2(n15884), .A(n15883), .B(n15882), .ZN(
        n15885) );
  OAI21_X1 U19470 ( .B1(n16121), .B2(n21105), .A(n15885), .ZN(P1_U2979) );
  NAND2_X1 U19471 ( .A1(n15887), .A2(n15886), .ZN(n15888) );
  XNOR2_X1 U19472 ( .A(n15889), .B(n15888), .ZN(n16131) );
  NOR2_X1 U19473 ( .A1(n21291), .A2(n15890), .ZN(n16124) );
  AOI21_X1 U19474 ( .B1(n18048), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n16124), .ZN(n15891) );
  OAI21_X1 U19475 ( .B1(n15892), .B2(n18056), .A(n15891), .ZN(n15893) );
  AOI21_X1 U19476 ( .B1(n15894), .B2(n18052), .A(n15893), .ZN(n15895) );
  OAI21_X1 U19477 ( .B1(n21105), .B2(n16131), .A(n15895), .ZN(P1_U2980) );
  NAND2_X1 U19478 ( .A1(n18072), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n16140) );
  OAI21_X1 U19479 ( .B1(n18061), .B2(n15896), .A(n16140), .ZN(n15900) );
  OAI21_X1 U19480 ( .B1(n15898), .B2(n15897), .A(n15870), .ZN(n16146) );
  NOR2_X1 U19481 ( .A1(n16146), .A2(n21105), .ZN(n15899) );
  AOI211_X1 U19482 ( .C1(n15997), .C2(n15901), .A(n15900), .B(n15899), .ZN(
        n15902) );
  OAI21_X1 U19483 ( .B1(n18057), .B2(n15903), .A(n15902), .ZN(P1_U2981) );
  NAND2_X1 U19484 ( .A1(n15909), .A2(n16162), .ZN(n15908) );
  INV_X1 U19485 ( .A(n15904), .ZN(n15905) );
  OAI21_X1 U19486 ( .B1(n15905), .B2(n15993), .A(n15952), .ZN(n15942) );
  OAI21_X1 U19487 ( .B1(n15942), .B2(n10290), .A(n15906), .ZN(n15907) );
  MUX2_X1 U19488 ( .A(n15909), .B(n15908), .S(n15907), .Z(n15910) );
  XNOR2_X1 U19489 ( .A(n15910), .B(n16147), .ZN(n16156) );
  NOR2_X1 U19490 ( .A1(n21291), .A2(n21770), .ZN(n16152) );
  NOR2_X1 U19491 ( .A1(n18061), .A2(n22100), .ZN(n15911) );
  AOI211_X1 U19492 ( .C1(n15997), .C2(n15912), .A(n16152), .B(n15911), .ZN(
        n15916) );
  INV_X1 U19493 ( .A(n15913), .ZN(n15914) );
  NAND2_X1 U19494 ( .A1(n15914), .A2(n18052), .ZN(n15915) );
  OAI211_X1 U19495 ( .C1(n16156), .C2(n21105), .A(n15916), .B(n15915), .ZN(
        P1_U2982) );
  INV_X1 U19496 ( .A(n15942), .ZN(n15918) );
  NOR2_X1 U19497 ( .A1(n15918), .A2(n15917), .ZN(n15927) );
  OAI21_X1 U19498 ( .B1(n15927), .B2(n10290), .A(n15930), .ZN(n15919) );
  XOR2_X1 U19499 ( .A(n15920), .B(n15919), .Z(n16167) );
  NAND2_X1 U19500 ( .A1(n15997), .A2(n15921), .ZN(n15922) );
  NAND2_X1 U19501 ( .A1(n18072), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n16157) );
  OAI211_X1 U19502 ( .C1(n18061), .C2(n15923), .A(n15922), .B(n16157), .ZN(
        n15924) );
  AOI21_X1 U19503 ( .B1(n15925), .B2(n18052), .A(n15924), .ZN(n15926) );
  OAI21_X1 U19504 ( .B1(n16167), .B2(n21105), .A(n15926), .ZN(P1_U2983) );
  INV_X1 U19505 ( .A(n15927), .ZN(n15929) );
  NAND2_X1 U19506 ( .A1(n15929), .A2(n15928), .ZN(n15933) );
  NAND2_X1 U19507 ( .A1(n15931), .A2(n15930), .ZN(n15932) );
  XNOR2_X1 U19508 ( .A(n15933), .B(n15932), .ZN(n16168) );
  NAND2_X1 U19509 ( .A1(n16168), .A2(n11864), .ZN(n15937) );
  NOR2_X1 U19510 ( .A1(n21291), .A2(n21860), .ZN(n16171) );
  NOR2_X1 U19511 ( .A1(n18056), .A2(n15934), .ZN(n15935) );
  AOI211_X1 U19512 ( .C1(n18048), .C2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16171), .B(n15935), .ZN(n15936) );
  OAI211_X1 U19513 ( .C1(n18057), .C2(n15938), .A(n15937), .B(n15936), .ZN(
        P1_U2984) );
  INV_X1 U19514 ( .A(n15939), .ZN(n15940) );
  AOI21_X1 U19515 ( .B1(n15942), .B2(n15941), .A(n15940), .ZN(n15944) );
  XNOR2_X1 U19516 ( .A(n15993), .B(n16176), .ZN(n15943) );
  XNOR2_X1 U19517 ( .A(n15944), .B(n15943), .ZN(n16183) );
  NAND2_X1 U19518 ( .A1(n18072), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n16179) );
  NAND2_X1 U19519 ( .A1(n18048), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15945) );
  OAI211_X1 U19520 ( .C1(n18056), .C2(n15946), .A(n16179), .B(n15945), .ZN(
        n15947) );
  AOI21_X1 U19521 ( .B1(n15948), .B2(n18052), .A(n15947), .ZN(n15949) );
  OAI21_X1 U19522 ( .B1(n16183), .B2(n21105), .A(n15949), .ZN(P1_U2985) );
  NOR2_X1 U19523 ( .A1(n21291), .A2(n22109), .ZN(n16188) );
  NOR2_X1 U19524 ( .A1(n18056), .A2(n15950), .ZN(n15951) );
  AOI211_X1 U19525 ( .C1(n18048), .C2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n16188), .B(n15951), .ZN(n15961) );
  INV_X1 U19526 ( .A(n15952), .ZN(n15978) );
  INV_X1 U19527 ( .A(n15953), .ZN(n15954) );
  AOI22_X1 U19528 ( .A1(n15978), .A2(n15955), .B1(n9784), .B2(n15954), .ZN(
        n15967) );
  INV_X1 U19529 ( .A(n15957), .ZN(n15956) );
  AOI21_X1 U19530 ( .B1(n15909), .B2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n15956), .ZN(n15966) );
  NAND2_X1 U19531 ( .A1(n15967), .A2(n15966), .ZN(n15965) );
  NAND2_X1 U19532 ( .A1(n15965), .A2(n15957), .ZN(n15958) );
  XOR2_X1 U19533 ( .A(n15959), .B(n15958), .Z(n16184) );
  NAND2_X1 U19534 ( .A1(n16184), .A2(n11864), .ZN(n15960) );
  OAI211_X1 U19535 ( .C1(n15962), .C2(n18057), .A(n15961), .B(n15960), .ZN(
        P1_U2986) );
  AND2_X1 U19536 ( .A1(n18072), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n16210) );
  NOR2_X1 U19537 ( .A1(n18056), .A2(n15963), .ZN(n15964) );
  AOI211_X1 U19538 ( .C1(n18048), .C2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16210), .B(n15964), .ZN(n15969) );
  OAI21_X1 U19539 ( .B1(n15967), .B2(n15966), .A(n15965), .ZN(n16196) );
  NAND2_X1 U19540 ( .A1(n16196), .A2(n11864), .ZN(n15968) );
  OAI211_X1 U19541 ( .C1(n15970), .C2(n18057), .A(n15969), .B(n15968), .ZN(
        P1_U2987) );
  NAND3_X1 U19542 ( .A1(n15978), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n15979), .ZN(n15971) );
  NAND2_X1 U19543 ( .A1(n15971), .A2(n15982), .ZN(n15972) );
  XNOR2_X1 U19544 ( .A(n15972), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16227) );
  NAND2_X1 U19545 ( .A1(n18072), .A2(P1_REIP_REG_11__SCAN_IN), .ZN(n16219) );
  NAND2_X1 U19546 ( .A1(n18048), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15973) );
  OAI211_X1 U19547 ( .C1(n18056), .C2(n15974), .A(n16219), .B(n15973), .ZN(
        n15975) );
  AOI21_X1 U19548 ( .B1(n15976), .B2(n18052), .A(n15975), .ZN(n15977) );
  OAI21_X1 U19549 ( .B1(n16227), .B2(n21105), .A(n15977), .ZN(P1_U2988) );
  XNOR2_X1 U19550 ( .A(n15978), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15980) );
  MUX2_X1 U19551 ( .A(n15981), .B(n15980), .S(n15979), .Z(n15983) );
  NAND2_X1 U19552 ( .A1(n15983), .A2(n15982), .ZN(n16228) );
  NAND2_X1 U19553 ( .A1(n16228), .A2(n11864), .ZN(n15989) );
  INV_X1 U19554 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n15984) );
  NOR2_X1 U19555 ( .A1(n21291), .A2(n15984), .ZN(n16232) );
  NOR2_X1 U19556 ( .A1(n18061), .A2(n15985), .ZN(n15986) );
  AOI211_X1 U19557 ( .C1(n15997), .C2(n15987), .A(n16232), .B(n15986), .ZN(
        n15988) );
  OAI211_X1 U19558 ( .C1(n18057), .C2(n15990), .A(n15989), .B(n15988), .ZN(
        P1_U2989) );
  XNOR2_X1 U19559 ( .A(n15993), .B(n15992), .ZN(n15994) );
  XNOR2_X1 U19560 ( .A(n15991), .B(n15994), .ZN(n16250) );
  NAND2_X1 U19561 ( .A1(n18072), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n16245) );
  OAI21_X1 U19562 ( .B1(n18061), .B2(n21130), .A(n16245), .ZN(n15996) );
  NOR2_X1 U19563 ( .A1(n21133), .A2(n18057), .ZN(n15995) );
  AOI211_X1 U19564 ( .C1(n15997), .C2(n21134), .A(n15996), .B(n15995), .ZN(
        n15998) );
  OAI21_X1 U19565 ( .B1(n21105), .B2(n16250), .A(n15998), .ZN(P1_U2990) );
  INV_X1 U19566 ( .A(n15999), .ZN(n16002) );
  AOI21_X1 U19567 ( .B1(n15999), .B2(n18069), .A(n16000), .ZN(n16001) );
  AOI21_X1 U19568 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16002), .A(
        n16001), .ZN(n16005) );
  XNOR2_X1 U19569 ( .A(n16003), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16004) );
  XNOR2_X1 U19570 ( .A(n16005), .B(n16004), .ZN(n16266) );
  INV_X1 U19571 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n16006) );
  NOR2_X1 U19572 ( .A1(n21291), .A2(n16006), .ZN(n16263) );
  AOI21_X1 U19573 ( .B1(n18048), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16263), .ZN(n16007) );
  OAI21_X1 U19574 ( .B1(n21145), .B2(n18056), .A(n16007), .ZN(n16008) );
  AOI21_X1 U19575 ( .B1(n21148), .B2(n18052), .A(n16008), .ZN(n16009) );
  OAI21_X1 U19576 ( .B1(n16266), .B2(n21105), .A(n16009), .ZN(P1_U2991) );
  INV_X1 U19577 ( .A(n16011), .ZN(n16016) );
  AOI21_X1 U19578 ( .B1(n16014), .B2(n16013), .A(n16012), .ZN(n16015) );
  AOI211_X1 U19579 ( .C1(n16017), .C2(n21282), .A(n16016), .B(n16015), .ZN(
        n16018) );
  OAI21_X1 U19580 ( .B1(n16010), .B2(n21294), .A(n16018), .ZN(P1_U3001) );
  NOR3_X1 U19581 ( .A1(n16030), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n10147), .ZN(n16019) );
  AOI211_X1 U19582 ( .C1(n16021), .C2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n16020), .B(n16019), .ZN(n16025) );
  INV_X1 U19583 ( .A(n16022), .ZN(n16023) );
  NAND2_X1 U19584 ( .A1(n16023), .A2(n21282), .ZN(n16024) );
  OAI211_X1 U19585 ( .C1(n16026), .C2(n21294), .A(n16025), .B(n16024), .ZN(
        P1_U3002) );
  NAND2_X1 U19586 ( .A1(n16027), .A2(n21286), .ZN(n16035) );
  INV_X1 U19587 ( .A(n16042), .ZN(n16033) );
  NOR3_X1 U19588 ( .A1(n16030), .A2(n16029), .A3(n16028), .ZN(n16031) );
  AOI211_X1 U19589 ( .C1(n16033), .C2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n16032), .B(n16031), .ZN(n16034) );
  OAI211_X1 U19590 ( .C1(n21293), .C2(n16036), .A(n16035), .B(n16034), .ZN(
        P1_U3003) );
  INV_X1 U19591 ( .A(n16037), .ZN(n16044) );
  NAND2_X1 U19592 ( .A1(n16038), .A2(n16041), .ZN(n16039) );
  OAI211_X1 U19593 ( .C1(n16042), .C2(n16041), .A(n16040), .B(n16039), .ZN(
        n16043) );
  AOI21_X1 U19594 ( .B1(n16044), .B2(n21282), .A(n16043), .ZN(n16045) );
  OAI21_X1 U19595 ( .B1(n16046), .B2(n21294), .A(n16045), .ZN(P1_U3004) );
  NOR2_X1 U19596 ( .A1(n16047), .A2(n21293), .ZN(n16054) );
  INV_X1 U19597 ( .A(n16079), .ZN(n16070) );
  NAND3_X1 U19598 ( .A1(n16070), .A2(n16048), .A3(n16060), .ZN(n16058) );
  AOI21_X1 U19599 ( .B1(n16061), .B2(n16058), .A(n16049), .ZN(n16053) );
  NOR3_X1 U19600 ( .A1(n16079), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n16050), .ZN(n16051) );
  NOR4_X1 U19601 ( .A1(n16054), .A2(n16053), .A3(n16052), .A4(n16051), .ZN(
        n16055) );
  OAI21_X1 U19602 ( .B1(n16056), .B2(n21294), .A(n16055), .ZN(P1_U3005) );
  INV_X1 U19603 ( .A(n16057), .ZN(n16063) );
  OAI211_X1 U19604 ( .C1(n16061), .C2(n16060), .A(n16059), .B(n16058), .ZN(
        n16062) );
  AOI21_X1 U19605 ( .B1(n16063), .B2(n21282), .A(n16062), .ZN(n16064) );
  OAI21_X1 U19606 ( .B1(n16065), .B2(n21294), .A(n16064), .ZN(P1_U3006) );
  NOR2_X1 U19607 ( .A1(n16066), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16067) );
  OAI21_X1 U19608 ( .B1(n16068), .B2(n16067), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16073) );
  NAND3_X1 U19609 ( .A1(n16070), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n16069), .ZN(n16071) );
  NAND3_X1 U19610 ( .A1(n16073), .A2(n16072), .A3(n16071), .ZN(n16074) );
  AOI21_X1 U19611 ( .B1(n16075), .B2(n21282), .A(n16074), .ZN(n16076) );
  OAI21_X1 U19612 ( .B1(n16077), .B2(n21294), .A(n16076), .ZN(P1_U3007) );
  NAND2_X1 U19613 ( .A1(n16078), .A2(n21286), .ZN(n16084) );
  NOR2_X1 U19614 ( .A1(n16079), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16080) );
  AOI211_X1 U19615 ( .C1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n16082), .A(
        n16081), .B(n16080), .ZN(n16083) );
  OAI211_X1 U19616 ( .C1(n21293), .C2(n16085), .A(n16084), .B(n16083), .ZN(
        P1_U3008) );
  NAND2_X1 U19617 ( .A1(n16198), .A2(n16134), .ZN(n16088) );
  INV_X1 U19618 ( .A(n16185), .ZN(n16133) );
  NAND3_X1 U19619 ( .A1(n16086), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n16133), .ZN(n16087) );
  NAND2_X1 U19620 ( .A1(n16089), .A2(n16133), .ZN(n16090) );
  NAND2_X1 U19621 ( .A1(n16190), .A2(n16090), .ZN(n16092) );
  NOR2_X1 U19622 ( .A1(n16093), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16095) );
  AOI21_X1 U19623 ( .B1(n16123), .B2(n16095), .A(n16094), .ZN(n16100) );
  AND2_X1 U19624 ( .A1(n16096), .A2(n16107), .ZN(n16097) );
  NAND2_X1 U19625 ( .A1(n16123), .A2(n16097), .ZN(n16105) );
  NAND2_X1 U19626 ( .A1(n16108), .A2(n16105), .ZN(n16098) );
  NAND2_X1 U19627 ( .A1(n16098), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16099) );
  OAI211_X1 U19628 ( .C1(n16101), .C2(n21293), .A(n16100), .B(n16099), .ZN(
        n16102) );
  INV_X1 U19629 ( .A(n16102), .ZN(n16103) );
  OAI21_X1 U19630 ( .B1(n16104), .B2(n21294), .A(n16103), .ZN(P1_U3009) );
  OAI211_X1 U19631 ( .C1(n16108), .C2(n16107), .A(n16106), .B(n16105), .ZN(
        n16109) );
  AOI21_X1 U19632 ( .B1(n16110), .B2(n21282), .A(n16109), .ZN(n16111) );
  OAI21_X1 U19633 ( .B1(n16112), .B2(n21294), .A(n16111), .ZN(P1_U3010) );
  AOI21_X1 U19634 ( .B1(n16123), .B2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16117) );
  NAND2_X1 U19635 ( .A1(n16186), .A2(n16190), .ZN(n16113) );
  AOI21_X1 U19636 ( .B1(n16114), .B2(n16113), .A(n16125), .ZN(n16116) );
  OAI21_X1 U19637 ( .B1(n16117), .B2(n16116), .A(n16115), .ZN(n16118) );
  AOI21_X1 U19638 ( .B1(n16119), .B2(n21282), .A(n16118), .ZN(n16120) );
  OAI21_X1 U19639 ( .B1(n16121), .B2(n21294), .A(n16120), .ZN(P1_U3011) );
  INV_X1 U19640 ( .A(n16122), .ZN(n16129) );
  INV_X1 U19641 ( .A(n16123), .ZN(n16127) );
  AOI21_X1 U19642 ( .B1(n16125), .B2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n16124), .ZN(n16126) );
  OAI21_X1 U19643 ( .B1(n16127), .B2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n16126), .ZN(n16128) );
  AOI21_X1 U19644 ( .B1(n16129), .B2(n21282), .A(n16128), .ZN(n16130) );
  OAI21_X1 U19645 ( .B1(n16131), .B2(n21294), .A(n16130), .ZN(P1_U3012) );
  INV_X1 U19646 ( .A(n16132), .ZN(n16144) );
  NAND2_X1 U19647 ( .A1(n16234), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16136) );
  AOI21_X1 U19648 ( .B1(n16134), .B2(n16252), .A(n16133), .ZN(n16135) );
  OAI21_X1 U19649 ( .B1(n16136), .B2(n16135), .A(n16240), .ZN(n16159) );
  OAI21_X1 U19650 ( .B1(n16137), .B2(n16138), .A(n16159), .ZN(n16154) );
  INV_X1 U19651 ( .A(n16154), .ZN(n16142) );
  NAND3_X1 U19652 ( .A1(n16161), .A2(n16138), .A3(n16141), .ZN(n16139) );
  OAI211_X1 U19653 ( .C1(n16142), .C2(n16141), .A(n16140), .B(n16139), .ZN(
        n16143) );
  AOI21_X1 U19654 ( .B1(n16144), .B2(n21282), .A(n16143), .ZN(n16145) );
  OAI21_X1 U19655 ( .B1(n16146), .B2(n21294), .A(n16145), .ZN(P1_U3013) );
  INV_X1 U19656 ( .A(n16161), .ZN(n16149) );
  OAI21_X1 U19657 ( .B1(n16149), .B2(n16148), .A(n16147), .ZN(n16153) );
  NOR2_X1 U19658 ( .A1(n16150), .A2(n21293), .ZN(n16151) );
  AOI211_X1 U19659 ( .C1(n16154), .C2(n16153), .A(n16152), .B(n16151), .ZN(
        n16155) );
  OAI21_X1 U19660 ( .B1(n16156), .B2(n21294), .A(n16155), .ZN(P1_U3014) );
  NAND4_X1 U19661 ( .A1(n16161), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A4(n16162), .ZN(n16158) );
  NAND2_X1 U19662 ( .A1(n16158), .A2(n16157), .ZN(n16164) );
  INV_X1 U19663 ( .A(n16159), .ZN(n16191) );
  AOI21_X1 U19664 ( .B1(n16176), .B2(n16257), .A(n16191), .ZN(n16175) );
  NOR2_X1 U19665 ( .A1(n16176), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16160) );
  NAND2_X1 U19666 ( .A1(n16161), .A2(n16160), .ZN(n16169) );
  AOI21_X1 U19667 ( .B1(n16175), .B2(n16169), .A(n16162), .ZN(n16163) );
  AOI211_X1 U19668 ( .C1(n21282), .C2(n16165), .A(n16164), .B(n16163), .ZN(
        n16166) );
  OAI21_X1 U19669 ( .B1(n16167), .B2(n21294), .A(n16166), .ZN(P1_U3015) );
  NAND2_X1 U19670 ( .A1(n16168), .A2(n21286), .ZN(n16174) );
  INV_X1 U19671 ( .A(n16169), .ZN(n16170) );
  AOI211_X1 U19672 ( .C1(n16172), .C2(n21282), .A(n16171), .B(n16170), .ZN(
        n16173) );
  OAI211_X1 U19673 ( .C1(n16175), .C2(n22124), .A(n16174), .B(n16173), .ZN(
        P1_U3016) );
  AND2_X1 U19674 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n16235) );
  NAND2_X1 U19675 ( .A1(n16207), .A2(n16235), .ZN(n16256) );
  NAND2_X1 U19676 ( .A1(n16256), .A2(n16203), .ZN(n16213) );
  NAND3_X1 U19677 ( .A1(n16213), .A2(n16177), .A3(n16176), .ZN(n16178) );
  OAI211_X1 U19678 ( .C1(n16180), .C2(n21293), .A(n16179), .B(n16178), .ZN(
        n16181) );
  AOI21_X1 U19679 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16191), .A(
        n16181), .ZN(n16182) );
  OAI21_X1 U19680 ( .B1(n16183), .B2(n21294), .A(n16182), .ZN(P1_U3017) );
  INV_X1 U19681 ( .A(n16184), .ZN(n16195) );
  NOR3_X1 U19682 ( .A1(n16186), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        n16185), .ZN(n16187) );
  AOI211_X1 U19683 ( .C1(n16189), .C2(n21282), .A(n16188), .B(n16187), .ZN(
        n16194) );
  INV_X1 U19684 ( .A(n16190), .ZN(n16192) );
  OAI21_X1 U19685 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16192), .A(
        n16191), .ZN(n16193) );
  OAI211_X1 U19686 ( .C1(n16195), .C2(n21294), .A(n16194), .B(n16193), .ZN(
        P1_U3018) );
  INV_X1 U19687 ( .A(n16196), .ZN(n16218) );
  INV_X1 U19688 ( .A(n16197), .ZN(n16211) );
  NAND2_X1 U19689 ( .A1(n16198), .A2(n16236), .ZN(n16199) );
  NAND2_X1 U19690 ( .A1(n16234), .A2(n16199), .ZN(n16253) );
  INV_X1 U19691 ( .A(n16200), .ZN(n16201) );
  NAND2_X1 U19692 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16201), .ZN(
        n16202) );
  NOR2_X1 U19693 ( .A1(n16222), .A2(n16202), .ZN(n16204) );
  OAI22_X1 U19694 ( .A1(n16252), .A2(n16204), .B1(n16215), .B2(n16203), .ZN(
        n16205) );
  OR2_X1 U19695 ( .A1(n16253), .A2(n16205), .ZN(n16225) );
  AOI21_X1 U19696 ( .B1(n16207), .B2(n16206), .A(n16225), .ZN(n16208) );
  NOR2_X1 U19697 ( .A1(n16208), .A2(n16214), .ZN(n16209) );
  AOI211_X1 U19698 ( .C1(n21282), .C2(n16211), .A(n16210), .B(n16209), .ZN(
        n16217) );
  NAND2_X1 U19699 ( .A1(n16213), .A2(n16212), .ZN(n21290) );
  NAND3_X1 U19700 ( .A1(n16221), .A2(n16215), .A3(n16214), .ZN(n16216) );
  OAI211_X1 U19701 ( .C1(n16218), .C2(n21294), .A(n16217), .B(n16216), .ZN(
        P1_U3019) );
  OAI21_X1 U19702 ( .B1(n16220), .B2(n21293), .A(n16219), .ZN(n16224) );
  NAND2_X1 U19703 ( .A1(n16221), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n18064) );
  NOR3_X1 U19704 ( .A1(n18064), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        n16222), .ZN(n16223) );
  AOI211_X1 U19705 ( .C1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n16225), .A(
        n16224), .B(n16223), .ZN(n16226) );
  OAI21_X1 U19706 ( .B1(n16227), .B2(n21294), .A(n16226), .ZN(P1_U3020) );
  INV_X1 U19707 ( .A(n16228), .ZN(n16244) );
  INV_X1 U19708 ( .A(n16229), .ZN(n16230) );
  NOR3_X1 U19709 ( .A1(n18064), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n16230), .ZN(n16231) );
  AOI211_X1 U19710 ( .C1(n21282), .C2(n16233), .A(n16232), .B(n16231), .ZN(
        n16243) );
  NOR3_X1 U19711 ( .A1(n18064), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        n16259), .ZN(n16246) );
  OAI21_X1 U19712 ( .B1(n16252), .B2(n16235), .A(n16234), .ZN(n21279) );
  INV_X1 U19713 ( .A(n16236), .ZN(n16238) );
  NAND3_X1 U19714 ( .A1(n16238), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        n16237), .ZN(n16239) );
  OR2_X1 U19715 ( .A1(n21279), .A2(n16239), .ZN(n16241) );
  AND2_X1 U19716 ( .A1(n16241), .A2(n16240), .ZN(n16248) );
  OAI21_X1 U19717 ( .B1(n16246), .B2(n16248), .A(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16242) );
  OAI211_X1 U19718 ( .C1(n16244), .C2(n21294), .A(n16243), .B(n16242), .ZN(
        P1_U3021) );
  OAI21_X1 U19719 ( .B1(n21127), .B2(n21293), .A(n16245), .ZN(n16247) );
  AOI211_X1 U19720 ( .C1(n16248), .C2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n16247), .B(n16246), .ZN(n16249) );
  OAI21_X1 U19721 ( .B1(n16250), .B2(n21294), .A(n16249), .ZN(P1_U3022) );
  INV_X1 U19722 ( .A(n21142), .ZN(n16264) );
  INV_X1 U19723 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16258) );
  NAND2_X1 U19724 ( .A1(n16251), .A2(n18080), .ZN(n18085) );
  INV_X1 U19725 ( .A(n16252), .ZN(n16254) );
  AOI21_X1 U19726 ( .B1(n16255), .B2(n16254), .A(n16253), .ZN(n18081) );
  OAI21_X1 U19727 ( .B1(n16256), .B2(n18085), .A(n18081), .ZN(n18074) );
  AOI21_X1 U19728 ( .B1(n16258), .B2(n16257), .A(n18074), .ZN(n18070) );
  INV_X1 U19729 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16261) );
  OAI21_X1 U19730 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16259), .ZN(n16260) );
  OAI22_X1 U19731 ( .A1(n18070), .A2(n16261), .B1(n18064), .B2(n16260), .ZN(
        n16262) );
  AOI211_X1 U19732 ( .C1(n21282), .C2(n16264), .A(n16263), .B(n16262), .ZN(
        n16265) );
  OAI21_X1 U19733 ( .B1(n21294), .B2(n16266), .A(n16265), .ZN(P1_U3023) );
  OAI21_X1 U19734 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n9707), .A(n21672), 
        .ZN(n16267) );
  OAI21_X1 U19735 ( .B1(n16268), .B2(n14754), .A(n16267), .ZN(n16269) );
  MUX2_X1 U19736 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n16269), .S(
        n21302), .Z(P1_U3477) );
  NOR2_X1 U19737 ( .A1(n10699), .A2(n13805), .ZN(n16276) );
  INV_X1 U19738 ( .A(n16276), .ZN(n16271) );
  OAI22_X1 U19739 ( .A1(n17995), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n16271), .B2(n16270), .ZN(n16272) );
  AOI21_X1 U19740 ( .B1(n21564), .B2(n16273), .A(n16272), .ZN(n17996) );
  AOI22_X1 U19741 ( .A1(n16277), .A2(n16276), .B1(n16275), .B2(n16274), .ZN(
        n16278) );
  OAI21_X1 U19742 ( .B1(n17996), .B2(n21802), .A(n16278), .ZN(n16279) );
  MUX2_X1 U19743 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n16279), .S(
        n18088), .Z(P1_U3473) );
  AOI21_X1 U19744 ( .B1(n21510), .B2(n16313), .A(n21528), .ZN(n16280) );
  NOR2_X1 U19745 ( .A1(n16280), .A2(n21667), .ZN(n16286) );
  NOR2_X1 U19746 ( .A1(n21479), .A2(n14754), .ZN(n16284) );
  INV_X1 U19747 ( .A(n21451), .ZN(n16281) );
  NOR2_X1 U19748 ( .A1(n16324), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21379) );
  INV_X1 U19749 ( .A(n16282), .ZN(n16283) );
  NOR2_X1 U19750 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n16283), .ZN(
        n16311) );
  INV_X1 U19751 ( .A(n16284), .ZN(n16285) );
  NOR2_X1 U19752 ( .A1(n21379), .A2(n10952), .ZN(n21376) );
  AOI21_X1 U19753 ( .B1(n16286), .B2(n16285), .A(n21376), .ZN(n16287) );
  OAI211_X1 U19754 ( .C1(n16311), .C2(n11673), .A(n21457), .B(n16287), .ZN(
        n16310) );
  AOI22_X1 U19755 ( .A1(n21670), .A2(n16311), .B1(
        P1_INSTQUEUE_REG_6__0__SCAN_IN), .B2(n16310), .ZN(n16288) );
  OAI21_X1 U19756 ( .B1(n16313), .B2(n21683), .A(n16288), .ZN(n16289) );
  AOI21_X1 U19757 ( .B1(n21498), .B2(n21680), .A(n16289), .ZN(n16290) );
  OAI21_X1 U19758 ( .B1(n16316), .B2(n16326), .A(n16290), .ZN(P1_U3081) );
  AOI22_X1 U19759 ( .A1(n21684), .A2(n16311), .B1(
        P1_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n16310), .ZN(n16291) );
  OAI21_X1 U19760 ( .B1(n16313), .B2(n21577), .A(n16291), .ZN(n16292) );
  AOI21_X1 U19761 ( .B1(n21498), .B2(n16351), .A(n16292), .ZN(n16293) );
  OAI21_X1 U19762 ( .B1(n16316), .B2(n16382), .A(n16293), .ZN(P1_U3082) );
  AOI22_X1 U19763 ( .A1(n21690), .A2(n16311), .B1(
        P1_INSTQUEUE_REG_6__2__SCAN_IN), .B2(n16310), .ZN(n16294) );
  OAI21_X1 U19764 ( .B1(n16313), .B2(n21695), .A(n16294), .ZN(n16295) );
  AOI21_X1 U19765 ( .B1(n21498), .B2(n21692), .A(n16295), .ZN(n16296) );
  OAI21_X1 U19766 ( .B1(n16316), .B2(n16356), .A(n16296), .ZN(P1_U3083) );
  AOI22_X1 U19767 ( .A1(n21696), .A2(n16311), .B1(
        P1_INSTQUEUE_REG_6__3__SCAN_IN), .B2(n16310), .ZN(n16297) );
  OAI21_X1 U19768 ( .B1(n16313), .B2(n21701), .A(n16297), .ZN(n16298) );
  AOI21_X1 U19769 ( .B1(n21498), .B2(n21698), .A(n16298), .ZN(n16299) );
  OAI21_X1 U19770 ( .B1(n16316), .B2(n16391), .A(n16299), .ZN(P1_U3084) );
  AOI22_X1 U19771 ( .A1(n21702), .A2(n16311), .B1(
        P1_INSTQUEUE_REG_6__4__SCAN_IN), .B2(n16310), .ZN(n16300) );
  OAI21_X1 U19772 ( .B1(n16313), .B2(n21646), .A(n16300), .ZN(n16301) );
  AOI21_X1 U19773 ( .B1(n21498), .B2(n21621), .A(n16301), .ZN(n16302) );
  OAI21_X1 U19774 ( .B1(n16316), .B2(n16303), .A(n16302), .ZN(P1_U3085) );
  AOI22_X1 U19775 ( .A1(n21708), .A2(n16311), .B1(
        P1_INSTQUEUE_REG_6__5__SCAN_IN), .B2(n16310), .ZN(n16304) );
  OAI21_X1 U19776 ( .B1(n16313), .B2(n21597), .A(n16304), .ZN(n16305) );
  AOI21_X1 U19777 ( .B1(n21498), .B2(n21546), .A(n16305), .ZN(n16306) );
  OAI21_X1 U19778 ( .B1(n16316), .B2(n16363), .A(n16306), .ZN(P1_U3086) );
  AOI22_X1 U19779 ( .A1(n21714), .A2(n16311), .B1(
        P1_INSTQUEUE_REG_6__6__SCAN_IN), .B2(n16310), .ZN(n16307) );
  OAI21_X1 U19780 ( .B1(n16313), .B2(n21631), .A(n16307), .ZN(n16308) );
  AOI21_X1 U19781 ( .B1(n21498), .B2(n21628), .A(n16308), .ZN(n16309) );
  OAI21_X1 U19782 ( .B1(n16316), .B2(n16405), .A(n16309), .ZN(P1_U3087) );
  AOI22_X1 U19783 ( .A1(n21723), .A2(n16311), .B1(
        P1_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n16310), .ZN(n16312) );
  OAI21_X1 U19784 ( .B1(n16313), .B2(n21732), .A(n16312), .ZN(n16314) );
  AOI21_X1 U19785 ( .B1(n21498), .B2(n21726), .A(n16314), .ZN(n16315) );
  OAI21_X1 U19786 ( .B1(n16316), .B2(n16410), .A(n16315), .ZN(P1_U3088) );
  INV_X1 U19787 ( .A(n21454), .ZN(n16318) );
  AOI21_X1 U19788 ( .B1(n21559), .B2(n16323), .A(n21528), .ZN(n16319) );
  AOI21_X1 U19789 ( .B1(n21565), .B2(n14754), .A(n16319), .ZN(n16320) );
  NOR2_X1 U19790 ( .A1(n16320), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n16322) );
  INV_X1 U19791 ( .A(n21560), .ZN(n21525) );
  NOR2_X1 U19792 ( .A1(n21525), .A2(n21453), .ZN(n21518) );
  NAND2_X1 U19793 ( .A1(n16321), .A2(n21451), .ZN(n21375) );
  NAND2_X1 U19794 ( .A1(n21521), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n16329) );
  NOR2_X1 U19795 ( .A1(n21564), .A2(n21667), .ZN(n21449) );
  AND2_X1 U19796 ( .A1(n21312), .A2(n16324), .ZN(n16344) );
  AOI22_X1 U19797 ( .A1(n21565), .A2(n21449), .B1(n16344), .B2(n16325), .ZN(
        n21511) );
  INV_X1 U19798 ( .A(n21518), .ZN(n16336) );
  OAI22_X1 U19799 ( .A1(n21511), .A2(n16326), .B1(n16336), .B2(n21639), .ZN(
        n16327) );
  AOI21_X1 U19800 ( .B1(n21520), .B2(n21680), .A(n16327), .ZN(n16328) );
  OAI211_X1 U19801 ( .C1(n21683), .C2(n21559), .A(n16329), .B(n16328), .ZN(
        P1_U3097) );
  NAND2_X1 U19802 ( .A1(n21521), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n16332) );
  OAI22_X1 U19803 ( .A1(n21511), .A2(n16382), .B1(n16336), .B2(n21576), .ZN(
        n16330) );
  AOI21_X1 U19804 ( .B1(n21520), .B2(n16351), .A(n16330), .ZN(n16331) );
  OAI211_X1 U19805 ( .C1(n21577), .C2(n21559), .A(n16332), .B(n16331), .ZN(
        P1_U3098) );
  NAND2_X1 U19806 ( .A1(n21521), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n16335) );
  OAI22_X1 U19807 ( .A1(n21511), .A2(n16356), .B1(n16336), .B2(n21581), .ZN(
        n16333) );
  AOI21_X1 U19808 ( .B1(n21520), .B2(n21692), .A(n16333), .ZN(n16334) );
  OAI211_X1 U19809 ( .C1(n21695), .C2(n21559), .A(n16335), .B(n16334), .ZN(
        P1_U3099) );
  NAND2_X1 U19810 ( .A1(n21521), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n16339) );
  OAI22_X1 U19811 ( .A1(n21511), .A2(n16363), .B1(n16336), .B2(n21593), .ZN(
        n16337) );
  AOI21_X1 U19812 ( .B1(n21520), .B2(n21546), .A(n16337), .ZN(n16338) );
  OAI211_X1 U19813 ( .C1(n21597), .C2(n21559), .A(n16339), .B(n16338), .ZN(
        P1_U3102) );
  NAND2_X1 U19814 ( .A1(n21653), .A2(n21647), .ZN(n16340) );
  NAND2_X1 U19815 ( .A1(n16340), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n16341) );
  NAND2_X1 U19816 ( .A1(n16341), .A2(n21679), .ZN(n16346) );
  OR2_X1 U19817 ( .A1(n21660), .A2(n21564), .ZN(n16343) );
  INV_X1 U19818 ( .A(n16344), .ZN(n16342) );
  OAI22_X1 U19819 ( .A1(n16346), .A2(n16343), .B1(n16342), .B2(n21451), .ZN(
        n21649) );
  NOR2_X1 U19820 ( .A1(n21664), .A2(n21453), .ZN(n21638) );
  INV_X1 U19821 ( .A(n16343), .ZN(n16345) );
  OAI22_X1 U19822 ( .A1(n16346), .A2(n16345), .B1(n16344), .B2(n10952), .ZN(
        n16347) );
  INV_X1 U19823 ( .A(n16347), .ZN(n16348) );
  OAI211_X1 U19824 ( .C1(n21638), .C2(n11673), .A(n21457), .B(n16348), .ZN(
        n21650) );
  AOI22_X1 U19825 ( .A1(n21684), .A2(n21638), .B1(
        P1_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n21650), .ZN(n16349) );
  OAI21_X1 U19826 ( .B1(n21647), .B2(n21577), .A(n16349), .ZN(n16350) );
  AOI21_X1 U19827 ( .B1(n21624), .B2(n16351), .A(n16350), .ZN(n16352) );
  OAI21_X1 U19828 ( .B1(n16370), .B2(n16382), .A(n16352), .ZN(P1_U3130) );
  AOI22_X1 U19829 ( .A1(n21690), .A2(n21638), .B1(
        P1_INSTQUEUE_REG_12__2__SCAN_IN), .B2(n21650), .ZN(n16353) );
  OAI21_X1 U19830 ( .B1(n21647), .B2(n21695), .A(n16353), .ZN(n16354) );
  AOI21_X1 U19831 ( .B1(n21624), .B2(n21692), .A(n16354), .ZN(n16355) );
  OAI21_X1 U19832 ( .B1(n16370), .B2(n16356), .A(n16355), .ZN(P1_U3131) );
  AOI22_X1 U19833 ( .A1(n21696), .A2(n21638), .B1(
        P1_INSTQUEUE_REG_12__3__SCAN_IN), .B2(n21650), .ZN(n16357) );
  OAI21_X1 U19834 ( .B1(n21647), .B2(n21701), .A(n16357), .ZN(n16358) );
  AOI21_X1 U19835 ( .B1(n21624), .B2(n21698), .A(n16358), .ZN(n16359) );
  OAI21_X1 U19836 ( .B1(n16370), .B2(n16391), .A(n16359), .ZN(P1_U3132) );
  AOI22_X1 U19837 ( .A1(n21708), .A2(n21638), .B1(
        P1_INSTQUEUE_REG_12__5__SCAN_IN), .B2(n21650), .ZN(n16360) );
  OAI21_X1 U19838 ( .B1(n21647), .B2(n21597), .A(n16360), .ZN(n16361) );
  AOI21_X1 U19839 ( .B1(n21624), .B2(n21546), .A(n16361), .ZN(n16362) );
  OAI21_X1 U19840 ( .B1(n16370), .B2(n16363), .A(n16362), .ZN(P1_U3134) );
  AOI22_X1 U19841 ( .A1(n21714), .A2(n21638), .B1(
        P1_INSTQUEUE_REG_12__6__SCAN_IN), .B2(n21650), .ZN(n16364) );
  OAI21_X1 U19842 ( .B1(n21647), .B2(n21631), .A(n16364), .ZN(n16365) );
  AOI21_X1 U19843 ( .B1(n21624), .B2(n21628), .A(n16365), .ZN(n16366) );
  OAI21_X1 U19844 ( .B1(n16370), .B2(n16405), .A(n16366), .ZN(P1_U3135) );
  AOI22_X1 U19845 ( .A1(n21723), .A2(n21638), .B1(
        P1_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n21650), .ZN(n16367) );
  OAI21_X1 U19846 ( .B1(n21647), .B2(n21732), .A(n16367), .ZN(n16368) );
  AOI21_X1 U19847 ( .B1(n21624), .B2(n21726), .A(n16368), .ZN(n16369) );
  OAI21_X1 U19848 ( .B1(n16370), .B2(n16410), .A(n16369), .ZN(P1_U3136) );
  INV_X1 U19849 ( .A(n21673), .ZN(n16372) );
  NAND2_X1 U19850 ( .A1(n21662), .A2(n21665), .ZN(n16377) );
  AOI21_X1 U19851 ( .B1(n16377), .B2(n21667), .A(n21484), .ZN(n16371) );
  OAI21_X1 U19852 ( .B1(n16372), .B2(n21667), .A(n16371), .ZN(n16375) );
  NOR2_X1 U19853 ( .A1(n21660), .A2(n16373), .ZN(n16374) );
  NOR3_X2 U19854 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21561), .A3(
        n21664), .ZN(n16411) );
  OAI21_X1 U19855 ( .B1(n16374), .B2(n16411), .A(n21679), .ZN(n16376) );
  INV_X1 U19856 ( .A(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n16381) );
  OAI21_X1 U19857 ( .B1(n16377), .B2(n10952), .A(n16376), .ZN(n16412) );
  AOI22_X1 U19858 ( .A1(n16412), .A2(n21671), .B1(n21670), .B2(n16411), .ZN(
        n16378) );
  OAI21_X1 U19859 ( .B1(n21647), .B2(n21643), .A(n16378), .ZN(n16379) );
  AOI21_X1 U19860 ( .B1(n10689), .B2(n21535), .A(n16379), .ZN(n16380) );
  OAI21_X1 U19861 ( .B1(n16417), .B2(n16381), .A(n16380), .ZN(P1_U3137) );
  INV_X1 U19862 ( .A(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n16386) );
  INV_X1 U19863 ( .A(n21577), .ZN(n21686) );
  AOI22_X1 U19864 ( .A1(n16412), .A2(n21685), .B1(n21684), .B2(n16411), .ZN(
        n16383) );
  OAI21_X1 U19865 ( .B1(n21647), .B2(n21689), .A(n16383), .ZN(n16384) );
  AOI21_X1 U19866 ( .B1(n10689), .B2(n21686), .A(n16384), .ZN(n16385) );
  OAI21_X1 U19867 ( .B1(n16417), .B2(n16386), .A(n16385), .ZN(P1_U3138) );
  INV_X1 U19868 ( .A(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n16390) );
  INV_X1 U19869 ( .A(n21695), .ZN(n21615) );
  AOI22_X1 U19870 ( .A1(n16412), .A2(n21691), .B1(n21690), .B2(n16411), .ZN(
        n16387) );
  OAI21_X1 U19871 ( .B1(n21647), .B2(n21618), .A(n16387), .ZN(n16388) );
  AOI21_X1 U19872 ( .B1(n10689), .B2(n21615), .A(n16388), .ZN(n16389) );
  OAI21_X1 U19873 ( .B1(n16417), .B2(n16390), .A(n16389), .ZN(P1_U3139) );
  INV_X1 U19874 ( .A(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16396) );
  INV_X1 U19875 ( .A(n21701), .ZN(n16394) );
  AOI22_X1 U19876 ( .A1(n16412), .A2(n21697), .B1(n21696), .B2(n16411), .ZN(
        n16392) );
  OAI21_X1 U19877 ( .B1(n21647), .B2(n21586), .A(n16392), .ZN(n16393) );
  AOI21_X1 U19878 ( .B1(n10689), .B2(n16394), .A(n16393), .ZN(n16395) );
  OAI21_X1 U19879 ( .B1(n16417), .B2(n16396), .A(n16395), .ZN(P1_U3140) );
  INV_X1 U19880 ( .A(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n16400) );
  INV_X1 U19881 ( .A(n21646), .ZN(n21704) );
  AOI22_X1 U19882 ( .A1(n16412), .A2(n21703), .B1(n21702), .B2(n16411), .ZN(
        n16397) );
  OAI21_X1 U19883 ( .B1(n21647), .B2(n21707), .A(n16397), .ZN(n16398) );
  AOI21_X1 U19884 ( .B1(n10689), .B2(n21704), .A(n16398), .ZN(n16399) );
  OAI21_X1 U19885 ( .B1(n16417), .B2(n16400), .A(n16399), .ZN(P1_U3141) );
  INV_X1 U19886 ( .A(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16404) );
  INV_X1 U19887 ( .A(n21597), .ZN(n21710) );
  AOI22_X1 U19888 ( .A1(n16412), .A2(n21709), .B1(n21708), .B2(n16411), .ZN(
        n16401) );
  OAI21_X1 U19889 ( .B1(n21647), .B2(n21713), .A(n16401), .ZN(n16402) );
  AOI21_X1 U19890 ( .B1(n10689), .B2(n21710), .A(n16402), .ZN(n16403) );
  OAI21_X1 U19891 ( .B1(n16417), .B2(n16404), .A(n16403), .ZN(P1_U3142) );
  INV_X1 U19892 ( .A(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16409) );
  INV_X1 U19893 ( .A(n21631), .ZN(n21716) );
  AOI22_X1 U19894 ( .A1(n16412), .A2(n21715), .B1(n21714), .B2(n16411), .ZN(
        n16406) );
  OAI21_X1 U19895 ( .B1(n21647), .B2(n21721), .A(n16406), .ZN(n16407) );
  AOI21_X1 U19896 ( .B1(n10689), .B2(n21716), .A(n16407), .ZN(n16408) );
  OAI21_X1 U19897 ( .B1(n16417), .B2(n16409), .A(n16408), .ZN(P1_U3143) );
  INV_X1 U19898 ( .A(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16416) );
  INV_X1 U19899 ( .A(n21732), .ZN(n21554) );
  AOI22_X1 U19900 ( .A1(n16412), .A2(n21724), .B1(n21723), .B2(n16411), .ZN(
        n16413) );
  OAI21_X1 U19901 ( .B1(n21647), .B2(n21610), .A(n16413), .ZN(n16414) );
  AOI21_X1 U19902 ( .B1(n10689), .B2(n21554), .A(n16414), .ZN(n16415) );
  OAI21_X1 U19903 ( .B1(n16417), .B2(n16416), .A(n16415), .ZN(P1_U3144) );
  AOI211_X1 U19904 ( .C1(n16419), .C2(n20712), .A(n20900), .B(n16418), .ZN(
        n16420) );
  NOR2_X1 U19905 ( .A1(n16420), .A2(n18138), .ZN(n16425) );
  AOI21_X1 U19906 ( .B1(n16421), .B2(n20834), .A(n21042), .ZN(n16422) );
  OAI211_X1 U19907 ( .C1(n20959), .C2(n20419), .A(n16423), .B(n16422), .ZN(
        n16424) );
  MUX2_X1 U19908 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .B(n16425), .S(n16424), 
        .Z(P2_U3610) );
  OAI22_X1 U19909 ( .A1(n22023), .A2(n20335), .B1(n20292), .B2(n21028), .ZN(
        n16427) );
  AOI21_X1 U19910 ( .B1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20262), .A(
        n16427), .ZN(n16428) );
  NOR2_X1 U19911 ( .A1(n16853), .A2(n20341), .ZN(n16429) );
  AOI21_X1 U19912 ( .B1(n16434), .B2(n20326), .A(n16692), .ZN(n16437) );
  NAND2_X1 U19913 ( .A1(n16431), .A2(n16736), .ZN(n16436) );
  OAI22_X1 U19914 ( .A1(n16432), .A2(n20335), .B1(n20292), .B2(n21026), .ZN(
        n16435) );
  INV_X1 U19915 ( .A(n16980), .ZN(n16433) );
  INV_X1 U19916 ( .A(n16438), .ZN(n16440) );
  OAI21_X1 U19917 ( .B1(n16440), .B2(n9897), .A(n16439), .ZN(n17253) );
  AOI21_X1 U19918 ( .B1(n16442), .B2(n16441), .A(n13205), .ZN(n17260) );
  NAND2_X1 U19919 ( .A1(n17260), .A2(n20329), .ZN(n16450) );
  XOR2_X1 U19920 ( .A(n16990), .B(n16443), .Z(n16448) );
  AOI22_X1 U19921 ( .A1(P2_EBX_REG_27__SCAN_IN), .A2(n20295), .B1(n20344), 
        .B2(P2_REIP_REG_27__SCAN_IN), .ZN(n16444) );
  OAI21_X1 U19922 ( .B1(n22083), .B2(n20339), .A(n16444), .ZN(n16447) );
  NOR2_X1 U19923 ( .A1(n16445), .A2(n20336), .ZN(n16446) );
  AOI211_X1 U19924 ( .C1(n20326), .C2(n16448), .A(n16447), .B(n16446), .ZN(
        n16449) );
  OAI211_X1 U19925 ( .C1(n20341), .C2(n17253), .A(n16450), .B(n16449), .ZN(
        P2_U2828) );
  OAI21_X1 U19926 ( .B1(n16451), .B2(n16452), .A(n16438), .ZN(n17272) );
  INV_X1 U19927 ( .A(n16453), .ZN(n16469) );
  INV_X1 U19928 ( .A(n16441), .ZN(n16454) );
  AOI21_X1 U19929 ( .B1(n16455), .B2(n16469), .A(n16454), .ZN(n17264) );
  NAND2_X1 U19930 ( .A1(n17264), .A2(n20329), .ZN(n16465) );
  INV_X1 U19931 ( .A(n12785), .ZN(n16463) );
  AOI21_X1 U19932 ( .B1(n16457), .B2(n20326), .A(n16692), .ZN(n16461) );
  OAI22_X1 U19933 ( .A1(n16767), .A2(n20335), .B1(n20292), .B2(n21023), .ZN(
        n16459) );
  INV_X1 U19934 ( .A(n17004), .ZN(n16456) );
  NOR3_X1 U19935 ( .A1(n16457), .A2(n16456), .A3(n16740), .ZN(n16458) );
  AOI211_X1 U19936 ( .C1(n20262), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n16459), .B(n16458), .ZN(n16460) );
  OAI21_X1 U19937 ( .B1(n16461), .B2(n17004), .A(n16460), .ZN(n16462) );
  AOI21_X1 U19938 ( .B1(n16463), .B2(n16736), .A(n16462), .ZN(n16464) );
  OAI211_X1 U19939 ( .C1(n20341), .C2(n17272), .A(n16465), .B(n16464), .ZN(
        P2_U2829) );
  NAND2_X1 U19940 ( .A1(n16466), .A2(n16467), .ZN(n16468) );
  NAND2_X1 U19941 ( .A1(n16469), .A2(n16468), .ZN(n17284) );
  XNOR2_X1 U19942 ( .A(n16470), .B(n17014), .ZN(n16473) );
  OAI22_X1 U19943 ( .A1(n10511), .A2(n20335), .B1(n20292), .B2(n21021), .ZN(
        n16471) );
  AOI21_X1 U19944 ( .B1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n20262), .A(
        n16471), .ZN(n16472) );
  OAI21_X1 U19945 ( .B1(n16473), .B2(n20351), .A(n16472), .ZN(n16479) );
  INV_X1 U19946 ( .A(n16451), .ZN(n16475) );
  OAI21_X1 U19947 ( .B1(n16477), .B2(n16476), .A(n16475), .ZN(n17279) );
  NOR2_X1 U19948 ( .A1(n17279), .A2(n20341), .ZN(n16478) );
  AOI211_X1 U19949 ( .C1(n16736), .C2(n16480), .A(n16479), .B(n16478), .ZN(
        n16481) );
  OAI21_X1 U19950 ( .B1(n17284), .B2(n20345), .A(n16481), .ZN(P2_U2830) );
  OAI21_X1 U19951 ( .B1(n16498), .B2(n16482), .A(n16466), .ZN(n17294) );
  XNOR2_X1 U19952 ( .A(n16496), .B(n16484), .ZN(n17293) );
  INV_X1 U19953 ( .A(n17293), .ZN(n16890) );
  NOR2_X1 U19954 ( .A1(n16485), .A2(n20336), .ZN(n16493) );
  AOI21_X1 U19955 ( .B1(n16487), .B2(n20326), .A(n16692), .ZN(n16491) );
  INV_X1 U19956 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n21019) );
  OAI22_X1 U19957 ( .A1(n12638), .A2(n20335), .B1(n20292), .B2(n21019), .ZN(
        n16489) );
  INV_X1 U19958 ( .A(n17022), .ZN(n16486) );
  NOR3_X1 U19959 ( .A1(n16487), .A2(n16486), .A3(n16740), .ZN(n16488) );
  AOI211_X1 U19960 ( .C1(n20262), .C2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n16489), .B(n16488), .ZN(n16490) );
  OAI21_X1 U19961 ( .B1(n16491), .B2(n17022), .A(n16490), .ZN(n16492) );
  AOI211_X1 U19962 ( .C1(n16890), .C2(n20330), .A(n16493), .B(n16492), .ZN(
        n16494) );
  OAI21_X1 U19963 ( .B1(n17294), .B2(n20345), .A(n16494), .ZN(P2_U2831) );
  INV_X1 U19964 ( .A(n16495), .ZN(n16497) );
  OAI21_X1 U19965 ( .B1(n16497), .B2(n9898), .A(n16496), .ZN(n17307) );
  AOI21_X1 U19966 ( .B1(n16499), .B2(n16511), .A(n16498), .ZN(n17310) );
  NAND2_X1 U19967 ( .A1(n17310), .A2(n20329), .ZN(n16508) );
  INV_X1 U19968 ( .A(n16500), .ZN(n16506) );
  XNOR2_X1 U19969 ( .A(n16501), .B(n17028), .ZN(n16504) );
  OAI22_X1 U19970 ( .A1(n12868), .A2(n20335), .B1(n20292), .B2(n21017), .ZN(
        n16502) );
  AOI21_X1 U19971 ( .B1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n20262), .A(
        n16502), .ZN(n16503) );
  OAI21_X1 U19972 ( .B1(n16504), .B2(n20351), .A(n16503), .ZN(n16505) );
  AOI21_X1 U19973 ( .B1(n16506), .B2(n16736), .A(n16505), .ZN(n16507) );
  OAI211_X1 U19974 ( .C1(n20341), .C2(n17307), .A(n16508), .B(n16507), .ZN(
        P2_U2832) );
  NAND2_X1 U19975 ( .A1(n13372), .A2(n16509), .ZN(n16510) );
  AND2_X1 U19976 ( .A1(n16511), .A2(n16510), .ZN(n17320) );
  OR2_X1 U19977 ( .A1(n13365), .A2(n16512), .ZN(n16513) );
  NAND2_X1 U19978 ( .A1(n16495), .A2(n16513), .ZN(n17318) );
  INV_X1 U19979 ( .A(n17318), .ZN(n16906) );
  NOR2_X1 U19980 ( .A1(n16514), .A2(n20336), .ZN(n16523) );
  AOI21_X1 U19981 ( .B1(n16517), .B2(n20326), .A(n16692), .ZN(n16521) );
  OAI22_X1 U19982 ( .A1(n16515), .A2(n20335), .B1(n20292), .B2(n21015), .ZN(
        n16519) );
  INV_X1 U19983 ( .A(n17043), .ZN(n16516) );
  NOR3_X1 U19984 ( .A1(n16517), .A2(n16516), .A3(n16740), .ZN(n16518) );
  AOI211_X1 U19985 ( .C1(n20262), .C2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n16519), .B(n16518), .ZN(n16520) );
  OAI21_X1 U19986 ( .B1(n16521), .B2(n17043), .A(n16520), .ZN(n16522) );
  AOI211_X1 U19987 ( .C1(n16906), .C2(n20330), .A(n16523), .B(n16522), .ZN(
        n16524) );
  OAI21_X1 U19988 ( .B1(n16791), .B2(n20345), .A(n16524), .ZN(P2_U2833) );
  XOR2_X1 U19989 ( .A(n17053), .B(n16544), .Z(n16527) );
  AOI22_X1 U19990 ( .A1(P2_EBX_REG_21__SCAN_IN), .A2(n20295), .B1(n20344), 
        .B2(P2_REIP_REG_21__SCAN_IN), .ZN(n16525) );
  OAI21_X1 U19991 ( .B1(n17049), .B2(n20339), .A(n16525), .ZN(n16526) );
  AOI21_X1 U19992 ( .B1(n16527), .B2(n20326), .A(n16526), .ZN(n16528) );
  OAI21_X1 U19993 ( .B1(n16529), .B2(n20336), .A(n16528), .ZN(n16530) );
  AOI21_X1 U19994 ( .B1(n16909), .B2(n20330), .A(n16530), .ZN(n16531) );
  OAI21_X1 U19995 ( .B1(n17050), .B2(n20345), .A(n16531), .ZN(P2_U2834) );
  NAND2_X1 U19996 ( .A1(n16929), .A2(n16533), .ZN(n16534) );
  NAND2_X1 U19997 ( .A1(n13364), .A2(n16534), .ZN(n17332) );
  INV_X1 U19998 ( .A(n13371), .ZN(n16536) );
  OAI21_X1 U19999 ( .B1(n16535), .B2(n16537), .A(n16536), .ZN(n17335) );
  INV_X1 U20000 ( .A(n17335), .ZN(n16538) );
  NAND2_X1 U20001 ( .A1(n16538), .A2(n20329), .ZN(n16550) );
  NOR2_X1 U20002 ( .A1(n20339), .A2(n16539), .ZN(n16543) );
  INV_X1 U20003 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n16541) );
  INV_X1 U20004 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n16540) );
  OAI22_X1 U20005 ( .A1(n16541), .A2(n20335), .B1(n20292), .B2(n16540), .ZN(
        n16542) );
  NOR2_X1 U20006 ( .A1(n16543), .A2(n16542), .ZN(n16546) );
  OAI211_X1 U20007 ( .C1(n20269), .C2(n17062), .A(n16544), .B(n20326), .ZN(
        n16545) );
  OAI211_X1 U20008 ( .C1(n16742), .C2(n17062), .A(n16546), .B(n16545), .ZN(
        n16547) );
  AOI21_X1 U20009 ( .B1(n16548), .B2(n16736), .A(n16547), .ZN(n16549) );
  OAI211_X1 U20010 ( .C1(n20341), .C2(n17332), .A(n16550), .B(n16549), .ZN(
        P2_U2835) );
  INV_X1 U20011 ( .A(n16552), .ZN(n16553) );
  AOI21_X1 U20012 ( .B1(n16554), .B2(n16551), .A(n16553), .ZN(n17080) );
  INV_X1 U20013 ( .A(n17080), .ZN(n17357) );
  OAI21_X1 U20014 ( .B1(n16559), .B2(n20351), .A(n16742), .ZN(n16555) );
  NAND2_X1 U20015 ( .A1(n16555), .A2(n10150), .ZN(n16562) );
  INV_X1 U20016 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n17081) );
  OR2_X1 U20017 ( .A1(n20292), .A2(n17081), .ZN(n16556) );
  OAI211_X1 U20018 ( .C1(n20335), .C2(n16557), .A(n16556), .B(n20260), .ZN(
        n16558) );
  AOI21_X1 U20019 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n20262), .A(
        n16558), .ZN(n16561) );
  NAND3_X1 U20020 ( .A1(n16706), .A2(n16559), .A3(n17084), .ZN(n16560) );
  NAND3_X1 U20021 ( .A1(n16562), .A2(n16561), .A3(n16560), .ZN(n16563) );
  AOI21_X1 U20022 ( .B1(n16564), .B2(n16736), .A(n16563), .ZN(n16569) );
  OR2_X1 U20023 ( .A1(n16573), .A2(n16566), .ZN(n16567) );
  AND2_X1 U20024 ( .A1(n16565), .A2(n16567), .ZN(n17353) );
  NAND2_X1 U20025 ( .A1(n17353), .A2(n20330), .ZN(n16568) );
  OAI211_X1 U20026 ( .C1(n17357), .C2(n20345), .A(n16569), .B(n16568), .ZN(
        P2_U2837) );
  OAI21_X1 U20027 ( .B1(n16586), .B2(n16570), .A(n16551), .ZN(n17370) );
  AND2_X1 U20028 ( .A1(n16589), .A2(n16571), .ZN(n16572) );
  NOR2_X1 U20029 ( .A1(n16573), .A2(n16572), .ZN(n17368) );
  NOR2_X1 U20030 ( .A1(n16574), .A2(n20336), .ZN(n16583) );
  AOI21_X1 U20031 ( .B1(n16577), .B2(n20326), .A(n16692), .ZN(n16581) );
  INV_X1 U20032 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n21007) );
  OAI21_X1 U20033 ( .B1(n21007), .B2(n20292), .A(n20260), .ZN(n16576) );
  NOR2_X1 U20034 ( .A1(n20339), .A2(n13232), .ZN(n16575) );
  AOI211_X1 U20035 ( .C1(n20295), .C2(P2_EBX_REG_17__SCAN_IN), .A(n16576), .B(
        n16575), .ZN(n16580) );
  INV_X1 U20036 ( .A(n16577), .ZN(n16578) );
  NAND3_X1 U20037 ( .A1(n16578), .A2(n16706), .A3(n17090), .ZN(n16579) );
  OAI211_X1 U20038 ( .C1(n16581), .C2(n17090), .A(n16580), .B(n16579), .ZN(
        n16582) );
  AOI211_X1 U20039 ( .C1(n17368), .C2(n20330), .A(n16583), .B(n16582), .ZN(
        n16584) );
  OAI21_X1 U20040 ( .B1(n17370), .B2(n20345), .A(n16584), .ZN(P2_U2838) );
  AND2_X1 U20041 ( .A1(n16824), .A2(n16585), .ZN(n16587) );
  OR2_X1 U20042 ( .A1(n16587), .A2(n16586), .ZN(n17374) );
  INV_X1 U20043 ( .A(n16589), .ZN(n16590) );
  AOI21_X1 U20044 ( .B1(n16591), .B2(n16588), .A(n16590), .ZN(n20364) );
  NOR2_X1 U20045 ( .A1(n16592), .A2(n20336), .ZN(n16600) );
  INV_X1 U20046 ( .A(n20283), .ZN(n16593) );
  AOI21_X1 U20047 ( .B1(n16593), .B2(n20326), .A(n16692), .ZN(n16598) );
  OAI21_X1 U20048 ( .B1(n12847), .B2(n20335), .A(n13139), .ZN(n16595) );
  NOR2_X1 U20049 ( .A1(n20292), .A2(n21005), .ZN(n16594) );
  AOI211_X1 U20050 ( .C1(n20262), .C2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n16595), .B(n16594), .ZN(n16597) );
  NAND3_X1 U20051 ( .A1(n20283), .A2(n16706), .A3(n17100), .ZN(n16596) );
  OAI211_X1 U20052 ( .C1(n16598), .C2(n17100), .A(n16597), .B(n16596), .ZN(
        n16599) );
  AOI211_X1 U20053 ( .C1(n20364), .C2(n20330), .A(n16600), .B(n16599), .ZN(
        n16601) );
  OAI21_X1 U20054 ( .B1(n17374), .B2(n20345), .A(n16601), .ZN(P2_U2839) );
  INV_X1 U20055 ( .A(n16602), .ZN(n17392) );
  NOR2_X1 U20056 ( .A1(n20299), .A2(n10160), .ZN(n16603) );
  XOR2_X1 U20057 ( .A(n17126), .B(n16603), .Z(n16610) );
  NAND2_X1 U20058 ( .A1(n16604), .A2(n16736), .ZN(n16609) );
  AOI21_X1 U20059 ( .B1(n20344), .B2(P2_REIP_REG_14__SCAN_IN), .A(n20343), 
        .ZN(n16605) );
  OAI21_X1 U20060 ( .B1(n16606), .B2(n20335), .A(n16605), .ZN(n16607) );
  AOI21_X1 U20061 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n20262), .A(
        n16607), .ZN(n16608) );
  OAI211_X1 U20062 ( .C1(n20351), .C2(n16610), .A(n16609), .B(n16608), .ZN(
        n16611) );
  AOI21_X1 U20063 ( .B1(n17392), .B2(n20330), .A(n16611), .ZN(n16612) );
  OAI21_X1 U20064 ( .B1(n17395), .B2(n20345), .A(n16612), .ZN(P2_U2841) );
  AND2_X1 U20065 ( .A1(n16613), .A2(n16614), .ZN(n16615) );
  OR2_X1 U20066 ( .A1(n16615), .A2(n14833), .ZN(n17148) );
  INV_X1 U20067 ( .A(n17413), .ZN(n16625) );
  AOI21_X1 U20068 ( .B1(n20326), .B2(n16619), .A(n16692), .ZN(n16623) );
  AOI22_X1 U20069 ( .A1(n16616), .A2(n16736), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n20262), .ZN(n16617) );
  OAI21_X1 U20070 ( .B1(n12832), .B2(n20335), .A(n16617), .ZN(n16618) );
  AOI211_X1 U20071 ( .C1(n20344), .C2(P2_REIP_REG_12__SCAN_IN), .A(n20343), 
        .B(n16618), .ZN(n16622) );
  INV_X1 U20072 ( .A(n16619), .ZN(n16620) );
  NAND3_X1 U20073 ( .A1(n16706), .A2(n17150), .A3(n16620), .ZN(n16621) );
  OAI211_X1 U20074 ( .C1(n16623), .C2(n17150), .A(n16622), .B(n16621), .ZN(
        n16624) );
  AOI21_X1 U20075 ( .B1(n16625), .B2(n20330), .A(n16624), .ZN(n16626) );
  OAI21_X1 U20076 ( .B1(n17148), .B2(n20345), .A(n16626), .ZN(P2_U2843) );
  NAND2_X1 U20077 ( .A1(n14883), .A2(n16627), .ZN(n16628) );
  AND2_X1 U20078 ( .A1(n16613), .A2(n16628), .ZN(n17163) );
  NAND2_X1 U20079 ( .A1(n16629), .A2(n16736), .ZN(n16639) );
  OAI21_X1 U20080 ( .B1(n12628), .B2(n20335), .A(n13139), .ZN(n16630) );
  INV_X1 U20081 ( .A(n16630), .ZN(n16631) );
  OAI21_X1 U20082 ( .B1(n20292), .B2(n17159), .A(n16631), .ZN(n16632) );
  AOI21_X1 U20083 ( .B1(n20262), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n16632), .ZN(n16638) );
  OAI21_X1 U20084 ( .B1(n20351), .B2(n16635), .A(n16742), .ZN(n16634) );
  NAND2_X1 U20085 ( .A1(n16634), .A2(n16633), .ZN(n16637) );
  NAND3_X1 U20086 ( .A1(n16706), .A2(n17161), .A3(n16635), .ZN(n16636) );
  NAND4_X1 U20087 ( .A1(n16639), .A2(n16638), .A3(n16637), .A4(n16636), .ZN(
        n16640) );
  AOI21_X1 U20088 ( .B1(n17427), .B2(n20330), .A(n16640), .ZN(n16641) );
  OAI21_X1 U20089 ( .B1(n17429), .B2(n20345), .A(n16641), .ZN(P2_U2844) );
  NAND2_X1 U20090 ( .A1(n20350), .A2(n20313), .ZN(n16642) );
  XOR2_X1 U20091 ( .A(n17174), .B(n16642), .Z(n16649) );
  OAI22_X1 U20092 ( .A1(n16643), .A2(n20336), .B1(n17172), .B2(n20339), .ZN(
        n16644) );
  INV_X1 U20093 ( .A(n16644), .ZN(n16645) );
  OAI211_X1 U20094 ( .C1(n16646), .C2(n20335), .A(n16645), .B(n13139), .ZN(
        n16647) );
  AOI21_X1 U20095 ( .B1(n20344), .B2(P2_REIP_REG_10__SCAN_IN), .A(n16647), 
        .ZN(n16648) );
  OAI21_X1 U20096 ( .B1(n16649), .B2(n20351), .A(n16648), .ZN(n16650) );
  AOI21_X1 U20097 ( .B1(n17441), .B2(n20330), .A(n16650), .ZN(n16651) );
  OAI21_X1 U20098 ( .B1(n17438), .B2(n20345), .A(n16651), .ZN(P2_U2845) );
  INV_X1 U20099 ( .A(n17463), .ZN(n16663) );
  NOR2_X1 U20100 ( .A1(n16652), .A2(n20336), .ZN(n16662) );
  AOI21_X1 U20101 ( .B1(n20326), .B2(n16655), .A(n16692), .ZN(n16653) );
  OR2_X1 U20102 ( .A1(n16653), .A2(n17200), .ZN(n16660) );
  OAI21_X1 U20103 ( .B1(n21858), .B2(n20335), .A(n13139), .ZN(n16654) );
  AOI21_X1 U20104 ( .B1(n20344), .B2(P2_REIP_REG_8__SCAN_IN), .A(n16654), .ZN(
        n16659) );
  INV_X1 U20105 ( .A(n16655), .ZN(n16656) );
  NAND3_X1 U20106 ( .A1(n16706), .A2(n17200), .A3(n16656), .ZN(n16658) );
  OR2_X1 U20107 ( .A1(n20339), .A2(n13265), .ZN(n16657) );
  NAND4_X1 U20108 ( .A1(n16660), .A2(n16659), .A3(n16658), .A4(n16657), .ZN(
        n16661) );
  AOI211_X1 U20109 ( .C1(n16663), .C2(n20330), .A(n16662), .B(n16661), .ZN(
        n16664) );
  OAI21_X1 U20110 ( .B1(n17461), .B2(n20345), .A(n16664), .ZN(P2_U2847) );
  AOI21_X1 U20111 ( .B1(n20326), .B2(n16667), .A(n16692), .ZN(n16672) );
  AOI22_X1 U20112 ( .A1(n20262), .A2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n16736), .B2(n16665), .ZN(n16666) );
  OAI211_X1 U20113 ( .C1(n20990), .C2(n20292), .A(n16666), .B(n13139), .ZN(
        n16670) );
  INV_X1 U20114 ( .A(n17212), .ZN(n16668) );
  NOR3_X1 U20115 ( .A1(n16740), .A2(n16668), .A3(n16667), .ZN(n16669) );
  AOI211_X1 U20116 ( .C1(n20295), .C2(P2_EBX_REG_7__SCAN_IN), .A(n16670), .B(
        n16669), .ZN(n16671) );
  OAI21_X1 U20117 ( .B1(n16672), .B2(n17212), .A(n16671), .ZN(n16673) );
  AOI21_X1 U20118 ( .B1(n20330), .B2(n17479), .A(n16673), .ZN(n16674) );
  OAI21_X1 U20119 ( .B1(n17476), .B2(n20345), .A(n16674), .ZN(P2_U2848) );
  INV_X1 U20120 ( .A(n16681), .ZN(n16675) );
  NOR2_X1 U20121 ( .A1(n18101), .A2(n16675), .ZN(n16680) );
  OAI21_X1 U20122 ( .B1(n12626), .B2(n20335), .A(n13139), .ZN(n16676) );
  INV_X1 U20123 ( .A(n16676), .ZN(n16678) );
  INV_X1 U20124 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n20988) );
  OR2_X1 U20125 ( .A1(n20292), .A2(n20988), .ZN(n16677) );
  OAI211_X1 U20126 ( .C1(n20339), .C2(n18113), .A(n16678), .B(n16677), .ZN(
        n16679) );
  AOI21_X1 U20127 ( .B1(n16706), .B2(n16680), .A(n16679), .ZN(n16685) );
  OAI21_X1 U20128 ( .B1(n16681), .B2(n20351), .A(n16742), .ZN(n16683) );
  AOI22_X1 U20129 ( .A1(n16683), .A2(n18101), .B1(n16682), .B2(n16736), .ZN(
        n16684) );
  OAI211_X1 U20130 ( .C1(n17495), .C2(n20341), .A(n16685), .B(n16684), .ZN(
        n16686) );
  AOI21_X1 U20131 ( .B1(n18106), .B2(n20329), .A(n16686), .ZN(n16687) );
  INV_X1 U20132 ( .A(n16687), .ZN(P2_U2849) );
  NAND2_X1 U20133 ( .A1(n21047), .A2(n20348), .ZN(n16704) );
  NAND2_X1 U20134 ( .A1(n16690), .A2(n16689), .ZN(n16691) );
  NAND2_X1 U20135 ( .A1(n16688), .A2(n16691), .ZN(n21051) );
  INV_X1 U20136 ( .A(n21051), .ZN(n20378) );
  AOI21_X1 U20137 ( .B1(n20326), .B2(n16697), .A(n16692), .ZN(n16701) );
  INV_X1 U20138 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n20983) );
  OAI22_X1 U20139 ( .A1(n12259), .A2(n20335), .B1(n20983), .B2(n20292), .ZN(
        n16693) );
  AOI21_X1 U20140 ( .B1(n20262), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n16693), .ZN(n16694) );
  OAI21_X1 U20141 ( .B1(n16695), .B2(n20336), .A(n16694), .ZN(n16696) );
  INV_X1 U20142 ( .A(n16696), .ZN(n16700) );
  INV_X1 U20143 ( .A(n16697), .ZN(n16698) );
  NAND3_X1 U20144 ( .A1(n16706), .A2(n17243), .A3(n16698), .ZN(n16699) );
  OAI211_X1 U20145 ( .C1(n16701), .C2(n17243), .A(n16700), .B(n16699), .ZN(
        n16702) );
  AOI21_X1 U20146 ( .B1(n20330), .B2(n20378), .A(n16702), .ZN(n16703) );
  OAI211_X1 U20147 ( .C1(n20345), .C2(n14288), .A(n16704), .B(n16703), .ZN(
        P2_U2852) );
  NAND2_X1 U20148 ( .A1(n16705), .A2(n20348), .ZN(n16717) );
  OAI21_X1 U20149 ( .B1(n20351), .B2(n16722), .A(n16742), .ZN(n16714) );
  NOR2_X1 U20150 ( .A1(n21056), .A2(n20341), .ZN(n16713) );
  NAND3_X1 U20151 ( .A1(n16706), .A2(n16722), .A3(n10154), .ZN(n16710) );
  OAI22_X1 U20152 ( .A1(n16707), .A2(n20335), .B1(n20981), .B2(n20292), .ZN(
        n16708) );
  AOI21_X1 U20153 ( .B1(n20262), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n16708), .ZN(n16709) );
  OAI211_X1 U20154 ( .C1(n20336), .C2(n16711), .A(n16710), .B(n16709), .ZN(
        n16712) );
  AOI211_X1 U20155 ( .C1(n16715), .C2(n16714), .A(n16713), .B(n16712), .ZN(
        n16716) );
  OAI211_X1 U20156 ( .C1(n20345), .C2(n12275), .A(n16717), .B(n16716), .ZN(
        P2_U2853) );
  NAND2_X1 U20157 ( .A1(n16718), .A2(n20329), .ZN(n16731) );
  INV_X1 U20158 ( .A(n16739), .ZN(n17536) );
  INV_X1 U20159 ( .A(n16719), .ZN(n16720) );
  NAND2_X1 U20160 ( .A1(n17536), .A2(n16720), .ZN(n16721) );
  AND2_X1 U20161 ( .A1(n16722), .A2(n16721), .ZN(n16723) );
  AND2_X1 U20162 ( .A1(n20350), .A2(n16723), .ZN(n17542) );
  OAI22_X1 U20163 ( .A1(n22096), .A2(n20335), .B1(n20336), .B2(n16724), .ZN(
        n16726) );
  NOR2_X1 U20164 ( .A1(n20292), .A2(n20979), .ZN(n16725) );
  NOR2_X1 U20165 ( .A1(n16726), .A2(n16725), .ZN(n16728) );
  NAND2_X1 U20166 ( .A1(n21067), .A2(n20330), .ZN(n16727) );
  OAI211_X1 U20167 ( .C1(n13229), .C2(n20339), .A(n16728), .B(n16727), .ZN(
        n16729) );
  AOI21_X1 U20168 ( .B1(n17542), .B2(n20326), .A(n16729), .ZN(n16730) );
  OAI211_X1 U20169 ( .C1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n16742), .A(
        n16731), .B(n16730), .ZN(n16732) );
  AOI21_X1 U20170 ( .B1(n21072), .B2(n20348), .A(n16732), .ZN(n16733) );
  INV_X1 U20171 ( .A(n16733), .ZN(P2_U2854) );
  INV_X1 U20172 ( .A(n20348), .ZN(n16746) );
  AOI22_X1 U20173 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(n20344), .B1(n20330), 
        .B2(n16734), .ZN(n16738) );
  AOI22_X1 U20174 ( .A1(P2_EBX_REG_0__SCAN_IN), .A2(n20295), .B1(n16736), .B2(
        n16735), .ZN(n16737) );
  OAI211_X1 U20175 ( .C1(n16740), .C2(n16739), .A(n16738), .B(n16737), .ZN(
        n16744) );
  AOI21_X1 U20176 ( .B1(n16742), .B2(n20339), .A(n16741), .ZN(n16743) );
  AOI211_X1 U20177 ( .C1(n20329), .C2(n13822), .A(n16744), .B(n16743), .ZN(
        n16745) );
  OAI21_X1 U20178 ( .B1(n21079), .B2(n16746), .A(n16745), .ZN(P2_U2855) );
  INV_X1 U20179 ( .A(n16747), .ZN(n16845) );
  NAND2_X1 U20180 ( .A1(n9862), .A2(n16748), .ZN(n16844) );
  NAND3_X1 U20181 ( .A1(n16845), .A2(n16830), .A3(n16844), .ZN(n16750) );
  NAND2_X1 U20182 ( .A1(n9713), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n16749) );
  OAI211_X1 U20183 ( .C1(n16970), .C2(n9713), .A(n16750), .B(n16749), .ZN(
        P2_U2858) );
  NAND2_X1 U20184 ( .A1(n16752), .A2(n16751), .ZN(n16754) );
  XNOR2_X1 U20185 ( .A(n16754), .B(n16753), .ZN(n16861) );
  NOR2_X1 U20186 ( .A1(n16984), .A2(n9713), .ZN(n16755) );
  AOI21_X1 U20187 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n9713), .A(n16755), .ZN(
        n16756) );
  OAI21_X1 U20188 ( .B1(n16861), .B2(n16840), .A(n16756), .ZN(P2_U2859) );
  INV_X1 U20189 ( .A(n17260), .ZN(n16761) );
  AOI21_X1 U20190 ( .B1(n16758), .B2(n16757), .A(n9839), .ZN(n16862) );
  NAND2_X1 U20191 ( .A1(n16862), .A2(n16830), .ZN(n16760) );
  NAND2_X1 U20192 ( .A1(n9713), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n16759) );
  OAI211_X1 U20193 ( .C1(n16761), .C2(n9713), .A(n16760), .B(n16759), .ZN(
        P2_U2860) );
  AOI21_X1 U20194 ( .B1(n16764), .B2(n16763), .A(n16762), .ZN(n16868) );
  NAND2_X1 U20195 ( .A1(n16868), .A2(n16830), .ZN(n16766) );
  NAND2_X1 U20196 ( .A1(n17264), .A2(n16835), .ZN(n16765) );
  OAI211_X1 U20197 ( .C1(n16835), .C2(n16767), .A(n16766), .B(n16765), .ZN(
        P2_U2861) );
  OAI21_X1 U20198 ( .B1(n16770), .B2(n16769), .A(n16768), .ZN(n16884) );
  NOR2_X1 U20199 ( .A1(n17284), .A2(n9713), .ZN(n16771) );
  AOI21_X1 U20200 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n9713), .A(n16771), .ZN(
        n16772) );
  OAI21_X1 U20201 ( .B1(n16840), .B2(n16884), .A(n16772), .ZN(P2_U2862) );
  XNOR2_X1 U20202 ( .A(n16773), .B(n16774), .ZN(n16785) );
  NOR2_X1 U20203 ( .A1(n12901), .A2(n16775), .ZN(n16784) );
  NAND2_X1 U20204 ( .A1(n16785), .A2(n16784), .ZN(n16783) );
  OAI21_X1 U20205 ( .B1(n16776), .B2(n16773), .A(n16783), .ZN(n16780) );
  XOR2_X1 U20206 ( .A(n16778), .B(n16777), .Z(n16779) );
  XNOR2_X1 U20207 ( .A(n16780), .B(n16779), .ZN(n16892) );
  NOR2_X1 U20208 ( .A1(n17294), .A2(n9713), .ZN(n16781) );
  AOI21_X1 U20209 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n9713), .A(n16781), .ZN(
        n16782) );
  OAI21_X1 U20210 ( .B1(n16892), .B2(n16840), .A(n16782), .ZN(P2_U2863) );
  OAI21_X1 U20211 ( .B1(n16785), .B2(n16784), .A(n16783), .ZN(n16900) );
  NAND2_X1 U20212 ( .A1(n17310), .A2(n16835), .ZN(n16787) );
  NAND2_X1 U20213 ( .A1(n9713), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n16786) );
  OAI211_X1 U20214 ( .C1(n16900), .C2(n16840), .A(n16787), .B(n16786), .ZN(
        P2_U2864) );
  OAI21_X1 U20215 ( .B1(n9864), .B2(n16788), .A(n16773), .ZN(n16908) );
  INV_X1 U20216 ( .A(n16908), .ZN(n16789) );
  AOI22_X1 U20217 ( .A1(n16789), .A2(n16830), .B1(P2_EBX_REG_22__SCAN_IN), 
        .B2(n9713), .ZN(n16790) );
  OAI21_X1 U20218 ( .B1(n16791), .B2(n9713), .A(n16790), .ZN(P2_U2865) );
  NAND2_X1 U20219 ( .A1(n9713), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n16795) );
  AND2_X1 U20220 ( .A1(n16797), .A2(n16792), .ZN(n16793) );
  NOR2_X1 U20221 ( .A1(n9864), .A2(n16793), .ZN(n16912) );
  NAND2_X1 U20222 ( .A1(n16912), .A2(n16830), .ZN(n16794) );
  OAI211_X1 U20223 ( .C1(n17050), .C2(n9713), .A(n16795), .B(n16794), .ZN(
        P2_U2866) );
  INV_X1 U20224 ( .A(n16796), .ZN(n16799) );
  INV_X1 U20225 ( .A(n16797), .ZN(n16798) );
  AOI21_X1 U20226 ( .B1(n16800), .B2(n16799), .A(n16798), .ZN(n16917) );
  AOI22_X1 U20227 ( .A1(n16917), .A2(n16830), .B1(P2_EBX_REG_20__SCAN_IN), 
        .B2(n9713), .ZN(n16801) );
  OAI21_X1 U20228 ( .B1(n17335), .B2(n9713), .A(n16801), .ZN(P2_U2867) );
  AND2_X1 U20229 ( .A1(n16552), .A2(n16802), .ZN(n16803) );
  OR2_X1 U20230 ( .A1(n16803), .A2(n16535), .ZN(n17347) );
  AOI21_X1 U20231 ( .B1(n16804), .B2(n16807), .A(n16796), .ZN(n16936) );
  AOI22_X1 U20232 ( .A1(n16936), .A2(n16830), .B1(P2_EBX_REG_19__SCAN_IN), 
        .B2(n9713), .ZN(n16805) );
  OAI21_X1 U20233 ( .B1(n17347), .B2(n9713), .A(n16805), .ZN(P2_U2868) );
  OAI21_X1 U20234 ( .B1(n16806), .B2(n16808), .A(n16807), .ZN(n16944) );
  INV_X1 U20235 ( .A(n16944), .ZN(n16809) );
  AOI22_X1 U20236 ( .A1(n16809), .A2(n16830), .B1(P2_EBX_REG_18__SCAN_IN), 
        .B2(n9713), .ZN(n16810) );
  OAI21_X1 U20237 ( .B1(n17357), .B2(n9713), .A(n16810), .ZN(P2_U2869) );
  NAND2_X1 U20238 ( .A1(n9713), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n16814) );
  AND2_X1 U20239 ( .A1(n16816), .A2(n16811), .ZN(n16812) );
  NOR2_X1 U20240 ( .A1(n16806), .A2(n16812), .ZN(n16948) );
  NAND2_X1 U20241 ( .A1(n16948), .A2(n16830), .ZN(n16813) );
  OAI211_X1 U20242 ( .C1(n17370), .C2(n9713), .A(n16814), .B(n16813), .ZN(
        P2_U2870) );
  INV_X1 U20243 ( .A(n16815), .ZN(n16820) );
  NOR2_X1 U20244 ( .A1(n16821), .A2(n16820), .ZN(n16818) );
  OAI21_X1 U20245 ( .B1(n16818), .B2(n16817), .A(n16816), .ZN(n20363) );
  MUX2_X1 U20246 ( .A(n17374), .B(n12847), .S(n9713), .Z(n16819) );
  OAI21_X1 U20247 ( .B1(n16840), .B2(n20363), .A(n16819), .ZN(P2_U2871) );
  XNOR2_X1 U20248 ( .A(n16821), .B(n16820), .ZN(n16827) );
  NAND2_X1 U20249 ( .A1(n14646), .A2(n16822), .ZN(n16823) );
  NAND2_X1 U20250 ( .A1(n16824), .A2(n16823), .ZN(n20288) );
  NOR2_X1 U20251 ( .A1(n20288), .A2(n9713), .ZN(n16825) );
  AOI21_X1 U20252 ( .B1(P2_EBX_REG_15__SCAN_IN), .B2(n9713), .A(n16825), .ZN(
        n16826) );
  OAI21_X1 U20253 ( .B1(n16827), .B2(n16840), .A(n16826), .ZN(P2_U2872) );
  INV_X1 U20254 ( .A(n16837), .ZN(n16828) );
  NOR2_X1 U20255 ( .A1(n16836), .A2(n16828), .ZN(n16832) );
  OAI211_X1 U20256 ( .C1(n16832), .C2(n16831), .A(n16830), .B(n16829), .ZN(
        n16834) );
  INV_X1 U20257 ( .A(n17148), .ZN(n17415) );
  NAND2_X1 U20258 ( .A1(n17415), .A2(n16835), .ZN(n16833) );
  OAI211_X1 U20259 ( .C1(n12832), .C2(n16835), .A(n16834), .B(n16833), .ZN(
        P2_U2875) );
  XOR2_X1 U20260 ( .A(n16837), .B(n16836), .Z(n16841) );
  NOR2_X1 U20261 ( .A1(n17429), .A2(n9713), .ZN(n16838) );
  AOI21_X1 U20262 ( .B1(P2_EBX_REG_11__SCAN_IN), .B2(n9713), .A(n16838), .ZN(
        n16839) );
  OAI21_X1 U20263 ( .B1(n16841), .B2(n16840), .A(n16839), .ZN(P2_U2876) );
  NAND2_X1 U20264 ( .A1(n15361), .A2(n20385), .ZN(n16843) );
  AOI22_X1 U20265 ( .A1(n20362), .A2(BUF2_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n16938), .ZN(n16842) );
  OAI211_X1 U20266 ( .C1(n18147), .C2(n16941), .A(n16843), .B(n16842), .ZN(
        P2_U2888) );
  NAND3_X1 U20267 ( .A1(n16845), .A2(n20373), .A3(n16844), .ZN(n16852) );
  INV_X1 U20268 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n16849) );
  NAND2_X1 U20269 ( .A1(n20361), .A2(BUF1_REG_29__SCAN_IN), .ZN(n16848) );
  AOI22_X1 U20270 ( .A1(n20360), .A2(n16846), .B1(P2_EAX_REG_29__SCAN_IN), 
        .B2(n16938), .ZN(n16847) );
  OAI211_X1 U20271 ( .C1(n16849), .C2(n16921), .A(n16848), .B(n16847), .ZN(
        n16850) );
  INV_X1 U20272 ( .A(n16850), .ZN(n16851) );
  OAI211_X1 U20273 ( .C1(n16853), .C2(n16934), .A(n16852), .B(n16851), .ZN(
        P2_U2890) );
  INV_X1 U20274 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n16857) );
  NAND2_X1 U20275 ( .A1(n20361), .A2(BUF1_REG_28__SCAN_IN), .ZN(n16856) );
  AOI22_X1 U20276 ( .A1(n20360), .A2(n16854), .B1(P2_EAX_REG_28__SCAN_IN), 
        .B2(n16938), .ZN(n16855) );
  OAI211_X1 U20277 ( .C1(n16857), .C2(n16921), .A(n16856), .B(n16855), .ZN(
        n16858) );
  AOI21_X1 U20278 ( .B1(n16859), .B2(n20385), .A(n16858), .ZN(n16860) );
  OAI21_X1 U20279 ( .B1(n16861), .B2(n20389), .A(n16860), .ZN(P2_U2891) );
  NAND2_X1 U20280 ( .A1(n16862), .A2(n20373), .ZN(n16867) );
  AOI22_X1 U20281 ( .A1(n20360), .A2(n16863), .B1(P2_EAX_REG_27__SCAN_IN), 
        .B2(n16938), .ZN(n16864) );
  OAI21_X1 U20282 ( .B1(n16941), .B2(n18153), .A(n16864), .ZN(n16865) );
  AOI21_X1 U20283 ( .B1(n20362), .B2(BUF2_REG_27__SCAN_IN), .A(n16865), .ZN(
        n16866) );
  OAI211_X1 U20284 ( .C1(n17253), .C2(n16934), .A(n16867), .B(n16866), .ZN(
        P2_U2892) );
  INV_X1 U20285 ( .A(n16868), .ZN(n16876) );
  INV_X1 U20286 ( .A(n17272), .ZN(n16874) );
  INV_X1 U20287 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n16872) );
  NAND2_X1 U20288 ( .A1(n20361), .A2(BUF1_REG_26__SCAN_IN), .ZN(n16871) );
  AOI22_X1 U20289 ( .A1(n20360), .A2(n16869), .B1(P2_EAX_REG_26__SCAN_IN), 
        .B2(n16938), .ZN(n16870) );
  OAI211_X1 U20290 ( .C1(n16872), .C2(n16921), .A(n16871), .B(n16870), .ZN(
        n16873) );
  AOI21_X1 U20291 ( .B1(n16874), .B2(n20385), .A(n16873), .ZN(n16875) );
  OAI21_X1 U20292 ( .B1(n16876), .B2(n20389), .A(n16875), .ZN(P2_U2893) );
  INV_X1 U20293 ( .A(n17279), .ZN(n16882) );
  INV_X1 U20294 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n16880) );
  NAND2_X1 U20295 ( .A1(n20361), .A2(BUF1_REG_25__SCAN_IN), .ZN(n16879) );
  AOI22_X1 U20296 ( .A1(n20360), .A2(n16877), .B1(P2_EAX_REG_25__SCAN_IN), 
        .B2(n16938), .ZN(n16878) );
  OAI211_X1 U20297 ( .C1(n16880), .C2(n16921), .A(n16879), .B(n16878), .ZN(
        n16881) );
  AOI21_X1 U20298 ( .B1(n16882), .B2(n20385), .A(n16881), .ZN(n16883) );
  OAI21_X1 U20299 ( .B1(n20389), .B2(n16884), .A(n16883), .ZN(P2_U2894) );
  INV_X1 U20300 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n16888) );
  NAND2_X1 U20301 ( .A1(n20361), .A2(BUF1_REG_24__SCAN_IN), .ZN(n16887) );
  AOI22_X1 U20302 ( .A1(n20360), .A2(n16885), .B1(P2_EAX_REG_24__SCAN_IN), 
        .B2(n16938), .ZN(n16886) );
  OAI211_X1 U20303 ( .C1(n16888), .C2(n16921), .A(n16887), .B(n16886), .ZN(
        n16889) );
  AOI21_X1 U20304 ( .B1(n16890), .B2(n20385), .A(n16889), .ZN(n16891) );
  OAI21_X1 U20305 ( .B1(n16892), .B2(n20389), .A(n16891), .ZN(P2_U2895) );
  INV_X1 U20306 ( .A(n17307), .ZN(n16898) );
  INV_X1 U20307 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n16896) );
  NAND2_X1 U20308 ( .A1(n20361), .A2(BUF1_REG_23__SCAN_IN), .ZN(n16895) );
  AOI22_X1 U20309 ( .A1(n20360), .A2(n16893), .B1(P2_EAX_REG_23__SCAN_IN), 
        .B2(n16938), .ZN(n16894) );
  OAI211_X1 U20310 ( .C1(n16896), .C2(n16921), .A(n16895), .B(n16894), .ZN(
        n16897) );
  AOI21_X1 U20311 ( .B1(n16898), .B2(n20385), .A(n16897), .ZN(n16899) );
  OAI21_X1 U20312 ( .B1(n20389), .B2(n16900), .A(n16899), .ZN(P2_U2896) );
  INV_X1 U20313 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n16904) );
  NAND2_X1 U20314 ( .A1(n20361), .A2(BUF1_REG_22__SCAN_IN), .ZN(n16903) );
  AOI22_X1 U20315 ( .A1(n20360), .A2(n16901), .B1(P2_EAX_REG_22__SCAN_IN), 
        .B2(n16938), .ZN(n16902) );
  OAI211_X1 U20316 ( .C1(n16904), .C2(n16921), .A(n16903), .B(n16902), .ZN(
        n16905) );
  AOI21_X1 U20317 ( .B1(n16906), .B2(n20385), .A(n16905), .ZN(n16907) );
  OAI21_X1 U20318 ( .B1(n20389), .B2(n16908), .A(n16907), .ZN(P2_U2897) );
  NAND2_X1 U20319 ( .A1(n16909), .A2(n20385), .ZN(n16916) );
  NAND2_X1 U20320 ( .A1(n16938), .A2(P2_EAX_REG_21__SCAN_IN), .ZN(n16910) );
  OAI21_X1 U20321 ( .B1(n16946), .B2(n20443), .A(n16910), .ZN(n16911) );
  AOI21_X1 U20322 ( .B1(n20361), .B2(BUF1_REG_21__SCAN_IN), .A(n16911), .ZN(
        n16915) );
  NAND2_X1 U20323 ( .A1(n16912), .A2(n20373), .ZN(n16914) );
  NAND2_X1 U20324 ( .A1(n20362), .A2(BUF2_REG_21__SCAN_IN), .ZN(n16913) );
  NAND4_X1 U20325 ( .A1(n16916), .A2(n16915), .A3(n16914), .A4(n16913), .ZN(
        P2_U2898) );
  INV_X1 U20326 ( .A(n16917), .ZN(n16926) );
  INV_X1 U20327 ( .A(n17332), .ZN(n16924) );
  INV_X1 U20328 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n16922) );
  NAND2_X1 U20329 ( .A1(n20361), .A2(BUF1_REG_20__SCAN_IN), .ZN(n16920) );
  AOI22_X1 U20330 ( .A1(n20360), .A2(n16918), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n16938), .ZN(n16919) );
  OAI211_X1 U20331 ( .C1(n16922), .C2(n16921), .A(n16920), .B(n16919), .ZN(
        n16923) );
  AOI21_X1 U20332 ( .B1(n16924), .B2(n20385), .A(n16923), .ZN(n16925) );
  OAI21_X1 U20333 ( .B1(n20389), .B2(n16926), .A(n16925), .ZN(P2_U2899) );
  NAND2_X1 U20334 ( .A1(n16565), .A2(n16927), .ZN(n16928) );
  NAND2_X1 U20335 ( .A1(n16929), .A2(n16928), .ZN(n20271) );
  NAND2_X1 U20336 ( .A1(n16938), .A2(P2_EAX_REG_19__SCAN_IN), .ZN(n16930) );
  OAI21_X1 U20337 ( .B1(n16946), .B2(n20437), .A(n16930), .ZN(n16931) );
  AOI21_X1 U20338 ( .B1(n20361), .B2(BUF1_REG_19__SCAN_IN), .A(n16931), .ZN(
        n16933) );
  NAND2_X1 U20339 ( .A1(n20362), .A2(BUF2_REG_19__SCAN_IN), .ZN(n16932) );
  OAI211_X1 U20340 ( .C1(n20271), .C2(n16934), .A(n16933), .B(n16932), .ZN(
        n16935) );
  AOI21_X1 U20341 ( .B1(n20373), .B2(n16936), .A(n16935), .ZN(n16937) );
  INV_X1 U20342 ( .A(n16937), .ZN(P2_U2900) );
  NAND2_X1 U20343 ( .A1(n20362), .A2(BUF2_REG_18__SCAN_IN), .ZN(n16940) );
  AOI22_X1 U20344 ( .A1(n20360), .A2(n20434), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n16938), .ZN(n16939) );
  OAI211_X1 U20345 ( .C1(n18168), .C2(n16941), .A(n16940), .B(n16939), .ZN(
        n16942) );
  AOI21_X1 U20346 ( .B1(n17353), .B2(n20385), .A(n16942), .ZN(n16943) );
  OAI21_X1 U20347 ( .B1(n20389), .B2(n16944), .A(n16943), .ZN(P2_U2901) );
  NAND2_X1 U20348 ( .A1(n17368), .A2(n20385), .ZN(n16952) );
  NAND2_X1 U20349 ( .A1(n16938), .A2(P2_EAX_REG_17__SCAN_IN), .ZN(n16945) );
  OAI21_X1 U20350 ( .B1(n16946), .B2(n20394), .A(n16945), .ZN(n16947) );
  AOI21_X1 U20351 ( .B1(n20361), .B2(BUF1_REG_17__SCAN_IN), .A(n16947), .ZN(
        n16951) );
  NAND2_X1 U20352 ( .A1(n16948), .A2(n20373), .ZN(n16950) );
  NAND2_X1 U20353 ( .A1(n20362), .A2(BUF2_REG_17__SCAN_IN), .ZN(n16949) );
  NAND4_X1 U20354 ( .A1(n16952), .A2(n16951), .A3(n16950), .A4(n16949), .ZN(
        P2_U2902) );
  OR2_X1 U20355 ( .A1(n14806), .A2(n16953), .ZN(n16954) );
  AND2_X1 U20356 ( .A1(n16588), .A2(n16954), .ZN(n20285) );
  INV_X1 U20357 ( .A(n20285), .ZN(n16956) );
  OAI222_X1 U20358 ( .A1(n16956), .A2(n16963), .B1(n16965), .B2(n20398), .C1(
        n16955), .C2(n20393), .ZN(P2_U2904) );
  AOI21_X1 U20359 ( .B1(n21056), .B2(n21058), .A(n16957), .ZN(n20381) );
  XOR2_X1 U20360 ( .A(n21051), .B(n21047), .Z(n20380) );
  NOR2_X1 U20361 ( .A1(n20381), .A2(n20380), .ZN(n20379) );
  NOR2_X1 U20362 ( .A1(n21047), .A2(n20378), .ZN(n16961) );
  NAND2_X1 U20363 ( .A1(n16688), .A2(n16959), .ZN(n16960) );
  NAND2_X1 U20364 ( .A1(n16958), .A2(n16960), .ZN(n20369) );
  OAI21_X1 U20365 ( .B1(n20379), .B2(n16961), .A(n20369), .ZN(n20371) );
  NAND3_X1 U20366 ( .A1(n20371), .A2(n20373), .A3(n20372), .ZN(n16969) );
  XOR2_X1 U20367 ( .A(n16958), .B(n16962), .Z(n20331) );
  INV_X1 U20368 ( .A(n16963), .ZN(n16967) );
  INV_X1 U20369 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n16964) );
  OAI22_X1 U20370 ( .A1(n20393), .A2(n20443), .B1(n16965), .B2(n16964), .ZN(
        n16966) );
  AOI21_X1 U20371 ( .B1(n20331), .B2(n16967), .A(n16966), .ZN(n16968) );
  NAND2_X1 U20372 ( .A1(n16969), .A2(n16968), .ZN(P2_U2914) );
  NOR2_X1 U20373 ( .A1(n18112), .A2(n16972), .ZN(n16973) );
  AOI211_X1 U20374 ( .C1(n16975), .C2(n18102), .A(n16974), .B(n16973), .ZN(
        n16976) );
  NOR2_X1 U20375 ( .A1(n17244), .A2(n16980), .ZN(n16981) );
  AOI211_X1 U20376 ( .C1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n17214), .A(
        n16982), .B(n16981), .ZN(n16983) );
  OAI21_X1 U20377 ( .B1(n16984), .B2(n17242), .A(n16983), .ZN(n16985) );
  AOI21_X1 U20378 ( .B1(n16986), .B2(n18108), .A(n16985), .ZN(n16987) );
  OAI21_X1 U20379 ( .B1(n16988), .B2(n17252), .A(n16987), .ZN(P2_U2986) );
  XNOR2_X1 U20380 ( .A(n16989), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17263) );
  NAND2_X1 U20381 ( .A1(n18102), .A2(n16990), .ZN(n16991) );
  NAND2_X1 U20382 ( .A1(n20343), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n17254) );
  OAI211_X1 U20383 ( .C1(n22083), .C2(n18112), .A(n16991), .B(n17254), .ZN(
        n16993) );
  OAI21_X1 U20384 ( .B1(n17263), .B2(n17252), .A(n16994), .ZN(P2_U2987) );
  INV_X1 U20385 ( .A(n17008), .ZN(n16995) );
  INV_X1 U20386 ( .A(n16997), .ZN(n16998) );
  NAND2_X1 U20387 ( .A1(n16999), .A2(n16998), .ZN(n17276) );
  AOI21_X1 U20388 ( .B1(n17267), .B2(n17000), .A(n17001), .ZN(n17274) );
  NAND2_X1 U20389 ( .A1(n17264), .A2(n18107), .ZN(n17003) );
  NOR2_X1 U20390 ( .A1(n13139), .A2(n21023), .ZN(n17269) );
  AOI21_X1 U20391 ( .B1(n17214), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n17269), .ZN(n17002) );
  OAI211_X1 U20392 ( .C1(n17244), .C2(n17004), .A(n17003), .B(n17002), .ZN(
        n17005) );
  AOI21_X1 U20393 ( .B1(n18108), .B2(n17274), .A(n17005), .ZN(n17006) );
  OAI21_X1 U20394 ( .B1(n17252), .B2(n17276), .A(n17006), .ZN(P2_U2988) );
  NAND2_X1 U20395 ( .A1(n17008), .A2(n17007), .ZN(n17009) );
  XNOR2_X1 U20396 ( .A(n17010), .B(n17009), .ZN(n17287) );
  NAND2_X1 U20397 ( .A1(n20343), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n17277) );
  OAI21_X1 U20398 ( .B1(n18112), .B2(n17012), .A(n17277), .ZN(n17013) );
  AOI21_X1 U20399 ( .B1(n18102), .B2(n17014), .A(n17013), .ZN(n17015) );
  OAI21_X1 U20400 ( .B1(n17284), .B2(n17242), .A(n17015), .ZN(n17016) );
  AOI21_X1 U20401 ( .B1(n17286), .B2(n18108), .A(n17016), .ZN(n17017) );
  OAI21_X1 U20402 ( .B1(n17252), .B2(n17287), .A(n17017), .ZN(P2_U2989) );
  XNOR2_X1 U20403 ( .A(n17018), .B(n10338), .ZN(n17019) );
  XNOR2_X1 U20404 ( .A(n17020), .B(n17019), .ZN(n17299) );
  NOR2_X1 U20405 ( .A1(n13139), .A2(n21019), .ZN(n17288) );
  NOR2_X1 U20406 ( .A1(n17244), .A2(n17022), .ZN(n17023) );
  AOI211_X1 U20407 ( .C1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(n17214), .A(
        n17288), .B(n17023), .ZN(n17024) );
  OAI21_X1 U20408 ( .B1(n17294), .B2(n17242), .A(n17024), .ZN(n17025) );
  OAI21_X1 U20409 ( .B1(n17034), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n17021), .ZN(n17312) );
  XNOR2_X1 U20410 ( .A(n17027), .B(n17026), .ZN(n17300) );
  NOR2_X1 U20411 ( .A1(n17300), .A2(n17252), .ZN(n17032) );
  NAND2_X1 U20412 ( .A1(n18102), .A2(n17028), .ZN(n17029) );
  NAND2_X1 U20413 ( .A1(n20343), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n17303) );
  OAI211_X1 U20414 ( .C1(n17030), .C2(n18112), .A(n17029), .B(n17303), .ZN(
        n17031) );
  AOI211_X1 U20415 ( .C1(n17310), .C2(n18107), .A(n17032), .B(n17031), .ZN(
        n17033) );
  OAI21_X1 U20416 ( .B1(n17218), .B2(n17312), .A(n17033), .ZN(P2_U2991) );
  AND2_X1 U20417 ( .A1(n17038), .A2(n17037), .ZN(n17039) );
  XNOR2_X1 U20418 ( .A(n17040), .B(n17039), .ZN(n17323) );
  NOR2_X1 U20419 ( .A1(n17323), .A2(n17252), .ZN(n17045) );
  NAND2_X1 U20420 ( .A1(n17320), .A2(n18107), .ZN(n17042) );
  NOR2_X1 U20421 ( .A1(n13139), .A2(n21015), .ZN(n17315) );
  AOI21_X1 U20422 ( .B1(n17214), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n17315), .ZN(n17041) );
  OAI211_X1 U20423 ( .C1(n17244), .C2(n17043), .A(n17042), .B(n17041), .ZN(
        n17044) );
  AOI211_X1 U20424 ( .C1(n17313), .C2(n18108), .A(n17045), .B(n17044), .ZN(
        n17046) );
  INV_X1 U20425 ( .A(n17046), .ZN(P2_U2992) );
  NAND2_X1 U20426 ( .A1(n17047), .A2(n18105), .ZN(n17055) );
  OAI21_X1 U20427 ( .B1(n18112), .B2(n17049), .A(n17048), .ZN(n17052) );
  NOR2_X1 U20428 ( .A1(n17050), .A2(n17242), .ZN(n17051) );
  AOI211_X1 U20429 ( .C1(n17053), .C2(n18102), .A(n17052), .B(n17051), .ZN(
        n17054) );
  OAI211_X1 U20430 ( .C1(n17218), .C2(n17056), .A(n17055), .B(n17054), .ZN(
        P2_U2993) );
  AND2_X1 U20431 ( .A1(n17058), .A2(n17057), .ZN(n17059) );
  OAI22_X1 U20432 ( .A1(n17060), .A2(n10603), .B1(n10388), .B2(n17059), .ZN(
        n17339) );
  NOR2_X1 U20433 ( .A1(n17335), .A2(n17242), .ZN(n17064) );
  NAND2_X1 U20434 ( .A1(n20343), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n17331) );
  NAND2_X1 U20435 ( .A1(n17214), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n17061) );
  OAI211_X1 U20436 ( .C1(n17244), .C2(n17062), .A(n17331), .B(n17061), .ZN(
        n17063) );
  OAI21_X1 U20437 ( .B1(n17339), .B2(n17252), .A(n17065), .ZN(P2_U2994) );
  NAND2_X1 U20438 ( .A1(n17067), .A2(n17066), .ZN(n17068) );
  INV_X1 U20439 ( .A(n17347), .ZN(n20274) );
  INV_X1 U20440 ( .A(n17069), .ZN(n20267) );
  NAND2_X1 U20441 ( .A1(n18102), .A2(n20267), .ZN(n17070) );
  OR2_X1 U20442 ( .A1(n13139), .A2(n21010), .ZN(n17342) );
  OAI211_X1 U20443 ( .C1(n17071), .C2(n18112), .A(n17070), .B(n17342), .ZN(
        n17073) );
  OAI21_X1 U20444 ( .B1(n17350), .B2(n17252), .A(n17074), .ZN(P2_U2995) );
  NAND2_X1 U20445 ( .A1(n17076), .A2(n17075), .ZN(n17077) );
  NAND2_X1 U20446 ( .A1(n17080), .A2(n18107), .ZN(n17083) );
  NOR2_X1 U20447 ( .A1(n13139), .A2(n17081), .ZN(n17352) );
  AOI21_X1 U20448 ( .B1(n17214), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n17352), .ZN(n17082) );
  OAI211_X1 U20449 ( .C1(n17244), .C2(n17084), .A(n17083), .B(n17082), .ZN(
        n17085) );
  AOI21_X1 U20450 ( .B1(n17359), .B2(n18108), .A(n17085), .ZN(n17086) );
  XOR2_X1 U20451 ( .A(n17088), .B(n17087), .Z(n17371) );
  INV_X1 U20452 ( .A(n17370), .ZN(n17092) );
  NOR2_X1 U20453 ( .A1(n13139), .A2(n21007), .ZN(n17367) );
  AOI21_X1 U20454 ( .B1(n17214), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n17367), .ZN(n17089) );
  OAI21_X1 U20455 ( .B1(n17244), .B2(n17090), .A(n17089), .ZN(n17091) );
  AOI21_X1 U20456 ( .B1(n17092), .B2(n18107), .A(n17091), .ZN(n17096) );
  AND2_X1 U20457 ( .A1(n17381), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17365) );
  INV_X1 U20458 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17376) );
  OAI211_X1 U20459 ( .C1(n17101), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n18108), .B(n17094), .ZN(n17095) );
  OAI211_X1 U20460 ( .C1(n17371), .C2(n17252), .A(n17096), .B(n17095), .ZN(
        P2_U2997) );
  XNOR2_X1 U20461 ( .A(n17098), .B(n17097), .ZN(n17378) );
  INV_X1 U20462 ( .A(n17374), .ZN(n17104) );
  NOR2_X1 U20463 ( .A1(n13139), .A2(n21005), .ZN(n17372) );
  AOI21_X1 U20464 ( .B1(n17214), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n17372), .ZN(n17099) );
  OAI21_X1 U20465 ( .B1(n17100), .B2(n17244), .A(n17099), .ZN(n17103) );
  AND2_X1 U20466 ( .A1(n17106), .A2(n17131), .ZN(n17119) );
  NOR2_X1 U20467 ( .A1(n17119), .A2(n17107), .ZN(n17124) );
  INV_X1 U20468 ( .A(n17123), .ZN(n17108) );
  NOR2_X1 U20469 ( .A1(n17124), .A2(n17108), .ZN(n17112) );
  NAND2_X1 U20470 ( .A1(n17110), .A2(n17109), .ZN(n17111) );
  XNOR2_X1 U20471 ( .A(n17112), .B(n17111), .ZN(n17387) );
  NOR2_X1 U20472 ( .A1(n13139), .A2(n21003), .ZN(n17382) );
  NOR2_X1 U20473 ( .A1(n18112), .A2(n20277), .ZN(n17114) );
  AOI211_X1 U20474 ( .C1(n20281), .C2(n18102), .A(n17382), .B(n17114), .ZN(
        n17115) );
  OAI21_X1 U20475 ( .B1(n20288), .B2(n17242), .A(n17115), .ZN(n17116) );
  OAI21_X1 U20476 ( .B1(n17387), .B2(n17252), .A(n17117), .ZN(P2_U2999) );
  OAI21_X1 U20477 ( .B1(n17137), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n17118), .ZN(n17400) );
  INV_X1 U20478 ( .A(n17119), .ZN(n17120) );
  AOI21_X1 U20479 ( .B1(n17121), .B2(n17123), .A(n17120), .ZN(n17122) );
  AOI21_X1 U20480 ( .B1(n17124), .B2(n17123), .A(n17122), .ZN(n17397) );
  NOR2_X1 U20481 ( .A1(n13139), .A2(n17125), .ZN(n17391) );
  NOR2_X1 U20482 ( .A1(n17244), .A2(n17126), .ZN(n17127) );
  AOI211_X1 U20483 ( .C1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .C2(n17214), .A(
        n17391), .B(n17127), .ZN(n17128) );
  OAI21_X1 U20484 ( .B1(n17395), .B2(n17242), .A(n17128), .ZN(n17129) );
  AOI21_X1 U20485 ( .B1(n17397), .B2(n18105), .A(n17129), .ZN(n17130) );
  OAI21_X1 U20486 ( .B1(n17400), .B2(n17218), .A(n17130), .ZN(P2_U3000) );
  NAND2_X1 U20487 ( .A1(n17132), .A2(n17131), .ZN(n17136) );
  INV_X1 U20488 ( .A(n17155), .ZN(n17133) );
  AOI21_X1 U20489 ( .B1(n17156), .B2(n17154), .A(n17133), .ZN(n17146) );
  INV_X1 U20490 ( .A(n17145), .ZN(n17134) );
  AOI21_X1 U20491 ( .B1(n17146), .B2(n17144), .A(n17134), .ZN(n17135) );
  XOR2_X1 U20492 ( .A(n17136), .B(n17135), .Z(n17411) );
  AOI21_X1 U20493 ( .B1(n17402), .B2(n17143), .A(n17137), .ZN(n17401) );
  NAND2_X1 U20494 ( .A1(n17401), .A2(n18108), .ZN(n17142) );
  INV_X1 U20495 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n21000) );
  NOR2_X1 U20496 ( .A1(n20260), .A2(n21000), .ZN(n17404) );
  AOI21_X1 U20497 ( .B1(n17214), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n17404), .ZN(n17138) );
  OAI21_X1 U20498 ( .B1(n17244), .B2(n20297), .A(n17138), .ZN(n17139) );
  AOI21_X1 U20499 ( .B1(n17140), .B2(n18107), .A(n17139), .ZN(n17141) );
  OAI21_X1 U20500 ( .B1(n17158), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n17143), .ZN(n17423) );
  NAND2_X1 U20501 ( .A1(n17145), .A2(n17144), .ZN(n17147) );
  XOR2_X1 U20502 ( .A(n17147), .B(n17146), .Z(n17421) );
  NOR2_X1 U20503 ( .A1(n17148), .A2(n17242), .ZN(n17152) );
  NAND2_X1 U20504 ( .A1(n20343), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n17412) );
  NAND2_X1 U20505 ( .A1(n17214), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17149) );
  OAI211_X1 U20506 ( .C1(n17244), .C2(n17150), .A(n17412), .B(n17149), .ZN(
        n17151) );
  AOI211_X1 U20507 ( .C1(n17421), .C2(n18105), .A(n17152), .B(n17151), .ZN(
        n17153) );
  OAI21_X1 U20508 ( .B1(n17423), .B2(n17218), .A(n17153), .ZN(P2_U3002) );
  NAND2_X1 U20509 ( .A1(n17155), .A2(n17154), .ZN(n17157) );
  XOR2_X1 U20510 ( .A(n17157), .B(n17156), .Z(n17436) );
  NAND2_X1 U20511 ( .A1(n17424), .A2(n18108), .ZN(n17165) );
  NOR2_X1 U20512 ( .A1(n20260), .A2(n17159), .ZN(n17426) );
  AOI21_X1 U20513 ( .B1(n17214), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n17426), .ZN(n17160) );
  OAI21_X1 U20514 ( .B1(n17244), .B2(n17161), .A(n17160), .ZN(n17162) );
  AOI21_X1 U20515 ( .B1(n17163), .B2(n18107), .A(n17162), .ZN(n17164) );
  OAI211_X1 U20516 ( .C1(n17436), .C2(n17252), .A(n17165), .B(n17164), .ZN(
        P2_U3003) );
  XNOR2_X1 U20517 ( .A(n17449), .B(n17432), .ZN(n17448) );
  NAND2_X1 U20518 ( .A1(n17166), .A2(n17183), .ZN(n17170) );
  NAND2_X1 U20519 ( .A1(n17168), .A2(n17167), .ZN(n17169) );
  XNOR2_X1 U20520 ( .A(n17170), .B(n17169), .ZN(n17446) );
  INV_X1 U20521 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n17171) );
  NOR2_X1 U20522 ( .A1(n20260), .A2(n17171), .ZN(n17440) );
  NOR2_X1 U20523 ( .A1(n18112), .A2(n17172), .ZN(n17173) );
  AOI211_X1 U20524 ( .C1(n17174), .C2(n18102), .A(n17440), .B(n17173), .ZN(
        n17175) );
  OAI21_X1 U20525 ( .B1(n17438), .B2(n17242), .A(n17175), .ZN(n17176) );
  AOI21_X1 U20526 ( .B1(n17446), .B2(n18105), .A(n17176), .ZN(n17177) );
  OAI21_X1 U20527 ( .B1(n17448), .B2(n17218), .A(n17177), .ZN(P2_U3004) );
  NAND2_X1 U20528 ( .A1(n17179), .A2(n17178), .ZN(n17211) );
  INV_X1 U20529 ( .A(n17180), .ZN(n17182) );
  OAI21_X1 U20530 ( .B1(n17211), .B2(n17182), .A(n17181), .ZN(n17186) );
  NAND2_X1 U20531 ( .A1(n17184), .A2(n17183), .ZN(n17185) );
  XNOR2_X1 U20532 ( .A(n17186), .B(n17185), .ZN(n17460) );
  INV_X1 U20533 ( .A(n17364), .ZN(n17187) );
  NAND2_X1 U20534 ( .A1(n17187), .A2(n17456), .ZN(n17450) );
  NAND3_X1 U20535 ( .A1(n17450), .A2(n18108), .A3(n17449), .ZN(n17191) );
  NAND2_X1 U20536 ( .A1(n20343), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n17452) );
  OAI21_X1 U20537 ( .B1(n18112), .B2(n20307), .A(n17452), .ZN(n17189) );
  NOR2_X1 U20538 ( .A1(n20316), .A2(n17242), .ZN(n17188) );
  AOI211_X1 U20539 ( .C1(n18102), .C2(n20311), .A(n17189), .B(n17188), .ZN(
        n17190) );
  OAI211_X1 U20540 ( .C1(n17252), .C2(n17460), .A(n17191), .B(n17190), .ZN(
        P2_U3005) );
  XNOR2_X1 U20541 ( .A(n17192), .B(n17193), .ZN(n17473) );
  NAND2_X1 U20542 ( .A1(n17195), .A2(n17194), .ZN(n17198) );
  INV_X1 U20543 ( .A(n17209), .ZN(n17196) );
  AOI21_X1 U20544 ( .B1(n17211), .B2(n17208), .A(n17196), .ZN(n17197) );
  XOR2_X1 U20545 ( .A(n17198), .B(n17197), .Z(n17471) );
  NOR2_X1 U20546 ( .A1(n17461), .A2(n17242), .ZN(n17202) );
  NAND2_X1 U20547 ( .A1(n20343), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n17462) );
  NAND2_X1 U20548 ( .A1(n17214), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17199) );
  OAI211_X1 U20549 ( .C1(n17244), .C2(n17200), .A(n17462), .B(n17199), .ZN(
        n17201) );
  AOI211_X1 U20550 ( .C1(n17471), .C2(n18105), .A(n17202), .B(n17201), .ZN(
        n17203) );
  OAI21_X1 U20551 ( .B1(n17473), .B2(n17218), .A(n17203), .ZN(P2_U3006) );
  XNOR2_X1 U20552 ( .A(n17206), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17207) );
  XNOR2_X1 U20553 ( .A(n17205), .B(n17207), .ZN(n17486) );
  NAND2_X1 U20554 ( .A1(n17209), .A2(n17208), .ZN(n17210) );
  XNOR2_X1 U20555 ( .A(n17211), .B(n17210), .ZN(n17484) );
  NOR2_X1 U20556 ( .A1(n20260), .A2(n20990), .ZN(n17478) );
  NOR2_X1 U20557 ( .A1(n17244), .A2(n17212), .ZN(n17213) );
  AOI211_X1 U20558 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n17214), .A(
        n17478), .B(n17213), .ZN(n17215) );
  OAI21_X1 U20559 ( .B1(n17476), .B2(n17242), .A(n17215), .ZN(n17216) );
  AOI21_X1 U20560 ( .B1(n17484), .B2(n18105), .A(n17216), .ZN(n17217) );
  OAI21_X1 U20561 ( .B1(n17486), .B2(n17218), .A(n17217), .ZN(P2_U3007) );
  XNOR2_X1 U20562 ( .A(n17220), .B(n17219), .ZN(n17514) );
  INV_X1 U20563 ( .A(n17221), .ZN(n17226) );
  AOI21_X1 U20564 ( .B1(n17225), .B2(n17223), .A(n17222), .ZN(n17224) );
  AOI21_X1 U20565 ( .B1(n17226), .B2(n17225), .A(n17224), .ZN(n17501) );
  NAND2_X1 U20566 ( .A1(n17501), .A2(n18108), .ZN(n17230) );
  INV_X1 U20567 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n22021) );
  OAI22_X1 U20568 ( .A1(n22021), .A2(n18112), .B1(n17244), .B2(n20324), .ZN(
        n17228) );
  NOR2_X1 U20569 ( .A1(n17507), .A2(n17242), .ZN(n17227) );
  AOI211_X1 U20570 ( .C1(n20343), .C2(P2_REIP_REG_5__SCAN_IN), .A(n17228), .B(
        n17227), .ZN(n17229) );
  OAI211_X1 U20571 ( .C1(n17252), .C2(n17514), .A(n17230), .B(n17229), .ZN(
        P2_U3009) );
  XOR2_X1 U20572 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n17231), .Z(
        n17241) );
  AOI22_X1 U20573 ( .A1(n17241), .A2(n17240), .B1(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n17231), .ZN(n17233) );
  XNOR2_X1 U20574 ( .A(n20337), .B(n22037), .ZN(n17232) );
  XNOR2_X1 U20575 ( .A(n17233), .B(n17232), .ZN(n17523) );
  XNOR2_X1 U20576 ( .A(n17235), .B(n22037), .ZN(n17521) );
  INV_X1 U20577 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n20984) );
  OAI22_X1 U20578 ( .A1(n20340), .A2(n18112), .B1(n20984), .B2(n13139), .ZN(
        n17236) );
  AOI21_X1 U20579 ( .B1(n18102), .B2(n20354), .A(n17236), .ZN(n17237) );
  OAI21_X1 U20580 ( .B1(n17242), .B2(n20346), .A(n17237), .ZN(n17238) );
  AOI21_X1 U20581 ( .B1(n17521), .B2(n18108), .A(n17238), .ZN(n17239) );
  OAI21_X1 U20582 ( .B1(n17523), .B2(n17252), .A(n17239), .ZN(P2_U3010) );
  XNOR2_X1 U20583 ( .A(n17241), .B(n17240), .ZN(n17535) );
  NOR2_X1 U20584 ( .A1(n14288), .A2(n17242), .ZN(n17247) );
  INV_X1 U20585 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17245) );
  OAI22_X1 U20586 ( .A1(n17245), .A2(n18112), .B1(n17244), .B2(n17243), .ZN(
        n17246) );
  AOI211_X1 U20587 ( .C1(n20343), .C2(P2_REIP_REG_3__SCAN_IN), .A(n17247), .B(
        n17246), .ZN(n17251) );
  NAND3_X1 U20588 ( .A1(n17248), .A2(n17531), .A3(n18108), .ZN(n17250) );
  OAI211_X1 U20589 ( .C1(n17535), .C2(n17252), .A(n17251), .B(n17250), .ZN(
        P2_U3011) );
  NOR2_X1 U20590 ( .A1(n17253), .A2(n18123), .ZN(n17259) );
  OAI211_X1 U20591 ( .C1(n17257), .C2(n17256), .A(n17255), .B(n17254), .ZN(
        n17258) );
  AOI211_X1 U20592 ( .C1(n17260), .C2(n18120), .A(n17259), .B(n17258), .ZN(
        n17262) );
  NAND2_X1 U20593 ( .A1(n17264), .A2(n18120), .ZN(n17271) );
  AOI211_X1 U20594 ( .C1(n17267), .C2(n17266), .A(n17265), .B(n17278), .ZN(
        n17268) );
  AOI211_X1 U20595 ( .C1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n17282), .A(
        n17269), .B(n17268), .ZN(n17270) );
  OAI211_X1 U20596 ( .C1(n18123), .C2(n17272), .A(n17271), .B(n17270), .ZN(
        n17273) );
  AOI21_X1 U20597 ( .B1(n18126), .B2(n17274), .A(n17273), .ZN(n17275) );
  OAI21_X1 U20598 ( .B1(n17534), .B2(n17276), .A(n17275), .ZN(P2_U3020) );
  OAI21_X1 U20599 ( .B1(n17278), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17277), .ZN(n17281) );
  NOR2_X1 U20600 ( .A1(n17279), .A2(n18123), .ZN(n17280) );
  AOI211_X1 U20601 ( .C1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n17282), .A(
        n17281), .B(n17280), .ZN(n17283) );
  OAI21_X1 U20602 ( .B1(n17518), .B2(n17284), .A(n17283), .ZN(n17285) );
  INV_X1 U20603 ( .A(n17502), .ZN(n17425) );
  NOR2_X1 U20604 ( .A1(n17425), .A2(n10338), .ZN(n17289) );
  AOI21_X1 U20605 ( .B1(n17290), .B2(n17289), .A(n17288), .ZN(n17292) );
  OAI211_X1 U20606 ( .C1(n17293), .C2(n18123), .A(n17292), .B(n17291), .ZN(
        n17296) );
  NOR2_X1 U20607 ( .A1(n17294), .A2(n17518), .ZN(n17295) );
  OAI21_X1 U20608 ( .B1(n17299), .B2(n17534), .A(n17298), .ZN(P2_U3022) );
  NOR2_X1 U20609 ( .A1(n17300), .A2(n17534), .ZN(n17309) );
  NAND2_X1 U20610 ( .A1(n17302), .A2(n17301), .ZN(n17316) );
  XNOR2_X1 U20611 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17304) );
  OAI21_X1 U20612 ( .B1(n9785), .B2(n17304), .A(n17303), .ZN(n17305) );
  AOI21_X1 U20613 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17316), .A(
        n17305), .ZN(n17306) );
  OAI21_X1 U20614 ( .B1(n17307), .B2(n18123), .A(n17306), .ZN(n17308) );
  AOI211_X1 U20615 ( .C1(n17310), .C2(n18120), .A(n17309), .B(n17308), .ZN(
        n17311) );
  OAI21_X1 U20616 ( .B1(n17500), .B2(n17312), .A(n17311), .ZN(P2_U3023) );
  NOR2_X1 U20617 ( .A1(n9785), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17314) );
  AOI211_X1 U20618 ( .C1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n17316), .A(
        n17315), .B(n17314), .ZN(n17317) );
  OAI21_X1 U20619 ( .B1(n18123), .B2(n17318), .A(n17317), .ZN(n17319) );
  AOI21_X1 U20620 ( .B1(n17320), .B2(n18120), .A(n17319), .ZN(n17321) );
  OAI211_X1 U20621 ( .C1(n17323), .C2(n17534), .A(n17322), .B(n17321), .ZN(
        P2_U3024) );
  NAND2_X1 U20622 ( .A1(n17453), .A2(n17381), .ZN(n17324) );
  NAND2_X1 U20623 ( .A1(n17324), .A2(n17502), .ZN(n17379) );
  OR2_X1 U20624 ( .A1(n18129), .A2(n17325), .ZN(n17326) );
  NAND2_X1 U20625 ( .A1(n17379), .A2(n17326), .ZN(n17354) );
  AND2_X1 U20626 ( .A1(n17457), .A2(n17327), .ZN(n17341) );
  AND2_X1 U20627 ( .A1(n17341), .A2(n17328), .ZN(n17351) );
  OR2_X1 U20628 ( .A1(n17354), .A2(n17351), .ZN(n17345) );
  OAI21_X1 U20629 ( .B1(n17328), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17329) );
  OAI211_X1 U20630 ( .C1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n17341), .B(n17329), .ZN(
        n17330) );
  OAI211_X1 U20631 ( .C1(n17332), .C2(n18123), .A(n17331), .B(n17330), .ZN(
        n17333) );
  AOI21_X1 U20632 ( .B1(n17345), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n17333), .ZN(n17334) );
  OAI21_X1 U20633 ( .B1(n17335), .B2(n17518), .A(n17334), .ZN(n17336) );
  AOI21_X1 U20634 ( .B1(n17337), .B2(n18126), .A(n17336), .ZN(n17338) );
  OAI21_X1 U20635 ( .B1(n17339), .B2(n17534), .A(n17338), .ZN(P2_U3026) );
  NAND3_X1 U20636 ( .A1(n17341), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n17340), .ZN(n17343) );
  OAI211_X1 U20637 ( .C1(n18123), .C2(n20271), .A(n17343), .B(n17342), .ZN(
        n17344) );
  AOI21_X1 U20638 ( .B1(n17345), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n17344), .ZN(n17346) );
  OAI21_X1 U20639 ( .B1(n17347), .B2(n17518), .A(n17346), .ZN(n17348) );
  OAI21_X1 U20640 ( .B1(n17350), .B2(n17534), .A(n17349), .ZN(P2_U3027) );
  AOI211_X1 U20641 ( .C1(n17505), .C2(n17353), .A(n17352), .B(n17351), .ZN(
        n17356) );
  NAND2_X1 U20642 ( .A1(n17354), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17355) );
  OAI211_X1 U20643 ( .C1(n17357), .C2(n17518), .A(n17356), .B(n17355), .ZN(
        n17358) );
  AOI21_X1 U20644 ( .B1(n17359), .B2(n18126), .A(n17358), .ZN(n17360) );
  INV_X1 U20645 ( .A(n17379), .ZN(n17362) );
  INV_X1 U20646 ( .A(n17365), .ZN(n17366) );
  AOI21_X1 U20647 ( .B1(n17368), .B2(n17505), .A(n17367), .ZN(n17369) );
  AOI21_X1 U20648 ( .B1(n20364), .B2(n17505), .A(n17372), .ZN(n17373) );
  OAI21_X1 U20649 ( .B1(n17374), .B2(n17518), .A(n17373), .ZN(n17375) );
  NOR2_X1 U20650 ( .A1(n17379), .A2(n17380), .ZN(n17386) );
  NAND3_X1 U20651 ( .A1(n17457), .A2(n17381), .A3(n17380), .ZN(n17384) );
  AOI21_X1 U20652 ( .B1(n20285), .B2(n17505), .A(n17382), .ZN(n17383) );
  OAI211_X1 U20653 ( .C1(n20288), .C2(n17518), .A(n17384), .B(n17383), .ZN(
        n17385) );
  NAND2_X1 U20654 ( .A1(n17457), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17444) );
  NOR2_X1 U20655 ( .A1(n17444), .A2(n17388), .ZN(n17403) );
  NAND2_X1 U20656 ( .A1(n17403), .A2(n17418), .ZN(n17417) );
  INV_X1 U20657 ( .A(n17388), .ZN(n17430) );
  NAND3_X1 U20658 ( .A1(n17453), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        n17430), .ZN(n17389) );
  NAND2_X1 U20659 ( .A1(n17389), .A2(n17502), .ZN(n17419) );
  NAND2_X1 U20660 ( .A1(n17417), .A2(n17419), .ZN(n17408) );
  OAI21_X1 U20661 ( .B1(n17418), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17390) );
  OAI211_X1 U20662 ( .C1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(n17403), .B(n17390), .ZN(
        n17394) );
  AOI21_X1 U20663 ( .B1(n17392), .B2(n17505), .A(n17391), .ZN(n17393) );
  OAI211_X1 U20664 ( .C1(n17395), .C2(n17518), .A(n17394), .B(n17393), .ZN(
        n17396) );
  AOI21_X1 U20665 ( .B1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17408), .A(
        n17396), .ZN(n17399) );
  NAND2_X1 U20666 ( .A1(n17397), .A2(n18118), .ZN(n17398) );
  OAI211_X1 U20667 ( .C1(n17400), .C2(n17500), .A(n17399), .B(n17398), .ZN(
        P2_U3032) );
  NAND2_X1 U20668 ( .A1(n17401), .A2(n18126), .ZN(n17410) );
  NAND3_X1 U20669 ( .A1(n17403), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        n17402), .ZN(n17406) );
  AOI21_X1 U20670 ( .B1(n20304), .B2(n17505), .A(n17404), .ZN(n17405) );
  OAI211_X1 U20671 ( .C1(n20301), .C2(n17518), .A(n17406), .B(n17405), .ZN(
        n17407) );
  AOI21_X1 U20672 ( .B1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n17408), .A(
        n17407), .ZN(n17409) );
  OAI21_X1 U20673 ( .B1(n17413), .B2(n18123), .A(n17412), .ZN(n17414) );
  AOI21_X1 U20674 ( .B1(n17415), .B2(n18120), .A(n17414), .ZN(n17416) );
  OAI211_X1 U20675 ( .C1(n17419), .C2(n17418), .A(n17417), .B(n17416), .ZN(
        n17420) );
  AOI21_X1 U20676 ( .B1(n17421), .B2(n18118), .A(n17420), .ZN(n17422) );
  OAI21_X1 U20677 ( .B1(n17423), .B2(n17500), .A(n17422), .ZN(P2_U3034) );
  AOI21_X1 U20678 ( .B1(n17453), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n17425), .ZN(n17437) );
  AOI21_X1 U20679 ( .B1(n17427), .B2(n17505), .A(n17426), .ZN(n17428) );
  OAI21_X1 U20680 ( .B1(n17429), .B2(n17518), .A(n17428), .ZN(n17434) );
  AOI211_X1 U20681 ( .C1(n17432), .C2(n17431), .A(n17430), .B(n17444), .ZN(
        n17433) );
  AOI211_X1 U20682 ( .C1(n17437), .C2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n17434), .B(n17433), .ZN(n17435) );
  NAND2_X1 U20683 ( .A1(n17437), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17443) );
  NOR2_X1 U20684 ( .A1(n17438), .A2(n17518), .ZN(n17439) );
  AOI211_X1 U20685 ( .C1(n17505), .C2(n17441), .A(n17440), .B(n17439), .ZN(
        n17442) );
  OAI211_X1 U20686 ( .C1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n17444), .A(
        n17443), .B(n17442), .ZN(n17445) );
  AOI21_X1 U20687 ( .B1(n17446), .B2(n18118), .A(n17445), .ZN(n17447) );
  OAI21_X1 U20688 ( .B1(n17448), .B2(n17500), .A(n17447), .ZN(P2_U3036) );
  NAND3_X1 U20689 ( .A1(n17450), .A2(n18126), .A3(n17449), .ZN(n17459) );
  NAND2_X1 U20690 ( .A1(n20319), .A2(n17505), .ZN(n17451) );
  OAI211_X1 U20691 ( .C1(n20316), .C2(n17518), .A(n17452), .B(n17451), .ZN(
        n17455) );
  NOR2_X1 U20692 ( .A1(n17453), .A2(n17456), .ZN(n17454) );
  AOI211_X1 U20693 ( .C1(n17457), .C2(n17456), .A(n17455), .B(n17454), .ZN(
        n17458) );
  OAI211_X1 U20694 ( .C1(n17460), .C2(n17534), .A(n17459), .B(n17458), .ZN(
        P2_U3037) );
  INV_X1 U20695 ( .A(n17461), .ZN(n17467) );
  OAI21_X1 U20696 ( .B1(n17463), .B2(n18123), .A(n17462), .ZN(n17466) );
  XNOR2_X1 U20697 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17464) );
  NOR2_X1 U20698 ( .A1(n17481), .A2(n17464), .ZN(n17465) );
  AOI211_X1 U20699 ( .C1(n17467), .C2(n18120), .A(n17466), .B(n17465), .ZN(
        n17468) );
  OAI21_X1 U20700 ( .B1(n17475), .B2(n17469), .A(n17468), .ZN(n17470) );
  AOI21_X1 U20701 ( .B1(n17471), .B2(n18118), .A(n17470), .ZN(n17472) );
  OAI21_X1 U20702 ( .B1(n17473), .B2(n17500), .A(n17472), .ZN(P2_U3038) );
  NOR2_X1 U20703 ( .A1(n17475), .A2(n17474), .ZN(n17483) );
  NOR2_X1 U20704 ( .A1(n17476), .A2(n17518), .ZN(n17477) );
  AOI211_X1 U20705 ( .C1(n17505), .C2(n17479), .A(n17478), .B(n17477), .ZN(
        n17480) );
  OAI21_X1 U20706 ( .B1(n17481), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n17480), .ZN(n17482) );
  AOI211_X1 U20707 ( .C1(n17484), .C2(n18118), .A(n17483), .B(n17482), .ZN(
        n17485) );
  OAI21_X1 U20708 ( .B1(n17486), .B2(n17500), .A(n17485), .ZN(P2_U3039) );
  XNOR2_X1 U20709 ( .A(n17488), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n18103) );
  XOR2_X1 U20710 ( .A(n17490), .B(n17489), .Z(n18104) );
  NAND2_X1 U20711 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n20343), .ZN(n17491) );
  OAI211_X1 U20712 ( .C1(n17494), .C2(n17493), .A(n17492), .B(n17491), .ZN(
        n17498) );
  OAI22_X1 U20713 ( .A1(n17496), .A2(n17518), .B1(n18123), .B2(n17495), .ZN(
        n17497) );
  AOI211_X1 U20714 ( .C1(n18104), .C2(n18118), .A(n17498), .B(n17497), .ZN(
        n17499) );
  OAI21_X1 U20715 ( .B1(n18103), .B2(n17500), .A(n17499), .ZN(P2_U3040) );
  NAND2_X1 U20716 ( .A1(n17501), .A2(n18126), .ZN(n17513) );
  INV_X1 U20717 ( .A(n17525), .ZN(n17503) );
  NAND2_X1 U20718 ( .A1(n17503), .A2(n17502), .ZN(n17516) );
  INV_X1 U20719 ( .A(n17516), .ZN(n17511) );
  INV_X1 U20720 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n20986) );
  NOR2_X1 U20721 ( .A1(n20986), .A2(n13139), .ZN(n17504) );
  AOI21_X1 U20722 ( .B1(n20331), .B2(n17505), .A(n17504), .ZN(n17506) );
  OAI21_X1 U20723 ( .B1(n17507), .B2(n17518), .A(n17506), .ZN(n17510) );
  AOI211_X1 U20724 ( .C1(n22037), .C2(n12506), .A(n17508), .B(n17517), .ZN(
        n17509) );
  AOI211_X1 U20725 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n17511), .A(
        n17510), .B(n17509), .ZN(n17512) );
  OAI211_X1 U20726 ( .C1(n17514), .C2(n17534), .A(n17513), .B(n17512), .ZN(
        P2_U3041) );
  NAND2_X1 U20727 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n20343), .ZN(n17515) );
  OAI221_X1 U20728 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n17517), .C1(
        n22037), .C2(n17516), .A(n17515), .ZN(n17520) );
  OAI22_X1 U20729 ( .A1(n20346), .A2(n17518), .B1(n18123), .B2(n20369), .ZN(
        n17519) );
  AOI211_X1 U20730 ( .C1(n17521), .C2(n18126), .A(n17520), .B(n17519), .ZN(
        n17522) );
  OAI21_X1 U20731 ( .B1(n17523), .B2(n17534), .A(n17522), .ZN(P2_U3042) );
  OAI22_X1 U20732 ( .A1(n18123), .A2(n21051), .B1(n20983), .B2(n20260), .ZN(
        n17529) );
  INV_X1 U20733 ( .A(n17524), .ZN(n17527) );
  AOI21_X1 U20734 ( .B1(n17527), .B2(n17526), .A(n17525), .ZN(n17528) );
  AOI211_X1 U20735 ( .C1(n18120), .C2(n17530), .A(n17529), .B(n17528), .ZN(
        n17533) );
  NAND3_X1 U20736 ( .A1(n17248), .A2(n17531), .A3(n18126), .ZN(n17532) );
  OAI211_X1 U20737 ( .C1(n17535), .C2(n17534), .A(n17533), .B(n17532), .ZN(
        P2_U3043) );
  MUX2_X1 U20738 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n17536), .S(
        n20350), .Z(n17541) );
  OAI222_X1 U20739 ( .A1(n18136), .A2(n17539), .B1(n17538), .B2(n17541), .C1(
        n17553), .C2(n17537), .ZN(n17540) );
  MUX2_X1 U20740 ( .A(n17540), .B(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .S(
        n17555), .Z(P2_U3601) );
  NAND2_X1 U20741 ( .A1(n17541), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n17551) );
  INV_X1 U20742 ( .A(n17551), .ZN(n17544) );
  AOI21_X1 U20743 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n10160), .A(
        n17542), .ZN(n17550) );
  INV_X1 U20744 ( .A(n18136), .ZN(n17543) );
  AOI222_X1 U20745 ( .A1(n17546), .A2(n17545), .B1(n17544), .B2(n17550), .C1(
        n17543), .C2(n21072), .ZN(n17548) );
  NAND2_X1 U20746 ( .A1(n17555), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n17547) );
  OAI21_X1 U20747 ( .B1(n17548), .B2(n17555), .A(n17547), .ZN(P2_U3600) );
  OAI222_X1 U20748 ( .A1(n21058), .A2(n18136), .B1(n17551), .B2(n17550), .C1(
        n17553), .C2(n17549), .ZN(n17552) );
  MUX2_X1 U20749 ( .A(n17552), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n17555), .Z(P2_U3599) );
  OAI22_X1 U20750 ( .A1(n20713), .A2(n18136), .B1(n17554), .B2(n17553), .ZN(
        n17556) );
  MUX2_X1 U20751 ( .A(n17556), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n17555), .Z(P2_U3596) );
  OR2_X2 U20752 ( .A1(n21058), .A2(n21045), .ZN(n20650) );
  NOR2_X4 U20753 ( .A1(n20722), .A2(n20650), .ZN(n20954) );
  INV_X1 U20754 ( .A(n21042), .ZN(n20717) );
  NOR3_X1 U20755 ( .A1(n20954), .A2(n20486), .A3(n20717), .ZN(n17557) );
  NOR2_X1 U20756 ( .A1(n20717), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20680) );
  NOR2_X1 U20757 ( .A1(n17557), .A2(n20680), .ZN(n17561) );
  INV_X1 U20758 ( .A(n17558), .ZN(n17559) );
  AND2_X1 U20759 ( .A1(n17559), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20950) );
  NAND2_X1 U20760 ( .A1(n21054), .A2(n21065), .ZN(n20520) );
  NOR2_X1 U20761 ( .A1(n20678), .A2(n20520), .ZN(n20451) );
  NOR2_X1 U20762 ( .A1(n20950), .A2(n20451), .ZN(n17564) );
  INV_X1 U20763 ( .A(n12433), .ZN(n17562) );
  OAI21_X1 U20764 ( .B1(n17562), .B2(n20451), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n17560) );
  INV_X1 U20765 ( .A(n20455), .ZN(n17577) );
  INV_X1 U20766 ( .A(n9708), .ZN(n17572) );
  INV_X1 U20767 ( .A(n20904), .ZN(n17588) );
  INV_X1 U20768 ( .A(n20451), .ZN(n17571) );
  OAI22_X1 U20769 ( .A1(n20587), .A2(n17572), .B1(n17588), .B2(n17571), .ZN(
        n17568) );
  INV_X1 U20770 ( .A(n17561), .ZN(n17565) );
  AOI211_X1 U20771 ( .C1(n17562), .C2(n20834), .A(n21042), .B(n20451), .ZN(
        n17563) );
  NOR2_X1 U20772 ( .A1(n20459), .A2(n17566), .ZN(n17567) );
  AOI211_X1 U20773 ( .C1(n20954), .C2(n20906), .A(n17568), .B(n17567), .ZN(
        n17569) );
  OAI21_X1 U20774 ( .B1(n20725), .B2(n17577), .A(n17569), .ZN(P2_U3048) );
  NOR2_X2 U20775 ( .A1(n20394), .A2(n20623), .ZN(n20912) );
  INV_X1 U20776 ( .A(n20912), .ZN(n20728) );
  AOI22_X1 U20777 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20454), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n20453), .ZN(n20846) );
  INV_X1 U20778 ( .A(n20846), .ZN(n20913) );
  AOI22_X1 U20779 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n20454), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n20453), .ZN(n20590) );
  NAND2_X1 U20780 ( .A1(n13145), .A2(n17570), .ZN(n20469) );
  OAI22_X1 U20781 ( .A1(n20590), .A2(n17572), .B1(n17571), .B2(n20469), .ZN(
        n17575) );
  NOR2_X1 U20782 ( .A1(n20459), .A2(n17573), .ZN(n17574) );
  AOI211_X1 U20783 ( .C1(n20954), .C2(n20913), .A(n17575), .B(n17574), .ZN(
        n17576) );
  OAI21_X1 U20784 ( .B1(n17577), .B2(n20728), .A(n17576), .ZN(P2_U3049) );
  NOR2_X4 U20785 ( .A1(n20722), .A2(n21062), .ZN(n20886) );
  NOR2_X4 U20786 ( .A1(n20753), .A2(n20650), .ZN(n20953) );
  NOR3_X1 U20787 ( .A1(n20886), .A2(n20953), .A3(n20717), .ZN(n17578) );
  NOR2_X1 U20788 ( .A1(n17578), .A2(n20680), .ZN(n17581) );
  NOR3_X2 U20789 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21054), .A3(
        n20892), .ZN(n20885) );
  NOR2_X1 U20790 ( .A1(n21083), .A2(n20836), .ZN(n20862) );
  NOR2_X1 U20791 ( .A1(n20885), .A2(n20862), .ZN(n17584) );
  INV_X1 U20792 ( .A(n17579), .ZN(n17582) );
  OAI21_X1 U20793 ( .B1(n17582), .B2(n20885), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n17580) );
  INV_X1 U20794 ( .A(n20887), .ZN(n17594) );
  INV_X1 U20795 ( .A(n17581), .ZN(n17585) );
  AOI211_X1 U20796 ( .C1(n17582), .C2(n20834), .A(n21042), .B(n20885), .ZN(
        n17583) );
  INV_X1 U20797 ( .A(n20891), .ZN(n17592) );
  INV_X1 U20798 ( .A(n20886), .ZN(n17586) );
  NOR2_X1 U20799 ( .A1(n20843), .A2(n17586), .ZN(n17591) );
  INV_X1 U20800 ( .A(n20953), .ZN(n17589) );
  INV_X1 U20801 ( .A(n20885), .ZN(n17587) );
  OAI22_X1 U20802 ( .A1(n20587), .A2(n17589), .B1(n17588), .B2(n17587), .ZN(
        n17590) );
  AOI211_X1 U20803 ( .C1(n17592), .C2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n17591), .B(n17590), .ZN(n17593) );
  OAI21_X1 U20804 ( .B1(n20725), .B2(n17594), .A(n17593), .ZN(P2_U3160) );
  AOI21_X1 U20805 ( .B1(n17595), .B2(n17597), .A(n20237), .ZN(n17600) );
  NAND2_X1 U20806 ( .A1(n18135), .A2(n20959), .ZN(n18137) );
  INV_X1 U20807 ( .A(n18137), .ZN(n17598) );
  NOR3_X1 U20808 ( .A1(n17597), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n17596), 
        .ZN(n18132) );
  OAI21_X1 U20809 ( .B1(n17598), .B2(n18132), .A(P2_STATE2_REG_1__SCAN_IN), 
        .ZN(n17599) );
  OAI211_X1 U20810 ( .C1(n18135), .C2(n17600), .A(n17599), .B(n20351), .ZN(
        P2_U3177) );
  INV_X1 U20811 ( .A(n18598), .ZN(n20113) );
  AOI21_X1 U20812 ( .B1(n10451), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n18584), .ZN(n18520) );
  INV_X1 U20813 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n18484) );
  OAI21_X1 U20814 ( .B1(n18484), .B2(n18525), .A(n18593), .ZN(n17602) );
  INV_X1 U20815 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n18810) );
  NAND2_X1 U20816 ( .A1(n18815), .A2(n18810), .ZN(n18581) );
  OAI21_X1 U20817 ( .B1(n18810), .B2(n18815), .A(n18581), .ZN(n18811) );
  OAI22_X1 U20818 ( .A1(n18522), .A2(n18810), .B1(n18579), .B2(n18811), .ZN(
        n17601) );
  AOI221_X1 U20819 ( .B1(n18520), .B2(n19347), .C1(n17602), .C2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n17601), .ZN(n17604) );
  NOR2_X1 U20820 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n18568), .ZN(n18588) );
  AOI21_X1 U20821 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n18589), .A(n18588), .ZN(
        n17603) );
  OAI211_X1 U20822 ( .C1(n18565), .C2(n17605), .A(n17604), .B(n17603), .ZN(
        P3_U2670) );
  AOI21_X1 U20823 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n18808), .A(n17606), .ZN(
        n17623) );
  OAI22_X1 U20824 ( .A1(n18636), .A2(n17608), .B1(n17607), .B2(n18640), .ZN(
        n17609) );
  INV_X1 U20825 ( .A(n17609), .ZN(n17613) );
  AOI22_X1 U20826 ( .A1(n18760), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n18616), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17612) );
  AOI22_X1 U20827 ( .A1(n13659), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14112), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17611) );
  AOI22_X1 U20828 ( .A1(n10682), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n18717), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17610) );
  AND4_X1 U20829 ( .A1(n17613), .A2(n17612), .A3(n17611), .A4(n17610), .ZN(
        n17622) );
  OAI22_X1 U20830 ( .A1(n18790), .A2(n17985), .B1(n9704), .B2(n17614), .ZN(
        n17618) );
  OAI22_X1 U20831 ( .A1(n17616), .A2(n18755), .B1(n18754), .B2(n17615), .ZN(
        n17617) );
  NOR2_X1 U20832 ( .A1(n17618), .A2(n17617), .ZN(n17621) );
  AOI22_X1 U20833 ( .A1(n18743), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18742), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17620) );
  AOI22_X1 U20834 ( .A1(n14951), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18646), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17619) );
  AND4_X1 U20835 ( .A1(n17622), .A2(n17621), .A3(n17620), .A4(n17619), .ZN(
        n18865) );
  OAI22_X1 U20836 ( .A1(n17623), .A2(n9866), .B1(n18865), .B2(n18808), .ZN(
        P3_U2681) );
  OAI21_X1 U20837 ( .B1(n9871), .B2(P3_EBX_REG_20__SCAN_IN), .A(n18808), .ZN(
        n17648) );
  AOI22_X1 U20838 ( .A1(n9712), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n14457), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17639) );
  OAI22_X1 U20839 ( .A1(n17625), .A2(n18613), .B1(n17695), .B2(n17624), .ZN(
        n17629) );
  OAI22_X1 U20840 ( .A1(n18715), .A2(n17627), .B1(n17698), .B2(n17626), .ZN(
        n17628) );
  NOR2_X1 U20841 ( .A1(n17629), .A2(n17628), .ZN(n17638) );
  AOI22_X1 U20842 ( .A1(n9705), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18652), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17637) );
  NAND2_X1 U20843 ( .A1(n18760), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n17635) );
  NAND2_X1 U20844 ( .A1(n17630), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n17634) );
  NAND2_X1 U20845 ( .A1(n17631), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n17633) );
  NAND2_X1 U20846 ( .A1(n17693), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n17632) );
  AND4_X1 U20847 ( .A1(n17635), .A2(n17634), .A3(n17633), .A4(n17632), .ZN(
        n17636) );
  NAND4_X1 U20848 ( .A1(n17639), .A2(n17638), .A3(n17637), .A4(n17636), .ZN(
        n17647) );
  NAND2_X1 U20849 ( .A1(n14951), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n17645) );
  NAND2_X1 U20850 ( .A1(n18646), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n17644) );
  OR2_X1 U20851 ( .A1(n18775), .A2(n17640), .ZN(n17643) );
  OR2_X1 U20852 ( .A1(n18773), .A2(n17641), .ZN(n17642) );
  NAND4_X1 U20853 ( .A1(n17645), .A2(n17644), .A3(n17643), .A4(n17642), .ZN(
        n17646) );
  NOR2_X1 U20854 ( .A1(n17647), .A2(n17646), .ZN(n17713) );
  OAI22_X1 U20855 ( .A1(n17648), .A2(n18706), .B1(n17713), .B2(n18808), .ZN(
        P3_U2683) );
  OAI21_X1 U20856 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17684), .A(n17649), .ZN(
        n17666) );
  NOR2_X1 U20857 ( .A1(n18754), .A2(n13897), .ZN(n17652) );
  OAI22_X1 U20858 ( .A1(n17650), .A2(n9704), .B1(n17985), .B2(n11994), .ZN(
        n17651) );
  AOI211_X1 U20859 ( .C1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .C2(n9706), .A(
        n17652), .B(n17651), .ZN(n17661) );
  AOI22_X1 U20860 ( .A1(n18759), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12013), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17660) );
  AOI22_X1 U20861 ( .A1(n14099), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18616), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17659) );
  OAI22_X1 U20862 ( .A1(n18613), .A2(n17654), .B1(n17695), .B2(n17653), .ZN(
        n17657) );
  OAI22_X1 U20863 ( .A1(n18715), .A2(n17655), .B1(n17698), .B2(n13896), .ZN(
        n17656) );
  NOR2_X1 U20864 ( .A1(n17657), .A2(n17656), .ZN(n17658) );
  AND4_X1 U20865 ( .A1(n17661), .A2(n17660), .A3(n17659), .A4(n17658), .ZN(
        n17664) );
  AOI22_X1 U20866 ( .A1(n18743), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18742), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17663) );
  AOI22_X1 U20867 ( .A1(n14951), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n18646), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17662) );
  NAND3_X1 U20868 ( .A1(n17664), .A2(n17663), .A3(n17662), .ZN(n17718) );
  NAND2_X1 U20869 ( .A1(n18812), .A2(n17718), .ZN(n17665) );
  OAI21_X1 U20870 ( .B1(n17666), .B2(n18812), .A(n17665), .ZN(P3_U2684) );
  NOR2_X1 U20871 ( .A1(n17985), .A2(n18807), .ZN(n17669) );
  INV_X1 U20872 ( .A(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17667) );
  OAI22_X1 U20873 ( .A1(n18755), .A2(n17667), .B1(n18754), .B2(n18735), .ZN(
        n17668) );
  AOI211_X1 U20874 ( .C1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .C2(n9712), .A(
        n17669), .B(n17668), .ZN(n17677) );
  AOI22_X1 U20875 ( .A1(n18759), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12013), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17676) );
  AOI22_X1 U20876 ( .A1(n14099), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18616), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17675) );
  OAI22_X1 U20877 ( .A1(n18763), .A2(n18733), .B1(n14983), .B2(n17670), .ZN(
        n17673) );
  OAI22_X1 U20878 ( .A1(n18715), .A2(n17671), .B1(n17698), .B2(n18734), .ZN(
        n17672) );
  NOR2_X1 U20879 ( .A1(n17673), .A2(n17672), .ZN(n17674) );
  NAND4_X1 U20880 ( .A1(n17677), .A2(n17676), .A3(n17675), .A4(n17674), .ZN(
        n17683) );
  INV_X1 U20881 ( .A(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17679) );
  OAI22_X1 U20882 ( .A1(n18775), .A2(n17679), .B1(n18773), .B2(n17678), .ZN(
        n17682) );
  INV_X1 U20883 ( .A(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n21988) );
  OAI22_X1 U20884 ( .A1(n13862), .A2(n17680), .B1(n18777), .B2(n21988), .ZN(
        n17681) );
  NOR3_X1 U20885 ( .A1(n17683), .A2(n17682), .A3(n17681), .ZN(n17723) );
  INV_X1 U20886 ( .A(n17684), .ZN(n17685) );
  OAI211_X1 U20887 ( .C1(n17686), .C2(P3_EBX_REG_18__SCAN_IN), .A(n18808), .B(
        n17685), .ZN(n17687) );
  OAI21_X1 U20888 ( .B1(n17723), .B2(n18808), .A(n17687), .ZN(P3_U2685) );
  OAI21_X1 U20889 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n18727), .A(n17688), .ZN(
        n17710) );
  NOR2_X1 U20890 ( .A1(n17985), .A2(n18809), .ZN(n17692) );
  OAI22_X1 U20891 ( .A1(n17690), .A2(n18755), .B1(n18754), .B2(n17689), .ZN(
        n17691) );
  AOI211_X1 U20892 ( .C1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .C2(n9712), .A(
        n17692), .B(n17691), .ZN(n17705) );
  AOI22_X1 U20893 ( .A1(n18759), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17693), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17704) );
  AOI22_X1 U20894 ( .A1(n18760), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17631), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17703) );
  OAI22_X1 U20895 ( .A1(n18613), .A2(n17696), .B1(n17695), .B2(n17694), .ZN(
        n17701) );
  OAI22_X1 U20896 ( .A1(n18715), .A2(n17699), .B1(n18764), .B2(n17697), .ZN(
        n17700) );
  NOR2_X1 U20897 ( .A1(n17701), .A2(n17700), .ZN(n17702) );
  AND4_X1 U20898 ( .A1(n17705), .A2(n17704), .A3(n17703), .A4(n17702), .ZN(
        n17708) );
  AOI22_X1 U20899 ( .A1(n18743), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n18742), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17707) );
  AOI22_X1 U20900 ( .A1(n14951), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n18646), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17706) );
  NAND3_X1 U20901 ( .A1(n17708), .A2(n17707), .A3(n17706), .ZN(n17729) );
  NAND2_X1 U20902 ( .A1(n18812), .A2(n17729), .ZN(n17709) );
  OAI21_X1 U20903 ( .B1(n17710), .B2(n18812), .A(n17709), .ZN(P3_U2686) );
  INV_X1 U20904 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n18938) );
  INV_X1 U20905 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n18940) );
  NOR2_X1 U20906 ( .A1(n18938), .A2(n18940), .ZN(n18817) );
  INV_X1 U20907 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n19023) );
  INV_X1 U20908 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n19018) );
  INV_X1 U20909 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n18951) );
  NAND3_X1 U20910 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_13__SCAN_IN), 
        .A3(P3_EAX_REG_11__SCAN_IN), .ZN(n17734) );
  NOR3_X1 U20911 ( .A1(n19018), .A2(n18951), .A3(n17734), .ZN(n18885) );
  NAND2_X1 U20912 ( .A1(n17711), .A2(n18885), .ZN(n17735) );
  INV_X1 U20913 ( .A(n18879), .ZN(n17712) );
  NAND2_X1 U20914 ( .A1(n17712), .A2(n18606), .ZN(n18861) );
  AOI21_X1 U20915 ( .B1(n18902), .B2(P3_EAX_REG_20__SCAN_IN), .A(n17721), .ZN(
        n17717) );
  NAND2_X1 U20916 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17721), .ZN(n18876) );
  INV_X1 U20917 ( .A(n18876), .ZN(n17716) );
  NAND2_X1 U20918 ( .A1(n19646), .A2(n18907), .ZN(n18872) );
  OAI22_X1 U20919 ( .A1(n18883), .A2(n17713), .B1(n18872), .B2(n19641), .ZN(
        n17714) );
  AOI21_X1 U20920 ( .B1(BUF2_REG_20__SCAN_IN), .B2(n18877), .A(n17714), .ZN(
        n17715) );
  OAI21_X1 U20921 ( .B1(n17717), .B2(n17716), .A(n17715), .ZN(P3_U2715) );
  AOI21_X1 U20922 ( .B1(P3_EAX_REG_19__SCAN_IN), .B2(n18902), .A(n17727), .ZN(
        n17722) );
  AOI22_X1 U20923 ( .A1(n18911), .A2(n17718), .B1(BUF2_REG_3__SCAN_IN), .B2(
        n18878), .ZN(n17720) );
  NAND2_X1 U20924 ( .A1(n18877), .A2(BUF2_REG_19__SCAN_IN), .ZN(n17719) );
  OAI211_X1 U20925 ( .C1(n17722), .C2(n17721), .A(n17720), .B(n17719), .ZN(
        P3_U2716) );
  AND2_X1 U20926 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n17728), .ZN(n17732) );
  AOI21_X1 U20927 ( .B1(n18902), .B2(P3_EAX_REG_18__SCAN_IN), .A(n17732), .ZN(
        n17726) );
  OAI22_X1 U20928 ( .A1(n18883), .A2(n17723), .B1(n18872), .B2(n19633), .ZN(
        n17724) );
  AOI21_X1 U20929 ( .B1(BUF2_REG_18__SCAN_IN), .B2(n18877), .A(n17724), .ZN(
        n17725) );
  OAI21_X1 U20930 ( .B1(n17727), .B2(n17726), .A(n17725), .ZN(P3_U2717) );
  AOI21_X1 U20931 ( .B1(P3_EAX_REG_17__SCAN_IN), .B2(n18902), .A(n17728), .ZN(
        n17733) );
  AOI22_X1 U20932 ( .A1(n18911), .A2(n17729), .B1(BUF2_REG_1__SCAN_IN), .B2(
        n18878), .ZN(n17731) );
  NAND2_X1 U20933 ( .A1(n18877), .A2(BUF2_REG_17__SCAN_IN), .ZN(n17730) );
  OAI211_X1 U20934 ( .C1(n17733), .C2(n17732), .A(n17731), .B(n17730), .ZN(
        P3_U2718) );
  NOR2_X1 U20935 ( .A1(n17734), .A2(n18895), .ZN(n17737) );
  NAND2_X1 U20936 ( .A1(n18902), .A2(n17735), .ZN(n18888) );
  INV_X1 U20937 ( .A(n18888), .ZN(n17736) );
  MUX2_X1 U20938 ( .A(n17737), .B(n17736), .S(P3_EAX_REG_14__SCAN_IN), .Z(
        n17738) );
  AOI21_X1 U20939 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n18900), .A(n17738), .ZN(
        n17739) );
  OAI21_X1 U20940 ( .B1(n17740), .B2(n18883), .A(n17739), .ZN(P3_U2721) );
  INV_X1 U20941 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n19014) );
  INV_X1 U20942 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n18949) );
  AOI21_X1 U20943 ( .B1(n18902), .B2(P3_EAX_REG_12__SCAN_IN), .A(n17746), .ZN(
        n17742) );
  NAND2_X1 U20944 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17746), .ZN(n18893) );
  INV_X1 U20945 ( .A(n18893), .ZN(n17741) );
  OAI222_X1 U20946 ( .A1(n18913), .A2(n19014), .B1(n18883), .B2(n17743), .C1(
        n17742), .C2(n17741), .ZN(P3_U2723) );
  INV_X1 U20947 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n19011) );
  INV_X1 U20948 ( .A(n17744), .ZN(n17748) );
  INV_X1 U20949 ( .A(n18895), .ZN(n17745) );
  AOI21_X1 U20950 ( .B1(n18902), .B2(P3_EAX_REG_11__SCAN_IN), .A(n17745), .ZN(
        n17747) );
  OAI222_X1 U20951 ( .A1(n18913), .A2(n19011), .B1(n18883), .B2(n17748), .C1(
        n17747), .C2(n17746), .ZN(P3_U2724) );
  INV_X1 U20952 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n21919) );
  INV_X1 U20953 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n18958) );
  NOR2_X1 U20954 ( .A1(n18958), .A2(n17749), .ZN(n17753) );
  AOI21_X1 U20955 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n18902), .A(n17753), .ZN(
        n17751) );
  OAI222_X1 U20956 ( .A1(n18883), .A2(n17778), .B1(n18913), .B2(n21919), .C1(
        n17751), .C2(n17750), .ZN(P3_U2728) );
  INV_X1 U20957 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n19649) );
  AOI21_X1 U20958 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n18902), .A(n17752), .ZN(
        n17754) );
  OAI222_X1 U20959 ( .A1(n18883), .A2(n17755), .B1(n18913), .B2(n19649), .C1(
        n17754), .C2(n17753), .ZN(P3_U2729) );
  NAND2_X1 U20960 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17964) );
  INV_X1 U20961 ( .A(n17964), .ZN(n17858) );
  NAND2_X1 U20962 ( .A1(n17858), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n19518) );
  NOR2_X1 U20963 ( .A1(n19518), .A2(n19524), .ZN(n19514) );
  NAND2_X1 U20964 ( .A1(n19514), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n19498) );
  AND2_X1 U20965 ( .A1(n19198), .A2(n17891), .ZN(n17756) );
  NOR2_X1 U20966 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n19259) );
  INV_X1 U20967 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17862) );
  NAND2_X1 U20968 ( .A1(n19259), .A2(n17862), .ZN(n19197) );
  INV_X1 U20969 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n19502) );
  INV_X1 U20970 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17843) );
  NAND4_X1 U20971 ( .A1(n19502), .A2(n17843), .A3(n19230), .A4(n19524), .ZN(
        n17757) );
  NAND2_X1 U20972 ( .A1(n19196), .A2(n17757), .ZN(n17758) );
  NAND2_X1 U20973 ( .A1(n19222), .A2(n17758), .ZN(n17760) );
  INV_X1 U20974 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n19464) );
  AND2_X1 U20975 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n19455) );
  NAND2_X1 U20976 ( .A1(n19175), .A2(n19455), .ZN(n19100) );
  INV_X1 U20977 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n21966) );
  INV_X1 U20978 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n19159) );
  NAND2_X1 U20979 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n19426) );
  NOR3_X1 U20980 ( .A1(n21966), .A2(n19159), .A3(n19426), .ZN(n19102) );
  AND2_X1 U20981 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n19102), .ZN(
        n19079) );
  AND2_X1 U20982 ( .A1(n19079), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17762) );
  AND2_X1 U20983 ( .A1(n17762), .A2(n19455), .ZN(n19073) );
  NAND2_X1 U20984 ( .A1(n19196), .A2(n19159), .ZN(n19158) );
  NOR2_X1 U20985 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n19158), .ZN(
        n19133) );
  INV_X1 U20986 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n19136) );
  NAND2_X1 U20987 ( .A1(n19133), .A2(n19136), .ZN(n19110) );
  NOR2_X1 U20988 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n19110), .ZN(
        n19101) );
  INV_X1 U20989 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n19394) );
  INV_X1 U20990 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n19419) );
  NAND3_X1 U20991 ( .A1(n19101), .A2(n19394), .A3(n19419), .ZN(n17763) );
  INV_X1 U20992 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n22049) );
  AND2_X1 U20993 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17901) );
  NAND2_X1 U20994 ( .A1(n17765), .A2(n10323), .ZN(n19060) );
  OAI21_X1 U20995 ( .B1(n17901), .B2(n19196), .A(n19060), .ZN(n17766) );
  AND2_X1 U20996 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17928) );
  AND2_X1 U20997 ( .A1(n17928), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17895) );
  INV_X1 U20998 ( .A(n17895), .ZN(n17903) );
  OAI21_X1 U20999 ( .B1(n17770), .B2(n19196), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n17769) );
  XNOR2_X1 U21000 ( .A(n19196), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n17772) );
  INV_X1 U21001 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n19034) );
  INV_X1 U21002 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17939) );
  NAND2_X1 U21003 ( .A1(n19196), .A2(n17939), .ZN(n17768) );
  INV_X1 U21004 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17932) );
  NAND2_X1 U21005 ( .A1(n17808), .A2(n17932), .ZN(n17794) );
  NAND2_X1 U21006 ( .A1(n17794), .A2(n19196), .ZN(n17771) );
  NAND3_X1 U21007 ( .A1(n17769), .A2(n17772), .A3(n17771), .ZN(n17777) );
  INV_X1 U21008 ( .A(n17770), .ZN(n17795) );
  NAND2_X1 U21009 ( .A1(n17775), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17902) );
  NAND3_X1 U21010 ( .A1(n17771), .A2(n17795), .A3(n17902), .ZN(n17774) );
  INV_X1 U21011 ( .A(n17772), .ZN(n17773) );
  OAI211_X1 U21012 ( .C1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n17775), .A(
        n17774), .B(n17773), .ZN(n17776) );
  NAND2_X1 U21013 ( .A1(n17777), .A2(n17776), .ZN(n17912) );
  INV_X1 U21014 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n19078) );
  INV_X1 U21015 ( .A(n19355), .ZN(n17913) );
  NAND2_X1 U21016 ( .A1(n17913), .A2(n17895), .ZN(n17919) );
  INV_X1 U21017 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n17779) );
  OAI21_X1 U21018 ( .B1(n17919), .B2(n17779), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n17780) );
  OAI21_X1 U21019 ( .B1(n17902), .B2(n17919), .A(n17780), .ZN(n17910) );
  INV_X2 U21020 ( .A(n19334), .ZN(n19340) );
  INV_X1 U21021 ( .A(n17891), .ZN(n19174) );
  NOR2_X1 U21022 ( .A1(n19403), .A2(n10016), .ZN(n19386) );
  INV_X1 U21023 ( .A(n19386), .ZN(n19064) );
  NOR2_X1 U21024 ( .A1(n19064), .A2(n19078), .ZN(n19049) );
  AND2_X1 U21025 ( .A1(n19049), .A2(n17901), .ZN(n19357) );
  INV_X1 U21026 ( .A(n19357), .ZN(n17916) );
  NOR2_X1 U21027 ( .A1(n17916), .A2(n17903), .ZN(n17921) );
  NAND2_X1 U21028 ( .A1(n17921), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17781) );
  XOR2_X1 U21029 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n17781), .Z(
        n17908) );
  NOR2_X1 U21030 ( .A1(n17908), .A2(n19208), .ZN(n17792) );
  INV_X1 U21031 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n19038) );
  NAND3_X1 U21032 ( .A1(n17782), .A2(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n19039) );
  NOR2_X1 U21033 ( .A1(n19038), .A2(n19039), .ZN(n17828) );
  NAND3_X1 U21034 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A3(n17828), .ZN(n17814) );
  NOR2_X1 U21035 ( .A1(n18263), .A2(n17814), .ZN(n17783) );
  NOR2_X1 U21036 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n20220) );
  NAND3_X1 U21037 ( .A1(n20107), .A2(n21986), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n19911) );
  NAND2_X1 U21038 ( .A1(n17783), .A2(n19212), .ZN(n17805) );
  XNOR2_X1 U21039 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n17790) );
  NOR2_X1 U21040 ( .A1(n18914), .A2(n20216), .ZN(n19307) );
  NOR2_X2 U21041 ( .A1(n19306), .A2(n19307), .ZN(n19348) );
  NOR2_X1 U21042 ( .A1(n19603), .A2(n20186), .ZN(n17905) );
  NOR2_X1 U21043 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n19082), .ZN(
        n17813) );
  INV_X1 U21044 ( .A(n19214), .ZN(n19142) );
  INV_X1 U21045 ( .A(n17783), .ZN(n17784) );
  AOI22_X1 U21046 ( .A1(n19142), .A2(n17785), .B1(n20002), .B2(n17784), .ZN(
        n17786) );
  NAND2_X1 U21047 ( .A1(n17786), .A2(n19313), .ZN(n17815) );
  NOR2_X1 U21048 ( .A1(n17813), .A2(n17815), .ZN(n17799) );
  NOR2_X1 U21049 ( .A1(n17787), .A2(n17799), .ZN(n17788) );
  AOI211_X1 U21050 ( .C1(n19236), .C2(n10451), .A(n17905), .B(n17788), .ZN(
        n17789) );
  OAI21_X1 U21051 ( .B1(n17805), .B2(n17790), .A(n17789), .ZN(n17791) );
  AOI211_X1 U21052 ( .C1(n17910), .C2(n19340), .A(n17792), .B(n17791), .ZN(
        n17793) );
  OAI21_X1 U21053 ( .B1(n17912), .B2(n19204), .A(n17793), .ZN(P3_U2799) );
  NAND2_X1 U21054 ( .A1(n17795), .A2(n17794), .ZN(n17796) );
  XNOR2_X1 U21055 ( .A(n17796), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17925) );
  OAI22_X1 U21056 ( .A1(n10312), .A2(n19334), .B1(n17921), .B2(n19208), .ZN(
        n17822) );
  NAND2_X1 U21057 ( .A1(n19455), .A2(n19102), .ZN(n19413) );
  NAND2_X1 U21058 ( .A1(n19188), .A2(n19340), .ZN(n17798) );
  INV_X2 U21059 ( .A(n19208), .ZN(n19065) );
  NAND2_X1 U21060 ( .A1(n19065), .A2(n19209), .ZN(n17797) );
  NOR2_X1 U21061 ( .A1(n19413), .A2(n19187), .ZN(n19106) );
  NAND2_X1 U21062 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n19106), .ZN(
        n19091) );
  NOR2_X1 U21063 ( .A1(n19394), .A2(n19078), .ZN(n19037) );
  NAND2_X1 U21064 ( .A1(n17901), .A2(n19037), .ZN(n19349) );
  NOR2_X1 U21065 ( .A1(n19091), .A2(n19349), .ZN(n19035) );
  NOR2_X1 U21066 ( .A1(n17903), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17918) );
  NAND2_X1 U21067 ( .A1(n19035), .A2(n17918), .ZN(n17804) );
  AND2_X1 U21068 ( .A1(n19566), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n17917) );
  NOR2_X1 U21069 ( .A1(n17800), .A2(n17799), .ZN(n17801) );
  AOI211_X1 U21070 ( .C1(n19236), .C2(n17802), .A(n17917), .B(n17801), .ZN(
        n17803) );
  OAI211_X1 U21071 ( .C1(n17805), .C2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n17804), .B(n17803), .ZN(n17806) );
  AOI21_X1 U21072 ( .B1(n17822), .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n17806), .ZN(n17807) );
  OAI21_X1 U21073 ( .B1(n17925), .B2(n19204), .A(n17807), .ZN(P3_U2800) );
  INV_X1 U21074 ( .A(n19027), .ZN(n17809) );
  AOI21_X1 U21075 ( .B1(n17809), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n17808), .ZN(n17810) );
  XNOR2_X1 U21076 ( .A(n17810), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17934) );
  INV_X1 U21077 ( .A(n17934), .ZN(n17824) );
  INV_X1 U21078 ( .A(n17921), .ZN(n17812) );
  INV_X1 U21079 ( .A(n17928), .ZN(n17811) );
  NOR2_X1 U21080 ( .A1(n17916), .A2(n17811), .ZN(n17951) );
  NAND3_X1 U21081 ( .A1(n17812), .A2(n19065), .A3(n17951), .ZN(n17819) );
  NAND2_X1 U21082 ( .A1(n19566), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n17931) );
  OAI21_X1 U21083 ( .B1(n19236), .B2(n17813), .A(n18261), .ZN(n17818) );
  NOR2_X1 U21084 ( .A1(n17814), .A2(n19863), .ZN(n17816) );
  OAI21_X1 U21085 ( .B1(n17816), .B2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n17815), .ZN(n17817) );
  NAND4_X1 U21086 ( .A1(n17819), .A2(n17931), .A3(n17818), .A4(n17817), .ZN(
        n17821) );
  NAND2_X1 U21087 ( .A1(n17913), .A2(n17928), .ZN(n17945) );
  NOR3_X1 U21088 ( .A1(n10312), .A2(n19334), .A3(n17945), .ZN(n17820) );
  AOI211_X1 U21089 ( .C1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n17822), .A(
        n17821), .B(n17820), .ZN(n17823) );
  OAI21_X1 U21090 ( .B1(n17824), .B2(n19204), .A(n17823), .ZN(P3_U2801) );
  XNOR2_X1 U21091 ( .A(n19196), .B(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n17954) );
  XNOR2_X1 U21092 ( .A(n17944), .B(n17954), .ZN(n17838) );
  NOR2_X1 U21093 ( .A1(n19340), .A2(n19065), .ZN(n19130) );
  OAI22_X1 U21094 ( .A1(n17913), .A2(n19334), .B1(n19357), .B2(n19208), .ZN(
        n19046) );
  NOR2_X1 U21095 ( .A1(n19034), .A2(n19046), .ZN(n17825) );
  NOR3_X1 U21096 ( .A1(n19130), .A2(n17825), .A3(n17939), .ZN(n17836) );
  OR2_X1 U21097 ( .A1(n19034), .A2(n19349), .ZN(n17938) );
  OR2_X1 U21098 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17938), .ZN(
        n17826) );
  NOR2_X1 U21099 ( .A1(n19091), .A2(n17826), .ZN(n17835) );
  INV_X1 U21100 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17830) );
  NAND2_X1 U21101 ( .A1(n17828), .A2(n19212), .ZN(n19032) );
  AOI221_X1 U21102 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C1(n19031), .C2(n17830), .A(
        n19032), .ZN(n17834) );
  INV_X1 U21103 ( .A(n19307), .ZN(n19140) );
  OR2_X1 U21104 ( .A1(n19214), .A2(n11873), .ZN(n17827) );
  OAI211_X1 U21105 ( .C1(n17828), .C2(n19140), .A(n19313), .B(n17827), .ZN(
        n19044) );
  AOI21_X1 U21106 ( .B1(n19123), .B2(n19038), .A(n19044), .ZN(n19030) );
  OAI22_X1 U21107 ( .A1(n19030), .A2(n17830), .B1(n19183), .B2(n17829), .ZN(
        n17832) );
  NAND2_X1 U21108 ( .A1(n19566), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17959) );
  INV_X1 U21109 ( .A(n17959), .ZN(n17831) );
  OR2_X1 U21110 ( .A1(n17832), .A2(n17831), .ZN(n17833) );
  NOR4_X1 U21111 ( .A1(n17836), .A2(n17835), .A3(n17834), .A4(n17833), .ZN(
        n17837) );
  OAI21_X1 U21112 ( .B1(n17838), .B2(n19204), .A(n17837), .ZN(P3_U2802) );
  AND2_X1 U21113 ( .A1(n11883), .A2(n19212), .ZN(n19179) );
  INV_X1 U21114 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18418) );
  INV_X1 U21115 ( .A(n11883), .ZN(n17839) );
  INV_X1 U21116 ( .A(n19348), .ZN(n17869) );
  OAI21_X1 U21117 ( .B1(n19306), .B2(n17839), .A(n17869), .ZN(n19193) );
  OAI21_X1 U21118 ( .B1(n17840), .B2(n19214), .A(n19193), .ZN(n19177) );
  OAI22_X1 U21119 ( .A1(n18418), .A2(n17840), .B1(n18428), .B2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18407) );
  INV_X1 U21120 ( .A(n18407), .ZN(n18405) );
  OAI22_X1 U21121 ( .A1(n19613), .A2(n20159), .B1(n19183), .B2(n18405), .ZN(
        n17841) );
  AOI221_X1 U21122 ( .B1(n19179), .B2(n18418), .C1(n19177), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17841), .ZN(n17853) );
  NAND2_X1 U21123 ( .A1(n19189), .A2(n17843), .ZN(n19490) );
  NOR2_X1 U21124 ( .A1(n19405), .A2(n19334), .ZN(n17851) );
  NAND2_X1 U21125 ( .A1(n19065), .A2(n19403), .ZN(n19092) );
  INV_X1 U21126 ( .A(n19476), .ZN(n17842) );
  OR2_X1 U21127 ( .A1(n17856), .A2(n17842), .ZN(n19202) );
  AND2_X1 U21128 ( .A1(n19202), .A2(n17843), .ZN(n19487) );
  NOR2_X1 U21129 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n19524), .ZN(
        n19520) );
  NOR2_X1 U21130 ( .A1(n17977), .A2(n19197), .ZN(n19237) );
  INV_X1 U21131 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n19230) );
  NAND2_X1 U21132 ( .A1(n19502), .A2(n19230), .ZN(n19190) );
  INV_X1 U21133 ( .A(n19190), .ZN(n17846) );
  NAND3_X1 U21134 ( .A1(n17844), .A2(n19514), .A3(n19198), .ZN(n19225) );
  NOR3_X1 U21135 ( .A1(n19196), .A2(n19502), .A3(n19225), .ZN(n17845) );
  AOI21_X1 U21136 ( .B1(n19237), .B2(n17846), .A(n17845), .ZN(n17847) );
  NOR2_X1 U21137 ( .A1(n19520), .A2(n17847), .ZN(n17848) );
  XOR2_X1 U21138 ( .A(n17848), .B(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .Z(
        n19488) );
  INV_X1 U21139 ( .A(n19488), .ZN(n17849) );
  OAI22_X1 U21140 ( .A1(n19092), .A2(n19487), .B1(n19204), .B2(n17849), .ZN(
        n17850) );
  AOI21_X1 U21141 ( .B1(n19490), .B2(n17851), .A(n17850), .ZN(n17852) );
  NAND2_X1 U21142 ( .A1(n17853), .A2(n17852), .ZN(P3_U2815) );
  INV_X1 U21143 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n19251) );
  INV_X1 U21144 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n21933) );
  NOR3_X1 U21145 ( .A1(n22115), .A2(n11890), .A3(n19863), .ZN(n19261) );
  NAND2_X1 U21146 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n19261), .ZN(
        n17882) );
  NOR2_X1 U21147 ( .A1(n21933), .A2(n17882), .ZN(n17868) );
  NAND2_X1 U21148 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17868), .ZN(
        n19252) );
  NOR2_X1 U21149 ( .A1(n19251), .A2(n19252), .ZN(n19250) );
  AOI21_X1 U21150 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17869), .A(
        n19250), .ZN(n17855) );
  INV_X1 U21151 ( .A(n17854), .ZN(n19217) );
  NOR2_X1 U21152 ( .A1(n19217), .A2(n19863), .ZN(n19192) );
  NOR2_X1 U21153 ( .A1(n17880), .A2(n18519), .ZN(n18483) );
  NAND2_X1 U21154 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n18483), .ZN(
        n18467) );
  NOR2_X1 U21155 ( .A1(n19251), .A2(n18467), .ZN(n18466) );
  NAND2_X1 U21156 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17854), .ZN(
        n18449) );
  OAI21_X1 U21157 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n18466), .A(
        n18449), .ZN(n18456) );
  OAI22_X1 U21158 ( .A1(n17855), .A2(n19192), .B1(n19309), .B2(n18456), .ZN(
        n17867) );
  AOI22_X1 U21159 ( .A1(n17857), .A2(n19340), .B1(n19065), .B2(n17856), .ZN(
        n19245) );
  NAND2_X1 U21160 ( .A1(n17873), .A2(n17964), .ZN(n19246) );
  AOI21_X1 U21161 ( .B1(n19245), .B2(n19246), .A(n17862), .ZN(n17866) );
  INV_X1 U21162 ( .A(n17873), .ZN(n19227) );
  NAND2_X1 U21163 ( .A1(n17858), .A2(n17862), .ZN(n17971) );
  INV_X1 U21164 ( .A(n19200), .ZN(n19239) );
  NOR2_X1 U21165 ( .A1(n19239), .A2(n17964), .ZN(n17979) );
  INV_X1 U21166 ( .A(n19259), .ZN(n17859) );
  NOR2_X1 U21167 ( .A1(n17977), .A2(n17859), .ZN(n17860) );
  NOR2_X1 U21168 ( .A1(n17979), .A2(n17860), .ZN(n17861) );
  XOR2_X1 U21169 ( .A(n17862), .B(n17861), .Z(n17968) );
  NOR2_X1 U21170 ( .A1(n19603), .A2(n20151), .ZN(n17863) );
  AOI21_X1 U21171 ( .B1(n19254), .B2(n17968), .A(n17863), .ZN(n17864) );
  OAI21_X1 U21172 ( .B1(n19227), .B2(n17971), .A(n17864), .ZN(n17865) );
  OR3_X1 U21173 ( .A1(n17867), .A2(n17866), .A3(n17865), .ZN(P3_U2819) );
  INV_X1 U21174 ( .A(n19252), .ZN(n17871) );
  AOI21_X1 U21175 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17869), .A(
        n17868), .ZN(n17870) );
  OAI21_X1 U21176 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18483), .A(
        n18467), .ZN(n18487) );
  OAI22_X1 U21177 ( .A1(n17871), .A2(n17870), .B1(n19309), .B2(n18487), .ZN(
        n17872) );
  AOI21_X1 U21178 ( .B1(n17974), .B2(n17873), .A(n17872), .ZN(n17877) );
  NOR2_X1 U21179 ( .A1(n19613), .A2(n14407), .ZN(n17874) );
  AOI21_X1 U21180 ( .B1(n19254), .B2(n17875), .A(n17874), .ZN(n17876) );
  OAI211_X1 U21181 ( .C1(n17974), .C2(n19245), .A(n17877), .B(n17876), .ZN(
        P3_U2821) );
  NOR2_X1 U21182 ( .A1(n19208), .A2(n17878), .ZN(n17885) );
  OAI21_X1 U21183 ( .B1(n17879), .B2(n19140), .A(n19313), .ZN(n19262) );
  AOI21_X1 U21184 ( .B1(n20002), .B2(n17880), .A(n19262), .ZN(n17883) );
  OAI221_X1 U21185 ( .B1(n17883), .B2(n21933), .C1(n17883), .C2(n17882), .A(
        n17881), .ZN(n17884) );
  AOI211_X1 U21186 ( .C1(n19254), .C2(n17886), .A(n17885), .B(n17884), .ZN(
        n17888) );
  INV_X1 U21187 ( .A(n18519), .ZN(n18507) );
  NAND2_X1 U21188 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n18507), .ZN(
        n18506) );
  AOI21_X1 U21189 ( .B1(n21933), .B2(n18506), .A(n18483), .ZN(n18496) );
  NAND2_X1 U21190 ( .A1(n19344), .A2(n18496), .ZN(n17887) );
  OAI211_X1 U21191 ( .C1(n17889), .C2(n19334), .A(n17888), .B(n17887), .ZN(
        P3_U2822) );
  INV_X1 U21192 ( .A(n19497), .ZN(n19565) );
  INV_X1 U21193 ( .A(n19455), .ZN(n19116) );
  NAND2_X1 U21194 ( .A1(n17891), .A2(n17890), .ZN(n17936) );
  NOR2_X1 U21195 ( .A1(n19116), .A2(n17936), .ZN(n19454) );
  NAND2_X1 U21196 ( .A1(n19079), .A2(n19454), .ZN(n19387) );
  INV_X1 U21197 ( .A(n19037), .ZN(n19352) );
  OR2_X1 U21198 ( .A1(n19387), .A2(n19352), .ZN(n17899) );
  INV_X1 U21199 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n19050) );
  AOI21_X1 U21200 ( .B1(n17899), .B2(n20058), .A(n19050), .ZN(n19372) );
  AND2_X1 U21201 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n19372), .ZN(
        n19353) );
  NAND2_X1 U21202 ( .A1(n17891), .A2(n19495), .ZN(n19474) );
  NOR2_X1 U21203 ( .A1(n19474), .A2(n19413), .ZN(n19351) );
  NAND2_X1 U21204 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n19351), .ZN(
        n17892) );
  OAI21_X1 U21205 ( .B1(n17892), .B2(n19349), .A(n19604), .ZN(n17894) );
  INV_X1 U21206 ( .A(n17892), .ZN(n17897) );
  NAND2_X1 U21207 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17897), .ZN(
        n19350) );
  OAI21_X1 U21208 ( .B1(n19350), .B2(n17938), .A(n19526), .ZN(n17893) );
  OAI211_X1 U21209 ( .C1(n19353), .C2(n19560), .A(n17894), .B(n17893), .ZN(
        n17948) );
  NAND2_X1 U21210 ( .A1(n17948), .A2(n19598), .ZN(n17920) );
  OAI21_X1 U21211 ( .B1(n17895), .B2(n19565), .A(n19564), .ZN(n17922) );
  INV_X1 U21212 ( .A(n17922), .ZN(n17896) );
  OAI211_X1 U21213 ( .C1(n19565), .C2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n17920), .B(n17896), .ZN(n17906) );
  NAND3_X1 U21214 ( .A1(n19037), .A2(n17897), .A3(n19593), .ZN(n17898) );
  OAI21_X1 U21215 ( .B1(n17899), .B2(n19560), .A(n17898), .ZN(n17900) );
  AND2_X1 U21216 ( .A1(n17900), .A2(n19598), .ZN(n19370) );
  NAND2_X1 U21217 ( .A1(n19370), .A2(n17901), .ZN(n17914) );
  NOR3_X1 U21218 ( .A1(n17914), .A2(n17903), .A3(n17902), .ZN(n17904) );
  AOI211_X1 U21219 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n17906), .A(
        n17905), .B(n17904), .ZN(n17907) );
  OAI21_X1 U21220 ( .B1(n17908), .B2(n19504), .A(n17907), .ZN(n17909) );
  AOI21_X1 U21221 ( .B1(n17910), .B2(n19610), .A(n17909), .ZN(n17911) );
  OAI21_X1 U21222 ( .B1(n17912), .B2(n19505), .A(n17911), .ZN(P3_U2831) );
  NAND2_X1 U21223 ( .A1(n17913), .A2(n19610), .ZN(n17915) );
  OAI211_X1 U21224 ( .C1(n19504), .C2(n17916), .A(n17915), .B(n17914), .ZN(
        n17929) );
  AOI21_X1 U21225 ( .B1(n17929), .B2(n17918), .A(n17917), .ZN(n17924) );
  OAI21_X1 U21226 ( .B1(n17926), .B2(n17922), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n17923) );
  OAI211_X1 U21227 ( .C1(n17925), .C2(n19505), .A(n17924), .B(n17923), .ZN(
        P3_U2832) );
  NOR2_X1 U21228 ( .A1(n19604), .A2(n20058), .ZN(n19516) );
  INV_X1 U21229 ( .A(n19516), .ZN(n17965) );
  NAND2_X1 U21230 ( .A1(n19034), .A2(n17965), .ZN(n17946) );
  OAI21_X1 U21231 ( .B1(n19575), .B2(n17946), .A(n19564), .ZN(n17927) );
  NAND3_X1 U21232 ( .A1(n17929), .A2(n17928), .A3(n17932), .ZN(n17930) );
  AOI21_X1 U21233 ( .B1(n19530), .B2(n17934), .A(n17933), .ZN(n17935) );
  INV_X1 U21234 ( .A(n17935), .ZN(P3_U2833) );
  INV_X1 U21235 ( .A(n19474), .ZN(n19453) );
  NOR2_X1 U21236 ( .A1(n19560), .A2(n17936), .ZN(n17937) );
  INV_X1 U21237 ( .A(n19405), .ZN(n19491) );
  INV_X1 U21238 ( .A(n20057), .ZN(n19404) );
  OAI22_X1 U21239 ( .A1(n19491), .A2(n19404), .B1(n19403), .B2(n19401), .ZN(
        n19451) );
  NOR2_X1 U21240 ( .A1(n19414), .A2(n19116), .ZN(n19420) );
  NOR3_X1 U21241 ( .A1(n19395), .A2(n17938), .A3(n19575), .ZN(n17941) );
  NOR2_X1 U21242 ( .A1(n19027), .A2(n19605), .ZN(n17940) );
  OAI21_X1 U21243 ( .B1(n17941), .B2(n17940), .A(n17939), .ZN(n17960) );
  NAND3_X1 U21244 ( .A1(n19027), .A2(n19587), .A3(n17942), .ZN(n17943) );
  AOI21_X1 U21245 ( .B1(n17954), .B2(n17944), .A(n17943), .ZN(n17953) );
  NAND2_X1 U21246 ( .A1(n17945), .A2(n20057), .ZN(n17950) );
  INV_X1 U21247 ( .A(n17946), .ZN(n17947) );
  NOR3_X1 U21248 ( .A1(n17948), .A2(n17947), .A3(n19575), .ZN(n17949) );
  OAI211_X1 U21249 ( .C1(n17951), .C2(n19401), .A(n17950), .B(n17949), .ZN(
        n17952) );
  OAI211_X1 U21250 ( .C1(n17953), .C2(n17952), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n19613), .ZN(n17958) );
  INV_X1 U21251 ( .A(n19026), .ZN(n17956) );
  INV_X1 U21252 ( .A(n17954), .ZN(n17955) );
  NAND3_X1 U21253 ( .A1(n17956), .A2(n19530), .A3(n17955), .ZN(n17957) );
  NAND4_X1 U21254 ( .A1(n17960), .A2(n17959), .A3(n17958), .A4(n17957), .ZN(
        P3_U2834) );
  NAND2_X1 U21255 ( .A1(n19404), .A2(n19401), .ZN(n19408) );
  AND2_X1 U21256 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n19495), .ZN(
        n17961) );
  AOI21_X1 U21257 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17961), .A(
        n17966), .ZN(n17963) );
  AOI211_X1 U21258 ( .C1(n17964), .C2(n19408), .A(n17963), .B(n17962), .ZN(
        n17972) );
  NOR2_X1 U21259 ( .A1(n19410), .A2(n19495), .ZN(n19472) );
  OAI21_X1 U21260 ( .B1(n19472), .B2(n19518), .A(n17965), .ZN(n19511) );
  OAI211_X1 U21261 ( .C1(n17966), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n17972), .B(n19511), .ZN(n17967) );
  NAND3_X1 U21262 ( .A1(n17967), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        n19603), .ZN(n17970) );
  AOI22_X1 U21263 ( .A1(n19530), .A2(n17968), .B1(n19566), .B2(
        P3_REIP_REG_11__SCAN_IN), .ZN(n17969) );
  OAI211_X1 U21264 ( .C1(n19519), .C2(n17971), .A(n17970), .B(n17969), .ZN(
        P3_U2851) );
  OR2_X1 U21265 ( .A1(n17974), .A2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17984) );
  OAI21_X1 U21266 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n19516), .A(
        n17972), .ZN(n17973) );
  OAI211_X1 U21267 ( .C1(n17973), .C2(n19472), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n19603), .ZN(n17983) );
  AOI21_X1 U21268 ( .B1(n19200), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17981) );
  NAND2_X1 U21269 ( .A1(n17975), .A2(n17974), .ZN(n17980) );
  INV_X1 U21270 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17976) );
  NOR3_X1 U21271 ( .A1(n17977), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        n17976), .ZN(n17978) );
  AOI211_X1 U21272 ( .C1(n17981), .C2(n17980), .A(n17979), .B(n17978), .ZN(
        n19255) );
  AOI22_X1 U21273 ( .A1(n19255), .A2(n19530), .B1(n19566), .B2(
        P3_REIP_REG_10__SCAN_IN), .ZN(n17982) );
  OAI211_X1 U21274 ( .C1(n19519), .C2(n17984), .A(n17983), .B(n17982), .ZN(
        P3_U2852) );
  NAND2_X1 U21275 ( .A1(n12089), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19618) );
  AND3_X1 U21276 ( .A1(n17985), .A2(n19614), .A3(n19616), .ZN(n17986) );
  OAI21_X1 U21277 ( .B1(n20198), .B2(n17986), .A(n19912), .ZN(n19623) );
  NAND2_X1 U21278 ( .A1(n19618), .A2(n19623), .ZN(n17989) );
  INV_X1 U21279 ( .A(n17989), .ZN(n17988) );
  OAI22_X1 U21280 ( .A1(n19307), .A2(n20211), .B1(n12089), .B2(n21986), .ZN(
        n17991) );
  NAND3_X1 U21281 ( .A1(n12088), .A2(n19623), .A3(n17991), .ZN(n17987) );
  OAI221_X1 U21282 ( .B1(n12088), .B2(n17988), .C1(n12088), .C2(n19911), .A(
        n17987), .ZN(P3_U2864) );
  NAND2_X1 U21283 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19839) );
  NOR2_X1 U21284 ( .A1(n19307), .A2(n20211), .ZN(n17990) );
  AOI221_X1 U21285 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n19839), .C1(n17990), 
        .C2(n19839), .A(n17989), .ZN(n19622) );
  INV_X1 U21286 ( .A(n19911), .ZN(n19967) );
  OAI221_X1 U21287 ( .B1(n19967), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n19967), .C2(n17991), .A(n19623), .ZN(n19620) );
  AOI22_X1 U21288 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19622), .B1(
        n19620), .B2(n20085), .ZN(P3_U2865) );
  NOR2_X1 U21289 ( .A1(n17992), .A2(n18030), .ZN(n18038) );
  INV_X1 U21290 ( .A(n17993), .ZN(n17994) );
  OAI211_X1 U21291 ( .C1(n10144), .C2(n17995), .A(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n17994), .ZN(n17999) );
  INV_X1 U21292 ( .A(n17996), .ZN(n17998) );
  OAI211_X1 U21293 ( .C1(n21665), .C2(n17999), .A(n17998), .B(n17997), .ZN(
        n18001) );
  NAND2_X1 U21294 ( .A1(n21665), .A2(n17999), .ZN(n18000) );
  NAND2_X1 U21295 ( .A1(n18001), .A2(n18000), .ZN(n18003) );
  INV_X1 U21296 ( .A(n18003), .ZN(n18002) );
  NOR2_X1 U21297 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18002), .ZN(
        n18004) );
  OAI22_X1 U21298 ( .A1(n18005), .A2(n18004), .B1(n18003), .B2(n21306), .ZN(
        n18008) );
  INV_X1 U21299 ( .A(n18006), .ZN(n18007) );
  AOI21_X1 U21300 ( .B1(n18008), .B2(n18007), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18010) );
  NOR2_X1 U21301 ( .A1(n18008), .A2(n18007), .ZN(n18009) );
  OAI21_X1 U21302 ( .B1(n18010), .B2(n18009), .A(n21303), .ZN(n18020) );
  NOR2_X1 U21303 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(P1_MORE_REG_SCAN_IN), .ZN(
        n18014) );
  OAI211_X1 U21304 ( .C1(n18014), .C2(n18013), .A(n18012), .B(n18011), .ZN(
        n18015) );
  OR2_X1 U21305 ( .A1(n18016), .A2(n18015), .ZN(n18017) );
  NOR2_X1 U21306 ( .A1(n18018), .A2(n18017), .ZN(n18019) );
  AND2_X1 U21307 ( .A1(n18020), .A2(n18019), .ZN(n18029) );
  OR2_X1 U21308 ( .A1(n18092), .A2(n18021), .ZN(n18027) );
  INV_X1 U21309 ( .A(n18022), .ZN(n18023) );
  NOR3_X1 U21310 ( .A1(n18025), .A2(n18024), .A3(n18023), .ZN(n18026) );
  AOI21_X1 U21311 ( .B1(n18028), .B2(n18027), .A(n18026), .ZN(n18094) );
  OAI221_X1 U21312 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n18029), 
        .A(n18094), .ZN(n18100) );
  NAND2_X1 U21313 ( .A1(n18100), .A2(n21733), .ZN(n18037) );
  INV_X1 U21314 ( .A(n18029), .ZN(n18033) );
  OAI211_X1 U21315 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n18092), .A(n18031), 
        .B(n18030), .ZN(n18032) );
  AOI21_X1 U21316 ( .B1(n18034), .B2(n18033), .A(n18032), .ZN(n18035) );
  AND2_X1 U21317 ( .A1(n18100), .A2(n18035), .ZN(n18036) );
  OAI22_X1 U21318 ( .A1(n18038), .A2(n18037), .B1(n18036), .B2(n21733), .ZN(
        P1_U3161) );
  INV_X1 U21319 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n21751) );
  INV_X1 U21320 ( .A(HOLD), .ZN(n21742) );
  NOR2_X1 U21321 ( .A1(n21751), .A2(n21742), .ZN(n21738) );
  AOI22_X1 U21322 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n18040) );
  NAND2_X1 U21323 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n21822), .ZN(n21741) );
  OAI211_X1 U21324 ( .C1(n21738), .C2(n18040), .A(n18039), .B(n21741), .ZN(
        P1_U3195) );
  INV_X1 U21325 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n18230) );
  NOR2_X1 U21326 ( .A1(n21237), .A2(n18230), .ZN(P1_U2905) );
  AOI21_X1 U21327 ( .B1(n18134), .B2(n12578), .A(n18041), .ZN(n18042) );
  OR2_X1 U21328 ( .A1(n20896), .A2(n18042), .ZN(n21084) );
  NOR2_X1 U21329 ( .A1(n18043), .A2(n21084), .ZN(P2_U3047) );
  AOI22_X1 U21330 ( .A1(n18048), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n18072), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n18047) );
  XNOR2_X1 U21331 ( .A(n18044), .B(n18069), .ZN(n18045) );
  XNOR2_X1 U21332 ( .A(n15999), .B(n18045), .ZN(n18066) );
  AOI22_X1 U21333 ( .A1(n18066), .A2(n11864), .B1(n18052), .B2(n21159), .ZN(
        n18046) );
  OAI211_X1 U21334 ( .C1(n18056), .C2(n21162), .A(n18047), .B(n18046), .ZN(
        P1_U2992) );
  AOI22_X1 U21335 ( .A1(n18048), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n18072), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n18054) );
  NAND2_X1 U21336 ( .A1(n9876), .A2(n18050), .ZN(n18051) );
  XNOR2_X1 U21337 ( .A(n18049), .B(n18051), .ZN(n18073) );
  AOI22_X1 U21338 ( .A1(n18073), .A2(n11864), .B1(n21169), .B2(n18052), .ZN(
        n18053) );
  OAI211_X1 U21339 ( .C1(n18056), .C2(n21172), .A(n18054), .B(n18053), .ZN(
        P1_U2993) );
  OAI22_X1 U21340 ( .A1(n21178), .A2(n18057), .B1(n21182), .B2(n18056), .ZN(
        n18058) );
  AOI21_X1 U21341 ( .B1(n18083), .B2(n11864), .A(n18058), .ZN(n18060) );
  INV_X1 U21342 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n21757) );
  NOR2_X1 U21343 ( .A1(n21291), .A2(n21757), .ZN(n18078) );
  INV_X1 U21344 ( .A(n18078), .ZN(n18059) );
  OAI211_X1 U21345 ( .C1(n18062), .C2(n18061), .A(n18060), .B(n18059), .ZN(
        P1_U2994) );
  INV_X1 U21346 ( .A(n18063), .ZN(n21152) );
  AOI22_X1 U21347 ( .A1(n21282), .A2(n21152), .B1(n18072), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n18068) );
  INV_X1 U21348 ( .A(n18064), .ZN(n18065) );
  AOI22_X1 U21349 ( .A1(n18066), .A2(n21286), .B1(n18069), .B2(n18065), .ZN(
        n18067) );
  OAI211_X1 U21350 ( .C1(n18070), .C2(n18069), .A(n18068), .B(n18067), .ZN(
        P1_U3024) );
  INV_X1 U21351 ( .A(n18071), .ZN(n21163) );
  AOI22_X1 U21352 ( .A1(n21282), .A2(n21163), .B1(n18072), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n18076) );
  AOI22_X1 U21353 ( .A1(n18074), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B1(
        n21286), .B2(n18073), .ZN(n18075) );
  OAI211_X1 U21354 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n18077), .A(
        n18076), .B(n18075), .ZN(P1_U3025) );
  AOI21_X1 U21355 ( .B1(n21282), .B2(n21175), .A(n18078), .ZN(n18079) );
  OAI21_X1 U21356 ( .B1(n18081), .B2(n18080), .A(n18079), .ZN(n18082) );
  AOI21_X1 U21357 ( .B1(n18083), .B2(n21286), .A(n18082), .ZN(n18084) );
  OAI21_X1 U21358 ( .B1(n21290), .B2(n18085), .A(n18084), .ZN(P1_U3026) );
  NAND3_X1 U21359 ( .A1(n21183), .A2(n18087), .A3(n18086), .ZN(n18090) );
  OAI22_X1 U21360 ( .A1(n18091), .A2(n18090), .B1(n18089), .B2(n18088), .ZN(
        P1_U3468) );
  NAND2_X1 U21361 ( .A1(n11673), .A2(n18092), .ZN(n18098) );
  AOI21_X1 U21362 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n18100), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n18097) );
  NOR2_X1 U21363 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21822), .ZN(n18093) );
  OAI221_X1 U21364 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(
        P1_STATEBS16_REG_SCAN_IN), .C1(n21733), .C2(n18093), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n21734) );
  AOI21_X1 U21365 ( .B1(n21734), .B2(n18095), .A(n18094), .ZN(n18096) );
  AOI211_X1 U21366 ( .C1(n21823), .C2(n18098), .A(n18097), .B(n18096), .ZN(
        P1_U3162) );
  OAI221_X1 U21367 ( .B1(n11673), .B2(P1_STATE2_REG_0__SCAN_IN), .C1(n11673), 
        .C2(n18100), .A(n18099), .ZN(P1_U3466) );
  AOI22_X1 U21368 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n20343), .B1(n18102), 
        .B2(n18101), .ZN(n18111) );
  INV_X1 U21369 ( .A(n18103), .ZN(n18109) );
  AOI222_X1 U21370 ( .A1(n18109), .A2(n18108), .B1(n18107), .B2(n18106), .C1(
        n18105), .C2(n18104), .ZN(n18110) );
  OAI211_X1 U21371 ( .C1(n18113), .C2(n18112), .A(n18111), .B(n18110), .ZN(
        P2_U3008) );
  INV_X1 U21372 ( .A(n18114), .ZN(n18117) );
  INV_X1 U21373 ( .A(n18115), .ZN(n18116) );
  AOI22_X1 U21374 ( .A1(n18118), .A2(n18117), .B1(n18116), .B2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18128) );
  AOI21_X1 U21375 ( .B1(n18120), .B2(n13822), .A(n18119), .ZN(n18121) );
  OAI21_X1 U21376 ( .B1(n18123), .B2(n18122), .A(n18121), .ZN(n18124) );
  AOI21_X1 U21377 ( .B1(n18126), .B2(n18125), .A(n18124), .ZN(n18127) );
  OAI211_X1 U21378 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n18129), .A(
        n18128), .B(n18127), .ZN(P2_U3046) );
  INV_X1 U21379 ( .A(n18130), .ZN(n18131) );
  AOI211_X1 U21380 ( .C1(n18134), .C2(n18133), .A(n18132), .B(n18131), .ZN(
        n18141) );
  MUX2_X1 U21381 ( .A(n18136), .B(n18135), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n18139) );
  OAI22_X1 U21382 ( .A1(n18139), .A2(n18138), .B1(n18137), .B2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n18140) );
  OAI211_X1 U21383 ( .C1(n18143), .C2(n18142), .A(n18141), .B(n18140), .ZN(
        P2_U3176) );
  NOR3_X1 U21384 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n18145) );
  NOR4_X1 U21385 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n18144) );
  NAND4_X1 U21386 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n18145), .A3(n18144), .A4(
        U215), .ZN(U213) );
  INV_X1 U21387 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n18229) );
  NOR2_X2 U21388 ( .A1(n18189), .A2(n18146), .ZN(n18191) );
  OAI222_X1 U21389 ( .A1(U212), .A2(n18229), .B1(n18195), .B2(n18147), .C1(
        U214), .C2(n18230), .ZN(U216) );
  AOI222_X1 U21390 ( .A1(n18193), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n18191), 
        .B2(BUF1_REG_30__SCAN_IN), .C1(n18189), .C2(P1_DATAO_REG_30__SCAN_IN), 
        .ZN(n18148) );
  INV_X1 U21391 ( .A(n18148), .ZN(U217) );
  INV_X1 U21392 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n18150) );
  AOI22_X1 U21393 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n18189), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n18193), .ZN(n18149) );
  OAI21_X1 U21394 ( .B1(n18150), .B2(n18195), .A(n18149), .ZN(U218) );
  AOI222_X1 U21395 ( .A1(n18193), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(n18191), 
        .B2(BUF1_REG_28__SCAN_IN), .C1(n18189), .C2(P1_DATAO_REG_28__SCAN_IN), 
        .ZN(n18151) );
  INV_X1 U21396 ( .A(n18151), .ZN(U219) );
  AOI22_X1 U21397 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n18189), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n18193), .ZN(n18152) );
  OAI21_X1 U21398 ( .B1(n18153), .B2(n18195), .A(n18152), .ZN(U220) );
  INV_X1 U21399 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n21983) );
  AOI22_X1 U21400 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n18189), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n18193), .ZN(n18154) );
  OAI21_X1 U21401 ( .B1(n21983), .B2(n18195), .A(n18154), .ZN(U221) );
  INV_X1 U21402 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n18156) );
  AOI22_X1 U21403 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n18189), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n18193), .ZN(n18155) );
  OAI21_X1 U21404 ( .B1(n18156), .B2(n18195), .A(n18155), .ZN(U222) );
  INV_X1 U21405 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n18158) );
  AOI22_X1 U21406 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n18189), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n18193), .ZN(n18157) );
  OAI21_X1 U21407 ( .B1(n18158), .B2(n18195), .A(n18157), .ZN(U223) );
  INV_X1 U21408 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n18160) );
  AOI22_X1 U21409 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n18189), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n18193), .ZN(n18159) );
  OAI21_X1 U21410 ( .B1(n18160), .B2(n18195), .A(n18159), .ZN(U224) );
  AOI222_X1 U21411 ( .A1(n18189), .A2(P1_DATAO_REG_22__SCAN_IN), .B1(n18191), 
        .B2(BUF1_REG_22__SCAN_IN), .C1(n18193), .C2(P2_DATAO_REG_22__SCAN_IN), 
        .ZN(n18161) );
  INV_X1 U21412 ( .A(n18161), .ZN(U225) );
  INV_X1 U21413 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n18163) );
  AOI22_X1 U21414 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n18189), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n18193), .ZN(n18162) );
  OAI21_X1 U21415 ( .B1(n18163), .B2(n18195), .A(n18162), .ZN(U226) );
  INV_X1 U21416 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n22130) );
  AOI22_X1 U21417 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n18189), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n18193), .ZN(n18164) );
  OAI21_X1 U21418 ( .B1(n22130), .B2(n18195), .A(n18164), .ZN(U227) );
  INV_X1 U21419 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n18166) );
  AOI22_X1 U21420 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n18189), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n18193), .ZN(n18165) );
  OAI21_X1 U21421 ( .B1(n18166), .B2(n18195), .A(n18165), .ZN(U228) );
  AOI22_X1 U21422 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n18189), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n18193), .ZN(n18167) );
  OAI21_X1 U21423 ( .B1(n18168), .B2(n18195), .A(n18167), .ZN(U229) );
  AOI222_X1 U21424 ( .A1(n18193), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n18191), 
        .B2(BUF1_REG_17__SCAN_IN), .C1(n18189), .C2(P1_DATAO_REG_17__SCAN_IN), 
        .ZN(n18169) );
  INV_X1 U21425 ( .A(n18169), .ZN(U230) );
  INV_X1 U21426 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n18171) );
  AOI22_X1 U21427 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n18189), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n18193), .ZN(n18170) );
  OAI21_X1 U21428 ( .B1(n18171), .B2(n18195), .A(n18170), .ZN(U231) );
  INV_X1 U21429 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n21227) );
  AOI22_X1 U21430 ( .A1(BUF1_REG_15__SCAN_IN), .A2(n18191), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n18193), .ZN(n18172) );
  OAI21_X1 U21431 ( .B1(n21227), .B2(U214), .A(n18172), .ZN(U232) );
  INV_X1 U21432 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n18174) );
  AOI22_X1 U21433 ( .A1(BUF1_REG_14__SCAN_IN), .A2(n18191), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n18189), .ZN(n18173) );
  OAI21_X1 U21434 ( .B1(n18174), .B2(U212), .A(n18173), .ZN(U233) );
  INV_X1 U21435 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n18176) );
  AOI22_X1 U21436 ( .A1(BUF1_REG_13__SCAN_IN), .A2(n18191), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n18189), .ZN(n18175) );
  OAI21_X1 U21437 ( .B1(n18176), .B2(U212), .A(n18175), .ZN(U234) );
  INV_X1 U21438 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n18208) );
  AOI22_X1 U21439 ( .A1(BUF1_REG_12__SCAN_IN), .A2(n18191), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n18189), .ZN(n18177) );
  OAI21_X1 U21440 ( .B1(n18208), .B2(U212), .A(n18177), .ZN(U235) );
  INV_X1 U21441 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n21856) );
  AOI22_X1 U21442 ( .A1(BUF1_REG_11__SCAN_IN), .A2(n18191), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n18193), .ZN(n18178) );
  OAI21_X1 U21443 ( .B1(n21856), .B2(U214), .A(n18178), .ZN(U236) );
  AOI22_X1 U21444 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n18189), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n18193), .ZN(n18179) );
  OAI21_X1 U21445 ( .B1(n18180), .B2(n18195), .A(n18179), .ZN(U237) );
  INV_X1 U21446 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n18205) );
  AOI22_X1 U21447 ( .A1(BUF1_REG_9__SCAN_IN), .A2(n18191), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n18189), .ZN(n18181) );
  OAI21_X1 U21448 ( .B1(n18205), .B2(U212), .A(n18181), .ZN(U238) );
  INV_X1 U21449 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n18183) );
  AOI22_X1 U21450 ( .A1(BUF1_REG_8__SCAN_IN), .A2(n18191), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n18189), .ZN(n18182) );
  OAI21_X1 U21451 ( .B1(n18183), .B2(U212), .A(n18182), .ZN(U239) );
  INV_X1 U21452 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n18203) );
  AOI22_X1 U21453 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n18191), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n18189), .ZN(n18184) );
  OAI21_X1 U21454 ( .B1(n18203), .B2(U212), .A(n18184), .ZN(U240) );
  INV_X1 U21455 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n18202) );
  AOI22_X1 U21456 ( .A1(BUF1_REG_6__SCAN_IN), .A2(n18191), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n18189), .ZN(n18185) );
  OAI21_X1 U21457 ( .B1(n18202), .B2(U212), .A(n18185), .ZN(U241) );
  AOI22_X1 U21458 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n18189), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n18193), .ZN(n18186) );
  OAI21_X1 U21459 ( .B1(n14574), .B2(n18195), .A(n18186), .ZN(U242) );
  AOI22_X1 U21460 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n18189), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n18193), .ZN(n18187) );
  OAI21_X1 U21461 ( .B1(n14259), .B2(n18195), .A(n18187), .ZN(U243) );
  INV_X1 U21462 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n18199) );
  AOI22_X1 U21463 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n18191), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n18189), .ZN(n18188) );
  OAI21_X1 U21464 ( .B1(n18199), .B2(U212), .A(n18188), .ZN(U244) );
  AOI22_X1 U21465 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n18189), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n18193), .ZN(n18190) );
  OAI21_X1 U21466 ( .B1(n13511), .B2(n18195), .A(n18190), .ZN(U245) );
  INV_X1 U21467 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n18197) );
  AOI22_X1 U21468 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n18191), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n18189), .ZN(n18192) );
  OAI21_X1 U21469 ( .B1(n18197), .B2(U212), .A(n18192), .ZN(U246) );
  AOI22_X1 U21470 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n18189), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n18193), .ZN(n18194) );
  OAI21_X1 U21471 ( .B1(n13524), .B2(n18195), .A(n18194), .ZN(U247) );
  OAI22_X1 U21472 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n18227), .ZN(n18196) );
  INV_X1 U21473 ( .A(n18196), .ZN(U251) );
  AOI22_X1 U21474 ( .A1(n18227), .A2(n18197), .B1(n21987), .B2(U215), .ZN(U252) );
  OAI22_X1 U21475 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n18218), .ZN(n18198) );
  INV_X1 U21476 ( .A(n18198), .ZN(U253) );
  AOI22_X1 U21477 ( .A1(n18227), .A2(n18199), .B1(n19637), .B2(U215), .ZN(U254) );
  OAI22_X1 U21478 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n18218), .ZN(n18200) );
  INV_X1 U21479 ( .A(n18200), .ZN(U255) );
  OAI22_X1 U21480 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n18218), .ZN(n18201) );
  INV_X1 U21481 ( .A(n18201), .ZN(U256) );
  AOI22_X1 U21482 ( .A1(n18227), .A2(n18202), .B1(n19649), .B2(U215), .ZN(U257) );
  AOI22_X1 U21483 ( .A1(n18227), .A2(n18203), .B1(n21919), .B2(U215), .ZN(U258) );
  OAI22_X1 U21484 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n18218), .ZN(n18204) );
  INV_X1 U21485 ( .A(n18204), .ZN(U259) );
  AOI22_X1 U21486 ( .A1(n18227), .A2(n18205), .B1(n19007), .B2(U215), .ZN(U260) );
  OAI22_X1 U21487 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n18218), .ZN(n18206) );
  INV_X1 U21488 ( .A(n18206), .ZN(U261) );
  OAI22_X1 U21489 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n18218), .ZN(n18207) );
  INV_X1 U21490 ( .A(n18207), .ZN(U262) );
  AOI22_X1 U21491 ( .A1(n18227), .A2(n18208), .B1(n19014), .B2(U215), .ZN(U263) );
  OAI22_X1 U21492 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n18218), .ZN(n18209) );
  INV_X1 U21493 ( .A(n18209), .ZN(U264) );
  OAI22_X1 U21494 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n18227), .ZN(n18210) );
  INV_X1 U21495 ( .A(n18210), .ZN(U265) );
  OAI22_X1 U21496 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n18218), .ZN(n18211) );
  INV_X1 U21497 ( .A(n18211), .ZN(U266) );
  OAI22_X1 U21498 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n18227), .ZN(n18212) );
  INV_X1 U21499 ( .A(n18212), .ZN(U267) );
  OAI22_X1 U21500 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n18218), .ZN(n18213) );
  INV_X1 U21501 ( .A(n18213), .ZN(U268) );
  OAI22_X1 U21502 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n18227), .ZN(n18214) );
  INV_X1 U21503 ( .A(n18214), .ZN(U269) );
  OAI22_X1 U21504 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n18227), .ZN(n18215) );
  INV_X1 U21505 ( .A(n18215), .ZN(U270) );
  OAI22_X1 U21506 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n18227), .ZN(n18216) );
  INV_X1 U21507 ( .A(n18216), .ZN(U271) );
  OAI22_X1 U21508 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n18227), .ZN(n18217) );
  INV_X1 U21509 ( .A(n18217), .ZN(U272) );
  INV_X1 U21510 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n22003) );
  AOI22_X1 U21511 ( .A1(n18227), .A2(n22003), .B1(n16904), .B2(U215), .ZN(U273) );
  OAI22_X1 U21512 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n18218), .ZN(n18219) );
  INV_X1 U21513 ( .A(n18219), .ZN(U274) );
  OAI22_X1 U21514 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n18227), .ZN(n18220) );
  INV_X1 U21515 ( .A(n18220), .ZN(U275) );
  OAI22_X1 U21516 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n18227), .ZN(n18221) );
  INV_X1 U21517 ( .A(n18221), .ZN(U276) );
  OAI22_X1 U21518 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n18227), .ZN(n18222) );
  INV_X1 U21519 ( .A(n18222), .ZN(U277) );
  OAI22_X1 U21520 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n18227), .ZN(n18223) );
  INV_X1 U21521 ( .A(n18223), .ZN(U278) );
  OAI22_X1 U21522 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n18227), .ZN(n18224) );
  INV_X1 U21523 ( .A(n18224), .ZN(U279) );
  OAI22_X1 U21524 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n18227), .ZN(n18225) );
  INV_X1 U21525 ( .A(n18225), .ZN(U280) );
  OAI22_X1 U21526 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n18227), .ZN(n18226) );
  INV_X1 U21527 ( .A(n18226), .ZN(U281) );
  INV_X1 U21528 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19656) );
  AOI22_X1 U21529 ( .A1(n18227), .A2(n18229), .B1(n19656), .B2(U215), .ZN(U282) );
  INV_X1 U21530 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n18228) );
  AOI222_X1 U21531 ( .A1(n18230), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n18229), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n18228), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n18231) );
  INV_X2 U21532 ( .A(n18233), .ZN(n18232) );
  INV_X1 U21533 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n20150) );
  INV_X1 U21534 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20996) );
  AOI22_X1 U21535 ( .A1(n18232), .A2(n20150), .B1(n20996), .B2(n18233), .ZN(
        U347) );
  INV_X1 U21536 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n20148) );
  INV_X1 U21537 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20995) );
  AOI22_X1 U21538 ( .A1(n18232), .A2(n20148), .B1(n20995), .B2(n18233), .ZN(
        U348) );
  INV_X1 U21539 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n20146) );
  INV_X1 U21540 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20993) );
  AOI22_X1 U21541 ( .A1(n18232), .A2(n20146), .B1(n20993), .B2(n18233), .ZN(
        U349) );
  INV_X1 U21542 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n20145) );
  INV_X1 U21543 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20991) );
  AOI22_X1 U21544 ( .A1(n18232), .A2(n20145), .B1(n20991), .B2(n18233), .ZN(
        U350) );
  INV_X1 U21545 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n20143) );
  INV_X1 U21546 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20989) );
  AOI22_X1 U21547 ( .A1(n18232), .A2(n20143), .B1(n20989), .B2(n18233), .ZN(
        U351) );
  INV_X1 U21548 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n20140) );
  INV_X1 U21549 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20987) );
  AOI22_X1 U21550 ( .A1(n18232), .A2(n20140), .B1(n20987), .B2(n18233), .ZN(
        U352) );
  INV_X1 U21551 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n21908) );
  INV_X1 U21552 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20985) );
  AOI22_X1 U21553 ( .A1(n18232), .A2(n21908), .B1(n20985), .B2(n18233), .ZN(
        U353) );
  INV_X1 U21554 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n20138) );
  INV_X1 U21555 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20982) );
  AOI22_X1 U21556 ( .A1(n18232), .A2(n20138), .B1(n20982), .B2(n18233), .ZN(
        U354) );
  INV_X1 U21557 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n20188) );
  INV_X1 U21558 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n21032) );
  AOI22_X1 U21559 ( .A1(n18232), .A2(n20188), .B1(n21032), .B2(n18233), .ZN(
        U355) );
  INV_X1 U21560 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n20184) );
  INV_X1 U21561 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n21029) );
  AOI22_X1 U21562 ( .A1(n18232), .A2(n20184), .B1(n21029), .B2(n18233), .ZN(
        U356) );
  INV_X1 U21563 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n20181) );
  INV_X1 U21564 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n21027) );
  AOI22_X1 U21565 ( .A1(n18232), .A2(n20181), .B1(n21027), .B2(n18233), .ZN(
        U357) );
  INV_X1 U21566 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n20180) );
  INV_X1 U21567 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n21025) );
  AOI22_X1 U21568 ( .A1(n18232), .A2(n20180), .B1(n21025), .B2(n18233), .ZN(
        U358) );
  INV_X1 U21569 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n20177) );
  INV_X1 U21570 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n21024) );
  AOI22_X1 U21571 ( .A1(n18232), .A2(n20177), .B1(n21024), .B2(n18233), .ZN(
        U359) );
  INV_X1 U21572 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n22040) );
  INV_X1 U21573 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n21022) );
  AOI22_X1 U21574 ( .A1(n18232), .A2(n22040), .B1(n21022), .B2(n18233), .ZN(
        U360) );
  INV_X1 U21575 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n20175) );
  INV_X1 U21576 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n21020) );
  AOI22_X1 U21577 ( .A1(n18232), .A2(n20175), .B1(n21020), .B2(n18233), .ZN(
        U361) );
  INV_X1 U21578 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n20174) );
  INV_X1 U21579 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n21018) );
  AOI22_X1 U21580 ( .A1(n18232), .A2(n20174), .B1(n21018), .B2(n18233), .ZN(
        U362) );
  INV_X1 U21581 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n20172) );
  INV_X1 U21582 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n21016) );
  AOI22_X1 U21583 ( .A1(n18232), .A2(n20172), .B1(n21016), .B2(n18233), .ZN(
        U363) );
  INV_X1 U21584 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n20170) );
  INV_X1 U21585 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n21014) );
  AOI22_X1 U21586 ( .A1(n18232), .A2(n20170), .B1(n21014), .B2(n18233), .ZN(
        U364) );
  INV_X1 U21587 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n20136) );
  INV_X1 U21588 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20980) );
  AOI22_X1 U21589 ( .A1(n18232), .A2(n20136), .B1(n20980), .B2(n18233), .ZN(
        U365) );
  INV_X1 U21590 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n20167) );
  INV_X1 U21591 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n21012) );
  AOI22_X1 U21592 ( .A1(n18232), .A2(n20167), .B1(n21012), .B2(n18233), .ZN(
        U366) );
  INV_X1 U21593 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n20166) );
  INV_X1 U21594 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n21011) );
  AOI22_X1 U21595 ( .A1(n18232), .A2(n20166), .B1(n21011), .B2(n18233), .ZN(
        U367) );
  INV_X1 U21596 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n20164) );
  INV_X1 U21597 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n21009) );
  AOI22_X1 U21598 ( .A1(n18232), .A2(n20164), .B1(n21009), .B2(n18233), .ZN(
        U368) );
  INV_X1 U21599 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n20161) );
  INV_X1 U21600 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n21008) );
  AOI22_X1 U21601 ( .A1(n18232), .A2(n20161), .B1(n21008), .B2(n18233), .ZN(
        U369) );
  INV_X1 U21602 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n22060) );
  INV_X1 U21603 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n21006) );
  AOI22_X1 U21604 ( .A1(n18232), .A2(n22060), .B1(n21006), .B2(n18233), .ZN(
        U370) );
  INV_X1 U21605 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n21876) );
  INV_X1 U21606 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n21004) );
  AOI22_X1 U21607 ( .A1(n18232), .A2(n21876), .B1(n21004), .B2(n18233), .ZN(
        U371) );
  INV_X1 U21608 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n20158) );
  INV_X1 U21609 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n21002) );
  AOI22_X1 U21610 ( .A1(n18232), .A2(n20158), .B1(n21002), .B2(n18233), .ZN(
        U372) );
  INV_X1 U21611 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n20156) );
  INV_X1 U21612 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n21001) );
  AOI22_X1 U21613 ( .A1(n18232), .A2(n20156), .B1(n21001), .B2(n18233), .ZN(
        U373) );
  INV_X1 U21614 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n20154) );
  INV_X1 U21615 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20999) );
  AOI22_X1 U21616 ( .A1(n18232), .A2(n20154), .B1(n20999), .B2(n18233), .ZN(
        U374) );
  INV_X1 U21617 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n20152) );
  INV_X1 U21618 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20997) );
  AOI22_X1 U21619 ( .A1(n18232), .A2(n20152), .B1(n20997), .B2(n18233), .ZN(
        U375) );
  INV_X1 U21620 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n20134) );
  AOI22_X1 U21621 ( .A1(n18232), .A2(n20134), .B1(n20978), .B2(n18233), .ZN(
        U376) );
  INV_X1 U21622 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n20133) );
  NAND2_X1 U21623 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n20133), .ZN(n20124) );
  AOI22_X1 U21624 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n20124), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n20131), .ZN(n20197) );
  AOI21_X1 U21625 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n20197), .ZN(n18234) );
  INV_X1 U21626 ( .A(n18234), .ZN(P3_U2633) );
  NAND2_X1 U21627 ( .A1(n20107), .A2(n21986), .ZN(n18238) );
  NOR2_X1 U21628 ( .A1(n18975), .A2(n18235), .ZN(n18236) );
  OAI21_X1 U21629 ( .B1(n18236), .B2(n18976), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n18237) );
  OAI21_X1 U21630 ( .B1(n18238), .B2(n20109), .A(n18237), .ZN(P3_U2634) );
  AOI21_X1 U21631 ( .B1(n20131), .B2(n20133), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n18239) );
  AOI22_X1 U21632 ( .A1(n20208), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n18239), 
        .B2(n20225), .ZN(P3_U2635) );
  OAI21_X1 U21633 ( .B1(n20118), .B2(BS16), .A(n20197), .ZN(n20195) );
  OAI21_X1 U21634 ( .B1(n20197), .B2(n20216), .A(n20195), .ZN(P3_U2636) );
  AOI211_X1 U21635 ( .C1(n18243), .C2(n18242), .A(n18241), .B(n18240), .ZN(
        n20066) );
  NOR2_X1 U21636 ( .A1(n20066), .A2(n20105), .ZN(n20209) );
  OAI21_X1 U21637 ( .B1(n20209), .B2(n19616), .A(n18244), .ZN(P3_U2637) );
  NOR4_X1 U21638 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18248) );
  NOR4_X1 U21639 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_14__SCAN_IN), .A3(P3_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18247) );
  NOR4_X1 U21640 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n18246) );
  NOR4_X1 U21641 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18245) );
  NAND4_X1 U21642 ( .A1(n18248), .A2(n18247), .A3(n18246), .A4(n18245), .ZN(
        n18254) );
  NOR4_X1 U21643 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_10__SCAN_IN), .A3(P3_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18252) );
  AOI211_X1 U21644 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_5__SCAN_IN), .B(
        P3_DATAWIDTH_REG_16__SCAN_IN), .ZN(n18251) );
  NOR4_X1 U21645 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_13__SCAN_IN), .ZN(n18250) );
  NOR4_X1 U21646 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n18249) );
  NAND4_X1 U21647 ( .A1(n18252), .A2(n18251), .A3(n18250), .A4(n18249), .ZN(
        n18253) );
  NOR2_X1 U21648 ( .A1(n18254), .A2(n18253), .ZN(n20204) );
  INV_X1 U21649 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18256) );
  NOR3_X1 U21650 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n18257) );
  OAI21_X1 U21651 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n18257), .A(n20204), .ZN(
        n18255) );
  OAI21_X1 U21652 ( .B1(n20204), .B2(n18256), .A(n18255), .ZN(P3_U2638) );
  INV_X1 U21653 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n20200) );
  INV_X1 U21654 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20196) );
  AOI21_X1 U21655 ( .B1(n20200), .B2(n20196), .A(n18257), .ZN(n18259) );
  INV_X1 U21656 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18258) );
  INV_X1 U21657 ( .A(n20204), .ZN(n20206) );
  AOI22_X1 U21658 ( .A1(n20204), .A2(n18259), .B1(n18258), .B2(n20206), .ZN(
        P3_U2639) );
  INV_X1 U21659 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n20183) );
  NAND3_X1 U21660 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n18283), .ZN(n18264) );
  OAI22_X1 U21661 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n18264), .B1(n18263), 
        .B2(n18593), .ZN(n18265) );
  INV_X1 U21662 ( .A(n18266), .ZN(n18267) );
  OAI21_X1 U21663 ( .B1(n18270), .B2(n18661), .A(n18267), .ZN(n18268) );
  AOI22_X1 U21664 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18481), .B1(
        n18596), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n18279) );
  AOI211_X1 U21665 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n18284), .A(n18270), .B(
        n18579), .ZN(n18275) );
  AOI211_X1 U21666 ( .C1(n18273), .C2(n18272), .A(n18271), .B(n18584), .ZN(
        n18274) );
  AOI211_X1 U21667 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n18296), .A(n18275), 
        .B(n18274), .ZN(n18278) );
  NAND2_X1 U21668 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n18276) );
  OAI211_X1 U21669 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n18283), .B(n18276), .ZN(n18277) );
  NAND3_X1 U21670 ( .A1(n18279), .A2(n18278), .A3(n18277), .ZN(P3_U2643) );
  INV_X1 U21671 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n20179) );
  AOI211_X1 U21672 ( .C1(n19028), .C2(n9850), .A(n18280), .B(n18584), .ZN(
        n18282) );
  OAI22_X1 U21673 ( .A1(n19031), .A2(n18593), .B1(n18522), .B2(n18669), .ZN(
        n18281) );
  AOI211_X1 U21674 ( .C1(n18283), .C2(n20179), .A(n18282), .B(n18281), .ZN(
        n18286) );
  OAI211_X1 U21675 ( .C1(n18290), .C2(n18669), .A(n18575), .B(n18284), .ZN(
        n18285) );
  OAI211_X1 U21676 ( .C1(n18287), .C2(n20179), .A(n18286), .B(n18285), .ZN(
        P3_U2644) );
  AOI22_X1 U21677 ( .A1(n18596), .A2(P3_EBX_REG_26__SCAN_IN), .B1(n18289), 
        .B2(n18288), .ZN(n18298) );
  AOI211_X1 U21678 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n18305), .A(n18290), .B(
        n18579), .ZN(n18295) );
  AOI211_X1 U21679 ( .C1(n18293), .C2(n18292), .A(n18291), .B(n18584), .ZN(
        n18294) );
  AOI211_X1 U21680 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n18296), .A(n18295), 
        .B(n18294), .ZN(n18297) );
  OAI211_X1 U21681 ( .C1(n19038), .C2(n18593), .A(n18298), .B(n18297), .ZN(
        P3_U2645) );
  INV_X1 U21682 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n22017) );
  OAI21_X1 U21683 ( .B1(n18311), .B2(n18568), .A(n18552), .ZN(n18325) );
  AOI21_X1 U21684 ( .B1(n18578), .B2(n22017), .A(n18325), .ZN(n18309) );
  AOI211_X1 U21685 ( .C1(n19058), .C2(n18300), .A(n18299), .B(n18584), .ZN(
        n18304) );
  NOR3_X1 U21686 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n18568), .A3(n18301), 
        .ZN(n18303) );
  OAI22_X1 U21687 ( .A1(n19056), .A2(n18593), .B1(n18522), .B2(n18306), .ZN(
        n18302) );
  NOR3_X1 U21688 ( .A1(n18304), .A2(n18303), .A3(n18302), .ZN(n18308) );
  OAI211_X1 U21689 ( .C1(n18312), .C2(n18306), .A(n18575), .B(n18305), .ZN(
        n18307) );
  OAI211_X1 U21690 ( .C1(n18309), .C2(n20176), .A(n18308), .B(n18307), .ZN(
        P3_U2646) );
  NOR2_X1 U21691 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n18568), .ZN(n18310) );
  AOI22_X1 U21692 ( .A1(n18596), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n18311), 
        .B2(n18310), .ZN(n18318) );
  AOI211_X1 U21693 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n18326), .A(n18312), .B(
        n18579), .ZN(n18316) );
  AOI211_X1 U21694 ( .C1(n19076), .C2(n18314), .A(n18313), .B(n18584), .ZN(
        n18315) );
  AOI211_X1 U21695 ( .C1(n18325), .C2(P3_REIP_REG_24__SCAN_IN), .A(n18316), 
        .B(n18315), .ZN(n18317) );
  OAI211_X1 U21696 ( .C1(n19068), .C2(n18593), .A(n18318), .B(n18317), .ZN(
        P3_U2647) );
  NAND2_X1 U21697 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n18319) );
  NAND2_X1 U21698 ( .A1(n18578), .A2(n18358), .ZN(n18369) );
  NOR2_X1 U21699 ( .A1(n18319), .A2(n18369), .ZN(n18354) );
  NAND2_X1 U21700 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n18354), .ZN(n18348) );
  OAI21_X1 U21701 ( .B1(n18337), .B2(n18348), .A(n20173), .ZN(n18324) );
  AOI211_X1 U21702 ( .C1(n19083), .C2(n18321), .A(n18320), .B(n18584), .ZN(
        n18323) );
  OAI22_X1 U21703 ( .A1(n19053), .A2(n18593), .B1(n18522), .B2(n21874), .ZN(
        n18322) );
  AOI211_X1 U21704 ( .C1(n18325), .C2(n18324), .A(n18323), .B(n18322), .ZN(
        n18328) );
  OAI211_X1 U21705 ( .C1(n18332), .C2(n21874), .A(n18575), .B(n18326), .ZN(
        n18327) );
  NAND2_X1 U21706 ( .A1(n18328), .A2(n18327), .ZN(P3_U2648) );
  INV_X1 U21707 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n20171) );
  AOI21_X1 U21708 ( .B1(n18578), .B2(n18329), .A(n18589), .ZN(n18351) );
  AOI211_X1 U21709 ( .C1(n19099), .C2(n18331), .A(n18330), .B(n18584), .ZN(
        n18336) );
  AOI211_X1 U21710 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n18343), .A(n18332), .B(
        n18579), .ZN(n18335) );
  AOI22_X1 U21711 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n18481), .B1(
        n18596), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n18333) );
  INV_X1 U21712 ( .A(n18333), .ZN(n18334) );
  NOR3_X1 U21713 ( .A1(n18336), .A2(n18335), .A3(n18334), .ZN(n18340) );
  INV_X1 U21714 ( .A(n18348), .ZN(n18338) );
  OAI211_X1 U21715 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(P3_REIP_REG_21__SCAN_IN), .A(n18338), .B(n18337), .ZN(n18339) );
  OAI211_X1 U21716 ( .C1(n20171), .C2(n18351), .A(n18340), .B(n18339), .ZN(
        P3_U2649) );
  INV_X1 U21717 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n20169) );
  AOI211_X1 U21718 ( .C1(n19115), .C2(n18342), .A(n18341), .B(n18584), .ZN(
        n18346) );
  OAI211_X1 U21719 ( .C1(n18349), .C2(n21897), .A(n18575), .B(n18343), .ZN(
        n18344) );
  OAI21_X1 U21720 ( .B1(n21897), .B2(n18522), .A(n18344), .ZN(n18345) );
  AOI211_X1 U21721 ( .C1(n18481), .C2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n18346), .B(n18345), .ZN(n18347) );
  OAI221_X1 U21722 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(n18348), .C1(n20169), 
        .C2(n18351), .A(n18347), .ZN(P3_U2650) );
  AOI211_X1 U21723 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n18365), .A(n18349), .B(
        n18579), .ZN(n18350) );
  AOI21_X1 U21724 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n18596), .A(n18350), .ZN(
        n18357) );
  INV_X1 U21725 ( .A(n18351), .ZN(n18355) );
  INV_X1 U21726 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n20168) );
  AOI211_X1 U21727 ( .C1(n19124), .C2(n18352), .A(n9874), .B(n18584), .ZN(
        n18353) );
  AOI221_X1 U21728 ( .B1(n18355), .B2(P3_REIP_REG_20__SCAN_IN), .C1(n18354), 
        .C2(n20168), .A(n18353), .ZN(n18356) );
  OAI211_X1 U21729 ( .C1(n19122), .C2(n18593), .A(n18357), .B(n18356), .ZN(
        P3_U2651) );
  NOR2_X1 U21730 ( .A1(n18358), .A2(n18568), .ZN(n18383) );
  NOR2_X1 U21731 ( .A1(n18589), .A2(n18383), .ZN(n18391) );
  OAI21_X1 U21732 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n18369), .A(n18391), 
        .ZN(n18364) );
  AOI211_X1 U21733 ( .C1(n19146), .C2(n18360), .A(n18359), .B(n18584), .ZN(
        n18363) );
  INV_X1 U21734 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n20163) );
  OR3_X1 U21735 ( .A1(n20163), .A2(n18369), .A3(P3_REIP_REG_19__SCAN_IN), .ZN(
        n18361) );
  OAI211_X1 U21736 ( .C1(n19143), .C2(n18593), .A(n19603), .B(n18361), .ZN(
        n18362) );
  AOI211_X1 U21737 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(n18364), .A(n18363), 
        .B(n18362), .ZN(n18367) );
  OAI211_X1 U21738 ( .C1(n18372), .C2(n18368), .A(n18575), .B(n18365), .ZN(
        n18366) );
  OAI211_X1 U21739 ( .C1(n18368), .C2(n18522), .A(n18367), .B(n18366), .ZN(
        P3_U2652) );
  AOI22_X1 U21740 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18481), .B1(
        n18596), .B2(P3_EBX_REG_18__SCAN_IN), .ZN(n18377) );
  NOR2_X1 U21741 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n18369), .ZN(n18375) );
  AOI211_X1 U21742 ( .C1(n19157), .C2(n18371), .A(n18370), .B(n18584), .ZN(
        n18374) );
  AOI211_X1 U21743 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n18381), .A(n18372), .B(
        n18579), .ZN(n18373) );
  NOR4_X1 U21744 ( .A1(n19556), .A2(n18375), .A3(n18374), .A4(n18373), .ZN(
        n18376) );
  OAI211_X1 U21745 ( .C1(n18391), .C2(n20163), .A(n18377), .B(n18376), .ZN(
        P3_U2653) );
  AOI211_X1 U21746 ( .C1(n18380), .C2(n18379), .A(n18378), .B(n18584), .ZN(
        n18389) );
  OAI211_X1 U21747 ( .C1(n18392), .C2(n18386), .A(n18575), .B(n18381), .ZN(
        n18382) );
  OAI21_X1 U21748 ( .B1(n18593), .B2(n19165), .A(n18382), .ZN(n18388) );
  INV_X1 U21749 ( .A(n18383), .ZN(n18384) );
  OAI22_X1 U21750 ( .A1(n18522), .A2(n18386), .B1(n18385), .B2(n18384), .ZN(
        n18387) );
  NOR4_X1 U21751 ( .A1(n19556), .A2(n18389), .A3(n18388), .A4(n18387), .ZN(
        n18390) );
  OAI21_X1 U21752 ( .B1(n18391), .B2(n20162), .A(n18390), .ZN(P3_U2654) );
  AOI22_X1 U21753 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n18481), .B1(
        n18596), .B2(P3_EBX_REG_16__SCAN_IN), .ZN(n18404) );
  NOR2_X1 U21754 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n18568), .ZN(n18394) );
  AOI211_X1 U21755 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n18414), .A(n18392), .B(
        n18579), .ZN(n18393) );
  AOI211_X1 U21756 ( .C1(n18395), .C2(n18394), .A(n19556), .B(n18393), .ZN(
        n18403) );
  AOI21_X1 U21757 ( .B1(n18421), .B2(n18578), .A(n18589), .ZN(n18432) );
  INV_X1 U21758 ( .A(n18432), .ZN(n18413) );
  NOR3_X1 U21759 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n18568), .A3(n18421), 
        .ZN(n18409) );
  OAI21_X1 U21760 ( .B1(n18413), .B2(n18409), .A(P3_REIP_REG_16__SCAN_IN), 
        .ZN(n18402) );
  NOR2_X1 U21761 ( .A1(n18418), .A2(n18428), .ZN(n18397) );
  OAI21_X1 U21762 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n18397), .A(
        n18396), .ZN(n19182) );
  OAI21_X1 U21763 ( .B1(n18418), .B2(n18398), .A(n10451), .ZN(n18400) );
  AOI21_X1 U21764 ( .B1(n19182), .B2(n18400), .A(n18584), .ZN(n18399) );
  OAI21_X1 U21765 ( .B1(n19182), .B2(n18400), .A(n18399), .ZN(n18401) );
  NAND4_X1 U21766 ( .A1(n18404), .A2(n18403), .A3(n18402), .A4(n18401), .ZN(
        P3_U2655) );
  INV_X1 U21767 ( .A(n18406), .ZN(n18408) );
  AOI221_X1 U21768 ( .B1(n18408), .B2(n18407), .C1(n18406), .C2(n18405), .A(
        n18584), .ZN(n18412) );
  AOI211_X1 U21769 ( .C1(n18596), .C2(P3_EBX_REG_15__SCAN_IN), .A(n19556), .B(
        n18409), .ZN(n18410) );
  INV_X1 U21770 ( .A(n18410), .ZN(n18411) );
  AOI211_X1 U21771 ( .C1(n18413), .C2(P3_REIP_REG_15__SCAN_IN), .A(n18412), 
        .B(n18411), .ZN(n18417) );
  OAI211_X1 U21772 ( .C1(n18419), .C2(n18415), .A(n18575), .B(n18414), .ZN(
        n18416) );
  OAI211_X1 U21773 ( .C1(n18593), .C2(n18418), .A(n18417), .B(n18416), .ZN(
        P3_U2656) );
  INV_X1 U21774 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n20157) );
  AOI211_X1 U21775 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n18437), .A(n18419), .B(
        n18579), .ZN(n18425) );
  NAND3_X1 U21776 ( .A1(n18421), .A2(n18420), .A3(n18578), .ZN(n18422) );
  OAI211_X1 U21777 ( .C1(n18522), .C2(n18423), .A(n19603), .B(n18422), .ZN(
        n18424) );
  AOI211_X1 U21778 ( .C1(n18481), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n18425), .B(n18424), .ZN(n18431) );
  AOI21_X1 U21779 ( .B1(n18426), .B2(n18527), .A(n10450), .ZN(n18450) );
  AOI21_X1 U21780 ( .B1(n10451), .B2(n18427), .A(n18450), .ZN(n18434) );
  INV_X1 U21781 ( .A(n18449), .ZN(n19215) );
  OAI221_X1 U21782 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19213), .C1(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .C2(n19215), .A(n18428), .ZN(
        n19195) );
  AOI21_X1 U21783 ( .B1(n18434), .B2(n19195), .A(n18584), .ZN(n18429) );
  OAI21_X1 U21784 ( .B1(n18434), .B2(n19195), .A(n18429), .ZN(n18430) );
  OAI211_X1 U21785 ( .C1(n18432), .C2(n20157), .A(n18431), .B(n18430), .ZN(
        P3_U2657) );
  INV_X1 U21786 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n19218) );
  NAND2_X1 U21787 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n19215), .ZN(
        n18433) );
  AOI22_X1 U21788 ( .A1(n19215), .A2(n19213), .B1(n19218), .B2(n18433), .ZN(
        n19221) );
  OR2_X1 U21789 ( .A1(n20113), .A2(n18434), .ZN(n18444) );
  NOR3_X1 U21790 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n18568), .A3(n18435), 
        .ZN(n18436) );
  AOI211_X1 U21791 ( .C1(n18596), .C2(P3_EBX_REG_13__SCAN_IN), .A(n19556), .B(
        n18436), .ZN(n18443) );
  OAI21_X1 U21792 ( .B1(n18448), .B2(n18568), .A(n18552), .ZN(n18458) );
  NOR2_X1 U21793 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n18568), .ZN(n18447) );
  OAI211_X1 U21794 ( .C1(n19218), .C2(n10450), .A(n19221), .B(n18520), .ZN(
        n18440) );
  OAI211_X1 U21795 ( .C1(n18445), .C2(n18438), .A(n18575), .B(n18437), .ZN(
        n18439) );
  OAI211_X1 U21796 ( .C1(n18593), .C2(n19218), .A(n18440), .B(n18439), .ZN(
        n18441) );
  AOI221_X1 U21797 ( .B1(n18458), .B2(P3_REIP_REG_13__SCAN_IN), .C1(n18447), 
        .C2(P3_REIP_REG_13__SCAN_IN), .A(n18441), .ZN(n18442) );
  OAI211_X1 U21798 ( .C1(n19221), .C2(n18444), .A(n18443), .B(n18442), .ZN(
        P3_U2658) );
  AOI211_X1 U21799 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n18460), .A(n18445), .B(
        n18579), .ZN(n18446) );
  AOI21_X1 U21800 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n18596), .A(n18446), .ZN(
        n18454) );
  AOI22_X1 U21801 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18481), .B1(
        n18448), .B2(n18447), .ZN(n18453) );
  INV_X1 U21802 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n19232) );
  AOI22_X1 U21803 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n19215), .B1(
        n18449), .B2(n19232), .ZN(n19235) );
  XOR2_X1 U21804 ( .A(n19235), .B(n18450), .Z(n18451) );
  AOI22_X1 U21805 ( .A1(n18598), .A2(n18451), .B1(P3_REIP_REG_12__SCAN_IN), 
        .B2(n18458), .ZN(n18452) );
  NAND4_X1 U21806 ( .A1(n18454), .A2(n18453), .A3(n18452), .A4(n19603), .ZN(
        P3_U2659) );
  AOI22_X1 U21807 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n18481), .B1(
        n18596), .B2(P3_EBX_REG_11__SCAN_IN), .ZN(n18464) );
  NAND3_X1 U21808 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n18483), .A3(
        n18484), .ZN(n18468) );
  OAI21_X1 U21809 ( .B1(n19251), .B2(n18468), .A(n10451), .ZN(n18455) );
  XOR2_X1 U21810 ( .A(n18456), .B(n18455), .Z(n18459) );
  NAND2_X1 U21811 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .ZN(n18515) );
  NOR3_X1 U21812 ( .A1(n18568), .A2(n18514), .A3(n18515), .ZN(n18498) );
  NAND2_X1 U21813 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n18498), .ZN(n18476) );
  OAI21_X1 U21814 ( .B1(n18477), .B2(n18476), .A(n20151), .ZN(n18457) );
  AOI22_X1 U21815 ( .A1(n18598), .A2(n18459), .B1(n18458), .B2(n18457), .ZN(
        n18463) );
  OAI211_X1 U21816 ( .C1(n18471), .C2(n18461), .A(n18575), .B(n18460), .ZN(
        n18462) );
  NAND4_X1 U21817 ( .A1(n18464), .A2(n18463), .A3(n19613), .A4(n18462), .ZN(
        P3_U2660) );
  INV_X1 U21818 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n20149) );
  AOI221_X1 U21819 ( .B1(n18514), .B2(n18578), .C1(n18465), .C2(n18578), .A(
        n18589), .ZN(n18482) );
  AOI21_X1 U21820 ( .B1(n19251), .B2(n18467), .A(n18466), .ZN(n19249) );
  NAND2_X1 U21821 ( .A1(n10451), .A2(n18468), .ZN(n18469) );
  INV_X1 U21822 ( .A(n18469), .ZN(n18485) );
  INV_X1 U21823 ( .A(n19249), .ZN(n18470) );
  AOI221_X1 U21824 ( .B1(n19249), .B2(n18485), .C1(n18470), .C2(n18469), .A(
        n18584), .ZN(n18475) );
  AOI211_X1 U21825 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n18472), .A(n18471), .B(
        n18579), .ZN(n18474) );
  OAI22_X1 U21826 ( .A1(n19251), .A2(n18593), .B1(n18522), .B2(n18751), .ZN(
        n18473) );
  NOR4_X1 U21827 ( .A1(n19556), .A2(n18475), .A3(n18474), .A4(n18473), .ZN(
        n18479) );
  INV_X1 U21828 ( .A(n18476), .ZN(n18490) );
  OAI211_X1 U21829 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(P3_REIP_REG_9__SCAN_IN), 
        .A(n18490), .B(n18477), .ZN(n18478) );
  OAI211_X1 U21830 ( .C1(n20149), .C2(n18482), .A(n18479), .B(n18478), .ZN(
        P3_U2661) );
  NOR2_X1 U21831 ( .A1(n18491), .A2(n18579), .ZN(n18499) );
  AOI22_X1 U21832 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n18481), .B1(
        n18499), .B2(n18480), .ZN(n18494) );
  INV_X1 U21833 ( .A(n18482), .ZN(n18497) );
  AND2_X1 U21834 ( .A1(n18484), .A2(n18483), .ZN(n18486) );
  OAI21_X1 U21835 ( .B1(n18486), .B2(n18487), .A(n18485), .ZN(n18488) );
  AOI221_X1 U21836 ( .B1(n10451), .B2(n18488), .C1(n18487), .C2(n18488), .A(
        n18584), .ZN(n18489) );
  AOI221_X1 U21837 ( .B1(n18497), .B2(P3_REIP_REG_9__SCAN_IN), .C1(n18490), 
        .C2(n14407), .A(n18489), .ZN(n18493) );
  OAI221_X1 U21838 ( .B1(n18596), .B2(n18575), .C1(n18596), .C2(n18491), .A(
        P3_EBX_REG_9__SCAN_IN), .ZN(n18492) );
  NAND4_X1 U21839 ( .A1(n18494), .A2(n18493), .A3(n19603), .A4(n18492), .ZN(
        P3_U2662) );
  AOI21_X1 U21840 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18527), .A(
        n10450), .ZN(n18495) );
  INV_X1 U21841 ( .A(n18495), .ZN(n18509) );
  XOR2_X1 U21842 ( .A(n18509), .B(n18496), .Z(n18505) );
  OAI21_X1 U21843 ( .B1(P3_REIP_REG_8__SCAN_IN), .B2(n18498), .A(n18497), .ZN(
        n18502) );
  INV_X1 U21844 ( .A(n18512), .ZN(n18500) );
  OAI21_X1 U21845 ( .B1(n18500), .B2(n18784), .A(n18499), .ZN(n18501) );
  OAI211_X1 U21846 ( .C1(n18593), .C2(n21933), .A(n18502), .B(n18501), .ZN(
        n18503) );
  AOI211_X1 U21847 ( .C1(n18596), .C2(P3_EBX_REG_8__SCAN_IN), .A(n19556), .B(
        n18503), .ZN(n18504) );
  OAI21_X1 U21848 ( .B1(n20113), .B2(n18505), .A(n18504), .ZN(P3_U2663) );
  AOI21_X1 U21849 ( .B1(n18578), .B2(n18514), .A(n18589), .ZN(n18537) );
  INV_X1 U21850 ( .A(n18537), .ZN(n18530) );
  OAI21_X1 U21851 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18507), .A(
        n18506), .ZN(n19272) );
  NOR3_X1 U21852 ( .A1(n18527), .A2(n10450), .A3(n19272), .ZN(n18508) );
  AOI211_X1 U21853 ( .C1(n19272), .C2(n18509), .A(n18508), .B(n18584), .ZN(
        n18511) );
  INV_X1 U21854 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n19260) );
  OAI22_X1 U21855 ( .A1(n19260), .A2(n18593), .B1(n18522), .B2(n18513), .ZN(
        n18510) );
  AOI211_X1 U21856 ( .C1(n18530), .C2(P3_REIP_REG_7__SCAN_IN), .A(n18511), .B(
        n18510), .ZN(n18518) );
  OAI211_X1 U21857 ( .C1(n18521), .C2(n18513), .A(n18575), .B(n18512), .ZN(
        n18517) );
  NOR2_X1 U21858 ( .A1(n18568), .A2(n18514), .ZN(n18529) );
  OAI211_X1 U21859 ( .C1(P3_REIP_REG_7__SCAN_IN), .C2(P3_REIP_REG_6__SCAN_IN), 
        .A(n18529), .B(n18515), .ZN(n18516) );
  NAND4_X1 U21860 ( .A1(n18518), .A2(n19603), .A3(n18517), .A4(n18516), .ZN(
        P3_U2664) );
  OAI21_X1 U21861 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18535), .A(
        n18519), .ZN(n19281) );
  OAI21_X1 U21862 ( .B1(n18535), .B2(n10450), .A(n18520), .ZN(n18533) );
  AOI211_X1 U21863 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n18540), .A(n18521), .B(
        n18579), .ZN(n18524) );
  OAI22_X1 U21864 ( .A1(n22115), .A2(n18593), .B1(n18522), .B2(n18788), .ZN(
        n18523) );
  NOR3_X1 U21865 ( .A1(n19556), .A2(n18524), .A3(n18523), .ZN(n18532) );
  INV_X1 U21866 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n20142) );
  INV_X1 U21867 ( .A(n19281), .ZN(n18526) );
  NOR3_X1 U21868 ( .A1(n18527), .A2(n18526), .A3(n18525), .ZN(n18528) );
  AOI221_X1 U21869 ( .B1(n18530), .B2(P3_REIP_REG_6__SCAN_IN), .C1(n18529), 
        .C2(n20142), .A(n18528), .ZN(n18531) );
  OAI211_X1 U21870 ( .C1(n19281), .C2(n18533), .A(n18532), .B(n18531), .ZN(
        P3_U2665) );
  INV_X1 U21871 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18544) );
  AND2_X1 U21872 ( .A1(n18578), .A2(n18553), .ZN(n18557) );
  AOI21_X1 U21873 ( .B1(P3_REIP_REG_4__SCAN_IN), .B2(n18557), .A(
        P3_REIP_REG_5__SCAN_IN), .ZN(n18538) );
  NAND2_X1 U21874 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18534), .ZN(
        n18546) );
  AOI21_X1 U21875 ( .B1(n18544), .B2(n18546), .A(n18535), .ZN(n19293) );
  OAI21_X1 U21876 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18546), .A(
        n10451), .ZN(n18547) );
  XOR2_X1 U21877 ( .A(n19293), .B(n18547), .Z(n18536) );
  OAI22_X1 U21878 ( .A1(n18538), .A2(n18537), .B1(n18584), .B2(n18536), .ZN(
        n18539) );
  AOI211_X1 U21879 ( .C1(n18596), .C2(P3_EBX_REG_5__SCAN_IN), .A(n19556), .B(
        n18539), .ZN(n18543) );
  OAI211_X1 U21880 ( .C1(n18550), .C2(n18541), .A(n18575), .B(n18540), .ZN(
        n18542) );
  OAI211_X1 U21881 ( .C1(n18593), .C2(n18544), .A(n18543), .B(n18542), .ZN(
        P3_U2666) );
  NOR2_X1 U21882 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18545), .ZN(
        n19301) );
  NOR2_X1 U21883 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19347), .ZN(
        n18600) );
  NOR2_X1 U21884 ( .A1(n19347), .A2(n18545), .ZN(n18563) );
  OAI21_X1 U21885 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n18563), .A(
        n18546), .ZN(n19308) );
  INV_X1 U21886 ( .A(n19308), .ZN(n18548) );
  OAI221_X1 U21887 ( .B1(n18548), .B2(n18547), .C1(n19308), .C2(n10451), .A(
        n19613), .ZN(n18549) );
  AOI21_X1 U21888 ( .B1(n19301), .B2(n18600), .A(n18549), .ZN(n18560) );
  AOI211_X1 U21889 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n18574), .A(n18550), .B(
        n18579), .ZN(n18551) );
  AOI21_X1 U21890 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n18596), .A(n18551), .ZN(
        n18559) );
  OAI21_X1 U21891 ( .B1(n18553), .B2(n18568), .A(n18552), .ZN(n18573) );
  INV_X1 U21892 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n20139) );
  NOR2_X1 U21893 ( .A1(n18646), .A2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n18555) );
  OAI22_X1 U21894 ( .A1(n18593), .A2(n18554), .B1(n18555), .B2(n18565), .ZN(
        n18556) );
  AOI221_X1 U21895 ( .B1(n18573), .B2(P3_REIP_REG_4__SCAN_IN), .C1(n18557), 
        .C2(n20139), .A(n18556), .ZN(n18558) );
  OAI211_X1 U21896 ( .C1(n18561), .C2(n18560), .A(n18559), .B(n18558), .ZN(
        P3_U2667) );
  INV_X1 U21897 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n19323) );
  AOI21_X1 U21898 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18600), .A(
        n10450), .ZN(n18597) );
  INV_X1 U21899 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18592) );
  NOR2_X1 U21900 ( .A1(n19347), .A2(n18592), .ZN(n18583) );
  INV_X1 U21901 ( .A(n18563), .ZN(n18564) );
  OAI21_X1 U21902 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n18583), .A(
        n18564), .ZN(n19314) );
  XOR2_X1 U21903 ( .A(n18597), .B(n19314), .Z(n18571) );
  INV_X1 U21904 ( .A(n18565), .ZN(n18587) );
  AOI22_X1 U21905 ( .A1(n18596), .A2(P3_EBX_REG_3__SCAN_IN), .B1(n18587), .B2(
        n18566), .ZN(n18570) );
  OR3_X1 U21906 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(n18568), .A3(n18567), .ZN(
        n18569) );
  OAI211_X1 U21907 ( .C1(n18571), .C2(n20113), .A(n18570), .B(n18569), .ZN(
        n18572) );
  AOI21_X1 U21908 ( .B1(P3_REIP_REG_3__SCAN_IN), .B2(n18573), .A(n18572), .ZN(
        n18577) );
  OAI211_X1 U21909 ( .C1(n18580), .C2(n18802), .A(n18575), .B(n18574), .ZN(
        n18576) );
  OAI211_X1 U21910 ( .C1(n18593), .C2(n19323), .A(n18577), .B(n18576), .ZN(
        P3_U2668) );
  NAND2_X1 U21911 ( .A1(n18578), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18603) );
  AOI211_X1 U21912 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n18581), .A(n18580), .B(
        n18579), .ZN(n18595) );
  INV_X1 U21913 ( .A(n18582), .ZN(n18586) );
  AOI21_X1 U21914 ( .B1(n19347), .B2(n18592), .A(n18583), .ZN(n19329) );
  NOR2_X1 U21915 ( .A1(n18584), .A2(n10451), .ZN(n18585) );
  AOI22_X1 U21916 ( .A1(n18587), .A2(n18586), .B1(n19329), .B2(n18585), .ZN(
        n18591) );
  OAI21_X1 U21917 ( .B1(n18589), .B2(n18588), .A(P3_REIP_REG_2__SCAN_IN), .ZN(
        n18590) );
  OAI211_X1 U21918 ( .C1(n18593), .C2(n18592), .A(n18591), .B(n18590), .ZN(
        n18594) );
  AOI211_X1 U21919 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n18596), .A(n18595), .B(
        n18594), .ZN(n18602) );
  INV_X1 U21920 ( .A(n19329), .ZN(n18599) );
  OAI211_X1 U21921 ( .C1(n18600), .C2(n18599), .A(n18598), .B(n18597), .ZN(
        n18601) );
  OAI211_X1 U21922 ( .C1(P3_REIP_REG_2__SCAN_IN), .C2(n18603), .A(n18602), .B(
        n18601), .ZN(P3_U2669) );
  NAND4_X1 U21923 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(P3_EBX_REG_24__SCAN_IN), .A4(n18604), .ZN(n18667) );
  NOR3_X1 U21924 ( .A1(n21874), .A2(n21897), .A3(n18667), .ZN(n18605) );
  NAND4_X1 U21925 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(n18706), .A4(n18605), .ZN(n18609) );
  NAND2_X1 U21926 ( .A1(n18808), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n18608) );
  NAND2_X1 U21927 ( .A1(n18660), .A2(n18606), .ZN(n18607) );
  OAI22_X1 U21928 ( .A1(n18660), .A2(n18608), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n18607), .ZN(P3_U2672) );
  NAND2_X1 U21929 ( .A1(n18610), .A2(n18609), .ZN(n18611) );
  NAND2_X1 U21930 ( .A1(n18611), .A2(n18808), .ZN(n18659) );
  OAI22_X1 U21931 ( .A1(n18614), .A2(n18613), .B1(n14983), .B2(n18612), .ZN(
        n18615) );
  INV_X1 U21932 ( .A(n18615), .ZN(n18623) );
  AOI22_X1 U21933 ( .A1(n18760), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n18616), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18622) );
  AOI22_X1 U21934 ( .A1(n18759), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18692), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n18621) );
  OAI22_X1 U21935 ( .A1(n18715), .A2(n18618), .B1(n18764), .B2(n18617), .ZN(
        n18619) );
  INV_X1 U21936 ( .A(n18619), .ZN(n18620) );
  AND4_X1 U21937 ( .A1(n18623), .A2(n18622), .A3(n18621), .A4(n18620), .ZN(
        n18634) );
  NAND2_X1 U21938 ( .A1(n18624), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n18630) );
  NAND2_X1 U21939 ( .A1(n18646), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n18629) );
  INV_X1 U21940 ( .A(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n18625) );
  OR2_X1 U21941 ( .A1(n18775), .A2(n18625), .ZN(n18628) );
  OR2_X1 U21942 ( .A1(n18773), .A2(n18626), .ZN(n18627) );
  AND4_X1 U21943 ( .A1(n18630), .A2(n18629), .A3(n18628), .A4(n18627), .ZN(
        n18633) );
  AOI22_X1 U21944 ( .A1(n9712), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n14457), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n18632) );
  AOI22_X1 U21945 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n9705), .B1(
        n18652), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n18631) );
  NAND4_X1 U21946 ( .A1(n18634), .A2(n18633), .A3(n18632), .A4(n18631), .ZN(
        n18658) );
  NOR2_X1 U21947 ( .A1(n18835), .A2(n18635), .ZN(n18662) );
  OAI22_X1 U21948 ( .A1(n18763), .A2(n18637), .B1(n14983), .B2(n18636), .ZN(
        n18638) );
  INV_X1 U21949 ( .A(n18638), .ZN(n18645) );
  AOI22_X1 U21950 ( .A1(n18760), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n18616), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18644) );
  AOI22_X1 U21951 ( .A1(n18759), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18692), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n18643) );
  OAI22_X1 U21952 ( .A1(n18715), .A2(n18640), .B1(n18764), .B2(n18639), .ZN(
        n18641) );
  INV_X1 U21953 ( .A(n18641), .ZN(n18642) );
  AND4_X1 U21954 ( .A1(n18645), .A2(n18644), .A3(n18643), .A4(n18642), .ZN(
        n18656) );
  NAND2_X1 U21955 ( .A1(n14951), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n18651) );
  NAND2_X1 U21956 ( .A1(n18646), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n18650) );
  OR2_X1 U21957 ( .A1(n18775), .A2(n14476), .ZN(n18649) );
  OR2_X1 U21958 ( .A1(n18773), .A2(n18647), .ZN(n18648) );
  AND4_X1 U21959 ( .A1(n18651), .A2(n18650), .A3(n18649), .A4(n18648), .ZN(
        n18655) );
  AOI22_X1 U21960 ( .A1(n9712), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14457), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n18654) );
  AOI22_X1 U21961 ( .A1(n9706), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18652), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n18653) );
  NAND4_X1 U21962 ( .A1(n18656), .A2(n18655), .A3(n18654), .A4(n18653), .ZN(
        n18663) );
  NAND2_X1 U21963 ( .A1(n18662), .A2(n18663), .ZN(n18657) );
  XOR2_X1 U21964 ( .A(n18658), .B(n18657), .Z(n18823) );
  OAI22_X1 U21965 ( .A1(n18660), .A2(n18659), .B1(n18823), .B2(n18808), .ZN(
        P3_U2673) );
  NAND2_X1 U21966 ( .A1(n9779), .A2(n18661), .ZN(n18666) );
  XOR2_X1 U21967 ( .A(n18663), .B(n18662), .Z(n18827) );
  AOI22_X1 U21968 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n18664), .B1(n18812), 
        .B2(n18827), .ZN(n18665) );
  OAI21_X1 U21969 ( .B1(n18667), .B2(n18666), .A(n18665), .ZN(P3_U2674) );
  OAI211_X1 U21970 ( .C1(n18837), .C2(n18836), .A(n18812), .B(n18835), .ZN(
        n18668) );
  OAI221_X1 U21971 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n18670), .C1(n18669), 
        .C2(n18674), .A(n18668), .ZN(P3_U2676) );
  INV_X1 U21972 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n18675) );
  AOI21_X1 U21973 ( .B1(n18671), .B2(n18676), .A(n18837), .ZN(n18842) );
  AOI22_X1 U21974 ( .A1(n18842), .A2(n18812), .B1(n18672), .B2(n18675), .ZN(
        n18673) );
  OAI21_X1 U21975 ( .B1(n18675), .B2(n18674), .A(n18673), .ZN(P3_U2677) );
  AOI21_X1 U21976 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n18808), .A(n9865), .ZN(
        n18678) );
  OAI21_X1 U21977 ( .B1(n18679), .B2(n18677), .A(n18676), .ZN(n18850) );
  OAI22_X1 U21978 ( .A1(n18672), .A2(n18678), .B1(n18808), .B2(n18850), .ZN(
        P3_U2678) );
  AOI21_X1 U21979 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n18808), .A(n9779), .ZN(
        n18682) );
  INV_X1 U21980 ( .A(n18679), .ZN(n18680) );
  OAI21_X1 U21981 ( .B1(n18683), .B2(n18681), .A(n18680), .ZN(n18855) );
  OAI22_X1 U21982 ( .A1(n9865), .A2(n18682), .B1(n18808), .B2(n18855), .ZN(
        P3_U2679) );
  AOI21_X1 U21983 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n18808), .A(n9866), .ZN(
        n18687) );
  AOI21_X1 U21984 ( .B1(n18685), .B2(n18684), .A(n18683), .ZN(n18686) );
  INV_X1 U21985 ( .A(n18686), .ZN(n18860) );
  OAI22_X1 U21986 ( .A1(n9779), .A2(n18687), .B1(n18808), .B2(n18860), .ZN(
        P3_U2680) );
  NOR2_X1 U21987 ( .A1(n18754), .A2(n18688), .ZN(n18691) );
  OAI22_X1 U21988 ( .A1(n9704), .A2(n18689), .B1(n17985), .B2(n18794), .ZN(
        n18690) );
  AOI211_X1 U21989 ( .C1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .C2(n9706), .A(
        n18691), .B(n18690), .ZN(n18702) );
  AOI22_X1 U21990 ( .A1(n18759), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n18692), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n18701) );
  AOI22_X1 U21991 ( .A1(n18760), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18616), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n18700) );
  OAI22_X1 U21992 ( .A1(n18763), .A2(n18694), .B1(n14983), .B2(n18693), .ZN(
        n18698) );
  OAI22_X1 U21993 ( .A1(n18715), .A2(n18696), .B1(n18764), .B2(n18695), .ZN(
        n18697) );
  NOR2_X1 U21994 ( .A1(n18698), .A2(n18697), .ZN(n18699) );
  AND4_X1 U21995 ( .A1(n18702), .A2(n18701), .A3(n18700), .A4(n18699), .ZN(
        n18705) );
  AOI22_X1 U21996 ( .A1(n18743), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n18742), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n18704) );
  AOI22_X1 U21997 ( .A1(n14951), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n18646), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n18703) );
  NAND3_X1 U21998 ( .A1(n18705), .A2(n18704), .A3(n18703), .ZN(n18870) );
  OAI21_X1 U21999 ( .B1(n18706), .B2(n21897), .A(n18808), .ZN(n18707) );
  OAI21_X1 U22000 ( .B1(n18808), .B2(n18870), .A(n18707), .ZN(n18708) );
  OAI21_X1 U22001 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n18709), .A(n18708), .ZN(
        P3_U2682) );
  AOI21_X1 U22002 ( .B1(n21981), .B2(n18710), .A(n18812), .ZN(n18711) );
  INV_X1 U22003 ( .A(n18711), .ZN(n18726) );
  AOI22_X1 U22004 ( .A1(n18743), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n18742), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n18713) );
  AOI22_X1 U22005 ( .A1(n14951), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n18646), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18712) );
  NAND2_X1 U22006 ( .A1(n18713), .A2(n18712), .ZN(n18725) );
  INV_X1 U22007 ( .A(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n18772) );
  INV_X1 U22008 ( .A(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n18774) );
  OAI22_X1 U22009 ( .A1(n9704), .A2(n18772), .B1(n18755), .B2(n18774), .ZN(
        n18724) );
  OAI22_X1 U22010 ( .A1(n19819), .A2(n18754), .B1(n17985), .B2(n12035), .ZN(
        n18723) );
  OAI22_X1 U22011 ( .A1(n18763), .A2(n18761), .B1(n18715), .B2(n18714), .ZN(
        n18716) );
  INV_X1 U22012 ( .A(n18716), .ZN(n18721) );
  AOI22_X1 U22013 ( .A1(n18760), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n18717), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18720) );
  AOI22_X1 U22014 ( .A1(n14112), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18616), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n18719) );
  AOI22_X1 U22015 ( .A1(n18759), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12013), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n18718) );
  NAND4_X1 U22016 ( .A1(n18721), .A2(n18720), .A3(n18719), .A4(n18718), .ZN(
        n18722) );
  NOR4_X1 U22017 ( .A1(n18725), .A2(n18724), .A3(n18723), .A4(n18722), .ZN(
        n18884) );
  OAI22_X1 U22018 ( .A1(n18727), .A2(n18726), .B1(n18884), .B2(n18808), .ZN(
        P3_U2687) );
  OAI22_X1 U22019 ( .A1(n9704), .A2(n18728), .B1(n17985), .B2(n14969), .ZN(
        n18732) );
  OAI22_X1 U22020 ( .A1(n18755), .A2(n18730), .B1(n18754), .B2(n18729), .ZN(
        n18731) );
  NOR2_X1 U22021 ( .A1(n18732), .A2(n18731), .ZN(n18741) );
  AOI22_X1 U22022 ( .A1(n18759), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12013), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n18740) );
  AOI22_X1 U22023 ( .A1(n18760), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18616), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n18739) );
  OAI22_X1 U22024 ( .A1(n18763), .A2(n18734), .B1(n14983), .B2(n18733), .ZN(
        n18737) );
  OAI22_X1 U22025 ( .A1(n18715), .A2(n21988), .B1(n18764), .B2(n18735), .ZN(
        n18736) );
  NOR2_X1 U22026 ( .A1(n18737), .A2(n18736), .ZN(n18738) );
  AND4_X1 U22027 ( .A1(n18741), .A2(n18740), .A3(n18739), .A4(n18738), .ZN(
        n18746) );
  AOI22_X1 U22028 ( .A1(n18743), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n18742), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18745) );
  AOI22_X1 U22029 ( .A1(n14951), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n18646), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n18744) );
  NAND3_X1 U22030 ( .A1(n18746), .A2(n18745), .A3(n18744), .ZN(n18894) );
  NOR3_X1 U22031 ( .A1(n18747), .A2(P3_EBX_REG_10__SCAN_IN), .A3(n19654), .ZN(
        n18748) );
  AOI21_X1 U22032 ( .B1(n18812), .B2(n18894), .A(n18748), .ZN(n18749) );
  OAI21_X1 U22033 ( .B1(n18751), .B2(n18750), .A(n18749), .ZN(P3_U2693) );
  NAND2_X1 U22034 ( .A1(n18808), .A2(n18781), .ZN(n18786) );
  OAI22_X1 U22035 ( .A1(n9704), .A2(n18752), .B1(n17985), .B2(n21925), .ZN(
        n18758) );
  OAI22_X1 U22036 ( .A1(n18756), .A2(n18755), .B1(n18754), .B2(n18753), .ZN(
        n18757) );
  NOR2_X1 U22037 ( .A1(n18758), .A2(n18757), .ZN(n18771) );
  AOI22_X1 U22038 ( .A1(n18759), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12013), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n18770) );
  AOI22_X1 U22039 ( .A1(n18760), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17631), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n18769) );
  OAI22_X1 U22040 ( .A1(n18763), .A2(n18762), .B1(n14983), .B2(n18761), .ZN(
        n18767) );
  OAI22_X1 U22041 ( .A1(n18715), .A2(n18765), .B1(n18764), .B2(n19819), .ZN(
        n18766) );
  NOR2_X1 U22042 ( .A1(n18767), .A2(n18766), .ZN(n18768) );
  NAND4_X1 U22043 ( .A1(n18771), .A2(n18770), .A3(n18769), .A4(n18768), .ZN(
        n18780) );
  OAI22_X1 U22044 ( .A1(n18775), .A2(n18774), .B1(n18773), .B2(n18772), .ZN(
        n18779) );
  OAI22_X1 U22045 ( .A1(n12035), .A2(n13862), .B1(n18777), .B2(n18776), .ZN(
        n18778) );
  OR3_X1 U22046 ( .A1(n18780), .A2(n18779), .A3(n18778), .ZN(n18899) );
  NOR3_X1 U22047 ( .A1(n18781), .A2(P3_EBX_REG_8__SCAN_IN), .A3(n19654), .ZN(
        n18782) );
  AOI21_X1 U22048 ( .B1(n18812), .B2(n18899), .A(n18782), .ZN(n18783) );
  OAI21_X1 U22049 ( .B1(n18784), .B2(n18786), .A(n18783), .ZN(P3_U2695) );
  NOR2_X1 U22050 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n9891), .ZN(n18787) );
  OAI22_X1 U22051 ( .A1(n18787), .A2(n18786), .B1(n18785), .B2(n18808), .ZN(
        P3_U2696) );
  AOI21_X1 U22052 ( .B1(n18788), .B2(n18792), .A(n18812), .ZN(n18789) );
  INV_X1 U22053 ( .A(n18789), .ZN(n18791) );
  OAI22_X1 U22054 ( .A1(n9891), .A2(n18791), .B1(n18790), .B2(n18808), .ZN(
        P3_U2697) );
  OAI21_X1 U22055 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n18798), .A(n18792), .ZN(
        n18793) );
  AOI22_X1 U22056 ( .A1(n18812), .A2(n18794), .B1(n18793), .B2(n18808), .ZN(
        P3_U2698) );
  AOI21_X1 U22057 ( .B1(n22097), .B2(n18795), .A(n18812), .ZN(n18796) );
  INV_X1 U22058 ( .A(n18796), .ZN(n18797) );
  OAI22_X1 U22059 ( .A1(n18798), .A2(n18797), .B1(n11975), .B2(n18808), .ZN(
        P3_U2699) );
  NOR2_X1 U22060 ( .A1(n18799), .A2(n18812), .ZN(n18804) );
  INV_X1 U22061 ( .A(n18799), .ZN(n18800) );
  OAI21_X1 U22062 ( .B1(n18800), .B2(n19654), .A(n18802), .ZN(n18801) );
  OAI21_X1 U22063 ( .B1(n18804), .B2(n18802), .A(n18801), .ZN(n18803) );
  OAI21_X1 U22064 ( .B1(n11994), .B2(n18808), .A(n18803), .ZN(P3_U2700) );
  OAI21_X1 U22065 ( .B1(P3_EBX_REG_2__SCAN_IN), .B2(n18805), .A(n18804), .ZN(
        n18806) );
  OAI21_X1 U22066 ( .B1(n18808), .B2(n18807), .A(n18806), .ZN(P3_U2701) );
  OAI222_X1 U22067 ( .A1(n18811), .A2(n18816), .B1(n18810), .B2(n18814), .C1(
        n18809), .C2(n18808), .ZN(P3_U2702) );
  NAND2_X1 U22068 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18812), .ZN(
        n18813) );
  OAI221_X1 U22069 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n18816), .C1(n18815), 
        .C2(n18814), .A(n18813), .ZN(P3_U2703) );
  INV_X1 U22070 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n18993) );
  INV_X1 U22071 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n18925) );
  INV_X1 U22072 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n18931) );
  NAND4_X1 U22073 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_21__SCAN_IN), 
        .A3(P3_EAX_REG_19__SCAN_IN), .A4(n18817), .ZN(n18862) );
  NAND2_X1 U22074 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n18852), .ZN(n18851) );
  NAND2_X1 U22075 ( .A1(n18824), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n18820) );
  OAI22_X1 U22076 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n18863), .B1(n18907), 
        .B2(n18824), .ZN(n18818) );
  AOI22_X1 U22077 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n18877), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n18818), .ZN(n18819) );
  OAI21_X1 U22078 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n18820), .A(n18819), .ZN(
        P3_U2704) );
  AOI22_X1 U22079 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18878), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n18877), .ZN(n18822) );
  OAI211_X1 U22080 ( .C1(n18824), .C2(P3_EAX_REG_30__SCAN_IN), .A(n18902), .B(
        n18820), .ZN(n18821) );
  OAI211_X1 U22081 ( .C1(n18823), .C2(n18883), .A(n18822), .B(n18821), .ZN(
        P3_U2705) );
  INV_X1 U22082 ( .A(n18824), .ZN(n18826) );
  OAI21_X1 U22083 ( .B1(n18907), .B2(n18993), .A(n18831), .ZN(n18825) );
  AOI22_X1 U22084 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18877), .B1(n18826), .B2(
        n18825), .ZN(n18829) );
  AOI22_X1 U22085 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18878), .B1(n18827), .B2(
        n18911), .ZN(n18828) );
  NAND2_X1 U22086 ( .A1(n18829), .A2(n18828), .ZN(P3_U2706) );
  AOI22_X1 U22087 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n18878), .B1(n18830), .B2(
        n18911), .ZN(n18834) );
  OAI211_X1 U22088 ( .C1(n18832), .C2(P3_EAX_REG_28__SCAN_IN), .A(n18902), .B(
        n18831), .ZN(n18833) );
  OAI211_X1 U22089 ( .C1(n18864), .C2(n16857), .A(n18834), .B(n18833), .ZN(
        P3_U2707) );
  OAI21_X1 U22090 ( .B1(n18837), .B2(n18836), .A(n18835), .ZN(n18841) );
  AOI22_X1 U22091 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18878), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n18877), .ZN(n18840) );
  OAI211_X1 U22092 ( .C1(n9867), .C2(P3_EAX_REG_27__SCAN_IN), .A(n18902), .B(
        n18838), .ZN(n18839) );
  OAI211_X1 U22093 ( .C1(n18883), .C2(n18841), .A(n18840), .B(n18839), .ZN(
        P3_U2708) );
  INV_X1 U22094 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n19009) );
  AOI22_X1 U22095 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18877), .B1(n18842), .B2(
        n18911), .ZN(n18845) );
  AOI211_X1 U22096 ( .C1(n18925), .C2(n18846), .A(n9867), .B(n18907), .ZN(
        n18843) );
  INV_X1 U22097 ( .A(n18843), .ZN(n18844) );
  OAI211_X1 U22098 ( .C1(n18872), .C2(n19009), .A(n18845), .B(n18844), .ZN(
        P3_U2709) );
  AOI22_X1 U22099 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18878), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n18877), .ZN(n18849) );
  OAI211_X1 U22100 ( .C1(n18847), .C2(P3_EAX_REG_25__SCAN_IN), .A(n18902), .B(
        n18846), .ZN(n18848) );
  OAI211_X1 U22101 ( .C1(n18883), .C2(n18850), .A(n18849), .B(n18848), .ZN(
        P3_U2710) );
  AOI22_X1 U22102 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18878), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n18877), .ZN(n18854) );
  OAI211_X1 U22103 ( .C1(n18852), .C2(P3_EAX_REG_24__SCAN_IN), .A(n18902), .B(
        n18851), .ZN(n18853) );
  OAI211_X1 U22104 ( .C1(n18883), .C2(n18855), .A(n18854), .B(n18853), .ZN(
        P3_U2711) );
  AOI22_X1 U22105 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18878), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n18877), .ZN(n18859) );
  OAI211_X1 U22106 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n18857), .A(n18902), .B(
        n18856), .ZN(n18858) );
  OAI211_X1 U22107 ( .C1(n18883), .C2(n18860), .A(n18859), .B(n18858), .ZN(
        P3_U2712) );
  NOR2_X1 U22108 ( .A1(n18862), .A2(n18861), .ZN(n18868) );
  NAND2_X1 U22109 ( .A1(n18902), .A2(n18876), .ZN(n18871) );
  OAI21_X1 U22110 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n18863), .A(n18871), .ZN(
        n18867) );
  OAI22_X1 U22111 ( .A1(n18865), .A2(n18883), .B1(n18864), .B2(n16904), .ZN(
        n18866) );
  AOI221_X1 U22112 ( .B1(n18868), .B2(n18931), .C1(n18867), .C2(
        P3_EAX_REG_22__SCAN_IN), .A(n18866), .ZN(n18869) );
  OAI21_X1 U22113 ( .B1(n19649), .B2(n18872), .A(n18869), .ZN(P3_U2713) );
  AOI22_X1 U22114 ( .A1(n18877), .A2(BUF2_REG_21__SCAN_IN), .B1(n18911), .B2(
        n18870), .ZN(n18875) );
  INV_X1 U22115 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n18933) );
  OAI22_X1 U22116 ( .A1(n19645), .A2(n18872), .B1(n18933), .B2(n18871), .ZN(
        n18873) );
  INV_X1 U22117 ( .A(n18873), .ZN(n18874) );
  OAI211_X1 U22118 ( .C1(P3_EAX_REG_21__SCAN_IN), .C2(n18876), .A(n18875), .B(
        n18874), .ZN(P3_U2714) );
  AOI22_X1 U22119 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n18878), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n18877), .ZN(n18882) );
  OAI211_X1 U22120 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n18880), .A(n18902), .B(
        n18879), .ZN(n18881) );
  OAI211_X1 U22121 ( .C1(n18884), .C2(n18883), .A(n18882), .B(n18881), .ZN(
        P3_U2719) );
  NAND2_X1 U22122 ( .A1(n18885), .A2(n18896), .ZN(n18889) );
  AOI22_X1 U22123 ( .A1(n18900), .A2(BUF2_REG_15__SCAN_IN), .B1(n18911), .B2(
        n18886), .ZN(n18887) );
  OAI221_X1 U22124 ( .B1(P3_EAX_REG_15__SCAN_IN), .B2(n18889), .C1(n19023), 
        .C2(n18888), .A(n18887), .ZN(P3_U2720) );
  NAND2_X1 U22125 ( .A1(n18893), .A2(P3_EAX_REG_13__SCAN_IN), .ZN(n18892) );
  AOI22_X1 U22126 ( .A1(n18900), .A2(BUF2_REG_13__SCAN_IN), .B1(n18911), .B2(
        n18890), .ZN(n18891) );
  OAI221_X1 U22127 ( .B1(n18893), .B2(P3_EAX_REG_13__SCAN_IN), .C1(n18892), 
        .C2(n18907), .A(n18891), .ZN(P3_U2722) );
  AOI22_X1 U22128 ( .A1(n18900), .A2(BUF2_REG_10__SCAN_IN), .B1(n18911), .B2(
        n18894), .ZN(n18898) );
  OAI211_X1 U22129 ( .C1(P3_EAX_REG_10__SCAN_IN), .C2(n18896), .A(n18902), .B(
        n18895), .ZN(n18897) );
  NAND2_X1 U22130 ( .A1(n18898), .A2(n18897), .ZN(P3_U2725) );
  AOI22_X1 U22131 ( .A1(n18900), .A2(BUF2_REG_8__SCAN_IN), .B1(n18911), .B2(
        n18899), .ZN(n18905) );
  OAI211_X1 U22132 ( .C1(P3_EAX_REG_8__SCAN_IN), .C2(n18903), .A(n18902), .B(
        n18901), .ZN(n18904) );
  NAND2_X1 U22133 ( .A1(n18905), .A2(n18904), .ZN(P3_U2727) );
  INV_X1 U22134 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n19641) );
  AOI211_X1 U22135 ( .C1(n18908), .C2(n18963), .A(n18907), .B(n18906), .ZN(
        n18909) );
  AOI21_X1 U22136 ( .B1(n18911), .B2(n18910), .A(n18909), .ZN(n18912) );
  OAI21_X1 U22137 ( .B1(n19641), .B2(n18913), .A(n18912), .ZN(P3_U2731) );
  NOR2_X2 U22138 ( .A1(n18914), .A2(n19214), .ZN(n20214) );
  INV_X1 U22139 ( .A(n18976), .ZN(n18916) );
  NOR2_X4 U22140 ( .A1(n20214), .A2(n18918), .ZN(n18961) );
  AND2_X1 U22141 ( .A1(n18961), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U22142 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n18995) );
  NAND2_X1 U22143 ( .A1(n18918), .A2(n18917), .ZN(n18942) );
  AOI22_X1 U22144 ( .A1(n20214), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n18961), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18919) );
  OAI21_X1 U22145 ( .B1(n18995), .B2(n18942), .A(n18919), .ZN(P3_U2737) );
  AOI22_X1 U22146 ( .A1(P3_DATAO_REG_29__SCAN_IN), .A2(n18961), .B1(n20214), 
        .B2(P3_UWORD_REG_13__SCAN_IN), .ZN(n18920) );
  OAI21_X1 U22147 ( .B1(n18993), .B2(n18942), .A(n18920), .ZN(P3_U2738) );
  INV_X1 U22148 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n18922) );
  AOI22_X1 U22149 ( .A1(n20214), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18961), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18921) );
  OAI21_X1 U22150 ( .B1(n18922), .B2(n18942), .A(n18921), .ZN(P3_U2739) );
  AOI22_X1 U22151 ( .A1(n20214), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n18961), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18923) );
  OAI21_X1 U22152 ( .B1(n10266), .B2(n18942), .A(n18923), .ZN(P3_U2740) );
  AOI22_X1 U22153 ( .A1(n20214), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n18961), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18924) );
  OAI21_X1 U22154 ( .B1(n18925), .B2(n18942), .A(n18924), .ZN(P3_U2741) );
  CLKBUF_X1 U22155 ( .A(n20214), .Z(n18967) );
  AOI22_X1 U22156 ( .A1(n18967), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18961), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18926) );
  OAI21_X1 U22157 ( .B1(n10265), .B2(n18942), .A(n18926), .ZN(P3_U2742) );
  INV_X1 U22158 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n18987) );
  AOI22_X1 U22159 ( .A1(n18967), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n18961), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18927) );
  OAI21_X1 U22160 ( .B1(n18987), .B2(n18942), .A(n18927), .ZN(P3_U2743) );
  INV_X1 U22161 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n18929) );
  AOI22_X1 U22162 ( .A1(n18967), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n18961), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18928) );
  OAI21_X1 U22163 ( .B1(n18929), .B2(n18942), .A(n18928), .ZN(P3_U2744) );
  AOI22_X1 U22164 ( .A1(n18967), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18961), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18930) );
  OAI21_X1 U22165 ( .B1(n18931), .B2(n18942), .A(n18930), .ZN(P3_U2745) );
  AOI22_X1 U22166 ( .A1(n18967), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n18961), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18932) );
  OAI21_X1 U22167 ( .B1(n18933), .B2(n18942), .A(n18932), .ZN(P3_U2746) );
  INV_X1 U22168 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n22101) );
  AOI22_X1 U22169 ( .A1(n18967), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18961), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18934) );
  OAI21_X1 U22170 ( .B1(n22101), .B2(n18942), .A(n18934), .ZN(P3_U2747) );
  INV_X1 U22171 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n18936) );
  AOI22_X1 U22172 ( .A1(n18967), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n18961), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18935) );
  OAI21_X1 U22173 ( .B1(n18936), .B2(n18942), .A(n18935), .ZN(P3_U2748) );
  AOI22_X1 U22174 ( .A1(n18967), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n18961), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18937) );
  OAI21_X1 U22175 ( .B1(n18938), .B2(n18942), .A(n18937), .ZN(P3_U2749) );
  AOI22_X1 U22176 ( .A1(n18967), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n18961), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18939) );
  OAI21_X1 U22177 ( .B1(n18940), .B2(n18942), .A(n18939), .ZN(P3_U2750) );
  INV_X1 U22178 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n18943) );
  AOI22_X1 U22179 ( .A1(n18967), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n18961), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18941) );
  OAI21_X1 U22180 ( .B1(n18943), .B2(n18942), .A(n18941), .ZN(P3_U2751) );
  AOI22_X1 U22181 ( .A1(n18967), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n18961), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18944) );
  OAI21_X1 U22182 ( .B1(n19023), .B2(n18971), .A(n18944), .ZN(P3_U2752) );
  AOI22_X1 U22183 ( .A1(n18967), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n18961), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18945) );
  OAI21_X1 U22184 ( .B1(n19018), .B2(n18971), .A(n18945), .ZN(P3_U2753) );
  INV_X1 U22185 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n19016) );
  AOI22_X1 U22186 ( .A1(n18967), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n18961), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18946) );
  OAI21_X1 U22187 ( .B1(n19016), .B2(n18971), .A(n18946), .ZN(P3_U2754) );
  INV_X1 U22188 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n21918) );
  AOI22_X1 U22189 ( .A1(n18967), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n18961), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18947) );
  OAI21_X1 U22190 ( .B1(n21918), .B2(n18971), .A(n18947), .ZN(P3_U2755) );
  AOI22_X1 U22191 ( .A1(n18967), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18961), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18948) );
  OAI21_X1 U22192 ( .B1(n18949), .B2(n18971), .A(n18948), .ZN(P3_U2756) );
  AOI22_X1 U22193 ( .A1(n18967), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18961), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18950) );
  OAI21_X1 U22194 ( .B1(n18951), .B2(n18971), .A(n18950), .ZN(P3_U2757) );
  AOI22_X1 U22195 ( .A1(n18967), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n18961), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18952) );
  OAI21_X1 U22196 ( .B1(n18953), .B2(n18971), .A(n18952), .ZN(P3_U2758) );
  INV_X1 U22197 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n19005) );
  AOI22_X1 U22198 ( .A1(n18967), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18961), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18954) );
  OAI21_X1 U22199 ( .B1(n19005), .B2(n18971), .A(n18954), .ZN(P3_U2759) );
  INV_X1 U22200 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n18956) );
  AOI22_X1 U22201 ( .A1(n18967), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n18961), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18955) );
  OAI21_X1 U22202 ( .B1(n18956), .B2(n18971), .A(n18955), .ZN(P3_U2760) );
  AOI22_X1 U22203 ( .A1(P3_DATAO_REG_6__SCAN_IN), .A2(n18961), .B1(n20214), 
        .B2(P3_LWORD_REG_6__SCAN_IN), .ZN(n18957) );
  OAI21_X1 U22204 ( .B1(n18958), .B2(n18971), .A(n18957), .ZN(P3_U2761) );
  INV_X1 U22205 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n18960) );
  AOI22_X1 U22206 ( .A1(n18967), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18961), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18959) );
  OAI21_X1 U22207 ( .B1(n18960), .B2(n18971), .A(n18959), .ZN(P3_U2762) );
  AOI22_X1 U22208 ( .A1(n18967), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18961), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18962) );
  OAI21_X1 U22209 ( .B1(n18963), .B2(n18971), .A(n18962), .ZN(P3_U2763) );
  INV_X1 U22210 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n18965) );
  AOI22_X1 U22211 ( .A1(n18967), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n18961), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18964) );
  OAI21_X1 U22212 ( .B1(n18965), .B2(n18971), .A(n18964), .ZN(P3_U2764) );
  INV_X1 U22213 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n22061) );
  AOI22_X1 U22214 ( .A1(n18967), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n18961), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18966) );
  OAI21_X1 U22215 ( .B1(n22061), .B2(n18971), .A(n18966), .ZN(P3_U2765) );
  AOI22_X1 U22216 ( .A1(n18967), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n18961), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18968) );
  OAI21_X1 U22217 ( .B1(n18969), .B2(n18971), .A(n18968), .ZN(P3_U2766) );
  AOI22_X1 U22218 ( .A1(P3_DATAO_REG_0__SCAN_IN), .A2(n18961), .B1(n20214), 
        .B2(P3_LWORD_REG_0__SCAN_IN), .ZN(n18970) );
  OAI21_X1 U22219 ( .B1(n18972), .B2(n18971), .A(n18970), .ZN(P3_U2767) );
  INV_X1 U22220 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n19624) );
  AOI21_X1 U22221 ( .B1(n18973), .B2(n20121), .A(n18976), .ZN(n18974) );
  NAND2_X2 U22222 ( .A1(n18975), .A2(n18974), .ZN(n19019) );
  OR2_X1 U22223 ( .A1(n19019), .A2(n20217), .ZN(n18985) );
  AOI22_X1 U22224 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n19012), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n19019), .ZN(n18977) );
  OAI21_X1 U22225 ( .B1(n19624), .B2(n18985), .A(n18977), .ZN(P3_U2768) );
  AOI22_X1 U22226 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n19012), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n19019), .ZN(n18978) );
  OAI21_X1 U22227 ( .B1(n21987), .B2(n18985), .A(n18978), .ZN(P3_U2769) );
  AOI22_X1 U22228 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n19012), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n19019), .ZN(n18979) );
  OAI21_X1 U22229 ( .B1(n19633), .B2(n18985), .A(n18979), .ZN(P3_U2770) );
  AOI22_X1 U22230 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n19012), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n19019), .ZN(n18980) );
  OAI21_X1 U22231 ( .B1(n19637), .B2(n18985), .A(n18980), .ZN(P3_U2771) );
  AOI22_X1 U22232 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n19012), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n19019), .ZN(n18981) );
  OAI21_X1 U22233 ( .B1(n19641), .B2(n18985), .A(n18981), .ZN(P3_U2772) );
  AOI22_X1 U22234 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n19012), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n19019), .ZN(n18982) );
  OAI21_X1 U22235 ( .B1(n19645), .B2(n18985), .A(n18982), .ZN(P3_U2773) );
  AOI22_X1 U22236 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n19012), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n19019), .ZN(n18983) );
  OAI21_X1 U22237 ( .B1(n19649), .B2(n18985), .A(n18983), .ZN(P3_U2774) );
  AOI22_X1 U22238 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n19012), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n19019), .ZN(n18984) );
  OAI21_X1 U22239 ( .B1(n21919), .B2(n18985), .A(n18984), .ZN(P3_U2775) );
  INV_X1 U22240 ( .A(n18985), .ZN(n19020) );
  AOI22_X1 U22241 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n19020), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n19019), .ZN(n18986) );
  OAI21_X1 U22242 ( .B1(n18987), .B2(n19022), .A(n18986), .ZN(P3_U2776) );
  AOI22_X1 U22243 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n19012), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n19019), .ZN(n18988) );
  OAI21_X1 U22244 ( .B1(n19007), .B2(n18985), .A(n18988), .ZN(P3_U2777) );
  AOI22_X1 U22245 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n19012), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n19019), .ZN(n18989) );
  OAI21_X1 U22246 ( .B1(n19009), .B2(n18985), .A(n18989), .ZN(P3_U2778) );
  AOI22_X1 U22247 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n19012), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n19019), .ZN(n18990) );
  OAI21_X1 U22248 ( .B1(n19011), .B2(n18985), .A(n18990), .ZN(P3_U2779) );
  AOI22_X1 U22249 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n19012), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n19019), .ZN(n18991) );
  OAI21_X1 U22250 ( .B1(n19014), .B2(n18985), .A(n18991), .ZN(P3_U2780) );
  AOI22_X1 U22251 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n19020), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n19019), .ZN(n18992) );
  OAI21_X1 U22252 ( .B1(n18993), .B2(n19022), .A(n18992), .ZN(P3_U2781) );
  AOI22_X1 U22253 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n19020), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n19019), .ZN(n18994) );
  OAI21_X1 U22254 ( .B1(n18995), .B2(n19022), .A(n18994), .ZN(P3_U2782) );
  AOI22_X1 U22255 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n19012), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n19019), .ZN(n18996) );
  OAI21_X1 U22256 ( .B1(n19624), .B2(n18985), .A(n18996), .ZN(P3_U2783) );
  AOI22_X1 U22257 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n19012), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n19019), .ZN(n18997) );
  OAI21_X1 U22258 ( .B1(n21987), .B2(n18985), .A(n18997), .ZN(P3_U2784) );
  AOI22_X1 U22259 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n19012), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n19019), .ZN(n18998) );
  OAI21_X1 U22260 ( .B1(n19633), .B2(n18985), .A(n18998), .ZN(P3_U2785) );
  AOI22_X1 U22261 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n19012), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n19019), .ZN(n18999) );
  OAI21_X1 U22262 ( .B1(n19637), .B2(n18985), .A(n18999), .ZN(P3_U2786) );
  AOI22_X1 U22263 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n19012), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n19019), .ZN(n19000) );
  OAI21_X1 U22264 ( .B1(n19641), .B2(n18985), .A(n19000), .ZN(P3_U2787) );
  AOI22_X1 U22265 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n19012), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n19019), .ZN(n19001) );
  OAI21_X1 U22266 ( .B1(n19645), .B2(n18985), .A(n19001), .ZN(P3_U2788) );
  AOI22_X1 U22267 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n19012), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n19019), .ZN(n19002) );
  OAI21_X1 U22268 ( .B1(n19649), .B2(n18985), .A(n19002), .ZN(P3_U2789) );
  AOI22_X1 U22269 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n19012), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n19019), .ZN(n19003) );
  OAI21_X1 U22270 ( .B1(n21919), .B2(n18985), .A(n19003), .ZN(P3_U2790) );
  AOI22_X1 U22271 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n19020), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n19019), .ZN(n19004) );
  OAI21_X1 U22272 ( .B1(n19005), .B2(n19022), .A(n19004), .ZN(P3_U2791) );
  AOI22_X1 U22273 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n19012), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n19019), .ZN(n19006) );
  OAI21_X1 U22274 ( .B1(n19007), .B2(n18985), .A(n19006), .ZN(P3_U2792) );
  AOI22_X1 U22275 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n19012), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n19019), .ZN(n19008) );
  OAI21_X1 U22276 ( .B1(n19009), .B2(n18985), .A(n19008), .ZN(P3_U2793) );
  AOI22_X1 U22277 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n19012), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n19019), .ZN(n19010) );
  OAI21_X1 U22278 ( .B1(n19011), .B2(n18985), .A(n19010), .ZN(P3_U2794) );
  AOI22_X1 U22279 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n19012), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n19019), .ZN(n19013) );
  OAI21_X1 U22280 ( .B1(n19014), .B2(n18985), .A(n19013), .ZN(P3_U2795) );
  AOI22_X1 U22281 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n19020), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n19019), .ZN(n19015) );
  OAI21_X1 U22282 ( .B1(n19016), .B2(n19022), .A(n19015), .ZN(P3_U2796) );
  AOI22_X1 U22283 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n19020), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n19019), .ZN(n19017) );
  OAI21_X1 U22284 ( .B1(n19018), .B2(n19022), .A(n19017), .ZN(P3_U2797) );
  AOI22_X1 U22285 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n19020), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n19019), .ZN(n19021) );
  OAI21_X1 U22286 ( .B1(n19023), .B2(n19022), .A(n19021), .ZN(P3_U2798) );
  INV_X1 U22287 ( .A(n19024), .ZN(n19025) );
  AOI22_X1 U22288 ( .A1(n19556), .A2(P3_REIP_REG_27__SCAN_IN), .B1(n19236), 
        .B2(n19028), .ZN(n19029) );
  OAI221_X1 U22289 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n19032), .C1(
        n19031), .C2(n19030), .A(n19029), .ZN(n19033) );
  AOI221_X1 U22290 ( .B1(n19035), .B2(n19034), .C1(n19046), .C2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n19033), .ZN(n19036) );
  OAI21_X1 U22291 ( .B1(n19362), .B2(n19204), .A(n19036), .ZN(P3_U2803) );
  NAND3_X1 U22292 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n19037), .A3(
        n22049), .ZN(n19364) );
  OAI21_X1 U22293 ( .B1(n19863), .B2(n19039), .A(n19038), .ZN(n19043) );
  AOI21_X1 U22294 ( .B1(n19183), .B2(n19082), .A(n19040), .ZN(n19042) );
  NAND2_X1 U22295 ( .A1(n19556), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n19368) );
  INV_X1 U22296 ( .A(n19368), .ZN(n19041) );
  AOI211_X1 U22297 ( .C1(n19044), .C2(n19043), .A(n19042), .B(n19041), .ZN(
        n19048) );
  XNOR2_X1 U22298 ( .A(n19045), .B(n22049), .ZN(n19366) );
  AOI22_X1 U22299 ( .A1(n19046), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B1(
        n19254), .B2(n19366), .ZN(n19047) );
  OAI211_X1 U22300 ( .C1(n19091), .C2(n19364), .A(n19048), .B(n19047), .ZN(
        P3_U2804) );
  XOR2_X1 U22301 ( .A(n19050), .B(n19049), .Z(n19380) );
  NOR2_X1 U22302 ( .A1(n19613), .A2(n20176), .ZN(n19375) );
  NAND2_X1 U22303 ( .A1(n19142), .A2(n19051), .ZN(n19052) );
  OAI211_X1 U22304 ( .C1(n17782), .C2(n19863), .A(n19313), .B(n19052), .ZN(
        n19084) );
  AOI21_X1 U22305 ( .B1(n19123), .B2(n19053), .A(n19084), .ZN(n19067) );
  NAND2_X1 U22306 ( .A1(n17782), .A2(n19212), .ZN(n19069) );
  OAI21_X1 U22307 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n19054), .ZN(n19055) );
  OAI22_X1 U22308 ( .A1(n19067), .A2(n19056), .B1(n19069), .B2(n19055), .ZN(
        n19057) );
  AOI211_X1 U22309 ( .C1(n19058), .C2(n19236), .A(n19375), .B(n19057), .ZN(
        n19063) );
  XOR2_X1 U22310 ( .A(n19059), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n19377) );
  NAND2_X1 U22311 ( .A1(n9859), .A2(n19060), .ZN(n19061) );
  XNOR2_X1 U22312 ( .A(n19061), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n19376) );
  AOI22_X1 U22313 ( .A1(n19340), .A2(n19377), .B1(n19254), .B2(n19376), .ZN(
        n19062) );
  OAI211_X1 U22314 ( .C1(n19208), .C2(n19380), .A(n19063), .B(n19062), .ZN(
        P3_U2805) );
  AOI22_X1 U22315 ( .A1(n19340), .A2(n19384), .B1(n19065), .B2(n19064), .ZN(
        n19090) );
  NAND2_X1 U22316 ( .A1(n19556), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n19066) );
  OAI221_X1 U22317 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n19069), .C1(
        n19068), .C2(n19067), .A(n19066), .ZN(n19075) );
  INV_X1 U22318 ( .A(n19070), .ZN(n19071) );
  AOI21_X1 U22319 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n19072), .A(
        n19071), .ZN(n19381) );
  NAND2_X1 U22320 ( .A1(n19073), .A2(n19078), .ZN(n19392) );
  OAI22_X1 U22321 ( .A1(n19381), .A2(n19204), .B1(n19187), .B2(n19392), .ZN(
        n19074) );
  AOI211_X1 U22322 ( .C1(n19236), .C2(n19076), .A(n19075), .B(n19074), .ZN(
        n19077) );
  OAI21_X1 U22323 ( .B1(n19090), .B2(n19078), .A(n19077), .ZN(P3_U2806) );
  INV_X1 U22324 ( .A(n19132), .ZN(n19104) );
  AOI21_X1 U22325 ( .B1(n19160), .B2(n19079), .A(n19101), .ZN(n19080) );
  AOI211_X1 U22326 ( .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n19196), .A(
        n19104), .B(n19080), .ZN(n19081) );
  XNOR2_X1 U22327 ( .A(n19081), .B(n19394), .ZN(n19398) );
  OAI21_X1 U22328 ( .B1(n19236), .B2(n19123), .A(n19083), .ZN(n19087) );
  INV_X1 U22329 ( .A(n11875), .ZN(n19085) );
  OAI221_X1 U22330 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n19085), .C1(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .C2(n20002), .A(n19084), .ZN(
        n19086) );
  OAI211_X1 U22331 ( .C1(n20173), .C2(n19613), .A(n19087), .B(n19086), .ZN(
        n19088) );
  AOI21_X1 U22332 ( .B1(n19254), .B2(n19398), .A(n19088), .ZN(n19089) );
  OAI221_X1 U22333 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n19091), 
        .C1(n19394), .C2(n19090), .A(n19089), .ZN(P3_U2807) );
  INV_X1 U22334 ( .A(n19413), .ZN(n19409) );
  OR2_X1 U22335 ( .A1(n19405), .A2(n19334), .ZN(n19093) );
  OAI21_X1 U22336 ( .B1(n19409), .B2(n19130), .A(n19186), .ZN(n19119) );
  INV_X1 U22337 ( .A(n19119), .ZN(n19109) );
  NAND2_X1 U22338 ( .A1(n11878), .A2(n19212), .ZN(n19113) );
  AOI221_X1 U22339 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C1(n21843), .C2(n19096), .A(
        n19113), .ZN(n19098) );
  NAND2_X1 U22340 ( .A1(n19142), .A2(n19094), .ZN(n19095) );
  OAI211_X1 U22341 ( .C1(n11878), .C2(n19140), .A(n19313), .B(n19095), .ZN(
        n19129) );
  AOI21_X1 U22342 ( .B1(n19123), .B2(n19122), .A(n19129), .ZN(n19112) );
  OAI22_X1 U22343 ( .A1(n19112), .A2(n19096), .B1(n19613), .B2(n20171), .ZN(
        n19097) );
  AOI211_X1 U22344 ( .C1(n19099), .C2(n19236), .A(n19098), .B(n19097), .ZN(
        n19108) );
  AOI21_X1 U22345 ( .B1(n10328), .B2(n19102), .A(n19101), .ZN(n19103) );
  NOR2_X1 U22346 ( .A1(n19104), .A2(n19103), .ZN(n19105) );
  XNOR2_X1 U22347 ( .A(n19105), .B(n19419), .ZN(n19400) );
  AOI22_X1 U22348 ( .A1(n19400), .A2(n19254), .B1(n19106), .B2(n19419), .ZN(
        n19107) );
  OAI211_X1 U22349 ( .C1(n19109), .C2(n19419), .A(n19108), .B(n19107), .ZN(
        P3_U2808) );
  NAND3_X1 U22350 ( .A1(n10328), .A2(n10323), .A3(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n19147) );
  OAI22_X1 U22351 ( .A1(n19160), .A2(n19110), .B1(n19426), .B2(n19147), .ZN(
        n19111) );
  XOR2_X1 U22352 ( .A(n21966), .B(n19111), .Z(n19434) );
  NAND2_X1 U22353 ( .A1(n19556), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n19432) );
  OAI221_X1 U22354 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n19113), .C1(
        n21843), .C2(n19112), .A(n19432), .ZN(n19114) );
  AOI21_X1 U22355 ( .B1(n19236), .B2(n19115), .A(n19114), .ZN(n19121) );
  NOR2_X1 U22356 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n19426), .ZN(
        n19431) );
  NOR2_X1 U22357 ( .A1(n19116), .A2(n19159), .ZN(n19421) );
  NAND2_X1 U22358 ( .A1(n19117), .A2(n19421), .ZN(n19152) );
  INV_X1 U22359 ( .A(n19152), .ZN(n19118) );
  AOI22_X1 U22360 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n19119), .B1(
        n19431), .B2(n19118), .ZN(n19120) );
  OAI211_X1 U22361 ( .C1(n19434), .C2(n19204), .A(n19121), .B(n19120), .ZN(
        P3_U2809) );
  NAND2_X1 U22362 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n19136), .ZN(
        n19442) );
  OAI21_X1 U22363 ( .B1(n11882), .B2(n19863), .A(n19122), .ZN(n19128) );
  NOR2_X1 U22364 ( .A1(n19603), .A2(n20168), .ZN(n19127) );
  INV_X1 U22365 ( .A(n19124), .ZN(n19125) );
  AOI21_X1 U22366 ( .B1(n19183), .B2(n19082), .A(n19125), .ZN(n19126) );
  AOI211_X1 U22367 ( .C1(n19129), .C2(n19128), .A(n19127), .B(n19126), .ZN(
        n19138) );
  NAND2_X1 U22368 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n19421), .ZN(
        n19406) );
  INV_X1 U22369 ( .A(n19406), .ZN(n19436) );
  OAI21_X1 U22370 ( .B1(n19130), .B2(n19436), .A(n19186), .ZN(n19149) );
  INV_X1 U22371 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n19131) );
  NOR2_X1 U22372 ( .A1(n19147), .A2(n19131), .ZN(n19134) );
  OAI21_X1 U22373 ( .B1(n19134), .B2(n19133), .A(n19132), .ZN(n19135) );
  XOR2_X1 U22374 ( .A(n19136), .B(n19135), .Z(n19435) );
  AOI22_X1 U22375 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n19149), .B1(
        n19254), .B2(n19435), .ZN(n19137) );
  OAI211_X1 U22376 ( .C1(n19442), .C2(n19152), .A(n19138), .B(n19137), .ZN(
        P3_U2810) );
  NAND2_X1 U22377 ( .A1(n19139), .A2(n19212), .ZN(n19155) );
  AOI221_X1 U22378 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C1(n19154), .C2(n19143), .A(
        n19155), .ZN(n19145) );
  OAI21_X1 U22379 ( .B1(n19139), .B2(n19140), .A(n19313), .ZN(n19167) );
  AOI21_X1 U22380 ( .B1(n19142), .B2(n19141), .A(n19167), .ZN(n19153) );
  NAND2_X1 U22381 ( .A1(n19556), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n19445) );
  OAI21_X1 U22382 ( .B1(n19153), .B2(n19143), .A(n19445), .ZN(n19144) );
  AOI211_X1 U22383 ( .C1(n19146), .C2(n19236), .A(n19145), .B(n19144), .ZN(
        n19151) );
  OAI21_X1 U22384 ( .B1(n19160), .B2(n19158), .A(n19147), .ZN(n19148) );
  XOR2_X1 U22385 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B(n19148), .Z(
        n19443) );
  AOI22_X1 U22386 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n19149), .B1(
        n19254), .B2(n19443), .ZN(n19150) );
  OAI211_X1 U22387 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n19152), .A(
        n19151), .B(n19150), .ZN(P3_U2811) );
  NAND2_X1 U22388 ( .A1(n19455), .A2(n19159), .ZN(n19463) );
  NAND2_X1 U22389 ( .A1(n19556), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n19461) );
  OAI221_X1 U22390 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n19155), .C1(
        n19154), .C2(n19153), .A(n19461), .ZN(n19156) );
  AOI21_X1 U22391 ( .B1(n19236), .B2(n19157), .A(n19156), .ZN(n19163) );
  OAI21_X1 U22392 ( .B1(n19455), .B2(n19187), .A(n19186), .ZN(n19170) );
  OAI21_X1 U22393 ( .B1(n19159), .B2(n19196), .A(n19158), .ZN(n19161) );
  XOR2_X1 U22394 ( .A(n19161), .B(n19160), .Z(n19458) );
  AOI22_X1 U22395 ( .A1(n19170), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B1(
        n19254), .B2(n19458), .ZN(n19162) );
  OAI211_X1 U22396 ( .C1(n19187), .C2(n19463), .A(n19163), .B(n19162), .ZN(
        P3_U2812) );
  OAI21_X1 U22397 ( .B1(n19164), .B2(n19863), .A(n19165), .ZN(n19166) );
  AOI22_X1 U22398 ( .A1(n19556), .A2(P3_REIP_REG_17__SCAN_IN), .B1(n19167), 
        .B2(n19166), .ZN(n19172) );
  OAI21_X1 U22399 ( .B1(n19187), .B2(n10428), .A(n19464), .ZN(n19169) );
  XNOR2_X1 U22400 ( .A(n9882), .B(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n19469) );
  INV_X1 U22401 ( .A(n19469), .ZN(n19168) );
  AOI22_X1 U22402 ( .A1(n19170), .A2(n19169), .B1(n19254), .B2(n19168), .ZN(
        n19171) );
  OAI211_X1 U22403 ( .C1(n19309), .C2(n19173), .A(n19172), .B(n19171), .ZN(
        P3_U2813) );
  OAI22_X1 U22404 ( .A1(n19175), .A2(n10323), .B1(n19239), .B2(n19174), .ZN(
        n19176) );
  XOR2_X1 U22405 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n19176), .Z(
        n19479) );
  AOI22_X1 U22406 ( .A1(n19556), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n19177), .ZN(n19181) );
  OAI211_X1 U22407 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n19179), .B(n19178), .ZN(n19180) );
  OAI211_X1 U22408 ( .C1(n19183), .C2(n19182), .A(n19181), .B(n19180), .ZN(
        n19184) );
  AOI21_X1 U22409 ( .B1(n19254), .B2(n19479), .A(n19184), .ZN(n19185) );
  OAI221_X1 U22410 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n19187), 
        .C1(n10428), .C2(n19186), .A(n19185), .ZN(P3_U2814) );
  NAND2_X1 U22411 ( .A1(n19514), .A2(n19188), .ZN(n19211) );
  INV_X1 U22412 ( .A(n19211), .ZN(n19191) );
  OAI211_X1 U22413 ( .C1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n19191), .A(
        n19190), .B(n19189), .ZN(n19510) );
  AOI21_X1 U22414 ( .B1(n19213), .B2(n19192), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n19194) );
  OAI22_X1 U22415 ( .A1(n19309), .A2(n19195), .B1(n19194), .B2(n19193), .ZN(
        n19206) );
  NAND2_X1 U22416 ( .A1(n19196), .A2(n19524), .ZN(n19224) );
  NOR4_X1 U22417 ( .A1(n19198), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        n19197), .A4(n19224), .ZN(n19199) );
  AOI21_X1 U22418 ( .B1(n19200), .B2(n19450), .A(n19199), .ZN(n19201) );
  XNOR2_X1 U22419 ( .A(n19201), .B(n19502), .ZN(n19506) );
  AND2_X1 U22420 ( .A1(n19209), .A2(n19450), .ZN(n19203) );
  OAI21_X1 U22421 ( .B1(n19203), .B2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n19202), .ZN(n19503) );
  OAI22_X1 U22422 ( .A1(n19506), .A2(n19204), .B1(n19208), .B2(n19503), .ZN(
        n19205) );
  AOI211_X1 U22423 ( .C1(n19556), .C2(P3_REIP_REG_14__SCAN_IN), .A(n19206), 
        .B(n19205), .ZN(n19207) );
  OAI21_X1 U22424 ( .B1(n19334), .B2(n19510), .A(n19207), .ZN(P3_U2816) );
  AOI21_X1 U22425 ( .B1(n19209), .B2(n19514), .A(n19208), .ZN(n19210) );
  AOI21_X1 U22426 ( .B1(n19340), .B2(n19211), .A(n19210), .ZN(n19244) );
  NAND2_X1 U22427 ( .A1(n17854), .A2(n19212), .ZN(n19233) );
  AOI211_X1 U22428 ( .C1(n19232), .C2(n19218), .A(n19213), .B(n19233), .ZN(
        n19220) );
  OAI21_X1 U22429 ( .B1(n19215), .B2(n19214), .A(n19313), .ZN(n19216) );
  AOI21_X1 U22430 ( .B1(n19307), .B2(n19217), .A(n19216), .ZN(n19231) );
  OAI22_X1 U22431 ( .A1(n19231), .A2(n19218), .B1(n19603), .B2(n20155), .ZN(
        n19219) );
  AOI211_X1 U22432 ( .C1(n19236), .C2(n19221), .A(n19220), .B(n19219), .ZN(
        n19229) );
  INV_X1 U22433 ( .A(n19222), .ZN(n19223) );
  AOI21_X1 U22434 ( .B1(n19225), .B2(n19224), .A(n19223), .ZN(n19226) );
  XNOR2_X1 U22435 ( .A(n19226), .B(n19230), .ZN(n19521) );
  NOR2_X1 U22436 ( .A1(n19227), .A2(n19518), .ZN(n19241) );
  AOI22_X1 U22437 ( .A1(n19254), .A2(n19521), .B1(n19520), .B2(n19241), .ZN(
        n19228) );
  OAI211_X1 U22438 ( .C1(n19244), .C2(n19230), .A(n19229), .B(n19228), .ZN(
        P3_U2817) );
  NAND2_X1 U22439 ( .A1(n19556), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n19531) );
  OAI221_X1 U22440 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19233), .C1(
        n19232), .C2(n19231), .A(n19531), .ZN(n19234) );
  AOI21_X1 U22441 ( .B1(n19236), .B2(n19235), .A(n19234), .ZN(n19243) );
  INV_X1 U22442 ( .A(n19237), .ZN(n19238) );
  OAI21_X1 U22443 ( .B1(n19518), .B2(n19239), .A(n19238), .ZN(n19240) );
  XOR2_X1 U22444 ( .A(n19240), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(
        n19529) );
  AOI22_X1 U22445 ( .A1(n19254), .A2(n19529), .B1(n19241), .B2(n19524), .ZN(
        n19242) );
  OAI211_X1 U22446 ( .C1(n19244), .C2(n19524), .A(n19243), .B(n19242), .ZN(
        P3_U2818) );
  INV_X1 U22447 ( .A(n19245), .ZN(n19248) );
  INV_X1 U22448 ( .A(n19246), .ZN(n19247) );
  AOI21_X1 U22449 ( .B1(n19248), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n19247), .ZN(n19258) );
  AOI22_X1 U22450 ( .A1(n19556), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n19249), 
        .B2(n19344), .ZN(n19257) );
  AOI211_X1 U22451 ( .C1(n19252), .C2(n19251), .A(n19348), .B(n19250), .ZN(
        n19253) );
  AOI21_X1 U22452 ( .B1(n19255), .B2(n19254), .A(n19253), .ZN(n19256) );
  OAI211_X1 U22453 ( .C1(n19259), .C2(n19258), .A(n19257), .B(n19256), .ZN(
        P3_U2820) );
  INV_X1 U22454 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n20144) );
  NOR2_X1 U22455 ( .A1(n19613), .A2(n20144), .ZN(n19537) );
  AOI221_X1 U22456 ( .B1(n19262), .B2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C1(
        n19261), .C2(n19260), .A(n19537), .ZN(n19271) );
  AOI21_X1 U22457 ( .B1(n19265), .B2(n19264), .A(n19263), .ZN(n19266) );
  XOR2_X1 U22458 ( .A(n19266), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n19539) );
  INV_X1 U22459 ( .A(n19342), .ZN(n19328) );
  OAI21_X1 U22460 ( .B1(n19268), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n19267), .ZN(n19269) );
  INV_X1 U22461 ( .A(n19269), .ZN(n19538) );
  AOI22_X1 U22462 ( .A1(n19539), .A2(n19340), .B1(n19328), .B2(n19538), .ZN(
        n19270) );
  OAI211_X1 U22463 ( .C1(n19309), .C2(n19272), .A(n19271), .B(n19270), .ZN(
        P3_U2823) );
  NOR2_X1 U22464 ( .A1(n11890), .A2(n19863), .ZN(n19278) );
  INV_X1 U22465 ( .A(n19278), .ZN(n19285) );
  NAND2_X1 U22466 ( .A1(n19274), .A2(n19273), .ZN(n19275) );
  NAND2_X1 U22467 ( .A1(n19276), .A2(n19275), .ZN(n19543) );
  OAI22_X1 U22468 ( .A1(n19342), .A2(n19543), .B1(n19613), .B2(n20142), .ZN(
        n19277) );
  INV_X1 U22469 ( .A(n19277), .ZN(n19284) );
  NOR2_X1 U22470 ( .A1(n19348), .A2(n19278), .ZN(n19294) );
  OAI21_X1 U22471 ( .B1(n19280), .B2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n19279), .ZN(n19551) );
  OAI22_X1 U22472 ( .A1(n19309), .A2(n19281), .B1(n19334), .B2(n19551), .ZN(
        n19282) );
  AOI21_X1 U22473 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n19294), .A(
        n19282), .ZN(n19283) );
  OAI211_X1 U22474 ( .C1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n19285), .A(
        n19284), .B(n19283), .ZN(P3_U2824) );
  XNOR2_X1 U22475 ( .A(n19286), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n19287) );
  XNOR2_X1 U22476 ( .A(n19288), .B(n19287), .ZN(n19552) );
  OAI21_X1 U22477 ( .B1(n19291), .B2(n19290), .A(n19289), .ZN(n19559) );
  INV_X1 U22478 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n20141) );
  OAI22_X1 U22479 ( .A1(n19334), .A2(n19559), .B1(n19603), .B2(n20141), .ZN(
        n19292) );
  AOI21_X1 U22480 ( .B1(n19293), .B2(n19344), .A(n19292), .ZN(n19296) );
  OAI221_X1 U22481 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n18534), .C1(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n19313), .A(n19294), .ZN(n19295) );
  OAI211_X1 U22482 ( .C1(n19342), .C2(n19552), .A(n19296), .B(n19295), .ZN(
        P3_U2825) );
  OAI21_X1 U22483 ( .B1(n19299), .B2(n19298), .A(n19297), .ZN(n19300) );
  XOR2_X1 U22484 ( .A(n19300), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(
        n19573) );
  AOI22_X1 U22485 ( .A1(n19566), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n20002), 
        .B2(n19301), .ZN(n19312) );
  OAI21_X1 U22486 ( .B1(n19304), .B2(n19303), .A(n19302), .ZN(n19305) );
  INV_X1 U22487 ( .A(n19305), .ZN(n19567) );
  AOI21_X1 U22488 ( .B1(n19307), .B2(n18545), .A(n19306), .ZN(n19324) );
  OAI22_X1 U22489 ( .A1(n19309), .A2(n19308), .B1(n19324), .B2(n18554), .ZN(
        n19310) );
  AOI21_X1 U22490 ( .B1(n19328), .B2(n19567), .A(n19310), .ZN(n19311) );
  OAI211_X1 U22491 ( .C1(n19334), .C2(n19573), .A(n19312), .B(n19311), .ZN(
        P3_U2826) );
  NAND2_X1 U22492 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n19313), .ZN(
        n19330) );
  INV_X1 U22493 ( .A(n19314), .ZN(n19321) );
  OAI21_X1 U22494 ( .B1(n19317), .B2(n19316), .A(n19315), .ZN(n19583) );
  XOR2_X1 U22495 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n19318), .Z(
        n19579) );
  NOR2_X1 U22496 ( .A1(n19603), .A2(n20137), .ZN(n19578) );
  AOI21_X1 U22497 ( .B1(n19328), .B2(n19579), .A(n19578), .ZN(n19319) );
  OAI21_X1 U22498 ( .B1(n19583), .B2(n19334), .A(n19319), .ZN(n19320) );
  AOI21_X1 U22499 ( .B1(n19344), .B2(n19321), .A(n19320), .ZN(n19322) );
  OAI221_X1 U22500 ( .B1(n19324), .B2(n19323), .C1(n19324), .C2(n19330), .A(
        n19322), .ZN(P3_U2827) );
  INV_X1 U22501 ( .A(n19327), .ZN(n19586) );
  AOI22_X1 U22502 ( .A1(n19344), .A2(n19329), .B1(n19328), .B2(n19586), .ZN(
        n19337) );
  OAI21_X1 U22503 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n20002), .A(
        n19330), .ZN(n19336) );
  NAND2_X1 U22504 ( .A1(n19556), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n19599) );
  OAI21_X1 U22505 ( .B1(n19333), .B2(n19332), .A(n19331), .ZN(n19601) );
  OR2_X1 U22506 ( .A1(n19334), .A2(n19601), .ZN(n19335) );
  NAND4_X1 U22507 ( .A1(n19337), .A2(n19336), .A3(n19599), .A4(n19335), .ZN(
        P3_U2828) );
  AOI21_X1 U22508 ( .B1(n19340), .B2(n19339), .A(n19338), .ZN(n19346) );
  NOR2_X1 U22509 ( .A1(n19342), .A2(n19341), .ZN(n19343) );
  AOI21_X1 U22510 ( .B1(n19344), .B2(n19347), .A(n19343), .ZN(n19345) );
  OAI211_X1 U22511 ( .C1(n19348), .C2(n19347), .A(n19346), .B(n19345), .ZN(
        P3_U2829) );
  NOR2_X1 U22512 ( .A1(n19349), .A2(n19395), .ZN(n19360) );
  OAI21_X1 U22513 ( .B1(n19419), .B2(n19526), .A(n19350), .ZN(n19411) );
  AOI21_X1 U22514 ( .B1(n19351), .B2(n19411), .A(n19561), .ZN(n19383) );
  AOI21_X1 U22515 ( .B1(n19352), .B2(n19589), .A(n19383), .ZN(n19373) );
  OAI22_X1 U22516 ( .A1(n19438), .A2(n19353), .B1(n19410), .B2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n19354) );
  AOI21_X1 U22517 ( .B1(n20057), .B2(n19355), .A(n19354), .ZN(n19356) );
  OAI211_X1 U22518 ( .C1(n19357), .C2(n19401), .A(n19373), .B(n19356), .ZN(
        n19363) );
  AOI21_X1 U22519 ( .B1(n19604), .B2(n22049), .A(n19363), .ZN(n19358) );
  INV_X1 U22520 ( .A(n19358), .ZN(n19359) );
  MUX2_X1 U22521 ( .A(n19360), .B(n19359), .S(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .Z(n19361) );
  INV_X1 U22522 ( .A(n19363), .ZN(n19365) );
  OAI22_X1 U22523 ( .A1(n19365), .A2(n22049), .B1(n19395), .B2(n19364), .ZN(
        n19367) );
  AOI22_X1 U22524 ( .A1(n19367), .A2(n19598), .B1(n19530), .B2(n19366), .ZN(
        n19369) );
  OAI211_X1 U22525 ( .C1(n19564), .C2(n22049), .A(n19369), .B(n19368), .ZN(
        P3_U2836) );
  AOI21_X1 U22526 ( .B1(n19598), .B2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n19370), .ZN(n19371) );
  AOI21_X1 U22527 ( .B1(n19373), .B2(n19372), .A(n19371), .ZN(n19374) );
  AOI211_X1 U22528 ( .C1(n19602), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n19375), .B(n19374), .ZN(n19379) );
  AOI22_X1 U22529 ( .A1(n19610), .A2(n19377), .B1(n19530), .B2(n19376), .ZN(
        n19378) );
  OAI211_X1 U22530 ( .C1(n19504), .C2(n19380), .A(n19379), .B(n19378), .ZN(
        P3_U2837) );
  NAND2_X1 U22531 ( .A1(n19598), .A2(n19420), .ZN(n19393) );
  INV_X1 U22532 ( .A(n19381), .ZN(n19382) );
  AOI22_X1 U22533 ( .A1(n19382), .A2(n19530), .B1(n19566), .B2(
        P3_REIP_REG_24__SCAN_IN), .ZN(n19391) );
  AOI211_X1 U22534 ( .C1(n20057), .C2(n19384), .A(n19602), .B(n19383), .ZN(
        n19385) );
  OAI21_X1 U22535 ( .B1(n19386), .B2(n19401), .A(n19385), .ZN(n19389) );
  AOI211_X1 U22536 ( .C1(n20058), .C2(n19387), .A(n19394), .B(n19389), .ZN(
        n19388) );
  NOR2_X1 U22537 ( .A1(n19556), .A2(n19388), .ZN(n19397) );
  OAI211_X1 U22538 ( .C1(n19477), .C2(n19389), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n19397), .ZN(n19390) );
  OAI211_X1 U22539 ( .C1(n19393), .C2(n19392), .A(n19391), .B(n19390), .ZN(
        P3_U2838) );
  OAI21_X1 U22540 ( .B1(n19602), .B2(n19395), .A(n19394), .ZN(n19396) );
  AOI22_X1 U22541 ( .A1(n19530), .A2(n19398), .B1(n19397), .B2(n19396), .ZN(
        n19399) );
  OAI21_X1 U22542 ( .B1(n19603), .B2(n20173), .A(n19399), .ZN(P3_U2839) );
  AOI22_X1 U22543 ( .A1(n19556), .A2(P3_REIP_REG_22__SCAN_IN), .B1(n19530), 
        .B2(n19400), .ZN(n19418) );
  INV_X1 U22544 ( .A(n19401), .ZN(n19402) );
  NAND2_X1 U22545 ( .A1(n19403), .A2(n19402), .ZN(n19486) );
  OAI21_X1 U22546 ( .B1(n19405), .B2(n19404), .A(n19486), .ZN(n19422) );
  OAI21_X1 U22547 ( .B1(n19474), .B2(n19406), .A(n19604), .ZN(n19407) );
  OAI221_X1 U22548 ( .B1(n19560), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), 
        .C1(n19560), .C2(n19454), .A(n19407), .ZN(n19423) );
  OAI22_X1 U22549 ( .A1(n19410), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n19409), .B2(n19513), .ZN(n19425) );
  AOI211_X1 U22550 ( .C1(n20058), .C2(n19426), .A(n19423), .B(n19425), .ZN(
        n19412) );
  OAI211_X1 U22551 ( .C1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n19516), .A(
        n19412), .B(n19411), .ZN(n19416) );
  OAI21_X1 U22552 ( .B1(n19414), .B2(n19413), .A(n19419), .ZN(n19415) );
  OAI211_X1 U22553 ( .C1(n19422), .C2(n19416), .A(n19598), .B(n19415), .ZN(
        n19417) );
  OAI211_X1 U22554 ( .C1(n19564), .C2(n19419), .A(n19418), .B(n19417), .ZN(
        P3_U2840) );
  NAND3_X1 U22555 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n19598), .A3(
        n19420), .ZN(n19447) );
  INV_X1 U22556 ( .A(n19447), .ZN(n19430) );
  NAND3_X1 U22557 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n19453), .A3(
        n19421), .ZN(n19424) );
  AOI21_X1 U22558 ( .B1(n19427), .B2(n19426), .A(n19425), .ZN(n19428) );
  AOI211_X1 U22559 ( .C1(n19437), .C2(n19428), .A(n19556), .B(n21966), .ZN(
        n19429) );
  AOI21_X1 U22560 ( .B1(n19431), .B2(n19430), .A(n19429), .ZN(n19433) );
  OAI211_X1 U22561 ( .C1(n19434), .C2(n19505), .A(n19433), .B(n19432), .ZN(
        P3_U2841) );
  AOI22_X1 U22562 ( .A1(n19556), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n19530), 
        .B2(n19435), .ZN(n19441) );
  AOI221_X1 U22563 ( .B1(n19513), .B2(n19437), .C1(n19436), .C2(n19437), .A(
        n19556), .ZN(n19444) );
  NOR3_X1 U22564 ( .A1(n19438), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n20107), .ZN(n19439) );
  OAI21_X1 U22565 ( .B1(n19444), .B2(n19439), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n19440) );
  OAI211_X1 U22566 ( .C1(n19447), .C2(n19442), .A(n19441), .B(n19440), .ZN(
        P3_U2842) );
  AOI22_X1 U22567 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n19444), .B1(
        n19530), .B2(n19443), .ZN(n19446) );
  OAI211_X1 U22568 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n19447), .A(
        n19446), .B(n19445), .ZN(P3_U2843) );
  NOR2_X1 U22569 ( .A1(n19576), .A2(n19448), .ZN(n19536) );
  NAND3_X1 U22570 ( .A1(n19450), .A2(n19449), .A3(n19536), .ZN(n19501) );
  NOR2_X1 U22571 ( .A1(n19502), .A2(n19501), .ZN(n19484) );
  OAI211_X1 U22572 ( .C1(n19451), .C2(n19484), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n19598), .ZN(n19482) );
  NAND3_X1 U22573 ( .A1(n19453), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n19452), .ZN(n19457) );
  OAI22_X1 U22574 ( .A1(n19455), .A2(n19513), .B1(n19454), .B2(n19560), .ZN(
        n19456) );
  AOI211_X1 U22575 ( .C1(n19589), .C2(n19457), .A(n19478), .B(n19456), .ZN(
        n19466) );
  OAI21_X1 U22576 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n19561), .A(
        n19466), .ZN(n19460) );
  NOR2_X1 U22577 ( .A1(n19566), .A2(n19159), .ZN(n19459) );
  AOI22_X1 U22578 ( .A1(n19460), .A2(n19459), .B1(n19530), .B2(n19458), .ZN(
        n19462) );
  OAI211_X1 U22579 ( .C1(n19463), .C2(n19482), .A(n19462), .B(n19461), .ZN(
        P3_U2844) );
  OR2_X1 U22580 ( .A1(n19556), .A2(n19464), .ZN(n19465) );
  OR2_X1 U22581 ( .A1(n19466), .A2(n19465), .ZN(n19468) );
  OR3_X1 U22582 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n10428), .A3(
        n19482), .ZN(n19467) );
  OAI211_X1 U22583 ( .C1(n19505), .C2(n19469), .A(n19468), .B(n19467), .ZN(
        n19470) );
  INV_X1 U22584 ( .A(n19470), .ZN(n19471) );
  OAI21_X1 U22585 ( .B1(n19603), .B2(n20162), .A(n19471), .ZN(P3_U2845) );
  NOR2_X1 U22586 ( .A1(n19473), .A2(n19472), .ZN(n19496) );
  OAI22_X1 U22587 ( .A1(n19526), .A2(n17843), .B1(n19606), .B2(n19474), .ZN(
        n19475) );
  OAI211_X1 U22588 ( .C1(n19476), .C2(n19516), .A(n19496), .B(n19475), .ZN(
        n19483) );
  OAI221_X1 U22589 ( .B1(n19478), .B2(n19477), .C1(n19478), .C2(n19483), .A(
        n19603), .ZN(n19481) );
  AOI22_X1 U22590 ( .A1(n19556), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n19530), 
        .B2(n19479), .ZN(n19480) );
  OAI221_X1 U22591 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n19482), 
        .C1(n10428), .C2(n19481), .A(n19480), .ZN(P3_U2846) );
  AOI22_X1 U22592 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n19602), .B1(
        n19556), .B2(P3_REIP_REG_15__SCAN_IN), .ZN(n19494) );
  OAI21_X1 U22593 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n19484), .A(
        n19483), .ZN(n19485) );
  OAI21_X1 U22594 ( .B1(n19487), .B2(n19486), .A(n19485), .ZN(n19489) );
  AOI22_X1 U22595 ( .A1(n19598), .A2(n19489), .B1(n19530), .B2(n19488), .ZN(
        n19493) );
  NAND3_X1 U22596 ( .A1(n19610), .A2(n19491), .A3(n19490), .ZN(n19492) );
  NAND3_X1 U22597 ( .A1(n19494), .A2(n19493), .A3(n19492), .ZN(P3_U2847) );
  NAND3_X1 U22598 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n19514), .A3(
        n19495), .ZN(n19527) );
  NAND2_X1 U22599 ( .A1(n19526), .A2(n19527), .ZN(n19515) );
  NAND3_X1 U22600 ( .A1(n19496), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n19515), .ZN(n19499) );
  AOI222_X1 U22601 ( .A1(n19499), .A2(n19598), .B1(n19602), .B2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C1(n19498), .C2(n19497), .ZN(
        n19500) );
  AOI21_X1 U22602 ( .B1(n19502), .B2(n19501), .A(n19500), .ZN(n19508) );
  OAI22_X1 U22603 ( .A1(n19506), .A2(n19505), .B1(n19504), .B2(n19503), .ZN(
        n19507) );
  AOI211_X1 U22604 ( .C1(P3_REIP_REG_14__SCAN_IN), .C2(n19556), .A(n19508), 
        .B(n19507), .ZN(n19509) );
  OAI21_X1 U22605 ( .B1(n10311), .B2(n19510), .A(n19509), .ZN(P3_U2848) );
  OAI211_X1 U22606 ( .C1(n19514), .C2(n19513), .A(n19512), .B(n19511), .ZN(
        n19525) );
  OAI211_X1 U22607 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n19516), .A(
        n19598), .B(n19515), .ZN(n19517) );
  OAI21_X1 U22608 ( .B1(n19525), .B2(n19517), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n19523) );
  NOR2_X1 U22609 ( .A1(n19519), .A2(n19518), .ZN(n19528) );
  AOI22_X1 U22610 ( .A1(n19530), .A2(n19521), .B1(n19520), .B2(n19528), .ZN(
        n19522) );
  OAI221_X1 U22611 ( .B1(n19556), .B2(n19523), .C1(n19603), .C2(n20155), .A(
        n19522), .ZN(P3_U2849) );
  AOI211_X1 U22612 ( .C1(n19527), .C2(n19526), .A(n19525), .B(n19524), .ZN(
        n19534) );
  AOI21_X1 U22613 ( .B1(n19598), .B2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n19528), .ZN(n19533) );
  AOI22_X1 U22614 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n19602), .B1(
        n19530), .B2(n19529), .ZN(n19532) );
  OAI211_X1 U22615 ( .C1(n19534), .C2(n19533), .A(n19532), .B(n19531), .ZN(
        P3_U2850) );
  OAI221_X1 U22616 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n19536), .A(n19535), .ZN(
        n19542) );
  AOI21_X1 U22617 ( .B1(n19602), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n19537), .ZN(n19541) );
  INV_X1 U22618 ( .A(n19605), .ZN(n19580) );
  AOI22_X1 U22619 ( .A1(n19539), .A2(n19610), .B1(n19580), .B2(n19538), .ZN(
        n19540) );
  OAI211_X1 U22620 ( .C1(n19575), .C2(n19542), .A(n19541), .B(n19540), .ZN(
        P3_U2855) );
  INV_X1 U22621 ( .A(n19543), .ZN(n19549) );
  OAI21_X1 U22622 ( .B1(n19575), .B2(n19544), .A(n19603), .ZN(n19553) );
  NAND2_X1 U22623 ( .A1(n19556), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n19545) );
  OAI221_X1 U22624 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n19547), .C1(
        n19546), .C2(n19553), .A(n19545), .ZN(n19548) );
  AOI21_X1 U22625 ( .B1(n19580), .B2(n19549), .A(n19548), .ZN(n19550) );
  OAI21_X1 U22626 ( .B1(n10311), .B2(n19551), .A(n19550), .ZN(P3_U2856) );
  NOR3_X1 U22627 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n10424), .A3(
        n19569), .ZN(n19555) );
  OAI22_X1 U22628 ( .A1(n10011), .A2(n19553), .B1(n19605), .B2(n19552), .ZN(
        n19554) );
  AOI21_X1 U22629 ( .B1(n19570), .B2(n19555), .A(n19554), .ZN(n19558) );
  NAND2_X1 U22630 ( .A1(n19556), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n19557) );
  OAI211_X1 U22631 ( .C1(n10311), .C2(n19559), .A(n19558), .B(n19557), .ZN(
        P3_U2857) );
  OAI22_X1 U22632 ( .A1(n19562), .A2(n19561), .B1(n19560), .B2(n19584), .ZN(
        n19563) );
  NOR3_X1 U22633 ( .A1(n19591), .A2(n10424), .A3(n19563), .ZN(n19574) );
  OAI21_X1 U22634 ( .B1(n19574), .B2(n19565), .A(n19564), .ZN(n19568) );
  AOI222_X1 U22635 ( .A1(n19568), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B1(
        n19580), .B2(n19567), .C1(P3_REIP_REG_4__SCAN_IN), .C2(n19566), .ZN(
        n19572) );
  NAND3_X1 U22636 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n19570), .A3(
        n19569), .ZN(n19571) );
  OAI211_X1 U22637 ( .C1(n19573), .C2(n10311), .A(n19572), .B(n19571), .ZN(
        P3_U2858) );
  AOI211_X1 U22638 ( .C1(n19576), .C2(n10424), .A(n19575), .B(n19574), .ZN(
        n19577) );
  AOI211_X1 U22639 ( .C1(n19580), .C2(n19579), .A(n19578), .B(n19577), .ZN(
        n19582) );
  NAND2_X1 U22640 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n19602), .ZN(
        n19581) );
  OAI211_X1 U22641 ( .C1(n19583), .C2(n10311), .A(n19582), .B(n19581), .ZN(
        P3_U2859) );
  NAND2_X1 U22642 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19585) );
  OAI21_X1 U22643 ( .B1(n19585), .B2(n19592), .A(n19584), .ZN(n19588) );
  AOI22_X1 U22644 ( .A1(n20058), .A2(n19588), .B1(n19587), .B2(n19586), .ZN(
        n19596) );
  OAI211_X1 U22645 ( .C1(n19591), .C2(n19590), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n19589), .ZN(n19595) );
  NAND3_X1 U22646 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n19593), .A3(
        n19592), .ZN(n19594) );
  NAND3_X1 U22647 ( .A1(n19596), .A2(n19595), .A3(n19594), .ZN(n19597) );
  AOI22_X1 U22648 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n19602), .B1(
        n19598), .B2(n19597), .ZN(n19600) );
  OAI211_X1 U22649 ( .C1(n10311), .C2(n19601), .A(n19600), .B(n19599), .ZN(
        P3_U2860) );
  AOI21_X1 U22650 ( .B1(n19604), .B2(n19603), .A(n19602), .ZN(n19607) );
  OAI22_X1 U22651 ( .A1(n19607), .A2(n19606), .B1(n19605), .B2(n19609), .ZN(
        n19608) );
  AOI21_X1 U22652 ( .B1(n19610), .B2(n19609), .A(n19608), .ZN(n19612) );
  OAI211_X1 U22653 ( .C1(n13938), .C2(n19613), .A(n19612), .B(n19611), .ZN(
        P3_U2862) );
  NAND2_X1 U22654 ( .A1(n17985), .A2(n19614), .ZN(n19617) );
  AOI21_X1 U22655 ( .B1(n19617), .B2(n19616), .A(n19615), .ZN(n20099) );
  INV_X1 U22656 ( .A(n19618), .ZN(n19661) );
  OAI21_X1 U22657 ( .B1(n20099), .B2(n19661), .A(n19623), .ZN(n19619) );
  OAI221_X1 U22658 ( .B1(n12089), .B2(n20211), .C1(n12089), .C2(n19623), .A(
        n19619), .ZN(P3_U2863) );
  INV_X1 U22659 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20087) );
  NAND2_X1 U22660 ( .A1(n20085), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19861) );
  INV_X1 U22661 ( .A(n19861), .ZN(n19887) );
  NAND2_X1 U22662 ( .A1(n20087), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19749) );
  INV_X1 U22663 ( .A(n19749), .ZN(n19794) );
  NOR2_X1 U22664 ( .A1(n19887), .A2(n19794), .ZN(n19621) );
  OAI22_X1 U22665 ( .A1(n19622), .A2(n20087), .B1(n19621), .B2(n19620), .ZN(
        P3_U2866) );
  NOR2_X1 U22666 ( .A1(n20088), .A2(n19623), .ZN(P3_U2867) );
  NAND2_X1 U22667 ( .A1(n20002), .A2(BUF2_REG_16__SCAN_IN), .ZN(n19972) );
  NOR2_X1 U22668 ( .A1(n20087), .A2(n19839), .ZN(n20000) );
  NAND2_X1 U22669 ( .A1(n20000), .A2(n12089), .ZN(n19996) );
  NAND2_X1 U22670 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n20002), .ZN(n20006) );
  NAND2_X1 U22671 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12088), .ZN(
        n19841) );
  NOR2_X1 U22672 ( .A1(n20085), .A2(n20087), .ZN(n19940) );
  INV_X1 U22673 ( .A(n19940), .ZN(n19938) );
  NOR2_X2 U22674 ( .A1(n19841), .A2(n19938), .ZN(n20048) );
  NOR2_X2 U22675 ( .A1(n19912), .A2(n19624), .ZN(n19997) );
  NOR2_X1 U22676 ( .A1(n12088), .A2(n12089), .ZN(n20075) );
  INV_X1 U22677 ( .A(n20075), .ZN(n19704) );
  NOR2_X2 U22678 ( .A1(n19704), .A2(n19938), .ZN(n20040) );
  INV_X1 U22679 ( .A(n20040), .ZN(n20055) );
  NAND2_X1 U22680 ( .A1(n12088), .A2(n12089), .ZN(n20081) );
  NOR2_X1 U22681 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19702) );
  NOR2_X2 U22682 ( .A1(n20081), .A2(n19703), .ZN(n19723) );
  AOI21_X1 U22683 ( .B1(n20055), .B2(n19718), .A(n20110), .ZN(n19657) );
  AOI22_X1 U22684 ( .A1(n19969), .A2(n20048), .B1(n19997), .B2(n19657), .ZN(
        n19630) );
  NAND2_X1 U22685 ( .A1(n19996), .A2(n20036), .ZN(n19968) );
  OAI21_X1 U22686 ( .B1(n12089), .B2(n21986), .A(n19862), .ZN(n19681) );
  AOI21_X1 U22687 ( .B1(n20055), .B2(n19718), .A(n19681), .ZN(n19683) );
  AOI21_X1 U22688 ( .B1(n20002), .B2(n19968), .A(n19683), .ZN(n19658) );
  INV_X1 U22689 ( .A(n19625), .ZN(n19626) );
  NAND2_X1 U22690 ( .A1(n19627), .A2(n19626), .ZN(n19653) );
  NOR2_X2 U22691 ( .A1(n19628), .A2(n19653), .ZN(n20003) );
  AOI22_X1 U22692 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19658), .B1(
        n20003), .B2(n19723), .ZN(n19629) );
  OAI211_X1 U22693 ( .C1(n19972), .C2(n19996), .A(n19630), .B(n19629), .ZN(
        P3_U2868) );
  NAND2_X1 U22694 ( .A1(n20002), .A2(BUF2_REG_17__SCAN_IN), .ZN(n20012) );
  NOR2_X2 U22695 ( .A1(n19912), .A2(n21987), .ZN(n20008) );
  NAND2_X1 U22696 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n20002), .ZN(n19976) );
  INV_X1 U22697 ( .A(n19976), .ZN(n20007) );
  AOI22_X1 U22698 ( .A1(n20008), .A2(n19657), .B1(n20007), .B2(n20048), .ZN(
        n19632) );
  NOR2_X2 U22699 ( .A1(n20217), .A2(n19653), .ZN(n20009) );
  AOI22_X1 U22700 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19658), .B1(
        n20009), .B2(n19723), .ZN(n19631) );
  OAI211_X1 U22701 ( .C1(n20012), .C2(n19996), .A(n19632), .B(n19631), .ZN(
        P3_U2869) );
  NAND2_X1 U22702 ( .A1(n20002), .A2(BUF2_REG_18__SCAN_IN), .ZN(n19949) );
  NOR2_X2 U22703 ( .A1(n19912), .A2(n19633), .ZN(n20013) );
  NAND2_X1 U22704 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n20002), .ZN(n20018) );
  AOI22_X1 U22705 ( .A1(n20013), .A2(n19657), .B1(n19946), .B2(n20048), .ZN(
        n19636) );
  NOR2_X2 U22706 ( .A1(n19634), .A2(n19653), .ZN(n20015) );
  AOI22_X1 U22707 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19658), .B1(
        n20015), .B2(n19723), .ZN(n19635) );
  OAI211_X1 U22708 ( .C1(n19949), .C2(n19996), .A(n19636), .B(n19635), .ZN(
        P3_U2870) );
  NAND2_X1 U22709 ( .A1(n20002), .A2(BUF2_REG_19__SCAN_IN), .ZN(n19953) );
  NAND2_X1 U22710 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n20002), .ZN(n20024) );
  INV_X1 U22711 ( .A(n20024), .ZN(n19950) );
  NOR2_X2 U22712 ( .A1(n19912), .A2(n19637), .ZN(n20019) );
  AOI22_X1 U22713 ( .A1(n19950), .A2(n20048), .B1(n20019), .B2(n19657), .ZN(
        n19640) );
  NOR2_X2 U22714 ( .A1(n19638), .A2(n19653), .ZN(n20021) );
  AOI22_X1 U22715 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19658), .B1(
        n20021), .B2(n19723), .ZN(n19639) );
  OAI211_X1 U22716 ( .C1(n19953), .C2(n19996), .A(n19640), .B(n19639), .ZN(
        P3_U2871) );
  NAND2_X1 U22717 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n20002), .ZN(n20030) );
  NAND2_X1 U22718 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n20002), .ZN(n19984) );
  INV_X1 U22719 ( .A(n19984), .ZN(n20026) );
  INV_X1 U22720 ( .A(n19996), .ZN(n19987) );
  NOR2_X2 U22721 ( .A1(n19641), .A2(n19912), .ZN(n20025) );
  AOI22_X1 U22722 ( .A1(n20026), .A2(n19987), .B1(n20025), .B2(n19657), .ZN(
        n19644) );
  NOR2_X2 U22723 ( .A1(n19642), .A2(n19653), .ZN(n20027) );
  AOI22_X1 U22724 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19658), .B1(
        n20027), .B2(n19723), .ZN(n19643) );
  OAI211_X1 U22725 ( .C1(n20030), .C2(n20036), .A(n19644), .B(n19643), .ZN(
        P3_U2872) );
  NAND2_X1 U22726 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n20002), .ZN(n19901) );
  NAND2_X1 U22727 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n20002), .ZN(n20037) );
  INV_X1 U22728 ( .A(n20037), .ZN(n19898) );
  NOR2_X2 U22729 ( .A1(n19645), .A2(n19912), .ZN(n20031) );
  AOI22_X1 U22730 ( .A1(n19898), .A2(n19987), .B1(n20031), .B2(n19657), .ZN(
        n19648) );
  NOR2_X2 U22731 ( .A1(n19646), .A2(n19653), .ZN(n20033) );
  AOI22_X1 U22732 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19658), .B1(
        n20033), .B2(n19723), .ZN(n19647) );
  OAI211_X1 U22733 ( .C1(n19901), .C2(n20036), .A(n19648), .B(n19647), .ZN(
        P3_U2873) );
  NAND2_X1 U22734 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n20002), .ZN(n20045) );
  NOR2_X2 U22735 ( .A1(n19649), .A2(n19912), .ZN(n20038) );
  AOI22_X1 U22736 ( .A1(n20039), .A2(n19987), .B1(n20038), .B2(n19657), .ZN(
        n19652) );
  NOR2_X2 U22737 ( .A1(n19650), .A2(n19653), .ZN(n20041) );
  AOI22_X1 U22738 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19658), .B1(
        n20041), .B2(n19723), .ZN(n19651) );
  OAI211_X1 U22739 ( .C1(n20045), .C2(n20036), .A(n19652), .B(n19651), .ZN(
        P3_U2874) );
  INV_X1 U22740 ( .A(n19653), .ZN(n19655) );
  NAND2_X1 U22741 ( .A1(n19655), .A2(n19654), .ZN(n20056) );
  NOR2_X2 U22742 ( .A1(n19656), .A2(n19863), .ZN(n20051) );
  NOR2_X2 U22743 ( .A1(n21919), .A2(n19912), .ZN(n20047) );
  AOI22_X1 U22744 ( .A1(n20051), .A2(n20048), .B1(n20047), .B2(n19657), .ZN(
        n19660) );
  AND2_X1 U22745 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n20002), .ZN(n20049) );
  AOI22_X1 U22746 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19658), .B1(
        n20049), .B2(n19987), .ZN(n19659) );
  OAI211_X1 U22747 ( .C1(n20056), .C2(n19718), .A(n19660), .B(n19659), .ZN(
        P3_U2875) );
  INV_X1 U22748 ( .A(n19972), .ZN(n19998) );
  NAND2_X1 U22749 ( .A1(n12088), .A2(n20102), .ZN(n19937) );
  NOR2_X1 U22750 ( .A1(n19703), .A2(n19937), .ZN(n19677) );
  AOI22_X1 U22751 ( .A1(n19998), .A2(n20040), .B1(n19997), .B2(n19677), .ZN(
        n19663) );
  NOR2_X1 U22752 ( .A1(n19912), .A2(n19661), .ZN(n19999) );
  INV_X1 U22753 ( .A(n19999), .ZN(n19792) );
  NOR2_X1 U22754 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19792), .ZN(
        n19939) );
  AOI22_X1 U22755 ( .A1(n20002), .A2(n20000), .B1(n19702), .B2(n19939), .ZN(
        n19678) );
  NOR2_X1 U22756 ( .A1(n19703), .A2(n19841), .ZN(n19676) );
  AOI22_X1 U22757 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19678), .B1(
        n19744), .B2(n20003), .ZN(n19662) );
  OAI211_X1 U22758 ( .C1(n20006), .C2(n19996), .A(n19663), .B(n19662), .ZN(
        P3_U2876) );
  INV_X1 U22759 ( .A(n20012), .ZN(n19973) );
  AOI22_X1 U22760 ( .A1(n19973), .A2(n20040), .B1(n20008), .B2(n19677), .ZN(
        n19665) );
  AOI22_X1 U22761 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19678), .B1(
        n19744), .B2(n20009), .ZN(n19664) );
  OAI211_X1 U22762 ( .C1(n19976), .C2(n19996), .A(n19665), .B(n19664), .ZN(
        P3_U2877) );
  AOI22_X1 U22763 ( .A1(n20013), .A2(n19677), .B1(n19946), .B2(n19987), .ZN(
        n19667) );
  AOI22_X1 U22764 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19678), .B1(
        n19744), .B2(n20015), .ZN(n19666) );
  OAI211_X1 U22765 ( .C1(n19949), .C2(n20055), .A(n19667), .B(n19666), .ZN(
        P3_U2878) );
  AOI22_X1 U22766 ( .A1(n19950), .A2(n19987), .B1(n20019), .B2(n19677), .ZN(
        n19669) );
  AOI22_X1 U22767 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19678), .B1(
        n19744), .B2(n20021), .ZN(n19668) );
  OAI211_X1 U22768 ( .C1(n19953), .C2(n20055), .A(n19669), .B(n19668), .ZN(
        P3_U2879) );
  INV_X1 U22769 ( .A(n20030), .ZN(n19981) );
  AOI22_X1 U22770 ( .A1(n20025), .A2(n19677), .B1(n19981), .B2(n19987), .ZN(
        n19671) );
  AOI22_X1 U22771 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19678), .B1(
        n19744), .B2(n20027), .ZN(n19670) );
  OAI211_X1 U22772 ( .C1(n19984), .C2(n20055), .A(n19671), .B(n19670), .ZN(
        P3_U2880) );
  INV_X1 U22773 ( .A(n19901), .ZN(n20032) );
  AOI22_X1 U22774 ( .A1(n20032), .A2(n19987), .B1(n20031), .B2(n19677), .ZN(
        n19673) );
  AOI22_X1 U22775 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19678), .B1(
        n19744), .B2(n20033), .ZN(n19672) );
  OAI211_X1 U22776 ( .C1(n20037), .C2(n20055), .A(n19673), .B(n19672), .ZN(
        P3_U2881) );
  AOI22_X1 U22777 ( .A1(n20039), .A2(n20040), .B1(n20038), .B2(n19677), .ZN(
        n19675) );
  AOI22_X1 U22778 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19678), .B1(
        n19744), .B2(n20041), .ZN(n19674) );
  OAI211_X1 U22779 ( .C1(n20045), .C2(n19996), .A(n19675), .B(n19674), .ZN(
        P3_U2882) );
  INV_X1 U22780 ( .A(n19676), .ZN(n19709) );
  AOI22_X1 U22781 ( .A1(n20051), .A2(n19987), .B1(n20047), .B2(n19677), .ZN(
        n19680) );
  AOI22_X1 U22782 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19678), .B1(
        n20049), .B2(n20040), .ZN(n19679) );
  OAI211_X1 U22783 ( .C1(n19709), .C2(n20056), .A(n19680), .B(n19679), .ZN(
        P3_U2883) );
  NOR2_X1 U22784 ( .A1(n12088), .A2(n19703), .ZN(n19748) );
  NAND2_X1 U22785 ( .A1(n19748), .A2(n12089), .ZN(n19764) );
  NAND2_X1 U22786 ( .A1(n19764), .A2(n19709), .ZN(n19682) );
  INV_X1 U22787 ( .A(n19682), .ZN(n19727) );
  NOR2_X1 U22788 ( .A1(n20110), .A2(n19727), .ZN(n19698) );
  AOI22_X1 U22789 ( .A1(n19998), .A2(n19723), .B1(n19997), .B2(n19698), .ZN(
        n19685) );
  INV_X1 U22790 ( .A(n19681), .ZN(n19965) );
  AOI22_X1 U22791 ( .A1(n19967), .A2(n19683), .B1(n19965), .B2(n19682), .ZN(
        n19699) );
  INV_X1 U22792 ( .A(n19764), .ZN(n19766) );
  AOI22_X1 U22793 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19699), .B1(
        n19766), .B2(n20003), .ZN(n19684) );
  OAI211_X1 U22794 ( .C1(n20006), .C2(n20055), .A(n19685), .B(n19684), .ZN(
        P3_U2884) );
  AOI22_X1 U22795 ( .A1(n19973), .A2(n19723), .B1(n20008), .B2(n19698), .ZN(
        n19687) );
  AOI22_X1 U22796 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19699), .B1(
        n19766), .B2(n20009), .ZN(n19686) );
  OAI211_X1 U22797 ( .C1(n19976), .C2(n20055), .A(n19687), .B(n19686), .ZN(
        P3_U2885) );
  AOI22_X1 U22798 ( .A1(n20013), .A2(n19698), .B1(n19946), .B2(n20040), .ZN(
        n19689) );
  AOI22_X1 U22799 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19699), .B1(
        n19766), .B2(n20015), .ZN(n19688) );
  OAI211_X1 U22800 ( .C1(n19949), .C2(n19718), .A(n19689), .B(n19688), .ZN(
        P3_U2886) );
  INV_X1 U22801 ( .A(n19953), .ZN(n20020) );
  AOI22_X1 U22802 ( .A1(n20020), .A2(n19723), .B1(n20019), .B2(n19698), .ZN(
        n19691) );
  AOI22_X1 U22803 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19699), .B1(
        n19766), .B2(n20021), .ZN(n19690) );
  OAI211_X1 U22804 ( .C1(n20024), .C2(n20055), .A(n19691), .B(n19690), .ZN(
        P3_U2887) );
  AOI22_X1 U22805 ( .A1(n20025), .A2(n19698), .B1(n19981), .B2(n20040), .ZN(
        n19693) );
  AOI22_X1 U22806 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19699), .B1(
        n19766), .B2(n20027), .ZN(n19692) );
  OAI211_X1 U22807 ( .C1(n19984), .C2(n19718), .A(n19693), .B(n19692), .ZN(
        P3_U2888) );
  AOI22_X1 U22808 ( .A1(n19898), .A2(n19723), .B1(n20031), .B2(n19698), .ZN(
        n19695) );
  AOI22_X1 U22809 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19699), .B1(
        n19766), .B2(n20033), .ZN(n19694) );
  OAI211_X1 U22810 ( .C1(n19901), .C2(n20055), .A(n19695), .B(n19694), .ZN(
        P3_U2889) );
  AOI22_X1 U22811 ( .A1(n20039), .A2(n19723), .B1(n20038), .B2(n19698), .ZN(
        n19697) );
  AOI22_X1 U22812 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19699), .B1(
        n19766), .B2(n20041), .ZN(n19696) );
  OAI211_X1 U22813 ( .C1(n20045), .C2(n20055), .A(n19697), .B(n19696), .ZN(
        P3_U2890) );
  AOI22_X1 U22814 ( .A1(n20049), .A2(n19723), .B1(n20047), .B2(n19698), .ZN(
        n19701) );
  AOI22_X1 U22815 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19699), .B1(
        n20051), .B2(n20040), .ZN(n19700) );
  OAI211_X1 U22816 ( .C1(n19764), .C2(n20056), .A(n19701), .B(n19700), .ZN(
        P3_U2891) );
  OAI211_X1 U22817 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n19967), .A(
        n19702), .B(n19999), .ZN(n19724) );
  INV_X1 U22818 ( .A(n19724), .ZN(n19721) );
  AND2_X1 U22819 ( .A1(n20102), .A2(n19748), .ZN(n19722) );
  AOI22_X1 U22820 ( .A1(n19969), .A2(n19723), .B1(n19997), .B2(n19722), .ZN(
        n19706) );
  NOR2_X2 U22821 ( .A1(n19704), .A2(n19703), .ZN(n19789) );
  AOI22_X1 U22822 ( .A1(n19998), .A2(n19744), .B1(n19789), .B2(n20003), .ZN(
        n19705) );
  OAI211_X1 U22823 ( .C1(n19721), .C2(n18714), .A(n19706), .B(n19705), .ZN(
        P3_U2892) );
  AOI22_X1 U22824 ( .A1(n20008), .A2(n19722), .B1(n20007), .B2(n19723), .ZN(
        n19708) );
  AOI22_X1 U22825 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19724), .B1(
        n19789), .B2(n20009), .ZN(n19707) );
  OAI211_X1 U22826 ( .C1(n19709), .C2(n20012), .A(n19708), .B(n19707), .ZN(
        P3_U2893) );
  INV_X1 U22827 ( .A(n19949), .ZN(n20014) );
  AOI22_X1 U22828 ( .A1(n19744), .A2(n20014), .B1(n20013), .B2(n19722), .ZN(
        n19711) );
  AOI22_X1 U22829 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19724), .B1(
        n19789), .B2(n20015), .ZN(n19710) );
  OAI211_X1 U22830 ( .C1(n20018), .C2(n19718), .A(n19711), .B(n19710), .ZN(
        P3_U2894) );
  AOI22_X1 U22831 ( .A1(n19744), .A2(n20020), .B1(n20019), .B2(n19722), .ZN(
        n19713) );
  AOI22_X1 U22832 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19724), .B1(
        n19789), .B2(n20021), .ZN(n19712) );
  OAI211_X1 U22833 ( .C1(n20024), .C2(n19718), .A(n19713), .B(n19712), .ZN(
        P3_U2895) );
  AOI22_X1 U22834 ( .A1(n19744), .A2(n20026), .B1(n20025), .B2(n19722), .ZN(
        n19715) );
  AOI22_X1 U22835 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19724), .B1(
        n19789), .B2(n20027), .ZN(n19714) );
  OAI211_X1 U22836 ( .C1(n20030), .C2(n19718), .A(n19715), .B(n19714), .ZN(
        P3_U2896) );
  AOI22_X1 U22837 ( .A1(n19744), .A2(n19898), .B1(n20031), .B2(n19722), .ZN(
        n19717) );
  AOI22_X1 U22838 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19724), .B1(
        n19789), .B2(n20033), .ZN(n19716) );
  OAI211_X1 U22839 ( .C1(n19901), .C2(n19718), .A(n19717), .B(n19716), .ZN(
        P3_U2897) );
  INV_X1 U22840 ( .A(n20045), .ZN(n19928) );
  AOI22_X1 U22841 ( .A1(n19928), .A2(n19723), .B1(n20038), .B2(n19722), .ZN(
        n19720) );
  AOI22_X1 U22842 ( .A1(n19789), .A2(n20041), .B1(n19744), .B2(n20039), .ZN(
        n19719) );
  OAI211_X1 U22843 ( .C1(n19721), .C2(n22118), .A(n19720), .B(n19719), .ZN(
        P3_U2898) );
  AOI22_X1 U22844 ( .A1(n20051), .A2(n19723), .B1(n20047), .B2(n19722), .ZN(
        n19726) );
  AOI22_X1 U22845 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19724), .B1(
        n19744), .B2(n20049), .ZN(n19725) );
  OAI211_X1 U22846 ( .C1(n19776), .C2(n20056), .A(n19726), .B(n19725), .ZN(
        P3_U2899) );
  NOR2_X2 U22847 ( .A1(n20081), .A2(n19749), .ZN(n19811) );
  AOI21_X1 U22848 ( .B1(n19807), .B2(n19776), .A(n20110), .ZN(n19743) );
  AOI22_X1 U22849 ( .A1(n19744), .A2(n19969), .B1(n19997), .B2(n19743), .ZN(
        n19730) );
  AOI221_X1 U22850 ( .B1(n19727), .B2(n19776), .C1(n19911), .C2(n19776), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n19728) );
  OAI21_X1 U22851 ( .B1(n19811), .B2(n19728), .A(n19862), .ZN(n19745) );
  AOI22_X1 U22852 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19745), .B1(
        n19811), .B2(n20003), .ZN(n19729) );
  OAI211_X1 U22853 ( .C1(n19972), .C2(n19764), .A(n19730), .B(n19729), .ZN(
        P3_U2900) );
  AOI22_X1 U22854 ( .A1(n19744), .A2(n20007), .B1(n19743), .B2(n20008), .ZN(
        n19732) );
  AOI22_X1 U22855 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19745), .B1(
        n19811), .B2(n20009), .ZN(n19731) );
  OAI211_X1 U22856 ( .C1(n19764), .C2(n20012), .A(n19732), .B(n19731), .ZN(
        P3_U2901) );
  AOI22_X1 U22857 ( .A1(n19744), .A2(n19946), .B1(n19743), .B2(n20013), .ZN(
        n19734) );
  AOI22_X1 U22858 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19745), .B1(
        n19811), .B2(n20015), .ZN(n19733) );
  OAI211_X1 U22859 ( .C1(n19764), .C2(n19949), .A(n19734), .B(n19733), .ZN(
        P3_U2902) );
  AOI22_X1 U22860 ( .A1(n19744), .A2(n19950), .B1(n19743), .B2(n20019), .ZN(
        n19736) );
  AOI22_X1 U22861 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19745), .B1(
        n19811), .B2(n20021), .ZN(n19735) );
  OAI211_X1 U22862 ( .C1(n19764), .C2(n19953), .A(n19736), .B(n19735), .ZN(
        P3_U2903) );
  AOI22_X1 U22863 ( .A1(n19744), .A2(n19981), .B1(n19743), .B2(n20025), .ZN(
        n19738) );
  AOI22_X1 U22864 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19745), .B1(
        n19811), .B2(n20027), .ZN(n19737) );
  OAI211_X1 U22865 ( .C1(n19764), .C2(n19984), .A(n19738), .B(n19737), .ZN(
        P3_U2904) );
  AOI22_X1 U22866 ( .A1(n19744), .A2(n20032), .B1(n19743), .B2(n20031), .ZN(
        n19740) );
  AOI22_X1 U22867 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19745), .B1(
        n19811), .B2(n20033), .ZN(n19739) );
  OAI211_X1 U22868 ( .C1(n19764), .C2(n20037), .A(n19740), .B(n19739), .ZN(
        P3_U2905) );
  INV_X1 U22869 ( .A(n20039), .ZN(n19931) );
  AOI22_X1 U22870 ( .A1(n19744), .A2(n19928), .B1(n19743), .B2(n20038), .ZN(
        n19742) );
  AOI22_X1 U22871 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19745), .B1(
        n19811), .B2(n20041), .ZN(n19741) );
  OAI211_X1 U22872 ( .C1(n19764), .C2(n19931), .A(n19742), .B(n19741), .ZN(
        P3_U2906) );
  AOI22_X1 U22873 ( .A1(n19766), .A2(n20049), .B1(n19743), .B2(n20047), .ZN(
        n19747) );
  AOI22_X1 U22874 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19745), .B1(
        n19744), .B2(n20051), .ZN(n19746) );
  OAI211_X1 U22875 ( .C1(n19807), .C2(n20056), .A(n19747), .B(n19746), .ZN(
        P3_U2907) );
  NOR2_X1 U22876 ( .A1(n19749), .A2(n19937), .ZN(n19765) );
  AOI22_X1 U22877 ( .A1(n19766), .A2(n19969), .B1(n19997), .B2(n19765), .ZN(
        n19751) );
  AOI22_X1 U22878 ( .A1(n20002), .A2(n19748), .B1(n19794), .B2(n19939), .ZN(
        n19767) );
  NOR2_X2 U22879 ( .A1(n19749), .A2(n19841), .ZN(n19835) );
  AOI22_X1 U22880 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19767), .B1(
        n20003), .B2(n19835), .ZN(n19750) );
  OAI211_X1 U22881 ( .C1(n19972), .C2(n19776), .A(n19751), .B(n19750), .ZN(
        P3_U2908) );
  AOI22_X1 U22882 ( .A1(n19789), .A2(n19973), .B1(n20008), .B2(n19765), .ZN(
        n19753) );
  AOI22_X1 U22883 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19767), .B1(
        n20009), .B2(n19835), .ZN(n19752) );
  OAI211_X1 U22884 ( .C1(n19764), .C2(n19976), .A(n19753), .B(n19752), .ZN(
        P3_U2909) );
  AOI22_X1 U22885 ( .A1(n19789), .A2(n20014), .B1(n20013), .B2(n19765), .ZN(
        n19755) );
  AOI22_X1 U22886 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19767), .B1(
        n20015), .B2(n19835), .ZN(n19754) );
  OAI211_X1 U22887 ( .C1(n19764), .C2(n20018), .A(n19755), .B(n19754), .ZN(
        P3_U2910) );
  AOI22_X1 U22888 ( .A1(n19789), .A2(n20020), .B1(n20019), .B2(n19765), .ZN(
        n19757) );
  AOI22_X1 U22889 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19767), .B1(
        n20021), .B2(n19835), .ZN(n19756) );
  OAI211_X1 U22890 ( .C1(n19764), .C2(n20024), .A(n19757), .B(n19756), .ZN(
        P3_U2911) );
  AOI22_X1 U22891 ( .A1(n19789), .A2(n20026), .B1(n20025), .B2(n19765), .ZN(
        n19759) );
  AOI22_X1 U22892 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19767), .B1(
        n20027), .B2(n19835), .ZN(n19758) );
  OAI211_X1 U22893 ( .C1(n19764), .C2(n20030), .A(n19759), .B(n19758), .ZN(
        P3_U2912) );
  AOI22_X1 U22894 ( .A1(n19789), .A2(n19898), .B1(n20031), .B2(n19765), .ZN(
        n19761) );
  AOI22_X1 U22895 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19767), .B1(
        n20033), .B2(n19835), .ZN(n19760) );
  OAI211_X1 U22896 ( .C1(n19764), .C2(n19901), .A(n19761), .B(n19760), .ZN(
        P3_U2913) );
  AOI22_X1 U22897 ( .A1(n19789), .A2(n20039), .B1(n20038), .B2(n19765), .ZN(
        n19763) );
  AOI22_X1 U22898 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19767), .B1(
        n20041), .B2(n19835), .ZN(n19762) );
  OAI211_X1 U22899 ( .C1(n19764), .C2(n20045), .A(n19763), .B(n19762), .ZN(
        P3_U2914) );
  AOI22_X1 U22900 ( .A1(n19766), .A2(n20051), .B1(n20047), .B2(n19765), .ZN(
        n19769) );
  AOI22_X1 U22901 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19767), .B1(
        n19789), .B2(n20049), .ZN(n19768) );
  OAI211_X1 U22902 ( .C1(n20056), .C2(n19833), .A(n19769), .B(n19768), .ZN(
        P3_U2915) );
  OR3_X1 U22903 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n19839), .ZN(n19846) );
  NAND2_X1 U22904 ( .A1(n19833), .A2(n19846), .ZN(n19771) );
  INV_X1 U22905 ( .A(n19771), .ZN(n19815) );
  NOR2_X1 U22906 ( .A1(n20110), .A2(n19815), .ZN(n19787) );
  AOI22_X1 U22907 ( .A1(n19998), .A2(n19811), .B1(n19997), .B2(n19787), .ZN(
        n19773) );
  NAND2_X1 U22908 ( .A1(n19807), .A2(n19776), .ZN(n19770) );
  OAI221_X1 U22909 ( .B1(n19771), .B2(n19967), .C1(n19771), .C2(n19770), .A(
        n19965), .ZN(n19788) );
  INV_X1 U22910 ( .A(n19846), .ZN(n19853) );
  AOI22_X1 U22911 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19788), .B1(
        n20003), .B2(n19853), .ZN(n19772) );
  OAI211_X1 U22912 ( .C1(n19776), .C2(n20006), .A(n19773), .B(n19772), .ZN(
        P3_U2916) );
  AOI22_X1 U22913 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19788), .B1(
        n20008), .B2(n19787), .ZN(n19775) );
  AOI22_X1 U22914 ( .A1(n19811), .A2(n19973), .B1(n20009), .B2(n19853), .ZN(
        n19774) );
  OAI211_X1 U22915 ( .C1(n19776), .C2(n19976), .A(n19775), .B(n19774), .ZN(
        P3_U2917) );
  AOI22_X1 U22916 ( .A1(n19789), .A2(n19946), .B1(n20013), .B2(n19787), .ZN(
        n19778) );
  AOI22_X1 U22917 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19788), .B1(
        n20015), .B2(n19853), .ZN(n19777) );
  OAI211_X1 U22918 ( .C1(n19807), .C2(n19949), .A(n19778), .B(n19777), .ZN(
        P3_U2918) );
  AOI22_X1 U22919 ( .A1(n19789), .A2(n19950), .B1(n20019), .B2(n19787), .ZN(
        n19780) );
  AOI22_X1 U22920 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19788), .B1(
        n20021), .B2(n19853), .ZN(n19779) );
  OAI211_X1 U22921 ( .C1(n19807), .C2(n19953), .A(n19780), .B(n19779), .ZN(
        P3_U2919) );
  AOI22_X1 U22922 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19788), .B1(
        n20025), .B2(n19787), .ZN(n19782) );
  AOI22_X1 U22923 ( .A1(n19789), .A2(n19981), .B1(n20027), .B2(n19853), .ZN(
        n19781) );
  OAI211_X1 U22924 ( .C1(n19807), .C2(n19984), .A(n19782), .B(n19781), .ZN(
        P3_U2920) );
  AOI22_X1 U22925 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19788), .B1(
        n20031), .B2(n19787), .ZN(n19784) );
  AOI22_X1 U22926 ( .A1(n19789), .A2(n20032), .B1(n20033), .B2(n19853), .ZN(
        n19783) );
  OAI211_X1 U22927 ( .C1(n19807), .C2(n20037), .A(n19784), .B(n19783), .ZN(
        P3_U2921) );
  AOI22_X1 U22928 ( .A1(n19789), .A2(n19928), .B1(n20038), .B2(n19787), .ZN(
        n19786) );
  AOI22_X1 U22929 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19788), .B1(
        n20041), .B2(n19853), .ZN(n19785) );
  OAI211_X1 U22930 ( .C1(n19807), .C2(n19931), .A(n19786), .B(n19785), .ZN(
        P3_U2922) );
  AOI22_X1 U22931 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19788), .B1(
        n20047), .B2(n19787), .ZN(n19791) );
  AOI22_X1 U22932 ( .A1(n19811), .A2(n20049), .B1(n19789), .B2(n20051), .ZN(
        n19790) );
  OAI211_X1 U22933 ( .C1(n20056), .C2(n19846), .A(n19791), .B(n19790), .ZN(
        P3_U2923) );
  AOI22_X1 U22934 ( .A1(n19998), .A2(n19835), .B1(n19997), .B2(n19810), .ZN(
        n19796) );
  AOI21_X1 U22935 ( .B1(n12088), .B2(n19911), .A(n19792), .ZN(n19793) );
  NAND2_X1 U22936 ( .A1(n19794), .A2(n19793), .ZN(n19812) );
  NAND2_X1 U22937 ( .A1(n20075), .A2(n19794), .ZN(n19880) );
  AOI22_X1 U22938 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19812), .B1(
        n20003), .B2(n19882), .ZN(n19795) );
  OAI211_X1 U22939 ( .C1(n19807), .C2(n20006), .A(n19796), .B(n19795), .ZN(
        P3_U2924) );
  AOI22_X1 U22940 ( .A1(n19973), .A2(n19835), .B1(n20008), .B2(n19810), .ZN(
        n19798) );
  AOI22_X1 U22941 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19812), .B1(
        n20009), .B2(n19882), .ZN(n19797) );
  OAI211_X1 U22942 ( .C1(n19807), .C2(n19976), .A(n19798), .B(n19797), .ZN(
        P3_U2925) );
  AOI22_X1 U22943 ( .A1(n19811), .A2(n19946), .B1(n20013), .B2(n19810), .ZN(
        n19800) );
  AOI22_X1 U22944 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19812), .B1(
        n20015), .B2(n19882), .ZN(n19799) );
  OAI211_X1 U22945 ( .C1(n19949), .C2(n19833), .A(n19800), .B(n19799), .ZN(
        P3_U2926) );
  AOI22_X1 U22946 ( .A1(n20020), .A2(n19835), .B1(n20019), .B2(n19810), .ZN(
        n19802) );
  AOI22_X1 U22947 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19812), .B1(
        n20021), .B2(n19882), .ZN(n19801) );
  OAI211_X1 U22948 ( .C1(n19807), .C2(n20024), .A(n19802), .B(n19801), .ZN(
        P3_U2927) );
  AOI22_X1 U22949 ( .A1(n20026), .A2(n19835), .B1(n20025), .B2(n19810), .ZN(
        n19804) );
  AOI22_X1 U22950 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19812), .B1(
        n20027), .B2(n19882), .ZN(n19803) );
  OAI211_X1 U22951 ( .C1(n19807), .C2(n20030), .A(n19804), .B(n19803), .ZN(
        P3_U2928) );
  AOI22_X1 U22952 ( .A1(n19898), .A2(n19835), .B1(n20031), .B2(n19810), .ZN(
        n19806) );
  AOI22_X1 U22953 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19812), .B1(
        n20033), .B2(n19882), .ZN(n19805) );
  OAI211_X1 U22954 ( .C1(n19807), .C2(n19901), .A(n19806), .B(n19805), .ZN(
        P3_U2929) );
  AOI22_X1 U22955 ( .A1(n19811), .A2(n19928), .B1(n20038), .B2(n19810), .ZN(
        n19809) );
  AOI22_X1 U22956 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19812), .B1(
        n20041), .B2(n19882), .ZN(n19808) );
  OAI211_X1 U22957 ( .C1(n19931), .C2(n19833), .A(n19809), .B(n19808), .ZN(
        P3_U2930) );
  AOI22_X1 U22958 ( .A1(n19811), .A2(n20051), .B1(n20047), .B2(n19810), .ZN(
        n19814) );
  AOI22_X1 U22959 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19812), .B1(
        n20049), .B2(n19835), .ZN(n19813) );
  OAI211_X1 U22960 ( .C1(n20056), .C2(n19880), .A(n19814), .B(n19813), .ZN(
        P3_U2931) );
  NOR2_X2 U22961 ( .A1(n20081), .A2(n19861), .ZN(n19906) );
  NOR2_X1 U22962 ( .A1(n19882), .A2(n19906), .ZN(n19864) );
  OAI21_X1 U22963 ( .B1(n19911), .B2(n19815), .A(n19864), .ZN(n19816) );
  OAI211_X1 U22964 ( .C1(n21986), .C2(n19906), .A(n19816), .B(n19862), .ZN(
        n19836) );
  INV_X1 U22965 ( .A(n19836), .ZN(n19826) );
  NOR2_X1 U22966 ( .A1(n20110), .A2(n19864), .ZN(n19834) );
  AOI22_X1 U22967 ( .A1(n19998), .A2(n19853), .B1(n19997), .B2(n19834), .ZN(
        n19818) );
  AOI22_X1 U22968 ( .A1(n20003), .A2(n19906), .B1(n19969), .B2(n19835), .ZN(
        n19817) );
  OAI211_X1 U22969 ( .C1(n19826), .C2(n19819), .A(n19818), .B(n19817), .ZN(
        P3_U2932) );
  AOI22_X1 U22970 ( .A1(n19973), .A2(n19853), .B1(n20008), .B2(n19834), .ZN(
        n19821) );
  AOI22_X1 U22971 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19836), .B1(
        n20009), .B2(n19906), .ZN(n19820) );
  OAI211_X1 U22972 ( .C1(n19976), .C2(n19833), .A(n19821), .B(n19820), .ZN(
        P3_U2933) );
  AOI22_X1 U22973 ( .A1(n20014), .A2(n19853), .B1(n20013), .B2(n19834), .ZN(
        n19823) );
  AOI22_X1 U22974 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19836), .B1(
        n20015), .B2(n19906), .ZN(n19822) );
  OAI211_X1 U22975 ( .C1(n20018), .C2(n19833), .A(n19823), .B(n19822), .ZN(
        P3_U2934) );
  AOI22_X1 U22976 ( .A1(n20020), .A2(n19853), .B1(n20019), .B2(n19834), .ZN(
        n19825) );
  AOI22_X1 U22977 ( .A1(n20021), .A2(n19906), .B1(n19950), .B2(n19835), .ZN(
        n19824) );
  OAI211_X1 U22978 ( .C1(n19826), .C2(n13897), .A(n19825), .B(n19824), .ZN(
        P3_U2935) );
  AOI22_X1 U22979 ( .A1(n20025), .A2(n19834), .B1(n19981), .B2(n19835), .ZN(
        n19828) );
  AOI22_X1 U22980 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19836), .B1(
        n20027), .B2(n19906), .ZN(n19827) );
  OAI211_X1 U22981 ( .C1(n19984), .C2(n19846), .A(n19828), .B(n19827), .ZN(
        P3_U2936) );
  AOI22_X1 U22982 ( .A1(n20032), .A2(n19835), .B1(n20031), .B2(n19834), .ZN(
        n19830) );
  AOI22_X1 U22983 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19836), .B1(
        n20033), .B2(n19906), .ZN(n19829) );
  OAI211_X1 U22984 ( .C1(n20037), .C2(n19846), .A(n19830), .B(n19829), .ZN(
        P3_U2937) );
  AOI22_X1 U22985 ( .A1(n20039), .A2(n19853), .B1(n20038), .B2(n19834), .ZN(
        n19832) );
  AOI22_X1 U22986 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19836), .B1(
        n20041), .B2(n19906), .ZN(n19831) );
  OAI211_X1 U22987 ( .C1(n20045), .C2(n19833), .A(n19832), .B(n19831), .ZN(
        P3_U2938) );
  INV_X1 U22988 ( .A(n19906), .ZN(n19904) );
  AOI22_X1 U22989 ( .A1(n20049), .A2(n19853), .B1(n20047), .B2(n19834), .ZN(
        n19838) );
  AOI22_X1 U22990 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19836), .B1(
        n20051), .B2(n19835), .ZN(n19837) );
  OAI211_X1 U22991 ( .C1(n20056), .C2(n19904), .A(n19838), .B(n19837), .ZN(
        P3_U2939) );
  NOR2_X1 U22992 ( .A1(n19861), .A2(n19937), .ZN(n19886) );
  AOI22_X1 U22993 ( .A1(n19969), .A2(n19853), .B1(n19997), .B2(n19886), .ZN(
        n19843) );
  NOR2_X1 U22994 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19839), .ZN(
        n19840) );
  AOI22_X1 U22995 ( .A1(n20002), .A2(n19840), .B1(n19887), .B2(n19939), .ZN(
        n19858) );
  AOI22_X1 U22996 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19858), .B1(
        n20003), .B2(n19933), .ZN(n19842) );
  OAI211_X1 U22997 ( .C1(n19972), .C2(n19880), .A(n19843), .B(n19842), .ZN(
        P3_U2940) );
  AOI22_X1 U22998 ( .A1(n19973), .A2(n19882), .B1(n20008), .B2(n19886), .ZN(
        n19845) );
  AOI22_X1 U22999 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19858), .B1(
        n20009), .B2(n19933), .ZN(n19844) );
  OAI211_X1 U23000 ( .C1(n19976), .C2(n19846), .A(n19845), .B(n19844), .ZN(
        P3_U2941) );
  AOI22_X1 U23001 ( .A1(n20013), .A2(n19886), .B1(n19946), .B2(n19853), .ZN(
        n19848) );
  AOI22_X1 U23002 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19858), .B1(
        n20015), .B2(n19933), .ZN(n19847) );
  OAI211_X1 U23003 ( .C1(n19949), .C2(n19880), .A(n19848), .B(n19847), .ZN(
        P3_U2942) );
  AOI22_X1 U23004 ( .A1(n19950), .A2(n19853), .B1(n20019), .B2(n19886), .ZN(
        n19850) );
  AOI22_X1 U23005 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19858), .B1(
        n20021), .B2(n19933), .ZN(n19849) );
  OAI211_X1 U23006 ( .C1(n19953), .C2(n19880), .A(n19850), .B(n19849), .ZN(
        P3_U2943) );
  AOI22_X1 U23007 ( .A1(n20025), .A2(n19886), .B1(n19981), .B2(n19853), .ZN(
        n19852) );
  AOI22_X1 U23008 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19858), .B1(
        n20027), .B2(n19933), .ZN(n19851) );
  OAI211_X1 U23009 ( .C1(n19984), .C2(n19880), .A(n19852), .B(n19851), .ZN(
        P3_U2944) );
  AOI22_X1 U23010 ( .A1(n20032), .A2(n19853), .B1(n20031), .B2(n19886), .ZN(
        n19855) );
  AOI22_X1 U23011 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19858), .B1(
        n20033), .B2(n19933), .ZN(n19854) );
  OAI211_X1 U23012 ( .C1(n20037), .C2(n19880), .A(n19855), .B(n19854), .ZN(
        P3_U2945) );
  AOI22_X1 U23013 ( .A1(n19928), .A2(n19853), .B1(n20038), .B2(n19886), .ZN(
        n19857) );
  AOI22_X1 U23014 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19858), .B1(
        n20041), .B2(n19933), .ZN(n19856) );
  OAI211_X1 U23015 ( .C1(n19931), .C2(n19880), .A(n19857), .B(n19856), .ZN(
        P3_U2946) );
  INV_X1 U23016 ( .A(n19933), .ZN(n19923) );
  AOI22_X1 U23017 ( .A1(n20051), .A2(n19853), .B1(n20047), .B2(n19886), .ZN(
        n19860) );
  AOI22_X1 U23018 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19858), .B1(
        n20049), .B2(n19882), .ZN(n19859) );
  OAI211_X1 U23019 ( .C1(n20056), .C2(n19923), .A(n19860), .B(n19859), .ZN(
        P3_U2947) );
  NOR2_X1 U23020 ( .A1(n12088), .A2(n19861), .ZN(n19941) );
  NAND2_X1 U23021 ( .A1(n19941), .A2(n12089), .ZN(n19960) );
  AOI21_X1 U23022 ( .B1(n19923), .B2(n19960), .A(n20110), .ZN(n19881) );
  AOI22_X1 U23023 ( .A1(n19998), .A2(n19906), .B1(n19997), .B2(n19881), .ZN(
        n19867) );
  INV_X1 U23024 ( .A(n19960), .ZN(n19961) );
  OAI21_X1 U23025 ( .B1(n19933), .B2(n19961), .A(n19862), .ZN(n19910) );
  OAI21_X1 U23026 ( .B1(n19864), .B2(n19863), .A(n19910), .ZN(n19865) );
  OAI21_X1 U23027 ( .B1(n19961), .B2(n21986), .A(n19865), .ZN(n19883) );
  AOI22_X1 U23028 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19883), .B1(
        n20003), .B2(n19961), .ZN(n19866) );
  OAI211_X1 U23029 ( .C1(n20006), .C2(n19880), .A(n19867), .B(n19866), .ZN(
        P3_U2948) );
  AOI22_X1 U23030 ( .A1(n20008), .A2(n19881), .B1(n20007), .B2(n19882), .ZN(
        n19869) );
  AOI22_X1 U23031 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19883), .B1(
        n20009), .B2(n19961), .ZN(n19868) );
  OAI211_X1 U23032 ( .C1(n20012), .C2(n19904), .A(n19869), .B(n19868), .ZN(
        P3_U2949) );
  AOI22_X1 U23033 ( .A1(n20014), .A2(n19906), .B1(n20013), .B2(n19881), .ZN(
        n19871) );
  AOI22_X1 U23034 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19883), .B1(
        n20015), .B2(n19961), .ZN(n19870) );
  OAI211_X1 U23035 ( .C1(n20018), .C2(n19880), .A(n19871), .B(n19870), .ZN(
        P3_U2950) );
  AOI22_X1 U23036 ( .A1(n19950), .A2(n19882), .B1(n20019), .B2(n19881), .ZN(
        n19873) );
  AOI22_X1 U23037 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19883), .B1(
        n20021), .B2(n19961), .ZN(n19872) );
  OAI211_X1 U23038 ( .C1(n19953), .C2(n19904), .A(n19873), .B(n19872), .ZN(
        P3_U2951) );
  AOI22_X1 U23039 ( .A1(n20026), .A2(n19906), .B1(n20025), .B2(n19881), .ZN(
        n19875) );
  AOI22_X1 U23040 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19883), .B1(
        n20027), .B2(n19961), .ZN(n19874) );
  OAI211_X1 U23041 ( .C1(n20030), .C2(n19880), .A(n19875), .B(n19874), .ZN(
        P3_U2952) );
  AOI22_X1 U23042 ( .A1(n19898), .A2(n19906), .B1(n20031), .B2(n19881), .ZN(
        n19877) );
  AOI22_X1 U23043 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19883), .B1(
        n20033), .B2(n19961), .ZN(n19876) );
  OAI211_X1 U23044 ( .C1(n19901), .C2(n19880), .A(n19877), .B(n19876), .ZN(
        P3_U2953) );
  AOI22_X1 U23045 ( .A1(n20039), .A2(n19906), .B1(n20038), .B2(n19881), .ZN(
        n19879) );
  AOI22_X1 U23046 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19883), .B1(
        n20041), .B2(n19961), .ZN(n19878) );
  OAI211_X1 U23047 ( .C1(n20045), .C2(n19880), .A(n19879), .B(n19878), .ZN(
        P3_U2954) );
  AOI22_X1 U23048 ( .A1(n20051), .A2(n19882), .B1(n20047), .B2(n19881), .ZN(
        n19885) );
  AOI22_X1 U23049 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19883), .B1(
        n20049), .B2(n19906), .ZN(n19884) );
  OAI211_X1 U23050 ( .C1(n20056), .C2(n19960), .A(n19885), .B(n19884), .ZN(
        P3_U2955) );
  AND2_X1 U23051 ( .A1(n20102), .A2(n19941), .ZN(n19905) );
  AOI22_X1 U23052 ( .A1(n19998), .A2(n19933), .B1(n19997), .B2(n19905), .ZN(
        n19889) );
  AOI22_X1 U23053 ( .A1(n20002), .A2(n19886), .B1(n19999), .B2(n19941), .ZN(
        n19907) );
  NAND2_X1 U23054 ( .A1(n20075), .A2(n19887), .ZN(n19990) );
  INV_X1 U23055 ( .A(n19990), .ZN(n19993) );
  AOI22_X1 U23056 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19907), .B1(
        n20003), .B2(n19993), .ZN(n19888) );
  OAI211_X1 U23057 ( .C1(n20006), .C2(n19904), .A(n19889), .B(n19888), .ZN(
        P3_U2956) );
  AOI22_X1 U23058 ( .A1(n20008), .A2(n19905), .B1(n20007), .B2(n19906), .ZN(
        n19891) );
  AOI22_X1 U23059 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19907), .B1(
        n20009), .B2(n19993), .ZN(n19890) );
  OAI211_X1 U23060 ( .C1(n20012), .C2(n19923), .A(n19891), .B(n19890), .ZN(
        P3_U2957) );
  AOI22_X1 U23061 ( .A1(n20013), .A2(n19905), .B1(n19946), .B2(n19906), .ZN(
        n19893) );
  AOI22_X1 U23062 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19907), .B1(
        n20015), .B2(n19993), .ZN(n19892) );
  OAI211_X1 U23063 ( .C1(n19949), .C2(n19923), .A(n19893), .B(n19892), .ZN(
        P3_U2958) );
  AOI22_X1 U23064 ( .A1(n20020), .A2(n19933), .B1(n20019), .B2(n19905), .ZN(
        n19895) );
  AOI22_X1 U23065 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19907), .B1(
        n20021), .B2(n19993), .ZN(n19894) );
  OAI211_X1 U23066 ( .C1(n20024), .C2(n19904), .A(n19895), .B(n19894), .ZN(
        P3_U2959) );
  AOI22_X1 U23067 ( .A1(n20026), .A2(n19933), .B1(n20025), .B2(n19905), .ZN(
        n19897) );
  AOI22_X1 U23068 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19907), .B1(
        n20027), .B2(n19993), .ZN(n19896) );
  OAI211_X1 U23069 ( .C1(n20030), .C2(n19904), .A(n19897), .B(n19896), .ZN(
        P3_U2960) );
  AOI22_X1 U23070 ( .A1(n19898), .A2(n19933), .B1(n20031), .B2(n19905), .ZN(
        n19900) );
  AOI22_X1 U23071 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19907), .B1(
        n20033), .B2(n19993), .ZN(n19899) );
  OAI211_X1 U23072 ( .C1(n19901), .C2(n19904), .A(n19900), .B(n19899), .ZN(
        P3_U2961) );
  AOI22_X1 U23073 ( .A1(n20039), .A2(n19933), .B1(n20038), .B2(n19905), .ZN(
        n19903) );
  AOI22_X1 U23074 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19907), .B1(
        n20041), .B2(n19993), .ZN(n19902) );
  OAI211_X1 U23075 ( .C1(n20045), .C2(n19904), .A(n19903), .B(n19902), .ZN(
        P3_U2962) );
  AOI22_X1 U23076 ( .A1(n20049), .A2(n19933), .B1(n20047), .B2(n19905), .ZN(
        n19909) );
  AOI22_X1 U23077 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19907), .B1(
        n20051), .B2(n19906), .ZN(n19908) );
  OAI211_X1 U23078 ( .C1(n20056), .C2(n19990), .A(n19909), .B(n19908), .ZN(
        P3_U2963) );
  NOR2_X2 U23079 ( .A1(n20081), .A2(n19938), .ZN(n20050) );
  INV_X1 U23080 ( .A(n20050), .ZN(n20044) );
  NAND2_X1 U23081 ( .A1(n19990), .A2(n20044), .ZN(n19966) );
  INV_X1 U23082 ( .A(n19966), .ZN(n19913) );
  NOR2_X1 U23083 ( .A1(n20110), .A2(n19913), .ZN(n19932) );
  AOI22_X1 U23084 ( .A1(n19969), .A2(n19933), .B1(n19997), .B2(n19932), .ZN(
        n19916) );
  OAI22_X1 U23085 ( .A1(n19913), .A2(n19912), .B1(n19911), .B2(n19910), .ZN(
        n19914) );
  OAI21_X1 U23086 ( .B1(n20050), .B2(n21986), .A(n19914), .ZN(n19934) );
  AOI22_X1 U23087 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19934), .B1(
        n20003), .B2(n20050), .ZN(n19915) );
  OAI211_X1 U23088 ( .C1(n19972), .C2(n19960), .A(n19916), .B(n19915), .ZN(
        P3_U2964) );
  AOI22_X1 U23089 ( .A1(n20008), .A2(n19932), .B1(n20007), .B2(n19933), .ZN(
        n19918) );
  AOI22_X1 U23090 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19934), .B1(
        n20009), .B2(n20050), .ZN(n19917) );
  OAI211_X1 U23091 ( .C1(n20012), .C2(n19960), .A(n19918), .B(n19917), .ZN(
        P3_U2965) );
  AOI22_X1 U23092 ( .A1(n20013), .A2(n19932), .B1(n19946), .B2(n19933), .ZN(
        n19920) );
  AOI22_X1 U23093 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19934), .B1(
        n20015), .B2(n20050), .ZN(n19919) );
  OAI211_X1 U23094 ( .C1(n19949), .C2(n19960), .A(n19920), .B(n19919), .ZN(
        P3_U2966) );
  AOI22_X1 U23095 ( .A1(n20020), .A2(n19961), .B1(n20019), .B2(n19932), .ZN(
        n19922) );
  AOI22_X1 U23096 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19934), .B1(
        n20021), .B2(n20050), .ZN(n19921) );
  OAI211_X1 U23097 ( .C1(n20024), .C2(n19923), .A(n19922), .B(n19921), .ZN(
        P3_U2967) );
  AOI22_X1 U23098 ( .A1(n20025), .A2(n19932), .B1(n19981), .B2(n19933), .ZN(
        n19925) );
  AOI22_X1 U23099 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19934), .B1(
        n20027), .B2(n20050), .ZN(n19924) );
  OAI211_X1 U23100 ( .C1(n19984), .C2(n19960), .A(n19925), .B(n19924), .ZN(
        P3_U2968) );
  AOI22_X1 U23101 ( .A1(n20032), .A2(n19933), .B1(n20031), .B2(n19932), .ZN(
        n19927) );
  AOI22_X1 U23102 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19934), .B1(
        n20033), .B2(n20050), .ZN(n19926) );
  OAI211_X1 U23103 ( .C1(n20037), .C2(n19960), .A(n19927), .B(n19926), .ZN(
        P3_U2969) );
  AOI22_X1 U23104 ( .A1(n19928), .A2(n19933), .B1(n20038), .B2(n19932), .ZN(
        n19930) );
  AOI22_X1 U23105 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19934), .B1(
        n20041), .B2(n20050), .ZN(n19929) );
  OAI211_X1 U23106 ( .C1(n19931), .C2(n19960), .A(n19930), .B(n19929), .ZN(
        P3_U2970) );
  AOI22_X1 U23107 ( .A1(n20049), .A2(n19961), .B1(n20047), .B2(n19932), .ZN(
        n19936) );
  AOI22_X1 U23108 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19934), .B1(
        n20051), .B2(n19933), .ZN(n19935) );
  OAI211_X1 U23109 ( .C1(n20056), .C2(n20044), .A(n19936), .B(n19935), .ZN(
        P3_U2971) );
  NOR2_X1 U23110 ( .A1(n19938), .A2(n19937), .ZN(n20001) );
  AOI22_X1 U23111 ( .A1(n19969), .A2(n19961), .B1(n19997), .B2(n20001), .ZN(
        n19943) );
  AOI22_X1 U23112 ( .A1(n20002), .A2(n19941), .B1(n19940), .B2(n19939), .ZN(
        n19962) );
  AOI22_X1 U23113 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19962), .B1(
        n20003), .B2(n20048), .ZN(n19942) );
  OAI211_X1 U23114 ( .C1(n19972), .C2(n19990), .A(n19943), .B(n19942), .ZN(
        P3_U2972) );
  AOI22_X1 U23115 ( .A1(n20008), .A2(n20001), .B1(n20007), .B2(n19961), .ZN(
        n19945) );
  AOI22_X1 U23116 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19962), .B1(
        n20009), .B2(n20048), .ZN(n19944) );
  OAI211_X1 U23117 ( .C1(n20012), .C2(n19990), .A(n19945), .B(n19944), .ZN(
        P3_U2973) );
  AOI22_X1 U23118 ( .A1(n20013), .A2(n20001), .B1(n19946), .B2(n19961), .ZN(
        n19948) );
  AOI22_X1 U23119 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19962), .B1(
        n20015), .B2(n20048), .ZN(n19947) );
  OAI211_X1 U23120 ( .C1(n19949), .C2(n19990), .A(n19948), .B(n19947), .ZN(
        P3_U2974) );
  AOI22_X1 U23121 ( .A1(n19950), .A2(n19961), .B1(n20019), .B2(n20001), .ZN(
        n19952) );
  AOI22_X1 U23122 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19962), .B1(
        n20021), .B2(n20048), .ZN(n19951) );
  OAI211_X1 U23123 ( .C1(n19953), .C2(n19990), .A(n19952), .B(n19951), .ZN(
        P3_U2975) );
  AOI22_X1 U23124 ( .A1(n20026), .A2(n19993), .B1(n20025), .B2(n20001), .ZN(
        n19955) );
  AOI22_X1 U23125 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19962), .B1(
        n20027), .B2(n20048), .ZN(n19954) );
  OAI211_X1 U23126 ( .C1(n20030), .C2(n19960), .A(n19955), .B(n19954), .ZN(
        P3_U2976) );
  AOI22_X1 U23127 ( .A1(n20032), .A2(n19961), .B1(n20031), .B2(n20001), .ZN(
        n19957) );
  AOI22_X1 U23128 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19962), .B1(
        n20033), .B2(n20048), .ZN(n19956) );
  OAI211_X1 U23129 ( .C1(n20037), .C2(n19990), .A(n19957), .B(n19956), .ZN(
        P3_U2977) );
  AOI22_X1 U23130 ( .A1(n20039), .A2(n19993), .B1(n20038), .B2(n20001), .ZN(
        n19959) );
  AOI22_X1 U23131 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19962), .B1(
        n20041), .B2(n20048), .ZN(n19958) );
  OAI211_X1 U23132 ( .C1(n20045), .C2(n19960), .A(n19959), .B(n19958), .ZN(
        P3_U2978) );
  AOI22_X1 U23133 ( .A1(n20049), .A2(n19993), .B1(n20047), .B2(n20001), .ZN(
        n19964) );
  AOI22_X1 U23134 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19962), .B1(
        n20051), .B2(n19961), .ZN(n19963) );
  OAI211_X1 U23135 ( .C1(n20056), .C2(n20036), .A(n19964), .B(n19963), .ZN(
        P3_U2979) );
  OAI221_X1 U23136 ( .B1(n19968), .B2(n19967), .C1(n19968), .C2(n19966), .A(
        n19965), .ZN(n19992) );
  AND2_X1 U23137 ( .A1(n20102), .A2(n19968), .ZN(n19991) );
  AOI22_X1 U23138 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19992), .B1(
        n19997), .B2(n19991), .ZN(n19971) );
  AOI22_X1 U23139 ( .A1(n20003), .A2(n19987), .B1(n19969), .B2(n19993), .ZN(
        n19970) );
  OAI211_X1 U23140 ( .C1(n19972), .C2(n20044), .A(n19971), .B(n19970), .ZN(
        P3_U2980) );
  AOI22_X1 U23141 ( .A1(n19973), .A2(n20050), .B1(n20008), .B2(n19991), .ZN(
        n19975) );
  AOI22_X1 U23142 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19992), .B1(
        n20009), .B2(n19987), .ZN(n19974) );
  OAI211_X1 U23143 ( .C1(n19976), .C2(n19990), .A(n19975), .B(n19974), .ZN(
        P3_U2981) );
  AOI22_X1 U23144 ( .A1(n20014), .A2(n20050), .B1(n20013), .B2(n19991), .ZN(
        n19978) );
  AOI22_X1 U23145 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19992), .B1(
        n20015), .B2(n19987), .ZN(n19977) );
  OAI211_X1 U23146 ( .C1(n20018), .C2(n19990), .A(n19978), .B(n19977), .ZN(
        P3_U2982) );
  AOI22_X1 U23147 ( .A1(n20020), .A2(n20050), .B1(n20019), .B2(n19991), .ZN(
        n19980) );
  AOI22_X1 U23148 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19992), .B1(
        n20021), .B2(n19987), .ZN(n19979) );
  OAI211_X1 U23149 ( .C1(n20024), .C2(n19990), .A(n19980), .B(n19979), .ZN(
        P3_U2983) );
  AOI22_X1 U23150 ( .A1(n20025), .A2(n19991), .B1(n19981), .B2(n19993), .ZN(
        n19983) );
  AOI22_X1 U23151 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19992), .B1(
        n20027), .B2(n19987), .ZN(n19982) );
  OAI211_X1 U23152 ( .C1(n19984), .C2(n20044), .A(n19983), .B(n19982), .ZN(
        P3_U2984) );
  AOI22_X1 U23153 ( .A1(n20032), .A2(n19993), .B1(n20031), .B2(n19991), .ZN(
        n19986) );
  AOI22_X1 U23154 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19992), .B1(
        n20033), .B2(n19987), .ZN(n19985) );
  OAI211_X1 U23155 ( .C1(n20037), .C2(n20044), .A(n19986), .B(n19985), .ZN(
        P3_U2985) );
  AOI22_X1 U23156 ( .A1(n20039), .A2(n20050), .B1(n20038), .B2(n19991), .ZN(
        n19989) );
  AOI22_X1 U23157 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19992), .B1(
        n20041), .B2(n19987), .ZN(n19988) );
  OAI211_X1 U23158 ( .C1(n20045), .C2(n19990), .A(n19989), .B(n19988), .ZN(
        P3_U2986) );
  AOI22_X1 U23159 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19992), .B1(
        n20047), .B2(n19991), .ZN(n19995) );
  AOI22_X1 U23160 ( .A1(n20051), .A2(n19993), .B1(n20049), .B2(n20050), .ZN(
        n19994) );
  OAI211_X1 U23161 ( .C1(n20056), .C2(n19996), .A(n19995), .B(n19994), .ZN(
        P3_U2987) );
  AND2_X1 U23162 ( .A1(n20102), .A2(n20000), .ZN(n20046) );
  AOI22_X1 U23163 ( .A1(n19998), .A2(n20048), .B1(n19997), .B2(n20046), .ZN(
        n20005) );
  AOI22_X1 U23164 ( .A1(n20002), .A2(n20001), .B1(n20000), .B2(n19999), .ZN(
        n20052) );
  AOI22_X1 U23165 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20052), .B1(
        n20003), .B2(n20040), .ZN(n20004) );
  OAI211_X1 U23166 ( .C1(n20006), .C2(n20044), .A(n20005), .B(n20004), .ZN(
        P3_U2988) );
  AOI22_X1 U23167 ( .A1(n20008), .A2(n20046), .B1(n20007), .B2(n20050), .ZN(
        n20011) );
  AOI22_X1 U23168 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20052), .B1(
        n20009), .B2(n20040), .ZN(n20010) );
  OAI211_X1 U23169 ( .C1(n20012), .C2(n20036), .A(n20011), .B(n20010), .ZN(
        P3_U2989) );
  AOI22_X1 U23170 ( .A1(n20014), .A2(n20048), .B1(n20013), .B2(n20046), .ZN(
        n20017) );
  AOI22_X1 U23171 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20052), .B1(
        n20015), .B2(n20040), .ZN(n20016) );
  OAI211_X1 U23172 ( .C1(n20018), .C2(n20044), .A(n20017), .B(n20016), .ZN(
        P3_U2990) );
  AOI22_X1 U23173 ( .A1(n20020), .A2(n20048), .B1(n20019), .B2(n20046), .ZN(
        n20023) );
  AOI22_X1 U23174 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20052), .B1(
        n20021), .B2(n20040), .ZN(n20022) );
  OAI211_X1 U23175 ( .C1(n20024), .C2(n20044), .A(n20023), .B(n20022), .ZN(
        P3_U2991) );
  AOI22_X1 U23176 ( .A1(n20026), .A2(n20048), .B1(n20025), .B2(n20046), .ZN(
        n20029) );
  AOI22_X1 U23177 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20052), .B1(
        n20027), .B2(n20040), .ZN(n20028) );
  OAI211_X1 U23178 ( .C1(n20030), .C2(n20044), .A(n20029), .B(n20028), .ZN(
        P3_U2992) );
  AOI22_X1 U23179 ( .A1(n20032), .A2(n20050), .B1(n20031), .B2(n20046), .ZN(
        n20035) );
  AOI22_X1 U23180 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20052), .B1(
        n20033), .B2(n20040), .ZN(n20034) );
  OAI211_X1 U23181 ( .C1(n20037), .C2(n20036), .A(n20035), .B(n20034), .ZN(
        P3_U2993) );
  AOI22_X1 U23182 ( .A1(n20039), .A2(n20048), .B1(n20038), .B2(n20046), .ZN(
        n20043) );
  AOI22_X1 U23183 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20052), .B1(
        n20041), .B2(n20040), .ZN(n20042) );
  OAI211_X1 U23184 ( .C1(n20045), .C2(n20044), .A(n20043), .B(n20042), .ZN(
        P3_U2994) );
  AOI22_X1 U23185 ( .A1(n20049), .A2(n20048), .B1(n20047), .B2(n20046), .ZN(
        n20054) );
  AOI22_X1 U23186 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20052), .B1(
        n20051), .B2(n20050), .ZN(n20053) );
  OAI211_X1 U23187 ( .C1(n20056), .C2(n20055), .A(n20054), .B(n20053), .ZN(
        P3_U2995) );
  NOR2_X1 U23188 ( .A1(n20058), .A2(n20057), .ZN(n20060) );
  OAI222_X1 U23189 ( .A1(n20064), .A2(n20063), .B1(n20062), .B2(n20061), .C1(
        n20060), .C2(n20059), .ZN(n20210) );
  INV_X1 U23190 ( .A(n20065), .ZN(n20068) );
  OAI21_X1 U23191 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n20066), .ZN(n20067) );
  OAI211_X1 U23192 ( .C1(n20073), .C2(n20069), .A(n20068), .B(n20067), .ZN(
        n20093) );
  OR2_X1 U23193 ( .A1(n20070), .A2(n20082), .ZN(n20072) );
  AOI22_X1 U23194 ( .A1(n20072), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n20073), .B2(n20071), .ZN(n20091) );
  MUX2_X1 U23195 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n20074), .S(
        n20073), .Z(n20086) );
  INV_X1 U23196 ( .A(n20076), .ZN(n20079) );
  NAND2_X1 U23197 ( .A1(n20076), .A2(n20075), .ZN(n20078) );
  AOI22_X1 U23198 ( .A1(n12088), .A2(n20079), .B1(n20078), .B2(n20077), .ZN(
        n20083) );
  NAND2_X1 U23199 ( .A1(n20086), .A2(n20085), .ZN(n20080) );
  OAI211_X1 U23200 ( .C1(n20083), .C2(n20082), .A(n20081), .B(n20080), .ZN(
        n20084) );
  OAI211_X1 U23201 ( .C1(n20085), .C2(n20086), .A(n20084), .B(n20088), .ZN(
        n20090) );
  AOI21_X1 U23202 ( .B1(n20088), .B2(n20087), .A(n20086), .ZN(n20089) );
  AOI222_X1 U23203 ( .A1(n20091), .A2(n20090), .B1(n20091), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n20090), .C2(n20089), .ZN(
        n20092) );
  NOR4_X1 U23204 ( .A1(n20094), .A2(n20210), .A3(n20093), .A4(n20092), .ZN(
        n20106) );
  AOI22_X1 U23205 ( .A1(n20095), .A2(n20220), .B1(n20121), .B2(n20214), .ZN(
        n20096) );
  INV_X1 U23206 ( .A(n20096), .ZN(n20101) );
  OAI211_X1 U23207 ( .C1(n20098), .C2(n20097), .A(n20212), .B(n20106), .ZN(
        n20199) );
  OAI21_X1 U23208 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n20218), .A(n20199), 
        .ZN(n20108) );
  NOR2_X1 U23209 ( .A1(n20099), .A2(n20108), .ZN(n20100) );
  MUX2_X1 U23210 ( .A(n20101), .B(n20100), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n20104) );
  OR2_X1 U23211 ( .A1(n20109), .A2(n20102), .ZN(n20103) );
  OAI211_X1 U23212 ( .C1(n20106), .C2(n20105), .A(n20104), .B(n20103), .ZN(
        P3_U2996) );
  NAND2_X1 U23213 ( .A1(n20121), .A2(n20214), .ZN(n20112) );
  NAND4_X1 U23214 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(n20121), .A4(n20107), .ZN(n20114) );
  OR3_X1 U23215 ( .A1(n20110), .A2(n20109), .A3(n20108), .ZN(n20111) );
  NAND4_X1 U23216 ( .A1(n20113), .A2(n20112), .A3(n20114), .A4(n20111), .ZN(
        P3_U2997) );
  AND4_X1 U23217 ( .A1(n20116), .A2(n20115), .A3(n20114), .A4(n20198), .ZN(
        P3_U2998) );
  AND2_X1 U23218 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n20117), .ZN(
        P3_U2999) );
  AND2_X1 U23219 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n20117), .ZN(
        P3_U3000) );
  AND2_X1 U23220 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n20117), .ZN(
        P3_U3001) );
  AND2_X1 U23221 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n20117), .ZN(
        P3_U3002) );
  AND2_X1 U23222 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n20117), .ZN(
        P3_U3003) );
  AND2_X1 U23223 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n20117), .ZN(
        P3_U3004) );
  INV_X1 U23224 ( .A(P3_DATAWIDTH_REG_25__SCAN_IN), .ZN(n22047) );
  NOR2_X1 U23225 ( .A1(n22047), .A2(n20197), .ZN(P3_U3005) );
  AND2_X1 U23226 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n20117), .ZN(
        P3_U3006) );
  AND2_X1 U23227 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n20117), .ZN(
        P3_U3007) );
  AND2_X1 U23228 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n20117), .ZN(
        P3_U3008) );
  AND2_X1 U23229 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n20117), .ZN(
        P3_U3009) );
  AND2_X1 U23230 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n20117), .ZN(
        P3_U3010) );
  AND2_X1 U23231 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n20117), .ZN(
        P3_U3011) );
  AND2_X1 U23232 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n20117), .ZN(
        P3_U3012) );
  AND2_X1 U23233 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n20117), .ZN(
        P3_U3013) );
  INV_X1 U23234 ( .A(P3_DATAWIDTH_REG_16__SCAN_IN), .ZN(n22093) );
  NOR2_X1 U23235 ( .A1(n22093), .A2(n20197), .ZN(P3_U3014) );
  AND2_X1 U23236 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n20117), .ZN(
        P3_U3015) );
  AND2_X1 U23237 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n20117), .ZN(
        P3_U3016) );
  AND2_X1 U23238 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n20117), .ZN(
        P3_U3017) );
  INV_X1 U23239 ( .A(P3_DATAWIDTH_REG_12__SCAN_IN), .ZN(n21864) );
  NOR2_X1 U23240 ( .A1(n21864), .A2(n20197), .ZN(P3_U3018) );
  AND2_X1 U23241 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n20117), .ZN(
        P3_U3019) );
  INV_X1 U23242 ( .A(P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n21871) );
  NOR2_X1 U23243 ( .A1(n21871), .A2(n20197), .ZN(P3_U3020) );
  AND2_X1 U23244 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n20117), .ZN(P3_U3021) );
  AND2_X1 U23245 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n20117), .ZN(P3_U3022) );
  AND2_X1 U23246 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n20117), .ZN(P3_U3023) );
  AND2_X1 U23247 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n20117), .ZN(P3_U3024) );
  INV_X1 U23248 ( .A(P3_DATAWIDTH_REG_5__SCAN_IN), .ZN(n22085) );
  NOR2_X1 U23249 ( .A1(n22085), .A2(n20197), .ZN(P3_U3025) );
  AND2_X1 U23250 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n20117), .ZN(P3_U3026) );
  AND2_X1 U23251 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n20117), .ZN(P3_U3027) );
  AND2_X1 U23252 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n20117), .ZN(P3_U3028) );
  OAI21_X1 U23253 ( .B1(n20118), .B2(n21742), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n20119) );
  AOI22_X1 U23254 ( .A1(n20131), .A2(n20133), .B1(n20225), .B2(n20119), .ZN(
        n20120) );
  NAND3_X1 U23255 ( .A1(NA), .A2(n20131), .A3(n22024), .ZN(n20126) );
  OAI211_X1 U23256 ( .C1(n20218), .C2(n20124), .A(n20120), .B(n20126), .ZN(
        P3_U3029) );
  NOR2_X1 U23257 ( .A1(n20133), .A2(n21742), .ZN(n20129) );
  NOR2_X1 U23258 ( .A1(n20131), .A2(n20129), .ZN(n20122) );
  NAND2_X1 U23259 ( .A1(n20121), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n20127) );
  INV_X1 U23260 ( .A(n20127), .ZN(n20125) );
  AOI21_X1 U23261 ( .B1(n20122), .B2(P3_REQUESTPENDING_REG_SCAN_IN), .A(n20125), .ZN(n20123) );
  OAI211_X1 U23262 ( .C1(n21742), .C2(n20124), .A(n20123), .B(n20215), .ZN(
        P3_U3030) );
  AOI21_X1 U23263 ( .B1(n20131), .B2(n20126), .A(n20125), .ZN(n20132) );
  OAI22_X1 U23264 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n20127), .ZN(n20128) );
  OAI22_X1 U23265 ( .A1(n20129), .A2(n20128), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n20130) );
  OAI22_X1 U23266 ( .A1(n20132), .A2(n20133), .B1(n20131), .B2(n20130), .ZN(
        P3_U3031) );
  INV_X1 U23267 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n20135) );
  OAI222_X1 U23268 ( .A1(n20200), .A2(n20189), .B1(n20134), .B2(n20187), .C1(
        n20135), .C2(n20185), .ZN(P3_U3032) );
  OAI222_X1 U23269 ( .A1(n20185), .A2(n20137), .B1(n20136), .B2(n20187), .C1(
        n20135), .C2(n20189), .ZN(P3_U3033) );
  OAI222_X1 U23270 ( .A1(n20185), .A2(n20139), .B1(n20138), .B2(n20187), .C1(
        n20137), .C2(n20189), .ZN(P3_U3034) );
  OAI222_X1 U23271 ( .A1(n20185), .A2(n20141), .B1(n21908), .B2(n20187), .C1(
        n20139), .C2(n20189), .ZN(P3_U3035) );
  OAI222_X1 U23272 ( .A1(n20141), .A2(n20189), .B1(n20140), .B2(n20187), .C1(
        n20142), .C2(n20185), .ZN(P3_U3036) );
  OAI222_X1 U23273 ( .A1(n20185), .A2(n20144), .B1(n20143), .B2(n20187), .C1(
        n20142), .C2(n20189), .ZN(P3_U3037) );
  INV_X1 U23274 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n20147) );
  OAI222_X1 U23275 ( .A1(n20185), .A2(n20147), .B1(n20145), .B2(n20208), .C1(
        n20144), .C2(n20189), .ZN(P3_U3038) );
  OAI222_X1 U23276 ( .A1(n20147), .A2(n20189), .B1(n20146), .B2(n20187), .C1(
        n14407), .C2(n20185), .ZN(P3_U3039) );
  OAI222_X1 U23277 ( .A1(n20185), .A2(n20149), .B1(n20148), .B2(n20208), .C1(
        n14407), .C2(n20189), .ZN(P3_U3040) );
  OAI222_X1 U23278 ( .A1(n20185), .A2(n20151), .B1(n20150), .B2(n20208), .C1(
        n20149), .C2(n20189), .ZN(P3_U3041) );
  INV_X1 U23279 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n20153) );
  OAI222_X1 U23280 ( .A1(n20185), .A2(n20153), .B1(n20152), .B2(n20208), .C1(
        n20151), .C2(n20189), .ZN(P3_U3042) );
  OAI222_X1 U23281 ( .A1(n20185), .A2(n20155), .B1(n20154), .B2(n20208), .C1(
        n20153), .C2(n20189), .ZN(P3_U3043) );
  OAI222_X1 U23282 ( .A1(n20185), .A2(n20157), .B1(n20156), .B2(n20208), .C1(
        n20155), .C2(n20189), .ZN(P3_U3044) );
  OAI222_X1 U23283 ( .A1(n20185), .A2(n20159), .B1(n20158), .B2(n20208), .C1(
        n20157), .C2(n20189), .ZN(P3_U3045) );
  INV_X1 U23284 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n20160) );
  OAI222_X1 U23285 ( .A1(n20185), .A2(n20160), .B1(n21876), .B2(n20208), .C1(
        n20159), .C2(n20189), .ZN(P3_U3046) );
  OAI222_X1 U23286 ( .A1(n20185), .A2(n20162), .B1(n22060), .B2(n20208), .C1(
        n20160), .C2(n20189), .ZN(P3_U3047) );
  OAI222_X1 U23287 ( .A1(n20162), .A2(n20189), .B1(n20161), .B2(n20208), .C1(
        n20163), .C2(n20185), .ZN(P3_U3048) );
  INV_X1 U23288 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n20165) );
  OAI222_X1 U23289 ( .A1(n20185), .A2(n20165), .B1(n20164), .B2(n20208), .C1(
        n20163), .C2(n20189), .ZN(P3_U3049) );
  OAI222_X1 U23290 ( .A1(n20185), .A2(n20168), .B1(n20166), .B2(n20208), .C1(
        n20165), .C2(n20189), .ZN(P3_U3050) );
  OAI222_X1 U23291 ( .A1(n20168), .A2(n20189), .B1(n20167), .B2(n20208), .C1(
        n20169), .C2(n20185), .ZN(P3_U3051) );
  OAI222_X1 U23292 ( .A1(n20185), .A2(n20171), .B1(n20170), .B2(n20208), .C1(
        n20169), .C2(n20189), .ZN(P3_U3052) );
  OAI222_X1 U23293 ( .A1(n20185), .A2(n20173), .B1(n20172), .B2(n20208), .C1(
        n20171), .C2(n20189), .ZN(P3_U3053) );
  OAI222_X1 U23294 ( .A1(n20185), .A2(n22017), .B1(n20174), .B2(n20187), .C1(
        n20173), .C2(n20189), .ZN(P3_U3054) );
  OAI222_X1 U23295 ( .A1(n20185), .A2(n20176), .B1(n20175), .B2(n20187), .C1(
        n22017), .C2(n20189), .ZN(P3_U3055) );
  INV_X1 U23296 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n20178) );
  OAI222_X1 U23297 ( .A1(n20185), .A2(n20178), .B1(n22040), .B2(n20187), .C1(
        n20176), .C2(n20189), .ZN(P3_U3056) );
  OAI222_X1 U23298 ( .A1(n20178), .A2(n20189), .B1(n20177), .B2(n20187), .C1(
        n20179), .C2(n20185), .ZN(P3_U3057) );
  INV_X1 U23299 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n20182) );
  OAI222_X1 U23300 ( .A1(n20185), .A2(n20182), .B1(n20180), .B2(n20187), .C1(
        n20179), .C2(n20189), .ZN(P3_U3058) );
  OAI222_X1 U23301 ( .A1(n20182), .A2(n20189), .B1(n20181), .B2(n20187), .C1(
        n20183), .C2(n20185), .ZN(P3_U3059) );
  OAI222_X1 U23302 ( .A1(n20185), .A2(n22051), .B1(n20184), .B2(n20187), .C1(
        n20183), .C2(n20189), .ZN(P3_U3060) );
  OAI222_X1 U23303 ( .A1(n20189), .A2(n22051), .B1(n20188), .B2(n20187), .C1(
        n20186), .C2(n20185), .ZN(P3_U3061) );
  OAI22_X1 U23304 ( .A1(n20225), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n20187), .ZN(n20190) );
  INV_X1 U23305 ( .A(n20190), .ZN(P3_U3274) );
  OAI22_X1 U23306 ( .A1(n20225), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n20187), .ZN(n20191) );
  INV_X1 U23307 ( .A(n20191), .ZN(P3_U3275) );
  OAI22_X1 U23308 ( .A1(n20225), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n20187), .ZN(n20192) );
  INV_X1 U23309 ( .A(n20192), .ZN(P3_U3276) );
  OAI22_X1 U23310 ( .A1(n20225), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n20187), .ZN(n20193) );
  INV_X1 U23311 ( .A(n20193), .ZN(P3_U3277) );
  OAI21_X1 U23312 ( .B1(n20197), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n20195), 
        .ZN(n20194) );
  INV_X1 U23313 ( .A(n20194), .ZN(P3_U3280) );
  OAI21_X1 U23314 ( .B1(n20197), .B2(n20196), .A(n20195), .ZN(P3_U3281) );
  OAI221_X1 U23315 ( .B1(n21986), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n21986), 
        .C2(n20199), .A(n20198), .ZN(P3_U3282) );
  AOI21_X1 U23316 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20201) );
  AOI22_X1 U23317 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n20201), .B2(n20200), .ZN(n20203) );
  INV_X1 U23318 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20202) );
  AOI22_X1 U23319 ( .A1(n20204), .A2(n20203), .B1(n20202), .B2(n20206), .ZN(
        P3_U3292) );
  INV_X1 U23320 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n22112) );
  NOR2_X1 U23321 ( .A1(n20206), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n20205) );
  AOI22_X1 U23322 ( .A1(n22112), .A2(n20206), .B1(n13938), .B2(n20205), .ZN(
        P3_U3293) );
  INV_X1 U23323 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n20207) );
  AOI22_X1 U23324 ( .A1(n20208), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n20207), 
        .B2(n20225), .ZN(P3_U3294) );
  MUX2_X1 U23325 ( .A(P3_MORE_REG_SCAN_IN), .B(n20210), .S(n20209), .Z(
        P3_U3295) );
  OAI21_X1 U23326 ( .B1(n20212), .B2(n20211), .A(n20229), .ZN(n20213) );
  AOI21_X1 U23327 ( .B1(n20214), .B2(n20218), .A(n20213), .ZN(n20224) );
  AOI21_X1 U23328 ( .B1(n20217), .B2(n20216), .A(n20215), .ZN(n20219) );
  OAI211_X1 U23329 ( .C1(n20226), .C2(n20219), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n20218), .ZN(n20221) );
  AOI21_X1 U23330 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n20221), .A(n20220), 
        .ZN(n20223) );
  NAND2_X1 U23331 ( .A1(n20224), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20222) );
  OAI21_X1 U23332 ( .B1(n20224), .B2(n20223), .A(n20222), .ZN(P3_U3296) );
  MUX2_X1 U23333 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .B(P3_M_IO_N_REG_SCAN_IN), 
        .S(n20225), .Z(P3_U3297) );
  INV_X1 U23334 ( .A(n20226), .ZN(n20228) );
  OAI21_X1 U23335 ( .B1(n20230), .B2(P3_READREQUEST_REG_SCAN_IN), .A(n20229), 
        .ZN(n20227) );
  OAI21_X1 U23336 ( .B1(n20229), .B2(n20228), .A(n20227), .ZN(P3_U3298) );
  NOR2_X1 U23337 ( .A1(n20230), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n20232)
         );
  OAI21_X1 U23338 ( .B1(n20233), .B2(n20232), .A(n20231), .ZN(P3_U3299) );
  INV_X1 U23339 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20977) );
  NAND2_X1 U23340 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20977), .ZN(n20969) );
  OR2_X1 U23341 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n20966) );
  OAI21_X1 U23342 ( .B1(n20965), .B2(n20969), .A(n20966), .ZN(n21040) );
  AOI21_X1 U23343 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n21040), .ZN(n20234) );
  INV_X1 U23344 ( .A(n20234), .ZN(P2_U2815) );
  AOI22_X1 U23345 ( .A1(P2_D_C_N_REG_SCAN_IN), .A2(n21095), .B1(n20236), .B2(
        n20965), .ZN(n20235) );
  OAI21_X1 U23346 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(n21095), .A(n20235), 
        .ZN(P2_U2817) );
  OAI21_X1 U23347 ( .B1(n20236), .B2(BS16), .A(n21040), .ZN(n21038) );
  OAI21_X1 U23348 ( .B1(n21040), .B2(n20712), .A(n21038), .ZN(P2_U2818) );
  AND2_X1 U23349 ( .A1(n20238), .A2(n20237), .ZN(n21092) );
  OAI21_X1 U23350 ( .B1(n21092), .B2(n12578), .A(n20239), .ZN(P2_U2819) );
  NOR4_X1 U23351 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n20249) );
  NOR4_X1 U23352 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_6__SCAN_IN), .A3(P2_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_8__SCAN_IN), .ZN(n20248) );
  AOI211_X1 U23353 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_3__SCAN_IN), .B(
        P2_DATAWIDTH_REG_4__SCAN_IN), .ZN(n20240) );
  INV_X1 U23354 ( .A(P2_DATAWIDTH_REG_9__SCAN_IN), .ZN(n21968) );
  INV_X1 U23355 ( .A(P2_DATAWIDTH_REG_25__SCAN_IN), .ZN(n22129) );
  NAND3_X1 U23356 ( .A1(n20240), .A2(n21968), .A3(n22129), .ZN(n20246) );
  NOR4_X1 U23357 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n20244) );
  NOR4_X1 U23358 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n20243) );
  NOR4_X1 U23359 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20242) );
  NOR4_X1 U23360 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20241) );
  NAND4_X1 U23361 ( .A1(n20244), .A2(n20243), .A3(n20242), .A4(n20241), .ZN(
        n20245) );
  NOR4_X1 U23362 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_2__SCAN_IN), .A3(n20246), .A4(n20245), .ZN(n20247) );
  NAND3_X1 U23363 ( .A1(n20249), .A2(n20248), .A3(n20247), .ZN(n20257) );
  NOR2_X1 U23364 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n20257), .ZN(n20252) );
  INV_X1 U23365 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20250) );
  AOI22_X1 U23366 ( .A1(n20252), .A2(n12235), .B1(n20257), .B2(n20250), .ZN(
        P2_U2820) );
  INV_X1 U23367 ( .A(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n21926) );
  INV_X1 U23368 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21039) );
  NAND3_X1 U23369 ( .A1(n12235), .A2(n21926), .A3(n21039), .ZN(n20256) );
  INV_X1 U23370 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20251) );
  AOI22_X1 U23371 ( .A1(n20252), .A2(n20256), .B1(n20257), .B2(n20251), .ZN(
        P2_U2821) );
  NAND2_X1 U23372 ( .A1(n20252), .A2(n21039), .ZN(n20255) );
  INV_X1 U23373 ( .A(n20257), .ZN(n20259) );
  OAI21_X1 U23374 ( .B1(n12235), .B2(n20979), .A(n20259), .ZN(n20253) );
  OAI21_X1 U23375 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n20259), .A(n20253), 
        .ZN(n20254) );
  OAI221_X1 U23376 ( .B1(n20255), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n20255), .C2(P2_REIP_REG_0__SCAN_IN), .A(n20254), .ZN(P2_U2822) );
  INV_X1 U23377 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20258) );
  OAI221_X1 U23378 ( .B1(n20259), .B2(n20258), .C1(n20257), .C2(n20256), .A(
        n20255), .ZN(P2_U2823) );
  OAI21_X1 U23379 ( .B1(n20292), .B2(n21010), .A(n20260), .ZN(n20261) );
  AOI21_X1 U23380 ( .B1(n20262), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n20261), .ZN(n20263) );
  OAI21_X1 U23381 ( .B1(n20264), .B2(n20336), .A(n20263), .ZN(n20265) );
  INV_X1 U23382 ( .A(n20265), .ZN(n20276) );
  NOR2_X1 U23383 ( .A1(n10160), .A2(n20266), .ZN(n20268) );
  MUX2_X1 U23384 ( .A(n10160), .B(n20268), .S(n20267), .Z(n20270) );
  NOR3_X1 U23385 ( .A1(n20270), .A2(n20269), .A3(n20351), .ZN(n20273) );
  NOR2_X1 U23386 ( .A1(n20271), .A2(n20341), .ZN(n20272) );
  AOI211_X1 U23387 ( .C1(n20274), .C2(n20329), .A(n20273), .B(n20272), .ZN(
        n20275) );
  OAI211_X1 U23388 ( .C1(n21989), .C2(n20335), .A(n20276), .B(n20275), .ZN(
        P2_U2836) );
  OAI22_X1 U23389 ( .A1(n20278), .A2(n20336), .B1(n20277), .B2(n20339), .ZN(
        n20279) );
  AOI211_X1 U23390 ( .C1(P2_REIP_REG_15__SCAN_IN), .C2(n20344), .A(n20343), 
        .B(n20279), .ZN(n20291) );
  NAND2_X1 U23391 ( .A1(n20280), .A2(n20350), .ZN(n20282) );
  MUX2_X1 U23392 ( .A(n20350), .B(n20282), .S(n20281), .Z(n20284) );
  NAND3_X1 U23393 ( .A1(n20284), .A2(n20326), .A3(n20283), .ZN(n20287) );
  NAND2_X1 U23394 ( .A1(n20285), .A2(n20330), .ZN(n20286) );
  OAI211_X1 U23395 ( .C1(n20288), .C2(n20345), .A(n20287), .B(n20286), .ZN(
        n20289) );
  INV_X1 U23396 ( .A(n20289), .ZN(n20290) );
  OAI211_X1 U23397 ( .C1(n22063), .C2(n20335), .A(n20291), .B(n20290), .ZN(
        P2_U2840) );
  OAI22_X1 U23398 ( .A1(n20293), .A2(n20336), .B1(n21000), .B2(n20292), .ZN(
        n20294) );
  AOI211_X1 U23399 ( .C1(P2_EBX_REG_13__SCAN_IN), .C2(n20295), .A(n20343), .B(
        n20294), .ZN(n20306) );
  NOR2_X1 U23400 ( .A1(n10160), .A2(n20296), .ZN(n20298) );
  MUX2_X1 U23401 ( .A(n20298), .B(n10160), .S(n20297), .Z(n20300) );
  NOR3_X1 U23402 ( .A1(n20300), .A2(n20299), .A3(n20351), .ZN(n20303) );
  NOR2_X1 U23403 ( .A1(n20301), .A2(n20345), .ZN(n20302) );
  AOI211_X1 U23404 ( .C1(n20330), .C2(n20304), .A(n20303), .B(n20302), .ZN(
        n20305) );
  OAI211_X1 U23405 ( .C1(n10500), .C2(n20339), .A(n20306), .B(n20305), .ZN(
        P2_U2842) );
  OAI22_X1 U23406 ( .A1(n20308), .A2(n20336), .B1(n20307), .B2(n20339), .ZN(
        n20309) );
  AOI211_X1 U23407 ( .C1(P2_REIP_REG_9__SCAN_IN), .C2(n20344), .A(n20343), .B(
        n20309), .ZN(n20321) );
  NOR2_X1 U23408 ( .A1(n10160), .A2(n20310), .ZN(n20312) );
  MUX2_X1 U23409 ( .A(n10160), .B(n20312), .S(n20311), .Z(n20315) );
  INV_X1 U23410 ( .A(n20313), .ZN(n20314) );
  NOR3_X1 U23411 ( .A1(n20315), .A2(n20314), .A3(n20351), .ZN(n20318) );
  NOR2_X1 U23412 ( .A1(n20316), .A2(n20345), .ZN(n20317) );
  AOI211_X1 U23413 ( .C1(n20330), .C2(n20319), .A(n20318), .B(n20317), .ZN(
        n20320) );
  OAI211_X1 U23414 ( .C1(n10510), .C2(n20335), .A(n20321), .B(n20320), .ZN(
        P2_U2846) );
  OAI22_X1 U23415 ( .A1(n20322), .A2(n20336), .B1(n20335), .B2(n22065), .ZN(
        n20323) );
  AOI211_X1 U23416 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n20344), .A(n20343), .B(
        n20323), .ZN(n20333) );
  NOR2_X1 U23417 ( .A1(n10160), .A2(n9799), .ZN(n20325) );
  XNOR2_X1 U23418 ( .A(n20325), .B(n20324), .ZN(n20327) );
  AOI222_X1 U23419 ( .A1(n20331), .A2(n20330), .B1(n20329), .B2(n20328), .C1(
        n20327), .C2(n20326), .ZN(n20332) );
  OAI211_X1 U23420 ( .C1(n22021), .C2(n20339), .A(n20333), .B(n20332), .ZN(
        P2_U2850) );
  OAI22_X1 U23421 ( .A1(n20337), .A2(n20336), .B1(n20335), .B2(n20334), .ZN(
        n20338) );
  INV_X1 U23422 ( .A(n20338), .ZN(n20358) );
  OAI22_X1 U23423 ( .A1(n20369), .A2(n20341), .B1(n20340), .B2(n20339), .ZN(
        n20342) );
  AOI211_X1 U23424 ( .C1(P2_REIP_REG_4__SCAN_IN), .C2(n20344), .A(n20343), .B(
        n20342), .ZN(n20357) );
  NOR2_X1 U23425 ( .A1(n20346), .A2(n20345), .ZN(n20347) );
  AOI21_X1 U23426 ( .B1(n20372), .B2(n20348), .A(n20347), .ZN(n20356) );
  AND2_X1 U23427 ( .A1(n20350), .A2(n20349), .ZN(n20353) );
  AOI21_X1 U23428 ( .B1(n20353), .B2(n20354), .A(n20351), .ZN(n20352) );
  OAI21_X1 U23429 ( .B1(n20354), .B2(n20353), .A(n20352), .ZN(n20355) );
  NAND4_X1 U23430 ( .A1(n20358), .A2(n20357), .A3(n20356), .A4(n20355), .ZN(
        P2_U2851) );
  AOI22_X1 U23431 ( .A1(n20360), .A2(n20359), .B1(P2_EAX_REG_16__SCAN_IN), 
        .B2(n16938), .ZN(n20368) );
  AOI22_X1 U23432 ( .A1(n20362), .A2(BUF2_REG_16__SCAN_IN), .B1(n20361), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n20367) );
  INV_X1 U23433 ( .A(n20363), .ZN(n20365) );
  AOI22_X1 U23434 ( .A1(n20365), .A2(n20373), .B1(n20364), .B2(n20385), .ZN(
        n20366) );
  NAND3_X1 U23435 ( .A1(n20368), .A2(n20367), .A3(n20366), .ZN(P2_U2903) );
  INV_X1 U23436 ( .A(n20369), .ZN(n20370) );
  AOI22_X1 U23437 ( .A1(n20385), .A2(n20370), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n16938), .ZN(n20376) );
  XOR2_X1 U23438 ( .A(n20372), .B(n20371), .Z(n20374) );
  NAND2_X1 U23439 ( .A1(n20374), .A2(n20373), .ZN(n20375) );
  OAI211_X1 U23440 ( .C1(n20377), .C2(n20393), .A(n20376), .B(n20375), .ZN(
        P2_U2915) );
  AOI22_X1 U23441 ( .A1(n20385), .A2(n20378), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n16938), .ZN(n20384) );
  AOI21_X1 U23442 ( .B1(n20381), .B2(n20380), .A(n20379), .ZN(n20382) );
  OR2_X1 U23443 ( .A1(n20382), .A2(n20389), .ZN(n20383) );
  OAI211_X1 U23444 ( .C1(n20437), .C2(n20393), .A(n20384), .B(n20383), .ZN(
        P2_U2916) );
  AOI22_X1 U23445 ( .A1(n20385), .A2(n21067), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n16938), .ZN(n20392) );
  AOI21_X1 U23446 ( .B1(n20388), .B2(n20387), .A(n20386), .ZN(n20390) );
  OR2_X1 U23447 ( .A1(n20390), .A2(n20389), .ZN(n20391) );
  OAI211_X1 U23448 ( .C1(n20394), .C2(n20393), .A(n20392), .B(n20391), .ZN(
        P2_U2918) );
  AND2_X1 U23449 ( .A1(n20425), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  INV_X1 U23450 ( .A(P2_UWORD_REG_10__SCAN_IN), .ZN(n22004) );
  AOI22_X1 U23451 ( .A1(n20425), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(n20395), 
        .B2(P2_EAX_REG_26__SCAN_IN), .ZN(n20396) );
  OAI21_X1 U23452 ( .B1(n22004), .B2(n20419), .A(n20396), .ZN(P2_U2925) );
  AOI22_X1 U23453 ( .A1(n20426), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n20425), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n20397) );
  OAI21_X1 U23454 ( .B1(n20398), .B2(n20428), .A(n20397), .ZN(P2_U2936) );
  AOI22_X1 U23455 ( .A1(n20426), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n20425), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n20399) );
  OAI21_X1 U23456 ( .B1(n20400), .B2(n20428), .A(n20399), .ZN(P2_U2937) );
  AOI22_X1 U23457 ( .A1(n20426), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n20425), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n20401) );
  OAI21_X1 U23458 ( .B1(n20402), .B2(n20428), .A(n20401), .ZN(P2_U2938) );
  AOI22_X1 U23459 ( .A1(n20426), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n20425), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n20403) );
  OAI21_X1 U23460 ( .B1(n20404), .B2(n20428), .A(n20403), .ZN(P2_U2939) );
  AOI22_X1 U23461 ( .A1(n20426), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n20425), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n20405) );
  OAI21_X1 U23462 ( .B1(n21936), .B2(n20428), .A(n20405), .ZN(P2_U2940) );
  AOI22_X1 U23463 ( .A1(n20426), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n20425), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n20406) );
  OAI21_X1 U23464 ( .B1(n20407), .B2(n20428), .A(n20406), .ZN(P2_U2941) );
  AOI22_X1 U23465 ( .A1(n20426), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n20425), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n20408) );
  OAI21_X1 U23466 ( .B1(n20409), .B2(n20428), .A(n20408), .ZN(P2_U2942) );
  AOI22_X1 U23467 ( .A1(n20426), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n20425), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n20410) );
  OAI21_X1 U23468 ( .B1(n20411), .B2(n20428), .A(n20410), .ZN(P2_U2943) );
  AOI22_X1 U23469 ( .A1(n20426), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n20425), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n20412) );
  OAI21_X1 U23470 ( .B1(n20413), .B2(n20428), .A(n20412), .ZN(P2_U2944) );
  AOI22_X1 U23471 ( .A1(n20426), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n20425), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n20414) );
  OAI21_X1 U23472 ( .B1(n20415), .B2(n20428), .A(n20414), .ZN(P2_U2945) );
  AOI22_X1 U23473 ( .A1(n20426), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n20425), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n20416) );
  OAI21_X1 U23474 ( .B1(n16964), .B2(n20428), .A(n20416), .ZN(P2_U2946) );
  INV_X1 U23475 ( .A(P2_LWORD_REG_4__SCAN_IN), .ZN(n21923) );
  AOI22_X1 U23476 ( .A1(P2_EAX_REG_4__SCAN_IN), .A2(n20417), .B1(n20425), .B2(
        P2_DATAO_REG_4__SCAN_IN), .ZN(n20418) );
  OAI21_X1 U23477 ( .B1(n21923), .B2(n20419), .A(n20418), .ZN(P2_U2947) );
  INV_X1 U23478 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n20421) );
  AOI22_X1 U23479 ( .A1(n20426), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n20425), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n20420) );
  OAI21_X1 U23480 ( .B1(n20421), .B2(n20428), .A(n20420), .ZN(P2_U2948) );
  AOI22_X1 U23481 ( .A1(n20426), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n20425), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n20422) );
  OAI21_X1 U23482 ( .B1(n20423), .B2(n20428), .A(n20422), .ZN(P2_U2949) );
  INV_X1 U23483 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n22005) );
  AOI22_X1 U23484 ( .A1(n20426), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n20425), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n20424) );
  OAI21_X1 U23485 ( .B1(n22005), .B2(n20428), .A(n20424), .ZN(P2_U2950) );
  AOI22_X1 U23486 ( .A1(n20426), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n20425), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n20427) );
  OAI21_X1 U23487 ( .B1(n12894), .B2(n20428), .A(n20427), .ZN(P2_U2951) );
  AOI21_X1 U23488 ( .B1(n20430), .B2(P2_EAX_REG_26__SCAN_IN), .A(n20429), .ZN(
        n20431) );
  OAI21_X1 U23489 ( .B1(n22004), .B2(n20432), .A(n20431), .ZN(P2_U2962) );
  AOI22_X1 U23490 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20454), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n20453), .ZN(n20849) );
  INV_X1 U23491 ( .A(n20849), .ZN(n20920) );
  NOR2_X2 U23492 ( .A1(n20433), .A2(n20450), .ZN(n20918) );
  AOI22_X1 U23493 ( .A1(n20920), .A2(n20954), .B1(n20451), .B2(n20918), .ZN(
        n20436) );
  AND2_X1 U23494 ( .A1(n20896), .A2(n20434), .ZN(n20919) );
  AOI22_X1 U23495 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20454), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n20453), .ZN(n20474) );
  AOI22_X1 U23496 ( .A1(n20919), .A2(n20455), .B1(n9708), .B2(n20921), .ZN(
        n20435) );
  OAI211_X1 U23497 ( .C1(n20459), .C2(n12991), .A(n20436), .B(n20435), .ZN(
        P2_U3050) );
  AOI22_X1 U23498 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20454), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n20453), .ZN(n20852) );
  INV_X1 U23499 ( .A(n20852), .ZN(n20927) );
  NOR2_X2 U23500 ( .A1(n12211), .A2(n20450), .ZN(n20925) );
  AOI22_X1 U23501 ( .A1(n20927), .A2(n20954), .B1(n20451), .B2(n20925), .ZN(
        n20439) );
  NOR2_X2 U23502 ( .A1(n20437), .A2(n20623), .ZN(n20926) );
  AOI22_X1 U23503 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20454), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n20453), .ZN(n20595) );
  AOI22_X1 U23504 ( .A1(n20926), .A2(n20455), .B1(n9708), .B2(n20928), .ZN(
        n20438) );
  OAI211_X1 U23505 ( .C1(n20459), .C2(n12301), .A(n20439), .B(n20438), .ZN(
        P2_U3051) );
  INV_X1 U23506 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n20442) );
  AOI22_X1 U23507 ( .A1(n20934), .A2(n20954), .B1(n20932), .B2(n20451), .ZN(
        n20441) );
  AOI22_X1 U23508 ( .A1(n20933), .A2(n20455), .B1(n9708), .B2(n20935), .ZN(
        n20440) );
  OAI211_X1 U23509 ( .C1(n20459), .C2(n20442), .A(n20441), .B(n20440), .ZN(
        P2_U3052) );
  AOI22_X1 U23510 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n20453), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n20454), .ZN(n20858) );
  INV_X1 U23511 ( .A(n20858), .ZN(n20940) );
  NOR2_X2 U23512 ( .A1(n12631), .A2(n20450), .ZN(n20938) );
  AOI22_X1 U23513 ( .A1(n20940), .A2(n20954), .B1(n20451), .B2(n20938), .ZN(
        n20445) );
  NOR2_X2 U23514 ( .A1(n20443), .A2(n20623), .ZN(n20939) );
  AOI22_X1 U23515 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n20454), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n20453), .ZN(n20602) );
  AOI22_X1 U23516 ( .A1(n20939), .A2(n20455), .B1(n9708), .B2(n20941), .ZN(
        n20444) );
  OAI211_X1 U23517 ( .C1(n20459), .C2(n14494), .A(n20445), .B(n20444), .ZN(
        P2_U3053) );
  AOI22_X1 U23518 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n20453), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n20454), .ZN(n20861) );
  INV_X1 U23519 ( .A(n20861), .ZN(n20946) );
  NOR2_X2 U23520 ( .A1(n9715), .A2(n20450), .ZN(n20944) );
  AOI22_X1 U23521 ( .A1(n20946), .A2(n20954), .B1(n20451), .B2(n20944), .ZN(
        n20448) );
  NOR2_X2 U23522 ( .A1(n20623), .A2(n20446), .ZN(n20945) );
  AOI22_X1 U23523 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20454), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n20453), .ZN(n20672) );
  AOI22_X1 U23524 ( .A1(n20945), .A2(n20455), .B1(n9708), .B2(n20947), .ZN(
        n20447) );
  OAI211_X1 U23525 ( .C1(n20459), .C2(n20449), .A(n20448), .B(n20447), .ZN(
        P2_U3054) );
  AOI22_X1 U23526 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n20454), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n20453), .ZN(n20868) );
  INV_X1 U23527 ( .A(n20868), .ZN(n21834) );
  NOR2_X2 U23528 ( .A1(n10206), .A2(n20450), .ZN(n21831) );
  AOI22_X1 U23529 ( .A1(n21834), .A2(n20954), .B1(n20451), .B2(n21831), .ZN(
        n20457) );
  NOR2_X2 U23530 ( .A1(n20623), .A2(n20452), .ZN(n20951) );
  AOI22_X1 U23531 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20454), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n20453), .ZN(n20611) );
  AOI22_X1 U23532 ( .A1(n20951), .A2(n20455), .B1(n9708), .B2(n21835), .ZN(
        n20456) );
  OAI211_X1 U23533 ( .C1(n20459), .C2(n20458), .A(n20457), .B(n20456), .ZN(
        P2_U3055) );
  NOR2_X1 U23534 ( .A1(n20520), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20466) );
  INV_X1 U23535 ( .A(n20466), .ZN(n20462) );
  INV_X1 U23536 ( .A(n20460), .ZN(n20461) );
  NAND2_X1 U23537 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20466), .ZN(
        n20464) );
  INV_X1 U23538 ( .A(n20464), .ZN(n20484) );
  NOR3_X1 U23539 ( .A1(n20461), .A2(n20484), .A3(n20900), .ZN(n20463) );
  AOI211_X2 U23540 ( .C1(n20462), .C2(n20900), .A(n20647), .B(n20463), .ZN(
        n20485) );
  AOI22_X1 U23541 ( .A1(n20485), .A2(n20905), .B1(n20904), .B2(n20484), .ZN(
        n20468) );
  AOI211_X1 U23542 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n20464), .A(n20623), 
        .B(n20463), .ZN(n20465) );
  OAI221_X1 U23543 ( .B1(n20466), .B2(n20714), .C1(n20466), .C2(n20651), .A(
        n20465), .ZN(n20487) );
  AOI22_X1 U23544 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20487), .B1(
        n9708), .B2(n20906), .ZN(n20467) );
  OAI211_X1 U23545 ( .C1(n20587), .C2(n20518), .A(n20468), .B(n20467), .ZN(
        P2_U3056) );
  AOI22_X1 U23546 ( .A1(n20485), .A2(n20912), .B1(n20911), .B2(n20484), .ZN(
        n20471) );
  AOI22_X1 U23547 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20487), .B1(
        n9708), .B2(n20913), .ZN(n20470) );
  OAI211_X1 U23548 ( .C1(n20590), .C2(n20518), .A(n20471), .B(n20470), .ZN(
        P2_U3057) );
  AOI22_X1 U23549 ( .A1(n20485), .A2(n20919), .B1(n20918), .B2(n20484), .ZN(
        n20473) );
  AOI22_X1 U23550 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20487), .B1(
        n9708), .B2(n20920), .ZN(n20472) );
  OAI211_X1 U23551 ( .C1(n20474), .C2(n20518), .A(n20473), .B(n20472), .ZN(
        P2_U3058) );
  AOI22_X1 U23552 ( .A1(n20485), .A2(n20926), .B1(n20925), .B2(n20484), .ZN(
        n20476) );
  AOI22_X1 U23553 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20487), .B1(
        n9708), .B2(n20927), .ZN(n20475) );
  OAI211_X1 U23554 ( .C1(n20595), .C2(n20518), .A(n20476), .B(n20475), .ZN(
        P2_U3059) );
  AOI22_X1 U23555 ( .A1(n20485), .A2(n20933), .B1(n20932), .B2(n20484), .ZN(
        n20478) );
  AOI22_X1 U23556 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20487), .B1(
        n9708), .B2(n20934), .ZN(n20477) );
  OAI211_X1 U23557 ( .C1(n20479), .C2(n20518), .A(n20478), .B(n20477), .ZN(
        P2_U3060) );
  AOI22_X1 U23558 ( .A1(n20485), .A2(n20939), .B1(n20938), .B2(n20484), .ZN(
        n20481) );
  AOI22_X1 U23559 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20487), .B1(
        n9708), .B2(n20940), .ZN(n20480) );
  OAI211_X1 U23560 ( .C1(n20602), .C2(n20518), .A(n20481), .B(n20480), .ZN(
        P2_U3061) );
  AOI22_X1 U23561 ( .A1(n20485), .A2(n20945), .B1(n20944), .B2(n20484), .ZN(
        n20483) );
  AOI22_X1 U23562 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20487), .B1(
        n9708), .B2(n20946), .ZN(n20482) );
  OAI211_X1 U23563 ( .C1(n20672), .C2(n20518), .A(n20483), .B(n20482), .ZN(
        P2_U3062) );
  AOI22_X1 U23564 ( .A1(n20485), .A2(n20951), .B1(n21831), .B2(n20484), .ZN(
        n20489) );
  AOI22_X1 U23565 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20487), .B1(
        n9708), .B2(n21834), .ZN(n20488) );
  OAI211_X1 U23566 ( .C1(n20611), .C2(n20518), .A(n20489), .B(n20488), .ZN(
        P2_U3063) );
  INV_X1 U23567 ( .A(n20494), .ZN(n20490) );
  NOR2_X1 U23568 ( .A1(n22046), .A2(n20520), .ZN(n20519) );
  AND2_X1 U23569 ( .A1(n21083), .A2(n20519), .ZN(n20513) );
  OAI21_X1 U23570 ( .B1(n20490), .B2(n20513), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20491) );
  OR2_X1 U23571 ( .A1(n20751), .A2(n20520), .ZN(n20492) );
  NAND2_X1 U23572 ( .A1(n20491), .A2(n20492), .ZN(n20514) );
  AOI22_X1 U23573 ( .A1(n20514), .A2(n20905), .B1(n20904), .B2(n20513), .ZN(
        n20500) );
  AOI21_X1 U23574 ( .B1(n20498), .B2(n20518), .A(n20712), .ZN(n20497) );
  NAND2_X1 U23575 ( .A1(n20492), .A2(n21042), .ZN(n20496) );
  INV_X1 U23576 ( .A(n20513), .ZN(n20493) );
  OAI211_X1 U23577 ( .C1(n20494), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20717), 
        .B(n20493), .ZN(n20495) );
  OAI211_X1 U23578 ( .C1(n20497), .C2(n20496), .A(n20896), .B(n20495), .ZN(
        n20515) );
  AOI22_X1 U23579 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20515), .B1(
        n21833), .B2(n20907), .ZN(n20499) );
  OAI211_X1 U23580 ( .C1(n20843), .C2(n20518), .A(n20500), .B(n20499), .ZN(
        P2_U3064) );
  AOI22_X1 U23581 ( .A1(n20514), .A2(n20912), .B1(n20911), .B2(n20513), .ZN(
        n20502) );
  AOI22_X1 U23582 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20515), .B1(
        n21833), .B2(n20914), .ZN(n20501) );
  OAI211_X1 U23583 ( .C1(n20846), .C2(n20518), .A(n20502), .B(n20501), .ZN(
        P2_U3065) );
  AOI22_X1 U23584 ( .A1(n20514), .A2(n20919), .B1(n20918), .B2(n20513), .ZN(
        n20504) );
  AOI22_X1 U23585 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20515), .B1(
        n21833), .B2(n20921), .ZN(n20503) );
  OAI211_X1 U23586 ( .C1(n20849), .C2(n20518), .A(n20504), .B(n20503), .ZN(
        P2_U3066) );
  AOI22_X1 U23587 ( .A1(n20514), .A2(n20926), .B1(n20925), .B2(n20513), .ZN(
        n20506) );
  AOI22_X1 U23588 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20515), .B1(
        n21833), .B2(n20928), .ZN(n20505) );
  OAI211_X1 U23589 ( .C1(n20852), .C2(n20518), .A(n20506), .B(n20505), .ZN(
        P2_U3067) );
  AOI22_X1 U23590 ( .A1(n20514), .A2(n20933), .B1(n20932), .B2(n20513), .ZN(
        n20508) );
  AOI22_X1 U23591 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20515), .B1(
        n21833), .B2(n20935), .ZN(n20507) );
  OAI211_X1 U23592 ( .C1(n20855), .C2(n20518), .A(n20508), .B(n20507), .ZN(
        P2_U3068) );
  AOI22_X1 U23593 ( .A1(n20514), .A2(n20939), .B1(n20938), .B2(n20513), .ZN(
        n20510) );
  AOI22_X1 U23594 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20515), .B1(
        n21833), .B2(n20941), .ZN(n20509) );
  OAI211_X1 U23595 ( .C1(n20858), .C2(n20518), .A(n20510), .B(n20509), .ZN(
        P2_U3069) );
  AOI22_X1 U23596 ( .A1(n20514), .A2(n20945), .B1(n20944), .B2(n20513), .ZN(
        n20512) );
  AOI22_X1 U23597 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20515), .B1(
        n21833), .B2(n20947), .ZN(n20511) );
  OAI211_X1 U23598 ( .C1(n20861), .C2(n20518), .A(n20512), .B(n20511), .ZN(
        P2_U3070) );
  AOI22_X1 U23599 ( .A1(n20514), .A2(n20951), .B1(n21831), .B2(n20513), .ZN(
        n20517) );
  AOI22_X1 U23600 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20515), .B1(
        n21833), .B2(n21835), .ZN(n20516) );
  OAI211_X1 U23601 ( .C1(n20868), .C2(n20518), .A(n20517), .B(n20516), .ZN(
        P2_U3071) );
  INV_X1 U23602 ( .A(n20519), .ZN(n20524) );
  NOR2_X1 U23603 ( .A1(n20717), .A2(n20524), .ZN(n20523) );
  NOR2_X1 U23604 ( .A1(n20521), .A2(n20520), .ZN(n21832) );
  INV_X1 U23605 ( .A(n21832), .ZN(n20525) );
  AOI21_X1 U23606 ( .B1(n20526), .B2(n20525), .A(n20900), .ZN(n20522) );
  AOI22_X1 U23607 ( .A1(n20907), .A2(n21836), .B1(n20904), .B2(n21832), .ZN(
        n20530) );
  INV_X1 U23608 ( .A(n20651), .ZN(n20576) );
  NOR2_X1 U23609 ( .A1(n20576), .A2(n20752), .ZN(n20528) );
  OAI211_X1 U23610 ( .C1(n20526), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20717), 
        .B(n20525), .ZN(n20527) );
  OAI211_X1 U23611 ( .C1(n20528), .C2(n20519), .A(n20896), .B(n20527), .ZN(
        n21837) );
  AOI22_X1 U23612 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n21837), .B1(
        n21833), .B2(n20906), .ZN(n20529) );
  OAI211_X1 U23613 ( .C1(n21841), .C2(n20725), .A(n20530), .B(n20529), .ZN(
        P2_U3072) );
  AOI22_X1 U23614 ( .A1(n20914), .A2(n21836), .B1(n21832), .B2(n20911), .ZN(
        n20532) );
  AOI22_X1 U23615 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n21837), .B1(
        n21833), .B2(n20913), .ZN(n20531) );
  OAI211_X1 U23616 ( .C1(n21841), .C2(n20728), .A(n20532), .B(n20531), .ZN(
        P2_U3073) );
  INV_X1 U23617 ( .A(n20919), .ZN(n20731) );
  AOI22_X1 U23618 ( .A1(n20921), .A2(n21836), .B1(n21832), .B2(n20918), .ZN(
        n20534) );
  AOI22_X1 U23619 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n21837), .B1(
        n21833), .B2(n20920), .ZN(n20533) );
  OAI211_X1 U23620 ( .C1(n21841), .C2(n20731), .A(n20534), .B(n20533), .ZN(
        P2_U3074) );
  INV_X1 U23621 ( .A(n20926), .ZN(n20734) );
  AOI22_X1 U23622 ( .A1(n20928), .A2(n21836), .B1(n21832), .B2(n20925), .ZN(
        n20536) );
  AOI22_X1 U23623 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n21837), .B1(
        n21833), .B2(n20927), .ZN(n20535) );
  OAI211_X1 U23624 ( .C1(n21841), .C2(n20734), .A(n20536), .B(n20535), .ZN(
        P2_U3075) );
  INV_X1 U23625 ( .A(n20933), .ZN(n20737) );
  AOI22_X1 U23626 ( .A1(n20934), .A2(n21833), .B1(n20932), .B2(n21832), .ZN(
        n20538) );
  AOI22_X1 U23627 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n21837), .B1(
        n21836), .B2(n20935), .ZN(n20537) );
  OAI211_X1 U23628 ( .C1(n21841), .C2(n20737), .A(n20538), .B(n20537), .ZN(
        P2_U3076) );
  INV_X1 U23629 ( .A(n20939), .ZN(n20740) );
  AOI22_X1 U23630 ( .A1(n20940), .A2(n21833), .B1(n21832), .B2(n20938), .ZN(
        n20540) );
  AOI22_X1 U23631 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n21837), .B1(
        n21836), .B2(n20941), .ZN(n20539) );
  OAI211_X1 U23632 ( .C1(n21841), .C2(n20740), .A(n20540), .B(n20539), .ZN(
        P2_U3077) );
  INV_X1 U23633 ( .A(n20945), .ZN(n20743) );
  AOI22_X1 U23634 ( .A1(n20946), .A2(n21833), .B1(n21832), .B2(n20944), .ZN(
        n20542) );
  AOI22_X1 U23635 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n21837), .B1(
        n21836), .B2(n20947), .ZN(n20541) );
  OAI211_X1 U23636 ( .C1(n21841), .C2(n20743), .A(n20542), .B(n20541), .ZN(
        P2_U3078) );
  INV_X1 U23637 ( .A(n20619), .ZN(n20543) );
  NOR2_X1 U23638 ( .A1(n20617), .A2(n20678), .ZN(n20570) );
  AOI22_X1 U23639 ( .A1(n20907), .A2(n20606), .B1(n20904), .B2(n20570), .ZN(
        n20557) );
  AOI21_X1 U23640 ( .B1(n20551), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20549) );
  AOI21_X1 U23641 ( .B1(n20575), .B2(n20599), .A(n20712), .ZN(n20544) );
  NOR2_X1 U23642 ( .A1(n20544), .A2(n20717), .ZN(n20550) );
  INV_X1 U23643 ( .A(n20545), .ZN(n20547) );
  NAND2_X1 U23644 ( .A1(n20547), .A2(n20546), .ZN(n20554) );
  NAND2_X1 U23645 ( .A1(n20550), .A2(n20554), .ZN(n20548) );
  OAI211_X1 U23646 ( .C1(n20570), .C2(n20549), .A(n20548), .B(n20896), .ZN(
        n20572) );
  INV_X1 U23647 ( .A(n20550), .ZN(n20555) );
  INV_X1 U23648 ( .A(n20551), .ZN(n20552) );
  OAI21_X1 U23649 ( .B1(n20552), .B2(n20570), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20553) );
  AOI22_X1 U23650 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20572), .B1(
        n20905), .B2(n20571), .ZN(n20556) );
  OAI211_X1 U23651 ( .C1(n20843), .C2(n20575), .A(n20557), .B(n20556), .ZN(
        P2_U3080) );
  AOI22_X1 U23652 ( .A1(n20914), .A2(n20606), .B1(n20570), .B2(n20911), .ZN(
        n20559) );
  AOI22_X1 U23653 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20572), .B1(
        n20912), .B2(n20571), .ZN(n20558) );
  OAI211_X1 U23654 ( .C1(n20846), .C2(n20575), .A(n20559), .B(n20558), .ZN(
        P2_U3081) );
  AOI22_X1 U23655 ( .A1(n20921), .A2(n20606), .B1(n20570), .B2(n20918), .ZN(
        n20561) );
  AOI22_X1 U23656 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20572), .B1(
        n20919), .B2(n20571), .ZN(n20560) );
  OAI211_X1 U23657 ( .C1(n20849), .C2(n20575), .A(n20561), .B(n20560), .ZN(
        P2_U3082) );
  AOI22_X1 U23658 ( .A1(n20927), .A2(n21836), .B1(n20570), .B2(n20925), .ZN(
        n20563) );
  AOI22_X1 U23659 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20572), .B1(
        n20926), .B2(n20571), .ZN(n20562) );
  OAI211_X1 U23660 ( .C1(n20595), .C2(n20599), .A(n20563), .B(n20562), .ZN(
        P2_U3083) );
  AOI22_X1 U23661 ( .A1(n20935), .A2(n20606), .B1(n20932), .B2(n20570), .ZN(
        n20565) );
  AOI22_X1 U23662 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20572), .B1(
        n20933), .B2(n20571), .ZN(n20564) );
  OAI211_X1 U23663 ( .C1(n20855), .C2(n20575), .A(n20565), .B(n20564), .ZN(
        P2_U3084) );
  AOI22_X1 U23664 ( .A1(n20941), .A2(n20606), .B1(n20570), .B2(n20938), .ZN(
        n20567) );
  AOI22_X1 U23665 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20572), .B1(
        n20939), .B2(n20571), .ZN(n20566) );
  OAI211_X1 U23666 ( .C1(n20858), .C2(n20575), .A(n20567), .B(n20566), .ZN(
        P2_U3085) );
  AOI22_X1 U23667 ( .A1(n20947), .A2(n20606), .B1(n20570), .B2(n20944), .ZN(
        n20569) );
  AOI22_X1 U23668 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20572), .B1(
        n20945), .B2(n20571), .ZN(n20568) );
  OAI211_X1 U23669 ( .C1(n20861), .C2(n20575), .A(n20569), .B(n20568), .ZN(
        P2_U3086) );
  AOI22_X1 U23670 ( .A1(n21835), .A2(n20606), .B1(n20570), .B2(n21831), .ZN(
        n20574) );
  AOI22_X1 U23671 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20572), .B1(
        n20951), .B2(n20571), .ZN(n20573) );
  OAI211_X1 U23672 ( .C1(n20868), .C2(n20575), .A(n20574), .B(n20573), .ZN(
        P2_U3087) );
  NOR2_X1 U23673 ( .A1(n20617), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20579) );
  INV_X1 U23674 ( .A(n20579), .ZN(n20583) );
  NOR2_X1 U23675 ( .A1(n21083), .A2(n20583), .ZN(n20605) );
  AOI22_X1 U23676 ( .A1(n20906), .A2(n20606), .B1(n20904), .B2(n20605), .ZN(
        n20586) );
  OAI21_X1 U23677 ( .B1(n20576), .B2(n21062), .A(n21042), .ZN(n20584) );
  INV_X1 U23678 ( .A(n20605), .ZN(n20577) );
  OAI211_X1 U23679 ( .C1(n20580), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20717), 
        .B(n20577), .ZN(n20578) );
  OAI211_X1 U23680 ( .C1(n20584), .C2(n20579), .A(n20896), .B(n20578), .ZN(
        n20608) );
  INV_X1 U23681 ( .A(n20580), .ZN(n20581) );
  OAI21_X1 U23682 ( .B1(n20581), .B2(n20605), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20582) );
  AOI22_X1 U23683 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20608), .B1(
        n20905), .B2(n20607), .ZN(n20585) );
  OAI211_X1 U23684 ( .C1(n20587), .C2(n20644), .A(n20586), .B(n20585), .ZN(
        P2_U3088) );
  AOI22_X1 U23685 ( .A1(n20913), .A2(n20606), .B1(n20605), .B2(n20911), .ZN(
        n20589) );
  AOI22_X1 U23686 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20608), .B1(
        n20912), .B2(n20607), .ZN(n20588) );
  OAI211_X1 U23687 ( .C1(n20590), .C2(n20644), .A(n20589), .B(n20588), .ZN(
        P2_U3089) );
  INV_X1 U23688 ( .A(n20644), .ZN(n20596) );
  AOI22_X1 U23689 ( .A1(n20921), .A2(n20596), .B1(n20605), .B2(n20918), .ZN(
        n20592) );
  AOI22_X1 U23690 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20608), .B1(
        n20919), .B2(n20607), .ZN(n20591) );
  OAI211_X1 U23691 ( .C1(n20849), .C2(n20599), .A(n20592), .B(n20591), .ZN(
        P2_U3090) );
  AOI22_X1 U23692 ( .A1(n20927), .A2(n20606), .B1(n20605), .B2(n20925), .ZN(
        n20594) );
  AOI22_X1 U23693 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20608), .B1(
        n20926), .B2(n20607), .ZN(n20593) );
  OAI211_X1 U23694 ( .C1(n20595), .C2(n20644), .A(n20594), .B(n20593), .ZN(
        P2_U3091) );
  AOI22_X1 U23695 ( .A1(n20935), .A2(n20596), .B1(n20932), .B2(n20605), .ZN(
        n20598) );
  AOI22_X1 U23696 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20608), .B1(
        n20933), .B2(n20607), .ZN(n20597) );
  OAI211_X1 U23697 ( .C1(n20855), .C2(n20599), .A(n20598), .B(n20597), .ZN(
        P2_U3092) );
  AOI22_X1 U23698 ( .A1(n20940), .A2(n20606), .B1(n20938), .B2(n20605), .ZN(
        n20601) );
  AOI22_X1 U23699 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20608), .B1(
        n20939), .B2(n20607), .ZN(n20600) );
  OAI211_X1 U23700 ( .C1(n20602), .C2(n20644), .A(n20601), .B(n20600), .ZN(
        P2_U3093) );
  AOI22_X1 U23701 ( .A1(n20946), .A2(n20606), .B1(n20944), .B2(n20605), .ZN(
        n20604) );
  AOI22_X1 U23702 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20608), .B1(
        n20945), .B2(n20607), .ZN(n20603) );
  OAI211_X1 U23703 ( .C1(n20672), .C2(n20644), .A(n20604), .B(n20603), .ZN(
        P2_U3094) );
  AOI22_X1 U23704 ( .A1(n21834), .A2(n20606), .B1(n21831), .B2(n20605), .ZN(
        n20610) );
  AOI22_X1 U23705 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20608), .B1(
        n20951), .B2(n20607), .ZN(n20609) );
  OAI211_X1 U23706 ( .C1(n20611), .C2(n20644), .A(n20610), .B(n20609), .ZN(
        P2_U3095) );
  NAND3_X1 U23707 ( .A1(n20613), .A2(n20834), .A3(n20612), .ZN(n20616) );
  INV_X1 U23708 ( .A(n20614), .ZN(n20615) );
  NOR3_X2 U23709 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n20892), .ZN(n20639) );
  NOR3_X1 U23710 ( .A1(n20615), .A2(n20639), .A3(n20900), .ZN(n20624) );
  AOI21_X1 U23711 ( .B1(n20900), .B2(n20616), .A(n20624), .ZN(n20640) );
  AOI22_X1 U23712 ( .A1(n20640), .A2(n20905), .B1(n20904), .B2(n20639), .ZN(
        n20626) );
  NOR2_X1 U23713 ( .A1(n20618), .A2(n20617), .ZN(n20621) );
  NOR2_X4 U23714 ( .A1(n20650), .A2(n20619), .ZN(n20669) );
  AOI21_X1 U23715 ( .B1(n20677), .B2(n20644), .A(n20712), .ZN(n20620) );
  OAI22_X1 U23716 ( .A1(n20621), .A2(n20620), .B1(n20639), .B2(n20834), .ZN(
        n20622) );
  AOI22_X1 U23717 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20641), .B1(
        n20669), .B2(n20907), .ZN(n20625) );
  OAI211_X1 U23718 ( .C1(n20843), .C2(n20644), .A(n20626), .B(n20625), .ZN(
        P2_U3096) );
  AOI22_X1 U23719 ( .A1(n20640), .A2(n20912), .B1(n20911), .B2(n20639), .ZN(
        n20628) );
  AOI22_X1 U23720 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20641), .B1(
        n20669), .B2(n20914), .ZN(n20627) );
  OAI211_X1 U23721 ( .C1(n20846), .C2(n20644), .A(n20628), .B(n20627), .ZN(
        P2_U3097) );
  AOI22_X1 U23722 ( .A1(n20640), .A2(n20919), .B1(n20918), .B2(n20639), .ZN(
        n20630) );
  AOI22_X1 U23723 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20641), .B1(
        n20669), .B2(n20921), .ZN(n20629) );
  OAI211_X1 U23724 ( .C1(n20849), .C2(n20644), .A(n20630), .B(n20629), .ZN(
        P2_U3098) );
  AOI22_X1 U23725 ( .A1(n20640), .A2(n20926), .B1(n20925), .B2(n20639), .ZN(
        n20632) );
  AOI22_X1 U23726 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20641), .B1(
        n20669), .B2(n20928), .ZN(n20631) );
  OAI211_X1 U23727 ( .C1(n20852), .C2(n20644), .A(n20632), .B(n20631), .ZN(
        P2_U3099) );
  AOI22_X1 U23728 ( .A1(n20640), .A2(n20933), .B1(n20932), .B2(n20639), .ZN(
        n20634) );
  AOI22_X1 U23729 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20641), .B1(
        n20669), .B2(n20935), .ZN(n20633) );
  OAI211_X1 U23730 ( .C1(n20855), .C2(n20644), .A(n20634), .B(n20633), .ZN(
        P2_U3100) );
  AOI22_X1 U23731 ( .A1(n20640), .A2(n20939), .B1(n20938), .B2(n20639), .ZN(
        n20636) );
  AOI22_X1 U23732 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20641), .B1(
        n20669), .B2(n20941), .ZN(n20635) );
  OAI211_X1 U23733 ( .C1(n20858), .C2(n20644), .A(n20636), .B(n20635), .ZN(
        P2_U3101) );
  AOI22_X1 U23734 ( .A1(n20640), .A2(n20945), .B1(n20944), .B2(n20639), .ZN(
        n20638) );
  AOI22_X1 U23735 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20641), .B1(
        n20669), .B2(n20947), .ZN(n20637) );
  OAI211_X1 U23736 ( .C1(n20861), .C2(n20644), .A(n20638), .B(n20637), .ZN(
        P2_U3102) );
  AOI22_X1 U23737 ( .A1(n20640), .A2(n20951), .B1(n21831), .B2(n20639), .ZN(
        n20643) );
  AOI22_X1 U23738 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20641), .B1(
        n20669), .B2(n21835), .ZN(n20642) );
  OAI211_X1 U23739 ( .C1(n20868), .C2(n20644), .A(n20643), .B(n20642), .ZN(
        P2_U3103) );
  NOR2_X1 U23740 ( .A1(n20892), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20655) );
  INV_X1 U23741 ( .A(n20655), .ZN(n20648) );
  AND2_X1 U23742 ( .A1(n20649), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20645) );
  AOI211_X2 U23743 ( .C1(n20648), .C2(n20900), .A(n20647), .B(n20653), .ZN(
        n20673) );
  INV_X1 U23744 ( .A(n20649), .ZN(n20684) );
  AOI22_X1 U23745 ( .A1(n20673), .A2(n20905), .B1(n20684), .B2(n20904), .ZN(
        n20658) );
  AND2_X1 U23746 ( .A1(n20651), .A2(n20893), .ZN(n21041) );
  OAI21_X1 U23747 ( .B1(n20684), .B2(n20834), .A(n20896), .ZN(n20652) );
  NOR2_X1 U23748 ( .A1(n20653), .A2(n20652), .ZN(n20654) );
  AOI22_X1 U23749 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20674), .B1(
        n20679), .B2(n20907), .ZN(n20657) );
  OAI211_X1 U23750 ( .C1(n20843), .C2(n20677), .A(n20658), .B(n20657), .ZN(
        P2_U3104) );
  AOI22_X1 U23751 ( .A1(n20673), .A2(n20912), .B1(n20684), .B2(n20911), .ZN(
        n20660) );
  AOI22_X1 U23752 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20674), .B1(
        n20679), .B2(n20914), .ZN(n20659) );
  OAI211_X1 U23753 ( .C1(n20846), .C2(n20677), .A(n20660), .B(n20659), .ZN(
        P2_U3105) );
  AOI22_X1 U23754 ( .A1(n20673), .A2(n20919), .B1(n20684), .B2(n20918), .ZN(
        n20662) );
  AOI22_X1 U23755 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20674), .B1(
        n20679), .B2(n20921), .ZN(n20661) );
  OAI211_X1 U23756 ( .C1(n20849), .C2(n20677), .A(n20662), .B(n20661), .ZN(
        P2_U3106) );
  AOI22_X1 U23757 ( .A1(n20673), .A2(n20926), .B1(n20684), .B2(n20925), .ZN(
        n20664) );
  AOI22_X1 U23758 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20674), .B1(
        n20679), .B2(n20928), .ZN(n20663) );
  OAI211_X1 U23759 ( .C1(n20852), .C2(n20677), .A(n20664), .B(n20663), .ZN(
        P2_U3107) );
  AOI22_X1 U23760 ( .A1(n20673), .A2(n20933), .B1(n20684), .B2(n20932), .ZN(
        n20666) );
  AOI22_X1 U23761 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20674), .B1(
        n20679), .B2(n20935), .ZN(n20665) );
  OAI211_X1 U23762 ( .C1(n20855), .C2(n20677), .A(n20666), .B(n20665), .ZN(
        P2_U3108) );
  AOI22_X1 U23763 ( .A1(n20673), .A2(n20939), .B1(n20684), .B2(n20938), .ZN(
        n20668) );
  AOI22_X1 U23764 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20674), .B1(
        n20679), .B2(n20941), .ZN(n20667) );
  OAI211_X1 U23765 ( .C1(n20858), .C2(n20677), .A(n20668), .B(n20667), .ZN(
        P2_U3109) );
  AOI22_X1 U23766 ( .A1(n20673), .A2(n20945), .B1(n20684), .B2(n20944), .ZN(
        n20671) );
  AOI22_X1 U23767 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20674), .B1(
        n20669), .B2(n20946), .ZN(n20670) );
  OAI211_X1 U23768 ( .C1(n20672), .C2(n20708), .A(n20671), .B(n20670), .ZN(
        P2_U3110) );
  AOI22_X1 U23769 ( .A1(n20673), .A2(n20951), .B1(n20684), .B2(n21831), .ZN(
        n20676) );
  AOI22_X1 U23770 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20674), .B1(
        n20679), .B2(n21835), .ZN(n20675) );
  OAI211_X1 U23771 ( .C1(n20868), .C2(n20677), .A(n20676), .B(n20675), .ZN(
        P2_U3111) );
  NOR2_X1 U23772 ( .A1(n21054), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20781) );
  INV_X1 U23773 ( .A(n20781), .ZN(n20783) );
  NOR2_X1 U23774 ( .A1(n20678), .A2(n20783), .ZN(n20703) );
  AOI22_X1 U23775 ( .A1(n20907), .A2(n20744), .B1(n20904), .B2(n20703), .ZN(
        n20690) );
  NOR2_X1 U23776 ( .A1(n20681), .A2(n20680), .ZN(n20688) );
  NOR2_X1 U23777 ( .A1(n20688), .A2(n20684), .ZN(n20682) );
  NOR2_X1 U23778 ( .A1(n20684), .A2(n20703), .ZN(n20687) );
  OAI21_X1 U23779 ( .B1(n20685), .B2(n20703), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20686) );
  AOI22_X1 U23780 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20705), .B1(
        n20905), .B2(n20704), .ZN(n20689) );
  OAI211_X1 U23781 ( .C1(n20843), .C2(n20708), .A(n20690), .B(n20689), .ZN(
        P2_U3112) );
  AOI22_X1 U23782 ( .A1(n20914), .A2(n20744), .B1(n20703), .B2(n20911), .ZN(
        n20692) );
  AOI22_X1 U23783 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20705), .B1(
        n20704), .B2(n20912), .ZN(n20691) );
  OAI211_X1 U23784 ( .C1(n20846), .C2(n20708), .A(n20692), .B(n20691), .ZN(
        P2_U3113) );
  AOI22_X1 U23785 ( .A1(n20921), .A2(n20744), .B1(n20918), .B2(n20703), .ZN(
        n20694) );
  AOI22_X1 U23786 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20705), .B1(
        n20704), .B2(n20919), .ZN(n20693) );
  OAI211_X1 U23787 ( .C1(n20849), .C2(n20708), .A(n20694), .B(n20693), .ZN(
        P2_U3114) );
  AOI22_X1 U23788 ( .A1(n20928), .A2(n20744), .B1(n20925), .B2(n20703), .ZN(
        n20696) );
  AOI22_X1 U23789 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20705), .B1(
        n20704), .B2(n20926), .ZN(n20695) );
  OAI211_X1 U23790 ( .C1(n20852), .C2(n20708), .A(n20696), .B(n20695), .ZN(
        P2_U3115) );
  AOI22_X1 U23791 ( .A1(n20935), .A2(n20744), .B1(n20932), .B2(n20703), .ZN(
        n20698) );
  AOI22_X1 U23792 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20705), .B1(
        n20704), .B2(n20933), .ZN(n20697) );
  OAI211_X1 U23793 ( .C1(n20855), .C2(n20708), .A(n20698), .B(n20697), .ZN(
        P2_U3116) );
  AOI22_X1 U23794 ( .A1(n20941), .A2(n20744), .B1(n20938), .B2(n20703), .ZN(
        n20700) );
  AOI22_X1 U23795 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20705), .B1(
        n20704), .B2(n20939), .ZN(n20699) );
  OAI211_X1 U23796 ( .C1(n20858), .C2(n20708), .A(n20700), .B(n20699), .ZN(
        P2_U3117) );
  AOI22_X1 U23797 ( .A1(n20947), .A2(n20744), .B1(n20944), .B2(n20703), .ZN(
        n20702) );
  AOI22_X1 U23798 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20705), .B1(
        n20704), .B2(n20945), .ZN(n20701) );
  OAI211_X1 U23799 ( .C1(n20861), .C2(n20708), .A(n20702), .B(n20701), .ZN(
        P2_U3118) );
  AOI22_X1 U23800 ( .A1(n21835), .A2(n20744), .B1(n21831), .B2(n20703), .ZN(
        n20707) );
  AOI22_X1 U23801 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20705), .B1(
        n20704), .B2(n20951), .ZN(n20706) );
  OAI211_X1 U23802 ( .C1(n20868), .C2(n20708), .A(n20707), .B(n20706), .ZN(
        P2_U3119) );
  NAND3_X1 U23803 ( .A1(n22046), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(
        n20781), .ZN(n20718) );
  NAND2_X1 U23804 ( .A1(n12429), .A2(n20718), .ZN(n20710) );
  NOR2_X1 U23805 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20783), .ZN(
        n20711) );
  AND2_X1 U23806 ( .A1(n20711), .A2(n21042), .ZN(n20709) );
  INV_X1 U23807 ( .A(n20718), .ZN(n20754) );
  AOI22_X1 U23808 ( .A1(n20906), .A2(n20744), .B1(n20904), .B2(n20754), .ZN(
        n20724) );
  INV_X1 U23809 ( .A(n20711), .ZN(n20716) );
  NAND2_X1 U23810 ( .A1(n20894), .A2(n20714), .ZN(n20715) );
  NAND2_X1 U23811 ( .A1(n20716), .A2(n20715), .ZN(n20720) );
  OAI211_X1 U23812 ( .C1(n12429), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20718), 
        .B(n20717), .ZN(n20719) );
  NAND3_X1 U23813 ( .A1(n20720), .A2(n20896), .A3(n20719), .ZN(n20745) );
  AOI22_X1 U23814 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20745), .B1(
        n20755), .B2(n20907), .ZN(n20723) );
  OAI211_X1 U23815 ( .C1(n20748), .C2(n20725), .A(n20724), .B(n20723), .ZN(
        P2_U3120) );
  AOI22_X1 U23816 ( .A1(n20913), .A2(n20744), .B1(n20754), .B2(n20911), .ZN(
        n20727) );
  AOI22_X1 U23817 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20745), .B1(
        n20755), .B2(n20914), .ZN(n20726) );
  OAI211_X1 U23818 ( .C1(n20748), .C2(n20728), .A(n20727), .B(n20726), .ZN(
        P2_U3121) );
  AOI22_X1 U23819 ( .A1(n20920), .A2(n20744), .B1(n20918), .B2(n20754), .ZN(
        n20730) );
  AOI22_X1 U23820 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20745), .B1(
        n20755), .B2(n20921), .ZN(n20729) );
  OAI211_X1 U23821 ( .C1(n20748), .C2(n20731), .A(n20730), .B(n20729), .ZN(
        P2_U3122) );
  AOI22_X1 U23822 ( .A1(n20927), .A2(n20744), .B1(n20925), .B2(n20754), .ZN(
        n20733) );
  AOI22_X1 U23823 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20745), .B1(
        n20755), .B2(n20928), .ZN(n20732) );
  OAI211_X1 U23824 ( .C1(n20748), .C2(n20734), .A(n20733), .B(n20732), .ZN(
        P2_U3123) );
  AOI22_X1 U23825 ( .A1(n20934), .A2(n20744), .B1(n20932), .B2(n20754), .ZN(
        n20736) );
  AOI22_X1 U23826 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20745), .B1(
        n20755), .B2(n20935), .ZN(n20735) );
  OAI211_X1 U23827 ( .C1(n20748), .C2(n20737), .A(n20736), .B(n20735), .ZN(
        P2_U3124) );
  AOI22_X1 U23828 ( .A1(n20941), .A2(n20755), .B1(n20754), .B2(n20938), .ZN(
        n20739) );
  AOI22_X1 U23829 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20745), .B1(
        n20744), .B2(n20940), .ZN(n20738) );
  OAI211_X1 U23830 ( .C1(n20748), .C2(n20740), .A(n20739), .B(n20738), .ZN(
        P2_U3125) );
  AOI22_X1 U23831 ( .A1(n20946), .A2(n20744), .B1(n20944), .B2(n20754), .ZN(
        n20742) );
  AOI22_X1 U23832 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20745), .B1(
        n20755), .B2(n20947), .ZN(n20741) );
  OAI211_X1 U23833 ( .C1(n20748), .C2(n20743), .A(n20742), .B(n20741), .ZN(
        P2_U3126) );
  INV_X1 U23834 ( .A(n20951), .ZN(n21840) );
  AOI22_X1 U23835 ( .A1(n21835), .A2(n20755), .B1(n20754), .B2(n21831), .ZN(
        n20747) );
  AOI22_X1 U23836 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20745), .B1(
        n20744), .B2(n21834), .ZN(n20746) );
  OAI211_X1 U23837 ( .C1(n20748), .C2(n21840), .A(n20747), .B(n20746), .ZN(
        P2_U3127) );
  INV_X1 U23838 ( .A(n20757), .ZN(n20749) );
  NOR3_X2 U23839 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22046), .A3(
        n20783), .ZN(n20773) );
  OAI21_X1 U23840 ( .B1(n20749), .B2(n20773), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20750) );
  AOI22_X1 U23841 ( .A1(n20774), .A2(n20905), .B1(n20904), .B2(n20773), .ZN(
        n20760) );
  AOI221_X1 U23842 ( .B1(n20779), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n20755), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n20754), .ZN(n20756) );
  AOI211_X1 U23843 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n20757), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n20756), .ZN(n20758) );
  OAI21_X1 U23844 ( .B1(n20758), .B2(n20773), .A(n20896), .ZN(n20775) );
  AOI22_X1 U23845 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20775), .B1(
        n20779), .B2(n20907), .ZN(n20759) );
  OAI211_X1 U23846 ( .C1(n20843), .C2(n20778), .A(n20760), .B(n20759), .ZN(
        P2_U3128) );
  AOI22_X1 U23847 ( .A1(n20774), .A2(n20912), .B1(n20911), .B2(n20773), .ZN(
        n20762) );
  AOI22_X1 U23848 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20775), .B1(
        n20779), .B2(n20914), .ZN(n20761) );
  OAI211_X1 U23849 ( .C1(n20846), .C2(n20778), .A(n20762), .B(n20761), .ZN(
        P2_U3129) );
  AOI22_X1 U23850 ( .A1(n20774), .A2(n20919), .B1(n20918), .B2(n20773), .ZN(
        n20764) );
  AOI22_X1 U23851 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20775), .B1(
        n20779), .B2(n20921), .ZN(n20763) );
  OAI211_X1 U23852 ( .C1(n20849), .C2(n20778), .A(n20764), .B(n20763), .ZN(
        P2_U3130) );
  AOI22_X1 U23853 ( .A1(n20774), .A2(n20926), .B1(n20925), .B2(n20773), .ZN(
        n20766) );
  AOI22_X1 U23854 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20775), .B1(
        n20779), .B2(n20928), .ZN(n20765) );
  OAI211_X1 U23855 ( .C1(n20852), .C2(n20778), .A(n20766), .B(n20765), .ZN(
        P2_U3131) );
  AOI22_X1 U23856 ( .A1(n20774), .A2(n20933), .B1(n20932), .B2(n20773), .ZN(
        n20768) );
  AOI22_X1 U23857 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20775), .B1(
        n20779), .B2(n20935), .ZN(n20767) );
  OAI211_X1 U23858 ( .C1(n20855), .C2(n20778), .A(n20768), .B(n20767), .ZN(
        P2_U3132) );
  AOI22_X1 U23859 ( .A1(n20774), .A2(n20939), .B1(n20938), .B2(n20773), .ZN(
        n20770) );
  AOI22_X1 U23860 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20775), .B1(
        n20779), .B2(n20941), .ZN(n20769) );
  OAI211_X1 U23861 ( .C1(n20858), .C2(n20778), .A(n20770), .B(n20769), .ZN(
        P2_U3133) );
  AOI22_X1 U23862 ( .A1(n20774), .A2(n20945), .B1(n20944), .B2(n20773), .ZN(
        n20772) );
  AOI22_X1 U23863 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20775), .B1(
        n20779), .B2(n20947), .ZN(n20771) );
  OAI211_X1 U23864 ( .C1(n20861), .C2(n20778), .A(n20772), .B(n20771), .ZN(
        P2_U3134) );
  AOI22_X1 U23865 ( .A1(n20774), .A2(n20951), .B1(n21831), .B2(n20773), .ZN(
        n20777) );
  AOI22_X1 U23866 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20775), .B1(
        n20779), .B2(n21835), .ZN(n20776) );
  OAI211_X1 U23867 ( .C1(n20868), .C2(n20778), .A(n20777), .B(n20776), .ZN(
        P2_U3135) );
  NAND2_X1 U23868 ( .A1(n20781), .A2(n20780), .ZN(n20786) );
  AND2_X1 U23869 ( .A1(n20786), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20782) );
  NAND2_X1 U23870 ( .A1(n12426), .A2(n20782), .ZN(n20787) );
  NOR2_X1 U23871 ( .A1(n22046), .A2(n20783), .ZN(n20790) );
  INV_X1 U23872 ( .A(n20790), .ZN(n20784) );
  OAI21_X1 U23873 ( .B1(n20784), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20900), 
        .ZN(n20785) );
  INV_X1 U23874 ( .A(n20786), .ZN(n20805) );
  AOI22_X1 U23875 ( .A1(n20806), .A2(n20905), .B1(n20904), .B2(n20805), .ZN(
        n20792) );
  OAI211_X1 U23876 ( .C1(n20805), .C2(n20834), .A(n20787), .B(n20896), .ZN(
        n20788) );
  INV_X1 U23877 ( .A(n20788), .ZN(n20789) );
  OAI221_X1 U23878 ( .B1(n20790), .B2(n21043), .C1(n20790), .C2(n20894), .A(
        n20789), .ZN(n20807) );
  AOI22_X1 U23879 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20807), .B1(
        n20824), .B2(n20907), .ZN(n20791) );
  OAI211_X1 U23880 ( .C1(n20843), .C2(n20810), .A(n20792), .B(n20791), .ZN(
        P2_U3136) );
  AOI22_X1 U23881 ( .A1(n20806), .A2(n20912), .B1(n20911), .B2(n20805), .ZN(
        n20794) );
  AOI22_X1 U23882 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20807), .B1(
        n20824), .B2(n20914), .ZN(n20793) );
  OAI211_X1 U23883 ( .C1(n20846), .C2(n20810), .A(n20794), .B(n20793), .ZN(
        P2_U3137) );
  AOI22_X1 U23884 ( .A1(n20806), .A2(n20919), .B1(n20918), .B2(n20805), .ZN(
        n20796) );
  AOI22_X1 U23885 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20807), .B1(
        n20824), .B2(n20921), .ZN(n20795) );
  OAI211_X1 U23886 ( .C1(n20849), .C2(n20810), .A(n20796), .B(n20795), .ZN(
        P2_U3138) );
  AOI22_X1 U23887 ( .A1(n20806), .A2(n20926), .B1(n20925), .B2(n20805), .ZN(
        n20798) );
  AOI22_X1 U23888 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20807), .B1(
        n20824), .B2(n20928), .ZN(n20797) );
  OAI211_X1 U23889 ( .C1(n20852), .C2(n20810), .A(n20798), .B(n20797), .ZN(
        P2_U3139) );
  AOI22_X1 U23890 ( .A1(n20806), .A2(n20933), .B1(n20932), .B2(n20805), .ZN(
        n20800) );
  AOI22_X1 U23891 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20807), .B1(
        n20824), .B2(n20935), .ZN(n20799) );
  OAI211_X1 U23892 ( .C1(n20855), .C2(n20810), .A(n20800), .B(n20799), .ZN(
        P2_U3140) );
  AOI22_X1 U23893 ( .A1(n20806), .A2(n20939), .B1(n20938), .B2(n20805), .ZN(
        n20802) );
  AOI22_X1 U23894 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20807), .B1(
        n20824), .B2(n20941), .ZN(n20801) );
  OAI211_X1 U23895 ( .C1(n20858), .C2(n20810), .A(n20802), .B(n20801), .ZN(
        P2_U3141) );
  AOI22_X1 U23896 ( .A1(n20806), .A2(n20945), .B1(n20944), .B2(n20805), .ZN(
        n20804) );
  AOI22_X1 U23897 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20807), .B1(
        n20824), .B2(n20947), .ZN(n20803) );
  OAI211_X1 U23898 ( .C1(n20861), .C2(n20810), .A(n20804), .B(n20803), .ZN(
        P2_U3142) );
  AOI22_X1 U23899 ( .A1(n20806), .A2(n20951), .B1(n21831), .B2(n20805), .ZN(
        n20809) );
  AOI22_X1 U23900 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20807), .B1(
        n20824), .B2(n21835), .ZN(n20808) );
  OAI211_X1 U23901 ( .C1(n20868), .C2(n20810), .A(n20809), .B(n20808), .ZN(
        P2_U3143) );
  AOI22_X1 U23902 ( .A1(n20823), .A2(n20912), .B1(n20822), .B2(n20911), .ZN(
        n20812) );
  AOI22_X1 U23903 ( .A1(n20829), .A2(n20914), .B1(n20824), .B2(n20913), .ZN(
        n20811) );
  OAI211_X1 U23904 ( .C1(n20828), .C2(n12327), .A(n20812), .B(n20811), .ZN(
        P2_U3145) );
  INV_X1 U23905 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n20815) );
  AOI22_X1 U23906 ( .A1(n20823), .A2(n20919), .B1(n20822), .B2(n20918), .ZN(
        n20814) );
  AOI22_X1 U23907 ( .A1(n20829), .A2(n20921), .B1(n20824), .B2(n20920), .ZN(
        n20813) );
  OAI211_X1 U23908 ( .C1(n20828), .C2(n20815), .A(n20814), .B(n20813), .ZN(
        P2_U3146) );
  AOI22_X1 U23909 ( .A1(n20823), .A2(n20926), .B1(n20822), .B2(n20925), .ZN(
        n20817) );
  AOI22_X1 U23910 ( .A1(n20829), .A2(n20928), .B1(n20824), .B2(n20927), .ZN(
        n20816) );
  OAI211_X1 U23911 ( .C1(n20828), .C2(n12284), .A(n20817), .B(n20816), .ZN(
        P2_U3147) );
  AOI22_X1 U23912 ( .A1(n20823), .A2(n20939), .B1(n20822), .B2(n20938), .ZN(
        n20819) );
  AOI22_X1 U23913 ( .A1(n20829), .A2(n20941), .B1(n20824), .B2(n20940), .ZN(
        n20818) );
  OAI211_X1 U23914 ( .C1(n20828), .C2(n12439), .A(n20819), .B(n20818), .ZN(
        P2_U3149) );
  AOI22_X1 U23915 ( .A1(n20823), .A2(n20945), .B1(n20822), .B2(n20944), .ZN(
        n20821) );
  AOI22_X1 U23916 ( .A1(n20829), .A2(n20947), .B1(n20824), .B2(n20946), .ZN(
        n20820) );
  OAI211_X1 U23917 ( .C1(n20828), .C2(n12472), .A(n20821), .B(n20820), .ZN(
        P2_U3150) );
  INV_X1 U23918 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n20827) );
  AOI22_X1 U23919 ( .A1(n20823), .A2(n20951), .B1(n20822), .B2(n21831), .ZN(
        n20826) );
  AOI22_X1 U23920 ( .A1(n20829), .A2(n21835), .B1(n20824), .B2(n21834), .ZN(
        n20825) );
  OAI211_X1 U23921 ( .C1(n20828), .C2(n20827), .A(n20826), .B(n20825), .ZN(
        P2_U3151) );
  INV_X1 U23922 ( .A(n20862), .ZN(n20830) );
  AND2_X1 U23923 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n20830), .ZN(n20831) );
  NAND2_X1 U23924 ( .A1(n20832), .A2(n20831), .ZN(n20838) );
  OAI21_X1 U23925 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20836), .A(n20900), 
        .ZN(n20833) );
  AOI22_X1 U23926 ( .A1(n20863), .A2(n20905), .B1(n20904), .B2(n20862), .ZN(
        n20842) );
  NAND3_X1 U23927 ( .A1(n20894), .A2(n20835), .A3(n20834), .ZN(n20837) );
  NAND2_X1 U23928 ( .A1(n20837), .A2(n20836), .ZN(n20840) );
  NAND4_X1 U23929 ( .A1(n20840), .A2(n20839), .A3(n20896), .A4(n20838), .ZN(
        n20864) );
  AOI22_X1 U23930 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20864), .B1(
        n20886), .B2(n20907), .ZN(n20841) );
  OAI211_X1 U23931 ( .C1(n20843), .C2(n20867), .A(n20842), .B(n20841), .ZN(
        P2_U3152) );
  AOI22_X1 U23932 ( .A1(n20863), .A2(n20912), .B1(n20911), .B2(n20862), .ZN(
        n20845) );
  AOI22_X1 U23933 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20864), .B1(
        n20886), .B2(n20914), .ZN(n20844) );
  OAI211_X1 U23934 ( .C1(n20846), .C2(n20867), .A(n20845), .B(n20844), .ZN(
        P2_U3153) );
  AOI22_X1 U23935 ( .A1(n20863), .A2(n20919), .B1(n20918), .B2(n20862), .ZN(
        n20848) );
  AOI22_X1 U23936 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20864), .B1(
        n20886), .B2(n20921), .ZN(n20847) );
  OAI211_X1 U23937 ( .C1(n20849), .C2(n20867), .A(n20848), .B(n20847), .ZN(
        P2_U3154) );
  AOI22_X1 U23938 ( .A1(n20863), .A2(n20926), .B1(n20925), .B2(n20862), .ZN(
        n20851) );
  AOI22_X1 U23939 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20864), .B1(
        n20886), .B2(n20928), .ZN(n20850) );
  OAI211_X1 U23940 ( .C1(n20852), .C2(n20867), .A(n20851), .B(n20850), .ZN(
        P2_U3155) );
  AOI22_X1 U23941 ( .A1(n20863), .A2(n20933), .B1(n20932), .B2(n20862), .ZN(
        n20854) );
  AOI22_X1 U23942 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20864), .B1(
        n20886), .B2(n20935), .ZN(n20853) );
  OAI211_X1 U23943 ( .C1(n20855), .C2(n20867), .A(n20854), .B(n20853), .ZN(
        P2_U3156) );
  AOI22_X1 U23944 ( .A1(n20863), .A2(n20939), .B1(n20938), .B2(n20862), .ZN(
        n20857) );
  AOI22_X1 U23945 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20864), .B1(
        n20886), .B2(n20941), .ZN(n20856) );
  OAI211_X1 U23946 ( .C1(n20858), .C2(n20867), .A(n20857), .B(n20856), .ZN(
        P2_U3157) );
  AOI22_X1 U23947 ( .A1(n20863), .A2(n20945), .B1(n20944), .B2(n20862), .ZN(
        n20860) );
  AOI22_X1 U23948 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20864), .B1(
        n20886), .B2(n20947), .ZN(n20859) );
  OAI211_X1 U23949 ( .C1(n20861), .C2(n20867), .A(n20860), .B(n20859), .ZN(
        P2_U3158) );
  AOI22_X1 U23950 ( .A1(n20863), .A2(n20951), .B1(n21831), .B2(n20862), .ZN(
        n20866) );
  AOI22_X1 U23951 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20864), .B1(
        n20886), .B2(n21835), .ZN(n20865) );
  OAI211_X1 U23952 ( .C1(n20868), .C2(n20867), .A(n20866), .B(n20865), .ZN(
        P2_U3159) );
  AOI22_X1 U23953 ( .A1(n20913), .A2(n20886), .B1(n20885), .B2(n20911), .ZN(
        n20870) );
  AOI22_X1 U23954 ( .A1(n20912), .A2(n20887), .B1(n20953), .B2(n20914), .ZN(
        n20869) );
  OAI211_X1 U23955 ( .C1(n20891), .C2(n12332), .A(n20870), .B(n20869), .ZN(
        P2_U3161) );
  INV_X1 U23956 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n20873) );
  AOI22_X1 U23957 ( .A1(n20921), .A2(n20953), .B1(n20885), .B2(n20918), .ZN(
        n20872) );
  AOI22_X1 U23958 ( .A1(n20919), .A2(n20887), .B1(n20886), .B2(n20920), .ZN(
        n20871) );
  OAI211_X1 U23959 ( .C1(n20891), .C2(n20873), .A(n20872), .B(n20871), .ZN(
        P2_U3162) );
  INV_X1 U23960 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n20876) );
  AOI22_X1 U23961 ( .A1(n20928), .A2(n20953), .B1(n20885), .B2(n20925), .ZN(
        n20875) );
  AOI22_X1 U23962 ( .A1(n20926), .A2(n20887), .B1(n20886), .B2(n20927), .ZN(
        n20874) );
  OAI211_X1 U23963 ( .C1(n20891), .C2(n20876), .A(n20875), .B(n20874), .ZN(
        P2_U3163) );
  AOI22_X1 U23964 ( .A1(n20934), .A2(n20886), .B1(n20932), .B2(n20885), .ZN(
        n20878) );
  AOI22_X1 U23965 ( .A1(n20933), .A2(n20887), .B1(n20953), .B2(n20935), .ZN(
        n20877) );
  OAI211_X1 U23966 ( .C1(n20891), .C2(n20879), .A(n20878), .B(n20877), .ZN(
        P2_U3164) );
  AOI22_X1 U23967 ( .A1(n20940), .A2(n20886), .B1(n20885), .B2(n20938), .ZN(
        n20881) );
  AOI22_X1 U23968 ( .A1(n20939), .A2(n20887), .B1(n20953), .B2(n20941), .ZN(
        n20880) );
  OAI211_X1 U23969 ( .C1(n20891), .C2(n12443), .A(n20881), .B(n20880), .ZN(
        P2_U3165) );
  INV_X1 U23970 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n20884) );
  AOI22_X1 U23971 ( .A1(n20947), .A2(n20953), .B1(n20885), .B2(n20944), .ZN(
        n20883) );
  AOI22_X1 U23972 ( .A1(n20945), .A2(n20887), .B1(n20886), .B2(n20946), .ZN(
        n20882) );
  OAI211_X1 U23973 ( .C1(n20891), .C2(n20884), .A(n20883), .B(n20882), .ZN(
        P2_U3166) );
  INV_X1 U23974 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n20890) );
  AOI22_X1 U23975 ( .A1(n21834), .A2(n20886), .B1(n20885), .B2(n21831), .ZN(
        n20889) );
  AOI22_X1 U23976 ( .A1(n20951), .A2(n20887), .B1(n20953), .B2(n21835), .ZN(
        n20888) );
  OAI211_X1 U23977 ( .C1(n20891), .C2(n20890), .A(n20889), .B(n20888), .ZN(
        P2_U3167) );
  NOR2_X1 U23978 ( .A1(n21054), .A2(n20892), .ZN(n20899) );
  AOI21_X1 U23979 ( .B1(n20894), .B2(n20893), .A(n20899), .ZN(n20898) );
  NOR2_X1 U23980 ( .A1(n20950), .A2(n20900), .ZN(n20895) );
  OAI211_X1 U23981 ( .C1(n20950), .C2(n20834), .A(n20903), .B(n20896), .ZN(
        n20897) );
  INV_X1 U23982 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n20910) );
  INV_X1 U23983 ( .A(n20899), .ZN(n20901) );
  OAI21_X1 U23984 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20901), .A(n20900), 
        .ZN(n20902) );
  AOI22_X1 U23985 ( .A1(n20952), .A2(n20905), .B1(n20904), .B2(n20950), .ZN(
        n20909) );
  AOI22_X1 U23986 ( .A1(n20954), .A2(n20907), .B1(n20953), .B2(n20906), .ZN(
        n20908) );
  OAI211_X1 U23987 ( .C1(n20957), .C2(n20910), .A(n20909), .B(n20908), .ZN(
        P2_U3168) );
  AOI22_X1 U23988 ( .A1(n20952), .A2(n20912), .B1(n20911), .B2(n20950), .ZN(
        n20916) );
  AOI22_X1 U23989 ( .A1(n20954), .A2(n20914), .B1(n20953), .B2(n20913), .ZN(
        n20915) );
  OAI211_X1 U23990 ( .C1(n20957), .C2(n20917), .A(n20916), .B(n20915), .ZN(
        P2_U3169) );
  INV_X1 U23991 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n20924) );
  AOI22_X1 U23992 ( .A1(n20952), .A2(n20919), .B1(n20918), .B2(n20950), .ZN(
        n20923) );
  AOI22_X1 U23993 ( .A1(n20954), .A2(n20921), .B1(n20953), .B2(n20920), .ZN(
        n20922) );
  OAI211_X1 U23994 ( .C1(n20957), .C2(n20924), .A(n20923), .B(n20922), .ZN(
        P2_U3170) );
  INV_X1 U23995 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n20931) );
  AOI22_X1 U23996 ( .A1(n20952), .A2(n20926), .B1(n20925), .B2(n20950), .ZN(
        n20930) );
  AOI22_X1 U23997 ( .A1(n20954), .A2(n20928), .B1(n20953), .B2(n20927), .ZN(
        n20929) );
  OAI211_X1 U23998 ( .C1(n20957), .C2(n20931), .A(n20930), .B(n20929), .ZN(
        P2_U3171) );
  AOI22_X1 U23999 ( .A1(n20952), .A2(n20933), .B1(n20932), .B2(n20950), .ZN(
        n20937) );
  AOI22_X1 U24000 ( .A1(n20954), .A2(n20935), .B1(n20953), .B2(n20934), .ZN(
        n20936) );
  OAI211_X1 U24001 ( .C1(n20957), .C2(n12406), .A(n20937), .B(n20936), .ZN(
        P2_U3172) );
  AOI22_X1 U24002 ( .A1(n20952), .A2(n20939), .B1(n20938), .B2(n20950), .ZN(
        n20943) );
  AOI22_X1 U24003 ( .A1(n20954), .A2(n20941), .B1(n20953), .B2(n20940), .ZN(
        n20942) );
  OAI211_X1 U24004 ( .C1(n20957), .C2(n12458), .A(n20943), .B(n20942), .ZN(
        P2_U3173) );
  AOI22_X1 U24005 ( .A1(n20952), .A2(n20945), .B1(n20944), .B2(n20950), .ZN(
        n20949) );
  AOI22_X1 U24006 ( .A1(n20954), .A2(n20947), .B1(n20953), .B2(n20946), .ZN(
        n20948) );
  OAI211_X1 U24007 ( .C1(n20957), .C2(n12491), .A(n20949), .B(n20948), .ZN(
        P2_U3174) );
  AOI22_X1 U24008 ( .A1(n20952), .A2(n20951), .B1(n21831), .B2(n20950), .ZN(
        n20956) );
  AOI22_X1 U24009 ( .A1(n20954), .A2(n21835), .B1(n20953), .B2(n21834), .ZN(
        n20955) );
  OAI211_X1 U24010 ( .C1(n20957), .C2(n15319), .A(n20956), .B(n20955), .ZN(
        P2_U3175) );
  AND2_X1 U24011 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n20958), .ZN(
        P2_U3179) );
  AND2_X1 U24012 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n20958), .ZN(
        P2_U3180) );
  AND2_X1 U24013 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n20958), .ZN(
        P2_U3181) );
  AND2_X1 U24014 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n20958), .ZN(
        P2_U3182) );
  AND2_X1 U24015 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n20958), .ZN(
        P2_U3183) );
  AND2_X1 U24016 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20958), .ZN(
        P2_U3184) );
  NOR2_X1 U24017 ( .A1(n22129), .A2(n21040), .ZN(P2_U3185) );
  AND2_X1 U24018 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n20958), .ZN(
        P2_U3186) );
  AND2_X1 U24019 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20958), .ZN(
        P2_U3187) );
  AND2_X1 U24020 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n20958), .ZN(
        P2_U3188) );
  AND2_X1 U24021 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20958), .ZN(
        P2_U3189) );
  AND2_X1 U24022 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20958), .ZN(
        P2_U3190) );
  AND2_X1 U24023 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20958), .ZN(
        P2_U3191) );
  AND2_X1 U24024 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n20958), .ZN(
        P2_U3192) );
  AND2_X1 U24025 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n20958), .ZN(
        P2_U3193) );
  AND2_X1 U24026 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n20958), .ZN(
        P2_U3194) );
  AND2_X1 U24027 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n20958), .ZN(
        P2_U3195) );
  AND2_X1 U24028 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n20958), .ZN(
        P2_U3196) );
  AND2_X1 U24029 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n20958), .ZN(
        P2_U3197) );
  AND2_X1 U24030 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n20958), .ZN(
        P2_U3198) );
  INV_X1 U24031 ( .A(P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n22128) );
  NOR2_X1 U24032 ( .A1(n22128), .A2(n21040), .ZN(P2_U3199) );
  AND2_X1 U24033 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n20958), .ZN(
        P2_U3200) );
  NOR2_X1 U24034 ( .A1(n21968), .A2(n21040), .ZN(P2_U3201) );
  AND2_X1 U24035 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n20958), .ZN(P2_U3202) );
  AND2_X1 U24036 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n20958), .ZN(P2_U3203) );
  AND2_X1 U24037 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20958), .ZN(P2_U3204) );
  AND2_X1 U24038 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n20958), .ZN(P2_U3205) );
  AND2_X1 U24039 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n20958), .ZN(P2_U3206) );
  AND2_X1 U24040 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n20958), .ZN(P2_U3207) );
  AND2_X1 U24041 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n20958), .ZN(P2_U3208) );
  INV_X1 U24042 ( .A(NA), .ZN(n21746) );
  OAI21_X1 U24043 ( .B1(n21746), .B2(n20966), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n20975) );
  INV_X1 U24044 ( .A(n20975), .ZN(n20963) );
  NAND2_X1 U24045 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20959), .ZN(n20973) );
  AND3_X1 U24046 ( .A1(n20973), .A2(P2_REQUESTPENDING_REG_SCAN_IN), .A3(
        P2_STATE_REG_0__SCAN_IN), .ZN(n20962) );
  INV_X1 U24047 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20960) );
  OAI211_X1 U24048 ( .C1(HOLD), .C2(n20960), .A(n21095), .B(n20970), .ZN(
        n20961) );
  OAI21_X1 U24049 ( .B1(n20963), .B2(n20962), .A(n20961), .ZN(P2_U3209) );
  AND2_X1 U24050 ( .A1(n20964), .A2(n20973), .ZN(n20968) );
  NOR2_X1 U24051 ( .A1(HOLD), .A2(n20965), .ZN(n20974) );
  OAI211_X1 U24052 ( .C1(n20974), .C2(n20977), .A(
        P2_REQUESTPENDING_REG_SCAN_IN), .B(n20966), .ZN(n20967) );
  OAI211_X1 U24053 ( .C1(n20969), .C2(n21742), .A(n20968), .B(n20967), .ZN(
        P2_U3210) );
  OAI22_X1 U24054 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n20970), .B1(NA), 
        .B2(n20973), .ZN(n20971) );
  OAI211_X1 U24055 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n20971), .ZN(n20972) );
  OAI221_X1 U24056 ( .B1(n20975), .B2(n20974), .C1(n20975), .C2(n20973), .A(
        n20972), .ZN(P2_U3211) );
  OAI222_X1 U24057 ( .A1(n21030), .A2(n20979), .B1(n20978), .B2(n20976), .C1(
        n20981), .C2(n21033), .ZN(P2_U3212) );
  OAI222_X1 U24058 ( .A1(n21030), .A2(n20981), .B1(n20980), .B2(n20976), .C1(
        n20983), .C2(n21033), .ZN(P2_U3213) );
  OAI222_X1 U24059 ( .A1(n21030), .A2(n20983), .B1(n20982), .B2(n20976), .C1(
        n20984), .C2(n21033), .ZN(P2_U3214) );
  OAI222_X1 U24060 ( .A1(n21033), .A2(n20986), .B1(n20985), .B2(n20976), .C1(
        n20984), .C2(n21030), .ZN(P2_U3215) );
  OAI222_X1 U24061 ( .A1(n21033), .A2(n20988), .B1(n20987), .B2(n20976), .C1(
        n20986), .C2(n21030), .ZN(P2_U3216) );
  OAI222_X1 U24062 ( .A1(n21033), .A2(n20990), .B1(n20989), .B2(n20976), .C1(
        n20988), .C2(n21030), .ZN(P2_U3217) );
  INV_X1 U24063 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n20992) );
  OAI222_X1 U24064 ( .A1(n21033), .A2(n20992), .B1(n20991), .B2(n20976), .C1(
        n20990), .C2(n21030), .ZN(P2_U3218) );
  INV_X1 U24065 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n20994) );
  OAI222_X1 U24066 ( .A1(n21033), .A2(n20994), .B1(n20993), .B2(n20976), .C1(
        n20992), .C2(n21030), .ZN(P2_U3219) );
  OAI222_X1 U24067 ( .A1(n21033), .A2(n17171), .B1(n20995), .B2(n20976), .C1(
        n20994), .C2(n21030), .ZN(P2_U3220) );
  OAI222_X1 U24068 ( .A1(n21033), .A2(n17159), .B1(n20996), .B2(n20976), .C1(
        n17171), .C2(n21030), .ZN(P2_U3221) );
  INV_X1 U24069 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n20998) );
  OAI222_X1 U24070 ( .A1(n21033), .A2(n20998), .B1(n20997), .B2(n20976), .C1(
        n17159), .C2(n21030), .ZN(P2_U3222) );
  OAI222_X1 U24071 ( .A1(n21033), .A2(n21000), .B1(n20999), .B2(n20976), .C1(
        n20998), .C2(n21030), .ZN(P2_U3223) );
  OAI222_X1 U24072 ( .A1(n21033), .A2(n17125), .B1(n21001), .B2(n20976), .C1(
        n21000), .C2(n21030), .ZN(P2_U3224) );
  OAI222_X1 U24073 ( .A1(n21033), .A2(n21003), .B1(n21002), .B2(n20976), .C1(
        n17125), .C2(n21030), .ZN(P2_U3225) );
  OAI222_X1 U24074 ( .A1(n21033), .A2(n21005), .B1(n21004), .B2(n20976), .C1(
        n21003), .C2(n21030), .ZN(P2_U3226) );
  OAI222_X1 U24075 ( .A1(n21033), .A2(n21007), .B1(n21006), .B2(n20976), .C1(
        n21005), .C2(n21030), .ZN(P2_U3227) );
  OAI222_X1 U24076 ( .A1(n21033), .A2(n17081), .B1(n21008), .B2(n20976), .C1(
        n21007), .C2(n21030), .ZN(P2_U3228) );
  OAI222_X1 U24077 ( .A1(n21033), .A2(n21010), .B1(n21009), .B2(n20976), .C1(
        n17081), .C2(n21030), .ZN(P2_U3229) );
  OAI222_X1 U24078 ( .A1(n21033), .A2(n16540), .B1(n21011), .B2(n20976), .C1(
        n21010), .C2(n21030), .ZN(P2_U3230) );
  INV_X1 U24079 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n21013) );
  OAI222_X1 U24080 ( .A1(n21033), .A2(n21013), .B1(n21012), .B2(n20976), .C1(
        n16540), .C2(n21030), .ZN(P2_U3231) );
  OAI222_X1 U24081 ( .A1(n21033), .A2(n21015), .B1(n21014), .B2(n20976), .C1(
        n21013), .C2(n21030), .ZN(P2_U3232) );
  OAI222_X1 U24082 ( .A1(n21033), .A2(n21017), .B1(n21016), .B2(n20976), .C1(
        n21015), .C2(n21030), .ZN(P2_U3233) );
  OAI222_X1 U24083 ( .A1(n21033), .A2(n21019), .B1(n21018), .B2(n20976), .C1(
        n21017), .C2(n21030), .ZN(P2_U3234) );
  OAI222_X1 U24084 ( .A1(n21033), .A2(n21021), .B1(n21020), .B2(n20976), .C1(
        n21019), .C2(n21030), .ZN(P2_U3235) );
  OAI222_X1 U24085 ( .A1(n21033), .A2(n21023), .B1(n21022), .B2(n20976), .C1(
        n21021), .C2(n21030), .ZN(P2_U3236) );
  OAI222_X1 U24086 ( .A1(n21033), .A2(n21967), .B1(n21024), .B2(n20976), .C1(
        n21023), .C2(n21030), .ZN(P2_U3237) );
  OAI222_X1 U24087 ( .A1(n21030), .A2(n21967), .B1(n21025), .B2(n20976), .C1(
        n21026), .C2(n21033), .ZN(P2_U3238) );
  OAI222_X1 U24088 ( .A1(n21033), .A2(n21028), .B1(n21027), .B2(n20976), .C1(
        n21026), .C2(n21030), .ZN(P2_U3239) );
  INV_X1 U24089 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n21031) );
  OAI222_X1 U24090 ( .A1(n21033), .A2(n21031), .B1(n21029), .B2(n20976), .C1(
        n21028), .C2(n21030), .ZN(P2_U3240) );
  OAI222_X1 U24091 ( .A1(n21033), .A2(n13395), .B1(n21032), .B2(n20976), .C1(
        n21031), .C2(n21030), .ZN(P2_U3241) );
  OAI22_X1 U24092 ( .A1(n21095), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n20976), .ZN(n21034) );
  INV_X1 U24093 ( .A(n21034), .ZN(P2_U3585) );
  MUX2_X1 U24094 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n21095), .Z(P2_U3586) );
  OAI22_X1 U24095 ( .A1(n21095), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n20976), .ZN(n21035) );
  INV_X1 U24096 ( .A(n21035), .ZN(P2_U3587) );
  OAI22_X1 U24097 ( .A1(n21095), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n20976), .ZN(n21036) );
  INV_X1 U24098 ( .A(n21036), .ZN(P2_U3588) );
  OAI21_X1 U24099 ( .B1(n21040), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n21038), 
        .ZN(n21037) );
  INV_X1 U24100 ( .A(n21037), .ZN(P2_U3591) );
  OAI21_X1 U24101 ( .B1(n21040), .B2(n21039), .A(n21038), .ZN(P2_U3592) );
  INV_X1 U24102 ( .A(n21084), .ZN(n21075) );
  NAND2_X1 U24103 ( .A1(n21041), .A2(n21042), .ZN(n21050) );
  AND2_X1 U24104 ( .A1(n21042), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n21066) );
  NAND2_X1 U24105 ( .A1(n21043), .A2(n21066), .ZN(n21061) );
  AND2_X1 U24106 ( .A1(n21055), .A2(n21044), .ZN(n21068) );
  AOI21_X1 U24107 ( .B1(n21045), .B2(n21055), .A(n21068), .ZN(n21046) );
  NAND2_X1 U24108 ( .A1(n21061), .A2(n21046), .ZN(n21048) );
  NAND2_X1 U24109 ( .A1(n21048), .A2(n21047), .ZN(n21049) );
  OAI211_X1 U24110 ( .C1(n21051), .C2(n20834), .A(n21050), .B(n21049), .ZN(
        n21052) );
  INV_X1 U24111 ( .A(n21052), .ZN(n21053) );
  AOI22_X1 U24112 ( .A1(n21075), .A2(n21054), .B1(n21053), .B2(n21084), .ZN(
        P2_U3602) );
  INV_X1 U24113 ( .A(n21055), .ZN(n21078) );
  INV_X1 U24114 ( .A(n21068), .ZN(n21057) );
  OAI22_X1 U24115 ( .A1(n21058), .A2(n21057), .B1(n21056), .B2(n20834), .ZN(
        n21059) );
  INV_X1 U24116 ( .A(n21059), .ZN(n21060) );
  OAI211_X1 U24117 ( .C1(n21078), .C2(n21062), .A(n21061), .B(n21060), .ZN(
        n21063) );
  INV_X1 U24118 ( .A(n21063), .ZN(n21064) );
  AOI22_X1 U24119 ( .A1(n21075), .A2(n21065), .B1(n21064), .B2(n21084), .ZN(
        P2_U3603) );
  INV_X1 U24120 ( .A(n21066), .ZN(n21071) );
  NAND2_X1 U24121 ( .A1(n21067), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n21070) );
  NAND2_X1 U24122 ( .A1(n21072), .A2(n21068), .ZN(n21069) );
  OAI211_X1 U24123 ( .C1(n21072), .C2(n21071), .A(n21070), .B(n21069), .ZN(
        n21073) );
  INV_X1 U24124 ( .A(n21073), .ZN(n21074) );
  AOI22_X1 U24125 ( .A1(n21075), .A2(n22046), .B1(n21074), .B2(n21084), .ZN(
        P2_U3604) );
  NAND3_X1 U24126 ( .A1(n21076), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n21077) );
  OAI21_X1 U24127 ( .B1(n21079), .B2(n21078), .A(n21077), .ZN(n21081) );
  OAI21_X1 U24128 ( .B1(n21081), .B2(n21080), .A(n21084), .ZN(n21082) );
  OAI21_X1 U24129 ( .B1(n21084), .B2(n21083), .A(n21082), .ZN(P2_U3605) );
  INV_X1 U24130 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n21085) );
  AOI22_X1 U24131 ( .A1(n20976), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n21085), 
        .B2(n21095), .ZN(P2_U3608) );
  INV_X1 U24132 ( .A(n21086), .ZN(n21091) );
  NAND3_X1 U24133 ( .A1(n21089), .A2(n21088), .A3(n21087), .ZN(n21090) );
  NAND2_X1 U24134 ( .A1(n21091), .A2(n21090), .ZN(n21093) );
  MUX2_X1 U24135 ( .A(P2_MORE_REG_SCAN_IN), .B(n21093), .S(n21092), .Z(
        P2_U3609) );
  OAI22_X1 U24136 ( .A1(n21095), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n20976), .ZN(n21096) );
  INV_X1 U24137 ( .A(n21096), .ZN(P2_U3611) );
  OAI21_X1 U24138 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(n21097), .A(
        P1_STATE_REG_0__SCAN_IN), .ZN(n21749) );
  NOR2_X2 U24139 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21097), .ZN(n21817) );
  INV_X2 U24140 ( .A(n21817), .ZN(n21815) );
  OAI21_X1 U24141 ( .B1(n21749), .B2(P1_ADS_N_REG_SCAN_IN), .A(n21815), .ZN(
        n21098) );
  INV_X1 U24142 ( .A(n21098), .ZN(P1_U2802) );
  OAI21_X1 U24143 ( .B1(n21100), .B2(n21099), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n21101) );
  OAI21_X1 U24144 ( .B1(n21102), .B2(n21733), .A(n21101), .ZN(P1_U2803) );
  NOR2_X1 U24145 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n21104) );
  OAI21_X1 U24146 ( .B1(n21104), .B2(P1_D_C_N_REG_SCAN_IN), .A(n21815), .ZN(
        n21103) );
  OAI21_X1 U24147 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n21815), .A(n21103), 
        .ZN(P1_U2804) );
  INV_X1 U24148 ( .A(n21736), .ZN(n21798) );
  OAI21_X1 U24149 ( .B1(BS16), .B2(n21104), .A(n21798), .ZN(n21796) );
  OAI21_X1 U24150 ( .B1(n21798), .B2(n21528), .A(n21796), .ZN(P1_U2805) );
  INV_X1 U24151 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n21106) );
  OAI21_X1 U24152 ( .B1(n21107), .B2(n21106), .A(n21105), .ZN(P1_U2806) );
  NOR4_X1 U24153 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_19__SCAN_IN), .A3(P1_DATAWIDTH_REG_20__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_21__SCAN_IN), .ZN(n21111) );
  NOR4_X1 U24154 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_15__SCAN_IN), .A3(P1_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_17__SCAN_IN), .ZN(n21110) );
  NOR4_X1 U24155 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n21109) );
  NOR4_X1 U24156 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_23__SCAN_IN), .A3(P1_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n21108) );
  NAND4_X1 U24157 ( .A1(n21111), .A2(n21110), .A3(n21109), .A4(n21108), .ZN(
        n21117) );
  NOR4_X1 U24158 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_3__SCAN_IN), .A3(P1_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_5__SCAN_IN), .ZN(n21115) );
  AOI211_X1 U24159 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_28__SCAN_IN), .B(
        P1_DATAWIDTH_REG_24__SCAN_IN), .ZN(n21114) );
  NOR4_X1 U24160 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_11__SCAN_IN), .A3(P1_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_13__SCAN_IN), .ZN(n21113) );
  NOR4_X1 U24161 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_7__SCAN_IN), .A3(P1_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_9__SCAN_IN), .ZN(n21112) );
  NAND4_X1 U24162 ( .A1(n21115), .A2(n21114), .A3(n21113), .A4(n21112), .ZN(
        n21116) );
  NOR2_X1 U24163 ( .A1(n21117), .A2(n21116), .ZN(n21810) );
  INV_X1 U24164 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n21119) );
  NOR3_X1 U24165 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n21120) );
  OAI21_X1 U24166 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n21120), .A(n21810), .ZN(
        n21118) );
  OAI21_X1 U24167 ( .B1(n21810), .B2(n21119), .A(n21118), .ZN(P1_U2807) );
  INV_X1 U24168 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21797) );
  AOI21_X1 U24169 ( .B1(n21806), .B2(n21797), .A(n21120), .ZN(n21122) );
  INV_X1 U24170 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21121) );
  INV_X1 U24171 ( .A(n21810), .ZN(n21813) );
  AOI22_X1 U24172 ( .A1(n21810), .A2(n21122), .B1(n21121), .B2(n21813), .ZN(
        P1_U2808) );
  NAND2_X1 U24173 ( .A1(n21210), .A2(n21125), .ZN(n21187) );
  NAND2_X1 U24174 ( .A1(n21187), .A2(n21123), .ZN(n21191) );
  AOI21_X1 U24175 ( .B1(n21210), .B2(n21124), .A(n21191), .ZN(n21151) );
  NOR2_X1 U24176 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n21124), .ZN(n21132) );
  NOR2_X1 U24177 ( .A1(n21126), .A2(n21125), .ZN(n21174) );
  INV_X1 U24178 ( .A(n21127), .ZN(n21128) );
  AOI22_X1 U24179 ( .A1(n21173), .A2(P1_EBX_REG_9__SCAN_IN), .B1(n21209), .B2(
        n21128), .ZN(n21129) );
  OAI211_X1 U24180 ( .C1(n21203), .C2(n21130), .A(n21129), .B(n21291), .ZN(
        n21131) );
  AOI21_X1 U24181 ( .B1(n21132), .B2(n21174), .A(n21131), .ZN(n21137) );
  INV_X1 U24182 ( .A(n21133), .ZN(n21135) );
  AOI22_X1 U24183 ( .A1(n21135), .A2(n21168), .B1(n21146), .B2(n21134), .ZN(
        n21136) );
  OAI211_X1 U24184 ( .C1(n21151), .C2(n21138), .A(n21137), .B(n21136), .ZN(
        P1_U2831) );
  NAND3_X1 U24185 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .ZN(n21139) );
  NOR2_X1 U24186 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n21139), .ZN(n21140) );
  AOI22_X1 U24187 ( .A1(n21174), .A2(n21140), .B1(P1_EBX_REG_8__SCAN_IN), .B2(
        n21173), .ZN(n21141) );
  OAI21_X1 U24188 ( .B1(n21143), .B2(n21142), .A(n21141), .ZN(n21144) );
  AOI211_X1 U24189 ( .C1(n21190), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n21189), .B(n21144), .ZN(n21150) );
  INV_X1 U24190 ( .A(n21145), .ZN(n21147) );
  AOI22_X1 U24191 ( .A1(n21148), .A2(n21168), .B1(n21147), .B2(n21146), .ZN(
        n21149) );
  OAI211_X1 U24192 ( .C1(n21151), .C2(n16006), .A(n21150), .B(n21149), .ZN(
        P1_U2832) );
  INV_X1 U24193 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n21759) );
  OR2_X1 U24194 ( .A1(n21759), .A2(n21757), .ZN(n21157) );
  NOR2_X1 U24195 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n21157), .ZN(n21156) );
  AOI22_X1 U24196 ( .A1(n21173), .A2(P1_EBX_REG_7__SCAN_IN), .B1(n21209), .B2(
        n21152), .ZN(n21153) );
  OAI211_X1 U24197 ( .C1(n21203), .C2(n21154), .A(n21153), .B(n21291), .ZN(
        n21155) );
  AOI21_X1 U24198 ( .B1(n21156), .B2(n21174), .A(n21155), .ZN(n21161) );
  AND2_X1 U24199 ( .A1(n21210), .A2(n21157), .ZN(n21158) );
  OR2_X1 U24200 ( .A1(n21191), .A2(n21158), .ZN(n21167) );
  AOI22_X1 U24201 ( .A1(n21159), .A2(n21168), .B1(P1_REIP_REG_7__SCAN_IN), 
        .B2(n21167), .ZN(n21160) );
  OAI211_X1 U24202 ( .C1(n21162), .C2(n9710), .A(n21161), .B(n21160), .ZN(
        P1_U2833) );
  NAND2_X1 U24203 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n21174), .ZN(n21165) );
  AOI22_X1 U24204 ( .A1(n21173), .A2(P1_EBX_REG_6__SCAN_IN), .B1(n21209), .B2(
        n21163), .ZN(n21164) );
  OAI21_X1 U24205 ( .B1(P1_REIP_REG_6__SCAN_IN), .B2(n21165), .A(n21164), .ZN(
        n21166) );
  AOI211_X1 U24206 ( .C1(n21190), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n21189), .B(n21166), .ZN(n21171) );
  AOI22_X1 U24207 ( .A1(n21169), .A2(n21168), .B1(P1_REIP_REG_6__SCAN_IN), 
        .B2(n21167), .ZN(n21170) );
  OAI211_X1 U24208 ( .C1(n21172), .C2(n9710), .A(n21171), .B(n21170), .ZN(
        P1_U2834) );
  AOI22_X1 U24209 ( .A1(n21174), .A2(n21757), .B1(n21173), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n21181) );
  AOI22_X1 U24210 ( .A1(n21209), .A2(n21175), .B1(P1_REIP_REG_5__SCAN_IN), 
        .B2(n21191), .ZN(n21177) );
  AOI21_X1 U24211 ( .B1(n21190), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n21189), .ZN(n21176) );
  OAI211_X1 U24212 ( .C1(n21215), .C2(n21178), .A(n21177), .B(n21176), .ZN(
        n21179) );
  INV_X1 U24213 ( .A(n21179), .ZN(n21180) );
  OAI211_X1 U24214 ( .C1(n21182), .C2(n9710), .A(n21181), .B(n21180), .ZN(
        P1_U2835) );
  NAND3_X1 U24215 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n21186) );
  INV_X1 U24216 ( .A(n21183), .ZN(n21185) );
  OAI22_X1 U24217 ( .A1(n21187), .A2(n21186), .B1(n21185), .B2(n21184), .ZN(
        n21188) );
  AOI211_X1 U24218 ( .C1(n21190), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n21189), .B(n21188), .ZN(n21199) );
  INV_X1 U24219 ( .A(n21191), .ZN(n21193) );
  INV_X1 U24220 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n22126) );
  OAI22_X1 U24221 ( .A1(n21193), .A2(n22126), .B1(n21192), .B2(n21205), .ZN(
        n21197) );
  OAI22_X1 U24222 ( .A1(n21195), .A2(n21215), .B1(n21194), .B2(n9710), .ZN(
        n21196) );
  AOI211_X1 U24223 ( .C1(n21209), .C2(n21281), .A(n21197), .B(n21196), .ZN(
        n21198) );
  NAND2_X1 U24224 ( .A1(n21199), .A2(n21198), .ZN(P1_U2836) );
  AOI221_X1 U24225 ( .B1(n21806), .B2(n21210), .C1(n21201), .C2(n21210), .A(
        n21200), .ZN(n21223) );
  INV_X1 U24226 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n21755) );
  OAI22_X1 U24227 ( .A1(n21205), .A2(n21204), .B1(n21203), .B2(n21202), .ZN(
        n21206) );
  INV_X1 U24228 ( .A(n21206), .ZN(n21214) );
  NAND2_X1 U24229 ( .A1(n21207), .A2(n21310), .ZN(n21213) );
  NAND2_X1 U24230 ( .A1(n21209), .A2(n21208), .ZN(n21212) );
  NAND4_X1 U24231 ( .A1(n21210), .A2(n21755), .A3(P1_REIP_REG_2__SCAN_IN), 
        .A4(P1_REIP_REG_1__SCAN_IN), .ZN(n21211) );
  AND4_X1 U24232 ( .A1(n21214), .A2(n21213), .A3(n21212), .A4(n21211), .ZN(
        n21222) );
  INV_X1 U24233 ( .A(n21215), .ZN(n21219) );
  NOR2_X1 U24234 ( .A1(n9710), .A2(n21216), .ZN(n21218) );
  AOI21_X1 U24235 ( .B1(n21220), .B2(n21219), .A(n21218), .ZN(n21221) );
  OAI211_X1 U24236 ( .C1(n21223), .C2(n21755), .A(n21222), .B(n21221), .ZN(
        P1_U2837) );
  INV_X1 U24237 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n21882) );
  AOI22_X1 U24238 ( .A1(n21225), .A2(P1_EAX_REG_30__SCAN_IN), .B1(n21254), 
        .B2(P1_UWORD_REG_14__SCAN_IN), .ZN(n21224) );
  OAI21_X1 U24239 ( .B1(n21882), .B2(n21237), .A(n21224), .ZN(P1_U2906) );
  INV_X1 U24240 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n22066) );
  AOI22_X1 U24241 ( .A1(n21225), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n21254), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n21226) );
  OAI21_X1 U24242 ( .B1(n22066), .B2(n21237), .A(n21226), .ZN(P1_U2919) );
  OAI222_X1 U24243 ( .A1(n21229), .A2(n21821), .B1(n21256), .B2(n21228), .C1(
        n21237), .C2(n21227), .ZN(P1_U2921) );
  AOI22_X1 U24244 ( .A1(n21234), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n21231), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n21230) );
  OAI21_X1 U24245 ( .B1(n15782), .B2(n21256), .A(n21230), .ZN(P1_U2922) );
  AOI22_X1 U24246 ( .A1(n21254), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n21231), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n21232) );
  OAI21_X1 U24247 ( .B1(n15784), .B2(n21256), .A(n21232), .ZN(P1_U2923) );
  AOI22_X1 U24248 ( .A1(n21254), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n21231), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n21233) );
  OAI21_X1 U24249 ( .B1(n15787), .B2(n21256), .A(n21233), .ZN(P1_U2924) );
  AOI22_X1 U24250 ( .A1(P1_EAX_REG_11__SCAN_IN), .A2(n21235), .B1(n21234), 
        .B2(P1_LWORD_REG_11__SCAN_IN), .ZN(n21236) );
  OAI21_X1 U24251 ( .B1(n21856), .B2(n21237), .A(n21236), .ZN(P1_U2925) );
  AOI22_X1 U24252 ( .A1(n21254), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n21231), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n21238) );
  OAI21_X1 U24253 ( .B1(n14891), .B2(n21256), .A(n21238), .ZN(P1_U2926) );
  AOI22_X1 U24254 ( .A1(n21254), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n21231), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n21239) );
  OAI21_X1 U24255 ( .B1(n14848), .B2(n21256), .A(n21239), .ZN(P1_U2927) );
  AOI22_X1 U24256 ( .A1(n21254), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n21231), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n21240) );
  OAI21_X1 U24257 ( .B1(n21241), .B2(n21256), .A(n21240), .ZN(P1_U2928) );
  AOI22_X1 U24258 ( .A1(n21254), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n21231), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n21242) );
  OAI21_X1 U24259 ( .B1(n22079), .B2(n21256), .A(n21242), .ZN(P1_U2929) );
  AOI22_X1 U24260 ( .A1(n21254), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n21231), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n21243) );
  OAI21_X1 U24261 ( .B1(n21244), .B2(n21256), .A(n21243), .ZN(P1_U2930) );
  AOI22_X1 U24262 ( .A1(n21254), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n21231), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n21245) );
  OAI21_X1 U24263 ( .B1(n21246), .B2(n21256), .A(n21245), .ZN(P1_U2931) );
  AOI22_X1 U24264 ( .A1(n21254), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n21231), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n21247) );
  OAI21_X1 U24265 ( .B1(n21248), .B2(n21256), .A(n21247), .ZN(P1_U2932) );
  AOI22_X1 U24266 ( .A1(n21254), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n21231), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n21249) );
  OAI21_X1 U24267 ( .B1(n14598), .B2(n21256), .A(n21249), .ZN(P1_U2933) );
  INV_X1 U24268 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n21251) );
  AOI22_X1 U24269 ( .A1(n21254), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n21231), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n21250) );
  OAI21_X1 U24270 ( .B1(n21251), .B2(n21256), .A(n21250), .ZN(P1_U2934) );
  AOI22_X1 U24271 ( .A1(n21254), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n21231), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n21252) );
  OAI21_X1 U24272 ( .B1(n21253), .B2(n21256), .A(n21252), .ZN(P1_U2935) );
  AOI22_X1 U24273 ( .A1(n21254), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n21231), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n21255) );
  OAI21_X1 U24274 ( .B1(n21257), .B2(n21256), .A(n21255), .ZN(P1_U2936) );
  AOI22_X1 U24275 ( .A1(n21275), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n21270), .ZN(n21261) );
  INV_X1 U24276 ( .A(n21258), .ZN(n21259) );
  NAND2_X1 U24277 ( .A1(n21260), .A2(n21259), .ZN(n21276) );
  NAND2_X1 U24278 ( .A1(n21261), .A2(n21276), .ZN(P1_U2951) );
  AOI22_X1 U24279 ( .A1(n9699), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n21270), .ZN(n21263) );
  NAND2_X1 U24280 ( .A1(n21263), .A2(n21262), .ZN(P1_U2961) );
  AOI22_X1 U24281 ( .A1(n9699), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n21270), .ZN(n21265) );
  NAND2_X1 U24282 ( .A1(n21265), .A2(n21264), .ZN(P1_U2962) );
  AOI22_X1 U24283 ( .A1(n9699), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n21270), .ZN(n21267) );
  NAND2_X1 U24284 ( .A1(n21267), .A2(n21266), .ZN(P1_U2963) );
  AOI22_X1 U24285 ( .A1(n9699), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n21270), .ZN(n21269) );
  NAND2_X1 U24286 ( .A1(n21269), .A2(n21268), .ZN(P1_U2964) );
  AOI22_X1 U24287 ( .A1(n9699), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n21270), .ZN(n21273) );
  NAND2_X1 U24288 ( .A1(n21273), .A2(n21272), .ZN(P1_U2965) );
  AOI22_X1 U24289 ( .A1(n21275), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n21274), .ZN(n21277) );
  NAND2_X1 U24290 ( .A1(n21277), .A2(n21276), .ZN(P1_U2966) );
  OAI21_X1 U24291 ( .B1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n21278), .ZN(n21289) );
  NOR2_X1 U24292 ( .A1(n21280), .A2(n21279), .ZN(n21301) );
  NAND2_X1 U24293 ( .A1(n21282), .A2(n21281), .ZN(n21284) );
  OAI211_X1 U24294 ( .C1(n14509), .C2(n21301), .A(n21284), .B(n21283), .ZN(
        n21285) );
  AOI21_X1 U24295 ( .B1(n21287), .B2(n21286), .A(n21285), .ZN(n21288) );
  OAI21_X1 U24296 ( .B1(n21290), .B2(n21289), .A(n21288), .ZN(P1_U3027) );
  INV_X1 U24297 ( .A(n21290), .ZN(n21298) );
  OAI22_X1 U24298 ( .A1(n21293), .A2(n21292), .B1(n21755), .B2(n21291), .ZN(
        n21297) );
  NOR2_X1 U24299 ( .A1(n21295), .A2(n21294), .ZN(n21296) );
  AOI211_X1 U24300 ( .C1(n21298), .C2(n21300), .A(n21297), .B(n21296), .ZN(
        n21299) );
  OAI21_X1 U24301 ( .B1(n21301), .B2(n21300), .A(n21299), .ZN(P1_U3028) );
  NOR2_X1 U24302 ( .A1(n21303), .A2(n21302), .ZN(P1_U3032) );
  NAND2_X1 U24303 ( .A1(n11533), .A2(n21306), .ZN(n21370) );
  OR2_X1 U24304 ( .A1(n21453), .A2(n21370), .ZN(n21337) );
  OAI22_X1 U24305 ( .A1(n21731), .A2(n21643), .B1(n21337), .B2(n21639), .ZN(
        n21307) );
  INV_X1 U24306 ( .A(n21307), .ZN(n21318) );
  OAI21_X1 U24307 ( .B1(n21365), .B2(n21717), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21308) );
  NAND2_X1 U24308 ( .A1(n21308), .A2(n21679), .ZN(n21316) );
  OR2_X1 U24309 ( .A1(n21310), .A2(n21309), .ZN(n21414) );
  NOR2_X1 U24310 ( .A1(n21414), .A2(n21564), .ZN(n21314) );
  OR2_X1 U24311 ( .A1(n21312), .A2(n21311), .ZN(n21450) );
  AOI22_X1 U24312 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21450), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n21337), .ZN(n21313) );
  INV_X1 U24313 ( .A(n21314), .ZN(n21315) );
  AOI22_X1 U24314 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n21340), .B1(
        n21671), .B2(n21339), .ZN(n21317) );
  OAI211_X1 U24315 ( .C1(n21683), .C2(n21362), .A(n21318), .B(n21317), .ZN(
        P1_U3033) );
  OAI22_X1 U24316 ( .A1(n21731), .A2(n21689), .B1(n21337), .B2(n21576), .ZN(
        n21319) );
  INV_X1 U24317 ( .A(n21319), .ZN(n21321) );
  AOI22_X1 U24318 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n21340), .B1(
        n21685), .B2(n21339), .ZN(n21320) );
  OAI211_X1 U24319 ( .C1(n21577), .C2(n21362), .A(n21321), .B(n21320), .ZN(
        P1_U3034) );
  OAI22_X1 U24320 ( .A1(n21731), .A2(n21618), .B1(n21337), .B2(n21581), .ZN(
        n21322) );
  INV_X1 U24321 ( .A(n21322), .ZN(n21324) );
  AOI22_X1 U24322 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n21340), .B1(
        n21691), .B2(n21339), .ZN(n21323) );
  OAI211_X1 U24323 ( .C1(n21695), .C2(n21362), .A(n21324), .B(n21323), .ZN(
        P1_U3035) );
  OAI22_X1 U24324 ( .A1(n21731), .A2(n21586), .B1(n21337), .B2(n21585), .ZN(
        n21325) );
  INV_X1 U24325 ( .A(n21325), .ZN(n21327) );
  AOI22_X1 U24326 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n21340), .B1(
        n21697), .B2(n21339), .ZN(n21326) );
  OAI211_X1 U24327 ( .C1(n21701), .C2(n21362), .A(n21327), .B(n21326), .ZN(
        P1_U3036) );
  OAI22_X1 U24328 ( .A1(n21731), .A2(n21707), .B1(n21337), .B2(n21644), .ZN(
        n21328) );
  INV_X1 U24329 ( .A(n21328), .ZN(n21330) );
  AOI22_X1 U24330 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n21340), .B1(
        n21703), .B2(n21339), .ZN(n21329) );
  OAI211_X1 U24331 ( .C1(n21646), .C2(n21362), .A(n21330), .B(n21329), .ZN(
        P1_U3037) );
  OAI22_X1 U24332 ( .A1(n21731), .A2(n21713), .B1(n21337), .B2(n21593), .ZN(
        n21331) );
  INV_X1 U24333 ( .A(n21331), .ZN(n21333) );
  AOI22_X1 U24334 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n21340), .B1(
        n21709), .B2(n21339), .ZN(n21332) );
  OAI211_X1 U24335 ( .C1(n21597), .C2(n21362), .A(n21333), .B(n21332), .ZN(
        P1_U3038) );
  OAI22_X1 U24336 ( .A1(n21731), .A2(n21721), .B1(n21337), .B2(n21598), .ZN(
        n21334) );
  INV_X1 U24337 ( .A(n21334), .ZN(n21336) );
  AOI22_X1 U24338 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n21340), .B1(
        n21715), .B2(n21339), .ZN(n21335) );
  OAI211_X1 U24339 ( .C1(n21631), .C2(n21362), .A(n21336), .B(n21335), .ZN(
        P1_U3039) );
  OAI22_X1 U24340 ( .A1(n21731), .A2(n21610), .B1(n21337), .B2(n21602), .ZN(
        n21338) );
  INV_X1 U24341 ( .A(n21338), .ZN(n21342) );
  AOI22_X1 U24342 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n21340), .B1(
        n21724), .B2(n21339), .ZN(n21341) );
  OAI211_X1 U24343 ( .C1(n21732), .C2(n21362), .A(n21342), .B(n21341), .ZN(
        P1_U3040) );
  INV_X1 U24344 ( .A(n21414), .ZN(n21343) );
  INV_X1 U24345 ( .A(n16373), .ZN(n21524) );
  NOR2_X1 U24346 ( .A1(n21370), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n21347) );
  INV_X1 U24347 ( .A(n21347), .ZN(n21344) );
  NOR2_X1 U24348 ( .A1(n21561), .A2(n21344), .ZN(n21363) );
  AOI21_X1 U24349 ( .B1(n21343), .B2(n21524), .A(n21363), .ZN(n21345) );
  OAI22_X1 U24350 ( .A1(n21345), .A2(n21667), .B1(n21344), .B2(n10952), .ZN(
        n21364) );
  AOI22_X1 U24351 ( .A1(n21364), .A2(n21671), .B1(n21670), .B2(n21363), .ZN(
        n21349) );
  OAI211_X1 U24352 ( .C1(n21413), .C2(n21528), .A(n21679), .B(n21345), .ZN(
        n21346) );
  OAI211_X1 U24353 ( .C1(n21679), .C2(n21347), .A(n21677), .B(n21346), .ZN(
        n21366) );
  AOI22_X1 U24354 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n21366), .B1(
        n21372), .B2(n21535), .ZN(n21348) );
  OAI211_X1 U24355 ( .C1(n21643), .C2(n21362), .A(n21349), .B(n21348), .ZN(
        P1_U3041) );
  AOI22_X1 U24356 ( .A1(n21364), .A2(n21685), .B1(n21684), .B2(n21363), .ZN(
        n21351) );
  AOI22_X1 U24357 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n21366), .B1(
        n21372), .B2(n21686), .ZN(n21350) );
  OAI211_X1 U24358 ( .C1(n21689), .C2(n21362), .A(n21351), .B(n21350), .ZN(
        P1_U3042) );
  AOI22_X1 U24359 ( .A1(n21364), .A2(n21691), .B1(n21690), .B2(n21363), .ZN(
        n21353) );
  AOI22_X1 U24360 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n21366), .B1(
        n21372), .B2(n21615), .ZN(n21352) );
  OAI211_X1 U24361 ( .C1(n21618), .C2(n21362), .A(n21353), .B(n21352), .ZN(
        P1_U3043) );
  AOI22_X1 U24362 ( .A1(n21364), .A2(n21697), .B1(n21696), .B2(n21363), .ZN(
        n21355) );
  AOI22_X1 U24363 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n21366), .B1(
        n21365), .B2(n21698), .ZN(n21354) );
  OAI211_X1 U24364 ( .C1(n21701), .C2(n21404), .A(n21355), .B(n21354), .ZN(
        P1_U3044) );
  AOI22_X1 U24365 ( .A1(n21364), .A2(n21703), .B1(n21702), .B2(n21363), .ZN(
        n21357) );
  AOI22_X1 U24366 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n21366), .B1(
        n21372), .B2(n21704), .ZN(n21356) );
  OAI211_X1 U24367 ( .C1(n21707), .C2(n21362), .A(n21357), .B(n21356), .ZN(
        P1_U3045) );
  AOI22_X1 U24368 ( .A1(n21364), .A2(n21709), .B1(n21708), .B2(n21363), .ZN(
        n21359) );
  AOI22_X1 U24369 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n21366), .B1(
        n21365), .B2(n21546), .ZN(n21358) );
  OAI211_X1 U24370 ( .C1(n21597), .C2(n21404), .A(n21359), .B(n21358), .ZN(
        P1_U3046) );
  AOI22_X1 U24371 ( .A1(n21364), .A2(n21715), .B1(n21714), .B2(n21363), .ZN(
        n21361) );
  AOI22_X1 U24372 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n21366), .B1(
        n21372), .B2(n21716), .ZN(n21360) );
  OAI211_X1 U24373 ( .C1(n21721), .C2(n21362), .A(n21361), .B(n21360), .ZN(
        P1_U3047) );
  AOI22_X1 U24374 ( .A1(n21364), .A2(n21724), .B1(n21723), .B2(n21363), .ZN(
        n21368) );
  AOI22_X1 U24375 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n21366), .B1(
        n21365), .B2(n21726), .ZN(n21367) );
  OAI211_X1 U24376 ( .C1(n21732), .C2(n21404), .A(n21368), .B(n21367), .ZN(
        P1_U3048) );
  INV_X1 U24377 ( .A(n21370), .ZN(n21411) );
  NAND2_X1 U24378 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21411), .ZN(
        n21419) );
  OR2_X1 U24379 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21419), .ZN(
        n21403) );
  OAI22_X1 U24380 ( .A1(n21443), .A2(n21683), .B1(n21639), .B2(n21403), .ZN(
        n21371) );
  INV_X1 U24381 ( .A(n21371), .ZN(n21384) );
  NOR2_X1 U24382 ( .A1(n21414), .A2(n14754), .ZN(n21378) );
  INV_X1 U24383 ( .A(n21443), .ZN(n21373) );
  OAI21_X1 U24384 ( .B1(n21373), .B2(n21372), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21374) );
  NAND2_X1 U24385 ( .A1(n21374), .A2(n21679), .ZN(n21382) );
  AOI211_X1 U24386 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n21403), .A(n21376), 
        .B(n21375), .ZN(n21377) );
  INV_X1 U24387 ( .A(n21378), .ZN(n21381) );
  INV_X1 U24388 ( .A(n21379), .ZN(n21380) );
  AOI22_X1 U24389 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n21407), .B1(
        n21671), .B2(n21406), .ZN(n21383) );
  OAI211_X1 U24390 ( .C1(n21643), .C2(n21404), .A(n21384), .B(n21383), .ZN(
        P1_U3049) );
  OAI22_X1 U24391 ( .A1(n21443), .A2(n21577), .B1(n21576), .B2(n21403), .ZN(
        n21385) );
  INV_X1 U24392 ( .A(n21385), .ZN(n21387) );
  AOI22_X1 U24393 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n21407), .B1(
        n21685), .B2(n21406), .ZN(n21386) );
  OAI211_X1 U24394 ( .C1(n21689), .C2(n21404), .A(n21387), .B(n21386), .ZN(
        P1_U3050) );
  OAI22_X1 U24395 ( .A1(n21443), .A2(n21695), .B1(n21581), .B2(n21403), .ZN(
        n21388) );
  INV_X1 U24396 ( .A(n21388), .ZN(n21390) );
  AOI22_X1 U24397 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n21407), .B1(
        n21691), .B2(n21406), .ZN(n21389) );
  OAI211_X1 U24398 ( .C1(n21618), .C2(n21404), .A(n21390), .B(n21389), .ZN(
        P1_U3051) );
  OAI22_X1 U24399 ( .A1(n21404), .A2(n21586), .B1(n21585), .B2(n21403), .ZN(
        n21391) );
  INV_X1 U24400 ( .A(n21391), .ZN(n21393) );
  AOI22_X1 U24401 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n21407), .B1(
        n21697), .B2(n21406), .ZN(n21392) );
  OAI211_X1 U24402 ( .C1(n21701), .C2(n21443), .A(n21393), .B(n21392), .ZN(
        P1_U3052) );
  OAI22_X1 U24403 ( .A1(n21404), .A2(n21707), .B1(n21644), .B2(n21403), .ZN(
        n21394) );
  INV_X1 U24404 ( .A(n21394), .ZN(n21396) );
  AOI22_X1 U24405 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n21407), .B1(
        n21703), .B2(n21406), .ZN(n21395) );
  OAI211_X1 U24406 ( .C1(n21646), .C2(n21443), .A(n21396), .B(n21395), .ZN(
        P1_U3053) );
  OAI22_X1 U24407 ( .A1(n21443), .A2(n21597), .B1(n21593), .B2(n21403), .ZN(
        n21397) );
  INV_X1 U24408 ( .A(n21397), .ZN(n21399) );
  AOI22_X1 U24409 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n21407), .B1(
        n21709), .B2(n21406), .ZN(n21398) );
  OAI211_X1 U24410 ( .C1(n21713), .C2(n21404), .A(n21399), .B(n21398), .ZN(
        P1_U3054) );
  OAI22_X1 U24411 ( .A1(n21404), .A2(n21721), .B1(n21598), .B2(n21403), .ZN(
        n21400) );
  INV_X1 U24412 ( .A(n21400), .ZN(n21402) );
  AOI22_X1 U24413 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n21407), .B1(
        n21715), .B2(n21406), .ZN(n21401) );
  OAI211_X1 U24414 ( .C1(n21631), .C2(n21443), .A(n21402), .B(n21401), .ZN(
        P1_U3055) );
  OAI22_X1 U24415 ( .A1(n21404), .A2(n21610), .B1(n21602), .B2(n21403), .ZN(
        n21405) );
  INV_X1 U24416 ( .A(n21405), .ZN(n21409) );
  AOI22_X1 U24417 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n21407), .B1(
        n21724), .B2(n21406), .ZN(n21408) );
  OAI211_X1 U24418 ( .C1(n21732), .C2(n21443), .A(n21409), .B(n21408), .ZN(
        P1_U3056) );
  NAND2_X1 U24419 ( .A1(n21661), .A2(n21411), .ZN(n21442) );
  OAI22_X1 U24420 ( .A1(n21471), .A2(n21683), .B1(n21442), .B2(n21639), .ZN(
        n21412) );
  INV_X1 U24421 ( .A(n21412), .ZN(n21423) );
  AOI21_X1 U24422 ( .B1(n21413), .B2(n21679), .A(n21672), .ZN(n21421) );
  OR2_X1 U24423 ( .A1(n21414), .A2(n21659), .ZN(n21415) );
  INV_X1 U24424 ( .A(n21420), .ZN(n21418) );
  AOI21_X1 U24425 ( .B1(n21667), .B2(n21419), .A(n21416), .ZN(n21417) );
  OAI22_X1 U24426 ( .A1(n21421), .A2(n21420), .B1(n10952), .B2(n21419), .ZN(
        n21445) );
  AOI22_X1 U24427 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n21446), .B1(
        n21671), .B2(n21445), .ZN(n21422) );
  OAI211_X1 U24428 ( .C1(n21643), .C2(n21443), .A(n21423), .B(n21422), .ZN(
        P1_U3057) );
  OAI22_X1 U24429 ( .A1(n21471), .A2(n21577), .B1(n21442), .B2(n21576), .ZN(
        n21424) );
  INV_X1 U24430 ( .A(n21424), .ZN(n21426) );
  AOI22_X1 U24431 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n21446), .B1(
        n21685), .B2(n21445), .ZN(n21425) );
  OAI211_X1 U24432 ( .C1(n21689), .C2(n21443), .A(n21426), .B(n21425), .ZN(
        P1_U3058) );
  OAI22_X1 U24433 ( .A1(n21443), .A2(n21618), .B1(n21581), .B2(n21442), .ZN(
        n21427) );
  INV_X1 U24434 ( .A(n21427), .ZN(n21429) );
  AOI22_X1 U24435 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n21446), .B1(
        n21691), .B2(n21445), .ZN(n21428) );
  OAI211_X1 U24436 ( .C1(n21695), .C2(n21471), .A(n21429), .B(n21428), .ZN(
        P1_U3059) );
  OAI22_X1 U24437 ( .A1(n21443), .A2(n21586), .B1(n21585), .B2(n21442), .ZN(
        n21430) );
  INV_X1 U24438 ( .A(n21430), .ZN(n21432) );
  AOI22_X1 U24439 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n21446), .B1(
        n21697), .B2(n21445), .ZN(n21431) );
  OAI211_X1 U24440 ( .C1(n21701), .C2(n21471), .A(n21432), .B(n21431), .ZN(
        P1_U3060) );
  OAI22_X1 U24441 ( .A1(n21443), .A2(n21707), .B1(n21644), .B2(n21442), .ZN(
        n21433) );
  INV_X1 U24442 ( .A(n21433), .ZN(n21435) );
  AOI22_X1 U24443 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n21446), .B1(
        n21703), .B2(n21445), .ZN(n21434) );
  OAI211_X1 U24444 ( .C1(n21646), .C2(n21471), .A(n21435), .B(n21434), .ZN(
        P1_U3061) );
  OAI22_X1 U24445 ( .A1(n21471), .A2(n21597), .B1(n21442), .B2(n21593), .ZN(
        n21436) );
  INV_X1 U24446 ( .A(n21436), .ZN(n21438) );
  AOI22_X1 U24447 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n21446), .B1(
        n21709), .B2(n21445), .ZN(n21437) );
  OAI211_X1 U24448 ( .C1(n21713), .C2(n21443), .A(n21438), .B(n21437), .ZN(
        P1_U3062) );
  OAI22_X1 U24449 ( .A1(n21443), .A2(n21721), .B1(n21598), .B2(n21442), .ZN(
        n21439) );
  INV_X1 U24450 ( .A(n21439), .ZN(n21441) );
  AOI22_X1 U24451 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n21446), .B1(
        n21715), .B2(n21445), .ZN(n21440) );
  OAI211_X1 U24452 ( .C1(n21631), .C2(n21471), .A(n21441), .B(n21440), .ZN(
        P1_U3063) );
  OAI22_X1 U24453 ( .A1(n21443), .A2(n21610), .B1(n21602), .B2(n21442), .ZN(
        n21444) );
  INV_X1 U24454 ( .A(n21444), .ZN(n21448) );
  AOI22_X1 U24455 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n21446), .B1(
        n21724), .B2(n21445), .ZN(n21447) );
  OAI211_X1 U24456 ( .C1(n21732), .C2(n21471), .A(n21448), .B(n21447), .ZN(
        P1_U3064) );
  INV_X1 U24457 ( .A(n21449), .ZN(n21452) );
  OAI22_X1 U24458 ( .A1(n21452), .A2(n21479), .B1(n21451), .B2(n21450), .ZN(
        n21474) );
  AOI22_X1 U24459 ( .A1(n21474), .A2(n21671), .B1(n21670), .B2(n10670), .ZN(
        n21460) );
  OAI21_X1 U24460 ( .B1(n21475), .B2(n21506), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21456) );
  OAI21_X1 U24461 ( .B1(n21564), .B2(n21479), .A(n21456), .ZN(n21458) );
  AOI22_X1 U24462 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n21476), .B1(
        n21506), .B2(n21535), .ZN(n21459) );
  OAI211_X1 U24463 ( .C1(n21643), .C2(n21471), .A(n21460), .B(n21459), .ZN(
        P1_U3065) );
  AOI22_X1 U24464 ( .A1(n21474), .A2(n21685), .B1(n21684), .B2(n10670), .ZN(
        n21462) );
  AOI22_X1 U24465 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n21476), .B1(
        n21506), .B2(n21686), .ZN(n21461) );
  OAI211_X1 U24466 ( .C1(n21689), .C2(n21471), .A(n21462), .B(n21461), .ZN(
        P1_U3066) );
  AOI22_X1 U24467 ( .A1(n21474), .A2(n21691), .B1(n21690), .B2(n10670), .ZN(
        n21464) );
  AOI22_X1 U24468 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n21476), .B1(
        n21506), .B2(n21615), .ZN(n21463) );
  OAI211_X1 U24469 ( .C1(n21618), .C2(n21471), .A(n21464), .B(n21463), .ZN(
        P1_U3067) );
  AOI22_X1 U24470 ( .A1(n21474), .A2(n21697), .B1(n21696), .B2(n10670), .ZN(
        n21466) );
  AOI22_X1 U24471 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n21476), .B1(
        n21475), .B2(n21698), .ZN(n21465) );
  OAI211_X1 U24472 ( .C1(n21701), .C2(n21501), .A(n21466), .B(n21465), .ZN(
        P1_U3068) );
  AOI22_X1 U24473 ( .A1(n21474), .A2(n21703), .B1(n21702), .B2(n10670), .ZN(
        n21468) );
  AOI22_X1 U24474 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n21476), .B1(
        n21475), .B2(n21621), .ZN(n21467) );
  OAI211_X1 U24475 ( .C1(n21646), .C2(n21501), .A(n21468), .B(n21467), .ZN(
        P1_U3069) );
  AOI22_X1 U24476 ( .A1(n21474), .A2(n21709), .B1(n21708), .B2(n10670), .ZN(
        n21470) );
  AOI22_X1 U24477 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n21476), .B1(
        n21506), .B2(n21710), .ZN(n21469) );
  OAI211_X1 U24478 ( .C1(n21713), .C2(n21471), .A(n21470), .B(n21469), .ZN(
        P1_U3070) );
  AOI22_X1 U24479 ( .A1(n21474), .A2(n21715), .B1(n21714), .B2(n10670), .ZN(
        n21473) );
  AOI22_X1 U24480 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n21476), .B1(
        n21475), .B2(n21628), .ZN(n21472) );
  OAI211_X1 U24481 ( .C1(n21631), .C2(n21501), .A(n21473), .B(n21472), .ZN(
        P1_U3071) );
  AOI22_X1 U24482 ( .A1(n21474), .A2(n21724), .B1(n21723), .B2(n10670), .ZN(
        n21478) );
  AOI22_X1 U24483 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n21476), .B1(
        n21475), .B2(n21726), .ZN(n21477) );
  OAI211_X1 U24484 ( .C1(n21732), .C2(n21501), .A(n21478), .B(n21477), .ZN(
        P1_U3072) );
  INV_X1 U24485 ( .A(n21479), .ZN(n21481) );
  NOR2_X1 U24486 ( .A1(n21480), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n21487) );
  INV_X1 U24487 ( .A(n21487), .ZN(n21482) );
  NOR2_X1 U24488 ( .A1(n21561), .A2(n21482), .ZN(n21504) );
  AOI21_X1 U24489 ( .B1(n21481), .B2(n21524), .A(n21504), .ZN(n21483) );
  OAI22_X1 U24490 ( .A1(n21483), .A2(n21667), .B1(n21482), .B2(n10952), .ZN(
        n21505) );
  AOI22_X1 U24491 ( .A1(n21505), .A2(n21671), .B1(n21670), .B2(n21504), .ZN(
        n21489) );
  OAI21_X1 U24492 ( .B1(n21485), .B2(n21484), .A(n21483), .ZN(n21486) );
  OAI211_X1 U24493 ( .C1(n21679), .C2(n21487), .A(n21677), .B(n21486), .ZN(
        n21507) );
  AOI22_X1 U24494 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n21507), .B1(
        n21498), .B2(n21535), .ZN(n21488) );
  OAI211_X1 U24495 ( .C1(n21643), .C2(n21501), .A(n21489), .B(n21488), .ZN(
        P1_U3073) );
  AOI22_X1 U24496 ( .A1(n21505), .A2(n21685), .B1(n21684), .B2(n21504), .ZN(
        n21491) );
  AOI22_X1 U24497 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n21507), .B1(
        n21498), .B2(n21686), .ZN(n21490) );
  OAI211_X1 U24498 ( .C1(n21689), .C2(n21501), .A(n21491), .B(n21490), .ZN(
        P1_U3074) );
  AOI22_X1 U24499 ( .A1(n21505), .A2(n21691), .B1(n21690), .B2(n21504), .ZN(
        n21493) );
  AOI22_X1 U24500 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n21507), .B1(
        n21498), .B2(n21615), .ZN(n21492) );
  OAI211_X1 U24501 ( .C1(n21618), .C2(n21501), .A(n21493), .B(n21492), .ZN(
        P1_U3075) );
  AOI22_X1 U24502 ( .A1(n21505), .A2(n21697), .B1(n21696), .B2(n21504), .ZN(
        n21495) );
  AOI22_X1 U24503 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n21507), .B1(
        n21506), .B2(n21698), .ZN(n21494) );
  OAI211_X1 U24504 ( .C1(n21701), .C2(n21510), .A(n21495), .B(n21494), .ZN(
        P1_U3076) );
  AOI22_X1 U24505 ( .A1(n21505), .A2(n21703), .B1(n21702), .B2(n21504), .ZN(
        n21497) );
  AOI22_X1 U24506 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n21507), .B1(
        n21506), .B2(n21621), .ZN(n21496) );
  OAI211_X1 U24507 ( .C1(n21646), .C2(n21510), .A(n21497), .B(n21496), .ZN(
        P1_U3077) );
  AOI22_X1 U24508 ( .A1(n21505), .A2(n21709), .B1(n21708), .B2(n21504), .ZN(
        n21500) );
  AOI22_X1 U24509 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n21507), .B1(
        n21498), .B2(n21710), .ZN(n21499) );
  OAI211_X1 U24510 ( .C1(n21713), .C2(n21501), .A(n21500), .B(n21499), .ZN(
        P1_U3078) );
  AOI22_X1 U24511 ( .A1(n21505), .A2(n21715), .B1(n21714), .B2(n21504), .ZN(
        n21503) );
  AOI22_X1 U24512 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n21507), .B1(
        n21506), .B2(n21628), .ZN(n21502) );
  OAI211_X1 U24513 ( .C1(n21631), .C2(n21510), .A(n21503), .B(n21502), .ZN(
        P1_U3079) );
  AOI22_X1 U24514 ( .A1(n21505), .A2(n21724), .B1(n21723), .B2(n21504), .ZN(
        n21509) );
  AOI22_X1 U24515 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n21507), .B1(
        n21506), .B2(n21726), .ZN(n21508) );
  OAI211_X1 U24516 ( .C1(n21732), .C2(n21510), .A(n21509), .B(n21508), .ZN(
        P1_U3080) );
  INV_X1 U24517 ( .A(n21511), .ZN(n21519) );
  AOI22_X1 U24518 ( .A1(n21519), .A2(n21697), .B1(n21518), .B2(n21696), .ZN(
        n21513) );
  AOI22_X1 U24519 ( .A1(n21521), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n21520), .B2(n21698), .ZN(n21512) );
  OAI211_X1 U24520 ( .C1(n21701), .C2(n21559), .A(n21513), .B(n21512), .ZN(
        P1_U3100) );
  AOI22_X1 U24521 ( .A1(n21519), .A2(n21703), .B1(n21518), .B2(n21702), .ZN(
        n21515) );
  AOI22_X1 U24522 ( .A1(n21521), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n21520), .B2(n21621), .ZN(n21514) );
  OAI211_X1 U24523 ( .C1(n21646), .C2(n21559), .A(n21515), .B(n21514), .ZN(
        P1_U3101) );
  AOI22_X1 U24524 ( .A1(n21519), .A2(n21715), .B1(n21518), .B2(n21714), .ZN(
        n21517) );
  AOI22_X1 U24525 ( .A1(n21521), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n21520), .B2(n21628), .ZN(n21516) );
  OAI211_X1 U24526 ( .C1(n21631), .C2(n21559), .A(n21517), .B(n21516), .ZN(
        P1_U3103) );
  AOI22_X1 U24527 ( .A1(n21519), .A2(n21724), .B1(n21518), .B2(n21723), .ZN(
        n21523) );
  AOI22_X1 U24528 ( .A1(n21521), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n21520), .B2(n21726), .ZN(n21522) );
  OAI211_X1 U24529 ( .C1(n21732), .C2(n21559), .A(n21523), .B(n21522), .ZN(
        P1_U3104) );
  NOR3_X2 U24530 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21561), .A3(
        n21525), .ZN(n21552) );
  AOI21_X1 U24531 ( .B1(n21565), .B2(n21524), .A(n21552), .ZN(n21527) );
  NOR2_X1 U24532 ( .A1(n21525), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n21531) );
  INV_X1 U24533 ( .A(n21531), .ZN(n21526) );
  OAI22_X1 U24534 ( .A1(n21527), .A2(n21667), .B1(n21526), .B2(n10952), .ZN(
        n21553) );
  AOI22_X1 U24535 ( .A1(n21553), .A2(n21671), .B1(n21670), .B2(n21552), .ZN(
        n21537) );
  OAI21_X1 U24536 ( .B1(n21529), .B2(n21528), .A(n21527), .ZN(n21530) );
  OAI221_X1 U24537 ( .B1(n21679), .B2(n21531), .C1(n21667), .C2(n21530), .A(
        n21677), .ZN(n21556) );
  INV_X1 U24538 ( .A(n21532), .ZN(n21533) );
  INV_X1 U24539 ( .A(n21609), .ZN(n21555) );
  AOI22_X1 U24540 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n21556), .B1(
        n21555), .B2(n21535), .ZN(n21536) );
  OAI211_X1 U24541 ( .C1(n21643), .C2(n21559), .A(n21537), .B(n21536), .ZN(
        P1_U3105) );
  AOI22_X1 U24542 ( .A1(n21553), .A2(n21685), .B1(n21684), .B2(n21552), .ZN(
        n21539) );
  AOI22_X1 U24543 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n21556), .B1(
        n21555), .B2(n21686), .ZN(n21538) );
  OAI211_X1 U24544 ( .C1(n21689), .C2(n21559), .A(n21539), .B(n21538), .ZN(
        P1_U3106) );
  AOI22_X1 U24545 ( .A1(n21553), .A2(n21691), .B1(n21690), .B2(n21552), .ZN(
        n21541) );
  INV_X1 U24546 ( .A(n21559), .ZN(n21547) );
  AOI22_X1 U24547 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n21556), .B1(
        n21547), .B2(n21692), .ZN(n21540) );
  OAI211_X1 U24548 ( .C1(n21695), .C2(n21609), .A(n21541), .B(n21540), .ZN(
        P1_U3107) );
  AOI22_X1 U24549 ( .A1(n21553), .A2(n21697), .B1(n21696), .B2(n21552), .ZN(
        n21543) );
  AOI22_X1 U24550 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n21556), .B1(
        n21547), .B2(n21698), .ZN(n21542) );
  OAI211_X1 U24551 ( .C1(n21701), .C2(n21609), .A(n21543), .B(n21542), .ZN(
        P1_U3108) );
  AOI22_X1 U24552 ( .A1(n21553), .A2(n21703), .B1(n21702), .B2(n21552), .ZN(
        n21545) );
  AOI22_X1 U24553 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n21556), .B1(
        n21547), .B2(n21621), .ZN(n21544) );
  OAI211_X1 U24554 ( .C1(n21646), .C2(n21609), .A(n21545), .B(n21544), .ZN(
        P1_U3109) );
  AOI22_X1 U24555 ( .A1(n21553), .A2(n21709), .B1(n21708), .B2(n21552), .ZN(
        n21549) );
  AOI22_X1 U24556 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n21556), .B1(
        n21547), .B2(n21546), .ZN(n21548) );
  OAI211_X1 U24557 ( .C1(n21597), .C2(n21609), .A(n21549), .B(n21548), .ZN(
        P1_U3110) );
  AOI22_X1 U24558 ( .A1(n21553), .A2(n21715), .B1(n21714), .B2(n21552), .ZN(
        n21551) );
  AOI22_X1 U24559 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n21556), .B1(
        n21555), .B2(n21716), .ZN(n21550) );
  OAI211_X1 U24560 ( .C1(n21721), .C2(n21559), .A(n21551), .B(n21550), .ZN(
        P1_U3111) );
  AOI22_X1 U24561 ( .A1(n21553), .A2(n21724), .B1(n21723), .B2(n21552), .ZN(
        n21558) );
  AOI22_X1 U24562 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n21556), .B1(
        n21555), .B2(n21554), .ZN(n21557) );
  OAI211_X1 U24563 ( .C1(n21610), .C2(n21559), .A(n21558), .B(n21557), .ZN(
        P1_U3112) );
  NAND3_X1 U24564 ( .A1(n21561), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(
        n21560), .ZN(n21603) );
  OAI22_X1 U24565 ( .A1(n21627), .A2(n21683), .B1(n21603), .B2(n21639), .ZN(
        n21562) );
  INV_X1 U24566 ( .A(n21562), .ZN(n21575) );
  NAND2_X1 U24567 ( .A1(n21627), .A2(n21609), .ZN(n21563) );
  AOI21_X1 U24568 ( .B1(n21563), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n21667), 
        .ZN(n21569) );
  NAND2_X1 U24569 ( .A1(n21565), .A2(n21564), .ZN(n21572) );
  AOI22_X1 U24570 ( .A1(n21569), .A2(n21572), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n21603), .ZN(n21567) );
  NAND3_X1 U24571 ( .A1(n21568), .A2(n21567), .A3(n21566), .ZN(n21606) );
  INV_X1 U24572 ( .A(n21569), .ZN(n21573) );
  AOI22_X1 U24573 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n21606), .B1(
        n21671), .B2(n21605), .ZN(n21574) );
  OAI211_X1 U24574 ( .C1(n21643), .C2(n21609), .A(n21575), .B(n21574), .ZN(
        P1_U3113) );
  OAI22_X1 U24575 ( .A1(n21627), .A2(n21577), .B1(n21603), .B2(n21576), .ZN(
        n21578) );
  INV_X1 U24576 ( .A(n21578), .ZN(n21580) );
  AOI22_X1 U24577 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n21606), .B1(
        n21685), .B2(n21605), .ZN(n21579) );
  OAI211_X1 U24578 ( .C1(n21689), .C2(n21609), .A(n21580), .B(n21579), .ZN(
        P1_U3114) );
  OAI22_X1 U24579 ( .A1(n21627), .A2(n21695), .B1(n21603), .B2(n21581), .ZN(
        n21582) );
  INV_X1 U24580 ( .A(n21582), .ZN(n21584) );
  AOI22_X1 U24581 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n21606), .B1(
        n21691), .B2(n21605), .ZN(n21583) );
  OAI211_X1 U24582 ( .C1(n21618), .C2(n21609), .A(n21584), .B(n21583), .ZN(
        P1_U3115) );
  OAI22_X1 U24583 ( .A1(n21609), .A2(n21586), .B1(n21603), .B2(n21585), .ZN(
        n21587) );
  INV_X1 U24584 ( .A(n21587), .ZN(n21589) );
  AOI22_X1 U24585 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n21606), .B1(
        n21697), .B2(n21605), .ZN(n21588) );
  OAI211_X1 U24586 ( .C1(n21701), .C2(n21627), .A(n21589), .B(n21588), .ZN(
        P1_U3116) );
  OAI22_X1 U24587 ( .A1(n21609), .A2(n21707), .B1(n21603), .B2(n21644), .ZN(
        n21590) );
  INV_X1 U24588 ( .A(n21590), .ZN(n21592) );
  AOI22_X1 U24589 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n21606), .B1(
        n21703), .B2(n21605), .ZN(n21591) );
  OAI211_X1 U24590 ( .C1(n21646), .C2(n21627), .A(n21592), .B(n21591), .ZN(
        P1_U3117) );
  OAI22_X1 U24591 ( .A1(n21609), .A2(n21713), .B1(n21603), .B2(n21593), .ZN(
        n21594) );
  INV_X1 U24592 ( .A(n21594), .ZN(n21596) );
  AOI22_X1 U24593 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n21606), .B1(
        n21709), .B2(n21605), .ZN(n21595) );
  OAI211_X1 U24594 ( .C1(n21597), .C2(n21627), .A(n21596), .B(n21595), .ZN(
        P1_U3118) );
  OAI22_X1 U24595 ( .A1(n21627), .A2(n21631), .B1(n21603), .B2(n21598), .ZN(
        n21599) );
  INV_X1 U24596 ( .A(n21599), .ZN(n21601) );
  AOI22_X1 U24597 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n21606), .B1(
        n21715), .B2(n21605), .ZN(n21600) );
  OAI211_X1 U24598 ( .C1(n21721), .C2(n21609), .A(n21601), .B(n21600), .ZN(
        P1_U3119) );
  OAI22_X1 U24599 ( .A1(n21627), .A2(n21732), .B1(n21603), .B2(n21602), .ZN(
        n21604) );
  INV_X1 U24600 ( .A(n21604), .ZN(n21608) );
  AOI22_X1 U24601 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n21606), .B1(
        n21724), .B2(n21605), .ZN(n21607) );
  OAI211_X1 U24602 ( .C1(n21610), .C2(n21609), .A(n21608), .B(n21607), .ZN(
        P1_U3120) );
  INV_X1 U24603 ( .A(n21612), .ZN(n21632) );
  AOI22_X1 U24604 ( .A1(n21633), .A2(n21685), .B1(n21684), .B2(n21632), .ZN(
        n21614) );
  AOI22_X1 U24605 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n21635), .B1(
        n21624), .B2(n21686), .ZN(n21613) );
  OAI211_X1 U24606 ( .C1(n21689), .C2(n21627), .A(n21614), .B(n21613), .ZN(
        P1_U3122) );
  AOI22_X1 U24607 ( .A1(n21633), .A2(n21691), .B1(n21690), .B2(n21632), .ZN(
        n21617) );
  AOI22_X1 U24608 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n21635), .B1(
        n21624), .B2(n21615), .ZN(n21616) );
  OAI211_X1 U24609 ( .C1(n21618), .C2(n21627), .A(n21617), .B(n21616), .ZN(
        P1_U3123) );
  AOI22_X1 U24610 ( .A1(n21633), .A2(n21697), .B1(n21696), .B2(n21632), .ZN(
        n21620) );
  INV_X1 U24611 ( .A(n21627), .ZN(n21634) );
  AOI22_X1 U24612 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n21635), .B1(
        n21634), .B2(n21698), .ZN(n21619) );
  OAI211_X1 U24613 ( .C1(n21701), .C2(n21653), .A(n21620), .B(n21619), .ZN(
        P1_U3124) );
  AOI22_X1 U24614 ( .A1(n21633), .A2(n21703), .B1(n21702), .B2(n21632), .ZN(
        n21623) );
  AOI22_X1 U24615 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n21635), .B1(
        n21634), .B2(n21621), .ZN(n21622) );
  OAI211_X1 U24616 ( .C1(n21646), .C2(n21653), .A(n21623), .B(n21622), .ZN(
        P1_U3125) );
  AOI22_X1 U24617 ( .A1(n21633), .A2(n21709), .B1(n21708), .B2(n21632), .ZN(
        n21626) );
  AOI22_X1 U24618 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n21635), .B1(
        n21624), .B2(n21710), .ZN(n21625) );
  OAI211_X1 U24619 ( .C1(n21713), .C2(n21627), .A(n21626), .B(n21625), .ZN(
        P1_U3126) );
  AOI22_X1 U24620 ( .A1(n21633), .A2(n21715), .B1(n21714), .B2(n21632), .ZN(
        n21630) );
  AOI22_X1 U24621 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n21635), .B1(
        n21634), .B2(n21628), .ZN(n21629) );
  OAI211_X1 U24622 ( .C1(n21631), .C2(n21653), .A(n21630), .B(n21629), .ZN(
        P1_U3127) );
  AOI22_X1 U24623 ( .A1(n21633), .A2(n21724), .B1(n21723), .B2(n21632), .ZN(
        n21637) );
  AOI22_X1 U24624 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n21635), .B1(
        n21634), .B2(n21726), .ZN(n21636) );
  OAI211_X1 U24625 ( .C1(n21732), .C2(n21653), .A(n21637), .B(n21636), .ZN(
        P1_U3128) );
  INV_X1 U24626 ( .A(n21638), .ZN(n21645) );
  OAI22_X1 U24627 ( .A1(n21647), .A2(n21683), .B1(n21645), .B2(n21639), .ZN(
        n21640) );
  INV_X1 U24628 ( .A(n21640), .ZN(n21642) );
  AOI22_X1 U24629 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n21650), .B1(
        n21671), .B2(n21649), .ZN(n21641) );
  OAI211_X1 U24630 ( .C1(n21643), .C2(n21653), .A(n21642), .B(n21641), .ZN(
        P1_U3129) );
  OAI22_X1 U24631 ( .A1(n21647), .A2(n21646), .B1(n21645), .B2(n21644), .ZN(
        n21648) );
  INV_X1 U24632 ( .A(n21648), .ZN(n21652) );
  AOI22_X1 U24633 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n21650), .B1(
        n21703), .B2(n21649), .ZN(n21651) );
  OAI211_X1 U24634 ( .C1(n21707), .C2(n21653), .A(n21652), .B(n21651), .ZN(
        P1_U3133) );
  AOI22_X1 U24635 ( .A1(n21655), .A2(n21697), .B1(n21696), .B2(n21654), .ZN(
        n21658) );
  AOI22_X1 U24636 ( .A1(n21656), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10689), .B2(n21698), .ZN(n21657) );
  OAI211_X1 U24637 ( .C1(n21701), .C2(n21720), .A(n21658), .B(n21657), .ZN(
        P1_U3148) );
  OR2_X1 U24638 ( .A1(n21660), .A2(n21659), .ZN(n21663) );
  NAND2_X1 U24639 ( .A1(n21662), .A2(n21661), .ZN(n21669) );
  NAND2_X1 U24640 ( .A1(n21663), .A2(n21669), .ZN(n21674) );
  INV_X1 U24641 ( .A(n21674), .ZN(n21668) );
  NOR2_X1 U24642 ( .A1(n21665), .A2(n21664), .ZN(n21678) );
  INV_X1 U24643 ( .A(n21678), .ZN(n21666) );
  OAI22_X1 U24644 ( .A1(n21668), .A2(n21667), .B1(n21666), .B2(n10952), .ZN(
        n21725) );
  INV_X1 U24645 ( .A(n21669), .ZN(n21722) );
  AOI22_X1 U24646 ( .A1(n21725), .A2(n21671), .B1(n21670), .B2(n21722), .ZN(
        n21682) );
  AOI21_X1 U24647 ( .B1(n21673), .B2(n21679), .A(n21672), .ZN(n21675) );
  OR2_X1 U24648 ( .A1(n21675), .A2(n21674), .ZN(n21676) );
  OAI211_X1 U24649 ( .C1(n21679), .C2(n21678), .A(n21677), .B(n21676), .ZN(
        n21728) );
  AOI22_X1 U24650 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n21728), .B1(
        n21727), .B2(n21680), .ZN(n21681) );
  OAI211_X1 U24651 ( .C1(n21683), .C2(n21731), .A(n21682), .B(n21681), .ZN(
        P1_U3153) );
  AOI22_X1 U24652 ( .A1(n21725), .A2(n21685), .B1(n21684), .B2(n21722), .ZN(
        n21688) );
  AOI22_X1 U24653 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n21728), .B1(
        n21717), .B2(n21686), .ZN(n21687) );
  OAI211_X1 U24654 ( .C1(n21689), .C2(n21720), .A(n21688), .B(n21687), .ZN(
        P1_U3154) );
  AOI22_X1 U24655 ( .A1(n21725), .A2(n21691), .B1(n21690), .B2(n21722), .ZN(
        n21694) );
  AOI22_X1 U24656 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n21728), .B1(
        n21727), .B2(n21692), .ZN(n21693) );
  OAI211_X1 U24657 ( .C1(n21695), .C2(n21731), .A(n21694), .B(n21693), .ZN(
        P1_U3155) );
  AOI22_X1 U24658 ( .A1(n21725), .A2(n21697), .B1(n21696), .B2(n21722), .ZN(
        n21700) );
  AOI22_X1 U24659 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n21728), .B1(
        n21727), .B2(n21698), .ZN(n21699) );
  OAI211_X1 U24660 ( .C1(n21701), .C2(n21731), .A(n21700), .B(n21699), .ZN(
        P1_U3156) );
  AOI22_X1 U24661 ( .A1(n21725), .A2(n21703), .B1(n21702), .B2(n21722), .ZN(
        n21706) );
  AOI22_X1 U24662 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n21728), .B1(
        n21717), .B2(n21704), .ZN(n21705) );
  OAI211_X1 U24663 ( .C1(n21707), .C2(n21720), .A(n21706), .B(n21705), .ZN(
        P1_U3157) );
  AOI22_X1 U24664 ( .A1(n21725), .A2(n21709), .B1(n21708), .B2(n21722), .ZN(
        n21712) );
  AOI22_X1 U24665 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n21728), .B1(
        n21717), .B2(n21710), .ZN(n21711) );
  OAI211_X1 U24666 ( .C1(n21713), .C2(n21720), .A(n21712), .B(n21711), .ZN(
        P1_U3158) );
  AOI22_X1 U24667 ( .A1(n21725), .A2(n21715), .B1(n21714), .B2(n21722), .ZN(
        n21719) );
  AOI22_X1 U24668 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n21728), .B1(
        n21717), .B2(n21716), .ZN(n21718) );
  OAI211_X1 U24669 ( .C1(n21721), .C2(n21720), .A(n21719), .B(n21718), .ZN(
        P1_U3159) );
  AOI22_X1 U24670 ( .A1(n21725), .A2(n21724), .B1(n21723), .B2(n21722), .ZN(
        n21730) );
  AOI22_X1 U24671 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n21728), .B1(
        n21727), .B2(n21726), .ZN(n21729) );
  OAI211_X1 U24672 ( .C1(n21732), .C2(n21731), .A(n21730), .B(n21729), .ZN(
        P1_U3160) );
  NOR2_X1 U24673 ( .A1(n21733), .A2(n15370), .ZN(n21735) );
  OAI21_X1 U24674 ( .B1(n21735), .B2(n10952), .A(n21734), .ZN(P1_U3163) );
  AND2_X1 U24675 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n21736), .ZN(
        P1_U3164) );
  AND2_X1 U24676 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n21736), .ZN(
        P1_U3165) );
  AND2_X1 U24677 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n21736), .ZN(
        P1_U3166) );
  INV_X1 U24678 ( .A(P1_DATAWIDTH_REG_28__SCAN_IN), .ZN(n21921) );
  NOR2_X1 U24679 ( .A1(n21798), .A2(n21921), .ZN(P1_U3167) );
  AND2_X1 U24680 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n21736), .ZN(
        P1_U3168) );
  AND2_X1 U24681 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n21736), .ZN(
        P1_U3169) );
  AND2_X1 U24682 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n21736), .ZN(
        P1_U3170) );
  INV_X1 U24683 ( .A(P1_DATAWIDTH_REG_24__SCAN_IN), .ZN(n22035) );
  NOR2_X1 U24684 ( .A1(n21798), .A2(n22035), .ZN(P1_U3171) );
  AND2_X1 U24685 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n21736), .ZN(
        P1_U3172) );
  AND2_X1 U24686 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n21736), .ZN(
        P1_U3173) );
  AND2_X1 U24687 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n21736), .ZN(
        P1_U3174) );
  AND2_X1 U24688 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n21736), .ZN(
        P1_U3175) );
  AND2_X1 U24689 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n21736), .ZN(
        P1_U3176) );
  AND2_X1 U24690 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n21736), .ZN(
        P1_U3177) );
  AND2_X1 U24691 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n21736), .ZN(
        P1_U3178) );
  AND2_X1 U24692 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n21736), .ZN(
        P1_U3179) );
  AND2_X1 U24693 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n21736), .ZN(
        P1_U3180) );
  AND2_X1 U24694 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n21736), .ZN(
        P1_U3181) );
  AND2_X1 U24695 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n21736), .ZN(
        P1_U3182) );
  AND2_X1 U24696 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n21736), .ZN(
        P1_U3183) );
  AND2_X1 U24697 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n21736), .ZN(
        P1_U3184) );
  AND2_X1 U24698 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n21736), .ZN(
        P1_U3185) );
  AND2_X1 U24699 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n21736), .ZN(P1_U3186) );
  AND2_X1 U24700 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n21736), .ZN(P1_U3187) );
  AND2_X1 U24701 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n21736), .ZN(P1_U3188) );
  AND2_X1 U24702 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n21736), .ZN(P1_U3189) );
  AND2_X1 U24703 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n21736), .ZN(P1_U3190) );
  AND2_X1 U24704 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n21736), .ZN(P1_U3191) );
  AND2_X1 U24705 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n21736), .ZN(P1_U3192) );
  AND2_X1 U24706 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n21736), .ZN(P1_U3193) );
  NAND2_X1 U24707 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21741), .ZN(n21745) );
  INV_X1 U24708 ( .A(n21745), .ZN(n21740) );
  OAI21_X1 U24709 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n21746), .A(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21737) );
  AOI211_X1 U24710 ( .C1(HOLD), .C2(P1_STATE_REG_1__SCAN_IN), .A(n21738), .B(
        n21737), .ZN(n21739) );
  OAI22_X1 U24711 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21740), .B1(n21817), 
        .B2(n21739), .ZN(P1_U3194) );
  INV_X1 U24712 ( .A(n21741), .ZN(n21744) );
  INV_X1 U24713 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21829) );
  AOI21_X1 U24714 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(n21751), .A(n21742), .ZN(n21743) );
  AOI21_X1 U24715 ( .B1(n21744), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .A(n21743), .ZN(n21750) );
  NAND3_X1 U24716 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21822), .A3(n21746), 
        .ZN(n21748) );
  OAI211_X1 U24717 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n21746), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n21745), .ZN(n21747) );
  OAI221_X1 U24718 ( .B1(n21750), .B2(n21749), .C1(n21750), .C2(n21748), .A(
        n21747), .ZN(P1_U3196) );
  NOR2_X1 U24719 ( .A1(n21815), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n21784) );
  CLKBUF_X1 U24720 ( .A(n21784), .Z(n21788) );
  AOI222_X1 U24721 ( .A1(n21788), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n21815), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n21789), .ZN(n21752) );
  INV_X1 U24722 ( .A(n21752), .ZN(P1_U3197) );
  AOI222_X1 U24723 ( .A1(n21789), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n21815), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n21784), .ZN(n21753) );
  INV_X1 U24724 ( .A(n21753), .ZN(P1_U3198) );
  INV_X1 U24725 ( .A(n21789), .ZN(n21780) );
  INV_X1 U24726 ( .A(n21784), .ZN(n21777) );
  OAI222_X1 U24727 ( .A1(n21780), .A2(n21755), .B1(n21754), .B2(n21817), .C1(
        n22126), .C2(n21777), .ZN(P1_U3199) );
  AOI222_X1 U24728 ( .A1(n21788), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n21815), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n21789), .ZN(n21756) );
  INV_X1 U24729 ( .A(n21756), .ZN(P1_U3200) );
  INV_X1 U24730 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n21905) );
  OAI222_X1 U24731 ( .A1(n21780), .A2(n21757), .B1(n21905), .B2(n21817), .C1(
        n21759), .C2(n21777), .ZN(P1_U3201) );
  AOI22_X1 U24732 ( .A1(P1_ADDRESS_REG_5__SCAN_IN), .A2(n21815), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n21784), .ZN(n21758) );
  OAI21_X1 U24733 ( .B1(n21759), .B2(n21780), .A(n21758), .ZN(P1_U3202) );
  AOI22_X1 U24734 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n21815), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n21789), .ZN(n21760) );
  OAI21_X1 U24735 ( .B1(n16006), .B2(n21777), .A(n21760), .ZN(P1_U3203) );
  AOI222_X1 U24736 ( .A1(n21789), .A2(P1_REIP_REG_8__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n21815), .C1(P1_REIP_REG_9__SCAN_IN), 
        .C2(n21784), .ZN(n21761) );
  INV_X1 U24737 ( .A(n21761), .ZN(P1_U3204) );
  AOI222_X1 U24738 ( .A1(n21789), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n21815), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n21788), .ZN(n21762) );
  INV_X1 U24739 ( .A(n21762), .ZN(P1_U3205) );
  INV_X1 U24740 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n21863) );
  INV_X1 U24741 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n21763) );
  OAI222_X1 U24742 ( .A1(n21780), .A2(n15984), .B1(n21863), .B2(n21817), .C1(
        n21763), .C2(n21777), .ZN(P1_U3206) );
  AOI222_X1 U24743 ( .A1(n21789), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n21815), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n21788), .ZN(n21764) );
  INV_X1 U24744 ( .A(n21764), .ZN(P1_U3207) );
  AOI222_X1 U24745 ( .A1(n21784), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n21815), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n21789), .ZN(n21765) );
  INV_X1 U24746 ( .A(n21765), .ZN(P1_U3208) );
  AOI222_X1 U24747 ( .A1(n21784), .A2(P1_REIP_REG_14__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n21815), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n21789), .ZN(n21766) );
  INV_X1 U24748 ( .A(n21766), .ZN(P1_U3209) );
  AOI222_X1 U24749 ( .A1(n21788), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n21815), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n21789), .ZN(n21767) );
  INV_X1 U24750 ( .A(n21767), .ZN(P1_U3210) );
  AOI222_X1 U24751 ( .A1(n21788), .A2(P1_REIP_REG_16__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n21815), .C1(P1_REIP_REG_15__SCAN_IN), 
        .C2(n21789), .ZN(n21768) );
  INV_X1 U24752 ( .A(n21768), .ZN(P1_U3211) );
  AOI222_X1 U24753 ( .A1(n21789), .A2(P1_REIP_REG_16__SCAN_IN), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n21815), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n21784), .ZN(n21769) );
  INV_X1 U24754 ( .A(n21769), .ZN(P1_U3212) );
  INV_X1 U24755 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n21910) );
  OAI222_X1 U24756 ( .A1(n21777), .A2(n21771), .B1(n21910), .B2(n21817), .C1(
        n21770), .C2(n21780), .ZN(P1_U3213) );
  AOI222_X1 U24757 ( .A1(n21789), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n21815), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n21784), .ZN(n21772) );
  INV_X1 U24758 ( .A(n21772), .ZN(P1_U3214) );
  AOI222_X1 U24759 ( .A1(n21789), .A2(P1_REIP_REG_19__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n21815), .C1(P1_REIP_REG_20__SCAN_IN), 
        .C2(n21788), .ZN(n21773) );
  INV_X1 U24760 ( .A(n21773), .ZN(P1_U3215) );
  AOI22_X1 U24761 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(n21815), .B1(
        P1_REIP_REG_21__SCAN_IN), .B2(n21788), .ZN(n21774) );
  OAI21_X1 U24762 ( .B1(n21775), .B2(n21780), .A(n21774), .ZN(P1_U3216) );
  AOI22_X1 U24763 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(n21815), .B1(
        P1_REIP_REG_21__SCAN_IN), .B2(n21789), .ZN(n21776) );
  OAI21_X1 U24764 ( .B1(n21971), .B2(n21777), .A(n21776), .ZN(P1_U3217) );
  INV_X1 U24765 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n21893) );
  OAI222_X1 U24766 ( .A1(n21780), .A2(n21971), .B1(n21893), .B2(n21817), .C1(
        n21779), .C2(n21777), .ZN(P1_U3218) );
  INV_X1 U24767 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n21778) );
  OAI222_X1 U24768 ( .A1(n21780), .A2(n21779), .B1(n21778), .B2(n21817), .C1(
        n22018), .C2(n21777), .ZN(P1_U3219) );
  AOI222_X1 U24769 ( .A1(n21789), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n21815), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n21788), .ZN(n21781) );
  INV_X1 U24770 ( .A(n21781), .ZN(P1_U3220) );
  AOI222_X1 U24771 ( .A1(n21789), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n21815), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n21784), .ZN(n21782) );
  INV_X1 U24772 ( .A(n21782), .ZN(P1_U3221) );
  AOI222_X1 U24773 ( .A1(n21789), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n21815), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n21784), .ZN(n21783) );
  INV_X1 U24774 ( .A(n21783), .ZN(P1_U3222) );
  AOI222_X1 U24775 ( .A1(n21784), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n21815), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n21789), .ZN(n21785) );
  INV_X1 U24776 ( .A(n21785), .ZN(P1_U3223) );
  AOI222_X1 U24777 ( .A1(n21789), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n21815), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n21788), .ZN(n21786) );
  INV_X1 U24778 ( .A(n21786), .ZN(P1_U3224) );
  AOI222_X1 U24779 ( .A1(n21789), .A2(P1_REIP_REG_29__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n21815), .C1(P1_REIP_REG_30__SCAN_IN), 
        .C2(n21788), .ZN(n21787) );
  INV_X1 U24780 ( .A(n21787), .ZN(P1_U3225) );
  AOI222_X1 U24781 ( .A1(n21789), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n21815), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n21788), .ZN(n21790) );
  INV_X1 U24782 ( .A(n21790), .ZN(P1_U3226) );
  OAI22_X1 U24783 ( .A1(n21815), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n21817), .ZN(n21791) );
  INV_X1 U24784 ( .A(n21791), .ZN(P1_U3458) );
  OAI22_X1 U24785 ( .A1(n21815), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n21817), .ZN(n21792) );
  INV_X1 U24786 ( .A(n21792), .ZN(P1_U3459) );
  OAI22_X1 U24787 ( .A1(n21815), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n21817), .ZN(n21793) );
  INV_X1 U24788 ( .A(n21793), .ZN(P1_U3460) );
  OAI22_X1 U24789 ( .A1(n21815), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n21817), .ZN(n21794) );
  INV_X1 U24790 ( .A(n21794), .ZN(P1_U3461) );
  OAI21_X1 U24791 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n21798), .A(n21796), 
        .ZN(n21795) );
  INV_X1 U24792 ( .A(n21795), .ZN(P1_U3464) );
  OAI21_X1 U24793 ( .B1(n21798), .B2(n21797), .A(n21796), .ZN(P1_U3465) );
  INV_X1 U24794 ( .A(n21799), .ZN(n21803) );
  OAI22_X1 U24795 ( .A1(n21803), .A2(n21802), .B1(n21801), .B2(n21800), .ZN(
        n21805) );
  MUX2_X1 U24796 ( .A(n21805), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n21804), .Z(P1_U3469) );
  AOI21_X1 U24797 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n21807) );
  AOI22_X1 U24798 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n21807), .B2(n21806), .ZN(n21809) );
  INV_X1 U24799 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21808) );
  AOI22_X1 U24800 ( .A1(n21810), .A2(n21809), .B1(n21808), .B2(n21813), .ZN(
        P1_U3481) );
  INV_X1 U24801 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21814) );
  NOR2_X1 U24802 ( .A1(n21813), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n21811) );
  AOI22_X1 U24803 ( .A1(n21814), .A2(n21813), .B1(n21812), .B2(n21811), .ZN(
        P1_U3482) );
  AOI22_X1 U24804 ( .A1(n21817), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21816), 
        .B2(n21815), .ZN(P1_U3483) );
  INV_X1 U24805 ( .A(n21818), .ZN(n21819) );
  OAI211_X1 U24806 ( .C1(n21822), .C2(n21821), .A(n21820), .B(n21819), .ZN(
        n21830) );
  NOR2_X1 U24807 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21823), .ZN(n21828) );
  OAI211_X1 U24808 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n21825), .A(n21824), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n21826) );
  NAND2_X1 U24809 ( .A1(n21830), .A2(n21826), .ZN(n21827) );
  OAI22_X1 U24810 ( .A1(n21830), .A2(n21829), .B1(n21828), .B2(n21827), .ZN(
        P1_U3485) );
  MUX2_X1 U24811 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(P1_M_IO_N_REG_SCAN_IN), 
        .S(n21815), .Z(P1_U3486) );
  AOI22_X1 U24812 ( .A1(n21834), .A2(n21833), .B1(n21832), .B2(n21831), .ZN(
        n21839) );
  AOI22_X1 U24813 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n21837), .B1(
        n21836), .B2(n21835), .ZN(n21838) );
  OAI211_X1 U24814 ( .C1(n21841), .C2(n21840), .A(n21839), .B(n21838), .ZN(
        n22149) );
  AOI22_X1 U24815 ( .A1(n21967), .A2(keyinput34), .B1(keyinput57), .B2(n21843), 
        .ZN(n21842) );
  OAI221_X1 U24816 ( .B1(n21967), .B2(keyinput34), .C1(n21843), .C2(keyinput57), .A(n21842), .ZN(n21854) );
  INV_X1 U24817 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n21845) );
  AOI22_X1 U24818 ( .A1(n16396), .A2(keyinput91), .B1(keyinput109), .B2(n21845), .ZN(n21844) );
  OAI221_X1 U24819 ( .B1(n16396), .B2(keyinput91), .C1(n21845), .C2(
        keyinput109), .A(n21844), .ZN(n21853) );
  INV_X1 U24820 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n21847) );
  AOI22_X1 U24821 ( .A1(n21848), .A2(keyinput64), .B1(n21847), .B2(keyinput16), 
        .ZN(n21846) );
  OAI221_X1 U24822 ( .B1(n21848), .B2(keyinput64), .C1(n21847), .C2(keyinput16), .A(n21846), .ZN(n21852) );
  XOR2_X1 U24823 ( .A(n21966), .B(keyinput31), .Z(n21850) );
  XNOR2_X1 U24824 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(keyinput108), 
        .ZN(n21849) );
  NAND2_X1 U24825 ( .A1(n21850), .A2(n21849), .ZN(n21851) );
  NOR4_X1 U24826 ( .A1(n21854), .A2(n21853), .A3(n21852), .A4(n21851), .ZN(
        n22147) );
  NAND2_X1 U24827 ( .A1(n21968), .A2(keyinput66), .ZN(n21855) );
  OAI221_X1 U24828 ( .B1(n21856), .B2(keyinput60), .C1(n21968), .C2(keyinput66), .A(n21855), .ZN(n21868) );
  AOI22_X1 U24829 ( .A1(n21971), .A2(keyinput97), .B1(n21858), .B2(keyinput105), .ZN(n21857) );
  OAI221_X1 U24830 ( .B1(n21971), .B2(keyinput97), .C1(n21858), .C2(
        keyinput105), .A(n21857), .ZN(n21867) );
  AOI22_X1 U24831 ( .A1(n21861), .A2(keyinput70), .B1(keyinput19), .B2(n21860), 
        .ZN(n21859) );
  OAI221_X1 U24832 ( .B1(n21861), .B2(keyinput70), .C1(n21860), .C2(keyinput19), .A(n21859), .ZN(n21866) );
  AOI22_X1 U24833 ( .A1(n21864), .A2(keyinput32), .B1(n21863), .B2(keyinput112), .ZN(n21862) );
  OAI221_X1 U24834 ( .B1(n21864), .B2(keyinput32), .C1(n21863), .C2(
        keyinput112), .A(n21862), .ZN(n21865) );
  NOR4_X1 U24835 ( .A1(n21868), .A2(n21867), .A3(n21866), .A4(n21865), .ZN(
        n22146) );
  INV_X1 U24836 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n21870) );
  AOI22_X1 U24837 ( .A1(n21871), .A2(keyinput116), .B1(n21870), .B2(
        keyinput100), .ZN(n21869) );
  OAI221_X1 U24838 ( .B1(n21871), .B2(keyinput116), .C1(n21870), .C2(
        keyinput100), .A(n21869), .ZN(n21950) );
  AOI22_X1 U24839 ( .A1(n21986), .A2(keyinput65), .B1(n21985), .B2(keyinput8), 
        .ZN(n21872) );
  OAI221_X1 U24840 ( .B1(n21986), .B2(keyinput65), .C1(n21985), .C2(keyinput8), 
        .A(n21872), .ZN(n21949) );
  OAI22_X1 U24841 ( .A1(n12357), .A2(keyinput27), .B1(n21874), .B2(keyinput72), 
        .ZN(n21873) );
  AOI221_X1 U24842 ( .B1(n12357), .B2(keyinput27), .C1(keyinput72), .C2(n21874), .A(n21873), .ZN(n21891) );
  INV_X1 U24843 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n21877) );
  OAI22_X1 U24844 ( .A1(n21877), .A2(keyinput93), .B1(n21876), .B2(keyinput41), 
        .ZN(n21875) );
  AOI221_X1 U24845 ( .B1(n21877), .B2(keyinput93), .C1(keyinput41), .C2(n21876), .A(n21875), .ZN(n21890) );
  AOI22_X1 U24846 ( .A1(n16540), .A2(keyinput3), .B1(n13229), .B2(keyinput28), 
        .ZN(n21878) );
  OAI221_X1 U24847 ( .B1(n16540), .B2(keyinput3), .C1(n13229), .C2(keyinput28), 
        .A(n21878), .ZN(n21888) );
  AOI22_X1 U24848 ( .A1(n14260), .A2(keyinput75), .B1(n21984), .B2(keyinput46), 
        .ZN(n21879) );
  OAI221_X1 U24849 ( .B1(n14260), .B2(keyinput75), .C1(n21984), .C2(keyinput46), .A(n21879), .ZN(n21887) );
  INV_X1 U24850 ( .A(P3_DATAO_REG_0__SCAN_IN), .ZN(n21881) );
  AOI22_X1 U24851 ( .A1(n21882), .A2(keyinput83), .B1(keyinput120), .B2(n21881), .ZN(n21880) );
  OAI221_X1 U24852 ( .B1(n21882), .B2(keyinput83), .C1(n21881), .C2(
        keyinput120), .A(n21880), .ZN(n21886) );
  INV_X1 U24853 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n21884) );
  AOI22_X1 U24854 ( .A1(n21884), .A2(keyinput33), .B1(n16409), .B2(keyinput44), 
        .ZN(n21883) );
  OAI221_X1 U24855 ( .B1(n21884), .B2(keyinput33), .C1(n16409), .C2(keyinput44), .A(n21883), .ZN(n21885) );
  NOR4_X1 U24856 ( .A1(n21888), .A2(n21887), .A3(n21886), .A4(n21885), .ZN(
        n21889) );
  NAND3_X1 U24857 ( .A1(n21891), .A2(n21890), .A3(n21889), .ZN(n21948) );
  AOI22_X1 U24858 ( .A1(n21894), .A2(keyinput111), .B1(keyinput98), .B2(n21893), .ZN(n21892) );
  OAI221_X1 U24859 ( .B1(n21894), .B2(keyinput111), .C1(n21893), .C2(
        keyinput98), .A(n21892), .ZN(n21903) );
  AOI22_X1 U24860 ( .A1(n21989), .A2(keyinput17), .B1(keyinput40), .B2(n14575), 
        .ZN(n21895) );
  OAI221_X1 U24861 ( .B1(n21989), .B2(keyinput17), .C1(n14575), .C2(keyinput40), .A(n21895), .ZN(n21902) );
  AOI22_X1 U24862 ( .A1(n21897), .A2(keyinput6), .B1(n21988), .B2(keyinput115), 
        .ZN(n21896) );
  OAI221_X1 U24863 ( .B1(n21897), .B2(keyinput6), .C1(n21988), .C2(keyinput115), .A(n21896), .ZN(n21901) );
  XOR2_X1 U24864 ( .A(n21987), .B(keyinput95), .Z(n21899) );
  XNOR2_X1 U24865 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B(keyinput5), .ZN(
        n21898) );
  NAND2_X1 U24866 ( .A1(n21899), .A2(n21898), .ZN(n21900) );
  NOR4_X1 U24867 ( .A1(n21903), .A2(n21902), .A3(n21901), .A4(n21900), .ZN(
        n21946) );
  AOI22_X1 U24868 ( .A1(n21906), .A2(keyinput68), .B1(keyinput86), .B2(n21905), 
        .ZN(n21904) );
  OAI221_X1 U24869 ( .B1(n21906), .B2(keyinput68), .C1(n21905), .C2(keyinput86), .A(n21904), .ZN(n21916) );
  AOI22_X1 U24870 ( .A1(n21983), .A2(keyinput48), .B1(keyinput87), .B2(n21908), 
        .ZN(n21907) );
  OAI221_X1 U24871 ( .B1(n21983), .B2(keyinput48), .C1(n21908), .C2(keyinput87), .A(n21907), .ZN(n21915) );
  AOI22_X1 U24872 ( .A1(n21910), .A2(keyinput22), .B1(keyinput59), .B2(n15984), 
        .ZN(n21909) );
  OAI221_X1 U24873 ( .B1(n21910), .B2(keyinput22), .C1(n15984), .C2(keyinput59), .A(n21909), .ZN(n21914) );
  AOI22_X1 U24874 ( .A1(n21981), .A2(keyinput56), .B1(n21912), .B2(keyinput62), 
        .ZN(n21911) );
  OAI221_X1 U24875 ( .B1(n21981), .B2(keyinput56), .C1(n21912), .C2(keyinput62), .A(n21911), .ZN(n21913) );
  NOR4_X1 U24876 ( .A1(n21916), .A2(n21915), .A3(n21914), .A4(n21913), .ZN(
        n21945) );
  AOI22_X1 U24877 ( .A1(n21919), .A2(keyinput127), .B1(keyinput114), .B2(
        n21918), .ZN(n21917) );
  OAI221_X1 U24878 ( .B1(n21919), .B2(keyinput127), .C1(n21918), .C2(
        keyinput114), .A(n21917), .ZN(n21930) );
  AOI22_X1 U24879 ( .A1(n15132), .A2(keyinput121), .B1(keyinput45), .B2(n21921), .ZN(n21920) );
  OAI221_X1 U24880 ( .B1(n15132), .B2(keyinput121), .C1(n21921), .C2(
        keyinput45), .A(n21920), .ZN(n21929) );
  AOI22_X1 U24881 ( .A1(n21923), .A2(keyinput26), .B1(n22005), .B2(keyinput125), .ZN(n21922) );
  OAI221_X1 U24882 ( .B1(n21923), .B2(keyinput26), .C1(n22005), .C2(
        keyinput125), .A(n21922), .ZN(n21928) );
  AOI22_X1 U24883 ( .A1(n21926), .A2(keyinput9), .B1(n21925), .B2(keyinput23), 
        .ZN(n21924) );
  OAI221_X1 U24884 ( .B1(n21926), .B2(keyinput9), .C1(n21925), .C2(keyinput23), 
        .A(n21924), .ZN(n21927) );
  NOR4_X1 U24885 ( .A1(n21930), .A2(n21929), .A3(n21928), .A4(n21927), .ZN(
        n21944) );
  AOI22_X1 U24886 ( .A1(n22004), .A2(keyinput38), .B1(keyinput101), .B2(n22003), .ZN(n21931) );
  OAI221_X1 U24887 ( .B1(n22004), .B2(keyinput38), .C1(n22003), .C2(
        keyinput101), .A(n21931), .ZN(n21942) );
  AOI22_X1 U24888 ( .A1(n21933), .A2(keyinput107), .B1(n11533), .B2(keyinput2), 
        .ZN(n21932) );
  OAI221_X1 U24889 ( .B1(n21933), .B2(keyinput107), .C1(n11533), .C2(keyinput2), .A(n21932), .ZN(n21941) );
  INV_X1 U24890 ( .A(DATAI_19_), .ZN(n21935) );
  AOI22_X1 U24891 ( .A1(n21935), .A2(keyinput58), .B1(n14509), .B2(keyinput113), .ZN(n21934) );
  OAI221_X1 U24892 ( .B1(n21935), .B2(keyinput58), .C1(n14509), .C2(
        keyinput113), .A(n21934), .ZN(n21940) );
  XOR2_X1 U24893 ( .A(n21936), .B(keyinput110), .Z(n21938) );
  XNOR2_X1 U24894 ( .A(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B(keyinput53), .ZN(
        n21937) );
  NAND2_X1 U24895 ( .A1(n21938), .A2(n21937), .ZN(n21939) );
  NOR4_X1 U24896 ( .A1(n21942), .A2(n21941), .A3(n21940), .A4(n21939), .ZN(
        n21943) );
  NAND4_X1 U24897 ( .A1(n21946), .A2(n21945), .A3(n21944), .A4(n21943), .ZN(
        n21947) );
  NOR4_X1 U24898 ( .A1(n21950), .A2(n21949), .A3(n21948), .A4(n21947), .ZN(
        n22145) );
  NOR4_X1 U24899 ( .A1(P2_EBX_REG_5__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_7__5__SCAN_IN), .A3(P3_ADDRESS_REG_15__SCAN_IN), .A4(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n21962) );
  NOR4_X1 U24900 ( .A1(P2_EBX_REG_6__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A3(P2_EBX_REG_15__SCAN_IN), .A4(
        P3_EAX_REG_2__SCAN_IN), .ZN(n21961) );
  NAND4_X1 U24901 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(P3_DATAO_REG_6__SCAN_IN), .A4(
        P3_EAX_REG_20__SCAN_IN), .ZN(n21953) );
  INV_X1 U24902 ( .A(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n21951) );
  NAND2_X1 U24903 ( .A1(n21951), .A2(P1_EAX_REG_7__SCAN_IN), .ZN(n21952) );
  NOR4_X1 U24904 ( .A1(n21953), .A2(n21952), .A3(n22083), .A4(
        P2_EAX_REG_16__SCAN_IN), .ZN(n21960) );
  NAND4_X1 U24905 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(
        P3_BYTEENABLE_REG_0__SCAN_IN), .A3(n22115), .A4(n22118), .ZN(n21958)
         );
  NAND4_X1 U24906 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n22100), .A3(n22099), .A4(
        n22110), .ZN(n21957) );
  NAND4_X1 U24907 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_DATAO_REG_28__SCAN_IN), 
        .A3(P2_DATAWIDTH_REG_25__SCAN_IN), .A4(n22124), .ZN(n21956) );
  INV_X1 U24908 ( .A(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n21954) );
  NAND4_X1 U24909 ( .A1(n21954), .A2(P2_EBX_REG_7__SCAN_IN), .A3(
        P1_INSTQUEUE_REG_5__3__SCAN_IN), .A4(n22130), .ZN(n21955) );
  NOR4_X1 U24910 ( .A1(n21958), .A2(n21957), .A3(n21956), .A4(n21955), .ZN(
        n21959) );
  NAND4_X1 U24911 ( .A1(n21962), .A2(n21961), .A3(n21960), .A4(n21959), .ZN(
        n22015) );
  INV_X1 U24912 ( .A(n13261), .ZN(n21963) );
  NOR4_X1 U24913 ( .A1(n21964), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A3(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A4(n21963), .ZN(n21965) );
  NAND3_X1 U24914 ( .A1(n21965), .A2(P2_DATAWIDTH_REG_11__SCAN_IN), .A3(n22093), .ZN(n21979) );
  NAND4_X1 U24915 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n21967), .A3(n16396), 
        .A4(n21966), .ZN(n21978) );
  NAND4_X1 U24916 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_12__SCAN_IN), .A4(
        n21968), .ZN(n21977) );
  INV_X1 U24917 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n22114) );
  NOR4_X1 U24918 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(
        P2_EBX_REG_1__SCAN_IN), .A3(n12440), .A4(n22114), .ZN(n21975) );
  NOR4_X1 U24919 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_14__0__SCAN_IN), .A3(P2_INSTQUEUE_REG_8__0__SCAN_IN), 
        .A4(n22046), .ZN(n21970) );
  NOR4_X1 U24920 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_4__6__SCAN_IN), .A3(P2_INSTQUEUE_REG_5__6__SCAN_IN), 
        .A4(n12452), .ZN(n21969) );
  NAND3_X1 U24921 ( .A1(n21971), .A2(n21970), .A3(n21969), .ZN(n21973) );
  NOR4_X1 U24922 ( .A1(n21973), .A2(n21972), .A3(P2_EBX_REG_8__SCAN_IN), .A4(
        BUF2_REG_7__SCAN_IN), .ZN(n21974) );
  NAND2_X1 U24923 ( .A1(n21975), .A2(n21974), .ZN(n21976) );
  NOR4_X1 U24924 ( .A1(n21979), .A2(n21978), .A3(n21977), .A4(n21976), .ZN(
        n22013) );
  NOR4_X1 U24925 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(P3_ADDRESS_REG_14__SCAN_IN), .A3(P1_DATAO_REG_30__SCAN_IN), .A4(P3_DATAO_REG_0__SCAN_IN), .ZN(n21980) );
  NAND3_X1 U24926 ( .A1(P2_UWORD_REG_1__SCAN_IN), .A2(n21980), .A3(n16540), 
        .ZN(n21997) );
  NAND4_X1 U24927 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(n15984), .A4(n21981), .ZN(
        n21982) );
  NOR3_X1 U24928 ( .A1(P3_ADDRESS_REG_3__SCAN_IN), .A2(n21983), .A3(n21982), 
        .ZN(n21995) );
  NAND4_X1 U24929 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_10__SCAN_IN), .A3(n14260), .A4(n21984), .ZN(n21993)
         );
  NAND4_X1 U24930 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A3(n21986), .A4(n21985), .ZN(
        n21992) );
  NAND4_X1 U24931 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_12__5__SCAN_IN), .A3(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A4(n21987), .ZN(n21991) );
  NAND4_X1 U24932 ( .A1(DATAI_5_), .A2(P3_EBX_REG_21__SCAN_IN), .A3(n21989), 
        .A4(n21988), .ZN(n21990) );
  NOR4_X1 U24933 ( .A1(n21993), .A2(n21992), .A3(n21991), .A4(n21990), .ZN(
        n21994) );
  NAND4_X1 U24934 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_ADDRESS_REG_4__SCAN_IN), .A3(n21995), .A4(n21994), .ZN(n21996) );
  NOR4_X1 U24935 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(
        P1_CODEFETCH_REG_SCAN_IN), .A3(n21997), .A4(n21996), .ZN(n22012) );
  NAND4_X1 U24936 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_EBX_REG_29__SCAN_IN), .A3(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A4(
        n22035), .ZN(n22002) );
  INV_X1 U24937 ( .A(P3_DATAO_REG_29__SCAN_IN), .ZN(n22039) );
  NAND4_X1 U24938 ( .A1(n22037), .A2(n22040), .A3(n22039), .A4(
        P3_REIP_REG_30__SCAN_IN), .ZN(n22001) );
  NAND4_X1 U24939 ( .A1(P1_EBX_REG_31__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(P3_DATAWIDTH_REG_25__SCAN_IN), 
        .A4(P1_UWORD_REG_12__SCAN_IN), .ZN(n22000) );
  INV_X1 U24940 ( .A(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n21998) );
  INV_X1 U24941 ( .A(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n22025) );
  NAND4_X1 U24942 ( .A1(n21998), .A2(P3_REIP_REG_24__SCAN_IN), .A3(n22025), 
        .A4(P3_STATE_REG_1__SCAN_IN), .ZN(n21999) );
  NOR4_X1 U24943 ( .A1(n22002), .A2(n22001), .A3(n22000), .A4(n21999), .ZN(
        n22011) );
  NAND4_X1 U24944 ( .A1(DATAI_19_), .A2(P1_DATAWIDTH_REG_28__SCAN_IN), .A3(
        n14509), .A4(n22003), .ZN(n22009) );
  NAND4_X1 U24945 ( .A1(P2_EAX_REG_11__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_4__3__SCAN_IN), .A3(n11533), .A4(n22004), .ZN(n22008)
         );
  INV_X1 U24946 ( .A(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n22020) );
  NAND4_X1 U24947 ( .A1(n22021), .A2(n22005), .A3(n22020), .A4(n22018), .ZN(
        n22007) );
  NAND4_X1 U24948 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(
        P3_EAX_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .A4(
        P2_LWORD_REG_4__SCAN_IN), .ZN(n22006) );
  NOR4_X1 U24949 ( .A1(n22009), .A2(n22008), .A3(n22007), .A4(n22006), .ZN(
        n22010) );
  NAND4_X1 U24950 ( .A1(n22013), .A2(n22012), .A3(n22011), .A4(n22010), .ZN(
        n22014) );
  OAI21_X1 U24951 ( .B1(n22015), .B2(n22014), .A(P1_DATAO_REG_11__SCAN_IN), 
        .ZN(n22143) );
  AOI22_X1 U24952 ( .A1(n22018), .A2(keyinput29), .B1(keyinput117), .B2(n22017), .ZN(n22016) );
  OAI221_X1 U24953 ( .B1(n22018), .B2(keyinput29), .C1(n22017), .C2(
        keyinput117), .A(n22016), .ZN(n22031) );
  AOI22_X1 U24954 ( .A1(n22021), .A2(keyinput96), .B1(keyinput77), .B2(n22020), 
        .ZN(n22019) );
  OAI221_X1 U24955 ( .B1(n22021), .B2(keyinput96), .C1(n22020), .C2(keyinput77), .A(n22019), .ZN(n22030) );
  AOI22_X1 U24956 ( .A1(n22024), .A2(keyinput30), .B1(n22023), .B2(keyinput25), 
        .ZN(n22022) );
  OAI221_X1 U24957 ( .B1(n22024), .B2(keyinput30), .C1(n22023), .C2(keyinput25), .A(n22022), .ZN(n22029) );
  XOR2_X1 U24958 ( .A(n22025), .B(keyinput118), .Z(n22027) );
  XNOR2_X1 U24959 ( .A(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B(keyinput71), .ZN(
        n22026) );
  NAND2_X1 U24960 ( .A1(n22027), .A2(n22026), .ZN(n22028) );
  NOR4_X1 U24961 ( .A1(n22031), .A2(n22030), .A3(n22029), .A4(n22028), .ZN(
        n22076) );
  AOI22_X1 U24962 ( .A1(n22033), .A2(keyinput50), .B1(n12440), .B2(keyinput21), 
        .ZN(n22032) );
  OAI221_X1 U24963 ( .B1(n22033), .B2(keyinput50), .C1(n12440), .C2(keyinput21), .A(n22032), .ZN(n22044) );
  AOI22_X1 U24964 ( .A1(n12475), .A2(keyinput124), .B1(keyinput73), .B2(n22035), .ZN(n22034) );
  OAI221_X1 U24965 ( .B1(n12475), .B2(keyinput124), .C1(n22035), .C2(
        keyinput73), .A(n22034), .ZN(n22043) );
  AOI22_X1 U24966 ( .A1(n13896), .A2(keyinput85), .B1(n22037), .B2(keyinput81), 
        .ZN(n22036) );
  OAI221_X1 U24967 ( .B1(n13896), .B2(keyinput85), .C1(n22037), .C2(keyinput81), .A(n22036), .ZN(n22042) );
  AOI22_X1 U24968 ( .A1(n22040), .A2(keyinput43), .B1(keyinput35), .B2(n22039), 
        .ZN(n22038) );
  OAI221_X1 U24969 ( .B1(n22040), .B2(keyinput43), .C1(n22039), .C2(keyinput35), .A(n22038), .ZN(n22041) );
  NOR4_X1 U24970 ( .A1(n22044), .A2(n22043), .A3(n22042), .A4(n22041), .ZN(
        n22075) );
  AOI22_X1 U24971 ( .A1(n22047), .A2(keyinput106), .B1(n22046), .B2(keyinput0), 
        .ZN(n22045) );
  OAI221_X1 U24972 ( .B1(n22047), .B2(keyinput106), .C1(n22046), .C2(keyinput0), .A(n22045), .ZN(n22058) );
  AOI22_X1 U24973 ( .A1(n22049), .A2(keyinput92), .B1(n13265), .B2(keyinput14), 
        .ZN(n22048) );
  OAI221_X1 U24974 ( .B1(n22049), .B2(keyinput92), .C1(n13265), .C2(keyinput14), .A(n22048), .ZN(n22057) );
  AOI22_X1 U24975 ( .A1(n22051), .A2(keyinput104), .B1(n11675), .B2(keyinput94), .ZN(n22050) );
  OAI221_X1 U24976 ( .B1(n22051), .B2(keyinput104), .C1(n11675), .C2(
        keyinput94), .A(n22050), .ZN(n22056) );
  XOR2_X1 U24977 ( .A(n22052), .B(keyinput63), .Z(n22054) );
  XNOR2_X1 U24978 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(keyinput89), 
        .ZN(n22053) );
  NAND2_X1 U24979 ( .A1(n22054), .A2(n22053), .ZN(n22055) );
  NOR4_X1 U24980 ( .A1(n22058), .A2(n22057), .A3(n22056), .A4(n22055), .ZN(
        n22074) );
  AOI22_X1 U24981 ( .A1(n22061), .A2(keyinput67), .B1(keyinput18), .B2(n22060), 
        .ZN(n22059) );
  OAI221_X1 U24982 ( .B1(n22061), .B2(keyinput67), .C1(n22060), .C2(keyinput18), .A(n22059), .ZN(n22072) );
  AOI22_X1 U24983 ( .A1(n22063), .A2(keyinput12), .B1(n12626), .B2(keyinput74), 
        .ZN(n22062) );
  OAI221_X1 U24984 ( .B1(n22063), .B2(keyinput12), .C1(n12626), .C2(keyinput74), .A(n22062), .ZN(n22071) );
  AOI22_X1 U24985 ( .A1(n22066), .A2(keyinput126), .B1(n22065), .B2(
        keyinput119), .ZN(n22064) );
  OAI221_X1 U24986 ( .B1(n22066), .B2(keyinput126), .C1(n22065), .C2(
        keyinput119), .A(n22064), .ZN(n22070) );
  XOR2_X1 U24987 ( .A(n12478), .B(keyinput84), .Z(n22068) );
  XNOR2_X1 U24988 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B(keyinput103), .ZN(
        n22067) );
  NAND2_X1 U24989 ( .A1(n22068), .A2(n22067), .ZN(n22069) );
  NOR4_X1 U24990 ( .A1(n22072), .A2(n22071), .A3(n22070), .A4(n22069), .ZN(
        n22073) );
  NAND4_X1 U24991 ( .A1(n22076), .A2(n22075), .A3(n22074), .A4(n22073), .ZN(
        n22142) );
  AOI22_X1 U24992 ( .A1(n22079), .A2(keyinput102), .B1(keyinput99), .B2(n22078), .ZN(n22077) );
  OAI221_X1 U24993 ( .B1(n22079), .B2(keyinput102), .C1(n22078), .C2(
        keyinput99), .A(n22077), .ZN(n22091) );
  AOI22_X1 U24994 ( .A1(n22081), .A2(keyinput78), .B1(n15141), .B2(keyinput15), 
        .ZN(n22080) );
  OAI221_X1 U24995 ( .B1(n22081), .B2(keyinput78), .C1(n15141), .C2(keyinput15), .A(n22080), .ZN(n22090) );
  INV_X1 U24996 ( .A(P3_DATAO_REG_6__SCAN_IN), .ZN(n22084) );
  AOI22_X1 U24997 ( .A1(n22084), .A2(keyinput4), .B1(n22083), .B2(keyinput51), 
        .ZN(n22082) );
  OAI221_X1 U24998 ( .B1(n22084), .B2(keyinput4), .C1(n22083), .C2(keyinput51), 
        .A(n22082), .ZN(n22089) );
  XOR2_X1 U24999 ( .A(n22085), .B(keyinput1), .Z(n22087) );
  XNOR2_X1 U25000 ( .A(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B(keyinput10), .ZN(
        n22086) );
  NAND2_X1 U25001 ( .A1(n22087), .A2(n22086), .ZN(n22088) );
  NOR4_X1 U25002 ( .A1(n22091), .A2(n22090), .A3(n22089), .A4(n22088), .ZN(
        n22140) );
  AOI22_X1 U25003 ( .A1(n22094), .A2(keyinput61), .B1(keyinput39), .B2(n22093), 
        .ZN(n22092) );
  OAI221_X1 U25004 ( .B1(n22094), .B2(keyinput61), .C1(n22093), .C2(keyinput39), .A(n22092), .ZN(n22107) );
  AOI22_X1 U25005 ( .A1(n22097), .A2(keyinput36), .B1(n22096), .B2(keyinput122), .ZN(n22095) );
  OAI221_X1 U25006 ( .B1(n22097), .B2(keyinput36), .C1(n22096), .C2(
        keyinput122), .A(n22095), .ZN(n22106) );
  AOI22_X1 U25007 ( .A1(n22100), .A2(keyinput47), .B1(keyinput37), .B2(n22099), 
        .ZN(n22098) );
  OAI221_X1 U25008 ( .B1(n22100), .B2(keyinput47), .C1(n22099), .C2(keyinput37), .A(n22098), .ZN(n22105) );
  XOR2_X1 U25009 ( .A(n22101), .B(keyinput20), .Z(n22103) );
  XNOR2_X1 U25010 ( .A(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B(keyinput52), .ZN(
        n22102) );
  NAND2_X1 U25011 ( .A1(n22103), .A2(n22102), .ZN(n22104) );
  NOR4_X1 U25012 ( .A1(n22107), .A2(n22106), .A3(n22105), .A4(n22104), .ZN(
        n22139) );
  AOI22_X1 U25013 ( .A1(n22110), .A2(keyinput54), .B1(keyinput7), .B2(n22109), 
        .ZN(n22108) );
  OAI221_X1 U25014 ( .B1(n22110), .B2(keyinput54), .C1(n22109), .C2(keyinput7), 
        .A(n22108), .ZN(n22122) );
  AOI22_X1 U25015 ( .A1(n22112), .A2(keyinput88), .B1(n12452), .B2(keyinput90), 
        .ZN(n22111) );
  OAI221_X1 U25016 ( .B1(n22112), .B2(keyinput88), .C1(n12452), .C2(keyinput90), .A(n22111), .ZN(n22121) );
  AOI22_X1 U25017 ( .A1(n22115), .A2(keyinput76), .B1(n22114), .B2(keyinput79), 
        .ZN(n22113) );
  OAI221_X1 U25018 ( .B1(n22115), .B2(keyinput76), .C1(n22114), .C2(keyinput79), .A(n22113), .ZN(n22120) );
  AOI22_X1 U25019 ( .A1(n22118), .A2(keyinput123), .B1(n22117), .B2(keyinput55), .ZN(n22116) );
  OAI221_X1 U25020 ( .B1(n22118), .B2(keyinput123), .C1(n22117), .C2(
        keyinput55), .A(n22116), .ZN(n22119) );
  NOR4_X1 U25021 ( .A1(n22122), .A2(n22121), .A3(n22120), .A4(n22119), .ZN(
        n22138) );
  AOI22_X1 U25022 ( .A1(n22124), .A2(keyinput69), .B1(keyinput11), .B2(n13791), 
        .ZN(n22123) );
  OAI221_X1 U25023 ( .B1(n22124), .B2(keyinput69), .C1(n13791), .C2(keyinput11), .A(n22123), .ZN(n22136) );
  AOI22_X1 U25024 ( .A1(n12815), .A2(keyinput80), .B1(keyinput42), .B2(n22126), 
        .ZN(n22125) );
  OAI221_X1 U25025 ( .B1(n12815), .B2(keyinput80), .C1(n22126), .C2(keyinput42), .A(n22125), .ZN(n22135) );
  AOI22_X1 U25026 ( .A1(n22129), .A2(keyinput24), .B1(n22128), .B2(keyinput82), 
        .ZN(n22127) );
  OAI221_X1 U25027 ( .B1(n22129), .B2(keyinput24), .C1(n22128), .C2(keyinput82), .A(n22127), .ZN(n22134) );
  XOR2_X1 U25028 ( .A(n22130), .B(keyinput49), .Z(n22132) );
  XNOR2_X1 U25029 ( .A(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B(keyinput13), .ZN(
        n22131) );
  NAND2_X1 U25030 ( .A1(n22132), .A2(n22131), .ZN(n22133) );
  NOR4_X1 U25031 ( .A1(n22136), .A2(n22135), .A3(n22134), .A4(n22133), .ZN(
        n22137) );
  NAND4_X1 U25032 ( .A1(n22140), .A2(n22139), .A3(n22138), .A4(n22137), .ZN(
        n22141) );
  AOI211_X1 U25033 ( .C1(keyinput60), .C2(n22143), .A(n22142), .B(n22141), 
        .ZN(n22144) );
  NAND4_X1 U25034 ( .A1(n22147), .A2(n22146), .A3(n22145), .A4(n22144), .ZN(
        n22148) );
  XNOR2_X1 U25035 ( .A(n22149), .B(n22148), .ZN(P2_U3079) );
  NOR2_X2 U11170 ( .A1(n11889), .A2(n22115), .ZN(n17879) );
  INV_X1 U15139 ( .A(n18427), .ZN(n19213) );
  NAND2_X1 U12706 ( .A1(n9733), .A2(n18398), .ZN(n18406) );
  NOR2_X1 U13731 ( .A1(n18299), .A2(n10450), .ZN(n18292) );
  NOR2_X1 U15189 ( .A1(n19099), .A2(n18331), .ZN(n18330) );
  NOR2_X1 U15191 ( .A1(n19076), .A2(n18314), .ZN(n18313) );
  NOR2_X1 U12467 ( .A1(n19083), .A2(n18321), .ZN(n18320) );
  NOR2_X1 U12691 ( .A1(n18262), .A2(n18261), .ZN(n18260) );
  NOR2_X1 U15192 ( .A1(n18273), .A2(n18272), .ZN(n18271) );
  NOR2_X1 U12702 ( .A1(n19157), .A2(n18371), .ZN(n18370) );
  NOR2_X1 U12697 ( .A1(n18342), .A2(n19115), .ZN(n18341) );
  OR2_X1 U11149 ( .A1(n18292), .A2(n10447), .ZN(n10445) );
  NAND2_X1 U13492 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18545) );
  INV_X1 U15289 ( .A(n9781), .ZN(n17631) );
  INV_X1 U11246 ( .A(n12206), .ZN(n12901) );
  INV_X1 U11159 ( .A(n14457), .ZN(n17985) );
  INV_X1 U13102 ( .A(n10450), .ZN(n10451) );
  AND2_X2 U11274 ( .A1(n9727), .A2(n12129), .ZN(n15177) );
  CLKBUF_X1 U11169 ( .A(n12177), .Z(n9726) );
  CLKBUF_X1 U11182 ( .A(n12245), .Z(n12254) );
  NOR2_X1 U11197 ( .A1(n11875), .A2(n10438), .ZN(n10437) );
  CLKBUF_X1 U11209 ( .A(n12248), .Z(n12857) );
  CLKBUF_X2 U11221 ( .A(n13223), .Z(n12812) );
  AND4_X1 U11222 ( .A1(n11867), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n18426) );
  AND2_X1 U11223 ( .A1(n11891), .A2(n11868), .ZN(n9737) );
  NAND2_X2 U11244 ( .A1(n10020), .A2(n14410), .ZN(n19198) );
  CLKBUF_X1 U11310 ( .A(n14384), .Z(n9707) );
  CLKBUF_X1 U11324 ( .A(n17113), .Z(n9701) );
  XNOR2_X1 U11341 ( .A(n11887), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11894) );
  CLKBUF_X1 U11561 ( .A(n20113), .Z(n18584) );
  MUX2_X1 U12243 ( .A(n15030), .B(n11654), .S(n15378), .Z(n11656) );
  CLKBUF_X1 U12473 ( .A(n12900), .Z(n14426) );
  CLKBUF_X1 U12696 ( .A(n14287), .Z(n17530) );
  CLKBUF_X1 U12711 ( .A(n12551), .Z(n15209) );
  CLKBUF_X1 U12788 ( .A(n20486), .Z(n9708) );
  CLKBUF_X1 U12840 ( .A(n18218), .Z(n18227) );
  CLKBUF_X3 U13211 ( .A(n12898), .Z(n9987) );
endmodule

