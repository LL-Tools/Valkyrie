

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput63, keyinput62, keyinput61, 
        keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, 
        keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, 
        keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, 
        keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, 
        keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, 
        keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, 
        keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, 
        keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, 
        keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, 
        keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, 
        keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput63, keyinput62,
         keyinput61, keyinput60, keyinput59, keyinput58, keyinput57,
         keyinput56, keyinput55, keyinput54, keyinput53, keyinput52,
         keyinput51, keyinput50, keyinput49, keyinput48, keyinput47,
         keyinput46, keyinput45, keyinput44, keyinput43, keyinput42,
         keyinput41, keyinput40, keyinput39, keyinput38, keyinput37,
         keyinput36, keyinput35, keyinput34, keyinput33, keyinput32,
         keyinput31, keyinput30, keyinput29, keyinput28, keyinput27,
         keyinput26, keyinput25, keyinput24, keyinput23, keyinput22,
         keyinput21, keyinput20, keyinput19, keyinput18, keyinput17,
         keyinput16, keyinput15, keyinput14, keyinput13, keyinput12,
         keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6,
         keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707;

  CLKBUF_X2 U3405 ( .A(n4116), .Z(n5555) );
  AND2_X1 U3406 ( .A1(n3118), .A2(n5313), .ZN(n5414) );
  INV_X2 U3407 ( .A(n5673), .ZN(n5409) );
  INV_X4 U3408 ( .A(n4079), .ZN(n5673) );
  OR2_X1 U3409 ( .A1(n4303), .A2(n3637), .ZN(n3639) );
  CLKBUF_X2 U3410 ( .A(n4003), .Z(n4749) );
  XNOR2_X1 U3411 ( .A(n3020), .B(n4222), .ZN(n4261) );
  AND2_X1 U3412 ( .A1(n3018), .A2(n3017), .ZN(n4222) );
  CLKBUF_X2 U3413 ( .A(n3583), .Z(n2957) );
  CLKBUF_X2 U3414 ( .A(n3585), .Z(n3942) );
  CLKBUF_X2 U3415 ( .A(n3274), .Z(n3941) );
  OR2_X2 U3416 ( .A1(n3012), .A2(n3011), .ZN(n4465) );
  BUF_X2 U3417 ( .A(n3238), .Z(n3940) );
  AND2_X1 U3418 ( .A1(n4337), .A2(n4366), .ZN(n3586) );
  INV_X1 U3419 ( .A(n4465), .ZN(n3514) );
  CLKBUF_X2 U3420 ( .A(n3238), .Z(n3782) );
  AND4_X1 U3421 ( .A1(n3130), .A2(n3129), .A3(n3128), .A4(n3127), .ZN(n3146)
         );
  AND2_X1 U3422 ( .A1(n4421), .A2(n4460), .ZN(n3019) );
  BUF_X1 U3423 ( .A(n3019), .Z(n4214) );
  INV_X1 U3425 ( .A(n5026), .ZN(n4631) );
  AND2_X1 U3426 ( .A1(n5123), .A2(n4842), .ZN(n6044) );
  OR2_X1 U3427 ( .A1(n5326), .A2(n5327), .ZN(n5491) );
  NAND2_X1 U3428 ( .A1(n3639), .A2(n4304), .ZN(n4302) );
  INV_X1 U3429 ( .A(n6044), .ZN(n6030) );
  XNOR2_X1 U3430 ( .A(n3126), .B(n3125), .ZN(n5701) );
  OR2_X1 U3431 ( .A1(n5345), .A2(n5344), .ZN(n5582) );
  INV_X1 U3432 ( .A(n3224), .ZN(n3381) );
  OAI211_X2 U3433 ( .C1(n4157), .C2(n3487), .A(n4248), .B(n5920), .ZN(n3484)
         );
  NAND2_X1 U3434 ( .A1(n3219), .A2(n4455), .ZN(n3248) );
  NAND2_X2 U3435 ( .A1(n3545), .A2(n3544), .ZN(n3548) );
  NOR2_X2 U3436 ( .A1(n5387), .A2(n4325), .ZN(n4405) );
  NOR2_X4 U3437 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n2976) );
  OAI21_X2 U3438 ( .B1(n5555), .B2(n5522), .A(n5655), .ZN(n5667) );
  OAI22_X1 U3439 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n5352), .B1(n5351), .B2(n5350), .ZN(n5353) );
  AOI211_X1 U3440 ( .C1(n5440), .C2(n5883), .A(n5435), .B(n5434), .ZN(n5436)
         );
  AOI211_X1 U3441 ( .C1(n5883), .C2(n5670), .A(n5669), .B(n5668), .ZN(n5671)
         );
  AND2_X1 U3442 ( .A1(n4101), .A2(n5662), .ZN(n5652) );
  OR2_X1 U3443 ( .A1(n5655), .A2(n5656), .ZN(n5653) );
  CLKBUF_X1 U3444 ( .A(n5220), .Z(n5237) );
  NAND2_X1 U34450 ( .A1(n5144), .A2(n5145), .ZN(n5148) );
  NOR2_X1 U34460 ( .A1(n3832), .A2(n3831), .ZN(n3833) );
  AND2_X1 U34470 ( .A1(n4838), .A2(n2960), .ZN(n5097) );
  CLKBUF_X1 U34480 ( .A(n4613), .Z(n4836) );
  NAND2_X1 U3449 ( .A1(n3731), .A2(n3730), .ZN(n4518) );
  AND2_X1 U3450 ( .A1(n5100), .A2(n5103), .ZN(n4082) );
  INV_X1 U34510 ( .A(n4323), .ZN(n3731) );
  INV_X1 U34520 ( .A(n4402), .ZN(n3730) );
  AND2_X1 U34530 ( .A1(n3684), .A2(n3714), .ZN(n4003) );
  NOR2_X1 U3454 ( .A1(n5242), .A2(n5243), .ZN(n5241) );
  INV_X1 U34550 ( .A(n3640), .ZN(n3681) );
  AND2_X1 U34560 ( .A1(n3612), .A2(n3611), .ZN(n3640) );
  CLKBUF_X1 U3457 ( .A(n4331), .Z(n6038) );
  NAND2_X2 U3458 ( .A1(n5562), .A2(n4289), .ZN(n5877) );
  NAND2_X1 U34590 ( .A1(n3643), .A2(n3642), .ZN(n4361) );
  NAND2_X1 U34600 ( .A1(n3563), .A2(n3562), .ZN(n3616) );
  AND2_X1 U34610 ( .A1(n3500), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3527) );
  AND2_X1 U34620 ( .A1(n3498), .A2(n4168), .ZN(n3523) );
  INV_X1 U34630 ( .A(n3486), .ZN(n4108) );
  INV_X2 U34640 ( .A(n4214), .ZN(n4260) );
  BUF_X1 U34650 ( .A(n3248), .Z(n4212) );
  INV_X1 U3466 ( .A(n3491), .ZN(n3481) );
  CLKBUF_X1 U3467 ( .A(n3219), .Z(n5309) );
  AND2_X1 U34680 ( .A1(n4058), .A2(n4237), .ZN(n4153) );
  NAND2_X1 U34690 ( .A1(n2965), .A2(n2966), .ZN(n3491) );
  INV_X1 U34700 ( .A(n4455), .ZN(n3518) );
  CLKBUF_X1 U34710 ( .A(n3231), .Z(n4474) );
  INV_X1 U34720 ( .A(n3245), .ZN(n4237) );
  BUF_X2 U34730 ( .A(n3245), .Z(n4479) );
  AND4_X1 U34740 ( .A1(n2986), .A2(n2985), .A3(n2984), .A4(n2983), .ZN(n3002)
         );
  AND4_X1 U3475 ( .A1(n3213), .A2(n3212), .A3(n3211), .A4(n3210), .ZN(n3218)
         );
  AND4_X1 U3476 ( .A1(n3138), .A2(n3137), .A3(n3136), .A4(n3135), .ZN(n3144)
         );
  BUF_X2 U3477 ( .A(n3592), .Z(n3939) );
  BUF_X2 U3478 ( .A(n3587), .Z(n3938) );
  BUF_X2 U3479 ( .A(n3593), .Z(n2958) );
  CLKBUF_X2 U3480 ( .A(n3593), .Z(n2959) );
  BUF_X2 U3481 ( .A(n3586), .Z(n3948) );
  BUF_X2 U3482 ( .A(n3273), .Z(n3947) );
  BUF_X2 U3483 ( .A(n3584), .Z(n3949) );
  BUF_X2 U3484 ( .A(n3594), .Z(n3952) );
  AND2_X2 U3485 ( .A1(n4192), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4164)
         );
  CLKBUF_X1 U3486 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n6552) );
  NOR2_X2 U3487 ( .A1(n5255), .A2(n5254), .ZN(n5291) );
  AND2_X4 U3488 ( .A1(n4164), .A2(n4337), .ZN(n3376) );
  NOR2_X2 U3489 ( .A1(n5908), .A2(n5909), .ZN(n5910) );
  NOR2_X2 U3490 ( .A1(n5992), .A2(n5993), .ZN(n5991) );
  AND2_X1 U3491 ( .A1(n4094), .A2(n5270), .ZN(n4095) );
  INV_X1 U3492 ( .A(n6552), .ZN(n3532) );
  OR2_X1 U3493 ( .A1(n3561), .A2(n3560), .ZN(n4016) );
  NAND2_X1 U3494 ( .A1(n4400), .A2(n4324), .ZN(n4323) );
  NAND2_X1 U3495 ( .A1(n3735), .A2(n3734), .ZN(n4059) );
  OR2_X1 U3496 ( .A1(n4069), .A2(n4068), .ZN(n4074) );
  AND2_X1 U3497 ( .A1(n3160), .A2(n4479), .ZN(n3736) );
  XNOR2_X1 U3498 ( .A(n4361), .B(n4716), .ZN(n4331) );
  NAND2_X1 U3499 ( .A1(n3921), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n2992) );
  AND4_X1 U3500 ( .A1(n3134), .A2(n3133), .A3(n3132), .A4(n3131), .ZN(n3145)
         );
  NAND2_X2 U3501 ( .A1(n3156), .A2(n3155), .ZN(n3231) );
  INV_X1 U3502 ( .A(n4869), .ZN(n4156) );
  NAND2_X1 U3503 ( .A1(n3244), .A2(n4460), .ZN(n4157) );
  BUF_X1 U3504 ( .A(n3483), .Z(n4179) );
  NAND2_X1 U3505 ( .A1(n4130), .A2(n4171), .ZN(n4869) );
  AND2_X1 U3506 ( .A1(n4237), .A2(n4455), .ZN(n4282) );
  INV_X1 U3507 ( .A(n3476), .ZN(n3474) );
  OAI21_X1 U3508 ( .B1(n4080), .B2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(n5673), 
        .ZN(n4084) );
  NAND2_X1 U3509 ( .A1(n4104), .A2(n4103), .ZN(n5644) );
  NAND2_X1 U3510 ( .A1(n6529), .A2(n4420), .ZN(n4754) );
  NAND2_X1 U3511 ( .A1(n5598), .A2(n3979), .ZN(n3993) );
  AND2_X1 U3512 ( .A1(n5562), .A2(n5310), .ZN(n6077) );
  OR2_X1 U3513 ( .A1(n4309), .A2(n6402), .ZN(n6166) );
  NAND2_X1 U3514 ( .A1(n3124), .A2(n3123), .ZN(n3126) );
  INV_X1 U3515 ( .A(n5420), .ZN(n3123) );
  NAND2_X1 U3516 ( .A1(n5352), .A2(n4106), .ZN(n4107) );
  NOR2_X1 U3517 ( .A1(n4421), .A2(n3480), .ZN(n3487) );
  CLKBUF_X1 U3518 ( .A(n3921), .Z(n3951) );
  NAND2_X1 U3519 ( .A1(n3625), .A2(n3995), .ZN(n3615) );
  NAND2_X1 U3520 ( .A1(n4495), .A2(n6529), .ZN(n3563) );
  OAI21_X1 U3521 ( .B1(n3533), .B2(n3532), .A(n3531), .ZN(n3642) );
  INV_X1 U3522 ( .A(n3644), .ZN(n3533) );
  NAND2_X1 U3523 ( .A1(n5222), .A2(n5221), .ZN(n5220) );
  BUF_X1 U3524 ( .A(n3518), .Z(n4241) );
  AND2_X1 U3525 ( .A1(n4214), .A2(n5530), .ZN(n3075) );
  CLKBUF_X1 U3526 ( .A(n3031), .Z(n3105) );
  NAND2_X1 U3527 ( .A1(n3510), .A2(n3509), .ZN(n3576) );
  XNOR2_X1 U3528 ( .A(n3641), .B(n3642), .ZN(n4345) );
  INV_X1 U3529 ( .A(n3581), .ZN(n3549) );
  AND3_X1 U3530 ( .A1(n3519), .A2(n3247), .A3(n5308), .ZN(n3494) );
  CLKBUF_X1 U3531 ( .A(n3527), .Z(n3644) );
  OAI21_X1 U3532 ( .B1(n6535), .B2(n4367), .A(n6550), .ZN(n4420) );
  NAND2_X1 U3533 ( .A1(n4331), .A2(n6529), .ZN(n3662) );
  INV_X1 U3534 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6399) );
  AND2_X2 U3535 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4359) );
  NAND2_X1 U3536 ( .A1(n3606), .A2(n3546), .ZN(n3737) );
  AND2_X1 U3537 ( .A1(n3204), .A2(n3203), .ZN(n3250) );
  CLKBUF_X1 U3538 ( .A(n4166), .Z(n4247) );
  INV_X1 U3539 ( .A(n6021), .ZN(n5118) );
  INV_X1 U3540 ( .A(n6523), .ZN(n4893) );
  OR2_X1 U3541 ( .A1(n4309), .A2(n4157), .ZN(n4263) );
  OR2_X1 U3542 ( .A1(n3267), .A2(n5465), .ZN(n3476) );
  AND2_X1 U3543 ( .A1(n5555), .A2(n5321), .ZN(n5377) );
  AND2_X1 U3544 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n3264), .ZN(n3393)
         );
  INV_X1 U3545 ( .A(n3413), .ZN(n3264) );
  NOR2_X1 U3546 ( .A1(n3862), .A2(n3861), .ZN(n3879) );
  OR2_X1 U3547 ( .A1(n3847), .A2(n5231), .ZN(n3862) );
  OR2_X2 U3548 ( .A1(n5220), .A2(n5238), .ZN(n5255) );
  NAND2_X1 U3549 ( .A1(n5148), .A2(n3846), .ZN(n5222) );
  AND2_X1 U3550 ( .A1(n3812), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3826)
         );
  OR2_X1 U3552 ( .A1(n3742), .A2(n3741), .ZN(n3757) );
  NOR2_X1 U3553 ( .A1(n6569), .A2(n3757), .ZN(n3776) );
  NOR2_X1 U3554 ( .A1(n3707), .A2(n4874), .ZN(n3725) );
  AOI21_X1 U3555 ( .B1(n4057), .B2(n3871), .A(n3729), .ZN(n4402) );
  NAND2_X1 U3556 ( .A1(n3710), .A2(n3709), .ZN(n4324) );
  NAND2_X1 U3557 ( .A1(n4046), .A2(n3871), .ZN(n3710) );
  BUF_X1 U3558 ( .A(n4323), .Z(n4403) );
  AND2_X1 U3559 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n3685), .ZN(n3687)
         );
  NAND2_X1 U3560 ( .A1(n3687), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3707)
         );
  NOR2_X2 U3561 ( .A1(n4302), .A2(n3692), .ZN(n4400) );
  NAND2_X1 U3562 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3631) );
  CLKBUF_X1 U3563 ( .A(n5326), .Z(n5373) );
  NOR2_X2 U3564 ( .A1(n5513), .A2(n5392), .ZN(n5394) );
  AND2_X1 U3565 ( .A1(n5241), .A2(n3090), .ZN(n5545) );
  OAI21_X1 U3566 ( .B1(n5661), .B2(n5663), .A(n4079), .ZN(n4101) );
  CLKBUF_X1 U3567 ( .A(n4104), .Z(n5650) );
  NAND2_X1 U3568 ( .A1(n5910), .A2(n5226), .ZN(n5242) );
  CLKBUF_X1 U3569 ( .A(n5241), .Z(n5773) );
  CLKBUF_X1 U3570 ( .A(n5112), .Z(n5163) );
  BUF_X1 U3571 ( .A(n5129), .Z(n5152) );
  BUF_X1 U3572 ( .A(n4958), .Z(n5101) );
  NOR2_X1 U3573 ( .A1(n4320), .A2(n4321), .ZN(n5385) );
  NAND2_X1 U3574 ( .A1(n5385), .A2(n5386), .ZN(n5387) );
  AND2_X1 U3575 ( .A1(n5822), .A2(n5819), .ZN(n5771) );
  NAND2_X1 U3576 ( .A1(n4236), .A2(n4235), .ZN(n4251) );
  XNOR2_X1 U3577 ( .A(n3682), .B(n3640), .ZN(n4010) );
  CLKBUF_X1 U3578 ( .A(n4345), .Z(n5117) );
  INV_X1 U3579 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n2969) );
  INV_X1 U3580 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n2971) );
  OR2_X1 U3581 ( .A1(n4190), .A2(n4286), .ZN(n6391) );
  INV_X1 U3582 ( .A(n4369), .ZN(n4600) );
  AND4_X1 U3583 ( .A1(n2990), .A2(n2989), .A3(n2988), .A4(n2987), .ZN(n3001)
         );
  AND4_X1 U3584 ( .A1(n2998), .A2(n2997), .A3(n2996), .A4(n2995), .ZN(n2999)
         );
  AND3_X1 U3585 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6529), .A3(n4420), .ZN(
        n4484) );
  INV_X1 U3586 ( .A(n6024), .ZN(n6033) );
  AND2_X1 U3587 ( .A1(n5123), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6008) );
  AND2_X1 U3588 ( .A1(n4219), .A2(n4284), .ZN(n6065) );
  CLKBUF_X1 U3589 ( .A(n5438), .Z(n5451) );
  NAND2_X1 U3590 ( .A1(n4287), .A2(n6143), .ZN(n5562) );
  OR2_X1 U3591 ( .A1(n3975), .A2(n6571), .ZN(n3977) );
  AOI21_X1 U3592 ( .B1(n5656), .B2(n5655), .A(n5654), .ZN(n5878) );
  CLKBUF_X1 U3593 ( .A(n5137), .Z(n5139) );
  INV_X1 U3594 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4874) );
  INV_X1 U3595 ( .A(n6242), .ZN(n6263) );
  NAND2_X2 U3596 ( .A1(n3625), .A2(n3624), .ZN(n5026) );
  CLKBUF_X1 U3597 ( .A(n3626), .Z(n4903) );
  INV_X1 U3598 ( .A(n4600), .ZN(n5830) );
  OAI21_X1 U3599 ( .B1(n5066), .B2(n6512), .A(n5060), .ZN(n5088) );
  OR2_X1 U3600 ( .A1(n4225), .A2(n6512), .ZN(n6550) );
  INV_X1 U3601 ( .A(n3262), .ZN(n3994) );
  OAI21_X1 U3602 ( .B1(n5845), .B2(n6164), .A(n4126), .ZN(n4127) );
  AND2_X2 U3603 ( .A1(n4171), .A2(n4460), .ZN(n3496) );
  INV_X2 U3605 ( .A(n3381), .ZN(n3915) );
  INV_X1 U3606 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6529) );
  NOR4_X2 U3607 ( .A1(n5942), .A2(n5941), .A3(n5940), .A4(n5939), .ZN(n6516)
         );
  INV_X1 U3608 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4344) );
  NOR2_X1 U3609 ( .A1(n5095), .A2(n4911), .ZN(n2960) );
  OR4_X1 U3610 ( .A1(n5459), .A2(REIP_REG_31__SCAN_IN), .A3(n6505), .A4(n6501), 
        .ZN(n2961) );
  AND2_X1 U3611 ( .A1(n4079), .A2(n5405), .ZN(n2962) );
  NAND2_X1 U3612 ( .A1(n5409), .A2(n4097), .ZN(n2963) );
  NAND2_X1 U3613 ( .A1(n5409), .A2(n4090), .ZN(n2964) );
  AND4_X1 U3614 ( .A1(n3236), .A2(n3235), .A3(n3234), .A4(n3233), .ZN(n2965)
         );
  OR2_X1 U3615 ( .A1(n5308), .A2(n6522), .ZN(n3930) );
  AND4_X1 U3616 ( .A1(n3242), .A2(n3241), .A3(n3240), .A4(n3239), .ZN(n2966)
         );
  AND4_X1 U3617 ( .A1(n3217), .A2(n3216), .A3(n3215), .A4(n3214), .ZN(n2967)
         );
  OR2_X1 U3618 ( .A1(n4079), .A2(n4086), .ZN(n2968) );
  INV_X1 U3619 ( .A(n4460), .ZN(n4130) );
  AOI21_X1 U3620 ( .B1(n3492), .B2(n4450), .A(n4421), .ZN(n3493) );
  BUF_X1 U3621 ( .A(n3650), .Z(n3937) );
  INV_X1 U3622 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n2970) );
  NAND2_X1 U3623 ( .A1(n3527), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3510) );
  AND2_X1 U3624 ( .A1(n3248), .A2(n5308), .ZN(n3485) );
  INV_X1 U3625 ( .A(n3119), .ZN(n3031) );
  NAND2_X1 U3626 ( .A1(n5097), .A2(n5110), .ZN(n3832) );
  OR2_X1 U3627 ( .A1(n3714), .A2(n3713), .ZN(n3732) );
  AND2_X1 U3628 ( .A1(n2964), .A2(n5280), .ZN(n4089) );
  INV_X1 U3629 ( .A(n3732), .ZN(n3735) );
  AOI21_X1 U3630 ( .B1(n3527), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n3504), 
        .ZN(n3503) );
  NOR2_X2 U3631 ( .A1(n2970), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4333)
         );
  OR2_X1 U3632 ( .A1(n4150), .A2(n3524), .ZN(n3577) );
  AND4_X1 U3633 ( .A1(n3142), .A2(n3141), .A3(n3140), .A4(n3139), .ZN(n3143)
         );
  NAND2_X1 U3634 ( .A1(n3481), .A2(n4465), .ZN(n4017) );
  NOR2_X1 U3635 ( .A1(n3392), .A2(n3265), .ZN(n3357) );
  INV_X1 U3636 ( .A(n3231), .ZN(n3219) );
  NOR2_X1 U3637 ( .A1(n4257), .A2(n3638), .ZN(n3637) );
  AND4_X1 U3638 ( .A1(n3154), .A2(n3153), .A3(n3152), .A4(n3151), .ZN(n3155)
         );
  AND2_X1 U3639 ( .A1(n4172), .A2(n4359), .ZN(n3592) );
  AND2_X1 U3640 ( .A1(n5269), .A2(n4087), .ZN(n4088) );
  OR2_X1 U3641 ( .A1(n3573), .A2(n3572), .ZN(n4070) );
  AND2_X1 U3642 ( .A1(n5887), .A2(n4091), .ZN(n4092) );
  AND2_X1 U3643 ( .A1(n5279), .A2(n4089), .ZN(n5269) );
  INV_X1 U3644 ( .A(n5102), .ZN(n4081) );
  OR2_X1 U3645 ( .A1(n3600), .A2(n3599), .ZN(n4024) );
  NAND2_X1 U3646 ( .A1(n3576), .A2(n3577), .ZN(n3581) );
  NAND3_X1 U3647 ( .A1(n3682), .A2(n3681), .A3(n4626), .ZN(n3714) );
  OR2_X1 U3648 ( .A1(n4479), .A2(n6529), .ZN(n3606) );
  NAND4_X1 U3649 ( .A1(n3146), .A2(n3145), .A3(n3144), .A4(n3143), .ZN(n3245)
         );
  AND2_X1 U3650 ( .A1(n3914), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3412)
         );
  AND2_X1 U3651 ( .A1(n5478), .A2(n5464), .ZN(n3118) );
  INV_X1 U3652 ( .A(n5552), .ZN(n3935) );
  XNOR2_X1 U3653 ( .A(n3706), .B(n3711), .ZN(n4046) );
  OR2_X1 U3654 ( .A1(n3449), .A2(n3448), .ZN(n3451) );
  NOR2_X1 U3655 ( .A1(n3894), .A2(n5294), .ZN(n3912) );
  OR2_X1 U3656 ( .A1(n3807), .A2(n3263), .ZN(n3781) );
  XNOR2_X1 U3657 ( .A(n4059), .B(n3740), .ZN(n4067) );
  OR2_X1 U3658 ( .A1(n4093), .A2(n4092), .ZN(n5270) );
  NOR2_X1 U3659 ( .A1(n5164), .A2(n5165), .ZN(n5112) );
  INV_X1 U3660 ( .A(n3075), .ZN(n3112) );
  AND2_X1 U3661 ( .A1(n4243), .A2(n4224), .ZN(n4245) );
  NAND2_X1 U3662 ( .A1(n4283), .A2(n4141), .ZN(n4248) );
  NAND2_X1 U3663 ( .A1(n3581), .A2(n3580), .ZN(n3626) );
  AND2_X1 U3664 ( .A1(n4528), .A2(n5829), .ZN(n4530) );
  NAND2_X1 U3665 ( .A1(n3649), .A2(n3648), .ZN(n4716) );
  NAND2_X1 U3666 ( .A1(n3662), .A2(n3661), .ZN(n4626) );
  NAND2_X1 U3667 ( .A1(n3207), .A2(n3206), .ZN(n3209) );
  NAND2_X1 U3668 ( .A1(n3393), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3392)
         );
  NAND2_X1 U3669 ( .A1(n3412), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3413)
         );
  INV_X1 U3670 ( .A(n6008), .ZN(n6036) );
  NAND2_X1 U3671 ( .A1(n4231), .A2(n3982), .ZN(n6021) );
  BUF_X1 U3672 ( .A(n3118), .Z(n5417) );
  NAND2_X1 U3673 ( .A1(n5291), .A2(n5290), .ZN(n4112) );
  AND4_X1 U3674 ( .A1(n2994), .A2(n2993), .A3(n2992), .A4(n2991), .ZN(n3000)
         );
  NAND2_X1 U3675 ( .A1(n3474), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n3975)
         );
  AND2_X1 U3676 ( .A1(n3912), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3914)
         );
  NOR2_X1 U3677 ( .A1(n3781), .A2(n5983), .ZN(n3812) );
  AOI21_X1 U3678 ( .B1(n4067), .B2(n3871), .A(n3746), .ZN(n4519) );
  INV_X1 U3679 ( .A(n3631), .ZN(n3685) );
  NOR2_X1 U3680 ( .A1(n5411), .A2(n5625), .ZN(n5618) );
  NAND2_X1 U3681 ( .A1(n5588), .A2(n5408), .ZN(n5411) );
  NAND2_X1 U3682 ( .A1(n5652), .A2(n5651), .ZN(n4104) );
  OR2_X1 U3683 ( .A1(n5557), .A2(n5556), .ZN(n5559) );
  CLKBUF_X1 U3684 ( .A(n4520), .Z(n4616) );
  NAND2_X1 U3685 ( .A1(n4015), .A2(n4014), .ZN(n6173) );
  OR2_X1 U3686 ( .A1(n3026), .A2(n3025), .ZN(n4306) );
  AND2_X2 U3687 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6549) );
  INV_X1 U3688 ( .A(n6038), .ZN(n5064) );
  OR2_X1 U3689 ( .A1(n4492), .A2(n5830), .ZN(n4721) );
  OR2_X1 U3690 ( .A1(n4492), .A2(n4600), .ZN(n6326) );
  INV_X1 U3691 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6393) );
  XNOR2_X1 U3692 ( .A(n3617), .B(n3616), .ZN(n4369) );
  AND2_X1 U3693 ( .A1(n3609), .A2(n3608), .ZN(n3625) );
  NAND2_X1 U3694 ( .A1(n3209), .A2(n3208), .ZN(n4225) );
  INV_X1 U3695 ( .A(n5985), .ZN(n3979) );
  OR2_X1 U3696 ( .A1(n6523), .A2(n3259), .ZN(n5123) );
  AND2_X1 U3697 ( .A1(n4849), .A2(n6523), .ZN(n6032) );
  NOR2_X1 U3698 ( .A1(n5489), .A2(n5477), .ZN(n5478) );
  INV_X1 U3699 ( .A(n4112), .ZN(n5553) );
  INV_X1 U3700 ( .A(n6055), .ZN(n6060) );
  XNOR2_X1 U3701 ( .A(n5433), .B(n5432), .ZN(n5438) );
  AND2_X1 U3702 ( .A1(n4115), .A2(n4114), .ZN(n5345) );
  AND2_X1 U3703 ( .A1(n5562), .A2(n4290), .ZN(n5245) );
  AND2_X1 U3704 ( .A1(n4313), .A2(n4312), .ZN(n6093) );
  INV_X1 U3705 ( .A(n4311), .ZN(n6144) );
  AOI21_X1 U3706 ( .B1(n5379), .B2(n5378), .A(n5377), .ZN(n5538) );
  INV_X1 U3707 ( .A(n5676), .ZN(n6066) );
  NAND2_X1 U3708 ( .A1(n3826), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3847)
         );
  NAND2_X1 U3709 ( .A1(n3725), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3742)
         );
  INV_X1 U3710 ( .A(n6182), .ZN(n5883) );
  OR2_X1 U3711 ( .A1(n4225), .A2(n6424), .ZN(n4309) );
  BUF_X1 U3712 ( .A(n5411), .Z(n5627) );
  OR2_X1 U3713 ( .A1(n6184), .A2(n5821), .ZN(n6186) );
  NOR2_X1 U3714 ( .A1(n5771), .A2(n4429), .ZN(n6254) );
  INV_X1 U3715 ( .A(n6246), .ZN(n6258) );
  AND2_X1 U3716 ( .A1(n5830), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5834) );
  INV_X1 U3717 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4198) );
  INV_X1 U3718 ( .A(n4721), .ZN(n6307) );
  AND2_X1 U3719 ( .A1(n5835), .A2(n4371), .ZN(n4723) );
  OR2_X1 U3720 ( .A1(n4443), .A2(n4442), .ZN(n4490) );
  INV_X1 U3721 ( .A(n4534), .ZN(n4552) );
  OR2_X1 U3722 ( .A1(n4684), .A2(n4683), .ZN(n4708) );
  INV_X1 U3723 ( .A(n4678), .ZN(n4712) );
  AND2_X1 U3724 ( .A1(n4562), .A2(n4631), .ZN(n4953) );
  AND2_X1 U3725 ( .A1(n4632), .A2(n4631), .ZN(n4789) );
  NAND2_X1 U3726 ( .A1(n4263), .A2(n4134), .ZN(n6523) );
  NAND2_X1 U3727 ( .A1(n3991), .A2(REIP_REG_31__SCAN_IN), .ZN(n3992) );
  NAND2_X1 U3728 ( .A1(n5123), .A2(n3978), .ZN(n5985) );
  AND2_X1 U3729 ( .A1(n5985), .A2(n4870), .ZN(n6041) );
  OAI21_X1 U3730 ( .B1(n5345), .B2(n4118), .A(n5378), .ZN(n5845) );
  OR2_X1 U3731 ( .A1(n6093), .A2(n6112), .ZN(n6095) );
  INV_X1 U3732 ( .A(n6093), .ZN(n6118) );
  OR3_X1 U3733 ( .A1(n4309), .A2(READY_N), .A3(n4265), .ZN(n6143) );
  OR2_X1 U3734 ( .A1(n4263), .A2(n4421), .ZN(n4311) );
  INV_X1 U3735 ( .A(n4127), .ZN(n4128) );
  OR2_X1 U3736 ( .A1(n6171), .A2(n4208), .ZN(n6182) );
  INV_X1 U3737 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6691) );
  INV_X1 U3738 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4970) );
  NAND2_X1 U3739 ( .A1(n4601), .A2(n5026), .ZN(n6291) );
  NAND2_X1 U3740 ( .A1(n4723), .A2(n4722), .ZN(n5094) );
  OR2_X1 U3741 ( .A1(n4525), .A2(n5830), .ZN(n4978) );
  OR2_X1 U3742 ( .A1(n4527), .A2(n4493), .ZN(n6385) );
  OR2_X1 U3743 ( .A1(n4525), .A2(n4600), .ZN(n6378) );
  AND2_X2 U3744 ( .A1(n2969), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4172)
         );
  AND2_X2 U3745 ( .A1(n4172), .A2(n2976), .ZN(n3650) );
  AOI22_X1 U3746 ( .A1(n3592), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3650), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n2975) );
  AND2_X2 U3747 ( .A1(n4333), .A2(n4172), .ZN(n3224) );
  INV_X2 U3748 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4192) );
  AND2_X4 U3749 ( .A1(n4164), .A2(n2976), .ZN(n3921) );
  AOI22_X1 U3750 ( .A1(n3224), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n2974) );
  NOR2_X4 U3751 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4366) );
  AND2_X2 U3752 ( .A1(n4333), .A2(n4366), .ZN(n3593) );
  NOR2_X4 U3753 ( .A1(n2971), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4337)
         );
  AND2_X2 U3754 ( .A1(n4337), .A2(n6549), .ZN(n3583) );
  AOI22_X1 U3755 ( .A1(n2958), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3583), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n2973) );
  AND2_X2 U3756 ( .A1(n4333), .A2(n6549), .ZN(n3587) );
  AND2_X2 U3757 ( .A1(n4366), .A2(n4359), .ZN(n3237) );
  AOI22_X1 U3758 ( .A1(n3587), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3237), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n2972) );
  NAND4_X1 U3759 ( .A1(n2975), .A2(n2974), .A3(n2973), .A4(n2972), .ZN(n2982)
         );
  AND2_X2 U3760 ( .A1(n4172), .A2(n4337), .ZN(n3273) );
  AOI22_X1 U3761 ( .A1(n3376), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n2980) );
  AND2_X2 U3762 ( .A1(n4333), .A2(n4164), .ZN(n3584) );
  AND2_X2 U3763 ( .A1(n4164), .A2(n4359), .ZN(n3585) );
  AOI22_X1 U3764 ( .A1(n3584), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3585), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n2979) );
  AND2_X2 U3765 ( .A1(n4366), .A2(n2976), .ZN(n3238) );
  AND2_X2 U3766 ( .A1(n4359), .A2(n6549), .ZN(n3594) );
  AOI22_X1 U3767 ( .A1(n3940), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3594), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n2978) );
  AND2_X2 U3768 ( .A1(n2976), .A2(n6549), .ZN(n3274) );
  AOI22_X1 U3769 ( .A1(n3586), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3274), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n2977) );
  NAND4_X1 U3770 ( .A1(n2980), .A2(n2979), .A3(n2978), .A4(n2977), .ZN(n2981)
         );
  OR2_X4 U3771 ( .A1(n2982), .A2(n2981), .ZN(n4421) );
  NAND2_X1 U3772 ( .A1(n3592), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n2986)
         );
  NAND2_X1 U3773 ( .A1(n3224), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n2985)
         );
  NAND2_X1 U3774 ( .A1(n3587), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n2984)
         );
  NAND2_X1 U3775 ( .A1(n3583), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n2983) );
  NAND2_X1 U3776 ( .A1(n3376), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n2990) );
  NAND2_X1 U3777 ( .A1(n3273), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n2989) );
  NAND2_X1 U3778 ( .A1(n3585), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n2988)
         );
  NAND2_X1 U3779 ( .A1(n3586), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n2987) );
  NAND2_X1 U3780 ( .A1(n3650), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n2994) );
  NAND2_X1 U3781 ( .A1(n2958), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n2993) );
  BUF_X2 U3782 ( .A(n3237), .Z(n3922) );
  NAND2_X1 U3783 ( .A1(n3922), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n2991)
         );
  NAND2_X1 U3784 ( .A1(n3584), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n2998) );
  NAND2_X1 U3785 ( .A1(n3594), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n2997)
         );
  NAND2_X1 U3786 ( .A1(n3940), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n2996) );
  NAND2_X1 U3787 ( .A1(n3274), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n2995) );
  NAND4_X4 U3788 ( .A1(n3002), .A2(n3001), .A3(n3000), .A4(n2999), .ZN(n4460)
         );
  AOI22_X1 U3789 ( .A1(n3592), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3650), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3006) );
  AOI22_X1 U3790 ( .A1(n3224), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3005) );
  AOI22_X1 U3791 ( .A1(n2959), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3583), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3004) );
  AOI22_X1 U3792 ( .A1(n3587), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3237), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3003) );
  NAND4_X1 U3793 ( .A1(n3006), .A2(n3005), .A3(n3004), .A4(n3003), .ZN(n3012)
         );
  AOI22_X1 U3794 ( .A1(n3376), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3010) );
  AOI22_X1 U3795 ( .A1(n3584), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3585), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3009) );
  AOI22_X1 U3796 ( .A1(n3940), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3594), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3008) );
  AOI22_X1 U3797 ( .A1(n3586), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3274), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3007) );
  NAND4_X1 U3798 ( .A1(n3010), .A2(n3009), .A3(n3008), .A4(n3007), .ZN(n3011)
         );
  AND2_X4 U3799 ( .A1(n4465), .A2(n4421), .ZN(n5774) );
  NAND2_X2 U3800 ( .A1(n3019), .A2(n5774), .ZN(n3119) );
  INV_X1 U3801 ( .A(EBX_REG_1__SCAN_IN), .ZN(n3013) );
  NAND2_X1 U3802 ( .A1(n3031), .A2(n3013), .ZN(n3016) );
  AND2_X4 U3803 ( .A1(n3514), .A2(n4460), .ZN(n3099) );
  NAND2_X1 U3804 ( .A1(n3019), .A2(n3013), .ZN(n3014) );
  INV_X4 U3805 ( .A(n5774), .ZN(n5530) );
  OAI211_X1 U3806 ( .C1(n3099), .C2(INSTADDRPOINTER_REG_1__SCAN_IN), .A(n3014), 
        .B(n5530), .ZN(n3015) );
  NAND2_X1 U3807 ( .A1(n3016), .A2(n3015), .ZN(n3020) );
  INV_X2 U3808 ( .A(n3099), .ZN(n3113) );
  NAND2_X1 U3809 ( .A1(n3113), .A2(EBX_REG_0__SCAN_IN), .ZN(n3018) );
  INV_X1 U3810 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4904) );
  NAND2_X1 U3811 ( .A1(n5530), .A2(n4904), .ZN(n3017) );
  NOR2_X1 U3812 ( .A1(n4261), .A2(n4260), .ZN(n3022) );
  INV_X1 U3813 ( .A(n3020), .ZN(n3021) );
  NOR2_X2 U3814 ( .A1(n3022), .A2(n3021), .ZN(n4305) );
  NAND2_X1 U3815 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n4260), .ZN(n3023)
         );
  OAI21_X1 U3816 ( .B1(n3119), .B2(EBX_REG_2__SCAN_IN), .A(n3023), .ZN(n3026)
         );
  NAND2_X1 U3817 ( .A1(n3099), .A2(n4260), .ZN(n3065) );
  NAND2_X1 U3818 ( .A1(n3099), .A2(EBX_REG_2__SCAN_IN), .ZN(n3024) );
  NAND2_X1 U3819 ( .A1(n3065), .A2(n3024), .ZN(n3025) );
  NAND2_X1 U3820 ( .A1(n4305), .A2(n4306), .ZN(n4320) );
  NAND2_X1 U3821 ( .A1(n5530), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3028)
         );
  INV_X1 U3822 ( .A(EBX_REG_3__SCAN_IN), .ZN(n6635) );
  NAND2_X1 U3823 ( .A1(n4214), .A2(n6635), .ZN(n3027) );
  NAND3_X1 U3824 ( .A1(n3113), .A2(n3028), .A3(n3027), .ZN(n3030) );
  NAND2_X1 U3825 ( .A1(n3075), .A2(n6635), .ZN(n3029) );
  NAND2_X1 U3826 ( .A1(n3030), .A2(n3029), .ZN(n4321) );
  INV_X1 U3827 ( .A(EBX_REG_4__SCAN_IN), .ZN(n3032) );
  NAND2_X1 U3828 ( .A1(n3105), .A2(n3032), .ZN(n3035) );
  NAND2_X1 U3829 ( .A1(n4214), .A2(n3032), .ZN(n3033) );
  OAI211_X1 U3830 ( .C1(n3099), .C2(INSTADDRPOINTER_REG_4__SCAN_IN), .A(n3033), 
        .B(n5530), .ZN(n3034) );
  NAND2_X1 U3831 ( .A1(n3035), .A2(n3034), .ZN(n5386) );
  NAND2_X1 U3832 ( .A1(n3113), .A2(n5530), .ZN(n4220) );
  NAND2_X1 U3833 ( .A1(n5774), .A2(EBX_REG_5__SCAN_IN), .ZN(n3037) );
  INV_X1 U3834 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4328) );
  NAND2_X1 U3835 ( .A1(n3075), .A2(n4328), .ZN(n3036) );
  OAI211_X1 U3836 ( .C1(n4220), .C2(INSTADDRPOINTER_REG_5__SCAN_IN), .A(n3037), 
        .B(n3036), .ZN(n4325) );
  INV_X1 U3837 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6006) );
  NAND2_X1 U3838 ( .A1(n3105), .A2(n6006), .ZN(n3040) );
  NAND2_X1 U3839 ( .A1(n4214), .A2(n6006), .ZN(n3038) );
  OAI211_X1 U3840 ( .C1(n3099), .C2(INSTADDRPOINTER_REG_6__SCAN_IN), .A(n3038), 
        .B(n5530), .ZN(n3039) );
  NAND2_X1 U3841 ( .A1(n3040), .A2(n3039), .ZN(n4406) );
  NAND2_X1 U3842 ( .A1(n4405), .A2(n4406), .ZN(n4521) );
  INV_X1 U3843 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6231) );
  INV_X1 U3844 ( .A(EBX_REG_7__SCAN_IN), .ZN(n4851) );
  NAND2_X1 U3845 ( .A1(n4214), .A2(n4851), .ZN(n3041) );
  OAI211_X1 U3846 ( .C1(n5774), .C2(n6231), .A(n3113), .B(n3041), .ZN(n3042)
         );
  OAI21_X1 U3847 ( .B1(n3112), .B2(EBX_REG_7__SCAN_IN), .A(n3042), .ZN(n4522)
         );
  NOR2_X2 U3848 ( .A1(n4521), .A2(n4522), .ZN(n4520) );
  INV_X1 U3849 ( .A(EBX_REG_8__SCAN_IN), .ZN(n3043) );
  NAND2_X1 U3850 ( .A1(n3105), .A2(n3043), .ZN(n3046) );
  NAND2_X1 U3851 ( .A1(n4214), .A2(n3043), .ZN(n3044) );
  OAI211_X1 U3852 ( .C1(n3099), .C2(INSTADDRPOINTER_REG_8__SCAN_IN), .A(n3044), 
        .B(n5530), .ZN(n3045) );
  NAND2_X1 U3853 ( .A1(n3046), .A2(n3045), .ZN(n4617) );
  NAND2_X1 U3854 ( .A1(n4520), .A2(n4617), .ZN(n5992) );
  INV_X1 U3855 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6195) );
  INV_X1 U3856 ( .A(EBX_REG_9__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U3857 ( .A1(n4214), .A2(n6064), .ZN(n3047) );
  OAI211_X1 U3858 ( .C1(n5774), .C2(n6195), .A(n3113), .B(n3047), .ZN(n3048)
         );
  OAI21_X1 U3859 ( .B1(n3112), .B2(EBX_REG_9__SCAN_IN), .A(n3048), .ZN(n5993)
         );
  NAND2_X1 U3860 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n4260), .ZN(n3049) );
  OAI21_X1 U3861 ( .B1(n3119), .B2(EBX_REG_10__SCAN_IN), .A(n3049), .ZN(n3052)
         );
  NAND2_X1 U3862 ( .A1(n3099), .A2(EBX_REG_10__SCAN_IN), .ZN(n3050) );
  NAND2_X1 U3863 ( .A1(n3065), .A2(n3050), .ZN(n3051) );
  OR2_X1 U3864 ( .A1(n3052), .A2(n3051), .ZN(n4967) );
  NAND2_X1 U3865 ( .A1(n5991), .A2(n4967), .ZN(n5164) );
  INV_X1 U3866 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6574) );
  INV_X1 U3867 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6059) );
  NAND2_X1 U3868 ( .A1(n4214), .A2(n6059), .ZN(n3053) );
  OAI211_X1 U3869 ( .C1(n5774), .C2(n6574), .A(n3113), .B(n3053), .ZN(n3055)
         );
  NAND2_X1 U3870 ( .A1(n3075), .A2(n6059), .ZN(n3054) );
  NAND2_X1 U3871 ( .A1(n3055), .A2(n3054), .ZN(n5165) );
  NAND2_X1 U3872 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n4260), .ZN(n3056) );
  OAI21_X1 U3873 ( .B1(n3119), .B2(EBX_REG_12__SCAN_IN), .A(n3056), .ZN(n3059)
         );
  NAND2_X1 U3874 ( .A1(n3099), .A2(EBX_REG_12__SCAN_IN), .ZN(n3057) );
  NAND2_X1 U3875 ( .A1(n3065), .A2(n3057), .ZN(n3058) );
  OR2_X1 U3876 ( .A1(n3059), .A2(n3058), .ZN(n5114) );
  NAND2_X1 U3877 ( .A1(n5112), .A2(n5114), .ZN(n5908) );
  INV_X1 U3878 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5354) );
  INV_X1 U3879 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6556) );
  NAND2_X1 U3880 ( .A1(n4214), .A2(n6556), .ZN(n3060) );
  OAI211_X1 U3881 ( .C1(n5774), .C2(n5354), .A(n3113), .B(n3060), .ZN(n3062)
         );
  NAND2_X1 U3882 ( .A1(n3075), .A2(n6556), .ZN(n3061) );
  NAND2_X1 U3883 ( .A1(n3062), .A2(n3061), .ZN(n5909) );
  NAND2_X1 U3884 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n4260), .ZN(n3063) );
  OAI21_X1 U3885 ( .B1(n3119), .B2(EBX_REG_14__SCAN_IN), .A(n3063), .ZN(n3067)
         );
  NAND2_X1 U3886 ( .A1(n3099), .A2(EBX_REG_14__SCAN_IN), .ZN(n3064) );
  NAND2_X1 U3887 ( .A1(n3065), .A2(n3064), .ZN(n3066) );
  OR2_X1 U3888 ( .A1(n3067), .A2(n3066), .ZN(n5226) );
  INV_X1 U3889 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5906) );
  INV_X1 U3890 ( .A(EBX_REG_15__SCAN_IN), .ZN(n3068) );
  NAND2_X1 U3891 ( .A1(n4214), .A2(n3068), .ZN(n3069) );
  OAI211_X1 U3892 ( .C1(n5774), .C2(n5906), .A(n3113), .B(n3069), .ZN(n3070)
         );
  OAI21_X1 U3893 ( .B1(n3112), .B2(EBX_REG_15__SCAN_IN), .A(n3070), .ZN(n5243)
         );
  INV_X1 U3894 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5525) );
  NAND2_X1 U3895 ( .A1(n3105), .A2(n5525), .ZN(n3074) );
  INV_X1 U3896 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5663) );
  NAND2_X1 U3897 ( .A1(n3113), .A2(n5663), .ZN(n3072) );
  NAND2_X1 U3898 ( .A1(n4214), .A2(n5525), .ZN(n3071) );
  NAND3_X1 U3899 ( .A1(n3072), .A2(n5530), .A3(n3071), .ZN(n3073) );
  AND2_X1 U3900 ( .A1(n3074), .A2(n3073), .ZN(n5532) );
  INV_X1 U3901 ( .A(n5532), .ZN(n3081) );
  INV_X1 U3902 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6615) );
  NAND2_X1 U3903 ( .A1(n3075), .A2(n6615), .ZN(n3078) );
  NAND2_X1 U3904 ( .A1(n5530), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3076) );
  OAI211_X1 U3905 ( .C1(n4260), .C2(EBX_REG_17__SCAN_IN), .A(n3113), .B(n3076), 
        .ZN(n3077) );
  AND2_X1 U3906 ( .A1(n3078), .A2(n3077), .ZN(n5299) );
  NAND2_X1 U3907 ( .A1(n4260), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3080) );
  NAND2_X1 U3908 ( .A1(n3099), .A2(EBX_REG_16__SCAN_IN), .ZN(n3079) );
  OAI211_X1 U3909 ( .C1(n3119), .C2(EBX_REG_16__SCAN_IN), .A(n3080), .B(n3079), 
        .ZN(n5257) );
  AND2_X1 U3910 ( .A1(n5299), .A2(n5257), .ZN(n5298) );
  AND2_X1 U3911 ( .A1(n3081), .A2(n5298), .ZN(n5772) );
  OR2_X1 U3912 ( .A1(n4220), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3084)
         );
  INV_X1 U3913 ( .A(EBX_REG_20__SCAN_IN), .ZN(n3082) );
  NAND2_X1 U3914 ( .A1(n4214), .A2(n3082), .ZN(n3083) );
  AND2_X1 U3915 ( .A1(n3084), .A2(n3083), .ZN(n5778) );
  OR2_X1 U3916 ( .A1(n4220), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3085)
         );
  INV_X1 U3917 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5561) );
  NAND2_X1 U3918 ( .A1(n4214), .A2(n5561), .ZN(n5528) );
  NAND2_X1 U3919 ( .A1(n3085), .A2(n5528), .ZN(n5776) );
  NAND2_X1 U3920 ( .A1(n5774), .A2(EBX_REG_20__SCAN_IN), .ZN(n3087) );
  NAND2_X1 U3921 ( .A1(n5776), .A2(n5530), .ZN(n3086) );
  OAI211_X1 U3922 ( .C1(n5778), .C2(n5776), .A(n3087), .B(n3086), .ZN(n3088)
         );
  INV_X1 U3923 ( .A(n3088), .ZN(n3089) );
  AND2_X1 U3924 ( .A1(n5772), .A2(n3089), .ZN(n3090) );
  OR2_X1 U3925 ( .A1(n4220), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3092)
         );
  NAND2_X1 U3926 ( .A1(n5774), .A2(EBX_REG_21__SCAN_IN), .ZN(n3091) );
  OAI211_X1 U3927 ( .C1(n3112), .C2(EBX_REG_21__SCAN_IN), .A(n3092), .B(n3091), 
        .ZN(n3093) );
  INV_X1 U3928 ( .A(n3093), .ZN(n5544) );
  NAND2_X1 U3929 ( .A1(n5545), .A2(n5544), .ZN(n5547) );
  AOI22_X1 U3930 ( .A1(n3099), .A2(EBX_REG_22__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n4260), .ZN(n3096) );
  INV_X1 U3931 ( .A(EBX_REG_22__SCAN_IN), .ZN(n3094) );
  NAND2_X1 U3932 ( .A1(n3105), .A2(n3094), .ZN(n3095) );
  AND2_X1 U3933 ( .A1(n3096), .A2(n3095), .ZN(n5511) );
  OR2_X2 U3934 ( .A1(n5547), .A2(n5511), .ZN(n5513) );
  NAND2_X1 U3935 ( .A1(n5530), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3097) );
  OAI211_X1 U3936 ( .C1(n4260), .C2(EBX_REG_23__SCAN_IN), .A(n3113), .B(n3097), 
        .ZN(n3098) );
  OAI21_X1 U3937 ( .B1(n3112), .B2(EBX_REG_23__SCAN_IN), .A(n3098), .ZN(n5392)
         );
  NAND2_X1 U3938 ( .A1(n4260), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3101) );
  NAND2_X1 U3939 ( .A1(n3099), .A2(EBX_REG_24__SCAN_IN), .ZN(n3100) );
  OAI211_X1 U3940 ( .C1(n3119), .C2(EBX_REG_24__SCAN_IN), .A(n3101), .B(n3100), 
        .ZN(n5371) );
  NAND2_X1 U3941 ( .A1(n5394), .A2(n5371), .ZN(n5326) );
  OR2_X1 U3942 ( .A1(n4220), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3103)
         );
  NAND2_X1 U3943 ( .A1(n5774), .A2(EBX_REG_25__SCAN_IN), .ZN(n3102) );
  OAI211_X1 U3944 ( .C1(n3112), .C2(EBX_REG_25__SCAN_IN), .A(n3103), .B(n3102), 
        .ZN(n5327) );
  INV_X1 U3945 ( .A(EBX_REG_26__SCAN_IN), .ZN(n3104) );
  NAND2_X1 U3946 ( .A1(n3105), .A2(n3104), .ZN(n3109) );
  INV_X1 U3947 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3106) );
  NAND2_X1 U3948 ( .A1(n3113), .A2(n3106), .ZN(n3107) );
  OAI211_X1 U3949 ( .C1(EBX_REG_26__SCAN_IN), .C2(n4260), .A(n3107), .B(n5530), 
        .ZN(n3108) );
  AND2_X1 U3950 ( .A1(n3109), .A2(n3108), .ZN(n5492) );
  OR2_X2 U3951 ( .A1(n5491), .A2(n5492), .ZN(n5489) );
  OR2_X1 U3952 ( .A1(n4220), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3111)
         );
  NAND2_X1 U3953 ( .A1(n5774), .A2(EBX_REG_27__SCAN_IN), .ZN(n3110) );
  OAI211_X1 U3954 ( .C1(n3112), .C2(EBX_REG_27__SCAN_IN), .A(n3111), .B(n3110), 
        .ZN(n5477) );
  INV_X1 U3955 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5610) );
  NAND2_X1 U3956 ( .A1(n3113), .A2(n5610), .ZN(n3114) );
  OAI211_X1 U3957 ( .C1(EBX_REG_28__SCAN_IN), .C2(n4260), .A(n3114), .B(n5530), 
        .ZN(n3115) );
  OAI21_X1 U3958 ( .B1(n3119), .B2(EBX_REG_28__SCAN_IN), .A(n3115), .ZN(n5464)
         );
  INV_X1 U3959 ( .A(n4220), .ZN(n3117) );
  INV_X1 U3960 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5589) );
  NOR2_X1 U3961 ( .A1(n4260), .A2(EBX_REG_29__SCAN_IN), .ZN(n3116) );
  AOI21_X1 U3962 ( .B1(n3117), .B2(n5589), .A(n3116), .ZN(n5313) );
  NAND2_X1 U3963 ( .A1(n5414), .A2(n5530), .ZN(n3121) );
  NOR2_X1 U3964 ( .A1(n3119), .A2(EBX_REG_29__SCAN_IN), .ZN(n5314) );
  NAND2_X1 U3965 ( .A1(n5417), .A2(n5314), .ZN(n3120) );
  NAND2_X1 U3966 ( .A1(n3121), .A2(n3120), .ZN(n5319) );
  AND2_X1 U3967 ( .A1(n4260), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3122)
         );
  AOI21_X1 U3968 ( .B1(n4220), .B2(EBX_REG_30__SCAN_IN), .A(n3122), .ZN(n5415)
         );
  NAND2_X1 U3969 ( .A1(n5319), .A2(n5415), .ZN(n3124) );
  NOR2_X1 U3970 ( .A1(n5414), .A2(n5774), .ZN(n5420) );
  OAI22_X1 U3971 ( .A1(n4220), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4260), .ZN(n3125) );
  INV_X1 U3972 ( .A(READY_N), .ZN(n6441) );
  INV_X1 U3973 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6527) );
  NAND2_X1 U3974 ( .A1(n6441), .A2(n6527), .ZN(n3980) );
  AND2_X1 U3975 ( .A1(n4460), .A2(n3980), .ZN(n4846) );
  NAND2_X1 U3976 ( .A1(n3587), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3130)
         );
  NAND2_X1 U3977 ( .A1(n3592), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3129)
         );
  NAND2_X1 U3978 ( .A1(n3650), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3128) );
  NAND2_X1 U3979 ( .A1(n3922), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3127)
         );
  NAND2_X1 U3980 ( .A1(n3224), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3134)
         );
  NAND2_X1 U3981 ( .A1(n3921), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3133) );
  NAND2_X1 U3982 ( .A1(n2958), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3132) );
  NAND2_X1 U3983 ( .A1(n3583), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3131) );
  NAND2_X1 U3984 ( .A1(n3376), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3138) );
  NAND2_X1 U3985 ( .A1(n3273), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3137) );
  NAND2_X1 U3986 ( .A1(n3594), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3136)
         );
  NAND2_X1 U3987 ( .A1(n3940), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3135) );
  NAND2_X1 U3988 ( .A1(n3584), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3142) );
  NAND2_X1 U3989 ( .A1(n3585), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3141)
         );
  NAND2_X1 U3990 ( .A1(n3586), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3140) );
  NAND2_X1 U3991 ( .A1(n3274), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3139) );
  AOI22_X1 U3992 ( .A1(n3592), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3650), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3150) );
  AOI22_X1 U3993 ( .A1(n3224), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3149) );
  AOI22_X1 U3994 ( .A1(n3593), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3583), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3148) );
  AOI22_X1 U3995 ( .A1(n3587), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3237), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3147) );
  AND4_X2 U3996 ( .A1(n3150), .A2(n3149), .A3(n3148), .A4(n3147), .ZN(n3156)
         );
  AOI22_X1 U3997 ( .A1(n3782), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3594), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3154) );
  AOI22_X1 U3998 ( .A1(n3376), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3153) );
  AOI22_X1 U3999 ( .A1(n3586), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3274), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3152) );
  AOI22_X1 U4000 ( .A1(n3584), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3585), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3151) );
  NAND2_X1 U4001 ( .A1(n4237), .A2(n4474), .ZN(n4110) );
  NAND2_X1 U4002 ( .A1(n6691), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3173) );
  OAI21_X1 U4003 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6691), .A(n3173), 
        .ZN(n3161) );
  INV_X1 U4004 ( .A(n3161), .ZN(n3158) );
  AND2_X1 U4005 ( .A1(n4460), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3160) );
  INV_X1 U4006 ( .A(n3160), .ZN(n3157) );
  AOI21_X1 U4007 ( .B1(n4110), .B2(n3158), .A(n3157), .ZN(n3165) );
  INV_X2 U4008 ( .A(n4421), .ZN(n4171) );
  NAND2_X1 U4009 ( .A1(n4171), .A2(n4474), .ZN(n3159) );
  NAND2_X1 U4010 ( .A1(n4869), .A2(n3159), .ZN(n3178) );
  OR2_X1 U4011 ( .A1(n4460), .A2(n6529), .ZN(n3546) );
  AOI21_X1 U4012 ( .B1(n3737), .B2(n4421), .A(n5309), .ZN(n3166) );
  XNOR2_X1 U4013 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3175) );
  XNOR2_X1 U4014 ( .A(n3175), .B(n3173), .ZN(n3252) );
  NAND2_X1 U4015 ( .A1(n3252), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3167) );
  NAND2_X1 U4016 ( .A1(n3166), .A2(n3167), .ZN(n3164) );
  INV_X1 U4017 ( .A(n3737), .ZN(n3162) );
  AND2_X2 U4018 ( .A1(n3231), .A2(n4421), .ZN(n4058) );
  NAND2_X1 U4019 ( .A1(n3736), .A2(n4058), .ZN(n3197) );
  OAI21_X1 U4020 ( .B1(n3162), .B2(n3161), .A(n3197), .ZN(n3163) );
  OAI211_X1 U4021 ( .C1(n3165), .C2(n3178), .A(n3164), .B(n3163), .ZN(n3172)
         );
  INV_X1 U4022 ( .A(n3166), .ZN(n3170) );
  INV_X1 U4023 ( .A(n3252), .ZN(n3169) );
  NAND2_X1 U4024 ( .A1(n3197), .A2(n3167), .ZN(n3168) );
  OAI21_X1 U4025 ( .B1(n3170), .B2(n3169), .A(n3168), .ZN(n3171) );
  NAND2_X1 U4026 ( .A1(n3172), .A2(n3171), .ZN(n3181) );
  INV_X1 U4027 ( .A(n3173), .ZN(n3174) );
  NAND2_X1 U4028 ( .A1(n3175), .A2(n3174), .ZN(n3177) );
  NAND2_X1 U4029 ( .A1(n6393), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3176) );
  NAND2_X1 U4030 ( .A1(n3177), .A2(n3176), .ZN(n3186) );
  XNOR2_X1 U4031 ( .A(n3532), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3184)
         );
  XNOR2_X1 U4032 ( .A(n3186), .B(n3184), .ZN(n3253) );
  OAI211_X1 U4033 ( .C1(n3181), .C2(n3178), .A(n3253), .B(n3737), .ZN(n3183)
         );
  INV_X1 U4034 ( .A(n3736), .ZN(n3194) );
  INV_X1 U4035 ( .A(n3178), .ZN(n3179) );
  OAI21_X1 U4036 ( .B1(n3253), .B2(n3194), .A(n3179), .ZN(n3180) );
  NAND2_X1 U4037 ( .A1(n3181), .A2(n3180), .ZN(n3182) );
  NAND2_X1 U4038 ( .A1(n3183), .A2(n3182), .ZN(n3196) );
  INV_X1 U4039 ( .A(n3184), .ZN(n3185) );
  NAND2_X1 U4040 ( .A1(n3186), .A2(n3185), .ZN(n3188) );
  NAND2_X1 U4041 ( .A1(n6399), .A2(n6552), .ZN(n3187) );
  NAND2_X1 U4042 ( .A1(n3188), .A2(n3187), .ZN(n3193) );
  XNOR2_X1 U4043 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3191) );
  NAND2_X1 U4044 ( .A1(n3193), .A2(n3191), .ZN(n3190) );
  NAND2_X1 U4045 ( .A1(n4970), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3189) );
  NAND2_X1 U4046 ( .A1(n3190), .A2(n3189), .ZN(n3202) );
  INV_X1 U4047 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5924) );
  NAND2_X1 U4048 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n5924), .ZN(n3203) );
  OR2_X1 U4049 ( .A1(n3202), .A2(n3203), .ZN(n3254) );
  INV_X1 U4050 ( .A(n3191), .ZN(n3192) );
  XNOR2_X1 U4051 ( .A(n3193), .B(n3192), .ZN(n3251) );
  NAND2_X1 U4052 ( .A1(n3254), .A2(n3251), .ZN(n3198) );
  NAND2_X1 U4053 ( .A1(n3194), .A2(n3198), .ZN(n3195) );
  NAND2_X1 U4054 ( .A1(n3196), .A2(n3195), .ZN(n3200) );
  INV_X1 U4055 ( .A(n3197), .ZN(n3205) );
  AOI22_X1 U4056 ( .A1(n3205), .A2(n3198), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6529), .ZN(n3199) );
  NAND2_X1 U4057 ( .A1(n3200), .A2(n3199), .ZN(n3207) );
  INV_X1 U4058 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6412) );
  AND2_X1 U4059 ( .A1(n6412), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3201)
         );
  OR2_X1 U4060 ( .A1(n3202), .A2(n3201), .ZN(n3204) );
  NAND2_X1 U4061 ( .A1(n3205), .A2(n3250), .ZN(n3206) );
  NAND2_X1 U4062 ( .A1(n3737), .A2(n3250), .ZN(n3208) );
  INV_X1 U4063 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n4364) );
  AND2_X1 U4064 ( .A1(n4364), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3508) );
  NAND2_X1 U4065 ( .A1(n3508), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6424) );
  AOI22_X1 U4066 ( .A1(n3592), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3650), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3213) );
  AOI22_X1 U4067 ( .A1(n3224), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3212) );
  AOI22_X1 U4068 ( .A1(n2959), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3583), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3211) );
  AOI22_X1 U4069 ( .A1(n3587), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3237), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3210) );
  AOI22_X1 U4070 ( .A1(n3376), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3217) );
  AOI22_X1 U4071 ( .A1(n3584), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3585), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3216) );
  AOI22_X1 U4072 ( .A1(n3238), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3594), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3215) );
  AOI22_X1 U4073 ( .A1(n3586), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3274), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3214) );
  NAND2_X2 U4074 ( .A1(n3218), .A2(n2967), .ZN(n4455) );
  AOI22_X1 U4075 ( .A1(n3587), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3650), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3223) );
  AOI22_X1 U4076 ( .A1(n3592), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3222) );
  AOI22_X1 U4077 ( .A1(n2958), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3583), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3221) );
  AOI22_X1 U4078 ( .A1(n3584), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3586), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3220) );
  NAND4_X1 U4079 ( .A1(n3223), .A2(n3222), .A3(n3221), .A4(n3220), .ZN(n3230)
         );
  AOI22_X1 U4080 ( .A1(n3376), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3228) );
  AOI22_X1 U4081 ( .A1(n3224), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3237), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3227) );
  AOI22_X1 U4082 ( .A1(n3585), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3274), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3226) );
  AOI22_X1 U4083 ( .A1(n3782), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3594), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3225) );
  NAND4_X1 U4084 ( .A1(n3228), .A2(n3227), .A3(n3226), .A4(n3225), .ZN(n3229)
         );
  OR2_X2 U4085 ( .A1(n3230), .A2(n3229), .ZN(n5308) );
  NAND2_X1 U4086 ( .A1(n3485), .A2(n4237), .ZN(n3497) );
  NAND2_X2 U4087 ( .A1(n3518), .A2(n3231), .ZN(n4288) );
  INV_X1 U4088 ( .A(n4288), .ZN(n3232) );
  NOR2_X2 U4089 ( .A1(n3497), .A2(n3232), .ZN(n4147) );
  AOI22_X1 U4090 ( .A1(n3224), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3587), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3236) );
  AOI22_X1 U4091 ( .A1(n3584), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3376), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3235) );
  AOI22_X1 U4092 ( .A1(n2959), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3583), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3234) );
  AOI22_X1 U4093 ( .A1(n3585), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3274), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3233) );
  AOI22_X1 U4094 ( .A1(n3592), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3242) );
  BUF_X4 U4095 ( .A(n3237), .Z(n3950) );
  AOI22_X1 U4096 ( .A1(n3650), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3241) );
  BUF_X2 U4097 ( .A(n3238), .Z(n3916) );
  AOI22_X1 U4098 ( .A1(n3273), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3240) );
  AOI22_X1 U4099 ( .A1(n3586), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3594), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3239) );
  NOR2_X1 U4100 ( .A1(n4017), .A2(n4455), .ZN(n3243) );
  NAND2_X1 U4101 ( .A1(n4147), .A2(n3243), .ZN(n4166) );
  INV_X1 U4102 ( .A(n4166), .ZN(n3244) );
  NAND2_X1 U4103 ( .A1(n4288), .A2(n4465), .ZN(n3519) );
  NAND2_X1 U4104 ( .A1(n3518), .A2(n3245), .ZN(n3246) );
  NAND3_X1 U4105 ( .A1(n3248), .A2(n3246), .A3(n3481), .ZN(n3247) );
  NAND2_X1 U4106 ( .A1(n4282), .A2(n4212), .ZN(n3492) );
  NOR2_X1 U4107 ( .A1(n3492), .A2(n4460), .ZN(n3249) );
  NAND2_X1 U4108 ( .A1(n3494), .A2(n3249), .ZN(n3483) );
  INV_X1 U4109 ( .A(n3250), .ZN(n3256) );
  NAND4_X1 U4110 ( .A1(n3254), .A2(n3253), .A3(n3252), .A4(n3251), .ZN(n3255)
         );
  NAND2_X1 U4111 ( .A1(n3256), .A2(n3255), .ZN(n4186) );
  NOR2_X1 U4112 ( .A1(n4179), .A2(n4186), .ZN(n4136) );
  INV_X1 U4113 ( .A(n6424), .ZN(n4284) );
  NAND2_X1 U4114 ( .A1(n4136), .A2(n4284), .ZN(n4134) );
  AND2_X1 U4115 ( .A1(EBX_REG_31__SCAN_IN), .A2(n6523), .ZN(n3260) );
  AND2_X1 U4116 ( .A1(n4421), .A2(n3260), .ZN(n3257) );
  NAND2_X1 U4117 ( .A1(n4846), .A2(n3257), .ZN(n6024) );
  INV_X1 U4118 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6512) );
  NOR2_X1 U4119 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6535) );
  INV_X1 U4120 ( .A(n6535), .ZN(n6431) );
  NOR3_X1 U4121 ( .A1(n6529), .A2(n6512), .A3(n6431), .ZN(n6418) );
  NOR2_X1 U4122 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n4201) );
  NOR2_X1 U4123 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6434) );
  AND2_X1 U4124 ( .A1(n4201), .A2(n6434), .ZN(n6018) );
  INV_X1 U4125 ( .A(n6018), .ZN(n4889) );
  INV_X1 U4126 ( .A(n4889), .ZN(n6189) );
  NOR2_X1 U4127 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4364), .ZN(n6525) );
  NOR2_X1 U4128 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3878) );
  INV_X1 U4129 ( .A(n3878), .ZN(n3963) );
  INV_X1 U4130 ( .A(n3963), .ZN(n3968) );
  AND2_X1 U4131 ( .A1(n6525), .A2(n3968), .ZN(n6426) );
  OR2_X1 U4132 ( .A1(n6189), .A2(n6426), .ZN(n3258) );
  OR2_X1 U4133 ( .A1(n6418), .A2(n3258), .ZN(n3259) );
  INV_X1 U4134 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6440) );
  XNOR2_X1 U4135 ( .A(n6440), .B(STATE_REG_2__SCAN_IN), .ZN(n3480) );
  INV_X1 U4136 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6442) );
  NAND2_X1 U4137 ( .A1(n3480), .A2(n6442), .ZN(n6528) );
  OR2_X1 U4138 ( .A1(n6528), .A2(n3980), .ZN(n6417) );
  AND2_X1 U4139 ( .A1(n3496), .A2(n6417), .ZN(n4845) );
  AOI22_X1 U4140 ( .A1(n6008), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .B1(n3260), 
        .B2(n4845), .ZN(n3261) );
  OAI21_X1 U4141 ( .B1(n5701), .B2(n6024), .A(n3261), .ZN(n3262) );
  INV_X1 U4142 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n6569) );
  INV_X1 U4143 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3741) );
  NAND2_X1 U4144 ( .A1(n3776), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3807)
         );
  INV_X1 U4145 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3263) );
  INV_X1 U4146 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5983) );
  INV_X1 U4147 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5231) );
  INV_X1 U4148 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3861) );
  NAND2_X1 U4149 ( .A1(n3879), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3894)
         );
  INV_X1 U4150 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5294) );
  NAND2_X1 U4151 ( .A1(PHYADDRPOINTER_REG_23__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3265) );
  NAND2_X1 U4152 ( .A1(n3357), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3449)
         );
  INV_X1 U4153 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3448) );
  INV_X1 U4154 ( .A(n3451), .ZN(n3266) );
  NAND2_X1 U4155 ( .A1(n3266), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n3267)
         );
  INV_X1 U4156 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5465) );
  NAND2_X1 U4157 ( .A1(n3267), .A2(n5465), .ZN(n3268) );
  NAND2_X1 U4158 ( .A1(n3476), .A2(n3268), .ZN(n5613) );
  AOI22_X1 U4159 ( .A1(n3938), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3939), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3272) );
  AOI22_X1 U4160 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n3915), .B1(n2957), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3271) );
  AOI22_X1 U4161 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n3942), .B1(n3948), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3270) );
  AOI22_X1 U4162 ( .A1(n3376), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3952), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3269) );
  NAND4_X1 U4163 ( .A1(n3272), .A2(n3271), .A3(n3270), .A4(n3269), .ZN(n3280)
         );
  AOI22_X1 U4164 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n3551), .B1(n3951), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3278) );
  AOI22_X1 U4165 ( .A1(n3937), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3277) );
  AOI22_X1 U4166 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n3947), .B1(n3940), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3276) );
  AOI22_X1 U4167 ( .A1(n3949), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3941), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3275) );
  NAND4_X1 U4168 ( .A1(n3278), .A2(n3277), .A3(n3276), .A4(n3275), .ZN(n3279)
         );
  NOR2_X1 U4169 ( .A1(n3280), .A2(n3279), .ZN(n3346) );
  AOI22_X1 U4170 ( .A1(n3939), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3284) );
  AOI22_X1 U4171 ( .A1(n3915), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3283) );
  AOI22_X1 U4172 ( .A1(n2958), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3282) );
  AOI22_X1 U4173 ( .A1(n3938), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3922), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3281) );
  NAND4_X1 U4174 ( .A1(n3284), .A2(n3283), .A3(n3282), .A4(n3281), .ZN(n3290)
         );
  AOI22_X1 U4175 ( .A1(n3769), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3947), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3288) );
  AOI22_X1 U4176 ( .A1(n3949), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3287) );
  AOI22_X1 U4177 ( .A1(n3782), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3952), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3286) );
  AOI22_X1 U4178 ( .A1(n3948), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3941), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3285) );
  NAND4_X1 U4179 ( .A1(n3288), .A2(n3287), .A3(n3286), .A4(n3285), .ZN(n3289)
         );
  NOR2_X1 U4180 ( .A1(n3290), .A2(n3289), .ZN(n3354) );
  AOI22_X1 U4181 ( .A1(n3951), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3551), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3294) );
  AOI22_X1 U4182 ( .A1(n3949), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3948), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3293) );
  AOI22_X1 U4183 ( .A1(n3947), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3292) );
  AOI22_X1 U4184 ( .A1(n3938), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3291) );
  NAND4_X1 U4185 ( .A1(n3294), .A2(n3293), .A3(n3292), .A4(n3291), .ZN(n3300)
         );
  AOI22_X1 U4186 ( .A1(n3939), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3298) );
  AOI22_X1 U4187 ( .A1(n3915), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3297) );
  AOI22_X1 U4188 ( .A1(n3376), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3952), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3296) );
  AOI22_X1 U4189 ( .A1(n3942), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3941), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3295) );
  NAND4_X1 U4190 ( .A1(n3298), .A2(n3297), .A3(n3296), .A4(n3295), .ZN(n3299)
         );
  NOR2_X1 U4191 ( .A1(n3300), .A2(n3299), .ZN(n3369) );
  AOI22_X1 U4192 ( .A1(n3915), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3304) );
  AOI22_X1 U4193 ( .A1(n3769), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3303) );
  AOI22_X1 U4194 ( .A1(n3938), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3302) );
  AOI22_X1 U4195 ( .A1(n3949), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3941), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3301) );
  NAND4_X1 U4196 ( .A1(n3304), .A2(n3303), .A3(n3302), .A4(n3301), .ZN(n3310)
         );
  AOI22_X1 U4197 ( .A1(n3939), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3308) );
  AOI22_X1 U4198 ( .A1(n3551), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3947), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3307) );
  AOI22_X1 U4199 ( .A1(n3942), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3948), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3306) );
  AOI22_X1 U4200 ( .A1(n3940), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3952), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3305) );
  NAND4_X1 U4201 ( .A1(n3308), .A2(n3307), .A3(n3306), .A4(n3305), .ZN(n3309)
         );
  NOR2_X1 U4202 ( .A1(n3310), .A2(n3309), .ZN(n3370) );
  NOR2_X1 U4203 ( .A1(n3369), .A2(n3370), .ZN(n3365) );
  AOI22_X1 U4204 ( .A1(n3939), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3314) );
  AOI22_X1 U4205 ( .A1(n3915), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3951), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3313) );
  AOI22_X1 U4206 ( .A1(n3551), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3312) );
  AOI22_X1 U4207 ( .A1(n3938), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3311) );
  NAND4_X1 U4208 ( .A1(n3314), .A2(n3313), .A3(n3312), .A4(n3311), .ZN(n3320)
         );
  AOI22_X1 U4209 ( .A1(n3769), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3947), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3318) );
  AOI22_X1 U4210 ( .A1(n3949), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3317) );
  AOI22_X1 U4211 ( .A1(n3940), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3952), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3316) );
  AOI22_X1 U4212 ( .A1(n3948), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3941), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3315) );
  NAND4_X1 U4213 ( .A1(n3318), .A2(n3317), .A3(n3316), .A4(n3315), .ZN(n3319)
         );
  OR2_X1 U4214 ( .A1(n3320), .A2(n3319), .ZN(n3364) );
  NAND2_X1 U4215 ( .A1(n3365), .A2(n3364), .ZN(n3353) );
  NOR2_X1 U4216 ( .A1(n3354), .A2(n3353), .ZN(n3453) );
  AOI22_X1 U4217 ( .A1(n3939), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3324) );
  AOI22_X1 U4218 ( .A1(n3915), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3951), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3323) );
  AOI22_X1 U4219 ( .A1(n2959), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3322) );
  AOI22_X1 U4220 ( .A1(n3938), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3321) );
  NAND4_X1 U4221 ( .A1(n3324), .A2(n3323), .A3(n3322), .A4(n3321), .ZN(n3330)
         );
  AOI22_X1 U4222 ( .A1(n3376), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3947), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3328) );
  AOI22_X1 U4223 ( .A1(n3949), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3327) );
  AOI22_X1 U4224 ( .A1(n3940), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3952), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3326) );
  AOI22_X1 U4225 ( .A1(n3948), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3941), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3325) );
  NAND4_X1 U4226 ( .A1(n3328), .A2(n3327), .A3(n3326), .A4(n3325), .ZN(n3329)
         );
  OR2_X1 U4227 ( .A1(n3330), .A2(n3329), .ZN(n3452) );
  NAND2_X1 U4228 ( .A1(n3453), .A2(n3452), .ZN(n3347) );
  NOR2_X1 U4229 ( .A1(n3346), .A2(n3347), .ZN(n3461) );
  AOI22_X1 U4230 ( .A1(n3939), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3650), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3334) );
  AOI22_X1 U4231 ( .A1(n3915), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3951), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3333) );
  AOI22_X1 U4232 ( .A1(n2958), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3332) );
  AOI22_X1 U4233 ( .A1(n3938), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3331) );
  NAND4_X1 U4234 ( .A1(n3334), .A2(n3333), .A3(n3332), .A4(n3331), .ZN(n3340)
         );
  AOI22_X1 U4235 ( .A1(n3376), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3947), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3338) );
  AOI22_X1 U4236 ( .A1(n3949), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3337) );
  AOI22_X1 U4237 ( .A1(n3940), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3952), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3336) );
  AOI22_X1 U4238 ( .A1(n3948), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3941), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3335) );
  NAND4_X1 U4239 ( .A1(n3338), .A2(n3337), .A3(n3336), .A4(n3335), .ZN(n3339)
         );
  OR2_X1 U4240 ( .A1(n3340), .A2(n3339), .ZN(n3460) );
  XNOR2_X1 U4241 ( .A(n3461), .B(n3460), .ZN(n3344) );
  NAND2_X1 U4242 ( .A1(n4479), .A2(n5308), .ZN(n3341) );
  OR2_X1 U4243 ( .A1(n4288), .A2(n3341), .ZN(n4173) );
  INV_X1 U4244 ( .A(n4173), .ZN(n4197) );
  NAND2_X1 U4245 ( .A1(n4197), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3966) );
  INV_X2 U4246 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6522) );
  AOI21_X1 U4247 ( .B1(PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6522), .A(n3968), 
        .ZN(n3343) );
  INV_X2 U4248 ( .A(n3930), .ZN(n3972) );
  NAND2_X1 U4249 ( .A1(n3972), .A2(EAX_REG_28__SCAN_IN), .ZN(n3342) );
  OAI211_X1 U4250 ( .C1(n3344), .C2(n3966), .A(n3343), .B(n3342), .ZN(n3345)
         );
  OAI21_X1 U4251 ( .B1(n3963), .B2(n5613), .A(n3345), .ZN(n5462) );
  XOR2_X1 U4252 ( .A(n3347), .B(n3346), .Z(n3348) );
  INV_X1 U4253 ( .A(n3966), .ZN(n3933) );
  NAND2_X1 U4254 ( .A1(n3348), .A2(n3933), .ZN(n3352) );
  INV_X1 U4255 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n3349) );
  NOR2_X1 U4256 ( .A1(n3349), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3350) );
  AOI211_X1 U4257 ( .C1(n3972), .C2(EAX_REG_27__SCAN_IN), .A(n3968), .B(n3350), 
        .ZN(n3351) );
  XNOR2_X1 U4258 ( .A(n3451), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5476)
         );
  AOI22_X1 U4259 ( .A1(n3352), .A2(n3351), .B1(n3968), .B2(n5476), .ZN(n5474)
         );
  XOR2_X1 U4260 ( .A(n3354), .B(n3353), .Z(n3355) );
  NAND2_X1 U4261 ( .A1(n3355), .A2(n3933), .ZN(n3361) );
  INV_X1 U4262 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n6659) );
  NOR2_X1 U4263 ( .A1(n6659), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3356) );
  AOI211_X1 U4264 ( .C1(n3972), .C2(EAX_REG_25__SCAN_IN), .A(n3878), .B(n3356), 
        .ZN(n3360) );
  INV_X1 U4265 ( .A(n3357), .ZN(n3358) );
  NAND2_X1 U4266 ( .A1(n3358), .A2(n6659), .ZN(n3359) );
  AND2_X1 U4267 ( .A1(n3449), .A2(n3359), .ZN(n5637) );
  AOI22_X1 U4268 ( .A1(n3361), .A2(n3360), .B1(n3968), .B2(n5637), .ZN(n5323)
         );
  INV_X1 U4269 ( .A(n3392), .ZN(n3362) );
  NAND2_X1 U4270 ( .A1(n3362), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3363)
         );
  XNOR2_X1 U4271 ( .A(n3363), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5505)
         );
  INV_X1 U4272 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5502) );
  NAND2_X1 U4273 ( .A1(n6522), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3828) );
  OAI22_X1 U4274 ( .A1(n5505), .A2(n3963), .B1(n5502), .B2(n3828), .ZN(n3368)
         );
  XNOR2_X1 U4275 ( .A(n3365), .B(n3364), .ZN(n3366) );
  NOR2_X1 U4276 ( .A1(n3366), .A2(n3966), .ZN(n3367) );
  AOI211_X1 U4277 ( .C1(n3972), .C2(EAX_REG_24__SCAN_IN), .A(n3368), .B(n3367), 
        .ZN(n5379) );
  INV_X1 U4278 ( .A(n5379), .ZN(n3447) );
  XNOR2_X1 U4279 ( .A(n3392), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5844)
         );
  XOR2_X1 U4280 ( .A(n3370), .B(n3369), .Z(n3374) );
  INV_X1 U4281 ( .A(EAX_REG_23__SCAN_IN), .ZN(n3372) );
  NAND2_X1 U4282 ( .A1(n6522), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3371)
         );
  OAI211_X1 U4283 ( .C1(n3930), .C2(n3372), .A(n3963), .B(n3371), .ZN(n3373)
         );
  AOI21_X1 U4284 ( .B1(n3933), .B2(n3374), .A(n3373), .ZN(n3375) );
  AOI21_X1 U4285 ( .B1(n3968), .B2(n5844), .A(n3375), .ZN(n4118) );
  AOI22_X1 U4286 ( .A1(n3938), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3380) );
  AOI22_X1 U4287 ( .A1(n3939), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3551), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3379) );
  AOI22_X1 U4289 ( .A1(n3769), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3947), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3378) );
  AOI22_X1 U4290 ( .A1(n3949), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3941), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3377) );
  NAND4_X1 U4291 ( .A1(n3380), .A2(n3379), .A3(n3378), .A4(n3377), .ZN(n3387)
         );
  AOI22_X1 U4292 ( .A1(n3915), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3385) );
  AOI22_X1 U4293 ( .A1(n3942), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3948), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3384) );
  AOI22_X1 U4294 ( .A1(n3951), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3383) );
  AOI22_X1 U4295 ( .A1(n3782), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3952), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3382) );
  NAND4_X1 U4296 ( .A1(n3385), .A2(n3384), .A3(n3383), .A4(n3382), .ZN(n3386)
         );
  NOR2_X1 U4297 ( .A1(n3387), .A2(n3386), .ZN(n3391) );
  NAND2_X1 U4298 ( .A1(n6522), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3388)
         );
  NAND2_X1 U4299 ( .A1(n3963), .A2(n3388), .ZN(n3389) );
  AOI21_X1 U4300 ( .B1(n3972), .B2(EAX_REG_22__SCAN_IN), .A(n3389), .ZN(n3390)
         );
  OAI21_X1 U4301 ( .B1(n3966), .B2(n3391), .A(n3390), .ZN(n3395) );
  OAI21_X1 U4302 ( .B1(n3393), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n3392), 
        .ZN(n5515) );
  OR2_X1 U4303 ( .A1(n5515), .A2(n3963), .ZN(n3394) );
  AND2_X1 U4304 ( .A1(n3395), .A2(n3394), .ZN(n5343) );
  INV_X1 U4305 ( .A(n5343), .ZN(n3429) );
  AOI22_X1 U4306 ( .A1(n3951), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3399) );
  AOI22_X1 U4307 ( .A1(n3551), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3922), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3398) );
  AOI22_X1 U4308 ( .A1(n3948), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3397) );
  AOI22_X1 U4309 ( .A1(n3939), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3941), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3396) );
  NAND4_X1 U4310 ( .A1(n3399), .A2(n3398), .A3(n3397), .A4(n3396), .ZN(n3407)
         );
  NAND2_X1 U4311 ( .A1(n3949), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3401)
         );
  NAND2_X1 U4312 ( .A1(n3937), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3400) );
  AND3_X1 U4313 ( .A1(n3401), .A2(n3400), .A3(n3963), .ZN(n3405) );
  AOI22_X1 U4314 ( .A1(n3915), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3404) );
  AOI22_X1 U4315 ( .A1(n3938), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3403) );
  AOI22_X1 U4316 ( .A1(n3947), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3952), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3402) );
  NAND4_X1 U4317 ( .A1(n3405), .A2(n3404), .A3(n3403), .A4(n3402), .ZN(n3406)
         );
  NAND2_X1 U4318 ( .A1(n3966), .A2(n3963), .ZN(n3910) );
  OAI21_X1 U4319 ( .B1(n3407), .B2(n3406), .A(n3910), .ZN(n3409) );
  AOI22_X1 U4320 ( .A1(n3972), .A2(EAX_REG_21__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6522), .ZN(n3408) );
  NAND2_X1 U4321 ( .A1(n3409), .A2(n3408), .ZN(n3411) );
  XNOR2_X1 U4322 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .B(n3413), .ZN(n5859)
         );
  NAND2_X1 U4323 ( .A1(n5859), .A2(n3878), .ZN(n3410) );
  NAND2_X1 U4324 ( .A1(n3411), .A2(n3410), .ZN(n5543) );
  OR2_X1 U4325 ( .A1(n3412), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3414)
         );
  NAND2_X1 U4326 ( .A1(n3414), .A2(n3413), .ZN(n5869) );
  AOI22_X1 U4327 ( .A1(n3938), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3418) );
  AOI22_X1 U4328 ( .A1(n3939), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3417) );
  AOI22_X1 U4329 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n3949), .B1(n3948), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3416) );
  AOI22_X1 U4330 ( .A1(n3947), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3952), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3415) );
  NAND4_X1 U4331 ( .A1(n3418), .A2(n3417), .A3(n3416), .A4(n3415), .ZN(n3424)
         );
  AOI22_X1 U4332 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n3551), .B1(n2957), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3422) );
  AOI22_X1 U4333 ( .A1(n3915), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3922), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3421) );
  AOI22_X1 U4334 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n3769), .B1(n3916), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3420) );
  AOI22_X1 U4335 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n3942), .B1(n3941), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3419) );
  NAND4_X1 U4336 ( .A1(n3422), .A2(n3421), .A3(n3420), .A4(n3419), .ZN(n3423)
         );
  NOR2_X1 U4337 ( .A1(n3424), .A2(n3423), .ZN(n3427) );
  OAI21_X1 U4338 ( .B1(PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6527), .A(n6522), 
        .ZN(n3426) );
  NAND2_X1 U4339 ( .A1(n3972), .A2(EAX_REG_20__SCAN_IN), .ZN(n3425) );
  OAI211_X1 U4340 ( .C1(n3966), .C2(n3427), .A(n3426), .B(n3425), .ZN(n3428)
         );
  OAI21_X1 U4341 ( .B1(n5869), .B2(n3963), .A(n3428), .ZN(n5656) );
  OR2_X1 U4342 ( .A1(n5543), .A2(n5656), .ZN(n5342) );
  NOR2_X1 U4343 ( .A1(n3429), .A2(n5342), .ZN(n4114) );
  AND2_X1 U4344 ( .A1(n4118), .A2(n4114), .ZN(n3446) );
  INV_X1 U4345 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5666) );
  XNOR2_X1 U4346 ( .A(n3914), .B(n5666), .ZN(n5670) );
  AOI22_X1 U4347 ( .A1(n3938), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3435) );
  AOI22_X1 U4348 ( .A1(n3769), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3434) );
  NAND2_X1 U4349 ( .A1(n3939), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3431) );
  NAND2_X1 U4350 ( .A1(n3948), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3430) );
  AND3_X1 U4351 ( .A1(n3431), .A2(n3430), .A3(n3963), .ZN(n3433) );
  AOI22_X1 U4352 ( .A1(n3551), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3432) );
  NAND4_X1 U4353 ( .A1(n3435), .A2(n3434), .A3(n3433), .A4(n3432), .ZN(n3441)
         );
  AOI22_X1 U4354 ( .A1(n3915), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3439) );
  AOI22_X1 U4355 ( .A1(n3947), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3941), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3438) );
  AOI22_X1 U4356 ( .A1(n3949), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3922), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3437) );
  AOI22_X1 U4357 ( .A1(n3951), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3952), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3436) );
  NAND4_X1 U4358 ( .A1(n3439), .A2(n3438), .A3(n3437), .A4(n3436), .ZN(n3440)
         );
  OR2_X1 U4359 ( .A1(n3441), .A2(n3440), .ZN(n3444) );
  INV_X1 U4360 ( .A(EAX_REG_19__SCAN_IN), .ZN(n3442) );
  OAI22_X1 U4361 ( .A1(n3930), .A2(n3442), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5666), .ZN(n3443) );
  AOI21_X1 U4362 ( .B1(n3910), .B2(n3444), .A(n3443), .ZN(n3445) );
  AOI21_X1 U4363 ( .B1(n5670), .B2(n3878), .A(n3445), .ZN(n5522) );
  AND2_X1 U4364 ( .A1(n3446), .A2(n5522), .ZN(n4117) );
  AND2_X1 U4365 ( .A1(n3447), .A2(n4117), .ZN(n5321) );
  AND2_X1 U4366 ( .A1(n5323), .A2(n5321), .ZN(n5322) );
  NAND2_X1 U4367 ( .A1(n3449), .A2(n3448), .ZN(n3450) );
  NAND2_X1 U4368 ( .A1(n3451), .A2(n3450), .ZN(n5630) );
  XNOR2_X1 U4369 ( .A(n3453), .B(n3452), .ZN(n3456) );
  AOI21_X1 U4370 ( .B1(PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n6522), .A(n3878), 
        .ZN(n3455) );
  NAND2_X1 U4371 ( .A1(n3972), .A2(EAX_REG_26__SCAN_IN), .ZN(n3454) );
  OAI211_X1 U4372 ( .C1(n3456), .C2(n3966), .A(n3455), .B(n3454), .ZN(n3457)
         );
  OAI21_X1 U4373 ( .B1(n3963), .B2(n5630), .A(n3457), .ZN(n5488) );
  INV_X1 U4374 ( .A(n5488), .ZN(n3458) );
  AND2_X1 U4375 ( .A1(n5322), .A2(n3458), .ZN(n5472) );
  AND2_X1 U4376 ( .A1(n5474), .A2(n5472), .ZN(n5460) );
  INV_X1 U4377 ( .A(n5460), .ZN(n3459) );
  NOR2_X1 U4378 ( .A1(n5462), .A2(n3459), .ZN(n5305) );
  NAND2_X1 U4379 ( .A1(n3461), .A2(n3460), .ZN(n3959) );
  AOI22_X1 U4380 ( .A1(n3915), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3947), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3465) );
  AOI22_X1 U4381 ( .A1(n3949), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3376), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3464) );
  AOI22_X1 U4382 ( .A1(n3951), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3463) );
  AOI22_X1 U4383 ( .A1(n3942), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3941), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3462) );
  NAND4_X1 U4384 ( .A1(n3465), .A2(n3464), .A3(n3463), .A4(n3462), .ZN(n3471)
         );
  AOI22_X1 U4385 ( .A1(n3938), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3650), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3469) );
  AOI22_X1 U4386 ( .A1(n3939), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3551), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3468) );
  AOI22_X1 U4387 ( .A1(n2957), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3467) );
  AOI22_X1 U4388 ( .A1(n3948), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3952), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3466) );
  NAND4_X1 U4389 ( .A1(n3469), .A2(n3468), .A3(n3467), .A4(n3466), .ZN(n3470)
         );
  NOR2_X1 U4390 ( .A1(n3471), .A2(n3470), .ZN(n3960) );
  XOR2_X1 U4391 ( .A(n3959), .B(n3960), .Z(n3472) );
  NAND2_X1 U4392 ( .A1(n3472), .A2(n3933), .ZN(n3479) );
  INV_X1 U4393 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n3475) );
  AOI21_X1 U4394 ( .B1(n3475), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3473) );
  AOI21_X1 U4395 ( .B1(n3972), .B2(EAX_REG_29__SCAN_IN), .A(n3473), .ZN(n3478)
         );
  NAND2_X1 U4396 ( .A1(n3476), .A2(n3475), .ZN(n3477) );
  AND2_X1 U4397 ( .A1(n3975), .A2(n3477), .ZN(n5453) );
  AOI22_X1 U4398 ( .A1(n3479), .A2(n3478), .B1(n3968), .B2(n5453), .ZN(n5306)
         );
  AND2_X1 U4399 ( .A1(n5305), .A2(n5306), .ZN(n3936) );
  NAND2_X1 U4400 ( .A1(n3514), .A2(n3481), .ZN(n3517) );
  NOR2_X1 U4401 ( .A1(n3517), .A2(n4474), .ZN(n3482) );
  AND2_X2 U4402 ( .A1(n4156), .A2(n3482), .ZN(n4283) );
  AND2_X1 U4403 ( .A1(n5308), .A2(n4455), .ZN(n4141) );
  OR2_X2 U4404 ( .A1(n3483), .A2(n4421), .ZN(n5920) );
  NAND2_X1 U4405 ( .A1(n3484), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3506) );
  NAND2_X1 U4406 ( .A1(n4288), .A2(n4460), .ZN(n4145) );
  OAI21_X1 U4407 ( .B1(n4479), .B2(n4288), .A(n3485), .ZN(n3486) );
  INV_X1 U4408 ( .A(n3487), .ZN(n3488) );
  AOI21_X1 U4409 ( .B1(n5309), .B2(n3488), .A(n4017), .ZN(n3489) );
  OAI211_X1 U4410 ( .C1(n4237), .C2(n4145), .A(n4108), .B(n3489), .ZN(n3490)
         );
  INV_X1 U4411 ( .A(n3490), .ZN(n3499) );
  NAND2_X1 U4412 ( .A1(n3494), .A2(n3493), .ZN(n3495) );
  NAND2_X1 U4413 ( .A1(n3495), .A2(n4130), .ZN(n3511) );
  NAND2_X1 U4414 ( .A1(n3497), .A2(n3496), .ZN(n3498) );
  NAND2_X1 U4415 ( .A1(n4153), .A2(n4465), .ZN(n4168) );
  NAND3_X1 U4416 ( .A1(n3499), .A2(n3511), .A3(n3523), .ZN(n3500) );
  NAND2_X1 U4417 ( .A1(n4201), .A2(n6529), .ZN(n4120) );
  INV_X1 U4418 ( .A(n4120), .ZN(n3647) );
  XNOR2_X1 U4419 ( .A(n6393), .B(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5177)
         );
  NAND2_X1 U4420 ( .A1(n3647), .A2(n5177), .ZN(n3502) );
  INV_X1 U4421 ( .A(n3508), .ZN(n3646) );
  NAND2_X1 U4422 ( .A1(n3646), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3501) );
  NAND2_X1 U4423 ( .A1(n3502), .A2(n3501), .ZN(n3504) );
  NAND2_X2 U4424 ( .A1(n3506), .A2(n3503), .ZN(n3525) );
  NOR2_X1 U4425 ( .A1(n3504), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3505)
         );
  OR2_X2 U4426 ( .A1(n3506), .A2(n3505), .ZN(n3507) );
  NAND2_X2 U4427 ( .A1(n3525), .A2(n3507), .ZN(n3550) );
  MUX2_X1 U4428 ( .A(n4120), .B(n3508), .S(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), 
        .Z(n3509) );
  OR2_X1 U4429 ( .A1(n3511), .A2(n4153), .ZN(n3513) );
  NAND2_X1 U4430 ( .A1(n4450), .A2(n4460), .ZN(n3512) );
  NAND2_X1 U4431 ( .A1(n3513), .A2(n3512), .ZN(n4150) );
  AOI21_X1 U4432 ( .B1(n4288), .B2(n4479), .A(n3514), .ZN(n3515) );
  NAND2_X1 U4433 ( .A1(n4108), .A2(n3515), .ZN(n3516) );
  NAND2_X1 U4434 ( .A1(n3516), .A2(n4421), .ZN(n3522) );
  INV_X1 U4435 ( .A(n3517), .ZN(n4216) );
  AND2_X1 U4436 ( .A1(n4216), .A2(n4130), .ZN(n4151) );
  NAND2_X1 U4437 ( .A1(n4201), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6425) );
  AOI21_X1 U4438 ( .B1(n4151), .B2(n4241), .A(n6425), .ZN(n3521) );
  NAND2_X1 U4439 ( .A1(n3519), .A2(n3496), .ZN(n3520) );
  NAND4_X1 U4440 ( .A1(n3523), .A2(n3522), .A3(n3521), .A4(n3520), .ZN(n3524)
         );
  OR2_X2 U4441 ( .A1(n3550), .A2(n3549), .ZN(n3526) );
  NAND2_X2 U4442 ( .A1(n3526), .A2(n3525), .ZN(n3641) );
  AND2_X1 U4443 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3528) );
  NAND2_X1 U4444 ( .A1(n3528), .A2(n6399), .ZN(n4594) );
  INV_X1 U4445 ( .A(n3528), .ZN(n3529) );
  NAND2_X1 U4446 ( .A1(n3529), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3530) );
  NAND2_X1 U4447 ( .A1(n4594), .A2(n3530), .ZN(n4447) );
  AOI22_X1 U4448 ( .A1(n3647), .A2(n4447), .B1(n3646), .B2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3531) );
  NAND2_X1 U4449 ( .A1(n4345), .A2(n6529), .ZN(n3545) );
  INV_X1 U4450 ( .A(n3606), .ZN(n3610) );
  INV_X1 U4451 ( .A(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n6683) );
  AOI22_X1 U4452 ( .A1(n3939), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3650), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3537) );
  AOI22_X1 U4453 ( .A1(n3915), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3536) );
  AOI22_X1 U4454 ( .A1(n3551), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3583), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3535) );
  AOI22_X1 U4455 ( .A1(n3938), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3534) );
  NAND4_X1 U4456 ( .A1(n3537), .A2(n3536), .A3(n3535), .A4(n3534), .ZN(n3543)
         );
  AOI22_X1 U4457 ( .A1(n3769), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3947), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3541) );
  AOI22_X1 U4458 ( .A1(n3949), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3540) );
  AOI22_X1 U4459 ( .A1(n3782), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3952), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3539) );
  AOI22_X1 U4460 ( .A1(n3948), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3941), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3538) );
  NAND4_X1 U4461 ( .A1(n3541), .A2(n3540), .A3(n3539), .A4(n3538), .ZN(n3542)
         );
  OR2_X1 U4462 ( .A1(n3543), .A2(n3542), .ZN(n3997) );
  NAND2_X1 U4463 ( .A1(n3610), .A2(n3997), .ZN(n3544) );
  INV_X1 U4464 ( .A(n3546), .ZN(n6533) );
  AOI22_X1 U4465 ( .A1(n3736), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n6533), 
        .B2(n3997), .ZN(n3547) );
  XNOR2_X2 U4466 ( .A(n3548), .B(n3547), .ZN(n3682) );
  XNOR2_X2 U4467 ( .A(n3550), .B(n3549), .ZN(n4495) );
  INV_X1 U4468 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n6632) );
  AOI22_X1 U4469 ( .A1(n3939), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3650), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3555) );
  AOI22_X1 U4470 ( .A1(n3915), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3554) );
  CLKBUF_X1 U4471 ( .A(n2959), .Z(n3551) );
  AOI22_X1 U4472 ( .A1(n3551), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3583), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3553) );
  AOI22_X1 U4473 ( .A1(n3938), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3552) );
  NAND4_X1 U4474 ( .A1(n3555), .A2(n3554), .A3(n3553), .A4(n3552), .ZN(n3561)
         );
  AOI22_X1 U4475 ( .A1(n3769), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3947), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3559) );
  AOI22_X1 U4476 ( .A1(n3949), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3558) );
  AOI22_X1 U4477 ( .A1(n3782), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3952), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3557) );
  AOI22_X1 U4478 ( .A1(n3948), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3941), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3556) );
  NAND4_X1 U4479 ( .A1(n3559), .A2(n3558), .A3(n3557), .A4(n3556), .ZN(n3560)
         );
  NAND2_X1 U4480 ( .A1(n3610), .A2(n4016), .ZN(n3562) );
  AOI22_X1 U4481 ( .A1(n3938), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3939), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3567) );
  AOI22_X1 U4482 ( .A1(n3551), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3583), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3566) );
  AOI22_X1 U4483 ( .A1(n3949), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3948), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3565) );
  AOI22_X1 U4484 ( .A1(n3376), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3952), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3564) );
  NAND4_X1 U4485 ( .A1(n3567), .A2(n3566), .A3(n3565), .A4(n3564), .ZN(n3573)
         );
  AOI22_X1 U4486 ( .A1(n3915), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3571) );
  AOI22_X1 U4487 ( .A1(n3937), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3570) );
  AOI22_X1 U4488 ( .A1(n3947), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3569) );
  AOI22_X1 U4489 ( .A1(n3942), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3941), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3568) );
  NAND4_X1 U4490 ( .A1(n3571), .A2(n3570), .A3(n3569), .A4(n3568), .ZN(n3572)
         );
  NAND2_X1 U4491 ( .A1(n3736), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3575) );
  NAND2_X1 U4492 ( .A1(n6533), .A2(n4016), .ZN(n3574) );
  OAI211_X1 U4493 ( .C1(n4070), .C2(n3606), .A(n3575), .B(n3574), .ZN(n3614)
         );
  INV_X1 U4494 ( .A(n3576), .ZN(n3579) );
  INV_X1 U4495 ( .A(n3577), .ZN(n3578) );
  NAND2_X1 U4496 ( .A1(n3579), .A2(n3578), .ZN(n3580) );
  INV_X1 U4497 ( .A(n3626), .ZN(n3582) );
  NAND2_X1 U4498 ( .A1(n3582), .A2(n6529), .ZN(n3609) );
  NAND2_X1 U4499 ( .A1(n3736), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3605) );
  INV_X1 U4500 ( .A(n4070), .ZN(n3602) );
  AOI22_X1 U4501 ( .A1(n3951), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3583), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3591) );
  AOI22_X1 U4502 ( .A1(n3949), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3947), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3590) );
  AOI22_X1 U4503 ( .A1(n3942), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3948), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3589) );
  AOI22_X1 U4504 ( .A1(n3938), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3588) );
  NAND4_X1 U4505 ( .A1(n3591), .A2(n3590), .A3(n3589), .A4(n3588), .ZN(n3600)
         );
  AOI22_X1 U4506 ( .A1(n3939), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3650), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3598) );
  AOI22_X1 U4507 ( .A1(n3915), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3551), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3597) );
  AOI22_X1 U4508 ( .A1(n3769), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3596) );
  AOI22_X1 U4509 ( .A1(n3941), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3952), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3595) );
  NAND4_X1 U4510 ( .A1(n3598), .A2(n3597), .A3(n3596), .A4(n3595), .ZN(n3599)
         );
  NAND2_X1 U4511 ( .A1(n4130), .A2(n4024), .ZN(n3601) );
  OAI211_X1 U4512 ( .C1(n3602), .C2(n4479), .A(STATE2_REG_0__SCAN_IN), .B(
        n3601), .ZN(n3603) );
  INV_X1 U4513 ( .A(n3603), .ZN(n3604) );
  NAND2_X1 U4514 ( .A1(n3605), .A2(n3604), .ZN(n3623) );
  XNOR2_X1 U4515 ( .A(n4024), .B(n4070), .ZN(n3607) );
  NOR2_X1 U4516 ( .A1(n3607), .A2(n3606), .ZN(n3622) );
  NAND2_X1 U4517 ( .A1(n3623), .A2(n3622), .ZN(n3608) );
  NAND2_X1 U4518 ( .A1(n3610), .A2(n4070), .ZN(n3995) );
  OAI21_X1 U4519 ( .B1(n3616), .B2(n3614), .A(n3615), .ZN(n3612) );
  NAND2_X1 U4520 ( .A1(n3616), .A2(n3614), .ZN(n3611) );
  NOR2_X2 U4522 ( .A1(n4455), .A2(n6522), .ZN(n3871) );
  NAND2_X1 U4523 ( .A1(n5835), .A2(n3871), .ZN(n3613) );
  NAND2_X1 U4524 ( .A1(n3613), .A2(n3828), .ZN(n4303) );
  XNOR2_X1 U4525 ( .A(n3615), .B(n3614), .ZN(n3617) );
  NAND2_X1 U4526 ( .A1(n4369), .A2(n3871), .ZN(n3621) );
  AOI22_X1 U4527 ( .A1(n3972), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6522), .ZN(n3619) );
  AND2_X1 U4528 ( .A1(n4141), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3630) );
  NAND2_X1 U4529 ( .A1(n3630), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3618) );
  AND2_X1 U4530 ( .A1(n3619), .A2(n3618), .ZN(n3620) );
  NAND2_X1 U4531 ( .A1(n3621), .A2(n3620), .ZN(n4259) );
  OR2_X1 U4532 ( .A1(n3623), .A2(n3622), .ZN(n3624) );
  AOI21_X1 U4533 ( .B1(n5026), .B2(n4241), .A(n6522), .ZN(n4207) );
  INV_X1 U4534 ( .A(n4903), .ZN(n5017) );
  INV_X1 U4535 ( .A(n3630), .ZN(n3690) );
  NAND2_X1 U4536 ( .A1(n3972), .A2(EAX_REG_0__SCAN_IN), .ZN(n3628) );
  NAND2_X1 U4537 ( .A1(n6522), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n3627)
         );
  OAI211_X1 U4538 ( .C1(n3690), .C2(n4198), .A(n3628), .B(n3627), .ZN(n3629)
         );
  AOI21_X1 U4539 ( .B1(n5017), .B2(n3871), .A(n3629), .ZN(n4206) );
  MUX2_X1 U4540 ( .A(n4207), .B(n3968), .S(n4206), .Z(n4258) );
  NAND2_X1 U4541 ( .A1(n4259), .A2(n4258), .ZN(n4257) );
  NAND2_X1 U4542 ( .A1(n3630), .A2(n6552), .ZN(n3636) );
  INV_X1 U4543 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3633) );
  OAI21_X1 U4544 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3631), .ZN(n6181) );
  NAND2_X1 U4545 ( .A1(n3968), .A2(n6181), .ZN(n3632) );
  OAI21_X1 U4546 ( .B1(n3633), .B2(n3828), .A(n3632), .ZN(n3634) );
  AOI21_X1 U4547 ( .B1(n3972), .B2(EAX_REG_2__SCAN_IN), .A(n3634), .ZN(n3635)
         );
  AND2_X1 U4548 ( .A1(n3636), .A2(n3635), .ZN(n3638) );
  NAND2_X1 U4549 ( .A1(n4257), .A2(n3638), .ZN(n4304) );
  INV_X1 U4550 ( .A(n3641), .ZN(n3643) );
  NAND2_X1 U4551 ( .A1(n3644), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3649) );
  NAND3_X1 U4552 ( .A1(n4970), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4809) );
  INV_X1 U4553 ( .A(n4809), .ZN(n4811) );
  NAND2_X1 U4554 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4811), .ZN(n6325) );
  NAND2_X1 U4555 ( .A1(n4970), .A2(n6325), .ZN(n3645) );
  NOR3_X1 U4556 ( .A1(n4970), .A2(n6399), .A3(n6393), .ZN(n4919) );
  NAND2_X1 U4557 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4919), .ZN(n4672) );
  AND2_X1 U4558 ( .A1(n3645), .A2(n4672), .ZN(n4753) );
  AOI22_X1 U4559 ( .A1(n3647), .A2(n4753), .B1(n3646), .B2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3648) );
  AOI22_X1 U4560 ( .A1(n3939), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3650), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3654) );
  AOI22_X1 U4561 ( .A1(n3915), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3653) );
  AOI22_X1 U4562 ( .A1(n3551), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3652) );
  AOI22_X1 U4563 ( .A1(n3938), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3651) );
  NAND4_X1 U4564 ( .A1(n3654), .A2(n3653), .A3(n3652), .A4(n3651), .ZN(n3660)
         );
  AOI22_X1 U4565 ( .A1(n3769), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3947), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3658) );
  AOI22_X1 U4566 ( .A1(n3949), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3657) );
  AOI22_X1 U4567 ( .A1(n3782), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3952), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3656) );
  AOI22_X1 U4568 ( .A1(n3948), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3941), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3655) );
  NAND4_X1 U4569 ( .A1(n3658), .A2(n3657), .A3(n3656), .A4(n3655), .ZN(n3659)
         );
  OR2_X1 U4570 ( .A1(n3660), .A2(n3659), .ZN(n4004) );
  AOI22_X1 U4571 ( .A1(n3736), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3737), 
        .B2(n4004), .ZN(n3661) );
  NAND2_X1 U4572 ( .A1(n3736), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3674) );
  AOI22_X1 U4573 ( .A1(n3939), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3666) );
  AOI22_X1 U4574 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n3915), .B1(n3921), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3665) );
  AOI22_X1 U4575 ( .A1(n3551), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3664) );
  AOI22_X1 U4576 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n3938), .B1(n3950), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3663) );
  NAND4_X1 U4577 ( .A1(n3666), .A2(n3665), .A3(n3664), .A4(n3663), .ZN(n3672)
         );
  AOI22_X1 U4578 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n3947), .B1(n3769), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3670) );
  AOI22_X1 U4579 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n3949), .B1(n3942), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3669) );
  AOI22_X1 U4580 ( .A1(n3782), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3952), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3668) );
  AOI22_X1 U4581 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n3948), .B1(n3941), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3667) );
  NAND4_X1 U4582 ( .A1(n3670), .A2(n3669), .A3(n3668), .A4(n3667), .ZN(n3671)
         );
  OR2_X1 U4583 ( .A1(n3672), .A2(n3671), .ZN(n4047) );
  NAND2_X1 U4584 ( .A1(n3737), .A2(n4047), .ZN(n3673) );
  NAND2_X1 U4585 ( .A1(n3674), .A2(n3673), .ZN(n3712) );
  XNOR2_X1 U4586 ( .A(n3714), .B(n3712), .ZN(n4040) );
  NAND2_X1 U4587 ( .A1(n6522), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3676)
         );
  NAND2_X1 U4588 ( .A1(n3972), .A2(EAX_REG_4__SCAN_IN), .ZN(n3675) );
  OAI211_X1 U4589 ( .C1(n3690), .C2(n5924), .A(n3676), .B(n3675), .ZN(n3677)
         );
  NAND2_X1 U4590 ( .A1(n3677), .A2(n3963), .ZN(n3679) );
  OAI21_X1 U4591 ( .B1(n3687), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n3707), 
        .ZN(n6170) );
  NAND2_X1 U4592 ( .A1(n6170), .A2(n3968), .ZN(n3678) );
  NAND2_X1 U4593 ( .A1(n3679), .A2(n3678), .ZN(n3680) );
  AOI21_X1 U4594 ( .B1(n4040), .B2(n3871), .A(n3680), .ZN(n4399) );
  NAND2_X1 U4595 ( .A1(n3682), .A2(n3681), .ZN(n3683) );
  INV_X1 U4596 ( .A(n4626), .ZN(n4371) );
  NAND2_X1 U4597 ( .A1(n3683), .A2(n4371), .ZN(n3684) );
  NOR2_X1 U4598 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n3685), .ZN(n3686)
         );
  NOR2_X1 U4599 ( .A1(n3687), .A2(n3686), .ZN(n6045) );
  INV_X1 U4600 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6035) );
  OAI22_X1 U4601 ( .A1(n6045), .A2(n3963), .B1(n3828), .B2(n6035), .ZN(n3688)
         );
  AOI21_X1 U4602 ( .B1(n3972), .B2(EAX_REG_3__SCAN_IN), .A(n3688), .ZN(n3689)
         );
  OAI21_X1 U4603 ( .B1(n4344), .B2(n3690), .A(n3689), .ZN(n3691) );
  AOI21_X1 U4604 ( .B1(n4749), .B2(n3871), .A(n3691), .ZN(n4317) );
  OR2_X2 U4605 ( .A1(n4399), .A2(n4317), .ZN(n3692) );
  INV_X1 U4606 ( .A(n3712), .ZN(n3693) );
  OR2_X1 U4607 ( .A1(n3714), .A2(n3693), .ZN(n3706) );
  NAND2_X1 U4608 ( .A1(n3736), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3705) );
  AOI22_X1 U4609 ( .A1(n3939), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3697) );
  AOI22_X1 U4610 ( .A1(n3915), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3696) );
  AOI22_X1 U4611 ( .A1(n3551), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3695) );
  AOI22_X1 U4612 ( .A1(n3938), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3694) );
  NAND4_X1 U4613 ( .A1(n3697), .A2(n3696), .A3(n3695), .A4(n3694), .ZN(n3703)
         );
  AOI22_X1 U4614 ( .A1(n3769), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3947), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3701) );
  INV_X1 U4615 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n6578) );
  AOI22_X1 U4616 ( .A1(n3949), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3700) );
  AOI22_X1 U4617 ( .A1(n3916), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3952), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3699) );
  AOI22_X1 U4618 ( .A1(n3948), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3941), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3698) );
  NAND4_X1 U4619 ( .A1(n3701), .A2(n3700), .A3(n3699), .A4(n3698), .ZN(n3702)
         );
  OR2_X1 U4620 ( .A1(n3703), .A2(n3702), .ZN(n4050) );
  NAND2_X1 U4621 ( .A1(n3737), .A2(n4050), .ZN(n3704) );
  NAND2_X1 U4622 ( .A1(n3705), .A2(n3704), .ZN(n3711) );
  XNOR2_X1 U4623 ( .A(n3707), .B(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4880) );
  OAI22_X1 U4624 ( .A1(n4880), .A2(n3963), .B1(n3828), .B2(n4874), .ZN(n3708)
         );
  AOI21_X1 U4625 ( .B1(n3972), .B2(EAX_REG_5__SCAN_IN), .A(n3708), .ZN(n3709)
         );
  NAND2_X1 U4626 ( .A1(n3712), .A2(n3711), .ZN(n3713) );
  AOI22_X1 U4627 ( .A1(n3939), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3718) );
  AOI22_X1 U4628 ( .A1(n3915), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3717) );
  AOI22_X1 U4629 ( .A1(n3551), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3716) );
  AOI22_X1 U4630 ( .A1(n3938), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3715) );
  NAND4_X1 U4631 ( .A1(n3718), .A2(n3717), .A3(n3716), .A4(n3715), .ZN(n3724)
         );
  AOI22_X1 U4632 ( .A1(n3769), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3947), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3722) );
  AOI22_X1 U4633 ( .A1(n3949), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3721) );
  AOI22_X1 U4634 ( .A1(n3782), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3952), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3720) );
  AOI22_X1 U4635 ( .A1(n3948), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3941), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3719) );
  NAND4_X1 U4636 ( .A1(n3722), .A2(n3721), .A3(n3720), .A4(n3719), .ZN(n3723)
         );
  OR2_X1 U4637 ( .A1(n3724), .A2(n3723), .ZN(n4060) );
  AOI22_X1 U4638 ( .A1(n3736), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3737), 
        .B2(n4060), .ZN(n3733) );
  NAND2_X1 U4639 ( .A1(n3732), .A2(n3733), .ZN(n4057) );
  INV_X1 U4640 ( .A(EAX_REG_6__SCAN_IN), .ZN(n3728) );
  OR2_X1 U4641 ( .A1(n3725), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3726) );
  NAND2_X1 U4642 ( .A1(n3742), .A2(n3726), .ZN(n6160) );
  INV_X1 U4643 ( .A(n3828), .ZN(n3971) );
  AOI22_X1 U4644 ( .A1(n6160), .A2(n3968), .B1(n3971), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3727) );
  OAI21_X1 U4645 ( .B1(n3930), .B2(n3728), .A(n3727), .ZN(n3729) );
  INV_X1 U4646 ( .A(n3733), .ZN(n3734) );
  NAND2_X1 U4647 ( .A1(n3736), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3739) );
  NAND2_X1 U4648 ( .A1(n3737), .A2(n4070), .ZN(n3738) );
  NAND2_X1 U4649 ( .A1(n3739), .A2(n3738), .ZN(n3740) );
  INV_X1 U4650 ( .A(EAX_REG_7__SCAN_IN), .ZN(n3745) );
  XNOR2_X1 U4651 ( .A(n3742), .B(n3741), .ZN(n4843) );
  NAND2_X1 U4652 ( .A1(n4843), .A2(n3878), .ZN(n3744) );
  NAND2_X1 U4653 ( .A1(n3971), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3743)
         );
  OAI211_X1 U4654 ( .C1(n3930), .C2(n3745), .A(n3744), .B(n3743), .ZN(n3746)
         );
  NOR2_X2 U4655 ( .A1(n4518), .A2(n4519), .ZN(n4615) );
  INV_X1 U4656 ( .A(n3871), .ZN(n3764) );
  AOI22_X1 U4657 ( .A1(n3939), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3750) );
  AOI22_X1 U4658 ( .A1(n3921), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3551), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3749) );
  AOI22_X1 U4659 ( .A1(n3949), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3948), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3748) );
  AOI22_X1 U4660 ( .A1(n3947), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3952), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3747) );
  NAND4_X1 U4661 ( .A1(n3750), .A2(n3749), .A3(n3748), .A4(n3747), .ZN(n3756)
         );
  AOI22_X1 U4662 ( .A1(n3915), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3754) );
  AOI22_X1 U4663 ( .A1(n3938), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3753) );
  AOI22_X1 U4664 ( .A1(n3769), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3752) );
  AOI22_X1 U4665 ( .A1(n3942), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3941), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3751) );
  NAND4_X1 U4666 ( .A1(n3754), .A2(n3753), .A3(n3752), .A4(n3751), .ZN(n3755)
         );
  NOR2_X1 U4667 ( .A1(n3756), .A2(n3755), .ZN(n3763) );
  NAND2_X1 U4668 ( .A1(n3757), .A2(n6569), .ZN(n3759) );
  INV_X1 U4669 ( .A(n3776), .ZN(n3758) );
  NAND2_X1 U4670 ( .A1(n3759), .A2(n3758), .ZN(n4963) );
  NOR2_X1 U4671 ( .A1(n3828), .A2(n6569), .ZN(n3760) );
  AOI21_X1 U4672 ( .B1(n4963), .B2(n3878), .A(n3760), .ZN(n3762) );
  NAND2_X1 U4673 ( .A1(n3972), .A2(EAX_REG_8__SCAN_IN), .ZN(n3761) );
  OAI211_X1 U4674 ( .C1(n3764), .C2(n3763), .A(n3762), .B(n3761), .ZN(n4614)
         );
  NAND2_X1 U4675 ( .A1(n4615), .A2(n4614), .ZN(n4613) );
  AOI22_X1 U4676 ( .A1(n3951), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3551), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3768) );
  AOI22_X1 U4677 ( .A1(n3942), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3948), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3767) );
  AOI22_X1 U4678 ( .A1(n3939), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3766) );
  AOI22_X1 U4679 ( .A1(n2957), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3952), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3765) );
  NAND4_X1 U4680 ( .A1(n3768), .A2(n3767), .A3(n3766), .A4(n3765), .ZN(n3775)
         );
  AOI22_X1 U4681 ( .A1(n3938), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3773) );
  AOI22_X1 U4682 ( .A1(n3915), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3947), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3772) );
  AOI22_X1 U4683 ( .A1(n3769), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3771) );
  AOI22_X1 U4684 ( .A1(n3949), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3941), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3770) );
  NAND4_X1 U4685 ( .A1(n3773), .A2(n3772), .A3(n3771), .A4(n3770), .ZN(n3774)
         );
  OAI21_X1 U4686 ( .B1(n3775), .B2(n3774), .A(n3871), .ZN(n3780) );
  NAND2_X1 U4687 ( .A1(n3972), .A2(EAX_REG_9__SCAN_IN), .ZN(n3779) );
  INV_X1 U4688 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5994) );
  XNOR2_X1 U4689 ( .A(n5994), .B(n3776), .ZN(n5998) );
  INV_X1 U4690 ( .A(n5998), .ZN(n3777) );
  AOI22_X1 U4691 ( .A1(n3971), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .B1(n3968), 
        .B2(n3777), .ZN(n3778) );
  AND3_X1 U4692 ( .A1(n3780), .A2(n3779), .A3(n3778), .ZN(n4837) );
  NOR2_X2 U4693 ( .A1(n4613), .A2(n4837), .ZN(n4838) );
  XNOR2_X1 U4694 ( .A(n5983), .B(n3781), .ZN(n6149) );
  AOI22_X1 U4695 ( .A1(n3915), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3551), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3786) );
  AOI22_X1 U4696 ( .A1(n3949), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3785) );
  AOI22_X1 U4697 ( .A1(n3769), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3784) );
  AOI22_X1 U4698 ( .A1(n3782), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3952), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3783) );
  NAND4_X1 U4699 ( .A1(n3786), .A2(n3785), .A3(n3784), .A4(n3783), .ZN(n3792)
         );
  AOI22_X1 U4700 ( .A1(n3939), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3790) );
  AOI22_X1 U4701 ( .A1(n3951), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3947), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3789) );
  AOI22_X1 U4702 ( .A1(n3938), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3788) );
  AOI22_X1 U4703 ( .A1(n3948), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3941), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3787) );
  NAND4_X1 U4704 ( .A1(n3790), .A2(n3789), .A3(n3788), .A4(n3787), .ZN(n3791)
         );
  OAI21_X1 U4705 ( .B1(n3792), .B2(n3791), .A(n3871), .ZN(n3795) );
  NAND2_X1 U4706 ( .A1(n3972), .A2(EAX_REG_11__SCAN_IN), .ZN(n3794) );
  NAND2_X1 U4707 ( .A1(n3971), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3793)
         );
  NAND3_X1 U4708 ( .A1(n3795), .A2(n3794), .A3(n3793), .ZN(n3796) );
  AOI21_X1 U4709 ( .B1(n6149), .B2(n3878), .A(n3796), .ZN(n5095) );
  AOI22_X1 U4710 ( .A1(n3915), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3800) );
  AOI22_X1 U4711 ( .A1(n3769), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3947), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3799) );
  AOI22_X1 U4712 ( .A1(n3551), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3798) );
  AOI22_X1 U4713 ( .A1(n3948), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3797) );
  NAND4_X1 U4714 ( .A1(n3800), .A2(n3799), .A3(n3798), .A4(n3797), .ZN(n3806)
         );
  AOI22_X1 U4715 ( .A1(n3939), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3804) );
  AOI22_X1 U4716 ( .A1(n3937), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3803) );
  AOI22_X1 U4717 ( .A1(n3942), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3941), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3802) );
  AOI22_X1 U4718 ( .A1(n3949), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3952), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3801) );
  NAND4_X1 U4719 ( .A1(n3804), .A2(n3803), .A3(n3802), .A4(n3801), .ZN(n3805)
         );
  OAI21_X1 U4720 ( .B1(n3806), .B2(n3805), .A(n3871), .ZN(n3811) );
  NAND2_X1 U4721 ( .A1(n3972), .A2(EAX_REG_10__SCAN_IN), .ZN(n3810) );
  INV_X1 U4722 ( .A(n3807), .ZN(n3808) );
  XNOR2_X1 U4723 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3808), .ZN(n5132)
         );
  AOI22_X1 U4724 ( .A1(n3968), .A2(n5132), .B1(n3971), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3809) );
  AND3_X1 U4725 ( .A1(n3811), .A2(n3810), .A3(n3809), .ZN(n4911) );
  AOI22_X1 U4726 ( .A1(n3972), .A2(EAX_REG_12__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n6522), .ZN(n3825) );
  XNOR2_X1 U4727 ( .A(n3812), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5974)
         );
  NAND2_X1 U4728 ( .A1(n5974), .A2(n3878), .ZN(n3824) );
  AOI22_X1 U4729 ( .A1(n3938), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3816) );
  AOI22_X1 U4730 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n3915), .B1(n3939), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3815) );
  AOI22_X1 U4731 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n2959), .B1(n2957), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3814) );
  AOI22_X1 U4732 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n3769), .B1(n3948), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3813) );
  NAND4_X1 U4733 ( .A1(n3816), .A2(n3815), .A3(n3814), .A4(n3813), .ZN(n3822)
         );
  AOI22_X1 U4734 ( .A1(n3951), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3820) );
  AOI22_X1 U4735 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n3947), .B1(n3916), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3819) );
  AOI22_X1 U4736 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n3942), .B1(n3941), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3818) );
  AOI22_X1 U4737 ( .A1(n3949), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3952), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3817) );
  NAND4_X1 U4738 ( .A1(n3820), .A2(n3819), .A3(n3818), .A4(n3817), .ZN(n3821)
         );
  OAI21_X1 U4739 ( .B1(n3822), .B2(n3821), .A(n3871), .ZN(n3823) );
  OAI211_X1 U4740 ( .C1(n3968), .C2(n3825), .A(n3824), .B(n3823), .ZN(n5110)
         );
  INV_X1 U4741 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3829) );
  OAI21_X1 U4742 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n3826), .A(n3847), 
        .ZN(n5969) );
  NAND2_X1 U4743 ( .A1(n5969), .A2(n3878), .ZN(n3827) );
  OAI21_X1 U4744 ( .B1(n3829), .B2(n3828), .A(n3827), .ZN(n3830) );
  AOI21_X1 U4745 ( .B1(n3972), .B2(EAX_REG_13__SCAN_IN), .A(n3830), .ZN(n3831)
         );
  NAND2_X1 U4746 ( .A1(n3832), .A2(n3831), .ZN(n3834) );
  INV_X1 U4747 ( .A(n3833), .ZN(n3846) );
  AND2_X2 U4748 ( .A1(n3834), .A2(n3846), .ZN(n5144) );
  AOI22_X1 U4749 ( .A1(n3938), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3838) );
  AOI22_X1 U4750 ( .A1(n3915), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3551), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3837) );
  AOI22_X1 U4751 ( .A1(n3942), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3952), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3836) );
  AOI22_X1 U4752 ( .A1(n3948), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3941), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3835) );
  NAND4_X1 U4753 ( .A1(n3838), .A2(n3837), .A3(n3836), .A4(n3835), .ZN(n3844)
         );
  AOI22_X1 U4754 ( .A1(n3769), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3947), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3842) );
  AOI22_X1 U4755 ( .A1(n3951), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3841) );
  AOI22_X1 U4756 ( .A1(n3949), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4757 ( .A1(n3939), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3922), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3839) );
  NAND4_X1 U4758 ( .A1(n3842), .A2(n3841), .A3(n3840), .A4(n3839), .ZN(n3843)
         );
  OR2_X1 U4759 ( .A1(n3844), .A2(n3843), .ZN(n3845) );
  AND2_X1 U4760 ( .A1(n3871), .A2(n3845), .ZN(n5145) );
  XOR2_X1 U4761 ( .A(n5231), .B(n3847), .Z(n5284) );
  AOI22_X1 U4762 ( .A1(n3915), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3851) );
  AOI22_X1 U4763 ( .A1(n3942), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3948), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3850) );
  AOI22_X1 U4764 ( .A1(n2958), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3849) );
  AOI22_X1 U4765 ( .A1(n3949), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3952), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3848) );
  NAND4_X1 U4766 ( .A1(n3851), .A2(n3850), .A3(n3849), .A4(n3848), .ZN(n3857)
         );
  AOI22_X1 U4767 ( .A1(n3939), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4768 ( .A1(n3947), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3854) );
  AOI22_X1 U4769 ( .A1(n3938), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3922), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3853) );
  AOI22_X1 U4770 ( .A1(n3769), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3941), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3852) );
  NAND4_X1 U4771 ( .A1(n3855), .A2(n3854), .A3(n3853), .A4(n3852), .ZN(n3856)
         );
  OR2_X1 U4772 ( .A1(n3857), .A2(n3856), .ZN(n3858) );
  AOI22_X1 U4773 ( .A1(n3871), .A2(n3858), .B1(n3971), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3860) );
  NAND2_X1 U4774 ( .A1(n3972), .A2(EAX_REG_14__SCAN_IN), .ZN(n3859) );
  OAI211_X1 U4775 ( .C1(n5284), .C2(n3963), .A(n3860), .B(n3859), .ZN(n5221)
         );
  XNOR2_X1 U4776 ( .A(n3862), .B(n3861), .ZN(n5274) );
  AOI22_X1 U4777 ( .A1(n3915), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3866) );
  AOI22_X1 U4778 ( .A1(n3769), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3865) );
  AOI22_X1 U4779 ( .A1(n3949), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3864) );
  AOI22_X1 U4780 ( .A1(n3948), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3941), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3863) );
  NAND4_X1 U4781 ( .A1(n3866), .A2(n3865), .A3(n3864), .A4(n3863), .ZN(n3873)
         );
  AOI22_X1 U4782 ( .A1(n3939), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3870) );
  AOI22_X1 U4783 ( .A1(n2959), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3947), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3869) );
  AOI22_X1 U4784 ( .A1(n3938), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3922), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3868) );
  AOI22_X1 U4785 ( .A1(n3942), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3952), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3867) );
  NAND4_X1 U4786 ( .A1(n3870), .A2(n3869), .A3(n3868), .A4(n3867), .ZN(n3872)
         );
  OAI21_X1 U4787 ( .B1(n3873), .B2(n3872), .A(n3871), .ZN(n3876) );
  NAND2_X1 U4788 ( .A1(n3972), .A2(EAX_REG_15__SCAN_IN), .ZN(n3875) );
  NAND2_X1 U4789 ( .A1(n3971), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3874)
         );
  NAND3_X1 U4790 ( .A1(n3876), .A2(n3875), .A3(n3874), .ZN(n3877) );
  AOI21_X1 U4791 ( .B1(n5274), .B2(n3878), .A(n3877), .ZN(n5238) );
  XOR2_X1 U4792 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n3879), .Z(n5687) );
  INV_X1 U4793 ( .A(n5687), .ZN(n3893) );
  AOI22_X1 U4794 ( .A1(n3939), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3883) );
  AOI22_X1 U4795 ( .A1(n3949), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3376), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3882) );
  AOI22_X1 U4796 ( .A1(n3915), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3881) );
  AOI22_X1 U4797 ( .A1(n3937), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3922), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3880) );
  NAND4_X1 U4798 ( .A1(n3883), .A2(n3882), .A3(n3881), .A4(n3880), .ZN(n3889)
         );
  AOI22_X1 U4799 ( .A1(n3938), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3551), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3887) );
  AOI22_X1 U4800 ( .A1(n3947), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3886) );
  AOI22_X1 U4801 ( .A1(n3948), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3941), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3885) );
  AOI22_X1 U4802 ( .A1(n3942), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3952), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3884) );
  NAND4_X1 U4803 ( .A1(n3887), .A2(n3886), .A3(n3885), .A4(n3884), .ZN(n3888)
         );
  NOR2_X1 U4804 ( .A1(n3889), .A2(n3888), .ZN(n3891) );
  AOI22_X1 U4805 ( .A1(n3972), .A2(EAX_REG_16__SCAN_IN), .B1(n3971), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3890) );
  OAI21_X1 U4806 ( .B1(n3966), .B2(n3891), .A(n3890), .ZN(n3892) );
  AOI21_X1 U4807 ( .B1(n3893), .B2(n3968), .A(n3892), .ZN(n5254) );
  XNOR2_X1 U4808 ( .A(n3894), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5882)
         );
  AOI22_X1 U4809 ( .A1(n3938), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n2959), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3900) );
  NAND2_X1 U4810 ( .A1(n3937), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3896) );
  NAND2_X1 U4811 ( .A1(n3948), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3895) );
  AND3_X1 U4812 ( .A1(n3896), .A2(n3895), .A3(n3963), .ZN(n3899) );
  AOI22_X1 U4813 ( .A1(n3942), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3898) );
  AOI22_X1 U4814 ( .A1(n3951), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3952), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3897) );
  NAND4_X1 U4815 ( .A1(n3900), .A2(n3899), .A3(n3898), .A4(n3897), .ZN(n3906)
         );
  AOI22_X1 U4816 ( .A1(n3915), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3376), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3904) );
  AOI22_X1 U4817 ( .A1(n3949), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3939), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3903) );
  AOI22_X1 U4818 ( .A1(n2957), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3922), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3902) );
  AOI22_X1 U4819 ( .A1(n3947), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3941), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3901) );
  NAND4_X1 U4820 ( .A1(n3904), .A2(n3903), .A3(n3902), .A4(n3901), .ZN(n3905)
         );
  OR2_X1 U4821 ( .A1(n3906), .A2(n3905), .ZN(n3909) );
  INV_X1 U4822 ( .A(EAX_REG_17__SCAN_IN), .ZN(n3907) );
  OAI22_X1 U4823 ( .A1(n3930), .A2(n3907), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5294), .ZN(n3908) );
  AOI21_X1 U4824 ( .B1(n3910), .B2(n3909), .A(n3908), .ZN(n3911) );
  AOI21_X1 U4825 ( .B1(n5882), .B2(n3968), .A(n3911), .ZN(n5290) );
  NOR2_X1 U4826 ( .A1(n3912), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3913)
         );
  OR2_X1 U4827 ( .A1(n3914), .A2(n3913), .ZN(n5678) );
  INV_X1 U4828 ( .A(n5678), .ZN(n5949) );
  AOI22_X1 U4829 ( .A1(n3915), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3650), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3920) );
  AOI22_X1 U4830 ( .A1(n3551), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3947), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3919) );
  AOI22_X1 U4831 ( .A1(n3942), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3918) );
  AOI22_X1 U4832 ( .A1(n3948), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3941), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3917) );
  NAND4_X1 U4833 ( .A1(n3920), .A2(n3919), .A3(n3918), .A4(n3917), .ZN(n3928)
         );
  AOI22_X1 U4834 ( .A1(n3939), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3926) );
  AOI22_X1 U4835 ( .A1(n3769), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3925) );
  AOI22_X1 U4836 ( .A1(n3938), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3922), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3924) );
  AOI22_X1 U4837 ( .A1(n3949), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3952), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3923) );
  NAND4_X1 U4838 ( .A1(n3926), .A2(n3925), .A3(n3924), .A4(n3923), .ZN(n3927)
         );
  OR2_X1 U4839 ( .A1(n3928), .A2(n3927), .ZN(n3932) );
  INV_X1 U4840 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4315) );
  NAND2_X1 U4841 ( .A1(n6522), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3929)
         );
  OAI211_X1 U4842 ( .C1(n3930), .C2(n4315), .A(n3963), .B(n3929), .ZN(n3931)
         );
  AOI21_X1 U4843 ( .B1(n3933), .B2(n3932), .A(n3931), .ZN(n3934) );
  AOI21_X1 U4844 ( .B1(n5949), .B2(n3968), .A(n3934), .ZN(n5552) );
  NAND2_X1 U4846 ( .A1(n3936), .A2(n4116), .ZN(n5433) );
  AOI22_X1 U4847 ( .A1(n3938), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3946) );
  AOI22_X1 U4848 ( .A1(n3915), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3939), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3945) );
  AOI22_X1 U4849 ( .A1(n2958), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3944) );
  AOI22_X1 U4850 ( .A1(n3942), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3941), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3943) );
  NAND4_X1 U4851 ( .A1(n3946), .A2(n3945), .A3(n3944), .A4(n3943), .ZN(n3958)
         );
  AOI22_X1 U4852 ( .A1(n3947), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n2957), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3956) );
  AOI22_X1 U4853 ( .A1(n3949), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3948), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3955) );
  AOI22_X1 U4854 ( .A1(n3951), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3950), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3954) );
  AOI22_X1 U4855 ( .A1(n3376), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3952), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3953) );
  NAND4_X1 U4856 ( .A1(n3956), .A2(n3955), .A3(n3954), .A4(n3953), .ZN(n3957)
         );
  NOR2_X1 U4857 ( .A1(n3958), .A2(n3957), .ZN(n3962) );
  NOR2_X1 U4858 ( .A1(n3960), .A2(n3959), .ZN(n3961) );
  XOR2_X1 U4859 ( .A(n3962), .B(n3961), .Z(n3967) );
  INV_X1 U4860 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n6571) );
  OAI21_X1 U4861 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6571), .A(n3963), .ZN(
        n3964) );
  AOI21_X1 U4862 ( .B1(n3972), .B2(EAX_REG_30__SCAN_IN), .A(n3964), .ZN(n3965)
         );
  OAI21_X1 U4863 ( .B1(n3967), .B2(n3966), .A(n3965), .ZN(n3970) );
  XNOR2_X1 U4864 ( .A(n3975), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5440)
         );
  NAND2_X1 U4865 ( .A1(n5440), .A2(n3968), .ZN(n3969) );
  NAND2_X1 U4866 ( .A1(n3970), .A2(n3969), .ZN(n5432) );
  NOR2_X1 U4867 ( .A1(n5433), .A2(n5432), .ZN(n3974) );
  AOI22_X1 U4868 ( .A1(n3972), .A2(EAX_REG_31__SCAN_IN), .B1(n3971), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n3973) );
  XNOR2_X1 U4869 ( .A(n3974), .B(n3973), .ZN(n5598) );
  INV_X1 U4870 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n3976) );
  XNOR2_X1 U4871 ( .A(n3977), .B(n3976), .ZN(n5596) );
  NOR2_X1 U4872 ( .A1(n5596), .A2(n4364), .ZN(n3978) );
  INV_X1 U4873 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6478) );
  INV_X1 U4874 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6673) );
  NAND2_X1 U4875 ( .A1(n4171), .A2(n6528), .ZN(n4231) );
  NOR2_X1 U4876 ( .A1(n4893), .A2(n3980), .ZN(n3981) );
  AND2_X1 U4877 ( .A1(n4460), .A2(n3981), .ZN(n3982) );
  INV_X1 U4878 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6470) );
  INV_X1 U4879 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6457) );
  INV_X1 U4880 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6456) );
  NAND3_X1 U4881 ( .A1(REIP_REG_2__SCAN_IN), .A2(REIP_REG_1__SCAN_IN), .A3(
        REIP_REG_3__SCAN_IN), .ZN(n6020) );
  OR2_X1 U4882 ( .A1(n6456), .A2(n6020), .ZN(n4875) );
  NOR2_X1 U4883 ( .A1(n6457), .A2(n4875), .ZN(n4844) );
  INV_X1 U4884 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6460) );
  INV_X1 U4885 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6459) );
  NOR2_X1 U4886 ( .A1(n6460), .A2(n6459), .ZN(n4862) );
  NAND2_X1 U4887 ( .A1(REIP_REG_8__SCAN_IN), .A2(n4862), .ZN(n4864) );
  INV_X1 U4888 ( .A(n4864), .ZN(n3983) );
  INV_X1 U4889 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6466) );
  NAND2_X1 U4890 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .ZN(
        n5990) );
  NOR2_X1 U4891 ( .A1(n6466), .A2(n5990), .ZN(n5956) );
  INV_X1 U4892 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6472) );
  INV_X1 U4893 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6469) );
  NOR2_X1 U4894 ( .A1(n6472), .A2(n6469), .ZN(n5955) );
  NAND4_X1 U4895 ( .A1(n4844), .A2(n3983), .A3(n5956), .A4(n5955), .ZN(n5227)
         );
  NOR2_X1 U4896 ( .A1(n6470), .A2(n5227), .ZN(n3987) );
  NAND2_X1 U4897 ( .A1(n5118), .A2(n3987), .ZN(n5249) );
  NOR2_X1 U4898 ( .A1(n6673), .A2(n5249), .ZN(n5260) );
  NAND2_X1 U4899 ( .A1(REIP_REG_16__SCAN_IN), .A2(n5260), .ZN(n5293) );
  NOR2_X1 U4900 ( .A1(n6478), .A2(n5293), .ZN(n5951) );
  NAND2_X1 U4901 ( .A1(REIP_REG_18__SCAN_IN), .A2(n5951), .ZN(n5866) );
  NAND2_X1 U4902 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .ZN(
        n3984) );
  NOR2_X1 U4903 ( .A1(n5866), .A2(n3984), .ZN(n5847) );
  NAND4_X1 U4904 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n5847), .ZN(n5508) );
  NAND3_X1 U4905 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n5475) );
  INV_X1 U4906 ( .A(n5475), .ZN(n3985) );
  NAND2_X1 U4907 ( .A1(REIP_REG_27__SCAN_IN), .A2(n3985), .ZN(n3986) );
  NOR2_X1 U4908 ( .A1(n5508), .A2(n3986), .ZN(n5469) );
  NAND2_X1 U4909 ( .A1(n5469), .A2(REIP_REG_28__SCAN_IN), .ZN(n5459) );
  INV_X1 U4910 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6505) );
  INV_X1 U4911 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6501) );
  NAND3_X1 U4912 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n3988) );
  INV_X1 U4913 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6480) );
  NAND2_X1 U4914 ( .A1(n3987), .A2(n5123), .ZN(n5225) );
  NOR2_X1 U4915 ( .A1(n6673), .A2(n5225), .ZN(n5263) );
  NAND3_X1 U4916 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        n5263), .ZN(n5296) );
  NOR2_X1 U4917 ( .A1(n6480), .A2(n5296), .ZN(n5523) );
  NAND3_X1 U4918 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        n5523), .ZN(n5510) );
  OR2_X1 U4919 ( .A1(n3988), .A2(n5510), .ZN(n5325) );
  NAND2_X1 U4920 ( .A1(n5123), .A2(n6021), .ZN(n6015) );
  OAI21_X1 U4921 ( .B1(n5325), .B2(n5475), .A(n6015), .ZN(n5495) );
  AND2_X1 U4922 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n3989) );
  OR2_X1 U4923 ( .A1(n6021), .A2(n3989), .ZN(n3990) );
  NAND2_X1 U4924 ( .A1(n5495), .A2(n3990), .ZN(n5468) );
  AOI21_X1 U4925 ( .B1(n5118), .B2(n6501), .A(n5468), .ZN(n5439) );
  OAI21_X1 U4926 ( .B1(REIP_REG_30__SCAN_IN), .B2(n6021), .A(n5439), .ZN(n3991) );
  NAND4_X1 U4927 ( .A1(n3994), .A2(n3993), .A3(n2961), .A4(n3992), .ZN(U2796)
         );
  INV_X1 U4928 ( .A(n4058), .ZN(n4068) );
  NOR2_X1 U4929 ( .A1(n3995), .A2(n4068), .ZN(n3996) );
  NAND2_X1 U4930 ( .A1(n4024), .A2(n4016), .ZN(n4012) );
  INV_X1 U4931 ( .A(n3997), .ZN(n4011) );
  NAND2_X1 U4932 ( .A1(n4012), .A2(n4011), .ZN(n4006) );
  NAND2_X1 U4933 ( .A1(n4006), .A2(n4004), .ZN(n4049) );
  NAND2_X1 U4934 ( .A1(n4047), .A2(n4050), .ZN(n3998) );
  OR2_X1 U4935 ( .A1(n4049), .A2(n3998), .ZN(n4061) );
  INV_X1 U4936 ( .A(n4061), .ZN(n3999) );
  NAND2_X1 U4937 ( .A1(n3999), .A2(n4060), .ZN(n4071) );
  INV_X1 U4938 ( .A(n4071), .ZN(n4000) );
  NAND3_X1 U4939 ( .A1(n4000), .A2(n3496), .A3(n4070), .ZN(n4001) );
  NAND2_X1 U4940 ( .A1(n4079), .A2(n4001), .ZN(n4077) );
  NAND2_X1 U4941 ( .A1(n4077), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5100)
         );
  OR2_X1 U4942 ( .A1(n5409), .A2(n6195), .ZN(n5103) );
  INV_X1 U4943 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4002) );
  AND2_X1 U4944 ( .A1(n4082), .A2(n4002), .ZN(n4078) );
  NAND2_X1 U4945 ( .A1(n4003), .A2(n4058), .ZN(n4009) );
  INV_X1 U4946 ( .A(n4004), .ZN(n4005) );
  XNOR2_X1 U4947 ( .A(n4006), .B(n4005), .ZN(n4007) );
  NAND2_X1 U4948 ( .A1(n4007), .A2(n3496), .ZN(n4008) );
  NAND2_X1 U4949 ( .A1(n4009), .A2(n4008), .ZN(n4038) );
  XNOR2_X1 U4950 ( .A(n4038), .B(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n5691)
         );
  INV_X1 U4951 ( .A(n5691), .ZN(n4037) );
  NAND2_X1 U4952 ( .A1(n4010), .A2(n4058), .ZN(n4015) );
  XNOR2_X1 U4953 ( .A(n4012), .B(n4011), .ZN(n4013) );
  AND2_X1 U4954 ( .A1(n4130), .A2(n4465), .ZN(n4152) );
  AOI21_X1 U4955 ( .B1(n4013), .B2(n3496), .A(n4152), .ZN(n4014) );
  NAND2_X1 U4956 ( .A1(n6173), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4033)
         );
  NAND2_X1 U4957 ( .A1(n4369), .A2(n4058), .ZN(n4022) );
  XNOR2_X1 U4958 ( .A(n4024), .B(n4016), .ZN(n4019) );
  INV_X1 U4959 ( .A(n3496), .ZN(n4246) );
  INV_X1 U4960 ( .A(n4017), .ZN(n4018) );
  OAI211_X1 U4961 ( .C1(n4019), .C2(n4246), .A(n4018), .B(n4474), .ZN(n4020)
         );
  INV_X1 U4962 ( .A(n4020), .ZN(n4021) );
  NAND2_X1 U4963 ( .A1(n4022), .A2(n4021), .ZN(n4295) );
  NAND2_X1 U4964 ( .A1(n4631), .A2(n4058), .ZN(n4027) );
  INV_X1 U4965 ( .A(n4152), .ZN(n4023) );
  OAI21_X1 U4966 ( .B1(n4246), .B2(n4024), .A(n4023), .ZN(n4025) );
  INV_X1 U4967 ( .A(n4025), .ZN(n4026) );
  NAND2_X1 U4968 ( .A1(n4027), .A2(n4026), .ZN(n4205) );
  NAND2_X1 U4969 ( .A1(n4205), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4028)
         );
  INV_X1 U4970 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5157) );
  NAND2_X1 U4971 ( .A1(n4028), .A2(n5157), .ZN(n4030) );
  AND2_X1 U4972 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4029) );
  NAND2_X1 U4973 ( .A1(n4205), .A2(n4029), .ZN(n4031) );
  AND2_X1 U4974 ( .A1(n4030), .A2(n4031), .ZN(n4296) );
  INV_X1 U4975 ( .A(n4031), .ZN(n4032) );
  AOI21_X1 U4976 ( .B1(n4295), .B2(n4296), .A(n4032), .ZN(n6172) );
  NAND2_X1 U4977 ( .A1(n4033), .A2(n6172), .ZN(n4035) );
  OR2_X1 U4978 ( .A1(n6173), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4034)
         );
  NAND2_X1 U4979 ( .A1(n4035), .A2(n4034), .ZN(n5690) );
  INV_X1 U4980 ( .A(n5690), .ZN(n4036) );
  NAND2_X1 U4981 ( .A1(n4037), .A2(n4036), .ZN(n6248) );
  NAND2_X1 U4982 ( .A1(n4038), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4039)
         );
  NAND2_X1 U4983 ( .A1(n6248), .A2(n4039), .ZN(n6163) );
  NAND2_X1 U4984 ( .A1(n4040), .A2(n4058), .ZN(n4043) );
  XNOR2_X1 U4985 ( .A(n4049), .B(n4047), .ZN(n4041) );
  NAND2_X1 U4986 ( .A1(n4041), .A2(n3496), .ZN(n4042) );
  NAND2_X1 U4987 ( .A1(n4043), .A2(n4042), .ZN(n4044) );
  INV_X1 U4988 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6241) );
  XNOR2_X1 U4989 ( .A(n4044), .B(n6241), .ZN(n6162) );
  NAND2_X1 U4990 ( .A1(n6163), .A2(n6162), .ZN(n6161) );
  NAND2_X1 U4991 ( .A1(n4044), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4045)
         );
  NAND2_X1 U4992 ( .A1(n6161), .A2(n4045), .ZN(n4428) );
  NAND2_X1 U4993 ( .A1(n4046), .A2(n4058), .ZN(n4054) );
  INV_X1 U4994 ( .A(n4047), .ZN(n4048) );
  OR2_X1 U4995 ( .A1(n4049), .A2(n4048), .ZN(n4051) );
  XNOR2_X1 U4996 ( .A(n4051), .B(n4050), .ZN(n4052) );
  NAND2_X1 U4997 ( .A1(n4052), .A2(n3496), .ZN(n4053) );
  NAND2_X1 U4998 ( .A1(n4054), .A2(n4053), .ZN(n4055) );
  INV_X1 U4999 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4432) );
  XNOR2_X1 U5000 ( .A(n4055), .B(n4432), .ZN(n4427) );
  NAND2_X1 U5001 ( .A1(n4428), .A2(n4427), .ZN(n4426) );
  NAND2_X1 U5002 ( .A1(n4055), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4056)
         );
  NAND2_X1 U5003 ( .A1(n4426), .A2(n4056), .ZN(n4888) );
  NAND3_X1 U5004 ( .A1(n4059), .A2(n4058), .A3(n4057), .ZN(n4064) );
  XNOR2_X1 U5005 ( .A(n4061), .B(n4060), .ZN(n4062) );
  NAND2_X1 U5006 ( .A1(n4062), .A2(n3496), .ZN(n4063) );
  NAND2_X1 U5007 ( .A1(n4064), .A2(n4063), .ZN(n4065) );
  INV_X1 U5008 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6655) );
  XNOR2_X1 U5009 ( .A(n4065), .B(n6655), .ZN(n4887) );
  NAND2_X1 U5010 ( .A1(n4888), .A2(n4887), .ZN(n4886) );
  NAND2_X1 U5011 ( .A1(n4065), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4066)
         );
  NAND2_X1 U5012 ( .A1(n4886), .A2(n4066), .ZN(n4801) );
  INV_X1 U5013 ( .A(n4067), .ZN(n4069) );
  XNOR2_X1 U5014 ( .A(n4071), .B(n4070), .ZN(n4072) );
  NAND2_X1 U5015 ( .A1(n4072), .A2(n3496), .ZN(n4073) );
  NAND2_X1 U5016 ( .A1(n4074), .A2(n4073), .ZN(n4075) );
  XNOR2_X1 U5017 ( .A(n4075), .B(n6231), .ZN(n4800) );
  NAND2_X1 U5018 ( .A1(n4801), .A2(n4800), .ZN(n4799) );
  NAND2_X1 U5019 ( .A1(n4075), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4076)
         );
  NAND2_X1 U5020 ( .A1(n4799), .A2(n4076), .ZN(n4960) );
  INV_X1 U5021 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6222) );
  XNOR2_X1 U5022 ( .A(n4077), .B(n6222), .ZN(n4959) );
  NAND2_X1 U5023 ( .A1(n4960), .A2(n4959), .ZN(n4958) );
  NAND2_X1 U5024 ( .A1(n4078), .A2(n4958), .ZN(n4080) );
  NAND2_X1 U5025 ( .A1(n4079), .A2(n6195), .ZN(n5102) );
  AOI21_X2 U5026 ( .B1(n4958), .B2(n4082), .A(n4081), .ZN(n5129) );
  NAND3_X1 U5027 ( .A1(n5129), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4083) );
  NAND2_X1 U5028 ( .A1(n4084), .A2(n4083), .ZN(n5137) );
  INV_X1 U5029 ( .A(n5137), .ZN(n4085) );
  INV_X1 U5030 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4086) );
  NAND2_X2 U5031 ( .A1(n4085), .A2(n2968), .ZN(n5268) );
  NAND2_X1 U5032 ( .A1(n5409), .A2(n4086), .ZN(n5279) );
  INV_X1 U5033 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4090) );
  NAND2_X1 U5034 ( .A1(n4079), .A2(n5354), .ZN(n5280) );
  NAND2_X1 U5035 ( .A1(n5409), .A2(n5906), .ZN(n4087) );
  NAND2_X1 U5036 ( .A1(n5268), .A2(n4088), .ZN(n4096) );
  OR2_X1 U5037 ( .A1(n4079), .A2(n5906), .ZN(n4094) );
  INV_X1 U5038 ( .A(n4089), .ZN(n4093) );
  XNOR2_X1 U5039 ( .A(n5409), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5887)
         );
  OR2_X1 U5040 ( .A1(n5409), .A2(n4090), .ZN(n4091) );
  NAND2_X2 U5041 ( .A1(n4096), .A2(n4095), .ZN(n5672) );
  NAND3_X1 U5042 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A3(INSTADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n4097) );
  NAND2_X2 U5043 ( .A1(n5672), .A2(n2963), .ZN(n5661) );
  INV_X1 U5044 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5898) );
  INV_X1 U5045 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5799) );
  INV_X1 U5046 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6629) );
  AND3_X1 U5047 ( .A1(n5898), .A2(n5799), .A3(n6629), .ZN(n4098) );
  OR2_X1 U5048 ( .A1(n5409), .A2(n4098), .ZN(n5660) );
  INV_X1 U5049 ( .A(n5660), .ZN(n4099) );
  NOR2_X1 U5050 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n4099), .ZN(n4100)
         );
  NAND2_X1 U5051 ( .A1(n5661), .A2(n4100), .ZN(n5662) );
  XNOR2_X1 U5052 ( .A(n4079), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5651)
         );
  INV_X1 U5053 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4102) );
  OR2_X1 U5054 ( .A1(n5409), .A2(n4102), .ZN(n4103) );
  INV_X1 U5055 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5758) );
  XNOR2_X1 U5056 ( .A(n4079), .B(n5758), .ZN(n5645) );
  NOR2_X2 U5057 ( .A1(n5644), .A2(n5645), .ZN(n5643) );
  NOR2_X1 U5058 ( .A1(n4079), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5340)
         );
  NAND2_X1 U5059 ( .A1(n5643), .A2(n5340), .ZN(n5352) );
  AND2_X1 U5060 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5750) );
  AND2_X1 U5061 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5783) );
  NAND2_X1 U5062 ( .A1(n5750), .A2(n5783), .ZN(n4105) );
  OR2_X1 U5063 ( .A1(n5650), .A2(n4105), .ZN(n4106) );
  INV_X1 U5064 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5400) );
  XNOR2_X1 U5065 ( .A(n4107), .B(n5400), .ZN(n5391) );
  AOI21_X1 U5066 ( .B1(n4173), .B2(n4130), .A(n4017), .ZN(n4109) );
  AND2_X1 U5067 ( .A1(n4108), .A2(n4109), .ZN(n4177) );
  INV_X1 U5068 ( .A(n4110), .ZN(n4111) );
  NAND2_X1 U5069 ( .A1(n4177), .A2(n4111), .ZN(n6402) );
  INV_X1 U5070 ( .A(n6166), .ZN(n6178) );
  NAND2_X1 U5071 ( .A1(n5391), .A2(n6178), .ZN(n4129) );
  AND2_X1 U5072 ( .A1(n5522), .A2(n5552), .ZN(n4113) );
  NAND2_X2 U5073 ( .A1(n5553), .A2(n4113), .ZN(n5655) );
  INV_X1 U5074 ( .A(n5655), .ZN(n4115) );
  NAND2_X1 U5075 ( .A1(n5555), .A2(n4117), .ZN(n5378) );
  NOR2_X2 U5076 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n5829) );
  NAND2_X1 U5077 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n6525), .ZN(n6432) );
  INV_X1 U5078 ( .A(n6432), .ZN(n4119) );
  NAND2_X1 U5079 ( .A1(n5829), .A2(n4119), .ZN(n6164) );
  INV_X1 U5080 ( .A(n5829), .ZN(n5838) );
  NAND2_X1 U5081 ( .A1(n5838), .A2(n4120), .ZN(n6524) );
  NAND2_X1 U5082 ( .A1(n6524), .A2(n6529), .ZN(n4121) );
  AND2_X2 U5083 ( .A1(n6166), .A2(n4121), .ZN(n6171) );
  NAND2_X1 U5084 ( .A1(n6529), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4123) );
  NAND2_X1 U5085 ( .A1(n6527), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4122) );
  AND2_X1 U5086 ( .A1(n4123), .A2(n4122), .ZN(n4208) );
  AND2_X1 U5087 ( .A1(n6189), .A2(REIP_REG_23__SCAN_IN), .ZN(n5396) );
  INV_X1 U5088 ( .A(n6171), .ZN(n5684) );
  INV_X1 U5089 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4124) );
  NOR2_X1 U5090 ( .A1(n5684), .A2(n4124), .ZN(n4125) );
  AOI211_X1 U5091 ( .C1(n5883), .C2(n5844), .A(n5396), .B(n4125), .ZN(n4126)
         );
  NAND2_X1 U5092 ( .A1(n4129), .A2(n4128), .ZN(U2963) );
  NAND2_X1 U5093 ( .A1(n5829), .A2(n4364), .ZN(n5928) );
  INV_X1 U5094 ( .A(n5928), .ZN(n4133) );
  NOR2_X1 U5095 ( .A1(n4133), .A2(READREQUEST_REG_SCAN_IN), .ZN(n4132) );
  NAND2_X1 U5096 ( .A1(n4130), .A2(n4421), .ZN(n4894) );
  NAND3_X1 U5097 ( .A1(n6523), .A2(n4246), .A3(n4894), .ZN(n4131) );
  OAI21_X1 U5098 ( .B1(n6523), .B2(n4132), .A(n4131), .ZN(U3474) );
  INV_X1 U5099 ( .A(n4263), .ZN(n4264) );
  AOI211_X1 U5100 ( .C1(MEMORYFETCH_REG_SCAN_IN), .C2(n4134), .A(n4133), .B(
        n4264), .ZN(n4135) );
  INV_X1 U5101 ( .A(n4135), .ZN(U2788) );
  INV_X1 U5102 ( .A(n4225), .ZN(n4138) );
  INV_X1 U5103 ( .A(n4157), .ZN(n4137) );
  OAI22_X1 U5104 ( .A1(n4138), .A2(n4156), .B1(n4137), .B2(n4136), .ZN(n5926)
         );
  NAND2_X1 U5105 ( .A1(n4421), .A2(n6528), .ZN(n6526) );
  OAI21_X1 U5106 ( .B1(n6526), .B2(n4460), .A(n6441), .ZN(n4139) );
  AOI21_X1 U5107 ( .B1(n3496), .B2(n6528), .A(n4139), .ZN(n4140) );
  NOR2_X1 U5108 ( .A1(n5926), .A2(n4140), .ZN(n6405) );
  OR2_X1 U5109 ( .A1(n6405), .A2(n6424), .ZN(n5932) );
  INV_X1 U5110 ( .A(n5932), .ZN(n4163) );
  INV_X1 U5111 ( .A(MORE_REG_SCAN_IN), .ZN(n4162) );
  NOR2_X1 U5112 ( .A1(n4894), .A2(n4450), .ZN(n4181) );
  OAI21_X1 U5113 ( .B1(n4181), .B2(n4220), .A(n4017), .ZN(n4143) );
  INV_X1 U5114 ( .A(n4141), .ZN(n5307) );
  NAND2_X1 U5115 ( .A1(n5307), .A2(n4450), .ZN(n4142) );
  OAI211_X1 U5116 ( .C1(n4108), .C2(n5530), .A(n4143), .B(n4142), .ZN(n4144)
         );
  INV_X1 U5117 ( .A(n4144), .ZN(n4148) );
  AND2_X1 U5118 ( .A1(n4246), .A2(n4145), .ZN(n4146) );
  OR2_X1 U5119 ( .A1(n4147), .A2(n4146), .ZN(n4178) );
  NAND2_X1 U5120 ( .A1(n4148), .A2(n4178), .ZN(n4149) );
  OR2_X1 U5121 ( .A1(n4150), .A2(n4149), .ZN(n4165) );
  NAND2_X1 U5122 ( .A1(n4197), .A2(n4151), .ZN(n4352) );
  NAND2_X1 U5123 ( .A1(n4153), .A2(n4152), .ZN(n4154) );
  NAND2_X1 U5124 ( .A1(n4352), .A2(n4154), .ZN(n4155) );
  NOR2_X1 U5125 ( .A1(n4165), .A2(n4155), .ZN(n4243) );
  NOR2_X1 U5126 ( .A1(n4173), .A2(n4171), .ZN(n4224) );
  INV_X1 U5127 ( .A(n4245), .ZN(n4335) );
  NAND2_X1 U5128 ( .A1(n4177), .A2(n4156), .ZN(n4334) );
  AND2_X1 U5129 ( .A1(n6402), .A2(n4334), .ZN(n4239) );
  NAND2_X1 U5130 ( .A1(n4239), .A2(n4157), .ZN(n4159) );
  INV_X1 U5131 ( .A(n4179), .ZN(n4158) );
  AOI22_X1 U5132 ( .A1(n4225), .A2(n4159), .B1(n4158), .B2(n4186), .ZN(n4160)
         );
  OAI21_X1 U5133 ( .B1(n4335), .B2(n4225), .A(n4160), .ZN(n6404) );
  NAND2_X1 U5134 ( .A1(n4163), .A2(n6404), .ZN(n4161) );
  OAI21_X1 U5135 ( .B1(n4163), .B2(n4162), .A(n4161), .ZN(U3471) );
  INV_X1 U5136 ( .A(n4164), .ZN(n4176) );
  INV_X1 U5137 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5698) );
  AOI22_X1 U5138 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n5698), .B2(n5157), .ZN(n6545)
         );
  NAND2_X1 U5139 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6541) );
  INV_X1 U5140 ( .A(n4201), .ZN(n6547) );
  INV_X1 U5141 ( .A(n4165), .ZN(n4170) );
  INV_X1 U5142 ( .A(n4283), .ZN(n4167) );
  AND4_X1 U5143 ( .A1(n4247), .A2(n5920), .A3(n4168), .A4(n4167), .ZN(n4169)
         );
  NAND2_X1 U5144 ( .A1(n4170), .A2(n4169), .ZN(n4355) );
  NOR2_X1 U5145 ( .A1(n4179), .A2(n4171), .ZN(n4347) );
  NAND2_X1 U5146 ( .A1(n4347), .A2(n4192), .ZN(n4348) );
  INV_X1 U5147 ( .A(n4348), .ZN(n4175) );
  INV_X1 U5148 ( .A(n4172), .ZN(n4193) );
  AOI21_X1 U5149 ( .B1(n4193), .B2(n4176), .A(n4173), .ZN(n4174) );
  AOI211_X1 U5150 ( .C1(n4495), .C2(n4355), .A(n4175), .B(n4174), .ZN(n6390)
         );
  OAI222_X1 U5151 ( .A1(n6550), .A2(n4176), .B1(n6545), .B2(n6541), .C1(n6547), 
        .C2(n6390), .ZN(n4195) );
  NAND2_X1 U5152 ( .A1(n4245), .A2(n4225), .ZN(n4218) );
  NAND2_X1 U5153 ( .A1(n4178), .A2(n4177), .ZN(n4180) );
  NAND2_X1 U5154 ( .A1(n4180), .A2(n4179), .ZN(n4228) );
  INV_X1 U5155 ( .A(n4181), .ZN(n4185) );
  INV_X1 U5156 ( .A(n6528), .ZN(n4312) );
  OAI21_X1 U5157 ( .B1(n3244), .B2(n4347), .A(n4312), .ZN(n4182) );
  OR2_X1 U5158 ( .A1(n4247), .A2(n4260), .ZN(n4265) );
  AND2_X1 U5159 ( .A1(n4182), .A2(n4265), .ZN(n4183) );
  OR3_X1 U5160 ( .A1(n4225), .A2(READY_N), .A3(n4183), .ZN(n4184) );
  NAND4_X1 U5161 ( .A1(n4218), .A2(n4228), .A3(n4185), .A4(n4184), .ZN(n4190)
         );
  OR2_X1 U5162 ( .A1(n4225), .A2(n4334), .ZN(n4189) );
  INV_X1 U5163 ( .A(n5920), .ZN(n4187) );
  NOR2_X1 U5164 ( .A1(READY_N), .A2(n4186), .ZN(n4226) );
  NAND2_X1 U5165 ( .A1(n4187), .A2(n4226), .ZN(n4188) );
  NAND2_X1 U5166 ( .A1(n4189), .A2(n4188), .ZN(n4286) );
  NOR2_X1 U5167 ( .A1(n4364), .A2(n6522), .ZN(n4367) );
  INV_X1 U5168 ( .A(n4367), .ZN(n4377) );
  NOR2_X1 U5169 ( .A1(n6529), .A2(n4377), .ZN(n6430) );
  AND2_X1 U5170 ( .A1(FLUSH_REG_SCAN_IN), .A2(n6430), .ZN(n4191) );
  AOI21_X1 U5171 ( .B1(n6391), .B2(n4284), .A(n4191), .ZN(n5921) );
  OAI21_X1 U5172 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n6512), .A(n5921), .ZN(
        n6553) );
  OAI22_X1 U5173 ( .A1(n6550), .A2(n4193), .B1(n6553), .B2(n4192), .ZN(n4194)
         );
  AOI21_X1 U5174 ( .B1(n4195), .B2(n6553), .A(n4194), .ZN(n4196) );
  INV_X1 U5175 ( .A(n4196), .ZN(U3460) );
  AOI22_X1 U5176 ( .A1(n5017), .A2(n4355), .B1(n4197), .B2(n4198), .ZN(n6387)
         );
  OAI21_X1 U5177 ( .B1(n6387), .B2(STATE2_REG_3__SCAN_IN), .A(n4364), .ZN(
        n4200) );
  INV_X1 U5178 ( .A(n6550), .ZN(n4199) );
  AOI22_X1 U5179 ( .A1(n4200), .A2(n6541), .B1(n4199), .B2(n4198), .ZN(n4204)
         );
  INV_X1 U5180 ( .A(n6553), .ZN(n4203) );
  AND2_X1 U5181 ( .A1(n4347), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6388)
         );
  AOI22_X1 U5182 ( .A1(n6388), .A2(n4201), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n4203), .ZN(n4202) );
  OAI21_X1 U5183 ( .B1(n4204), .B2(n4203), .A(n4202), .ZN(U3461) );
  XNOR2_X1 U5184 ( .A(n4205), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4256)
         );
  XNOR2_X1 U5185 ( .A(n4207), .B(n4206), .ZN(n4223) );
  INV_X2 U5186 ( .A(n6164), .ZN(n6176) );
  NAND2_X1 U5187 ( .A1(n4223), .A2(n6176), .ZN(n4211) );
  NAND2_X1 U5188 ( .A1(n5684), .A2(n4208), .ZN(n4209) );
  AOI22_X1 U5189 ( .A1(n4209), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .B1(n6018), 
        .B2(REIP_REG_0__SCAN_IN), .ZN(n4210) );
  OAI211_X1 U5190 ( .C1(n4256), .C2(n6166), .A(n4211), .B(n4210), .ZN(U2986)
         );
  INV_X1 U5191 ( .A(n4212), .ZN(n4215) );
  NOR2_X1 U5192 ( .A1(n5308), .A2(n4479), .ZN(n4213) );
  NAND4_X1 U5193 ( .A1(n4216), .A2(n4215), .A3(n4214), .A4(n4213), .ZN(n4217)
         );
  NAND2_X1 U5194 ( .A1(n4218), .A2(n4217), .ZN(n4219) );
  INV_X1 U5195 ( .A(n5308), .ZN(n5563) );
  NAND2_X1 U5196 ( .A1(n6065), .A2(n5563), .ZN(n6055) );
  NOR2_X1 U5197 ( .A1(n4220), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4221)
         );
  NOR2_X1 U5198 ( .A1(n4222), .A2(n4221), .ZN(n4254) );
  INV_X1 U5199 ( .A(n4254), .ZN(n4905) );
  AND2_X1 U5200 ( .A1(n6065), .A2(n5308), .ZN(n6061) );
  INV_X2 U5201 ( .A(n6061), .ZN(n6056) );
  INV_X1 U5202 ( .A(n4223), .ZN(n4910) );
  OAI222_X1 U5203 ( .A1(n6055), .A2(n4905), .B1(n4904), .B2(n6065), .C1(n6056), 
        .C2(n4910), .ZN(U2859) );
  NAND2_X1 U5204 ( .A1(n4225), .A2(n4224), .ZN(n4229) );
  NAND3_X1 U5205 ( .A1(n6526), .A2(n4226), .A3(n4450), .ZN(n4227) );
  NAND3_X1 U5206 ( .A1(n4229), .A2(n4228), .A3(n4227), .ZN(n4230) );
  NAND2_X1 U5207 ( .A1(n4230), .A2(n4284), .ZN(n4236) );
  NAND2_X1 U5208 ( .A1(n4231), .A2(n6441), .ZN(n4232) );
  OAI211_X1 U5209 ( .C1(n4247), .C2(n4232), .A(n4460), .B(n5307), .ZN(n4233)
         );
  INV_X1 U5210 ( .A(n4233), .ZN(n4234) );
  OR3_X1 U5211 ( .A1(n4309), .A2(n4234), .A3(n4450), .ZN(n4235) );
  OR2_X1 U5212 ( .A1(n4248), .A2(n4237), .ZN(n4238) );
  NAND4_X1 U5213 ( .A1(n4239), .A2(n5920), .A3(n4265), .A4(n4238), .ZN(n4240)
         );
  NAND2_X1 U5214 ( .A1(n4251), .A2(n4240), .ZN(n6242) );
  INV_X1 U5215 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4430) );
  NAND2_X1 U5216 ( .A1(n4283), .A2(n4241), .ZN(n4242) );
  NAND2_X1 U5217 ( .A1(n4243), .A2(n4242), .ZN(n4244) );
  NAND2_X1 U5218 ( .A1(n4251), .A2(n4244), .ZN(n5822) );
  NAND2_X1 U5219 ( .A1(n4251), .A2(n4245), .ZN(n6199) );
  NAND2_X1 U5220 ( .A1(n5822), .A2(n6199), .ZN(n5817) );
  NAND2_X1 U5221 ( .A1(n4430), .A2(n5817), .ZN(n4294) );
  OR2_X1 U5222 ( .A1(n4247), .A2(n4246), .ZN(n6416) );
  OAI21_X1 U5223 ( .B1(n4248), .B2(n4479), .A(n6416), .ZN(n4249) );
  NAND2_X1 U5224 ( .A1(n4251), .A2(n4249), .ZN(n6246) );
  INV_X1 U5225 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6518) );
  NOR2_X1 U5226 ( .A1(n4889), .A2(n6518), .ZN(n4253) );
  INV_X1 U5227 ( .A(n4251), .ZN(n4250) );
  NAND2_X1 U5228 ( .A1(n4250), .A2(n4889), .ZN(n4293) );
  NAND2_X1 U5229 ( .A1(n4251), .A2(n4347), .ZN(n5819) );
  AOI21_X1 U5230 ( .B1(n4293), .B2(n5819), .A(n4430), .ZN(n4252) );
  AOI211_X1 U5231 ( .C1(n6258), .C2(n4254), .A(n4253), .B(n4252), .ZN(n4255)
         );
  OAI211_X1 U5232 ( .C1(n4256), .C2(n6242), .A(n4294), .B(n4255), .ZN(U3018)
         );
  OAI21_X1 U5233 ( .B1(n4259), .B2(n4258), .A(n4257), .ZN(n4902) );
  XNOR2_X1 U5234 ( .A(n4261), .B(n4260), .ZN(n4895) );
  INV_X1 U5235 ( .A(n6065), .ZN(n5549) );
  AOI22_X1 U5236 ( .A1(n6060), .A2(n4895), .B1(n5549), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4262) );
  OAI21_X1 U5237 ( .B1(n4902), .B2(n6056), .A(n4262), .ZN(U2858) );
  INV_X1 U5238 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4384) );
  OAI21_X1 U5239 ( .B1(n3496), .B2(n6441), .A(n4264), .ZN(n6139) );
  INV_X1 U5240 ( .A(n6139), .ZN(n6120) );
  NAND2_X1 U5241 ( .A1(n6139), .A2(UWORD_REG_12__SCAN_IN), .ZN(n4266) );
  INV_X1 U5242 ( .A(n6143), .ZN(n6146) );
  NAND2_X1 U5243 ( .A1(n6146), .A2(DATAI_12_), .ZN(n4270) );
  OAI211_X1 U5244 ( .C1(n4384), .C2(n4311), .A(n4266), .B(n4270), .ZN(U2936)
         );
  INV_X1 U5245 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4391) );
  NAND2_X1 U5246 ( .A1(n6139), .A2(UWORD_REG_9__SCAN_IN), .ZN(n4267) );
  NAND2_X1 U5247 ( .A1(n6146), .A2(DATAI_9_), .ZN(n4273) );
  OAI211_X1 U5248 ( .C1(n4391), .C2(n4311), .A(n4267), .B(n4273), .ZN(U2933)
         );
  INV_X1 U5249 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4395) );
  NAND2_X1 U5250 ( .A1(n6145), .A2(UWORD_REG_8__SCAN_IN), .ZN(n4268) );
  NAND2_X1 U5251 ( .A1(n6146), .A2(DATAI_8_), .ZN(n4275) );
  OAI211_X1 U5252 ( .C1(n4395), .C2(n4311), .A(n4268), .B(n4275), .ZN(U2932)
         );
  INV_X1 U5253 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6088) );
  NAND2_X1 U5254 ( .A1(n6145), .A2(LWORD_REG_14__SCAN_IN), .ZN(n4269) );
  NAND2_X1 U5255 ( .A1(n6146), .A2(DATAI_14_), .ZN(n4292) );
  OAI211_X1 U5256 ( .C1(n6088), .C2(n4311), .A(n4269), .B(n4292), .ZN(U2953)
         );
  INV_X1 U5257 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6092) );
  NAND2_X1 U5258 ( .A1(n6145), .A2(LWORD_REG_12__SCAN_IN), .ZN(n4271) );
  OAI211_X1 U5259 ( .C1(n6092), .C2(n4311), .A(n4271), .B(n4270), .ZN(U2951)
         );
  INV_X1 U5260 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6090) );
  NAND2_X1 U5261 ( .A1(n6145), .A2(LWORD_REG_13__SCAN_IN), .ZN(n4272) );
  NAND2_X1 U5262 ( .A1(n6146), .A2(DATAI_13_), .ZN(n4277) );
  OAI211_X1 U5263 ( .C1(n6090), .C2(n4311), .A(n4272), .B(n4277), .ZN(U2952)
         );
  INV_X1 U5264 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6099) );
  NAND2_X1 U5265 ( .A1(n6145), .A2(LWORD_REG_9__SCAN_IN), .ZN(n4274) );
  OAI211_X1 U5266 ( .C1(n6099), .C2(n4311), .A(n4274), .B(n4273), .ZN(U2948)
         );
  INV_X1 U5267 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6101) );
  NAND2_X1 U5268 ( .A1(n6145), .A2(LWORD_REG_8__SCAN_IN), .ZN(n4276) );
  OAI211_X1 U5269 ( .C1(n6101), .C2(n4311), .A(n4276), .B(n4275), .ZN(U2947)
         );
  INV_X1 U5270 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4386) );
  NAND2_X1 U5271 ( .A1(n6145), .A2(UWORD_REG_13__SCAN_IN), .ZN(n4278) );
  OAI211_X1 U5272 ( .C1(n4386), .C2(n4311), .A(n4278), .B(n4277), .ZN(U2937)
         );
  INV_X1 U5273 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4388) );
  AOI22_X1 U5274 ( .A1(n6139), .A2(UWORD_REG_11__SCAN_IN), .B1(n6146), .B2(
        DATAI_11_), .ZN(n4279) );
  OAI21_X1 U5275 ( .B1(n4388), .B2(n4311), .A(n4279), .ZN(U2935) );
  INV_X1 U5276 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4393) );
  AOI22_X1 U5277 ( .A1(n6139), .A2(UWORD_REG_0__SCAN_IN), .B1(n6146), .B2(
        DATAI_0_), .ZN(n4280) );
  OAI21_X1 U5278 ( .B1(n4393), .B2(n4311), .A(n4280), .ZN(U2924) );
  INV_X1 U5279 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6086) );
  AOI22_X1 U5280 ( .A1(n6139), .A2(LWORD_REG_15__SCAN_IN), .B1(n6146), .B2(
        DATAI_15_), .ZN(n4281) );
  OAI21_X1 U5281 ( .B1(n6086), .B2(n4311), .A(n4281), .ZN(U2954) );
  AND3_X1 U5282 ( .A1(n4283), .A2(n5563), .A3(n4282), .ZN(n4285) );
  OAI21_X1 U5283 ( .B1(n4286), .B2(n4285), .A(n4284), .ZN(n4287) );
  NAND2_X1 U5284 ( .A1(n4288), .A2(n5308), .ZN(n4289) );
  INV_X1 U5285 ( .A(n4289), .ZN(n4290) );
  INV_X1 U5286 ( .A(n5245), .ZN(n4410) );
  INV_X1 U5287 ( .A(DATAI_0_), .ZN(n6130) );
  INV_X1 U5288 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6119) );
  OAI222_X1 U5289 ( .A1(n5877), .A2(n4910), .B1(n4410), .B2(n6130), .C1(n5562), 
        .C2(n6119), .ZN(U2891) );
  INV_X1 U5290 ( .A(DATAI_1_), .ZN(n6602) );
  INV_X1 U5291 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6114) );
  OAI222_X1 U5292 ( .A1(n4902), .A2(n5877), .B1(n4410), .B2(n6602), .C1(n5562), 
        .C2(n6114), .ZN(U2890) );
  INV_X1 U5293 ( .A(UWORD_REG_14__SCAN_IN), .ZN(n6643) );
  NAND2_X1 U5294 ( .A1(n6144), .A2(EAX_REG_30__SCAN_IN), .ZN(n4291) );
  OAI211_X1 U5295 ( .C1(n6120), .C2(n6643), .A(n4292), .B(n4291), .ZN(U2938)
         );
  NAND2_X1 U5296 ( .A1(n4294), .A2(n4293), .ZN(n5158) );
  INV_X1 U5297 ( .A(n5158), .ZN(n4301) );
  XOR2_X1 U5298 ( .A(n4296), .B(n4295), .Z(n4834) );
  NAND2_X1 U5299 ( .A1(n5771), .A2(n6199), .ZN(n6201) );
  INV_X1 U5300 ( .A(n6201), .ZN(n6203) );
  AND2_X1 U5301 ( .A1(n5819), .A2(n4430), .ZN(n4429) );
  NOR3_X1 U5302 ( .A1(n6203), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n4429), 
        .ZN(n4299) );
  INV_X1 U5303 ( .A(n4895), .ZN(n4297) );
  INV_X1 U5304 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6513) );
  OAI22_X1 U5305 ( .A1(n6246), .A2(n4297), .B1(n6513), .B2(n4889), .ZN(n4298)
         );
  AOI211_X1 U5306 ( .C1(n4834), .C2(n6263), .A(n4299), .B(n4298), .ZN(n4300)
         );
  OAI21_X1 U5307 ( .B1(n4301), .B2(n5157), .A(n4300), .ZN(U3017) );
  OAI21_X1 U5308 ( .B1(n4304), .B2(n4303), .A(n4302), .ZN(n6175) );
  XOR2_X1 U5309 ( .A(n4306), .B(n4305), .Z(n6259) );
  AOI22_X1 U5310 ( .A1(n6259), .A2(n6060), .B1(EBX_REG_2__SCAN_IN), .B2(n5549), 
        .ZN(n4307) );
  OAI21_X1 U5311 ( .B1(n6175), .B2(n6056), .A(n4307), .ZN(U2857) );
  INV_X1 U5312 ( .A(UWORD_REG_2__SCAN_IN), .ZN(n4316) );
  NOR2_X1 U5313 ( .A1(n4377), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6116) );
  INV_X1 U5314 ( .A(n6116), .ZN(n6413) );
  INV_X1 U5315 ( .A(n4347), .ZN(n4308) );
  OR2_X1 U5316 ( .A1(n4309), .A2(n4308), .ZN(n4310) );
  NAND2_X1 U5317 ( .A1(n4311), .A2(n4310), .ZN(n4313) );
  NAND2_X1 U5318 ( .A1(n6093), .A2(n4460), .ZN(n4397) );
  INV_X1 U5319 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n4314) );
  INV_X1 U5320 ( .A(n6413), .ZN(n6112) );
  OAI222_X1 U5321 ( .A1(n4316), .A2(n6413), .B1(n4397), .B2(n4315), .C1(n4314), 
        .C2(n6095), .ZN(U2905) );
  INV_X1 U5322 ( .A(n4302), .ZN(n4319) );
  INV_X1 U5323 ( .A(n4317), .ZN(n4318) );
  NAND2_X1 U5324 ( .A1(n4319), .A2(n4318), .ZN(n4398) );
  OAI21_X1 U5325 ( .B1(n4319), .B2(n4318), .A(n4398), .ZN(n6042) );
  AOI21_X1 U5326 ( .B1(n4321), .B2(n4320), .A(n5385), .ZN(n6244) );
  AOI22_X1 U5327 ( .A1(n6060), .A2(n6244), .B1(n5549), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4322) );
  OAI21_X1 U5328 ( .B1(n6042), .B2(n6056), .A(n4322), .ZN(U2856) );
  INV_X1 U5329 ( .A(DATAI_2_), .ZN(n6584) );
  INV_X1 U5330 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6111) );
  OAI222_X1 U5331 ( .A1(n6175), .A2(n5877), .B1(n4410), .B2(n6584), .C1(n5562), 
        .C2(n6111), .ZN(U2889) );
  INV_X1 U5332 ( .A(DATAI_3_), .ZN(n6134) );
  INV_X1 U5333 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6109) );
  OAI222_X1 U5334 ( .A1(n6042), .A2(n5877), .B1(n4410), .B2(n6134), .C1(n5562), 
        .C2(n6109), .ZN(U2888) );
  OAI21_X1 U5335 ( .B1(n4400), .B2(n4324), .A(n4403), .ZN(n4882) );
  NAND2_X1 U5336 ( .A1(n4325), .A2(n5387), .ZN(n4327) );
  INV_X1 U5337 ( .A(n4405), .ZN(n4326) );
  NAND2_X1 U5338 ( .A1(n4327), .A2(n4326), .ZN(n4871) );
  OAI222_X1 U5339 ( .A1(n4882), .A2(n6056), .B1(n4328), .B2(n6065), .C1(n4871), 
        .C2(n6055), .ZN(U2854) );
  INV_X1 U5340 ( .A(DATAI_5_), .ZN(n6137) );
  INV_X1 U5341 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6105) );
  OAI222_X1 U5342 ( .A1(n4882), .A2(n5877), .B1(n4410), .B2(n6137), .C1(n5562), 
        .C2(n6105), .ZN(U2886) );
  INV_X1 U5343 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n4330) );
  INV_X1 U5344 ( .A(n4397), .ZN(n6083) );
  AOI22_X1 U5345 ( .A1(n6083), .A2(EAX_REG_20__SCAN_IN), .B1(n6112), .B2(
        UWORD_REG_4__SCAN_IN), .ZN(n4329) );
  OAI21_X1 U5346 ( .B1(n6095), .B2(n4330), .A(n4329), .ZN(U2903) );
  NOR2_X1 U5347 ( .A1(FLUSH_REG_SCAN_IN), .A2(n4364), .ZN(n4363) );
  AOI21_X1 U5348 ( .B1(n6549), .B2(n6552), .A(n4344), .ZN(n4332) );
  NOR2_X1 U5349 ( .A1(n2957), .A2(n4332), .ZN(n5841) );
  MUX2_X1 U5350 ( .A(n4333), .B(n4344), .S(n6549), .Z(n4336) );
  NAND2_X1 U5351 ( .A1(n4335), .A2(n4334), .ZN(n4346) );
  OAI21_X1 U5352 ( .B1(n4337), .B2(n4336), .A(n4346), .ZN(n4342) );
  NAND2_X1 U5353 ( .A1(n6552), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4338) );
  INV_X1 U5354 ( .A(n4338), .ZN(n4339) );
  MUX2_X1 U5355 ( .A(n4339), .B(n4338), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4340) );
  NAND2_X1 U5356 ( .A1(n4347), .A2(n4340), .ZN(n4341) );
  OAI211_X1 U5357 ( .C1(n5841), .C2(n4352), .A(n4342), .B(n4341), .ZN(n4343)
         );
  AOI21_X1 U5358 ( .B1(n6038), .B2(n4355), .A(n4343), .ZN(n5842) );
  MUX2_X1 U5359 ( .A(n4344), .B(n5842), .S(n6391), .Z(n6401) );
  XNOR2_X1 U5360 ( .A(n6549), .B(n6552), .ZN(n4353) );
  NAND2_X1 U5361 ( .A1(n4346), .A2(n4353), .ZN(n4351) );
  NAND2_X1 U5362 ( .A1(n4347), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4349) );
  MUX2_X1 U5363 ( .A(n4349), .B(n4348), .S(n6552), .Z(n4350) );
  OAI211_X1 U5364 ( .C1(n4353), .C2(n4352), .A(n4351), .B(n4350), .ZN(n4354)
         );
  AOI21_X1 U5365 ( .B1(n5117), .B2(n4355), .A(n4354), .ZN(n6548) );
  NOR2_X1 U5366 ( .A1(n6391), .A2(n6552), .ZN(n4356) );
  AOI21_X1 U5367 ( .B1(n6548), .B2(n6391), .A(n4356), .ZN(n6398) );
  INV_X1 U5368 ( .A(n6398), .ZN(n4357) );
  NOR3_X1 U5369 ( .A1(n6401), .A2(n4357), .A3(STATE2_REG_1__SCAN_IN), .ZN(
        n4358) );
  AOI21_X1 U5370 ( .B1(n4363), .B2(n4359), .A(n4358), .ZN(n6409) );
  INV_X1 U5371 ( .A(n4716), .ZN(n4360) );
  NOR2_X1 U5372 ( .A1(n4361), .A2(n4360), .ZN(n4362) );
  XNOR2_X1 U5373 ( .A(n4362), .B(n5924), .ZN(n6019) );
  INV_X1 U5374 ( .A(n6019), .ZN(n5922) );
  OAI22_X1 U5375 ( .A1(n5922), .A2(n5920), .B1(n5924), .B2(n6391), .ZN(n4365)
         );
  AOI22_X1 U5376 ( .A1(n4365), .A2(n4364), .B1(n4363), .B2(
        INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6408) );
  OAI21_X1 U5377 ( .B1(n6409), .B2(n4366), .A(n6408), .ZN(n4378) );
  OAI21_X1 U5378 ( .B1(n4378), .B2(FLUSH_REG_SCAN_IN), .A(n6430), .ZN(n4368)
         );
  NAND2_X1 U5379 ( .A1(n4368), .A2(n4754), .ZN(n6268) );
  AND2_X1 U5380 ( .A1(n4600), .A2(n4626), .ZN(n4370) );
  AND2_X1 U5381 ( .A1(n5835), .A2(n4370), .ZN(n4562) );
  NAND2_X1 U5382 ( .A1(n4562), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4556) );
  INV_X1 U5383 ( .A(n5835), .ZN(n4590) );
  NAND2_X1 U5384 ( .A1(n4590), .A2(n4749), .ZN(n4527) );
  NAND2_X1 U5385 ( .A1(n4556), .A2(n4527), .ZN(n4592) );
  INV_X1 U5386 ( .A(n4592), .ZN(n4372) );
  NAND2_X1 U5387 ( .A1(n4723), .A2(n5834), .ZN(n4806) );
  AOI21_X1 U5388 ( .B1(n4372), .B2(n4806), .A(n5838), .ZN(n4375) );
  INV_X1 U5389 ( .A(n4749), .ZN(n4373) );
  NAND2_X1 U5390 ( .A1(n5829), .A2(n6527), .ZN(n5169) );
  AND2_X1 U5391 ( .A1(n6512), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5836) );
  OAI22_X1 U5392 ( .A1(n4373), .A2(n5169), .B1(n5064), .B2(n5836), .ZN(n4374)
         );
  OAI21_X1 U5393 ( .B1(n4375), .B2(n4374), .A(n6268), .ZN(n4376) );
  OAI21_X1 U5394 ( .B1(n6268), .B2(n4970), .A(n4376), .ZN(U3462) );
  NOR2_X1 U5395 ( .A1(n4378), .A2(n4377), .ZN(n6419) );
  OAI22_X1 U5396 ( .A1(n5026), .A2(n5838), .B1(n4903), .B2(n5836), .ZN(n4379)
         );
  OAI21_X1 U5397 ( .B1(n6419), .B2(n4379), .A(n6268), .ZN(n4380) );
  OAI21_X1 U5398 ( .B1(n6268), .B2(n6691), .A(n4380), .ZN(U3465) );
  INV_X1 U5399 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4382) );
  INV_X2 U5400 ( .A(n6095), .ZN(n6115) );
  AOI22_X1 U5401 ( .A1(n6112), .A2(UWORD_REG_10__SCAN_IN), .B1(n6115), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4381) );
  OAI21_X1 U5402 ( .B1(n4382), .B2(n4397), .A(n4381), .ZN(U2897) );
  AOI22_X1 U5403 ( .A1(n6112), .A2(UWORD_REG_12__SCAN_IN), .B1(n6115), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4383) );
  OAI21_X1 U5404 ( .B1(n4384), .B2(n4397), .A(n4383), .ZN(U2895) );
  AOI22_X1 U5405 ( .A1(n6112), .A2(UWORD_REG_13__SCAN_IN), .B1(n6115), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4385) );
  OAI21_X1 U5406 ( .B1(n4386), .B2(n4397), .A(n4385), .ZN(U2894) );
  AOI22_X1 U5407 ( .A1(n6112), .A2(UWORD_REG_11__SCAN_IN), .B1(n6115), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4387) );
  OAI21_X1 U5408 ( .B1(n4388), .B2(n4397), .A(n4387), .ZN(U2896) );
  AOI22_X1 U5409 ( .A1(n6116), .A2(UWORD_REG_7__SCAN_IN), .B1(n6115), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4389) );
  OAI21_X1 U5410 ( .B1(n3372), .B2(n4397), .A(n4389), .ZN(U2900) );
  AOI22_X1 U5411 ( .A1(n6116), .A2(UWORD_REG_9__SCAN_IN), .B1(n6115), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4390) );
  OAI21_X1 U5412 ( .B1(n4391), .B2(n4397), .A(n4390), .ZN(U2898) );
  AOI22_X1 U5413 ( .A1(n6116), .A2(UWORD_REG_0__SCAN_IN), .B1(n6115), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4392) );
  OAI21_X1 U5414 ( .B1(n4393), .B2(n4397), .A(n4392), .ZN(U2907) );
  AOI22_X1 U5415 ( .A1(n6116), .A2(UWORD_REG_8__SCAN_IN), .B1(n6115), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4394) );
  OAI21_X1 U5416 ( .B1(n4395), .B2(n4397), .A(n4394), .ZN(U2899) );
  AOI22_X1 U5417 ( .A1(n6116), .A2(UWORD_REG_3__SCAN_IN), .B1(n6115), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4396) );
  OAI21_X1 U5418 ( .B1(n3442), .B2(n4397), .A(n4396), .ZN(U2904) );
  AND2_X1 U5419 ( .A1(n4399), .A2(n4398), .ZN(n4401) );
  OR2_X1 U5420 ( .A1(n4401), .A2(n4400), .ZN(n6165) );
  INV_X1 U5421 ( .A(DATAI_4_), .ZN(n6634) );
  INV_X1 U5422 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6107) );
  OAI222_X1 U5423 ( .A1(n6165), .A2(n5877), .B1(n4410), .B2(n6634), .C1(n5562), 
        .C2(n6107), .ZN(U2887) );
  NAND2_X1 U5424 ( .A1(n4403), .A2(n4402), .ZN(n4404) );
  AND2_X1 U5425 ( .A1(n4518), .A2(n4404), .ZN(n6156) );
  INV_X1 U5426 ( .A(n6156), .ZN(n4411) );
  OR2_X1 U5427 ( .A1(n4406), .A2(n4405), .ZN(n4407) );
  NAND2_X1 U5428 ( .A1(n4407), .A2(n4521), .ZN(n6004) );
  INV_X1 U5429 ( .A(n6004), .ZN(n4408) );
  AOI22_X1 U5430 ( .A1(n6060), .A2(n4408), .B1(n5549), .B2(EBX_REG_6__SCAN_IN), 
        .ZN(n4409) );
  OAI21_X1 U5431 ( .B1(n4411), .B2(n6056), .A(n4409), .ZN(U2853) );
  INV_X1 U5432 ( .A(DATAI_6_), .ZN(n6600) );
  OAI222_X1 U5433 ( .A1(n4411), .A2(n5877), .B1(n4410), .B2(n6600), .C1(n5562), 
        .C2(n3728), .ZN(U2885) );
  NAND3_X1 U5434 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6399), .ZN(n4974) );
  INV_X1 U5435 ( .A(n4527), .ZN(n4412) );
  NAND2_X1 U5436 ( .A1(n4412), .A2(n5834), .ZN(n4417) );
  INV_X1 U5437 ( .A(n4495), .ZN(n5831) );
  NOR2_X1 U5438 ( .A1(n5117), .A2(n5831), .ZN(n4593) );
  AND2_X1 U5439 ( .A1(n4593), .A2(n6038), .ZN(n4972) );
  INV_X1 U5440 ( .A(n4972), .ZN(n4975) );
  INV_X1 U5441 ( .A(n4594), .ZN(n4413) );
  NAND2_X1 U5442 ( .A1(n4413), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6375) );
  OAI21_X1 U5443 ( .B1(n4975), .B2(n4903), .A(n6375), .ZN(n4415) );
  NAND3_X1 U5444 ( .A1(n4417), .A2(n5829), .A3(n4415), .ZN(n4414) );
  OAI21_X1 U5445 ( .B1(n4974), .B2(n6522), .A(n4414), .ZN(n6380) );
  INV_X1 U5446 ( .A(n6380), .ZN(n4425) );
  NOR2_X1 U5447 ( .A1(n6602), .A2(n4754), .ZN(n6318) );
  INV_X1 U5448 ( .A(n6318), .ZN(n5198) );
  INV_X1 U5449 ( .A(n4974), .ZN(n4419) );
  INV_X1 U5450 ( .A(n4415), .ZN(n4416) );
  NAND3_X1 U5451 ( .A1(n4417), .A2(n5829), .A3(n4416), .ZN(n4418) );
  AOI21_X1 U5452 ( .B1(n6691), .B2(STATE2_REG_3__SCAN_IN), .A(n4754), .ZN(
        n5021) );
  OAI211_X1 U5453 ( .C1(n5829), .C2(n4419), .A(n4418), .B(n5021), .ZN(n6382)
         );
  NAND2_X1 U5454 ( .A1(n5830), .A2(n5026), .ZN(n4493) );
  NAND2_X1 U5455 ( .A1(n6176), .A2(DATAI_25_), .ZN(n6321) );
  NAND2_X1 U5456 ( .A1(n4484), .A2(n4421), .ZN(n6315) );
  OAI22_X1 U5457 ( .A1(n6385), .A2(n6321), .B1(n6315), .B2(n6375), .ZN(n4423)
         );
  OR2_X1 U5458 ( .A1(n4527), .A2(n5026), .ZN(n4525) );
  NAND2_X1 U5459 ( .A1(n6176), .A2(DATAI_17_), .ZN(n6316) );
  NOR2_X1 U5460 ( .A1(n6378), .A2(n6316), .ZN(n4422) );
  AOI211_X1 U5461 ( .C1(INSTQUEUE_REG_11__1__SCAN_IN), .C2(n6382), .A(n4423), 
        .B(n4422), .ZN(n4424) );
  OAI21_X1 U5462 ( .B1(n4425), .B2(n5198), .A(n4424), .ZN(U3109) );
  OAI21_X1 U5463 ( .B1(n4428), .B2(n4427), .A(n4426), .ZN(n4624) );
  INV_X1 U5464 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6252) );
  NOR2_X1 U5465 ( .A1(n6252), .A2(n6241), .ZN(n6234) );
  NAND3_X1 U5466 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n6254), .ZN(n5161) );
  INV_X1 U5467 ( .A(n5161), .ZN(n4883) );
  NAND3_X1 U5468 ( .A1(n6234), .A2(n4883), .A3(n4432), .ZN(n4438) );
  INV_X1 U5469 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6257) );
  OAI21_X1 U5470 ( .B1(n5157), .B2(n4430), .A(n6257), .ZN(n6255) );
  NAND2_X1 U5471 ( .A1(n6234), .A2(n6255), .ZN(n4433) );
  NOR2_X1 U5472 ( .A1(n6257), .A2(n5157), .ZN(n4431) );
  NAND2_X1 U5473 ( .A1(n6199), .A2(n5158), .ZN(n5769) );
  OAI21_X1 U5474 ( .B1(n5771), .B2(n4431), .A(n5769), .ZN(n6262) );
  AOI221_X1 U5475 ( .B1(n4432), .B2(n6201), .C1(n4433), .C2(n6201), .A(n6262), 
        .ZN(n4884) );
  INV_X1 U5476 ( .A(n4884), .ZN(n4436) );
  OAI21_X1 U5477 ( .B1(n6199), .B2(n4433), .A(n4432), .ZN(n4435) );
  OAI22_X1 U5478 ( .A1(n6246), .A2(n4871), .B1(n6457), .B2(n4889), .ZN(n4434)
         );
  AOI21_X1 U5479 ( .B1(n4436), .B2(n4435), .A(n4434), .ZN(n4437) );
  OAI211_X1 U5480 ( .C1(n4624), .C2(n6242), .A(n4438), .B(n4437), .ZN(U3013)
         );
  NAND2_X1 U5481 ( .A1(n4723), .A2(n4631), .ZN(n4492) );
  NOR2_X1 U5482 ( .A1(n5830), .A2(n4631), .ZN(n4722) );
  INV_X1 U5483 ( .A(n4722), .ZN(n4439) );
  OR2_X1 U5484 ( .A1(n4527), .A2(n4439), .ZN(n4534) );
  NAND3_X1 U5485 ( .A1(n6326), .A2(n5829), .A3(n4534), .ZN(n4440) );
  NOR2_X1 U5486 ( .A1(n5117), .A2(n4495), .ZN(n4752) );
  AND2_X1 U5487 ( .A1(n4752), .A2(n6038), .ZN(n4444) );
  AOI21_X1 U5488 ( .B1(n4440), .B2(n5169), .A(n4444), .ZN(n4443) );
  NAND3_X1 U5489 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6399), .A3(n6393), .ZN(n4531) );
  NOR2_X1 U5490 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4531), .ZN(n4485)
         );
  AND2_X1 U5491 ( .A1(n4447), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5063) );
  INV_X1 U5492 ( .A(n5063), .ZN(n4916) );
  INV_X1 U5493 ( .A(n4753), .ZN(n4441) );
  OR2_X1 U5494 ( .A1(n4441), .A2(n5177), .ZN(n4446) );
  AOI21_X1 U5495 ( .B1(n4446), .B2(STATE2_REG_2__SCAN_IN), .A(n4754), .ZN(
        n4682) );
  OAI211_X1 U5496 ( .C1(n6512), .C2(n4485), .A(n4916), .B(n4682), .ZN(n4442)
         );
  NAND2_X1 U5497 ( .A1(n6176), .A2(DATAI_26_), .ZN(n6346) );
  NOR2_X1 U5498 ( .A1(n6584), .A2(n4754), .ZN(n6343) );
  INV_X1 U5499 ( .A(n4444), .ZN(n4445) );
  OR2_X1 U5500 ( .A1(n4445), .A2(n5838), .ZN(n4449) );
  INV_X1 U5501 ( .A(n4446), .ZN(n4685) );
  NOR2_X1 U5502 ( .A1(n4447), .A2(n6522), .ZN(n5058) );
  NAND2_X1 U5503 ( .A1(n4685), .A2(n5058), .ZN(n4448) );
  NAND2_X1 U5504 ( .A1(n4449), .A2(n4448), .ZN(n4486) );
  NAND2_X1 U5505 ( .A1(n4484), .A2(n4450), .ZN(n6340) );
  INV_X1 U5506 ( .A(n6340), .ZN(n6300) );
  AOI22_X1 U5507 ( .A1(n6343), .A2(n4486), .B1(n6300), .B2(n4485), .ZN(n4452)
         );
  NAND2_X1 U5508 ( .A1(n6176), .A2(DATAI_18_), .ZN(n6341) );
  OR2_X1 U5509 ( .A1(n4534), .A2(n6341), .ZN(n4451) );
  OAI211_X1 U5510 ( .C1(n6326), .C2(n6346), .A(n4452), .B(n4451), .ZN(n4453)
         );
  AOI21_X1 U5511 ( .B1(n4490), .B2(INSTQUEUE_REG_8__2__SCAN_IN), .A(n4453), 
        .ZN(n4454) );
  INV_X1 U5512 ( .A(n4454), .ZN(U3086) );
  NAND2_X1 U5513 ( .A1(n6176), .A2(DATAI_30_), .ZN(n6374) );
  NOR2_X1 U5514 ( .A1(n6600), .A2(n4754), .ZN(n6371) );
  NAND2_X1 U5515 ( .A1(n4484), .A2(n4455), .ZN(n6368) );
  INV_X1 U5516 ( .A(n6368), .ZN(n6279) );
  AOI22_X1 U5517 ( .A1(n6371), .A2(n4486), .B1(n6279), .B2(n4485), .ZN(n4457)
         );
  NAND2_X1 U5518 ( .A1(n6176), .A2(DATAI_22_), .ZN(n6369) );
  OR2_X1 U5519 ( .A1(n4534), .A2(n6369), .ZN(n4456) );
  OAI211_X1 U5520 ( .C1(n6326), .C2(n6374), .A(n4457), .B(n4456), .ZN(n4458)
         );
  AOI21_X1 U5521 ( .B1(n4490), .B2(INSTQUEUE_REG_8__6__SCAN_IN), .A(n4458), 
        .ZN(n4459) );
  INV_X1 U5522 ( .A(n4459), .ZN(U3090) );
  NAND2_X1 U5523 ( .A1(n6176), .A2(DATAI_24_), .ZN(n6339) );
  NOR2_X1 U5524 ( .A1(n6130), .A2(n4754), .ZN(n6336) );
  NAND2_X1 U5525 ( .A1(n4484), .A2(n4460), .ZN(n6333) );
  INV_X1 U5526 ( .A(n6333), .ZN(n6292) );
  AOI22_X1 U5527 ( .A1(n6336), .A2(n4486), .B1(n6292), .B2(n4485), .ZN(n4462)
         );
  NAND2_X1 U5528 ( .A1(n6176), .A2(DATAI_16_), .ZN(n6334) );
  OR2_X1 U5529 ( .A1(n4534), .A2(n6334), .ZN(n4461) );
  OAI211_X1 U5530 ( .C1(n6326), .C2(n6339), .A(n4462), .B(n4461), .ZN(n4463)
         );
  AOI21_X1 U5531 ( .B1(n4490), .B2(INSTQUEUE_REG_8__0__SCAN_IN), .A(n4463), 
        .ZN(n4464) );
  INV_X1 U5532 ( .A(n4464), .ZN(U3084) );
  NAND2_X1 U5533 ( .A1(n6176), .A2(DATAI_27_), .ZN(n6353) );
  NOR2_X1 U5534 ( .A1(n6134), .A2(n4754), .ZN(n6350) );
  NAND2_X1 U5535 ( .A1(n4484), .A2(n4465), .ZN(n6347) );
  INV_X1 U5536 ( .A(n6347), .ZN(n6305) );
  AOI22_X1 U5537 ( .A1(n6350), .A2(n4486), .B1(n6305), .B2(n4485), .ZN(n4467)
         );
  NAND2_X1 U5538 ( .A1(n6176), .A2(DATAI_19_), .ZN(n6348) );
  OR2_X1 U5539 ( .A1(n4534), .A2(n6348), .ZN(n4466) );
  OAI211_X1 U5540 ( .C1(n6326), .C2(n6353), .A(n4467), .B(n4466), .ZN(n4468)
         );
  AOI21_X1 U5541 ( .B1(n4490), .B2(INSTQUEUE_REG_8__3__SCAN_IN), .A(n4468), 
        .ZN(n4469) );
  INV_X1 U5542 ( .A(n4469), .ZN(U3087) );
  INV_X1 U5543 ( .A(n6315), .ZN(n6296) );
  AOI22_X1 U5544 ( .A1(n6318), .A2(n4486), .B1(n6296), .B2(n4485), .ZN(n4471)
         );
  OR2_X1 U5545 ( .A1(n4534), .A2(n6316), .ZN(n4470) );
  OAI211_X1 U5546 ( .C1(n6326), .C2(n6321), .A(n4471), .B(n4470), .ZN(n4472)
         );
  AOI21_X1 U5547 ( .B1(n4490), .B2(INSTQUEUE_REG_8__1__SCAN_IN), .A(n4472), 
        .ZN(n4473) );
  INV_X1 U5548 ( .A(n4473), .ZN(U3085) );
  NAND2_X1 U5549 ( .A1(n6176), .A2(DATAI_29_), .ZN(n6367) );
  NOR2_X1 U5550 ( .A1(n6137), .A2(n4754), .ZN(n6364) );
  NAND2_X1 U5551 ( .A1(n4484), .A2(n4474), .ZN(n6361) );
  INV_X1 U5552 ( .A(n6361), .ZN(n5039) );
  AOI22_X1 U5553 ( .A1(n6364), .A2(n4486), .B1(n5039), .B2(n4485), .ZN(n4476)
         );
  NAND2_X1 U5554 ( .A1(n6176), .A2(DATAI_21_), .ZN(n6362) );
  OR2_X1 U5555 ( .A1(n4534), .A2(n6362), .ZN(n4475) );
  OAI211_X1 U5556 ( .C1(n6326), .C2(n6367), .A(n4476), .B(n4475), .ZN(n4477)
         );
  AOI21_X1 U5557 ( .B1(n4490), .B2(INSTQUEUE_REG_8__5__SCAN_IN), .A(n4477), 
        .ZN(n4478) );
  INV_X1 U5558 ( .A(n4478), .ZN(U3089) );
  NAND2_X1 U5559 ( .A1(n6176), .A2(DATAI_28_), .ZN(n6360) );
  NOR2_X1 U5560 ( .A1(n6634), .A2(n4754), .ZN(n6357) );
  NAND2_X1 U5561 ( .A1(n4484), .A2(n4479), .ZN(n6354) );
  INV_X1 U5562 ( .A(n6354), .ZN(n6275) );
  AOI22_X1 U5563 ( .A1(n6357), .A2(n4486), .B1(n6275), .B2(n4485), .ZN(n4481)
         );
  NAND2_X1 U5564 ( .A1(n6176), .A2(DATAI_20_), .ZN(n6355) );
  OR2_X1 U5565 ( .A1(n4534), .A2(n6355), .ZN(n4480) );
  OAI211_X1 U5566 ( .C1(n6326), .C2(n6360), .A(n4481), .B(n4480), .ZN(n4482)
         );
  AOI21_X1 U5567 ( .B1(n4490), .B2(INSTQUEUE_REG_8__4__SCAN_IN), .A(n4482), 
        .ZN(n4483) );
  INV_X1 U5568 ( .A(n4483), .ZN(U3088) );
  NAND2_X1 U5569 ( .A1(n6176), .A2(DATAI_31_), .ZN(n6386) );
  INV_X1 U5570 ( .A(DATAI_7_), .ZN(n6141) );
  NOR2_X1 U5571 ( .A1(n6141), .A2(n4754), .ZN(n6381) );
  NAND2_X1 U5572 ( .A1(n4484), .A2(n5308), .ZN(n6376) );
  INV_X1 U5573 ( .A(n6376), .ZN(n6284) );
  AOI22_X1 U5574 ( .A1(n6381), .A2(n4486), .B1(n6284), .B2(n4485), .ZN(n4488)
         );
  NAND2_X1 U5575 ( .A1(n6176), .A2(DATAI_23_), .ZN(n6377) );
  OR2_X1 U5576 ( .A1(n4534), .A2(n6377), .ZN(n4487) );
  OAI211_X1 U5577 ( .C1(n6326), .C2(n6386), .A(n4488), .B(n4487), .ZN(n4489)
         );
  AOI21_X1 U5578 ( .B1(n4490), .B2(INSTQUEUE_REG_8__7__SCAN_IN), .A(n4489), 
        .ZN(n4491) );
  INV_X1 U5579 ( .A(n4491), .ZN(U3091) );
  INV_X1 U5580 ( .A(n4493), .ZN(n4494) );
  NAND2_X1 U5581 ( .A1(n4723), .A2(n4494), .ZN(n6332) );
  AOI21_X1 U5582 ( .B1(n4721), .B2(n6332), .A(n6527), .ZN(n4500) );
  NAND2_X1 U5583 ( .A1(n5117), .A2(n4495), .ZN(n4923) );
  OR2_X1 U5584 ( .A1(n4923), .A2(n4716), .ZN(n4807) );
  NAND2_X1 U5585 ( .A1(n4807), .A2(n5829), .ZN(n4499) );
  INV_X1 U5586 ( .A(n4754), .ZN(n4496) );
  OAI21_X1 U5587 ( .B1(n5177), .B2(n6522), .A(n4496), .ZN(n4973) );
  NOR2_X1 U5588 ( .A1(n5058), .A2(n4973), .ZN(n4927) );
  NOR2_X1 U5589 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4809), .ZN(n6304)
         );
  OAI21_X1 U5590 ( .B1(n6512), .B2(n6304), .A(n4970), .ZN(n4497) );
  INV_X1 U5591 ( .A(n4497), .ZN(n4498) );
  OAI211_X1 U5592 ( .C1(n4500), .C2(n4499), .A(n4927), .B(n4498), .ZN(n6309)
         );
  OR2_X1 U5593 ( .A1(n4923), .A2(n5838), .ZN(n4915) );
  NAND3_X1 U5594 ( .A1(n5063), .A2(n5177), .A3(n4970), .ZN(n4501) );
  OAI21_X1 U5595 ( .B1(n4915), .B2(n6038), .A(n4501), .ZN(n6306) );
  AOI22_X1 U5596 ( .A1(n6371), .A2(n6306), .B1(n6279), .B2(n6304), .ZN(n4503)
         );
  OR2_X1 U5597 ( .A1(n6332), .A2(n6369), .ZN(n4502) );
  OAI211_X1 U5598 ( .C1(n4721), .C2(n6374), .A(n4503), .B(n4502), .ZN(n4504)
         );
  AOI21_X1 U5599 ( .B1(n6309), .B2(INSTQUEUE_REG_6__6__SCAN_IN), .A(n4504), 
        .ZN(n4505) );
  INV_X1 U5600 ( .A(n4505), .ZN(U3074) );
  AOI22_X1 U5601 ( .A1(n6381), .A2(n6306), .B1(n6284), .B2(n6304), .ZN(n4507)
         );
  OR2_X1 U5602 ( .A1(n6332), .A2(n6377), .ZN(n4506) );
  OAI211_X1 U5603 ( .C1(n4721), .C2(n6386), .A(n4507), .B(n4506), .ZN(n4508)
         );
  AOI21_X1 U5604 ( .B1(n6309), .B2(INSTQUEUE_REG_6__7__SCAN_IN), .A(n4508), 
        .ZN(n4509) );
  INV_X1 U5605 ( .A(n4509), .ZN(U3075) );
  AOI22_X1 U5606 ( .A1(n6364), .A2(n6306), .B1(n5039), .B2(n6304), .ZN(n4511)
         );
  OR2_X1 U5607 ( .A1(n6332), .A2(n6362), .ZN(n4510) );
  OAI211_X1 U5608 ( .C1(n4721), .C2(n6367), .A(n4511), .B(n4510), .ZN(n4512)
         );
  AOI21_X1 U5609 ( .B1(n6309), .B2(INSTQUEUE_REG_6__5__SCAN_IN), .A(n4512), 
        .ZN(n4513) );
  INV_X1 U5610 ( .A(n4513), .ZN(U3073) );
  AOI22_X1 U5611 ( .A1(n6357), .A2(n6306), .B1(n6275), .B2(n6304), .ZN(n4515)
         );
  OR2_X1 U5612 ( .A1(n6332), .A2(n6355), .ZN(n4514) );
  OAI211_X1 U5613 ( .C1(n4721), .C2(n6360), .A(n4515), .B(n4514), .ZN(n4516)
         );
  AOI21_X1 U5614 ( .B1(n6309), .B2(INSTQUEUE_REG_6__4__SCAN_IN), .A(n4516), 
        .ZN(n4517) );
  INV_X1 U5615 ( .A(n4517), .ZN(U3072) );
  XOR2_X1 U5616 ( .A(n4519), .B(n4518), .Z(n4804) );
  INV_X1 U5617 ( .A(n4804), .ZN(n4859) );
  AOI21_X1 U5618 ( .B1(n4522), .B2(n4521), .A(n4616), .ZN(n6225) );
  AOI22_X1 U5619 ( .A1(n6060), .A2(n6225), .B1(n5549), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n4523) );
  OAI21_X1 U5620 ( .B1(n4859), .B2(n6056), .A(n4523), .ZN(U2852) );
  INV_X2 U5621 ( .A(n5562), .ZN(n6076) );
  AOI22_X1 U5622 ( .A1(n5245), .A2(DATAI_7_), .B1(n6076), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n4524) );
  OAI21_X1 U5623 ( .B1(n4859), .B2(n5877), .A(n4524), .ZN(U2884) );
  NOR2_X1 U5624 ( .A1(n5830), .A2(n6527), .ZN(n4715) );
  INV_X1 U5625 ( .A(n4715), .ZN(n4526) );
  OR2_X1 U5626 ( .A1(n4527), .A2(n4526), .ZN(n4528) );
  NAND2_X1 U5627 ( .A1(n6038), .A2(n5017), .ZN(n4625) );
  INV_X1 U5628 ( .A(n4625), .ZN(n4555) );
  NOR2_X1 U5629 ( .A1(n6691), .A2(n4531), .ZN(n4551) );
  AOI21_X1 U5630 ( .B1(n4555), .B2(n4752), .A(n4551), .ZN(n4533) );
  AOI22_X1 U5631 ( .A1(n4530), .A2(n4533), .B1(n5838), .B2(n4531), .ZN(n4529)
         );
  NAND2_X1 U5632 ( .A1(n5021), .A2(n4529), .ZN(n4550) );
  INV_X1 U5633 ( .A(n4530), .ZN(n4532) );
  OAI22_X1 U5634 ( .A1(n4533), .A2(n4532), .B1(n6522), .B2(n4531), .ZN(n4549)
         );
  AOI22_X1 U5635 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4550), .B1(n6371), 
        .B2(n4549), .ZN(n4536) );
  INV_X1 U5636 ( .A(n6374), .ZN(n5217) );
  AOI22_X1 U5637 ( .A1(n4552), .A2(n5217), .B1(n6279), .B2(n4551), .ZN(n4535)
         );
  OAI211_X1 U5638 ( .C1(n4978), .C2(n6369), .A(n4536), .B(n4535), .ZN(U3098)
         );
  AOI22_X1 U5639 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4550), .B1(n6336), 
        .B2(n4549), .ZN(n4538) );
  INV_X1 U5640 ( .A(n6339), .ZN(n6293) );
  AOI22_X1 U5641 ( .A1(n4552), .A2(n6293), .B1(n6292), .B2(n4551), .ZN(n4537)
         );
  OAI211_X1 U5642 ( .C1(n4978), .C2(n6334), .A(n4538), .B(n4537), .ZN(U3092)
         );
  AOI22_X1 U5643 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4550), .B1(n6318), 
        .B2(n4549), .ZN(n4540) );
  INV_X1 U5644 ( .A(n6321), .ZN(n6297) );
  AOI22_X1 U5645 ( .A1(n4552), .A2(n6297), .B1(n6296), .B2(n4551), .ZN(n4539)
         );
  OAI211_X1 U5646 ( .C1(n4978), .C2(n6316), .A(n4540), .B(n4539), .ZN(U3093)
         );
  AOI22_X1 U5647 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4550), .B1(n6381), 
        .B2(n4549), .ZN(n4542) );
  INV_X1 U5648 ( .A(n6386), .ZN(n5208) );
  AOI22_X1 U5649 ( .A1(n4552), .A2(n5208), .B1(n6284), .B2(n4551), .ZN(n4541)
         );
  OAI211_X1 U5650 ( .C1(n4978), .C2(n6377), .A(n4542), .B(n4541), .ZN(U3099)
         );
  AOI22_X1 U5651 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4550), .B1(n6357), 
        .B2(n4549), .ZN(n4544) );
  INV_X1 U5652 ( .A(n6360), .ZN(n5187) );
  AOI22_X1 U5653 ( .A1(n4552), .A2(n5187), .B1(n6275), .B2(n4551), .ZN(n4543)
         );
  OAI211_X1 U5654 ( .C1(n4978), .C2(n6355), .A(n4544), .B(n4543), .ZN(U3096)
         );
  AOI22_X1 U5655 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4550), .B1(n6343), 
        .B2(n4549), .ZN(n4546) );
  INV_X1 U5656 ( .A(n6346), .ZN(n6301) );
  AOI22_X1 U5657 ( .A1(n4552), .A2(n6301), .B1(n6300), .B2(n4551), .ZN(n4545)
         );
  OAI211_X1 U5658 ( .C1(n4978), .C2(n6341), .A(n4546), .B(n4545), .ZN(U3094)
         );
  AOI22_X1 U5659 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4550), .B1(n6364), 
        .B2(n4549), .ZN(n4548) );
  INV_X1 U5660 ( .A(n6367), .ZN(n5182) );
  AOI22_X1 U5661 ( .A1(n4552), .A2(n5182), .B1(n5039), .B2(n4551), .ZN(n4547)
         );
  OAI211_X1 U5662 ( .C1(n4978), .C2(n6362), .A(n4548), .B(n4547), .ZN(U3097)
         );
  AOI22_X1 U5663 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4550), .B1(n6350), 
        .B2(n4549), .ZN(n4554) );
  INV_X1 U5664 ( .A(n6353), .ZN(n6308) );
  AOI22_X1 U5665 ( .A1(n4552), .A2(n6308), .B1(n6305), .B2(n4551), .ZN(n4553)
         );
  OAI211_X1 U5666 ( .C1(n4978), .C2(n6348), .A(n4554), .B(n4553), .ZN(U3095)
         );
  NAND2_X1 U5667 ( .A1(n6393), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4718) );
  NOR2_X1 U5668 ( .A1(n4970), .A2(n4718), .ZN(n4681) );
  INV_X1 U5669 ( .A(n4681), .ZN(n4559) );
  NAND2_X1 U5670 ( .A1(n5117), .A2(n5831), .ZN(n4717) );
  INV_X1 U5671 ( .A(n4717), .ZN(n4680) );
  AND2_X1 U5672 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4681), .ZN(n4584)
         );
  AOI21_X1 U5673 ( .B1(n4555), .B2(n4680), .A(n4584), .ZN(n4561) );
  NAND2_X1 U5674 ( .A1(n4561), .A2(n4556), .ZN(n4557) );
  NOR2_X1 U5675 ( .A1(n5838), .A2(n4557), .ZN(n4558) );
  INV_X1 U5676 ( .A(n5021), .ZN(n4596) );
  AOI211_X2 U5677 ( .C1(n5838), .C2(n4559), .A(n4558), .B(n4596), .ZN(n4589)
         );
  INV_X1 U5678 ( .A(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4565) );
  NAND2_X1 U5679 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4560) );
  OAI22_X1 U5680 ( .A1(n4561), .A2(n5838), .B1(n4560), .B2(n4718), .ZN(n4585)
         );
  AOI22_X1 U5681 ( .A1(n6364), .A2(n4585), .B1(n5039), .B2(n4584), .ZN(n4564)
         );
  NAND2_X1 U5682 ( .A1(n4562), .A2(n5026), .ZN(n4678) );
  INV_X1 U5683 ( .A(n6362), .ZN(n5040) );
  AOI22_X1 U5684 ( .A1(n4712), .A2(n5182), .B1(n4953), .B2(n5040), .ZN(n4563)
         );
  OAI211_X1 U5685 ( .C1(n4589), .C2(n4565), .A(n4564), .B(n4563), .ZN(U3129)
         );
  INV_X1 U5686 ( .A(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4568) );
  AOI22_X1 U5687 ( .A1(n6336), .A2(n4585), .B1(n6292), .B2(n4584), .ZN(n4567)
         );
  INV_X1 U5688 ( .A(n6334), .ZN(n5043) );
  AOI22_X1 U5689 ( .A1(n4712), .A2(n6293), .B1(n4953), .B2(n5043), .ZN(n4566)
         );
  OAI211_X1 U5690 ( .C1(n4589), .C2(n4568), .A(n4567), .B(n4566), .ZN(U3124)
         );
  INV_X1 U5691 ( .A(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4571) );
  AOI22_X1 U5692 ( .A1(n6371), .A2(n4585), .B1(n6279), .B2(n4584), .ZN(n4570)
         );
  INV_X1 U5693 ( .A(n6369), .ZN(n6280) );
  AOI22_X1 U5694 ( .A1(n4712), .A2(n5217), .B1(n4953), .B2(n6280), .ZN(n4569)
         );
  OAI211_X1 U5695 ( .C1(n4589), .C2(n4571), .A(n4570), .B(n4569), .ZN(U3130)
         );
  INV_X1 U5696 ( .A(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4574) );
  AOI22_X1 U5697 ( .A1(n6381), .A2(n4585), .B1(n6284), .B2(n4584), .ZN(n4573)
         );
  INV_X1 U5698 ( .A(n6377), .ZN(n6285) );
  AOI22_X1 U5699 ( .A1(n4712), .A2(n5208), .B1(n4953), .B2(n6285), .ZN(n4572)
         );
  OAI211_X1 U5700 ( .C1(n4589), .C2(n4574), .A(n4573), .B(n4572), .ZN(U3131)
         );
  INV_X1 U5701 ( .A(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4577) );
  AOI22_X1 U5702 ( .A1(n6343), .A2(n4585), .B1(n6300), .B2(n4584), .ZN(n4576)
         );
  INV_X1 U5703 ( .A(n6341), .ZN(n6272) );
  AOI22_X1 U5704 ( .A1(n4712), .A2(n6301), .B1(n4953), .B2(n6272), .ZN(n4575)
         );
  OAI211_X1 U5705 ( .C1(n4589), .C2(n4577), .A(n4576), .B(n4575), .ZN(U3126)
         );
  INV_X1 U5706 ( .A(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4580) );
  AOI22_X1 U5707 ( .A1(n6350), .A2(n4585), .B1(n6305), .B2(n4584), .ZN(n4579)
         );
  INV_X1 U5708 ( .A(n6348), .ZN(n5032) );
  AOI22_X1 U5709 ( .A1(n4712), .A2(n6308), .B1(n4953), .B2(n5032), .ZN(n4578)
         );
  OAI211_X1 U5710 ( .C1(n4589), .C2(n4580), .A(n4579), .B(n4578), .ZN(U3127)
         );
  INV_X1 U5711 ( .A(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4583) );
  AOI22_X1 U5712 ( .A1(n6357), .A2(n4585), .B1(n6275), .B2(n4584), .ZN(n4582)
         );
  INV_X1 U5713 ( .A(n6355), .ZN(n6276) );
  AOI22_X1 U5714 ( .A1(n4712), .A2(n5187), .B1(n4953), .B2(n6276), .ZN(n4581)
         );
  OAI211_X1 U5715 ( .C1(n4589), .C2(n4583), .A(n4582), .B(n4581), .ZN(U3128)
         );
  INV_X1 U5716 ( .A(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4588) );
  AOI22_X1 U5717 ( .A1(n6318), .A2(n4585), .B1(n6296), .B2(n4584), .ZN(n4587)
         );
  INV_X1 U5718 ( .A(n6316), .ZN(n6269) );
  AOI22_X1 U5719 ( .A1(n4712), .A2(n6297), .B1(n4953), .B2(n6269), .ZN(n4586)
         );
  OAI211_X1 U5720 ( .C1(n4589), .C2(n4588), .A(n4587), .B(n4586), .ZN(U3125)
         );
  NAND2_X1 U5721 ( .A1(n4590), .A2(n5834), .ZN(n4591) );
  OAI21_X1 U5722 ( .B1(n4592), .B2(n4591), .A(n5829), .ZN(n4599) );
  AND2_X1 U5723 ( .A1(n5064), .A2(n4593), .ZN(n5178) );
  NOR2_X1 U5724 ( .A1(n4594), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6283)
         );
  AOI21_X1 U5725 ( .B1(n5178), .B2(n5017), .A(n6283), .ZN(n4595) );
  NAND3_X1 U5726 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n4970), .A3(n6399), .ZN(n5168) );
  OAI22_X1 U5727 ( .A1(n4599), .A2(n4595), .B1(n5168), .B2(n6522), .ZN(n6287)
         );
  INV_X1 U5728 ( .A(n6287), .ZN(n4612) );
  INV_X1 U5729 ( .A(n6350), .ZN(n5190) );
  INV_X1 U5730 ( .A(n4595), .ZN(n4598) );
  AOI21_X1 U5731 ( .B1(n5838), .B2(n5168), .A(n4596), .ZN(n4597) );
  OAI21_X1 U5732 ( .B1(n4599), .B2(n4598), .A(n4597), .ZN(n6288) );
  OR3_X1 U5733 ( .A1(n4749), .A2(n5835), .A3(n4600), .ZN(n4602) );
  INV_X1 U5734 ( .A(n4602), .ZN(n4601) );
  NOR2_X2 U5735 ( .A1(n4602), .A2(n5026), .ZN(n6286) );
  AOI22_X1 U5736 ( .A1(n6286), .A2(n5032), .B1(n6305), .B2(n6283), .ZN(n4603)
         );
  OAI21_X1 U5737 ( .B1(n6353), .B2(n6291), .A(n4603), .ZN(n4604) );
  AOI21_X1 U5738 ( .B1(n6288), .B2(INSTQUEUE_REG_3__3__SCAN_IN), .A(n4604), 
        .ZN(n4605) );
  OAI21_X1 U5739 ( .B1(n4612), .B2(n5190), .A(n4605), .ZN(U3047) );
  INV_X1 U5740 ( .A(n6336), .ZN(n5202) );
  AOI22_X1 U5741 ( .A1(n6286), .A2(n5043), .B1(n6292), .B2(n6283), .ZN(n4606)
         );
  OAI21_X1 U5742 ( .B1(n6339), .B2(n6291), .A(n4606), .ZN(n4607) );
  AOI21_X1 U5743 ( .B1(n6288), .B2(INSTQUEUE_REG_3__0__SCAN_IN), .A(n4607), 
        .ZN(n4608) );
  OAI21_X1 U5744 ( .B1(n4612), .B2(n5202), .A(n4608), .ZN(U3044) );
  INV_X1 U5745 ( .A(n6364), .ZN(n5180) );
  AOI22_X1 U5746 ( .A1(n6286), .A2(n5040), .B1(n5039), .B2(n6283), .ZN(n4609)
         );
  OAI21_X1 U5747 ( .B1(n6367), .B2(n6291), .A(n4609), .ZN(n4610) );
  AOI21_X1 U5748 ( .B1(n6288), .B2(INSTQUEUE_REG_3__5__SCAN_IN), .A(n4610), 
        .ZN(n4611) );
  OAI21_X1 U5749 ( .B1(n4612), .B2(n5180), .A(n4611), .ZN(U3049) );
  OAI21_X1 U5750 ( .B1(n4615), .B2(n4614), .A(n4836), .ZN(n4961) );
  OR2_X1 U5751 ( .A1(n4617), .A2(n4616), .ZN(n4618) );
  AND2_X1 U5752 ( .A1(n4618), .A2(n5992), .ZN(n6218) );
  AOI22_X1 U5753 ( .A1(n6060), .A2(n6218), .B1(n5549), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n4619) );
  OAI21_X1 U5754 ( .B1(n4961), .B2(n6056), .A(n4619), .ZN(U2851) );
  AOI22_X1 U5755 ( .A1(n5245), .A2(DATAI_8_), .B1(n6076), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n4620) );
  OAI21_X1 U5756 ( .B1(n4961), .B2(n5877), .A(n4620), .ZN(U2883) );
  OAI22_X1 U5757 ( .A1(n5684), .A2(n4874), .B1(n4889), .B2(n6457), .ZN(n4622)
         );
  NOR2_X1 U5758 ( .A1(n4882), .A2(n6164), .ZN(n4621) );
  AOI211_X1 U5759 ( .C1(n5883), .C2(n4880), .A(n4622), .B(n4621), .ZN(n4623)
         );
  OAI21_X1 U5760 ( .B1(n6166), .B2(n4624), .A(n4623), .ZN(U2981) );
  OAI21_X1 U5761 ( .B1(n4625), .B2(n4923), .A(n4672), .ZN(n4633) );
  INV_X1 U5762 ( .A(n4633), .ZN(n4630) );
  AND2_X1 U5763 ( .A1(n4626), .A2(n5830), .ZN(n4627) );
  AND2_X1 U5764 ( .A1(n5835), .A2(n4627), .ZN(n4632) );
  OAI21_X1 U5765 ( .B1(n4632), .B2(n6164), .A(n5169), .ZN(n4629) );
  OAI21_X1 U5766 ( .B1(n4919), .B2(n5829), .A(n5021), .ZN(n4628) );
  AOI21_X1 U5767 ( .B1(n4630), .B2(n4629), .A(n4628), .ZN(n4677) );
  INV_X1 U5768 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4640) );
  NAND2_X1 U5769 ( .A1(n4632), .A2(n5026), .ZN(n4957) );
  NOR2_X1 U5770 ( .A1(n4957), .A2(n6367), .ZN(n4638) );
  NAND2_X1 U5771 ( .A1(n4633), .A2(n5829), .ZN(n4635) );
  NAND2_X1 U5772 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n4919), .ZN(n4634) );
  NAND2_X1 U5773 ( .A1(n4635), .A2(n4634), .ZN(n4670) );
  NAND2_X1 U5774 ( .A1(n6364), .A2(n4670), .ZN(n4636) );
  OAI21_X1 U5775 ( .B1(n6361), .B2(n4672), .A(n4636), .ZN(n4637) );
  AOI211_X1 U5776 ( .C1(n4789), .C2(n5040), .A(n4638), .B(n4637), .ZN(n4639)
         );
  OAI21_X1 U5777 ( .B1(n4677), .B2(n4640), .A(n4639), .ZN(U3145) );
  INV_X1 U5778 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4645) );
  NOR2_X1 U5779 ( .A1(n4957), .A2(n6346), .ZN(n4643) );
  NAND2_X1 U5780 ( .A1(n6343), .A2(n4670), .ZN(n4641) );
  OAI21_X1 U5781 ( .B1(n6340), .B2(n4672), .A(n4641), .ZN(n4642) );
  AOI211_X1 U5782 ( .C1(n4789), .C2(n6272), .A(n4643), .B(n4642), .ZN(n4644)
         );
  OAI21_X1 U5783 ( .B1(n4677), .B2(n4645), .A(n4644), .ZN(U3142) );
  INV_X1 U5784 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4650) );
  NOR2_X1 U5785 ( .A1(n4957), .A2(n6339), .ZN(n4648) );
  NAND2_X1 U5786 ( .A1(n6336), .A2(n4670), .ZN(n4646) );
  OAI21_X1 U5787 ( .B1(n6333), .B2(n4672), .A(n4646), .ZN(n4647) );
  AOI211_X1 U5788 ( .C1(n4789), .C2(n5043), .A(n4648), .B(n4647), .ZN(n4649)
         );
  OAI21_X1 U5789 ( .B1(n4677), .B2(n4650), .A(n4649), .ZN(U3140) );
  INV_X1 U5790 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4655) );
  NOR2_X1 U5791 ( .A1(n4957), .A2(n6353), .ZN(n4653) );
  NAND2_X1 U5792 ( .A1(n6350), .A2(n4670), .ZN(n4651) );
  OAI21_X1 U5793 ( .B1(n6347), .B2(n4672), .A(n4651), .ZN(n4652) );
  AOI211_X1 U5794 ( .C1(n4789), .C2(n5032), .A(n4653), .B(n4652), .ZN(n4654)
         );
  OAI21_X1 U5795 ( .B1(n4677), .B2(n4655), .A(n4654), .ZN(U3143) );
  INV_X1 U5796 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4660) );
  NOR2_X1 U5797 ( .A1(n4957), .A2(n6386), .ZN(n4658) );
  NAND2_X1 U5798 ( .A1(n6381), .A2(n4670), .ZN(n4656) );
  OAI21_X1 U5799 ( .B1(n6376), .B2(n4672), .A(n4656), .ZN(n4657) );
  AOI211_X1 U5800 ( .C1(n4789), .C2(n6285), .A(n4658), .B(n4657), .ZN(n4659)
         );
  OAI21_X1 U5801 ( .B1(n4677), .B2(n4660), .A(n4659), .ZN(U3147) );
  INV_X1 U5802 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4665) );
  NOR2_X1 U5803 ( .A1(n4957), .A2(n6374), .ZN(n4663) );
  NAND2_X1 U5804 ( .A1(n6371), .A2(n4670), .ZN(n4661) );
  OAI21_X1 U5805 ( .B1(n6368), .B2(n4672), .A(n4661), .ZN(n4662) );
  AOI211_X1 U5806 ( .C1(n4789), .C2(n6280), .A(n4663), .B(n4662), .ZN(n4664)
         );
  OAI21_X1 U5807 ( .B1(n4677), .B2(n4665), .A(n4664), .ZN(U3146) );
  NOR2_X1 U5808 ( .A1(n4957), .A2(n6321), .ZN(n4668) );
  NAND2_X1 U5809 ( .A1(n6318), .A2(n4670), .ZN(n4666) );
  OAI21_X1 U5810 ( .B1(n6315), .B2(n4672), .A(n4666), .ZN(n4667) );
  AOI211_X1 U5811 ( .C1(n4789), .C2(n6269), .A(n4668), .B(n4667), .ZN(n4669)
         );
  OAI21_X1 U5812 ( .B1(n4677), .B2(n6632), .A(n4669), .ZN(U3141) );
  INV_X1 U5813 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4676) );
  NOR2_X1 U5814 ( .A1(n4957), .A2(n6360), .ZN(n4674) );
  NAND2_X1 U5815 ( .A1(n6357), .A2(n4670), .ZN(n4671) );
  OAI21_X1 U5816 ( .B1(n6354), .B2(n4672), .A(n4671), .ZN(n4673) );
  AOI211_X1 U5817 ( .C1(n4789), .C2(n6276), .A(n4674), .B(n4673), .ZN(n4675)
         );
  OAI21_X1 U5818 ( .B1(n4677), .B2(n4676), .A(n4675), .ZN(U3144) );
  AOI21_X1 U5819 ( .B1(n6378), .B2(n4678), .A(n6527), .ZN(n4679) );
  AOI211_X1 U5820 ( .C1(n4680), .C2(n4716), .A(n5838), .B(n4679), .ZN(n4684)
         );
  AND2_X1 U5821 ( .A1(n6691), .A2(n4681), .ZN(n4686) );
  INV_X1 U5822 ( .A(n5058), .ZN(n5175) );
  OAI211_X1 U5823 ( .C1(n6512), .C2(n4686), .A(n5175), .B(n4682), .ZN(n4683)
         );
  NAND2_X1 U5824 ( .A1(n4708), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4689)
         );
  INV_X1 U5825 ( .A(n6357), .ZN(n5185) );
  NOR2_X1 U5826 ( .A1(n4717), .A2(n5838), .ZN(n5065) );
  AOI22_X1 U5827 ( .A1(n5065), .A2(n6038), .B1(n4685), .B2(n5063), .ZN(n4710)
         );
  INV_X1 U5828 ( .A(n4686), .ZN(n4709) );
  OAI22_X1 U5829 ( .A1(n5185), .A2(n4710), .B1(n6354), .B2(n4709), .ZN(n4687)
         );
  AOI21_X1 U5830 ( .B1(n6276), .B2(n4712), .A(n4687), .ZN(n4688) );
  OAI211_X1 U5831 ( .C1(n6378), .C2(n6360), .A(n4689), .B(n4688), .ZN(U3120)
         );
  NAND2_X1 U5832 ( .A1(n4708), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4692)
         );
  INV_X1 U5833 ( .A(n6343), .ZN(n5194) );
  OAI22_X1 U5834 ( .A1(n5194), .A2(n4710), .B1(n6340), .B2(n4709), .ZN(n4690)
         );
  AOI21_X1 U5835 ( .B1(n6272), .B2(n4712), .A(n4690), .ZN(n4691) );
  OAI211_X1 U5836 ( .C1(n6378), .C2(n6346), .A(n4692), .B(n4691), .ZN(U3118)
         );
  NAND2_X1 U5837 ( .A1(n4708), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4695)
         );
  OAI22_X1 U5838 ( .A1(n5202), .A2(n4710), .B1(n6333), .B2(n4709), .ZN(n4693)
         );
  AOI21_X1 U5839 ( .B1(n5043), .B2(n4712), .A(n4693), .ZN(n4694) );
  OAI211_X1 U5840 ( .C1(n6378), .C2(n6339), .A(n4695), .B(n4694), .ZN(U3116)
         );
  NAND2_X1 U5841 ( .A1(n4708), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4698)
         );
  INV_X1 U5842 ( .A(n6381), .ZN(n5206) );
  OAI22_X1 U5843 ( .A1(n5206), .A2(n4710), .B1(n6376), .B2(n4709), .ZN(n4696)
         );
  AOI21_X1 U5844 ( .B1(n6285), .B2(n4712), .A(n4696), .ZN(n4697) );
  OAI211_X1 U5845 ( .C1(n6378), .C2(n6386), .A(n4698), .B(n4697), .ZN(U3123)
         );
  NAND2_X1 U5846 ( .A1(n4708), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4701)
         );
  OAI22_X1 U5847 ( .A1(n5198), .A2(n4710), .B1(n6315), .B2(n4709), .ZN(n4699)
         );
  AOI21_X1 U5848 ( .B1(n6269), .B2(n4712), .A(n4699), .ZN(n4700) );
  OAI211_X1 U5849 ( .C1(n6378), .C2(n6321), .A(n4701), .B(n4700), .ZN(U3117)
         );
  NAND2_X1 U5850 ( .A1(n4708), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4704)
         );
  INV_X1 U5851 ( .A(n6371), .ZN(n5214) );
  OAI22_X1 U5852 ( .A1(n5214), .A2(n4710), .B1(n6368), .B2(n4709), .ZN(n4702)
         );
  AOI21_X1 U5853 ( .B1(n6280), .B2(n4712), .A(n4702), .ZN(n4703) );
  OAI211_X1 U5854 ( .C1(n6378), .C2(n6374), .A(n4704), .B(n4703), .ZN(U3122)
         );
  NAND2_X1 U5855 ( .A1(n4708), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4707)
         );
  OAI22_X1 U5856 ( .A1(n5190), .A2(n4710), .B1(n6347), .B2(n4709), .ZN(n4705)
         );
  AOI21_X1 U5857 ( .B1(n5032), .B2(n4712), .A(n4705), .ZN(n4706) );
  OAI211_X1 U5858 ( .C1(n6378), .C2(n6353), .A(n4707), .B(n4706), .ZN(U3119)
         );
  NAND2_X1 U5859 ( .A1(n4708), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4714)
         );
  OAI22_X1 U5860 ( .A1(n5180), .A2(n4710), .B1(n6361), .B2(n4709), .ZN(n4711)
         );
  AOI21_X1 U5861 ( .B1(n5040), .B2(n4712), .A(n4711), .ZN(n4713) );
  OAI211_X1 U5862 ( .C1(n6378), .C2(n6367), .A(n4714), .B(n4713), .ZN(U3121)
         );
  AOI21_X1 U5863 ( .B1(n4723), .B2(n4715), .A(n5838), .ZN(n4726) );
  OR2_X1 U5864 ( .A1(n4717), .A2(n4716), .ZN(n5054) );
  OR2_X1 U5865 ( .A1(n4718), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5052)
         );
  NOR2_X1 U5866 ( .A1(n6691), .A2(n5052), .ZN(n4794) );
  INV_X1 U5867 ( .A(n4794), .ZN(n4719) );
  OAI21_X1 U5868 ( .B1(n5054), .B2(n4903), .A(n4719), .ZN(n4724) );
  INV_X1 U5869 ( .A(n5052), .ZN(n4720) );
  AOI22_X1 U5870 ( .A1(n4726), .A2(n4724), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4720), .ZN(n4798) );
  INV_X1 U5871 ( .A(n4724), .ZN(n4725) );
  AOI22_X1 U5872 ( .A1(n4726), .A2(n4725), .B1(n5052), .B2(n5838), .ZN(n4727)
         );
  NAND2_X1 U5873 ( .A1(n5021), .A2(n4727), .ZN(n4793) );
  AOI22_X1 U5874 ( .A1(n6279), .A2(n4794), .B1(INSTQUEUE_REG_5__6__SCAN_IN), 
        .B2(n4793), .ZN(n4728) );
  OAI21_X1 U5875 ( .B1(n6374), .B2(n5094), .A(n4728), .ZN(n4729) );
  AOI21_X1 U5876 ( .B1(n6280), .B2(n6307), .A(n4729), .ZN(n4730) );
  OAI21_X1 U5877 ( .B1(n4798), .B2(n5214), .A(n4730), .ZN(U3066) );
  AOI22_X1 U5878 ( .A1(n6284), .A2(n4794), .B1(INSTQUEUE_REG_5__7__SCAN_IN), 
        .B2(n4793), .ZN(n4731) );
  OAI21_X1 U5879 ( .B1(n6386), .B2(n5094), .A(n4731), .ZN(n4732) );
  AOI21_X1 U5880 ( .B1(n6285), .B2(n6307), .A(n4732), .ZN(n4733) );
  OAI21_X1 U5881 ( .B1(n4798), .B2(n5206), .A(n4733), .ZN(U3067) );
  AOI22_X1 U5882 ( .A1(n6292), .A2(n4794), .B1(INSTQUEUE_REG_5__0__SCAN_IN), 
        .B2(n4793), .ZN(n4734) );
  OAI21_X1 U5883 ( .B1(n6339), .B2(n5094), .A(n4734), .ZN(n4735) );
  AOI21_X1 U5884 ( .B1(n5043), .B2(n6307), .A(n4735), .ZN(n4736) );
  OAI21_X1 U5885 ( .B1(n4798), .B2(n5202), .A(n4736), .ZN(U3060) );
  AOI22_X1 U5886 ( .A1(n6305), .A2(n4794), .B1(INSTQUEUE_REG_5__3__SCAN_IN), 
        .B2(n4793), .ZN(n4737) );
  OAI21_X1 U5887 ( .B1(n6353), .B2(n5094), .A(n4737), .ZN(n4738) );
  AOI21_X1 U5888 ( .B1(n5032), .B2(n6307), .A(n4738), .ZN(n4739) );
  OAI21_X1 U5889 ( .B1(n4798), .B2(n5190), .A(n4739), .ZN(U3063) );
  AOI22_X1 U5890 ( .A1(n5039), .A2(n4794), .B1(INSTQUEUE_REG_5__5__SCAN_IN), 
        .B2(n4793), .ZN(n4740) );
  OAI21_X1 U5891 ( .B1(n6367), .B2(n5094), .A(n4740), .ZN(n4741) );
  AOI21_X1 U5892 ( .B1(n5040), .B2(n6307), .A(n4741), .ZN(n4742) );
  OAI21_X1 U5893 ( .B1(n4798), .B2(n5180), .A(n4742), .ZN(U3065) );
  AOI22_X1 U5894 ( .A1(n6275), .A2(n4794), .B1(INSTQUEUE_REG_5__4__SCAN_IN), 
        .B2(n4793), .ZN(n4743) );
  OAI21_X1 U5895 ( .B1(n6360), .B2(n5094), .A(n4743), .ZN(n4744) );
  AOI21_X1 U5896 ( .B1(n6276), .B2(n6307), .A(n4744), .ZN(n4745) );
  OAI21_X1 U5897 ( .B1(n4798), .B2(n5185), .A(n4745), .ZN(U3064) );
  AOI22_X1 U5898 ( .A1(n6300), .A2(n4794), .B1(INSTQUEUE_REG_5__2__SCAN_IN), 
        .B2(n4793), .ZN(n4746) );
  OAI21_X1 U5899 ( .B1(n6346), .B2(n5094), .A(n4746), .ZN(n4747) );
  AOI21_X1 U5900 ( .B1(n6272), .B2(n6307), .A(n4747), .ZN(n4748) );
  OAI21_X1 U5901 ( .B1(n4798), .B2(n5194), .A(n4748), .ZN(U3062) );
  OR3_X1 U5902 ( .A1(n4749), .A2(n5835), .A3(n5830), .ZN(n5027) );
  INV_X1 U5903 ( .A(n5027), .ZN(n5019) );
  NAND2_X1 U5904 ( .A1(n5019), .A2(n5026), .ZN(n5051) );
  INV_X1 U5905 ( .A(n4789), .ZN(n4750) );
  NAND3_X1 U5906 ( .A1(n5051), .A2(n5829), .A3(n4750), .ZN(n4751) );
  NAND2_X1 U5907 ( .A1(n4751), .A2(n5169), .ZN(n4756) );
  NAND2_X1 U5908 ( .A1(n5064), .A2(n4752), .ZN(n5016) );
  NAND3_X1 U5909 ( .A1(n4970), .A2(n6399), .A3(n6393), .ZN(n5023) );
  NOR2_X1 U5910 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5023), .ZN(n4785)
         );
  OR2_X1 U5911 ( .A1(n4753), .A2(n5177), .ZN(n5061) );
  AOI21_X1 U5912 ( .B1(n5061), .B2(STATE2_REG_2__SCAN_IN), .A(n4754), .ZN(
        n5056) );
  OAI211_X1 U5913 ( .C1(n6512), .C2(n4785), .A(n4916), .B(n5056), .ZN(n4755)
         );
  AOI21_X1 U5914 ( .B1(n4756), .B2(n5016), .A(n4755), .ZN(n4792) );
  INV_X1 U5915 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4760) );
  OAI22_X1 U5916 ( .A1(n5016), .A2(n5838), .B1(n5175), .B2(n5061), .ZN(n4786)
         );
  AOI22_X1 U5917 ( .A1(n6336), .A2(n4786), .B1(n6292), .B2(n4785), .ZN(n4757)
         );
  OAI21_X1 U5918 ( .B1(n6334), .B2(n5051), .A(n4757), .ZN(n4758) );
  AOI21_X1 U5919 ( .B1(n6293), .B2(n4789), .A(n4758), .ZN(n4759) );
  OAI21_X1 U5920 ( .B1(n4792), .B2(n4760), .A(n4759), .ZN(U3020) );
  INV_X1 U5921 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4764) );
  AOI22_X1 U5922 ( .A1(n6318), .A2(n4786), .B1(n6296), .B2(n4785), .ZN(n4761)
         );
  OAI21_X1 U5923 ( .B1(n6316), .B2(n5051), .A(n4761), .ZN(n4762) );
  AOI21_X1 U5924 ( .B1(n6297), .B2(n4789), .A(n4762), .ZN(n4763) );
  OAI21_X1 U5925 ( .B1(n4792), .B2(n4764), .A(n4763), .ZN(U3021) );
  INV_X1 U5926 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4768) );
  AOI22_X1 U5927 ( .A1(n6350), .A2(n4786), .B1(n6305), .B2(n4785), .ZN(n4765)
         );
  OAI21_X1 U5928 ( .B1(n6348), .B2(n5051), .A(n4765), .ZN(n4766) );
  AOI21_X1 U5929 ( .B1(n6308), .B2(n4789), .A(n4766), .ZN(n4767) );
  OAI21_X1 U5930 ( .B1(n4792), .B2(n4768), .A(n4767), .ZN(U3023) );
  INV_X1 U5931 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4772) );
  AOI22_X1 U5932 ( .A1(n6357), .A2(n4786), .B1(n6275), .B2(n4785), .ZN(n4769)
         );
  OAI21_X1 U5933 ( .B1(n6355), .B2(n5051), .A(n4769), .ZN(n4770) );
  AOI21_X1 U5934 ( .B1(n5187), .B2(n4789), .A(n4770), .ZN(n4771) );
  OAI21_X1 U5935 ( .B1(n4792), .B2(n4772), .A(n4771), .ZN(U3024) );
  INV_X1 U5936 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4776) );
  AOI22_X1 U5937 ( .A1(n6343), .A2(n4786), .B1(n6300), .B2(n4785), .ZN(n4773)
         );
  OAI21_X1 U5938 ( .B1(n6341), .B2(n5051), .A(n4773), .ZN(n4774) );
  AOI21_X1 U5939 ( .B1(n6301), .B2(n4789), .A(n4774), .ZN(n4775) );
  OAI21_X1 U5940 ( .B1(n4792), .B2(n4776), .A(n4775), .ZN(U3022) );
  INV_X1 U5941 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4780) );
  AOI22_X1 U5942 ( .A1(n6371), .A2(n4786), .B1(n6279), .B2(n4785), .ZN(n4777)
         );
  OAI21_X1 U5943 ( .B1(n6369), .B2(n5051), .A(n4777), .ZN(n4778) );
  AOI21_X1 U5944 ( .B1(n5217), .B2(n4789), .A(n4778), .ZN(n4779) );
  OAI21_X1 U5945 ( .B1(n4792), .B2(n4780), .A(n4779), .ZN(U3026) );
  INV_X1 U5946 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4784) );
  AOI22_X1 U5947 ( .A1(n6381), .A2(n4786), .B1(n6284), .B2(n4785), .ZN(n4781)
         );
  OAI21_X1 U5948 ( .B1(n6377), .B2(n5051), .A(n4781), .ZN(n4782) );
  AOI21_X1 U5949 ( .B1(n5208), .B2(n4789), .A(n4782), .ZN(n4783) );
  OAI21_X1 U5950 ( .B1(n4792), .B2(n4784), .A(n4783), .ZN(U3027) );
  INV_X1 U5951 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4791) );
  AOI22_X1 U5952 ( .A1(n6364), .A2(n4786), .B1(n5039), .B2(n4785), .ZN(n4787)
         );
  OAI21_X1 U5953 ( .B1(n6362), .B2(n5051), .A(n4787), .ZN(n4788) );
  AOI21_X1 U5954 ( .B1(n5182), .B2(n4789), .A(n4788), .ZN(n4790) );
  OAI21_X1 U5955 ( .B1(n4792), .B2(n4791), .A(n4790), .ZN(U3025) );
  AOI22_X1 U5956 ( .A1(n6296), .A2(n4794), .B1(INSTQUEUE_REG_5__1__SCAN_IN), 
        .B2(n4793), .ZN(n4795) );
  OAI21_X1 U5957 ( .B1(n6321), .B2(n5094), .A(n4795), .ZN(n4796) );
  AOI21_X1 U5958 ( .B1(n6269), .B2(n6307), .A(n4796), .ZN(n4797) );
  OAI21_X1 U5959 ( .B1(n4798), .B2(n5198), .A(n4797), .ZN(U3061) );
  OAI21_X1 U5960 ( .B1(n4801), .B2(n4800), .A(n4799), .ZN(n6226) );
  NAND2_X1 U5961 ( .A1(n6018), .A2(REIP_REG_7__SCAN_IN), .ZN(n6223) );
  NAND2_X1 U5962 ( .A1(n6171), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4802)
         );
  OAI211_X1 U5963 ( .C1(n6182), .C2(n4843), .A(n6223), .B(n4802), .ZN(n4803)
         );
  AOI21_X1 U5964 ( .B1(n4804), .B2(n6176), .A(n4803), .ZN(n4805) );
  OAI21_X1 U5965 ( .B1(n6226), .B2(n6166), .A(n4805), .ZN(U2979) );
  NAND2_X1 U5966 ( .A1(n4806), .A2(n5829), .ZN(n4813) );
  INV_X1 U5967 ( .A(n4807), .ZN(n4808) );
  INV_X1 U5968 ( .A(n6325), .ZN(n4825) );
  AOI21_X1 U5969 ( .B1(n4808), .B2(n5017), .A(n4825), .ZN(n4810) );
  OAI22_X1 U5970 ( .A1(n4813), .A2(n4810), .B1(n4809), .B2(n6522), .ZN(n6328)
         );
  INV_X1 U5971 ( .A(n6328), .ZN(n4830) );
  INV_X1 U5972 ( .A(n6326), .ZN(n4828) );
  INV_X1 U5973 ( .A(n4810), .ZN(n4812) );
  OAI22_X1 U5974 ( .A1(n4813), .A2(n4812), .B1(n5829), .B2(n4811), .ZN(n4814)
         );
  INV_X1 U5975 ( .A(n4814), .ZN(n4815) );
  NAND2_X1 U5976 ( .A1(n5021), .A2(n4815), .ZN(n6329) );
  AOI22_X1 U5977 ( .A1(n6284), .A2(n4825), .B1(INSTQUEUE_REG_7__7__SCAN_IN), 
        .B2(n6329), .ZN(n4816) );
  OAI21_X1 U5978 ( .B1(n6386), .B2(n6332), .A(n4816), .ZN(n4817) );
  AOI21_X1 U5979 ( .B1(n6285), .B2(n4828), .A(n4817), .ZN(n4818) );
  OAI21_X1 U5980 ( .B1(n4830), .B2(n5206), .A(n4818), .ZN(U3083) );
  AOI22_X1 U5981 ( .A1(n5039), .A2(n4825), .B1(INSTQUEUE_REG_7__5__SCAN_IN), 
        .B2(n6329), .ZN(n4819) );
  OAI21_X1 U5982 ( .B1(n6367), .B2(n6332), .A(n4819), .ZN(n4820) );
  AOI21_X1 U5983 ( .B1(n5040), .B2(n4828), .A(n4820), .ZN(n4821) );
  OAI21_X1 U5984 ( .B1(n4830), .B2(n5180), .A(n4821), .ZN(U3081) );
  AOI22_X1 U5985 ( .A1(n6305), .A2(n4825), .B1(INSTQUEUE_REG_7__3__SCAN_IN), 
        .B2(n6329), .ZN(n4822) );
  OAI21_X1 U5986 ( .B1(n6353), .B2(n6332), .A(n4822), .ZN(n4823) );
  AOI21_X1 U5987 ( .B1(n5032), .B2(n4828), .A(n4823), .ZN(n4824) );
  OAI21_X1 U5988 ( .B1(n4830), .B2(n5190), .A(n4824), .ZN(U3079) );
  AOI22_X1 U5989 ( .A1(n6300), .A2(n4825), .B1(INSTQUEUE_REG_7__2__SCAN_IN), 
        .B2(n6329), .ZN(n4826) );
  OAI21_X1 U5990 ( .B1(n6346), .B2(n6332), .A(n4826), .ZN(n4827) );
  AOI21_X1 U5991 ( .B1(n6272), .B2(n4828), .A(n4827), .ZN(n4829) );
  OAI21_X1 U5992 ( .B1(n4830), .B2(n5194), .A(n4829), .ZN(U3078) );
  AOI22_X1 U5993 ( .A1(n6171), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6018), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n4832) );
  INV_X1 U5994 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4897) );
  NAND2_X1 U5995 ( .A1(n5883), .A2(n4897), .ZN(n4831) );
  OAI211_X1 U5996 ( .C1(n4902), .C2(n6164), .A(n4832), .B(n4831), .ZN(n4833)
         );
  AOI21_X1 U5997 ( .B1(n6178), .B2(n4834), .A(n4833), .ZN(n4835) );
  INV_X1 U5998 ( .A(n4835), .ZN(U2985) );
  INV_X1 U5999 ( .A(n4836), .ZN(n4840) );
  INV_X1 U6000 ( .A(n4837), .ZN(n4839) );
  INV_X1 U6001 ( .A(n4838), .ZN(n4912) );
  OAI21_X1 U6002 ( .B1(n4840), .B2(n4839), .A(n4912), .ZN(n5997) );
  AOI22_X1 U6003 ( .A1(n5245), .A2(DATAI_9_), .B1(n6076), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n4841) );
  OAI21_X1 U6004 ( .B1(n5997), .B2(n5877), .A(n4841), .ZN(U2882) );
  AND2_X1 U6005 ( .A1(n5596), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4842) );
  INV_X1 U6006 ( .A(n4843), .ZN(n4857) );
  NAND2_X1 U6007 ( .A1(n4844), .A2(n5123), .ZN(n4863) );
  NAND2_X1 U6008 ( .A1(n4863), .A2(n6015), .ZN(n6012) );
  INV_X1 U6009 ( .A(n4845), .ZN(n4848) );
  INV_X1 U6010 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5430) );
  NAND2_X1 U6011 ( .A1(n4846), .A2(n5430), .ZN(n4847) );
  NAND2_X1 U6012 ( .A1(n4848), .A2(n4847), .ZN(n4849) );
  INV_X1 U6013 ( .A(n6032), .ZN(n6005) );
  NAND2_X1 U6014 ( .A1(n6225), .A2(n6033), .ZN(n4850) );
  OAI211_X1 U6015 ( .C1(n4851), .C2(n6005), .A(n4850), .B(n4889), .ZN(n4852)
         );
  AOI21_X1 U6016 ( .B1(n6008), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n4852), 
        .ZN(n4855) );
  NOR3_X1 U6017 ( .A1(n6021), .A2(n6457), .A3(n4875), .ZN(n6009) );
  INV_X1 U6018 ( .A(n4862), .ZN(n4853) );
  OAI211_X1 U6019 ( .C1(REIP_REG_7__SCAN_IN), .C2(REIP_REG_6__SCAN_IN), .A(
        n6009), .B(n4853), .ZN(n4854) );
  OAI211_X1 U6020 ( .C1(n6012), .C2(n6460), .A(n4855), .B(n4854), .ZN(n4856)
         );
  AOI21_X1 U6021 ( .B1(n6044), .B2(n4857), .A(n4856), .ZN(n4858) );
  OAI21_X1 U6022 ( .B1(n4859), .B2(n5985), .A(n4858), .ZN(U2820) );
  INV_X1 U6023 ( .A(n4963), .ZN(n4867) );
  AOI21_X1 U6024 ( .B1(n6032), .B2(EBX_REG_8__SCAN_IN), .A(n6018), .ZN(n4861)
         );
  NAND2_X1 U6025 ( .A1(n6218), .A2(n6033), .ZN(n4860) );
  OAI211_X1 U6026 ( .C1(n6036), .C2(n6569), .A(n4861), .B(n4860), .ZN(n4866)
         );
  INV_X1 U6027 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6462) );
  NAND2_X1 U6028 ( .A1(n4862), .A2(n6009), .ZN(n5007) );
  OAI21_X1 U6029 ( .B1(n4864), .B2(n4863), .A(n6015), .ZN(n5959) );
  AOI21_X1 U6030 ( .B1(n6462), .B2(n5007), .A(n5959), .ZN(n4865) );
  AOI211_X1 U6031 ( .C1(n6044), .C2(n4867), .A(n4866), .B(n4865), .ZN(n4868)
         );
  OAI21_X1 U6032 ( .B1(n5985), .B2(n4961), .A(n4868), .ZN(U2819) );
  OR2_X1 U6033 ( .A1(n4869), .A2(n4893), .ZN(n4870) );
  INV_X1 U6034 ( .A(n4871), .ZN(n4872) );
  AOI22_X1 U6035 ( .A1(n6033), .A2(n4872), .B1(n6032), .B2(EBX_REG_5__SCAN_IN), 
        .ZN(n4873) );
  OAI211_X1 U6036 ( .C1(n6036), .C2(n4874), .A(n4873), .B(n4889), .ZN(n4879)
         );
  INV_X1 U6037 ( .A(n4875), .ZN(n4876) );
  NAND2_X1 U6038 ( .A1(n5118), .A2(n4876), .ZN(n4877) );
  AOI21_X1 U6039 ( .B1(n6457), .B2(n4877), .A(n6012), .ZN(n4878) );
  AOI211_X1 U6040 ( .C1(n6044), .C2(n4880), .A(n4879), .B(n4878), .ZN(n4881)
         );
  OAI21_X1 U6041 ( .B1(n6041), .B2(n4882), .A(n4881), .ZN(U2822) );
  NAND2_X1 U6043 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6234), .ZN(n5156)
         );
  INV_X1 U6044 ( .A(n6199), .ZN(n6260) );
  OAI21_X1 U6045 ( .B1(n6260), .B2(n4883), .A(n6255), .ZN(n6253) );
  OAI33_X1 U6046 ( .A1(1'b0), .A2(n4884), .A3(n6655), .B1(
        INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n5156), .B3(n6253), .ZN(n4892) );
  OAI21_X1 U6047 ( .B1(n4888), .B2(n4887), .A(n4886), .ZN(n6155) );
  NOR2_X1 U6048 ( .A1(n6155), .A2(n6242), .ZN(n4891) );
  OAI22_X1 U6049 ( .A1(n6246), .A2(n6004), .B1(n4889), .B2(n6459), .ZN(n4890)
         );
  OR3_X1 U6050 ( .A1(n4892), .A2(n4891), .A3(n4890), .ZN(U3012) );
  INV_X1 U6051 ( .A(n5123), .ZN(n6016) );
  AOI22_X1 U6052 ( .A1(EBX_REG_1__SCAN_IN), .A2(n6032), .B1(n6016), .B2(
        REIP_REG_1__SCAN_IN), .ZN(n4901) );
  NOR2_X1 U6053 ( .A1(n4894), .A2(n4893), .ZN(n6039) );
  INV_X1 U6054 ( .A(n6039), .ZN(n5121) );
  AOI22_X1 U6055 ( .A1(n4895), .A2(n6033), .B1(n5118), .B2(n6513), .ZN(n4896)
         );
  OAI21_X1 U6056 ( .B1(n5831), .B2(n5121), .A(n4896), .ZN(n4899) );
  NOR2_X1 U6057 ( .A1(n6036), .A2(n4897), .ZN(n4898) );
  AOI211_X1 U6058 ( .C1(n6044), .C2(n4897), .A(n4899), .B(n4898), .ZN(n4900)
         );
  OAI211_X1 U6059 ( .C1(n6041), .C2(n4902), .A(n4901), .B(n4900), .ZN(U2826)
         );
  NOR2_X1 U6060 ( .A1(n4903), .A2(n5121), .ZN(n4907) );
  OAI22_X1 U6061 ( .A1(n4905), .A2(n6024), .B1(n6005), .B2(n4904), .ZN(n4906)
         );
  AOI211_X1 U6062 ( .C1(n6015), .C2(REIP_REG_0__SCAN_IN), .A(n4907), .B(n4906), 
        .ZN(n4909) );
  OAI21_X1 U6063 ( .B1(n6008), .B2(n6044), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4908) );
  OAI211_X1 U6064 ( .C1(n4910), .C2(n6041), .A(n4909), .B(n4908), .ZN(U2827)
         );
  OR2_X1 U6065 ( .A1(n4912), .A2(n4911), .ZN(n5096) );
  NAND2_X1 U6066 ( .A1(n4912), .A2(n4911), .ZN(n4913) );
  NAND2_X1 U6067 ( .A1(n5096), .A2(n4913), .ZN(n5136) );
  AOI22_X1 U6068 ( .A1(n5245), .A2(DATAI_10_), .B1(n6076), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n4914) );
  OAI21_X1 U6069 ( .B1(n5136), .B2(n5877), .A(n4914), .ZN(U2881) );
  INV_X1 U6070 ( .A(n4915), .ZN(n4918) );
  NOR2_X1 U6071 ( .A1(n4916), .A2(n4970), .ZN(n4917) );
  AOI22_X1 U6072 ( .A1(n4918), .A2(n6038), .B1(n5177), .B2(n4917), .ZN(n4951)
         );
  INV_X1 U6073 ( .A(n4919), .ZN(n4920) );
  NOR2_X1 U6074 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4920), .ZN(n4924)
         );
  INV_X1 U6075 ( .A(n4924), .ZN(n4950) );
  OAI22_X1 U6076 ( .A1(n5190), .A2(n4951), .B1(n6347), .B2(n4950), .ZN(n4921)
         );
  AOI21_X1 U6077 ( .B1(n6308), .B2(n4953), .A(n4921), .ZN(n4931) );
  INV_X1 U6078 ( .A(n4953), .ZN(n4922) );
  AOI21_X1 U6079 ( .B1(n4922), .B2(n4957), .A(n6527), .ZN(n4929) );
  NAND2_X1 U6080 ( .A1(n5829), .A2(n4923), .ZN(n4928) );
  OAI21_X1 U6081 ( .B1(n6512), .B2(n4924), .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .ZN(n4925) );
  INV_X1 U6082 ( .A(n4925), .ZN(n4926) );
  OAI211_X1 U6083 ( .C1(n4929), .C2(n4928), .A(n4927), .B(n4926), .ZN(n4954)
         );
  NAND2_X1 U6084 ( .A1(n4954), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4930)
         );
  OAI211_X1 U6085 ( .C1(n4957), .C2(n6348), .A(n4931), .B(n4930), .ZN(U3135)
         );
  OAI22_X1 U6086 ( .A1(n5194), .A2(n4951), .B1(n6340), .B2(n4950), .ZN(n4932)
         );
  AOI21_X1 U6087 ( .B1(n6301), .B2(n4953), .A(n4932), .ZN(n4934) );
  NAND2_X1 U6088 ( .A1(n4954), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4933)
         );
  OAI211_X1 U6089 ( .C1(n4957), .C2(n6341), .A(n4934), .B(n4933), .ZN(U3134)
         );
  OAI22_X1 U6090 ( .A1(n5180), .A2(n4951), .B1(n6361), .B2(n4950), .ZN(n4935)
         );
  AOI21_X1 U6091 ( .B1(n5182), .B2(n4953), .A(n4935), .ZN(n4937) );
  NAND2_X1 U6092 ( .A1(n4954), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4936)
         );
  OAI211_X1 U6093 ( .C1(n4957), .C2(n6362), .A(n4937), .B(n4936), .ZN(U3137)
         );
  OAI22_X1 U6094 ( .A1(n5185), .A2(n4951), .B1(n6354), .B2(n4950), .ZN(n4938)
         );
  AOI21_X1 U6095 ( .B1(n5187), .B2(n4953), .A(n4938), .ZN(n4940) );
  NAND2_X1 U6096 ( .A1(n4954), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4939)
         );
  OAI211_X1 U6097 ( .C1(n4957), .C2(n6355), .A(n4940), .B(n4939), .ZN(U3136)
         );
  OAI22_X1 U6098 ( .A1(n5206), .A2(n4951), .B1(n6376), .B2(n4950), .ZN(n4941)
         );
  AOI21_X1 U6099 ( .B1(n5208), .B2(n4953), .A(n4941), .ZN(n4943) );
  NAND2_X1 U6100 ( .A1(n4954), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4942)
         );
  OAI211_X1 U6101 ( .C1(n4957), .C2(n6377), .A(n4943), .B(n4942), .ZN(U3139)
         );
  OAI22_X1 U6102 ( .A1(n5214), .A2(n4951), .B1(n6368), .B2(n4950), .ZN(n4944)
         );
  AOI21_X1 U6103 ( .B1(n5217), .B2(n4953), .A(n4944), .ZN(n4946) );
  NAND2_X1 U6104 ( .A1(n4954), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4945)
         );
  OAI211_X1 U6105 ( .C1(n4957), .C2(n6369), .A(n4946), .B(n4945), .ZN(U3138)
         );
  OAI22_X1 U6106 ( .A1(n5202), .A2(n4951), .B1(n6333), .B2(n4950), .ZN(n4947)
         );
  AOI21_X1 U6107 ( .B1(n6293), .B2(n4953), .A(n4947), .ZN(n4949) );
  NAND2_X1 U6108 ( .A1(n4954), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4948)
         );
  OAI211_X1 U6109 ( .C1(n4957), .C2(n6334), .A(n4949), .B(n4948), .ZN(U3132)
         );
  OAI22_X1 U6110 ( .A1(n5198), .A2(n4951), .B1(n6315), .B2(n4950), .ZN(n4952)
         );
  AOI21_X1 U6111 ( .B1(n6297), .B2(n4953), .A(n4952), .ZN(n4956) );
  NAND2_X1 U6112 ( .A1(n4954), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4955)
         );
  OAI211_X1 U6113 ( .C1(n4957), .C2(n6316), .A(n4956), .B(n4955), .ZN(U3133)
         );
  OAI21_X1 U6114 ( .B1(n4960), .B2(n4959), .A(n5101), .ZN(n6216) );
  INV_X1 U6115 ( .A(n4961), .ZN(n4965) );
  AOI22_X1 U6116 ( .A1(n6171), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n6018), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n4962) );
  OAI21_X1 U6117 ( .B1(n6182), .B2(n4963), .A(n4962), .ZN(n4964) );
  AOI21_X1 U6118 ( .B1(n4965), .B2(n6176), .A(n4964), .ZN(n4966) );
  OAI21_X1 U6119 ( .B1(n6216), .B2(n6166), .A(n4966), .ZN(U2978) );
  INV_X1 U6120 ( .A(EBX_REG_10__SCAN_IN), .ZN(n4968) );
  XNOR2_X1 U6121 ( .A(n4967), .B(n5991), .ZN(n6196) );
  OAI222_X1 U6122 ( .A1(n6056), .A2(n5136), .B1(n4968), .B2(n6065), .C1(n6055), 
        .C2(n6196), .ZN(U2849) );
  AOI21_X1 U6123 ( .B1(n4978), .B2(n6385), .A(n6527), .ZN(n4969) );
  NOR2_X1 U6124 ( .A1(n4969), .A2(n5838), .ZN(n4976) );
  NOR2_X1 U6125 ( .A1(n5175), .A2(n4970), .ZN(n4971) );
  AOI22_X1 U6126 ( .A1(n4976), .A2(n4972), .B1(n5177), .B2(n4971), .ZN(n5006)
         );
  NOR2_X1 U6127 ( .A1(n5063), .A2(n4973), .ZN(n5173) );
  OR2_X1 U6128 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4974), .ZN(n5001)
         );
  AOI22_X1 U6129 ( .A1(n4976), .A2(n4975), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n5001), .ZN(n4977) );
  OAI211_X1 U6130 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6522), .A(n5173), .B(n4977), .ZN(n5000) );
  NAND2_X1 U6131 ( .A1(n5000), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4981)
         );
  INV_X1 U6132 ( .A(n4978), .ZN(n5003) );
  OAI22_X1 U6133 ( .A1(n6385), .A2(n6348), .B1(n5001), .B2(n6347), .ZN(n4979)
         );
  AOI21_X1 U6134 ( .B1(n5003), .B2(n6308), .A(n4979), .ZN(n4980) );
  OAI211_X1 U6135 ( .C1(n5006), .C2(n5190), .A(n4981), .B(n4980), .ZN(U3103)
         );
  NAND2_X1 U6136 ( .A1(n5000), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4984)
         );
  OAI22_X1 U6137 ( .A1(n6385), .A2(n6334), .B1(n5001), .B2(n6333), .ZN(n4982)
         );
  AOI21_X1 U6138 ( .B1(n5003), .B2(n6293), .A(n4982), .ZN(n4983) );
  OAI211_X1 U6139 ( .C1(n5006), .C2(n5202), .A(n4984), .B(n4983), .ZN(U3100)
         );
  NAND2_X1 U6140 ( .A1(n5000), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4987)
         );
  OAI22_X1 U6141 ( .A1(n6385), .A2(n6362), .B1(n5001), .B2(n6361), .ZN(n4985)
         );
  AOI21_X1 U6142 ( .B1(n5003), .B2(n5182), .A(n4985), .ZN(n4986) );
  OAI211_X1 U6143 ( .C1(n5006), .C2(n5180), .A(n4987), .B(n4986), .ZN(U3105)
         );
  NAND2_X1 U6144 ( .A1(n5000), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4990)
         );
  OAI22_X1 U6145 ( .A1(n6385), .A2(n6377), .B1(n5001), .B2(n6376), .ZN(n4988)
         );
  AOI21_X1 U6146 ( .B1(n5003), .B2(n5208), .A(n4988), .ZN(n4989) );
  OAI211_X1 U6147 ( .C1(n5006), .C2(n5206), .A(n4990), .B(n4989), .ZN(U3107)
         );
  NAND2_X1 U6148 ( .A1(n5000), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4993)
         );
  OAI22_X1 U6149 ( .A1(n6385), .A2(n6341), .B1(n5001), .B2(n6340), .ZN(n4991)
         );
  AOI21_X1 U6150 ( .B1(n5003), .B2(n6301), .A(n4991), .ZN(n4992) );
  OAI211_X1 U6151 ( .C1(n5006), .C2(n5194), .A(n4993), .B(n4992), .ZN(U3102)
         );
  NAND2_X1 U6152 ( .A1(n5000), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4996)
         );
  OAI22_X1 U6153 ( .A1(n6385), .A2(n6355), .B1(n5001), .B2(n6354), .ZN(n4994)
         );
  AOI21_X1 U6154 ( .B1(n5003), .B2(n5187), .A(n4994), .ZN(n4995) );
  OAI211_X1 U6155 ( .C1(n5006), .C2(n5185), .A(n4996), .B(n4995), .ZN(U3104)
         );
  NAND2_X1 U6156 ( .A1(n5000), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4999)
         );
  OAI22_X1 U6157 ( .A1(n6385), .A2(n6316), .B1(n5001), .B2(n6315), .ZN(n4997)
         );
  AOI21_X1 U6158 ( .B1(n5003), .B2(n6297), .A(n4997), .ZN(n4998) );
  OAI211_X1 U6159 ( .C1(n5006), .C2(n5198), .A(n4999), .B(n4998), .ZN(U3101)
         );
  NAND2_X1 U6160 ( .A1(n5000), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5005)
         );
  OAI22_X1 U6161 ( .A1(n6385), .A2(n6369), .B1(n5001), .B2(n6368), .ZN(n5002)
         );
  AOI21_X1 U6162 ( .B1(n5003), .B2(n5217), .A(n5002), .ZN(n5004) );
  OAI211_X1 U6163 ( .C1(n5006), .C2(n5214), .A(n5005), .B(n5004), .ZN(U3106)
         );
  INV_X1 U6164 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6464) );
  NOR2_X1 U6165 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6464), .ZN(n5014) );
  NOR2_X1 U6166 ( .A1(n6462), .A2(n5007), .ZN(n6000) );
  INV_X1 U6167 ( .A(n6015), .ZN(n5524) );
  OAI21_X1 U6168 ( .B1(REIP_REG_9__SCAN_IN), .B2(n5524), .A(n5959), .ZN(n5999)
         );
  AOI22_X1 U6169 ( .A1(EBX_REG_10__SCAN_IN), .A2(n6032), .B1(
        REIP_REG_10__SCAN_IN), .B2(n5999), .ZN(n5012) );
  INV_X1 U6170 ( .A(n5132), .ZN(n5009) );
  OAI21_X1 U6171 ( .B1(n6196), .B2(n6024), .A(n4889), .ZN(n5008) );
  AOI21_X1 U6172 ( .B1(n6044), .B2(n5009), .A(n5008), .ZN(n5011) );
  NAND2_X1 U6173 ( .A1(n6008), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5010)
         );
  NAND3_X1 U6174 ( .A1(n5012), .A2(n5011), .A3(n5010), .ZN(n5013) );
  AOI21_X1 U6175 ( .B1(n5014), .B2(n6000), .A(n5013), .ZN(n5015) );
  OAI21_X1 U6176 ( .B1(n5985), .B2(n5136), .A(n5015), .ZN(U2817) );
  INV_X1 U6177 ( .A(n5016), .ZN(n5018) );
  NOR2_X1 U6178 ( .A1(n6691), .A2(n5023), .ZN(n5048) );
  AOI21_X1 U6179 ( .B1(n5018), .B2(n5017), .A(n5048), .ZN(n5024) );
  AOI21_X1 U6180 ( .B1(n5019), .B2(STATEBS16_REG_SCAN_IN), .A(n5838), .ZN(
        n5022) );
  AOI22_X1 U6181 ( .A1(n5024), .A2(n5022), .B1(n5838), .B2(n5023), .ZN(n5020)
         );
  NAND2_X1 U6182 ( .A1(n5021), .A2(n5020), .ZN(n5047) );
  INV_X1 U6183 ( .A(n5022), .ZN(n5025) );
  OAI22_X1 U6184 ( .A1(n5025), .A2(n5024), .B1(n6522), .B2(n5023), .ZN(n5046)
         );
  AOI22_X1 U6185 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n5047), .B1(n6343), 
        .B2(n5046), .ZN(n5029) );
  NOR2_X2 U6186 ( .A1(n5027), .A2(n5026), .ZN(n5216) );
  AOI22_X1 U6187 ( .A1(n5216), .A2(n6272), .B1(n6300), .B2(n5048), .ZN(n5028)
         );
  OAI211_X1 U6188 ( .C1(n6346), .C2(n5051), .A(n5029), .B(n5028), .ZN(U3030)
         );
  AOI22_X1 U6189 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n5047), .B1(n6371), 
        .B2(n5046), .ZN(n5031) );
  AOI22_X1 U6190 ( .A1(n5216), .A2(n6280), .B1(n6279), .B2(n5048), .ZN(n5030)
         );
  OAI211_X1 U6191 ( .C1(n6374), .C2(n5051), .A(n5031), .B(n5030), .ZN(U3034)
         );
  AOI22_X1 U6192 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n5047), .B1(n6350), 
        .B2(n5046), .ZN(n5034) );
  AOI22_X1 U6193 ( .A1(n5216), .A2(n5032), .B1(n6305), .B2(n5048), .ZN(n5033)
         );
  OAI211_X1 U6194 ( .C1(n6353), .C2(n5051), .A(n5034), .B(n5033), .ZN(U3031)
         );
  AOI22_X1 U6195 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n5047), .B1(n6357), 
        .B2(n5046), .ZN(n5036) );
  AOI22_X1 U6196 ( .A1(n5216), .A2(n6276), .B1(n6275), .B2(n5048), .ZN(n5035)
         );
  OAI211_X1 U6197 ( .C1(n6360), .C2(n5051), .A(n5036), .B(n5035), .ZN(U3032)
         );
  AOI22_X1 U6198 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n5047), .B1(n6381), 
        .B2(n5046), .ZN(n5038) );
  AOI22_X1 U6199 ( .A1(n5216), .A2(n6285), .B1(n6284), .B2(n5048), .ZN(n5037)
         );
  OAI211_X1 U6200 ( .C1(n6386), .C2(n5051), .A(n5038), .B(n5037), .ZN(U3035)
         );
  AOI22_X1 U6201 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n5047), .B1(n6364), 
        .B2(n5046), .ZN(n5042) );
  AOI22_X1 U6202 ( .A1(n5216), .A2(n5040), .B1(n5039), .B2(n5048), .ZN(n5041)
         );
  OAI211_X1 U6203 ( .C1(n6367), .C2(n5051), .A(n5042), .B(n5041), .ZN(U3033)
         );
  AOI22_X1 U6204 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n5047), .B1(n6336), 
        .B2(n5046), .ZN(n5045) );
  AOI22_X1 U6205 ( .A1(n5216), .A2(n5043), .B1(n6292), .B2(n5048), .ZN(n5044)
         );
  OAI211_X1 U6206 ( .C1(n6339), .C2(n5051), .A(n5045), .B(n5044), .ZN(U3028)
         );
  AOI22_X1 U6207 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n5047), .B1(n6318), 
        .B2(n5046), .ZN(n5050) );
  AOI22_X1 U6208 ( .A1(n5216), .A2(n6269), .B1(n6296), .B2(n5048), .ZN(n5049)
         );
  OAI211_X1 U6209 ( .C1(n6321), .C2(n5051), .A(n5050), .B(n5049), .ZN(U3029)
         );
  NOR2_X1 U6210 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5052), .ZN(n5066)
         );
  INV_X1 U6211 ( .A(n5094), .ZN(n5053) );
  OAI21_X1 U6212 ( .B1(n6286), .B2(n5053), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5055) );
  AND2_X1 U6213 ( .A1(n5055), .A2(n5054), .ZN(n5059) );
  INV_X1 U6214 ( .A(n5056), .ZN(n5057) );
  AOI211_X1 U6215 ( .C1(n5829), .C2(n5059), .A(n5058), .B(n5057), .ZN(n5060)
         );
  NAND2_X1 U6216 ( .A1(n5088), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n5069) );
  INV_X1 U6217 ( .A(n5061), .ZN(n5062) );
  AOI22_X1 U6218 ( .A1(n5065), .A2(n5064), .B1(n5063), .B2(n5062), .ZN(n5090)
         );
  INV_X1 U6219 ( .A(n5066), .ZN(n5089) );
  OAI22_X1 U6220 ( .A1(n5202), .A2(n5090), .B1(n6333), .B2(n5089), .ZN(n5067)
         );
  AOI21_X1 U6221 ( .B1(n6293), .B2(n6286), .A(n5067), .ZN(n5068) );
  OAI211_X1 U6222 ( .C1(n6334), .C2(n5094), .A(n5069), .B(n5068), .ZN(U3052)
         );
  NAND2_X1 U6223 ( .A1(n5088), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5072) );
  OAI22_X1 U6224 ( .A1(n5214), .A2(n5090), .B1(n6368), .B2(n5089), .ZN(n5070)
         );
  AOI21_X1 U6225 ( .B1(n5217), .B2(n6286), .A(n5070), .ZN(n5071) );
  OAI211_X1 U6226 ( .C1(n5094), .C2(n6369), .A(n5072), .B(n5071), .ZN(U3058)
         );
  NAND2_X1 U6227 ( .A1(n5088), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n5075) );
  OAI22_X1 U6228 ( .A1(n5198), .A2(n5090), .B1(n6315), .B2(n5089), .ZN(n5073)
         );
  AOI21_X1 U6229 ( .B1(n6297), .B2(n6286), .A(n5073), .ZN(n5074) );
  OAI211_X1 U6230 ( .C1(n5094), .C2(n6316), .A(n5075), .B(n5074), .ZN(U3053)
         );
  NAND2_X1 U6231 ( .A1(n5088), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5078) );
  OAI22_X1 U6232 ( .A1(n5180), .A2(n5090), .B1(n6361), .B2(n5089), .ZN(n5076)
         );
  AOI21_X1 U6233 ( .B1(n5182), .B2(n6286), .A(n5076), .ZN(n5077) );
  OAI211_X1 U6234 ( .C1(n5094), .C2(n6362), .A(n5078), .B(n5077), .ZN(U3057)
         );
  NAND2_X1 U6235 ( .A1(n5088), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n5081) );
  OAI22_X1 U6236 ( .A1(n5190), .A2(n5090), .B1(n6347), .B2(n5089), .ZN(n5079)
         );
  AOI21_X1 U6237 ( .B1(n6308), .B2(n6286), .A(n5079), .ZN(n5080) );
  OAI211_X1 U6238 ( .C1(n5094), .C2(n6348), .A(n5081), .B(n5080), .ZN(U3055)
         );
  NAND2_X1 U6239 ( .A1(n5088), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5084) );
  OAI22_X1 U6240 ( .A1(n5185), .A2(n5090), .B1(n6354), .B2(n5089), .ZN(n5082)
         );
  AOI21_X1 U6241 ( .B1(n5187), .B2(n6286), .A(n5082), .ZN(n5083) );
  OAI211_X1 U6242 ( .C1(n5094), .C2(n6355), .A(n5084), .B(n5083), .ZN(U3056)
         );
  NAND2_X1 U6243 ( .A1(n5088), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5087) );
  OAI22_X1 U6244 ( .A1(n5194), .A2(n5090), .B1(n6340), .B2(n5089), .ZN(n5085)
         );
  AOI21_X1 U6245 ( .B1(n6301), .B2(n6286), .A(n5085), .ZN(n5086) );
  OAI211_X1 U6246 ( .C1(n5094), .C2(n6341), .A(n5087), .B(n5086), .ZN(U3054)
         );
  NAND2_X1 U6247 ( .A1(n5088), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5093) );
  OAI22_X1 U6248 ( .A1(n5206), .A2(n5090), .B1(n6376), .B2(n5089), .ZN(n5091)
         );
  AOI21_X1 U6249 ( .B1(n5208), .B2(n6286), .A(n5091), .ZN(n5092) );
  OAI211_X1 U6250 ( .C1(n5094), .C2(n6377), .A(n5093), .B(n5092), .ZN(U3059)
         );
  AND2_X1 U6251 ( .A1(n5096), .A2(n5095), .ZN(n5098) );
  OR2_X1 U6252 ( .A1(n5098), .A2(n5109), .ZN(n6150) );
  AOI22_X1 U6253 ( .A1(n5245), .A2(DATAI_11_), .B1(n6076), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n5099) );
  OAI21_X1 U6254 ( .B1(n6150), .B2(n5877), .A(n5099), .ZN(U2880) );
  NAND2_X1 U6255 ( .A1(n5101), .A2(n5100), .ZN(n5105) );
  NAND2_X1 U6256 ( .A1(n5103), .A2(n5102), .ZN(n5104) );
  XNOR2_X1 U6257 ( .A(n5105), .B(n5104), .ZN(n6212) );
  NAND2_X1 U6258 ( .A1(n6212), .A2(n6178), .ZN(n5108) );
  NAND2_X1 U6259 ( .A1(n6189), .A2(REIP_REG_9__SCAN_IN), .ZN(n6208) );
  OAI21_X1 U6260 ( .B1(n5684), .B2(n5994), .A(n6208), .ZN(n5106) );
  AOI21_X1 U6261 ( .B1(n5883), .B2(n5998), .A(n5106), .ZN(n5107) );
  OAI211_X1 U6262 ( .C1(n6164), .C2(n5997), .A(n5108), .B(n5107), .ZN(U2977)
         );
  XOR2_X1 U6263 ( .A(n5110), .B(n5109), .Z(n5976) );
  INV_X1 U6264 ( .A(n5976), .ZN(n5116) );
  AOI22_X1 U6265 ( .A1(n5245), .A2(DATAI_12_), .B1(n6076), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n5111) );
  OAI21_X1 U6266 ( .B1(n5116), .B2(n5877), .A(n5111), .ZN(U2879) );
  INV_X1 U6267 ( .A(n5163), .ZN(n5113) );
  XNOR2_X1 U6268 ( .A(n5114), .B(n5113), .ZN(n6187) );
  AOI22_X1 U6269 ( .A1(n6060), .A2(n6187), .B1(EBX_REG_12__SCAN_IN), .B2(n5549), .ZN(n5115) );
  OAI21_X1 U6270 ( .B1(n5116), .B2(n6056), .A(n5115), .ZN(U2847) );
  INV_X1 U6271 ( .A(n5117), .ZN(n5837) );
  NAND2_X1 U6272 ( .A1(n6032), .A2(EBX_REG_2__SCAN_IN), .ZN(n5120) );
  INV_X1 U6273 ( .A(REIP_REG_2__SCAN_IN), .ZN(n5124) );
  NAND3_X1 U6274 ( .A1(n5118), .A2(REIP_REG_1__SCAN_IN), .A3(n5124), .ZN(n5119) );
  OAI211_X1 U6275 ( .C1(n5837), .C2(n5121), .A(n5120), .B(n5119), .ZN(n5126)
         );
  OR2_X1 U6276 ( .A1(n6021), .A2(REIP_REG_1__SCAN_IN), .ZN(n5122) );
  AND2_X1 U6277 ( .A1(n5123), .A2(n5122), .ZN(n6031) );
  OAI22_X1 U6278 ( .A1(n6030), .A2(n6181), .B1(n6031), .B2(n5124), .ZN(n5125)
         );
  AOI211_X1 U6279 ( .C1(PHYADDRPOINTER_REG_2__SCAN_IN), .C2(n6008), .A(n5126), 
        .B(n5125), .ZN(n5128) );
  NAND2_X1 U6280 ( .A1(n6259), .A2(n6033), .ZN(n5127) );
  OAI211_X1 U6281 ( .C1(n6175), .C2(n6041), .A(n5128), .B(n5127), .ZN(U2825)
         );
  XNOR2_X1 U6282 ( .A(n5673), .B(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5130)
         );
  XNOR2_X1 U6283 ( .A(n5152), .B(n5130), .ZN(n6204) );
  NAND2_X1 U6284 ( .A1(n6204), .A2(n6178), .ZN(n5135) );
  INV_X1 U6285 ( .A(REIP_REG_10__SCAN_IN), .ZN(n5131) );
  NOR2_X1 U6286 ( .A1(n4889), .A2(n5131), .ZN(n6197) );
  NOR2_X1 U6287 ( .A1(n6182), .A2(n5132), .ZN(n5133) );
  AOI211_X1 U6288 ( .C1(n6171), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6197), 
        .B(n5133), .ZN(n5134) );
  OAI211_X1 U6289 ( .C1(n6164), .C2(n5136), .A(n5135), .B(n5134), .ZN(U2976)
         );
  NAND2_X1 U6290 ( .A1(n2968), .A2(n5279), .ZN(n5138) );
  XNOR2_X1 U6291 ( .A(n5139), .B(n5138), .ZN(n6188) );
  INV_X1 U6292 ( .A(n6188), .ZN(n5143) );
  AOI22_X1 U6293 ( .A1(n6171), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .B1(n6189), 
        .B2(REIP_REG_12__SCAN_IN), .ZN(n5140) );
  OAI21_X1 U6294 ( .B1(n6182), .B2(n5974), .A(n5140), .ZN(n5141) );
  AOI21_X1 U6295 ( .B1(n5976), .B2(n6176), .A(n5141), .ZN(n5142) );
  OAI21_X1 U6296 ( .B1(n5143), .B2(n6166), .A(n5142), .ZN(U2974) );
  INV_X1 U6297 ( .A(n5144), .ZN(n5147) );
  INV_X1 U6298 ( .A(n5145), .ZN(n5146) );
  NAND2_X1 U6299 ( .A1(n5147), .A2(n5146), .ZN(n5149) );
  AND2_X1 U6300 ( .A1(n5149), .A2(n5148), .ZN(n6051) );
  INV_X1 U6301 ( .A(n6051), .ZN(n5151) );
  AOI22_X1 U6302 ( .A1(n5245), .A2(DATAI_13_), .B1(n6076), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n5150) );
  OAI21_X1 U6303 ( .B1(n5151), .B2(n5877), .A(n5150), .ZN(U2878) );
  OR2_X1 U6304 ( .A1(n5152), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5153)
         );
  AOI22_X1 U6305 ( .A1(n5153), .A2(n5673), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n5152), .ZN(n5155) );
  XNOR2_X1 U6306 ( .A(n5673), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5154)
         );
  XNOR2_X1 U6307 ( .A(n5155), .B(n5154), .ZN(n6154) );
  NOR2_X1 U6308 ( .A1(n6655), .A2(n5156), .ZN(n6194) );
  NAND2_X1 U6309 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6219) );
  INV_X1 U6310 ( .A(n6219), .ZN(n6202) );
  NAND4_X1 U6311 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n6194), .A4(n6202), .ZN(n5162)
         );
  NOR3_X1 U6312 ( .A1(n6257), .A2(n5157), .A3(n5162), .ZN(n5360) );
  NOR2_X1 U6313 ( .A1(n5158), .A2(n6260), .ZN(n5359) );
  INV_X1 U6314 ( .A(n6255), .ZN(n5159) );
  NOR2_X1 U6315 ( .A1(n5159), .A2(n5162), .ZN(n5355) );
  INV_X1 U6316 ( .A(n5355), .ZN(n5160) );
  NOR2_X1 U6317 ( .A1(n6199), .A2(n5160), .ZN(n5821) );
  OAI22_X1 U6318 ( .A1(n5771), .A2(n5360), .B1(n5359), .B2(n5821), .ZN(n6183)
         );
  NOR2_X1 U6319 ( .A1(n5162), .A2(n5161), .ZN(n6184) );
  AOI22_X1 U6320 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n6183), .B1(n6186), .B2(n6574), .ZN(n5167) );
  AOI21_X1 U6321 ( .B1(n5165), .B2(n5164), .A(n5163), .ZN(n6053) );
  AOI22_X1 U6322 ( .A1(n6258), .A2(n6053), .B1(n6018), .B2(
        REIP_REG_11__SCAN_IN), .ZN(n5166) );
  OAI211_X1 U6323 ( .C1(n6154), .C2(n6242), .A(n5167), .B(n5166), .ZN(U3007)
         );
  NOR2_X1 U6324 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5168), .ZN(n5179)
         );
  INV_X1 U6325 ( .A(n6291), .ZN(n5170) );
  OAI21_X1 U6326 ( .B1(n5170), .B2(n5216), .A(n5169), .ZN(n5172) );
  INV_X1 U6327 ( .A(n5178), .ZN(n5171) );
  NAND2_X1 U6328 ( .A1(n5172), .A2(n5171), .ZN(n5174) );
  OAI221_X1 U6329 ( .B1(n5179), .B2(n6512), .C1(n5179), .C2(n5174), .A(n5173), 
        .ZN(n5211) );
  NAND2_X1 U6330 ( .A1(n5211), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5184) );
  NOR2_X1 U6331 ( .A1(n5175), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5176)
         );
  AOI22_X1 U6332 ( .A1(n5178), .A2(n5829), .B1(n5177), .B2(n5176), .ZN(n5213)
         );
  INV_X1 U6333 ( .A(n5179), .ZN(n5212) );
  OAI22_X1 U6334 ( .A1(n5180), .A2(n5213), .B1(n6361), .B2(n5212), .ZN(n5181)
         );
  AOI21_X1 U6335 ( .B1(n5182), .B2(n5216), .A(n5181), .ZN(n5183) );
  OAI211_X1 U6336 ( .C1(n6291), .C2(n6362), .A(n5184), .B(n5183), .ZN(U3041)
         );
  NAND2_X1 U6337 ( .A1(n5211), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5189) );
  OAI22_X1 U6338 ( .A1(n5185), .A2(n5213), .B1(n6354), .B2(n5212), .ZN(n5186)
         );
  AOI21_X1 U6339 ( .B1(n5187), .B2(n5216), .A(n5186), .ZN(n5188) );
  OAI211_X1 U6340 ( .C1(n6291), .C2(n6355), .A(n5189), .B(n5188), .ZN(U3040)
         );
  NAND2_X1 U6341 ( .A1(n5211), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5193) );
  OAI22_X1 U6342 ( .A1(n5190), .A2(n5213), .B1(n6347), .B2(n5212), .ZN(n5191)
         );
  AOI21_X1 U6343 ( .B1(n6308), .B2(n5216), .A(n5191), .ZN(n5192) );
  OAI211_X1 U6344 ( .C1(n6291), .C2(n6348), .A(n5193), .B(n5192), .ZN(U3039)
         );
  NAND2_X1 U6345 ( .A1(n5211), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5197) );
  OAI22_X1 U6346 ( .A1(n5194), .A2(n5213), .B1(n6340), .B2(n5212), .ZN(n5195)
         );
  AOI21_X1 U6347 ( .B1(n6301), .B2(n5216), .A(n5195), .ZN(n5196) );
  OAI211_X1 U6348 ( .C1(n6291), .C2(n6341), .A(n5197), .B(n5196), .ZN(U3038)
         );
  NAND2_X1 U6349 ( .A1(n5211), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5201) );
  OAI22_X1 U6350 ( .A1(n5198), .A2(n5213), .B1(n6315), .B2(n5212), .ZN(n5199)
         );
  AOI21_X1 U6351 ( .B1(n6297), .B2(n5216), .A(n5199), .ZN(n5200) );
  OAI211_X1 U6352 ( .C1(n6291), .C2(n6316), .A(n5201), .B(n5200), .ZN(U3037)
         );
  NAND2_X1 U6353 ( .A1(n5211), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5205) );
  OAI22_X1 U6354 ( .A1(n5202), .A2(n5213), .B1(n6333), .B2(n5212), .ZN(n5203)
         );
  AOI21_X1 U6355 ( .B1(n6293), .B2(n5216), .A(n5203), .ZN(n5204) );
  OAI211_X1 U6356 ( .C1(n6334), .C2(n6291), .A(n5205), .B(n5204), .ZN(U3036)
         );
  NAND2_X1 U6357 ( .A1(n5211), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5210) );
  OAI22_X1 U6358 ( .A1(n5206), .A2(n5213), .B1(n6376), .B2(n5212), .ZN(n5207)
         );
  AOI21_X1 U6359 ( .B1(n5208), .B2(n5216), .A(n5207), .ZN(n5209) );
  OAI211_X1 U6360 ( .C1(n6291), .C2(n6377), .A(n5210), .B(n5209), .ZN(U3043)
         );
  NAND2_X1 U6361 ( .A1(n5211), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5219) );
  OAI22_X1 U6362 ( .A1(n5214), .A2(n5213), .B1(n6368), .B2(n5212), .ZN(n5215)
         );
  AOI21_X1 U6363 ( .B1(n5217), .B2(n5216), .A(n5215), .ZN(n5218) );
  OAI211_X1 U6364 ( .C1(n6291), .C2(n6369), .A(n5219), .B(n5218), .ZN(U3042)
         );
  OR2_X1 U6365 ( .A1(n5222), .A2(n5221), .ZN(n5223) );
  NAND2_X1 U6366 ( .A1(n5237), .A2(n5223), .ZN(n5287) );
  AOI22_X1 U6367 ( .A1(n5245), .A2(DATAI_14_), .B1(n6076), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5224) );
  OAI21_X1 U6368 ( .B1(n5287), .B2(n5877), .A(n5224), .ZN(U2877) );
  NAND2_X1 U6369 ( .A1(n6015), .A2(n5225), .ZN(n5248) );
  INV_X1 U6370 ( .A(n5248), .ZN(n5234) );
  OAI21_X1 U6371 ( .B1(n5226), .B2(n5910), .A(n5242), .ZN(n5815) );
  NAND2_X1 U6372 ( .A1(n6044), .A2(n5284), .ZN(n5230) );
  NOR3_X1 U6373 ( .A1(n6021), .A2(REIP_REG_14__SCAN_IN), .A3(n5227), .ZN(n5228) );
  AOI21_X1 U6374 ( .B1(n6032), .B2(EBX_REG_14__SCAN_IN), .A(n5228), .ZN(n5229)
         );
  OAI211_X1 U6375 ( .C1(n5815), .C2(n6024), .A(n5230), .B(n5229), .ZN(n5233)
         );
  OAI21_X1 U6376 ( .B1(n6036), .B2(n5231), .A(n4889), .ZN(n5232) );
  AOI211_X1 U6377 ( .C1(n5234), .C2(REIP_REG_14__SCAN_IN), .A(n5233), .B(n5232), .ZN(n5235) );
  OAI21_X1 U6378 ( .B1(n5287), .B2(n5985), .A(n5235), .ZN(U2813) );
  INV_X1 U6379 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5236) );
  OAI222_X1 U6380 ( .A1(n5287), .A2(n6056), .B1(n5236), .B2(n6065), .C1(n5815), 
        .C2(n6055), .ZN(U2845) );
  INV_X1 U6381 ( .A(n5237), .ZN(n5240) );
  INV_X1 U6382 ( .A(n5238), .ZN(n5239) );
  OAI21_X1 U6383 ( .B1(n5240), .B2(n5239), .A(n5255), .ZN(n5278) );
  AOI21_X1 U6384 ( .B1(n5243), .B2(n5242), .A(n5773), .ZN(n5900) );
  AOI22_X1 U6385 ( .A1(n6060), .A2(n5900), .B1(n5549), .B2(EBX_REG_15__SCAN_IN), .ZN(n5244) );
  OAI21_X1 U6386 ( .B1(n5278), .B2(n6056), .A(n5244), .ZN(U2844) );
  AOI22_X1 U6387 ( .A1(n5245), .A2(DATAI_15_), .B1(n6076), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5246) );
  OAI21_X1 U6388 ( .B1(n5278), .B2(n5877), .A(n5246), .ZN(U2876) );
  AOI21_X1 U6389 ( .B1(n6008), .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n6018), 
        .ZN(n5247) );
  OAI221_X1 U6390 ( .B1(REIP_REG_15__SCAN_IN), .B2(n5249), .C1(n6673), .C2(
        n5248), .A(n5247), .ZN(n5252) );
  AOI22_X1 U6391 ( .A1(n5900), .A2(n6033), .B1(n6032), .B2(EBX_REG_15__SCAN_IN), .ZN(n5250) );
  OAI21_X1 U6392 ( .B1(n6030), .B2(n5274), .A(n5250), .ZN(n5251) );
  NOR2_X1 U6393 ( .A1(n5252), .A2(n5251), .ZN(n5253) );
  OAI21_X1 U6394 ( .B1(n5278), .B2(n5985), .A(n5253), .ZN(U2812) );
  AND2_X1 U6395 ( .A1(n5255), .A2(n5254), .ZN(n5256) );
  OR2_X1 U6396 ( .A1(n5256), .A2(n5291), .ZN(n6072) );
  AND2_X1 U6397 ( .A1(n5257), .A2(n5773), .ZN(n5300) );
  NOR2_X1 U6398 ( .A1(n5257), .A2(n5773), .ZN(n5258) );
  OR2_X1 U6399 ( .A1(n5300), .A2(n5258), .ZN(n5891) );
  NAND2_X1 U6400 ( .A1(n6008), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5259)
         );
  OAI211_X1 U6401 ( .C1(n5891), .C2(n6024), .A(n5259), .B(n4889), .ZN(n5265)
         );
  NAND2_X1 U6402 ( .A1(n6015), .A2(REIP_REG_16__SCAN_IN), .ZN(n5262) );
  INV_X1 U6403 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6476) );
  AOI22_X1 U6404 ( .A1(EBX_REG_16__SCAN_IN), .A2(n6032), .B1(n5260), .B2(n6476), .ZN(n5261) );
  OAI21_X1 U6405 ( .B1(n5263), .B2(n5262), .A(n5261), .ZN(n5264) );
  AOI211_X1 U6406 ( .C1(n5687), .C2(n6044), .A(n5265), .B(n5264), .ZN(n5266)
         );
  OAI21_X1 U6407 ( .B1(n6072), .B2(n5985), .A(n5266), .ZN(U2811) );
  INV_X1 U6408 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5267) );
  OAI222_X1 U6409 ( .A1(n6072), .A2(n6056), .B1(n5267), .B2(n6065), .C1(n6055), 
        .C2(n5891), .ZN(U2843) );
  NAND2_X1 U6410 ( .A1(n5268), .A2(n5269), .ZN(n5271) );
  NAND2_X1 U6411 ( .A1(n5271), .A2(n5270), .ZN(n5273) );
  XNOR2_X1 U6412 ( .A(n4079), .B(n5906), .ZN(n5272) );
  XNOR2_X1 U6413 ( .A(n5273), .B(n5272), .ZN(n5903) );
  NAND2_X1 U6414 ( .A1(n5903), .A2(n6178), .ZN(n5277) );
  NOR2_X1 U6415 ( .A1(n4889), .A2(n6673), .ZN(n5899) );
  NOR2_X1 U6416 ( .A1(n6182), .A2(n5274), .ZN(n5275) );
  AOI211_X1 U6417 ( .C1(n6171), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n5899), 
        .B(n5275), .ZN(n5276) );
  OAI211_X1 U6418 ( .C1(n6164), .C2(n5278), .A(n5277), .B(n5276), .ZN(U2971)
         );
  NAND2_X1 U6419 ( .A1(n5268), .A2(n5279), .ZN(n5888) );
  NAND2_X1 U6420 ( .A1(n5888), .A2(n5887), .ZN(n5281) );
  NAND2_X1 U6421 ( .A1(n5281), .A2(n5280), .ZN(n5283) );
  XNOR2_X1 U6422 ( .A(n4079), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5282)
         );
  XNOR2_X1 U6423 ( .A(n5283), .B(n5282), .ZN(n5814) );
  AOI22_X1 U6424 ( .A1(n6171), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n6018), 
        .B2(REIP_REG_14__SCAN_IN), .ZN(n5286) );
  NAND2_X1 U6425 ( .A1(n5883), .A2(n5284), .ZN(n5285) );
  OAI211_X1 U6426 ( .C1(n5287), .C2(n6164), .A(n5286), .B(n5285), .ZN(n5288)
         );
  AOI21_X1 U6427 ( .B1(n5814), .B2(n6178), .A(n5288), .ZN(n5289) );
  INV_X1 U6428 ( .A(n5289), .ZN(U2972) );
  NOR2_X1 U6429 ( .A1(n5291), .A2(n5290), .ZN(n5292) );
  OR2_X1 U6430 ( .A1(n5553), .A2(n5292), .ZN(n5881) );
  AOI21_X1 U6431 ( .B1(n6478), .B2(n5293), .A(n5524), .ZN(n5297) );
  OAI22_X1 U6432 ( .A1(n6615), .A2(n6005), .B1(n5294), .B2(n6036), .ZN(n5295)
         );
  AOI211_X1 U6433 ( .C1(n5297), .C2(n5296), .A(n6018), .B(n5295), .ZN(n5304)
         );
  NAND2_X1 U6434 ( .A1(n5773), .A2(n5298), .ZN(n5556) );
  OR2_X1 U6435 ( .A1(n5300), .A2(n5299), .ZN(n5301) );
  NAND2_X1 U6436 ( .A1(n5556), .A2(n5301), .ZN(n5808) );
  INV_X1 U6437 ( .A(n5808), .ZN(n5302) );
  AOI22_X1 U6438 ( .A1(n6044), .A2(n5882), .B1(n5302), .B2(n6033), .ZN(n5303)
         );
  OAI211_X1 U6439 ( .C1(n5881), .C2(n5985), .A(n5304), .B(n5303), .ZN(U2810)
         );
  OAI222_X1 U6440 ( .A1(n5881), .A2(n6056), .B1(n6615), .B2(n6065), .C1(n5808), 
        .C2(n6055), .ZN(U2842) );
  AND2_X1 U6441 ( .A1(n5305), .A2(n5555), .ZN(n5461) );
  OAI21_X1 U6442 ( .B1(n5461), .B2(n5306), .A(n5433), .ZN(n5452) );
  NOR2_X2 U6443 ( .A1(n6076), .A2(n5307), .ZN(n6073) );
  AOI22_X1 U6444 ( .A1(n6073), .A2(DATAI_29_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n6076), .ZN(n5312) );
  AND2_X1 U6445 ( .A1(n5309), .A2(n5308), .ZN(n5310) );
  NAND2_X1 U6446 ( .A1(n6077), .A2(DATAI_13_), .ZN(n5311) );
  OAI211_X1 U6447 ( .C1(n5452), .C2(n5877), .A(n5312), .B(n5311), .ZN(U2862)
         );
  NAND2_X1 U6448 ( .A1(n5313), .A2(n5530), .ZN(n5316) );
  INV_X1 U6449 ( .A(n5314), .ZN(n5315) );
  NAND2_X1 U6450 ( .A1(n5316), .A2(n5315), .ZN(n5317) );
  NOR2_X1 U6451 ( .A1(n5417), .A2(n5317), .ZN(n5318) );
  NOR2_X1 U6452 ( .A1(n5319), .A2(n5318), .ZN(n5708) );
  AOI22_X1 U6453 ( .A1(n5708), .A2(n6060), .B1(EBX_REG_29__SCAN_IN), .B2(n5549), .ZN(n5320) );
  OAI21_X1 U6454 ( .B1(n5452), .B2(n6056), .A(n5320), .ZN(U2830) );
  NAND2_X1 U6455 ( .A1(n5555), .A2(n5322), .ZN(n5487) );
  OAI21_X1 U6456 ( .B1(n5377), .B2(n5323), .A(n5487), .ZN(n5338) );
  INV_X1 U6457 ( .A(n5338), .ZN(n5641) );
  XNOR2_X1 U6458 ( .A(REIP_REG_24__SCAN_IN), .B(REIP_REG_25__SCAN_IN), .ZN(
        n5324) );
  NOR2_X1 U6459 ( .A1(n5508), .A2(n5324), .ZN(n5333) );
  NAND2_X1 U6460 ( .A1(n5325), .A2(n6015), .ZN(n5850) );
  INV_X1 U6461 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6492) );
  NAND2_X1 U6462 ( .A1(n5373), .A2(n5327), .ZN(n5328) );
  NAND2_X1 U6463 ( .A1(n5491), .A2(n5328), .ZN(n5740) );
  INV_X1 U6464 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5335) );
  OAI22_X1 U6465 ( .A1(n5740), .A2(n6024), .B1(n6005), .B2(n5335), .ZN(n5329)
         );
  AOI21_X1 U6466 ( .B1(n5637), .B2(n6044), .A(n5329), .ZN(n5331) );
  NAND2_X1 U6467 ( .A1(n6008), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5330)
         );
  OAI211_X1 U6468 ( .C1(n5850), .C2(n6492), .A(n5331), .B(n5330), .ZN(n5332)
         );
  AOI211_X1 U6469 ( .C1(n5641), .C2(n3979), .A(n5333), .B(n5332), .ZN(n5334)
         );
  INV_X1 U6470 ( .A(n5334), .ZN(U2802) );
  OAI222_X1 U6471 ( .A1(n5338), .A2(n6056), .B1(n5335), .B2(n6065), .C1(n5740), 
        .C2(n6055), .ZN(U2834) );
  AOI22_X1 U6472 ( .A1(n6073), .A2(DATAI_25_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n6076), .ZN(n5337) );
  NAND2_X1 U6473 ( .A1(n6077), .A2(DATAI_9_), .ZN(n5336) );
  OAI211_X1 U6474 ( .C1(n5338), .C2(n5877), .A(n5337), .B(n5336), .ZN(U2866)
         );
  INV_X1 U6475 ( .A(n5643), .ZN(n5339) );
  OAI21_X1 U6476 ( .B1(n5673), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5339), 
        .ZN(n5351) );
  AOI21_X1 U6477 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n4079), .A(n5340), 
        .ZN(n5341) );
  XNOR2_X1 U6478 ( .A(n5351), .B(n5341), .ZN(n5757) );
  NOR2_X1 U6479 ( .A1(n5655), .A2(n5342), .ZN(n5542) );
  NOR2_X1 U6480 ( .A1(n5542), .A2(n5343), .ZN(n5344) );
  INV_X1 U6481 ( .A(n5582), .ZN(n5348) );
  NAND2_X1 U6482 ( .A1(n6018), .A2(REIP_REG_22__SCAN_IN), .ZN(n5752) );
  NAND2_X1 U6483 ( .A1(n6171), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5346)
         );
  OAI211_X1 U6484 ( .C1(n6182), .C2(n5515), .A(n5752), .B(n5346), .ZN(n5347)
         );
  AOI21_X1 U6485 ( .B1(n5348), .B2(n6176), .A(n5347), .ZN(n5349) );
  OAI21_X1 U6486 ( .B1(n5757), .B2(n6166), .A(n5349), .ZN(U2964) );
  NAND3_X1 U6487 ( .A1(n5409), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5350) );
  XNOR2_X1 U6488 ( .A(n5353), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5384)
         );
  NAND2_X1 U6489 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6185) );
  NOR2_X1 U6490 ( .A1(n5354), .A2(n6185), .ZN(n5820) );
  NAND2_X1 U6491 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5820), .ZN(n5901) );
  NAND2_X1 U6492 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5894) );
  NOR2_X1 U6493 ( .A1(n5901), .A2(n5894), .ZN(n5781) );
  NAND2_X1 U6494 ( .A1(n5781), .A2(n5355), .ZN(n5767) );
  INV_X1 U6495 ( .A(n5767), .ZN(n5357) );
  NAND4_X1 U6496 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A3(INSTADDRPOINTER_REG_19__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5361) );
  INV_X1 U6497 ( .A(n5361), .ZN(n5356) );
  NAND2_X1 U6498 ( .A1(n5357), .A2(n5356), .ZN(n5358) );
  NOR2_X1 U6499 ( .A1(n6199), .A2(n5358), .ZN(n5368) );
  OR2_X1 U6500 ( .A1(n5359), .A2(n5368), .ZN(n5363) );
  NAND2_X1 U6501 ( .A1(n5360), .A2(n5781), .ZN(n5766) );
  NOR2_X1 U6502 ( .A1(n5766), .A2(n5361), .ZN(n5367) );
  OR2_X1 U6503 ( .A1(n5771), .A2(n5367), .ZN(n5362) );
  NAND2_X1 U6504 ( .A1(n5363), .A2(n5362), .ZN(n5763) );
  INV_X1 U6505 ( .A(n5750), .ZN(n5364) );
  AND2_X1 U6506 ( .A1(n6201), .A2(n5364), .ZN(n5365) );
  NOR2_X1 U6507 ( .A1(n5763), .A2(n5365), .ZN(n5399) );
  AND2_X1 U6508 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5404) );
  INV_X1 U6509 ( .A(n5404), .ZN(n5421) );
  OAI21_X1 U6510 ( .B1(n6254), .B2(n6260), .A(n5421), .ZN(n5366) );
  NAND2_X1 U6511 ( .A1(n5399), .A2(n5366), .ZN(n5746) );
  NAND2_X1 U6512 ( .A1(n6254), .A2(n5367), .ZN(n5370) );
  INV_X1 U6513 ( .A(n5368), .ZN(n5369) );
  NAND2_X1 U6514 ( .A1(n5370), .A2(n5369), .ZN(n5759) );
  NAND2_X1 U6515 ( .A1(n5759), .A2(n5750), .ZN(n5422) );
  INV_X1 U6516 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5401) );
  OAI21_X1 U6517 ( .B1(n5422), .B2(n5400), .A(n5401), .ZN(n5375) );
  OR2_X1 U6518 ( .A1(n5394), .A2(n5371), .ZN(n5372) );
  NAND2_X1 U6519 ( .A1(n5373), .A2(n5372), .ZN(n5539) );
  NAND2_X1 U6520 ( .A1(n6189), .A2(REIP_REG_24__SCAN_IN), .ZN(n5380) );
  OAI21_X1 U6521 ( .B1(n5539), .B2(n6246), .A(n5380), .ZN(n5374) );
  AOI21_X1 U6522 ( .B1(n5746), .B2(n5375), .A(n5374), .ZN(n5376) );
  OAI21_X1 U6523 ( .B1(n5384), .B2(n6242), .A(n5376), .ZN(U2994) );
  NAND2_X1 U6524 ( .A1(n5883), .A2(n5505), .ZN(n5381) );
  OAI211_X1 U6525 ( .C1(n5502), .C2(n5684), .A(n5381), .B(n5380), .ZN(n5382)
         );
  AOI21_X1 U6526 ( .B1(n5538), .B2(n6176), .A(n5382), .ZN(n5383) );
  OAI21_X1 U6527 ( .B1(n5384), .B2(n6166), .A(n5383), .ZN(U2962) );
  OR2_X1 U6528 ( .A1(n5386), .A2(n5385), .ZN(n5388) );
  NAND2_X1 U6529 ( .A1(n5388), .A2(n5387), .ZN(n6236) );
  INV_X1 U6530 ( .A(n6236), .ZN(n5389) );
  AOI22_X1 U6531 ( .A1(n6060), .A2(n5389), .B1(n5549), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n5390) );
  OAI21_X1 U6532 ( .B1(n6165), .B2(n6056), .A(n5390), .ZN(U2855) );
  NAND2_X1 U6533 ( .A1(n5391), .A2(n6263), .ZN(n5398) );
  AND2_X1 U6534 ( .A1(n5513), .A2(n5392), .ZN(n5393) );
  NOR2_X1 U6535 ( .A1(n5394), .A2(n5393), .ZN(n5848) );
  NOR2_X1 U6536 ( .A1(n5422), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5395)
         );
  AOI211_X1 U6537 ( .C1(n6258), .C2(n5848), .A(n5396), .B(n5395), .ZN(n5397)
         );
  OAI211_X1 U6538 ( .C1(n5399), .C2(n5400), .A(n5398), .B(n5397), .ZN(U2995)
         );
  NOR2_X1 U6539 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5782) );
  NOR2_X1 U6540 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5749) );
  NAND4_X1 U6541 ( .A1(n5782), .A2(n5749), .A3(n5401), .A4(n5400), .ZN(n5402)
         );
  NAND2_X1 U6542 ( .A1(n5673), .A2(n5402), .ZN(n5403) );
  AND2_X1 U6543 ( .A1(n5660), .A2(n5403), .ZN(n5406) );
  NAND3_X1 U6544 ( .A1(n5404), .A2(n5750), .A3(n5783), .ZN(n5405) );
  AOI21_X2 U6545 ( .B1(n5661), .B2(n5406), .A(n2962), .ZN(n5635) );
  INV_X1 U6546 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5407) );
  XNOR2_X1 U6547 ( .A(n4079), .B(n5407), .ZN(n5636) );
  OR2_X2 U6548 ( .A1(n5635), .A2(n5636), .ZN(n5588) );
  NAND2_X1 U6549 ( .A1(n4079), .A2(n5407), .ZN(n5408) );
  OR2_X1 U6550 ( .A1(n5409), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5626)
         );
  INV_X1 U6551 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5716) );
  NAND2_X1 U6552 ( .A1(n5610), .A2(n5716), .ZN(n5410) );
  NOR2_X1 U6553 ( .A1(n5626), .A2(n5410), .ZN(n5591) );
  NAND2_X1 U6554 ( .A1(n5627), .A2(n5591), .ZN(n5600) );
  NAND2_X1 U6555 ( .A1(n4079), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5625) );
  AND2_X1 U6556 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5424) );
  NAND2_X1 U6557 ( .A1(n5618), .A2(n5424), .ZN(n5601) );
  MUX2_X2 U6558 ( .A(n5600), .B(n5601), .S(INSTADDRPOINTER_REG_29__SCAN_IN), 
        .Z(n5412) );
  INV_X1 U6559 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5590) );
  XNOR2_X1 U6560 ( .A(n5412), .B(n5590), .ZN(n5437) );
  NAND2_X1 U6561 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5423) );
  AOI21_X1 U6562 ( .B1(n6201), .B2(n5423), .A(n5746), .ZN(n5720) );
  OAI21_X1 U6563 ( .B1(n6203), .B2(n5424), .A(n5720), .ZN(n5712) );
  AOI21_X1 U6564 ( .B1(n6201), .B2(n5589), .A(n5712), .ZN(n5697) );
  INV_X1 U6565 ( .A(n5697), .ZN(n5428) );
  INV_X1 U6566 ( .A(n5417), .ZN(n5463) );
  INV_X1 U6567 ( .A(n5415), .ZN(n5413) );
  OAI21_X1 U6568 ( .B1(n5414), .B2(n5463), .A(n5413), .ZN(n5419) );
  INV_X1 U6569 ( .A(n5414), .ZN(n5416) );
  OAI211_X1 U6570 ( .C1(n5417), .C2(n5530), .A(n5416), .B(n5415), .ZN(n5418)
         );
  OAI21_X1 U6571 ( .B1(n5420), .B2(n5419), .A(n5418), .ZN(n5449) );
  OR2_X1 U6572 ( .A1(n5422), .A2(n5421), .ZN(n5744) );
  OR2_X1 U6573 ( .A1(n5744), .A2(n5423), .ZN(n5721) );
  INV_X1 U6574 ( .A(n5424), .ZN(n5425) );
  NOR2_X1 U6575 ( .A1(n5721), .A2(n5425), .ZN(n5706) );
  NAND3_X1 U6576 ( .A1(n5706), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5590), .ZN(n5426) );
  NAND2_X1 U6577 ( .A1(n6018), .A2(REIP_REG_30__SCAN_IN), .ZN(n5431) );
  OAI211_X1 U6578 ( .C1(n6246), .C2(n5449), .A(n5426), .B(n5431), .ZN(n5427)
         );
  AOI21_X1 U6579 ( .B1(n5428), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5427), 
        .ZN(n5429) );
  OAI21_X1 U6580 ( .B1(n5437), .B2(n6242), .A(n5429), .ZN(U2988) );
  OAI22_X1 U6581 ( .A1(n5701), .A2(n6055), .B1(n6065), .B2(n5430), .ZN(U2828)
         );
  OAI21_X1 U6582 ( .B1(n5684), .B2(n6571), .A(n5431), .ZN(n5435) );
  NOR2_X1 U6583 ( .A1(n5438), .A2(n6164), .ZN(n5434) );
  OAI21_X1 U6584 ( .B1(n5437), .B2(n6166), .A(n5436), .ZN(U2956) );
  INV_X1 U6585 ( .A(n5439), .ZN(n5445) );
  AOI22_X1 U6586 ( .A1(n6008), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .B1(
        EBX_REG_30__SCAN_IN), .B2(n6032), .ZN(n5442) );
  NAND2_X1 U6587 ( .A1(n6044), .A2(n5440), .ZN(n5441) );
  OAI211_X1 U6588 ( .C1(n5449), .C2(n6024), .A(n5442), .B(n5441), .ZN(n5444)
         );
  NOR3_X1 U6589 ( .A1(n5459), .A2(REIP_REG_30__SCAN_IN), .A3(n6501), .ZN(n5443) );
  AOI211_X1 U6590 ( .C1(REIP_REG_30__SCAN_IN), .C2(n5445), .A(n5444), .B(n5443), .ZN(n5446) );
  OAI21_X1 U6591 ( .B1(n5451), .B2(n5985), .A(n5446), .ZN(U2797) );
  AOI22_X1 U6592 ( .A1(n6073), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n6076), .ZN(n5448) );
  NAND2_X1 U6593 ( .A1(n6077), .A2(DATAI_14_), .ZN(n5447) );
  OAI211_X1 U6594 ( .C1(n5451), .C2(n5877), .A(n5448), .B(n5447), .ZN(U2861)
         );
  INV_X1 U6595 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5450) );
  OAI222_X1 U6596 ( .A1(n6056), .A2(n5451), .B1(n5450), .B2(n6065), .C1(n5449), 
        .C2(n6055), .ZN(U2829) );
  INV_X1 U6597 ( .A(n5452), .ZN(n5606) );
  NAND2_X1 U6598 ( .A1(n5606), .A2(n3979), .ZN(n5458) );
  INV_X1 U6599 ( .A(n5453), .ZN(n5604) );
  NAND2_X1 U6600 ( .A1(n5708), .A2(n6033), .ZN(n5455) );
  AOI22_X1 U6601 ( .A1(n6008), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .B1(n6032), 
        .B2(EBX_REG_29__SCAN_IN), .ZN(n5454) );
  OAI211_X1 U6602 ( .C1(n6030), .C2(n5604), .A(n5455), .B(n5454), .ZN(n5456)
         );
  AOI21_X1 U6603 ( .B1(n5468), .B2(REIP_REG_29__SCAN_IN), .A(n5456), .ZN(n5457) );
  OAI211_X1 U6604 ( .C1(REIP_REG_29__SCAN_IN), .C2(n5459), .A(n5458), .B(n5457), .ZN(U2798) );
  NAND2_X1 U6605 ( .A1(n5555), .A2(n5460), .ZN(n5473) );
  AOI21_X1 U6606 ( .B1(n5462), .B2(n5473), .A(n5461), .ZN(n5615) );
  INV_X1 U6607 ( .A(n5615), .ZN(n5568) );
  OAI21_X1 U6608 ( .B1(n5478), .B2(n5464), .A(n5463), .ZN(n5715) );
  INV_X1 U6609 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5535) );
  OAI22_X1 U6610 ( .A1(n5715), .A2(n6024), .B1(n6005), .B2(n5535), .ZN(n5467)
         );
  OAI22_X1 U6611 ( .A1(n5465), .A2(n6036), .B1(n6030), .B2(n5613), .ZN(n5466)
         );
  AOI211_X1 U6612 ( .C1(n5468), .C2(REIP_REG_28__SCAN_IN), .A(n5467), .B(n5466), .ZN(n5471) );
  INV_X1 U6613 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6499) );
  NAND2_X1 U6614 ( .A1(n5469), .A2(n6499), .ZN(n5470) );
  OAI211_X1 U6615 ( .C1(n5568), .C2(n5985), .A(n5471), .B(n5470), .ZN(U2799)
         );
  AND2_X1 U6616 ( .A1(n5555), .A2(n5472), .ZN(n5486) );
  OAI21_X1 U6617 ( .B1(n5486), .B2(n5474), .A(n5473), .ZN(n5571) );
  INV_X1 U6618 ( .A(n5571), .ZN(n5623) );
  NOR3_X1 U6619 ( .A1(n5508), .A2(REIP_REG_27__SCAN_IN), .A3(n5475), .ZN(n5484) );
  INV_X1 U6620 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6497) );
  INV_X1 U6621 ( .A(n5476), .ZN(n5621) );
  NOR2_X1 U6622 ( .A1(n6030), .A2(n5621), .ZN(n5481) );
  AND2_X1 U6623 ( .A1(n5489), .A2(n5477), .ZN(n5479) );
  OR2_X1 U6624 ( .A1(n5479), .A2(n5478), .ZN(n5725) );
  INV_X1 U6625 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5536) );
  OAI22_X1 U6626 ( .A1(n5725), .A2(n6024), .B1(n6005), .B2(n5536), .ZN(n5480)
         );
  AOI211_X1 U6627 ( .C1(n6008), .C2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5481), 
        .B(n5480), .ZN(n5482) );
  OAI21_X1 U6628 ( .B1(n5495), .B2(n6497), .A(n5482), .ZN(n5483) );
  AOI211_X1 U6629 ( .C1(n5623), .C2(n3979), .A(n5484), .B(n5483), .ZN(n5485)
         );
  INV_X1 U6630 ( .A(n5485), .ZN(U2800) );
  AOI21_X1 U6631 ( .B1(n5488), .B2(n5487), .A(n5486), .ZN(n5632) );
  INV_X1 U6632 ( .A(n5632), .ZN(n5574) );
  INV_X1 U6633 ( .A(n5489), .ZN(n5490) );
  AOI21_X1 U6634 ( .B1(n5492), .B2(n5491), .A(n5490), .ZN(n5734) );
  AOI22_X1 U6635 ( .A1(n5734), .A2(n6033), .B1(n6032), .B2(EBX_REG_26__SCAN_IN), .ZN(n5493) );
  OAI21_X1 U6636 ( .B1(n5630), .B2(n6030), .A(n5493), .ZN(n5494) );
  AOI21_X1 U6637 ( .B1(PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n6008), .A(n5494), 
        .ZN(n5499) );
  INV_X1 U6638 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6490) );
  NOR3_X1 U6639 ( .A1(n5508), .A2(n6490), .A3(n6492), .ZN(n5497) );
  INV_X1 U6640 ( .A(n5495), .ZN(n5496) );
  OAI21_X1 U6641 ( .B1(n5497), .B2(REIP_REG_26__SCAN_IN), .A(n5496), .ZN(n5498) );
  OAI211_X1 U6642 ( .C1(n5574), .C2(n5985), .A(n5499), .B(n5498), .ZN(U2801)
         );
  NAND2_X1 U6643 ( .A1(n5538), .A2(n3979), .ZN(n5507) );
  INV_X1 U6644 ( .A(n5539), .ZN(n5500) );
  AOI22_X1 U6645 ( .A1(n5500), .A2(n6033), .B1(EBX_REG_24__SCAN_IN), .B2(n6032), .ZN(n5501) );
  OAI21_X1 U6646 ( .B1(n6036), .B2(n5502), .A(n5501), .ZN(n5504) );
  NOR2_X1 U6647 ( .A1(n5850), .A2(n6490), .ZN(n5503) );
  AOI211_X1 U6648 ( .C1(n6044), .C2(n5505), .A(n5504), .B(n5503), .ZN(n5506)
         );
  OAI211_X1 U6649 ( .C1(REIP_REG_24__SCAN_IN), .C2(n5508), .A(n5507), .B(n5506), .ZN(U2803) );
  INV_X1 U6650 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6487) );
  INV_X1 U6651 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6484) );
  INV_X1 U6652 ( .A(n5847), .ZN(n5865) );
  NOR2_X1 U6653 ( .A1(n6487), .A2(n6484), .ZN(n5846) );
  AOI211_X1 U6654 ( .C1(n6487), .C2(n6484), .A(n5865), .B(n5846), .ZN(n5509)
         );
  INV_X1 U6655 ( .A(n5509), .ZN(n5521) );
  NAND2_X1 U6656 ( .A1(n6015), .A2(n5510), .ZN(n5873) );
  NAND2_X1 U6657 ( .A1(n5547), .A2(n5511), .ZN(n5512) );
  NAND2_X1 U6658 ( .A1(n5513), .A2(n5512), .ZN(n5753) );
  OAI22_X1 U6659 ( .A1(n5753), .A2(n6024), .B1(n3094), .B2(n6005), .ZN(n5514)
         );
  AOI21_X1 U6660 ( .B1(n6008), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n5514), 
        .ZN(n5518) );
  INV_X1 U6661 ( .A(n5515), .ZN(n5516) );
  NAND2_X1 U6662 ( .A1(n6044), .A2(n5516), .ZN(n5517) );
  OAI211_X1 U6663 ( .C1(n5873), .C2(n6487), .A(n5518), .B(n5517), .ZN(n5519)
         );
  INV_X1 U6664 ( .A(n5519), .ZN(n5520) );
  OAI211_X1 U6665 ( .C1(n5582), .C2(n5985), .A(n5521), .B(n5520), .ZN(U2805)
         );
  NOR2_X1 U6666 ( .A1(n5524), .A2(n5523), .ZN(n5950) );
  OAI21_X1 U6667 ( .B1(n6036), .B2(n5666), .A(n4889), .ZN(n5527) );
  OAI22_X1 U6668 ( .A1(REIP_REG_19__SCAN_IN), .A2(n5866), .B1(n5525), .B2(
        n6005), .ZN(n5526) );
  AOI211_X1 U6669 ( .C1(REIP_REG_19__SCAN_IN), .C2(n5950), .A(n5527), .B(n5526), .ZN(n5534) );
  INV_X1 U6670 ( .A(n5776), .ZN(n5531) );
  NOR2_X1 U6671 ( .A1(n5530), .A2(n5528), .ZN(n5529) );
  AOI21_X1 U6672 ( .B1(n5531), .B2(n5530), .A(n5529), .ZN(n5557) );
  XNOR2_X1 U6673 ( .A(n5559), .B(n5532), .ZN(n5789) );
  INV_X1 U6674 ( .A(n5789), .ZN(n5550) );
  AOI22_X1 U6675 ( .A1(n5670), .A2(n6044), .B1(n6033), .B2(n5550), .ZN(n5533)
         );
  OAI211_X1 U6676 ( .C1(n5667), .C2(n5985), .A(n5534), .B(n5533), .ZN(U2808)
         );
  OAI222_X1 U6677 ( .A1(n6056), .A2(n5568), .B1(n5535), .B2(n6065), .C1(n5715), 
        .C2(n6055), .ZN(U2831) );
  OAI222_X1 U6678 ( .A1(n6056), .A2(n5571), .B1(n5536), .B2(n6065), .C1(n5725), 
        .C2(n6055), .ZN(U2832) );
  AOI22_X1 U6679 ( .A1(n5734), .A2(n6060), .B1(EBX_REG_26__SCAN_IN), .B2(n5549), .ZN(n5537) );
  OAI21_X1 U6680 ( .B1(n5574), .B2(n6056), .A(n5537), .ZN(U2833) );
  INV_X1 U6681 ( .A(n5538), .ZN(n5577) );
  INV_X1 U6682 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5540) );
  OAI222_X1 U6683 ( .A1(n6056), .A2(n5577), .B1(n6065), .B2(n5540), .C1(n5539), 
        .C2(n6055), .ZN(U2835) );
  AOI22_X1 U6684 ( .A1(n6060), .A2(n5848), .B1(EBX_REG_23__SCAN_IN), .B2(n5549), .ZN(n5541) );
  OAI21_X1 U6685 ( .B1(n5845), .B2(n6056), .A(n5541), .ZN(U2836) );
  OAI222_X1 U6686 ( .A1(n6056), .A2(n5582), .B1(n6065), .B2(n3094), .C1(n5753), 
        .C2(n6055), .ZN(U2837) );
  AOI21_X1 U6687 ( .B1(n5543), .B2(n5653), .A(n5542), .ZN(n5862) );
  INV_X1 U6688 ( .A(n5862), .ZN(n5585) );
  INV_X1 U6689 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5548) );
  OR2_X1 U6690 ( .A1(n5545), .A2(n5544), .ZN(n5546) );
  NAND2_X1 U6691 ( .A1(n5547), .A2(n5546), .ZN(n5860) );
  OAI222_X1 U6692 ( .A1(n5585), .A2(n6056), .B1(n5548), .B2(n6065), .C1(n6055), 
        .C2(n5860), .ZN(U2838) );
  AOI22_X1 U6693 ( .A1(n6060), .A2(n5550), .B1(EBX_REG_19__SCAN_IN), .B2(n5549), .ZN(n5551) );
  OAI21_X1 U6694 ( .B1(n5667), .B2(n6056), .A(n5551), .ZN(U2840) );
  NOR2_X1 U6695 ( .A1(n5553), .A2(n5552), .ZN(n5554) );
  OR2_X1 U6696 ( .A1(n5555), .A2(n5554), .ZN(n5676) );
  NAND2_X1 U6697 ( .A1(n5557), .A2(n5556), .ZN(n5558) );
  AND2_X1 U6698 ( .A1(n5559), .A2(n5558), .ZN(n5948) );
  INV_X1 U6699 ( .A(n5948), .ZN(n5560) );
  OAI222_X1 U6700 ( .A1(n5676), .A2(n6056), .B1(n5561), .B2(n6065), .C1(n6055), 
        .C2(n5560), .ZN(U2841) );
  NAND3_X1 U6701 ( .A1(n5598), .A2(n5563), .A3(n5562), .ZN(n5565) );
  AOI22_X1 U6702 ( .A1(n6073), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6076), .ZN(n5564) );
  NAND2_X1 U6703 ( .A1(n5565), .A2(n5564), .ZN(U2860) );
  AOI22_X1 U6704 ( .A1(n6073), .A2(DATAI_28_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n6076), .ZN(n5567) );
  NAND2_X1 U6705 ( .A1(n6077), .A2(DATAI_12_), .ZN(n5566) );
  OAI211_X1 U6706 ( .C1(n5568), .C2(n5877), .A(n5567), .B(n5566), .ZN(U2863)
         );
  AOI22_X1 U6707 ( .A1(n6073), .A2(DATAI_27_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n6076), .ZN(n5570) );
  NAND2_X1 U6708 ( .A1(n6077), .A2(DATAI_11_), .ZN(n5569) );
  OAI211_X1 U6709 ( .C1(n5571), .C2(n5877), .A(n5570), .B(n5569), .ZN(U2864)
         );
  AOI22_X1 U6710 ( .A1(n6073), .A2(DATAI_26_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n6076), .ZN(n5573) );
  NAND2_X1 U6711 ( .A1(n6077), .A2(DATAI_10_), .ZN(n5572) );
  OAI211_X1 U6712 ( .C1(n5574), .C2(n5877), .A(n5573), .B(n5572), .ZN(U2865)
         );
  AOI22_X1 U6713 ( .A1(n6073), .A2(DATAI_24_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n6076), .ZN(n5576) );
  NAND2_X1 U6714 ( .A1(n6077), .A2(DATAI_8_), .ZN(n5575) );
  OAI211_X1 U6715 ( .C1(n5577), .C2(n5877), .A(n5576), .B(n5575), .ZN(U2867)
         );
  AOI22_X1 U6716 ( .A1(n6073), .A2(DATAI_23_), .B1(EAX_REG_23__SCAN_IN), .B2(
        n6076), .ZN(n5579) );
  NAND2_X1 U6717 ( .A1(n6077), .A2(DATAI_7_), .ZN(n5578) );
  OAI211_X1 U6718 ( .C1(n5845), .C2(n5877), .A(n5579), .B(n5578), .ZN(U2868)
         );
  AOI22_X1 U6719 ( .A1(n6073), .A2(DATAI_22_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n6076), .ZN(n5581) );
  NAND2_X1 U6720 ( .A1(n6077), .A2(DATAI_6_), .ZN(n5580) );
  OAI211_X1 U6721 ( .C1(n5582), .C2(n5877), .A(n5581), .B(n5580), .ZN(U2869)
         );
  AOI22_X1 U6722 ( .A1(n6073), .A2(DATAI_21_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n6076), .ZN(n5584) );
  NAND2_X1 U6723 ( .A1(n6077), .A2(DATAI_5_), .ZN(n5583) );
  OAI211_X1 U6724 ( .C1(n5585), .C2(n5877), .A(n5584), .B(n5583), .ZN(U2870)
         );
  AOI22_X1 U6725 ( .A1(n6073), .A2(DATAI_19_), .B1(EAX_REG_19__SCAN_IN), .B2(
        n6076), .ZN(n5587) );
  NAND2_X1 U6726 ( .A1(n6077), .A2(DATAI_3_), .ZN(n5586) );
  OAI211_X1 U6727 ( .C1(n5667), .C2(n5877), .A(n5587), .B(n5586), .ZN(U2872)
         );
  NAND2_X1 U6728 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5593) );
  INV_X1 U6729 ( .A(n5588), .ZN(n5634) );
  NAND4_X1 U6730 ( .A1(n5634), .A2(n5591), .A3(n5590), .A4(n5589), .ZN(n5592)
         );
  OAI21_X1 U6731 ( .B1(n5601), .B2(n5593), .A(n5592), .ZN(n5594) );
  XNOR2_X1 U6732 ( .A(n5594), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5705)
         );
  NAND2_X1 U6733 ( .A1(n6018), .A2(REIP_REG_31__SCAN_IN), .ZN(n5700) );
  NAND2_X1 U6734 ( .A1(n6171), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5595)
         );
  OAI211_X1 U6735 ( .C1(n6182), .C2(n5596), .A(n5700), .B(n5595), .ZN(n5597)
         );
  AOI21_X1 U6736 ( .B1(n5598), .B2(n6176), .A(n5597), .ZN(n5599) );
  OAI21_X1 U6737 ( .B1(n5705), .B2(n6166), .A(n5599), .ZN(U2955) );
  NAND2_X1 U6738 ( .A1(n5601), .A2(n5600), .ZN(n5602) );
  XNOR2_X1 U6739 ( .A(n5602), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5714)
         );
  AND2_X1 U6740 ( .A1(n6018), .A2(REIP_REG_29__SCAN_IN), .ZN(n5707) );
  AOI21_X1 U6741 ( .B1(n6171), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5707), 
        .ZN(n5603) );
  OAI21_X1 U6742 ( .B1(n6182), .B2(n5604), .A(n5603), .ZN(n5605) );
  AOI21_X1 U6743 ( .B1(n5606), .B2(n6176), .A(n5605), .ZN(n5607) );
  OAI21_X1 U6744 ( .B1(n5714), .B2(n6166), .A(n5607), .ZN(U2957) );
  NOR3_X1 U6745 ( .A1(n5627), .A2(n5673), .A3(n5716), .ZN(n5609) );
  OR2_X1 U6746 ( .A1(n5626), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5608)
         );
  NOR2_X1 U6747 ( .A1(n5635), .A2(n5608), .ZN(n5617) );
  OAI22_X1 U6748 ( .A1(n5609), .A2(n5617), .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n5716), .ZN(n5611) );
  XNOR2_X1 U6749 ( .A(n5611), .B(n5610), .ZN(n5724) );
  AND2_X1 U6750 ( .A1(n6189), .A2(REIP_REG_28__SCAN_IN), .ZN(n5718) );
  AOI21_X1 U6751 ( .B1(n6171), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5718), 
        .ZN(n5612) );
  OAI21_X1 U6752 ( .B1(n6182), .B2(n5613), .A(n5612), .ZN(n5614) );
  AOI21_X1 U6753 ( .B1(n5615), .B2(n6176), .A(n5614), .ZN(n5616) );
  OAI21_X1 U6754 ( .B1(n6166), .B2(n5724), .A(n5616), .ZN(U2958) );
  NOR2_X1 U6755 ( .A1(n5618), .A2(n5617), .ZN(n5619) );
  XNOR2_X1 U6756 ( .A(n5619), .B(n5716), .ZN(n5732) );
  AND2_X1 U6757 ( .A1(n6189), .A2(REIP_REG_27__SCAN_IN), .ZN(n5727) );
  AOI21_X1 U6758 ( .B1(n6171), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5727), 
        .ZN(n5620) );
  OAI21_X1 U6759 ( .B1(n6182), .B2(n5621), .A(n5620), .ZN(n5622) );
  AOI21_X1 U6760 ( .B1(n5623), .B2(n6176), .A(n5622), .ZN(n5624) );
  OAI21_X1 U6761 ( .B1(n5732), .B2(n6166), .A(n5624), .ZN(U2959) );
  NAND2_X1 U6762 ( .A1(n5626), .A2(n5625), .ZN(n5628) );
  XOR2_X1 U6763 ( .A(n5628), .B(n5627), .Z(n5739) );
  AND2_X1 U6764 ( .A1(n6189), .A2(REIP_REG_26__SCAN_IN), .ZN(n5733) );
  AOI21_X1 U6765 ( .B1(n6171), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5733), 
        .ZN(n5629) );
  OAI21_X1 U6766 ( .B1(n6182), .B2(n5630), .A(n5629), .ZN(n5631) );
  AOI21_X1 U6767 ( .B1(n5632), .B2(n6176), .A(n5631), .ZN(n5633) );
  OAI21_X1 U6768 ( .B1(n5739), .B2(n6166), .A(n5633), .ZN(U2960) );
  AOI21_X1 U6769 ( .B1(n5636), .B2(n5635), .A(n5634), .ZN(n5748) );
  INV_X1 U6770 ( .A(n5637), .ZN(n5639) );
  AND2_X1 U6771 ( .A1(n6189), .A2(REIP_REG_25__SCAN_IN), .ZN(n5741) );
  AOI21_X1 U6772 ( .B1(n6171), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n5741), 
        .ZN(n5638) );
  OAI21_X1 U6773 ( .B1(n6182), .B2(n5639), .A(n5638), .ZN(n5640) );
  AOI21_X1 U6774 ( .B1(n5641), .B2(n6176), .A(n5640), .ZN(n5642) );
  OAI21_X1 U6775 ( .B1(n5748), .B2(n6166), .A(n5642), .ZN(U2961) );
  AOI21_X1 U6776 ( .B1(n5645), .B2(n5644), .A(n5643), .ZN(n5765) );
  INV_X1 U6777 ( .A(n5859), .ZN(n5647) );
  NAND2_X1 U6778 ( .A1(n6171), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5646)
         );
  NAND2_X1 U6779 ( .A1(n6018), .A2(REIP_REG_21__SCAN_IN), .ZN(n5760) );
  OAI211_X1 U6780 ( .C1(n6182), .C2(n5647), .A(n5646), .B(n5760), .ZN(n5648)
         );
  AOI21_X1 U6781 ( .B1(n5862), .B2(n6176), .A(n5648), .ZN(n5649) );
  OAI21_X1 U6782 ( .B1(n5765), .B2(n6166), .A(n5649), .ZN(U2965) );
  OAI21_X1 U6783 ( .B1(n5652), .B2(n5651), .A(n5650), .ZN(n5787) );
  INV_X1 U6784 ( .A(n5653), .ZN(n5654) );
  NAND2_X1 U6785 ( .A1(n6018), .A2(REIP_REG_20__SCAN_IN), .ZN(n5780) );
  NAND2_X1 U6786 ( .A1(n6171), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5657)
         );
  OAI211_X1 U6787 ( .C1(n5869), .C2(n6182), .A(n5780), .B(n5657), .ZN(n5658)
         );
  AOI21_X1 U6788 ( .B1(n5878), .B2(n6176), .A(n5658), .ZN(n5659) );
  OAI21_X1 U6789 ( .B1(n5787), .B2(n6166), .A(n5659), .ZN(U2966) );
  AND2_X1 U6790 ( .A1(n5661), .A2(n5660), .ZN(n5664) );
  OAI21_X1 U6791 ( .B1(n5664), .B2(n5663), .A(n5662), .ZN(n5665) );
  XNOR2_X1 U6792 ( .A(n5665), .B(n4079), .ZN(n5795) );
  NAND2_X1 U6793 ( .A1(n6189), .A2(REIP_REG_19__SCAN_IN), .ZN(n5788) );
  OAI21_X1 U6794 ( .B1(n5684), .B2(n5666), .A(n5788), .ZN(n5669) );
  NOR2_X1 U6795 ( .A1(n5667), .A2(n6164), .ZN(n5668) );
  OAI21_X1 U6796 ( .B1(n6166), .B2(n5795), .A(n5671), .ZN(U2967) );
  INV_X1 U6797 ( .A(n5672), .ZN(n5682) );
  NAND3_X1 U6798 ( .A1(n5682), .A2(n5673), .A3(n5898), .ZN(n5804) );
  NOR3_X1 U6799 ( .A1(n5682), .A2(n5673), .A3(n5898), .ZN(n5806) );
  NAND2_X1 U6800 ( .A1(n5806), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5674) );
  OAI21_X1 U6801 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5804), .A(n5674), 
        .ZN(n5675) );
  XNOR2_X1 U6802 ( .A(n5675), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5803)
         );
  AND2_X1 U6803 ( .A1(n6189), .A2(REIP_REG_18__SCAN_IN), .ZN(n5798) );
  AOI21_X1 U6804 ( .B1(n6171), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n5798), 
        .ZN(n5677) );
  OAI21_X1 U6805 ( .B1(n5678), .B2(n6182), .A(n5677), .ZN(n5679) );
  AOI21_X1 U6806 ( .B1(n6066), .B2(n6176), .A(n5679), .ZN(n5680) );
  OAI21_X1 U6807 ( .B1(n5803), .B2(n6166), .A(n5680), .ZN(U2968) );
  XNOR2_X1 U6808 ( .A(n4079), .B(n5898), .ZN(n5681) );
  XNOR2_X1 U6809 ( .A(n5682), .B(n5681), .ZN(n5892) );
  INV_X1 U6810 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5683) );
  OAI22_X1 U6811 ( .A1(n5684), .A2(n5683), .B1(n4889), .B2(n6476), .ZN(n5686)
         );
  NOR2_X1 U6812 ( .A1(n6072), .A2(n6164), .ZN(n5685) );
  AOI211_X1 U6813 ( .C1(n5883), .C2(n5687), .A(n5686), .B(n5685), .ZN(n5688)
         );
  OAI21_X1 U6814 ( .B1(n6166), .B2(n5892), .A(n5688), .ZN(U2970) );
  INV_X1 U6815 ( .A(n6042), .ZN(n5689) );
  NAND2_X1 U6816 ( .A1(n5689), .A2(n6176), .ZN(n5696) );
  AOI22_X1 U6817 ( .A1(n6171), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .B1(n6018), 
        .B2(REIP_REG_3__SCAN_IN), .ZN(n5695) );
  AND2_X1 U6818 ( .A1(n5691), .A2(n5690), .ZN(n6243) );
  INV_X1 U6819 ( .A(n6243), .ZN(n5692) );
  NAND3_X1 U6820 ( .A1(n5692), .A2(n6178), .A3(n6248), .ZN(n5694) );
  NAND2_X1 U6821 ( .A1(n5883), .A2(n6045), .ZN(n5693) );
  NAND4_X1 U6822 ( .A1(n5696), .A2(n5695), .A3(n5694), .A4(n5693), .ZN(U2983)
         );
  OAI21_X1 U6823 ( .B1(n6203), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5697), 
        .ZN(n5703) );
  NAND4_X1 U6824 ( .A1(n5706), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_30__SCAN_IN), .A4(n5698), .ZN(n5699) );
  OAI211_X1 U6825 ( .C1(n5701), .C2(n6246), .A(n5700), .B(n5699), .ZN(n5702)
         );
  AOI21_X1 U6826 ( .B1(n5703), .B2(INSTADDRPOINTER_REG_31__SCAN_IN), .A(n5702), 
        .ZN(n5704) );
  OAI21_X1 U6827 ( .B1(n5705), .B2(n6242), .A(n5704), .ZN(U2987) );
  INV_X1 U6828 ( .A(n5706), .ZN(n5710) );
  AOI21_X1 U6829 ( .B1(n5708), .B2(n6258), .A(n5707), .ZN(n5709) );
  OAI21_X1 U6830 ( .B1(n5710), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5709), 
        .ZN(n5711) );
  AOI21_X1 U6831 ( .B1(n5712), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5711), 
        .ZN(n5713) );
  OAI21_X1 U6832 ( .B1(n5714), .B2(n6242), .A(n5713), .ZN(U2989) );
  INV_X1 U6833 ( .A(n5715), .ZN(n5719) );
  NOR3_X1 U6834 ( .A1(n5721), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .A3(n5716), 
        .ZN(n5717) );
  AOI211_X1 U6835 ( .C1(n6258), .C2(n5719), .A(n5718), .B(n5717), .ZN(n5723)
         );
  INV_X1 U6836 ( .A(n5720), .ZN(n5729) );
  NOR2_X1 U6837 ( .A1(n5721), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5726)
         );
  OAI21_X1 U6838 ( .B1(n5729), .B2(n5726), .A(INSTADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n5722) );
  OAI211_X1 U6839 ( .C1(n5724), .C2(n6242), .A(n5723), .B(n5722), .ZN(U2990)
         );
  INV_X1 U6840 ( .A(n5725), .ZN(n5728) );
  AOI211_X1 U6841 ( .C1(n6258), .C2(n5728), .A(n5727), .B(n5726), .ZN(n5731)
         );
  NAND2_X1 U6842 ( .A1(n5729), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5730) );
  OAI211_X1 U6843 ( .C1(n5732), .C2(n6242), .A(n5731), .B(n5730), .ZN(U2991)
         );
  XNOR2_X1 U6844 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .B(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5736) );
  AOI21_X1 U6845 ( .B1(n5734), .B2(n6258), .A(n5733), .ZN(n5735) );
  OAI21_X1 U6846 ( .B1(n5744), .B2(n5736), .A(n5735), .ZN(n5737) );
  AOI21_X1 U6847 ( .B1(n5746), .B2(INSTADDRPOINTER_REG_26__SCAN_IN), .A(n5737), 
        .ZN(n5738) );
  OAI21_X1 U6848 ( .B1(n5739), .B2(n6242), .A(n5738), .ZN(U2992) );
  INV_X1 U6849 ( .A(n5740), .ZN(n5742) );
  AOI21_X1 U6850 ( .B1(n5742), .B2(n6258), .A(n5741), .ZN(n5743) );
  OAI21_X1 U6851 ( .B1(n5744), .B2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5743), 
        .ZN(n5745) );
  AOI21_X1 U6852 ( .B1(n5746), .B2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5745), 
        .ZN(n5747) );
  OAI21_X1 U6853 ( .B1(n5748), .B2(n6242), .A(n5747), .ZN(U2993) );
  INV_X1 U6854 ( .A(n5759), .ZN(n5751) );
  NOR3_X1 U6855 ( .A1(n5751), .A2(n5750), .A3(n5749), .ZN(n5755) );
  OAI21_X1 U6856 ( .B1(n6246), .B2(n5753), .A(n5752), .ZN(n5754) );
  AOI211_X1 U6857 ( .C1(n5763), .C2(INSTADDRPOINTER_REG_22__SCAN_IN), .A(n5755), .B(n5754), .ZN(n5756) );
  OAI21_X1 U6858 ( .B1(n5757), .B2(n6242), .A(n5756), .ZN(U2996) );
  NAND2_X1 U6859 ( .A1(n5759), .A2(n5758), .ZN(n5761) );
  OAI211_X1 U6860 ( .C1(n6246), .C2(n5860), .A(n5761), .B(n5760), .ZN(n5762)
         );
  AOI21_X1 U6861 ( .B1(n5763), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5762), 
        .ZN(n5764) );
  OAI21_X1 U6862 ( .B1(n5765), .B2(n6242), .A(n5764), .ZN(U2997) );
  INV_X1 U6863 ( .A(n5766), .ZN(n5770) );
  OAI21_X1 U6864 ( .B1(n6629), .B2(n5767), .A(n6260), .ZN(n5768) );
  OAI211_X1 U6865 ( .C1(n5771), .C2(n5770), .A(n5769), .B(n5768), .ZN(n5812)
         );
  AOI21_X1 U6866 ( .B1(n6254), .B2(n6629), .A(n5812), .ZN(n5796) );
  OAI21_X1 U6867 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n6203), .A(n5796), 
        .ZN(n5793) );
  NAND2_X1 U6868 ( .A1(n5773), .A2(n5772), .ZN(n5777) );
  NAND2_X1 U6869 ( .A1(n5777), .A2(n5774), .ZN(n5775) );
  OAI21_X1 U6870 ( .B1(n5777), .B2(n5776), .A(n5775), .ZN(n5779) );
  XNOR2_X1 U6871 ( .A(n5779), .B(n5778), .ZN(n5868) );
  OAI21_X1 U6872 ( .B1(n6246), .B2(n5868), .A(n5780), .ZN(n5785) );
  NAND2_X1 U6873 ( .A1(n6186), .A2(n5781), .ZN(n5809) );
  INV_X1 U6874 ( .A(n5809), .ZN(n5800) );
  NAND3_X1 U6875 ( .A1(n5800), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5790) );
  NOR3_X1 U6876 ( .A1(n5790), .A2(n5783), .A3(n5782), .ZN(n5784) );
  AOI211_X1 U6877 ( .C1(INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n5793), .A(n5785), .B(n5784), .ZN(n5786) );
  OAI21_X1 U6878 ( .B1(n5787), .B2(n6242), .A(n5786), .ZN(U2998) );
  OAI21_X1 U6879 ( .B1(n6246), .B2(n5789), .A(n5788), .ZN(n5792) );
  NOR2_X1 U6880 ( .A1(n5790), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5791)
         );
  AOI211_X1 U6881 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n5793), .A(n5792), .B(n5791), .ZN(n5794) );
  OAI21_X1 U6882 ( .B1(n5795), .B2(n6242), .A(n5794), .ZN(U2999) );
  NOR2_X1 U6883 ( .A1(n5796), .A2(n5799), .ZN(n5797) );
  AOI211_X1 U6884 ( .C1(n6258), .C2(n5948), .A(n5798), .B(n5797), .ZN(n5802)
         );
  NAND3_X1 U6885 ( .A1(n5800), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n5799), .ZN(n5801) );
  OAI211_X1 U6886 ( .C1(n5803), .C2(n6242), .A(n5802), .B(n5801), .ZN(U3000)
         );
  INV_X1 U6887 ( .A(n5804), .ZN(n5805) );
  NOR2_X1 U6888 ( .A1(n5806), .A2(n5805), .ZN(n5807) );
  XNOR2_X1 U6889 ( .A(n5807), .B(n6629), .ZN(n5886) );
  OAI22_X1 U6890 ( .A1(n6246), .A2(n5808), .B1(n4889), .B2(n6478), .ZN(n5811)
         );
  NOR2_X1 U6891 ( .A1(n5809), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5810)
         );
  AOI211_X1 U6892 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n5812), .A(n5811), .B(n5810), .ZN(n5813) );
  OAI21_X1 U6893 ( .B1(n5886), .B2(n6242), .A(n5813), .ZN(U3001) );
  NAND2_X1 U6894 ( .A1(n5814), .A2(n6263), .ZN(n5828) );
  NAND3_X1 U6895 ( .A1(n5820), .A2(n4090), .A3(n6186), .ZN(n5827) );
  OAI22_X1 U6896 ( .A1(n6246), .A2(n5815), .B1(n6470), .B2(n4889), .ZN(n5816)
         );
  INV_X1 U6897 ( .A(n5816), .ZN(n5826) );
  AOI21_X1 U6898 ( .B1(n6185), .B2(n5817), .A(n6183), .ZN(n5818) );
  OAI21_X1 U6899 ( .B1(n5820), .B2(n5819), .A(n5818), .ZN(n5914) );
  INV_X1 U6900 ( .A(n5821), .ZN(n5823) );
  AOI21_X1 U6901 ( .B1(n5823), .B2(n5822), .A(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n5824) );
  OAI21_X1 U6902 ( .B1(n5914), .B2(n5824), .A(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n5825) );
  NAND4_X1 U6903 ( .A1(n5828), .A2(n5827), .A3(n5826), .A4(n5825), .ZN(U3004)
         );
  OAI21_X1 U6904 ( .B1(n5830), .B2(STATEBS16_REG_SCAN_IN), .A(n5829), .ZN(
        n5832) );
  OAI22_X1 U6905 ( .A1(n5832), .A2(n5834), .B1(n5831), .B2(n5836), .ZN(n5833)
         );
  MUX2_X1 U6906 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5833), .S(n6268), 
        .Z(U3464) );
  XNOR2_X1 U6907 ( .A(n5835), .B(n5834), .ZN(n5839) );
  OAI22_X1 U6908 ( .A1(n5839), .A2(n5838), .B1(n5837), .B2(n5836), .ZN(n5840)
         );
  MUX2_X1 U6909 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5840), .S(n6268), 
        .Z(U3463) );
  OAI22_X1 U6910 ( .A1(n5842), .A2(n6547), .B1(n5841), .B2(n6550), .ZN(n5843)
         );
  MUX2_X1 U6911 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5843), .S(n6553), 
        .Z(U3456) );
  AND2_X1 U6912 ( .A1(n6115), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  INV_X1 U6913 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5856) );
  AOI22_X1 U6914 ( .A1(PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n6008), .B1(n5844), 
        .B2(n6044), .ZN(n5855) );
  INV_X1 U6915 ( .A(n5845), .ZN(n5853) );
  AOI21_X1 U6916 ( .B1(n5847), .B2(n5846), .A(REIP_REG_23__SCAN_IN), .ZN(n5851) );
  INV_X1 U6917 ( .A(n5848), .ZN(n5849) );
  OAI22_X1 U6918 ( .A1(n5851), .A2(n5850), .B1(n5849), .B2(n6024), .ZN(n5852)
         );
  AOI21_X1 U6919 ( .B1(n5853), .B2(n3979), .A(n5852), .ZN(n5854) );
  OAI211_X1 U6920 ( .C1(n5856), .C2(n6005), .A(n5855), .B(n5854), .ZN(U2804)
         );
  AOI22_X1 U6921 ( .A1(EBX_REG_21__SCAN_IN), .A2(n6032), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6008), .ZN(n5857) );
  OAI21_X1 U6922 ( .B1(n6484), .B2(n5873), .A(n5857), .ZN(n5858) );
  AOI21_X1 U6923 ( .B1(n5859), .B2(n6044), .A(n5858), .ZN(n5864) );
  INV_X1 U6924 ( .A(n5860), .ZN(n5861) );
  AOI22_X1 U6925 ( .A1(n5862), .A2(n3979), .B1(n6033), .B2(n5861), .ZN(n5863)
         );
  OAI211_X1 U6926 ( .C1(REIP_REG_21__SCAN_IN), .C2(n5865), .A(n5864), .B(n5863), .ZN(U2806) );
  INV_X1 U6927 ( .A(n5866), .ZN(n5867) );
  AOI21_X1 U6928 ( .B1(n5867), .B2(REIP_REG_19__SCAN_IN), .A(
        REIP_REG_20__SCAN_IN), .ZN(n5874) );
  INV_X1 U6929 ( .A(n5868), .ZN(n5875) );
  AOI22_X1 U6930 ( .A1(n5878), .A2(n3979), .B1(n6033), .B2(n5875), .ZN(n5872)
         );
  OAI22_X1 U6931 ( .A1(n3082), .A2(n6005), .B1(n5869), .B2(n6030), .ZN(n5870)
         );
  AOI21_X1 U6932 ( .B1(PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6008), .A(n5870), 
        .ZN(n5871) );
  OAI211_X1 U6933 ( .C1(n5874), .C2(n5873), .A(n5872), .B(n5871), .ZN(U2807)
         );
  AOI22_X1 U6934 ( .A1(n5878), .A2(n6061), .B1(n6060), .B2(n5875), .ZN(n5876)
         );
  OAI21_X1 U6935 ( .B1(n6065), .B2(n3082), .A(n5876), .ZN(U2839) );
  INV_X1 U6936 ( .A(n5877), .ZN(n6074) );
  AOI22_X1 U6937 ( .A1(n5878), .A2(n6074), .B1(n6073), .B2(DATAI_20_), .ZN(
        n5880) );
  AOI22_X1 U6938 ( .A1(n6077), .A2(DATAI_4_), .B1(n6076), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5879) );
  NAND2_X1 U6939 ( .A1(n5880), .A2(n5879), .ZN(U2871) );
  AOI22_X1 U6940 ( .A1(n6189), .A2(REIP_REG_17__SCAN_IN), .B1(n6171), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5885) );
  INV_X1 U6941 ( .A(n5881), .ZN(n6069) );
  AOI22_X1 U6942 ( .A1(n6069), .A2(n6176), .B1(n5883), .B2(n5882), .ZN(n5884)
         );
  OAI211_X1 U6943 ( .C1(n5886), .C2(n6166), .A(n5885), .B(n5884), .ZN(U2969)
         );
  AOI22_X1 U6944 ( .A1(n6189), .A2(REIP_REG_13__SCAN_IN), .B1(n6171), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5890) );
  XNOR2_X1 U6945 ( .A(n5888), .B(n5887), .ZN(n5915) );
  AOI22_X1 U6946 ( .A1(n5915), .A2(n6178), .B1(n6176), .B2(n6051), .ZN(n5889)
         );
  OAI211_X1 U6947 ( .C1(n6182), .C2(n5969), .A(n5890), .B(n5889), .ZN(U2973)
         );
  AOI21_X1 U6948 ( .B1(n5901), .B2(n6201), .A(n6183), .ZN(n5907) );
  INV_X1 U6949 ( .A(n6186), .ZN(n5919) );
  AOI211_X1 U6950 ( .C1(n5906), .C2(n5898), .A(n5919), .B(n5901), .ZN(n5895)
         );
  OAI22_X1 U6951 ( .A1(n5892), .A2(n6242), .B1(n6246), .B2(n5891), .ZN(n5893)
         );
  AOI21_X1 U6952 ( .B1(n5895), .B2(n5894), .A(n5893), .ZN(n5897) );
  NAND2_X1 U6953 ( .A1(n6189), .A2(REIP_REG_16__SCAN_IN), .ZN(n5896) );
  OAI211_X1 U6954 ( .C1(n5907), .C2(n5898), .A(n5897), .B(n5896), .ZN(U3002)
         );
  AOI21_X1 U6955 ( .B1(n6258), .B2(n5900), .A(n5899), .ZN(n5905) );
  NOR2_X1 U6956 ( .A1(n5919), .A2(n5901), .ZN(n5902) );
  AOI22_X1 U6957 ( .A1(n5903), .A2(n6263), .B1(n5902), .B2(n5906), .ZN(n5904)
         );
  OAI211_X1 U6958 ( .C1(n5907), .C2(n5906), .A(n5905), .B(n5904), .ZN(U3003)
         );
  OR2_X1 U6959 ( .A1(n6185), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5918)
         );
  NAND2_X1 U6960 ( .A1(n5909), .A2(n5908), .ZN(n5912) );
  INV_X1 U6961 ( .A(n5910), .ZN(n5911) );
  NAND2_X1 U6962 ( .A1(n5912), .A2(n5911), .ZN(n6049) );
  INV_X1 U6963 ( .A(n6049), .ZN(n5913) );
  AOI22_X1 U6964 ( .A1(n6258), .A2(n5913), .B1(n6018), .B2(
        REIP_REG_13__SCAN_IN), .ZN(n5917) );
  AOI22_X1 U6965 ( .A1(n5915), .A2(n6263), .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5914), .ZN(n5916) );
  OAI211_X1 U6966 ( .C1(n5919), .C2(n5918), .A(n5917), .B(n5916), .ZN(U3005)
         );
  OR4_X1 U6967 ( .A1(n5922), .A2(n5921), .A3(n5920), .A4(n6547), .ZN(n5923) );
  OAI21_X1 U6968 ( .B1(n6553), .B2(n5924), .A(n5923), .ZN(U3455) );
  INV_X1 U6969 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6450) );
  AOI21_X1 U6970 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6450), .A(n6442), .ZN(n5930) );
  INV_X1 U6971 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5925) );
  AND2_X1 U6972 ( .A1(n6442), .A2(STATE_REG_1__SCAN_IN), .ZN(n6471) );
  AOI21_X1 U6973 ( .B1(n5930), .B2(n5925), .A(n6471), .ZN(U2789) );
  OAI21_X1 U6974 ( .B1(n5926), .B2(n6424), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5927) );
  OAI21_X1 U6975 ( .B1(n5928), .B2(n6529), .A(n5927), .ZN(U2790) );
  INV_X2 U6976 ( .A(n6471), .ZN(n6540) );
  NOR2_X1 U6977 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n5931) );
  OAI21_X1 U6978 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5931), .A(n6540), .ZN(n5929)
         );
  OAI21_X1 U6979 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6540), .A(n5929), .ZN(
        U2791) );
  NOR2_X1 U6980 ( .A1(n6471), .A2(n5930), .ZN(n6509) );
  OAI21_X1 U6981 ( .B1(BS16_N), .B2(n5931), .A(n6509), .ZN(n6507) );
  OAI21_X1 U6982 ( .B1(n6509), .B2(n6527), .A(n6507), .ZN(U2792) );
  AOI21_X1 U6983 ( .B1(n5932), .B2(FLUSH_REG_SCAN_IN), .A(n6178), .ZN(n5933)
         );
  INV_X1 U6984 ( .A(n5933), .ZN(U2793) );
  NOR2_X1 U6985 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(
        DATAWIDTH_REG_30__SCAN_IN), .ZN(n6686) );
  AOI211_X1 U6986 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_14__SCAN_IN), .B(
        DATAWIDTH_REG_2__SCAN_IN), .ZN(n5934) );
  INV_X1 U6987 ( .A(DATAWIDTH_REG_17__SCAN_IN), .ZN(n6660) );
  INV_X1 U6988 ( .A(DATAWIDTH_REG_5__SCAN_IN), .ZN(n6646) );
  NAND4_X1 U6989 ( .A1(n6686), .A2(n5934), .A3(n6660), .A4(n6646), .ZN(n5942)
         );
  OR4_X1 U6990 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(DATAWIDTH_REG_9__SCAN_IN), 
        .A3(DATAWIDTH_REG_10__SCAN_IN), .A4(DATAWIDTH_REG_11__SCAN_IN), .ZN(
        n5941) );
  OR4_X1 U6991 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), 
        .A3(DATAWIDTH_REG_6__SCAN_IN), .A4(DATAWIDTH_REG_7__SCAN_IN), .ZN(
        n5940) );
  NOR4_X1 U6992 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(
        DATAWIDTH_REG_19__SCAN_IN), .A3(DATAWIDTH_REG_20__SCAN_IN), .A4(
        DATAWIDTH_REG_22__SCAN_IN), .ZN(n5938) );
  NOR4_X1 U6993 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(
        DATAWIDTH_REG_12__SCAN_IN), .A3(DATAWIDTH_REG_13__SCAN_IN), .A4(
        DATAWIDTH_REG_16__SCAN_IN), .ZN(n5937) );
  NOR4_X1 U6994 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(
        DATAWIDTH_REG_27__SCAN_IN), .A3(DATAWIDTH_REG_28__SCAN_IN), .A4(
        DATAWIDTH_REG_29__SCAN_IN), .ZN(n5936) );
  NOR4_X1 U6995 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(
        DATAWIDTH_REG_24__SCAN_IN), .A3(DATAWIDTH_REG_25__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5935) );
  NAND4_X1 U6996 ( .A1(n5938), .A2(n5937), .A3(n5936), .A4(n5935), .ZN(n5939)
         );
  INV_X1 U6997 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n5944) );
  NOR3_X1 U6998 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5945) );
  OAI21_X1 U6999 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5945), .A(n6516), .ZN(n5943)
         );
  OAI21_X1 U7000 ( .B1(n6516), .B2(n5944), .A(n5943), .ZN(U2794) );
  INV_X1 U7001 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6508) );
  AOI21_X1 U7002 ( .B1(n6513), .B2(n6508), .A(n5945), .ZN(n5947) );
  INV_X1 U7003 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n5946) );
  INV_X1 U7004 ( .A(n6516), .ZN(n6519) );
  AOI22_X1 U7005 ( .A1(n6516), .A2(n5947), .B1(n5946), .B2(n6519), .ZN(U2795)
         );
  AOI22_X1 U7006 ( .A1(EBX_REG_18__SCAN_IN), .A2(n6032), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6008), .ZN(n5954) );
  AOI222_X1 U7007 ( .A1(n6066), .A2(n3979), .B1(n5949), .B2(n6044), .C1(n6033), 
        .C2(n5948), .ZN(n5953) );
  OAI21_X1 U7008 ( .B1(REIP_REG_18__SCAN_IN), .B2(n5951), .A(n5950), .ZN(n5952) );
  NAND4_X1 U7009 ( .A1(n5954), .A2(n5953), .A3(n4889), .A4(n5952), .ZN(U2809)
         );
  NAND2_X1 U7010 ( .A1(n5956), .A2(n6000), .ZN(n5979) );
  AOI211_X1 U7011 ( .C1(n6472), .C2(n6469), .A(n5955), .B(n5979), .ZN(n5966)
         );
  INV_X1 U7012 ( .A(n5956), .ZN(n5957) );
  NAND2_X1 U7013 ( .A1(n6015), .A2(n5957), .ZN(n5958) );
  NAND2_X1 U7014 ( .A1(n5959), .A2(n5958), .ZN(n5980) );
  NAND2_X1 U7015 ( .A1(n5980), .A2(REIP_REG_13__SCAN_IN), .ZN(n5964) );
  NAND2_X1 U7016 ( .A1(n6032), .A2(EBX_REG_13__SCAN_IN), .ZN(n5961) );
  AOI21_X1 U7017 ( .B1(n6008), .B2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6018), 
        .ZN(n5960) );
  OAI211_X1 U7018 ( .C1(n6049), .C2(n6024), .A(n5961), .B(n5960), .ZN(n5962)
         );
  INV_X1 U7019 ( .A(n5962), .ZN(n5963) );
  NAND2_X1 U7020 ( .A1(n5964), .A2(n5963), .ZN(n5965) );
  OR2_X1 U7021 ( .A1(n5966), .A2(n5965), .ZN(n5967) );
  AOI21_X1 U7022 ( .B1(n6051), .B2(n3979), .A(n5967), .ZN(n5968) );
  OAI21_X1 U7023 ( .B1(n5969), .B2(n6030), .A(n5968), .ZN(U2814) );
  AOI22_X1 U7024 ( .A1(EBX_REG_12__SCAN_IN), .A2(n6032), .B1(
        REIP_REG_12__SCAN_IN), .B2(n5980), .ZN(n5970) );
  NAND2_X1 U7025 ( .A1(n4889), .A2(n5970), .ZN(n5973) );
  INV_X1 U7026 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5971) );
  NOR2_X1 U7027 ( .A1(n6036), .A2(n5971), .ZN(n5972) );
  AOI211_X1 U7028 ( .C1(n6033), .C2(n6187), .A(n5973), .B(n5972), .ZN(n5978)
         );
  INV_X1 U7029 ( .A(n5974), .ZN(n5975) );
  AOI22_X1 U7030 ( .A1(n5976), .A2(n3979), .B1(n5975), .B2(n6044), .ZN(n5977)
         );
  OAI211_X1 U7031 ( .C1(REIP_REG_12__SCAN_IN), .C2(n5979), .A(n5978), .B(n5977), .ZN(U2815) );
  NAND2_X1 U7032 ( .A1(n6000), .A2(n6466), .ZN(n5989) );
  AOI22_X1 U7033 ( .A1(EBX_REG_11__SCAN_IN), .A2(n6032), .B1(
        REIP_REG_11__SCAN_IN), .B2(n5980), .ZN(n5982) );
  AOI21_X1 U7034 ( .B1(n6053), .B2(n6033), .A(n6018), .ZN(n5981) );
  OAI211_X1 U7035 ( .C1(n5983), .C2(n6036), .A(n5982), .B(n5981), .ZN(n5984)
         );
  INV_X1 U7036 ( .A(n5984), .ZN(n5988) );
  OAI22_X1 U7037 ( .A1(n6150), .A2(n5985), .B1(n6030), .B2(n6149), .ZN(n5986)
         );
  INV_X1 U7038 ( .A(n5986), .ZN(n5987) );
  OAI211_X1 U7039 ( .C1(n5990), .C2(n5989), .A(n5988), .B(n5987), .ZN(U2816)
         );
  AOI21_X1 U7040 ( .B1(n5993), .B2(n5992), .A(n5991), .ZN(n6210) );
  OAI21_X1 U7041 ( .B1(n6005), .B2(n6064), .A(n4889), .ZN(n5996) );
  NOR2_X1 U7042 ( .A1(n6036), .A2(n5994), .ZN(n5995) );
  AOI211_X1 U7043 ( .C1(n6210), .C2(n6033), .A(n5996), .B(n5995), .ZN(n6003)
         );
  INV_X1 U7044 ( .A(n5997), .ZN(n6062) );
  AOI22_X1 U7045 ( .A1(n6062), .A2(n3979), .B1(n6044), .B2(n5998), .ZN(n6002)
         );
  OAI21_X1 U7046 ( .B1(REIP_REG_9__SCAN_IN), .B2(n6000), .A(n5999), .ZN(n6001)
         );
  NAND3_X1 U7047 ( .A1(n6003), .A2(n6002), .A3(n6001), .ZN(U2818) );
  OAI22_X1 U7048 ( .A1(n6006), .A2(n6005), .B1(n6024), .B2(n6004), .ZN(n6007)
         );
  AOI211_X1 U7049 ( .C1(n6008), .C2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6018), 
        .B(n6007), .ZN(n6011) );
  NAND2_X1 U7050 ( .A1(n6009), .A2(n6459), .ZN(n6010) );
  OAI211_X1 U7051 ( .C1(n6012), .C2(n6459), .A(n6011), .B(n6010), .ZN(n6013)
         );
  AOI21_X1 U7052 ( .B1(n6156), .B2(n3979), .A(n6013), .ZN(n6014) );
  OAI21_X1 U7053 ( .B1(n6160), .B2(n6030), .A(n6014), .ZN(U2821) );
  INV_X1 U7054 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6631) );
  OAI21_X1 U7055 ( .B1(n6016), .B2(n6020), .A(n6015), .ZN(n6048) );
  OAI22_X1 U7056 ( .A1(n6631), .A2(n6036), .B1(n6456), .B2(n6048), .ZN(n6017)
         );
  AOI211_X1 U7057 ( .C1(n6019), .C2(n6039), .A(n6018), .B(n6017), .ZN(n6029)
         );
  INV_X1 U7058 ( .A(n6165), .ZN(n6027) );
  INV_X1 U7059 ( .A(n6041), .ZN(n6026) );
  NOR3_X1 U7060 ( .A1(n6021), .A2(REIP_REG_4__SCAN_IN), .A3(n6020), .ZN(n6022)
         );
  AOI21_X1 U7061 ( .B1(n6032), .B2(EBX_REG_4__SCAN_IN), .A(n6022), .ZN(n6023)
         );
  OAI21_X1 U7062 ( .B1(n6024), .B2(n6236), .A(n6023), .ZN(n6025) );
  AOI21_X1 U7063 ( .B1(n6027), .B2(n6026), .A(n6025), .ZN(n6028) );
  OAI211_X1 U7064 ( .C1(n6170), .C2(n6030), .A(n6029), .B(n6028), .ZN(U2823)
         );
  INV_X1 U7065 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6454) );
  NAND2_X1 U7066 ( .A1(n6031), .A2(REIP_REG_2__SCAN_IN), .ZN(n6047) );
  AOI22_X1 U7067 ( .A1(n6244), .A2(n6033), .B1(n6032), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n6034) );
  OAI21_X1 U7068 ( .B1(n6036), .B2(n6035), .A(n6034), .ZN(n6037) );
  AOI21_X1 U7069 ( .B1(n6039), .B2(n6038), .A(n6037), .ZN(n6040) );
  OAI21_X1 U7070 ( .B1(n6042), .B2(n6041), .A(n6040), .ZN(n6043) );
  AOI21_X1 U7071 ( .B1(n6045), .B2(n6044), .A(n6043), .ZN(n6046) );
  OAI221_X1 U7072 ( .B1(n6048), .B2(n6454), .C1(n6048), .C2(n6047), .A(n6046), 
        .ZN(U2824) );
  NOR2_X1 U7073 ( .A1(n6055), .A2(n6049), .ZN(n6050) );
  AOI21_X1 U7074 ( .B1(n6051), .B2(n6061), .A(n6050), .ZN(n6052) );
  OAI21_X1 U7075 ( .B1(n6065), .B2(n6556), .A(n6052), .ZN(U2846) );
  INV_X1 U7076 ( .A(n6053), .ZN(n6054) );
  OAI22_X1 U7077 ( .A1(n6150), .A2(n6056), .B1(n6055), .B2(n6054), .ZN(n6057)
         );
  INV_X1 U7078 ( .A(n6057), .ZN(n6058) );
  OAI21_X1 U7079 ( .B1(n6065), .B2(n6059), .A(n6058), .ZN(U2848) );
  AOI22_X1 U7080 ( .A1(n6062), .A2(n6061), .B1(n6060), .B2(n6210), .ZN(n6063)
         );
  OAI21_X1 U7081 ( .B1(n6065), .B2(n6064), .A(n6063), .ZN(U2850) );
  AOI22_X1 U7082 ( .A1(n6066), .A2(n6074), .B1(n6073), .B2(DATAI_18_), .ZN(
        n6068) );
  AOI22_X1 U7083 ( .A1(n6077), .A2(DATAI_2_), .B1(n6076), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6067) );
  NAND2_X1 U7084 ( .A1(n6068), .A2(n6067), .ZN(U2873) );
  AOI22_X1 U7085 ( .A1(n6069), .A2(n6074), .B1(n6073), .B2(DATAI_17_), .ZN(
        n6071) );
  AOI22_X1 U7086 ( .A1(n6077), .A2(DATAI_1_), .B1(n6076), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6070) );
  NAND2_X1 U7087 ( .A1(n6071), .A2(n6070), .ZN(U2874) );
  INV_X1 U7088 ( .A(n6072), .ZN(n6075) );
  AOI22_X1 U7089 ( .A1(n6075), .A2(n6074), .B1(n6073), .B2(DATAI_16_), .ZN(
        n6079) );
  AOI22_X1 U7090 ( .A1(n6077), .A2(DATAI_0_), .B1(n6076), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6078) );
  NAND2_X1 U7091 ( .A1(n6079), .A2(n6078), .ZN(U2875) );
  AOI22_X1 U7092 ( .A1(n6115), .A2(DATAO_REG_30__SCAN_IN), .B1(n6083), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n6080) );
  OAI21_X1 U7093 ( .B1(n6413), .B2(n6643), .A(n6080), .ZN(U2893) );
  INV_X1 U7094 ( .A(UWORD_REG_6__SCAN_IN), .ZN(n6627) );
  AOI22_X1 U7095 ( .A1(n6115), .A2(DATAO_REG_22__SCAN_IN), .B1(n6083), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n6081) );
  OAI21_X1 U7096 ( .B1(n6413), .B2(n6627), .A(n6081), .ZN(U2901) );
  INV_X1 U7097 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n6597) );
  AOI22_X1 U7098 ( .A1(n6083), .A2(EAX_REG_21__SCAN_IN), .B1(n6112), .B2(
        UWORD_REG_5__SCAN_IN), .ZN(n6082) );
  OAI21_X1 U7099 ( .B1(n6597), .B2(n6095), .A(n6082), .ZN(U2902) );
  INV_X1 U7100 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n6557) );
  AOI22_X1 U7101 ( .A1(n6083), .A2(EAX_REG_17__SCAN_IN), .B1(n6112), .B2(
        UWORD_REG_1__SCAN_IN), .ZN(n6084) );
  OAI21_X1 U7102 ( .B1(n6557), .B2(n6095), .A(n6084), .ZN(U2906) );
  AOI22_X1 U7103 ( .A1(n6116), .A2(LWORD_REG_15__SCAN_IN), .B1(n6115), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6085) );
  OAI21_X1 U7104 ( .B1(n6086), .B2(n6118), .A(n6085), .ZN(U2908) );
  AOI22_X1 U7105 ( .A1(n6116), .A2(LWORD_REG_14__SCAN_IN), .B1(n6115), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6087) );
  OAI21_X1 U7106 ( .B1(n6088), .B2(n6118), .A(n6087), .ZN(U2909) );
  AOI22_X1 U7107 ( .A1(n6116), .A2(LWORD_REG_13__SCAN_IN), .B1(n6115), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6089) );
  OAI21_X1 U7108 ( .B1(n6090), .B2(n6118), .A(n6089), .ZN(U2910) );
  AOI22_X1 U7109 ( .A1(n6112), .A2(LWORD_REG_12__SCAN_IN), .B1(n6115), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6091) );
  OAI21_X1 U7110 ( .B1(n6092), .B2(n6118), .A(n6091), .ZN(U2911) );
  INV_X1 U7111 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n6560) );
  AOI22_X1 U7112 ( .A1(EAX_REG_11__SCAN_IN), .A2(n6093), .B1(n6116), .B2(
        LWORD_REG_11__SCAN_IN), .ZN(n6094) );
  OAI21_X1 U7113 ( .B1(n6560), .B2(n6095), .A(n6094), .ZN(U2912) );
  INV_X1 U7114 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6097) );
  AOI22_X1 U7115 ( .A1(n6112), .A2(LWORD_REG_10__SCAN_IN), .B1(n6115), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6096) );
  OAI21_X1 U7116 ( .B1(n6097), .B2(n6118), .A(n6096), .ZN(U2913) );
  AOI22_X1 U7117 ( .A1(n6112), .A2(LWORD_REG_9__SCAN_IN), .B1(n6115), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6098) );
  OAI21_X1 U7118 ( .B1(n6099), .B2(n6118), .A(n6098), .ZN(U2914) );
  AOI22_X1 U7119 ( .A1(n6112), .A2(LWORD_REG_8__SCAN_IN), .B1(n6115), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6100) );
  OAI21_X1 U7120 ( .B1(n6101), .B2(n6118), .A(n6100), .ZN(U2915) );
  AOI22_X1 U7121 ( .A1(n6112), .A2(LWORD_REG_7__SCAN_IN), .B1(n6115), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6102) );
  OAI21_X1 U7122 ( .B1(n3745), .B2(n6118), .A(n6102), .ZN(U2916) );
  AOI22_X1 U7123 ( .A1(n6112), .A2(LWORD_REG_6__SCAN_IN), .B1(n6115), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6103) );
  OAI21_X1 U7124 ( .B1(n3728), .B2(n6118), .A(n6103), .ZN(U2917) );
  AOI22_X1 U7125 ( .A1(n6112), .A2(LWORD_REG_5__SCAN_IN), .B1(n6115), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6104) );
  OAI21_X1 U7126 ( .B1(n6105), .B2(n6118), .A(n6104), .ZN(U2918) );
  AOI22_X1 U7127 ( .A1(n6112), .A2(LWORD_REG_4__SCAN_IN), .B1(n6115), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6106) );
  OAI21_X1 U7128 ( .B1(n6107), .B2(n6118), .A(n6106), .ZN(U2919) );
  AOI22_X1 U7129 ( .A1(n6112), .A2(LWORD_REG_3__SCAN_IN), .B1(n6115), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6108) );
  OAI21_X1 U7130 ( .B1(n6109), .B2(n6118), .A(n6108), .ZN(U2920) );
  AOI22_X1 U7131 ( .A1(n6112), .A2(LWORD_REG_2__SCAN_IN), .B1(n6115), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6110) );
  OAI21_X1 U7132 ( .B1(n6111), .B2(n6118), .A(n6110), .ZN(U2921) );
  AOI22_X1 U7133 ( .A1(n6112), .A2(LWORD_REG_1__SCAN_IN), .B1(n6115), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6113) );
  OAI21_X1 U7134 ( .B1(n6114), .B2(n6118), .A(n6113), .ZN(U2922) );
  AOI22_X1 U7135 ( .A1(n6116), .A2(LWORD_REG_0__SCAN_IN), .B1(n6115), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6117) );
  OAI21_X1 U7136 ( .B1(n6119), .B2(n6118), .A(n6117), .ZN(U2923) );
  INV_X1 U7137 ( .A(n6120), .ZN(n6145) );
  AOI22_X1 U7138 ( .A1(UWORD_REG_1__SCAN_IN), .A2(n6145), .B1(n6144), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6121) );
  OAI21_X1 U7139 ( .B1(n6143), .B2(n6602), .A(n6121), .ZN(U2925) );
  AOI22_X1 U7140 ( .A1(UWORD_REG_2__SCAN_IN), .A2(n6145), .B1(n6144), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6122) );
  OAI21_X1 U7141 ( .B1(n6143), .B2(n6584), .A(n6122), .ZN(U2926) );
  AOI22_X1 U7142 ( .A1(UWORD_REG_3__SCAN_IN), .A2(n6145), .B1(n6144), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n6123) );
  OAI21_X1 U7143 ( .B1(n6143), .B2(n6134), .A(n6123), .ZN(U2927) );
  AOI22_X1 U7144 ( .A1(UWORD_REG_4__SCAN_IN), .A2(n6145), .B1(n6144), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n6124) );
  OAI21_X1 U7145 ( .B1(n6143), .B2(n6634), .A(n6124), .ZN(U2928) );
  AOI22_X1 U7146 ( .A1(UWORD_REG_5__SCAN_IN), .A2(n6145), .B1(n6144), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n6125) );
  OAI21_X1 U7147 ( .B1(n6143), .B2(n6137), .A(n6125), .ZN(U2929) );
  AOI22_X1 U7148 ( .A1(UWORD_REG_6__SCAN_IN), .A2(n6145), .B1(n6144), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n6126) );
  OAI21_X1 U7149 ( .B1(n6143), .B2(n6600), .A(n6126), .ZN(U2930) );
  AOI22_X1 U7150 ( .A1(UWORD_REG_7__SCAN_IN), .A2(n6145), .B1(n6144), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n6127) );
  OAI21_X1 U7151 ( .B1(n6143), .B2(n6141), .A(n6127), .ZN(U2931) );
  INV_X1 U7152 ( .A(DATAI_10_), .ZN(n6585) );
  AOI22_X1 U7153 ( .A1(UWORD_REG_10__SCAN_IN), .A2(n6145), .B1(n6144), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n6128) );
  OAI21_X1 U7154 ( .B1(n6143), .B2(n6585), .A(n6128), .ZN(U2934) );
  AOI22_X1 U7155 ( .A1(LWORD_REG_0__SCAN_IN), .A2(n6145), .B1(n6144), .B2(
        EAX_REG_0__SCAN_IN), .ZN(n6129) );
  OAI21_X1 U7156 ( .B1(n6143), .B2(n6130), .A(n6129), .ZN(U2939) );
  AOI22_X1 U7157 ( .A1(LWORD_REG_1__SCAN_IN), .A2(n6145), .B1(n6144), .B2(
        EAX_REG_1__SCAN_IN), .ZN(n6131) );
  OAI21_X1 U7158 ( .B1(n6143), .B2(n6602), .A(n6131), .ZN(U2940) );
  AOI22_X1 U7159 ( .A1(LWORD_REG_2__SCAN_IN), .A2(n6145), .B1(n6144), .B2(
        EAX_REG_2__SCAN_IN), .ZN(n6132) );
  OAI21_X1 U7160 ( .B1(n6143), .B2(n6584), .A(n6132), .ZN(U2941) );
  AOI22_X1 U7161 ( .A1(LWORD_REG_3__SCAN_IN), .A2(n6139), .B1(n6144), .B2(
        EAX_REG_3__SCAN_IN), .ZN(n6133) );
  OAI21_X1 U7162 ( .B1(n6143), .B2(n6134), .A(n6133), .ZN(U2942) );
  AOI22_X1 U7163 ( .A1(LWORD_REG_4__SCAN_IN), .A2(n6139), .B1(n6144), .B2(
        EAX_REG_4__SCAN_IN), .ZN(n6135) );
  OAI21_X1 U7164 ( .B1(n6143), .B2(n6634), .A(n6135), .ZN(U2943) );
  AOI22_X1 U7165 ( .A1(LWORD_REG_5__SCAN_IN), .A2(n6139), .B1(n6144), .B2(
        EAX_REG_5__SCAN_IN), .ZN(n6136) );
  OAI21_X1 U7166 ( .B1(n6143), .B2(n6137), .A(n6136), .ZN(U2944) );
  AOI22_X1 U7167 ( .A1(LWORD_REG_6__SCAN_IN), .A2(n6139), .B1(n6144), .B2(
        EAX_REG_6__SCAN_IN), .ZN(n6138) );
  OAI21_X1 U7168 ( .B1(n6143), .B2(n6600), .A(n6138), .ZN(U2945) );
  AOI22_X1 U7169 ( .A1(LWORD_REG_7__SCAN_IN), .A2(n6139), .B1(n6144), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n6140) );
  OAI21_X1 U7170 ( .B1(n6143), .B2(n6141), .A(n6140), .ZN(U2946) );
  AOI22_X1 U7171 ( .A1(LWORD_REG_10__SCAN_IN), .A2(n6145), .B1(n6144), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n6142) );
  OAI21_X1 U7172 ( .B1(n6143), .B2(n6585), .A(n6142), .ZN(U2949) );
  AOI22_X1 U7173 ( .A1(LWORD_REG_11__SCAN_IN), .A2(n6145), .B1(n6144), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n6148) );
  NAND2_X1 U7174 ( .A1(n6146), .A2(DATAI_11_), .ZN(n6147) );
  NAND2_X1 U7175 ( .A1(n6148), .A2(n6147), .ZN(U2950) );
  AOI22_X1 U7176 ( .A1(n6189), .A2(REIP_REG_11__SCAN_IN), .B1(n6171), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6153) );
  OAI22_X1 U7177 ( .A1(n6150), .A2(n6164), .B1(n6182), .B2(n6149), .ZN(n6151)
         );
  INV_X1 U7178 ( .A(n6151), .ZN(n6152) );
  OAI211_X1 U7179 ( .C1(n6154), .C2(n6166), .A(n6153), .B(n6152), .ZN(U2975)
         );
  AOI22_X1 U7180 ( .A1(n6189), .A2(REIP_REG_6__SCAN_IN), .B1(n6171), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6159) );
  INV_X1 U7181 ( .A(n6155), .ZN(n6157) );
  AOI22_X1 U7182 ( .A1(n6157), .A2(n6178), .B1(n6176), .B2(n6156), .ZN(n6158)
         );
  OAI211_X1 U7183 ( .C1(n6182), .C2(n6160), .A(n6159), .B(n6158), .ZN(U2980)
         );
  AOI22_X1 U7184 ( .A1(n6189), .A2(REIP_REG_4__SCAN_IN), .B1(n6171), .B2(
        PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6169) );
  OAI21_X1 U7185 ( .B1(n6163), .B2(n6162), .A(n6161), .ZN(n6235) );
  OAI22_X1 U7186 ( .A1(n6235), .A2(n6166), .B1(n6165), .B2(n6164), .ZN(n6167)
         );
  INV_X1 U7187 ( .A(n6167), .ZN(n6168) );
  OAI211_X1 U7188 ( .C1(n6182), .C2(n6170), .A(n6169), .B(n6168), .ZN(U2982)
         );
  AOI22_X1 U7189 ( .A1(n6189), .A2(REIP_REG_2__SCAN_IN), .B1(n6171), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6180) );
  XOR2_X1 U7190 ( .A(n6172), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n6174) );
  XNOR2_X1 U7191 ( .A(n6174), .B(n6173), .ZN(n6264) );
  INV_X1 U7192 ( .A(n6175), .ZN(n6177) );
  AOI22_X1 U7193 ( .A1(n6178), .A2(n6264), .B1(n6177), .B2(n6176), .ZN(n6179)
         );
  OAI211_X1 U7194 ( .C1(n6182), .C2(n6181), .A(n6180), .B(n6179), .ZN(U2984)
         );
  AOI221_X1 U7195 ( .B1(n6260), .B2(n6185), .C1(n6184), .C2(n6185), .A(n6183), 
        .ZN(n6193) );
  AOI21_X1 U7196 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6186), .A(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6192) );
  AOI22_X1 U7197 ( .A1(n6188), .A2(n6263), .B1(n6258), .B2(n6187), .ZN(n6191)
         );
  NAND2_X1 U7198 ( .A1(n6189), .A2(REIP_REG_12__SCAN_IN), .ZN(n6190) );
  OAI211_X1 U7199 ( .C1(n6193), .C2(n6192), .A(n6191), .B(n6190), .ZN(U3006)
         );
  INV_X1 U7200 ( .A(n6194), .ZN(n6200) );
  NOR2_X1 U7201 ( .A1(n6200), .A2(n6253), .ZN(n6227) );
  NAND2_X1 U7202 ( .A1(n6202), .A2(n6227), .ZN(n6215) );
  AOI22_X1 U7203 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n4002), .B1(
        INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6195), .ZN(n6207) );
  INV_X1 U7204 ( .A(n6196), .ZN(n6198) );
  AOI21_X1 U7205 ( .B1(n6258), .B2(n6198), .A(n6197), .ZN(n6206) );
  NOR2_X1 U7206 ( .A1(n6199), .A2(n6255), .ZN(n6233) );
  AOI211_X1 U7207 ( .C1(n6201), .C2(n6200), .A(n6233), .B(n6262), .ZN(n6232)
         );
  OAI21_X1 U7208 ( .B1(n6203), .B2(n6202), .A(n6232), .ZN(n6211) );
  AOI22_X1 U7209 ( .A1(n6204), .A2(n6263), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6211), .ZN(n6205) );
  OAI211_X1 U7210 ( .C1(n6215), .C2(n6207), .A(n6206), .B(n6205), .ZN(U3008)
         );
  INV_X1 U7211 ( .A(n6208), .ZN(n6209) );
  AOI21_X1 U7212 ( .B1(n6258), .B2(n6210), .A(n6209), .ZN(n6214) );
  AOI22_X1 U7213 ( .A1(n6212), .A2(n6263), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n6211), .ZN(n6213) );
  OAI211_X1 U7214 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6215), .A(n6214), 
        .B(n6213), .ZN(U3009) );
  INV_X1 U7215 ( .A(n6216), .ZN(n6217) );
  AOI222_X1 U7216 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6189), .B1(n6258), .B2(
        n6218), .C1(n6263), .C2(n6217), .ZN(n6221) );
  OAI211_X1 U7217 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n6227), .B(n6219), .ZN(n6220) );
  OAI211_X1 U7218 ( .C1(n6232), .C2(n6222), .A(n6221), .B(n6220), .ZN(U3010)
         );
  INV_X1 U7219 ( .A(n6223), .ZN(n6224) );
  AOI21_X1 U7220 ( .B1(n6258), .B2(n6225), .A(n6224), .ZN(n6230) );
  INV_X1 U7221 ( .A(n6226), .ZN(n6228) );
  AOI22_X1 U7222 ( .A1(n6228), .A2(n6263), .B1(n6227), .B2(n6231), .ZN(n6229)
         );
  OAI211_X1 U7223 ( .C1(n6232), .C2(n6231), .A(n6230), .B(n6229), .ZN(U3011)
         );
  NOR2_X1 U7224 ( .A1(n6233), .A2(n6262), .ZN(n6251) );
  AOI211_X1 U7225 ( .C1(n6252), .C2(n6241), .A(n6234), .B(n6253), .ZN(n6239)
         );
  NOR2_X1 U7226 ( .A1(n6235), .A2(n6242), .ZN(n6238) );
  OAI22_X1 U7227 ( .A1(n6246), .A2(n6236), .B1(n6456), .B2(n4889), .ZN(n6237)
         );
  NOR3_X1 U7228 ( .A1(n6239), .A2(n6238), .A3(n6237), .ZN(n6240) );
  OAI21_X1 U7229 ( .B1(n6251), .B2(n6241), .A(n6240), .ZN(U3014) );
  NOR2_X1 U7230 ( .A1(n6243), .A2(n6242), .ZN(n6249) );
  INV_X1 U7231 ( .A(n6244), .ZN(n6245) );
  OAI22_X1 U7232 ( .A1(n6246), .A2(n6245), .B1(n6454), .B2(n4889), .ZN(n6247)
         );
  AOI21_X1 U7233 ( .B1(n6249), .B2(n6248), .A(n6247), .ZN(n6250) );
  OAI221_X1 U7234 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n6253), .C1(n6252), .C2(n6251), .A(n6250), .ZN(U3015) );
  NAND2_X1 U7235 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6254), .ZN(n6267)
         );
  NAND2_X1 U7236 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6256) );
  OAI21_X1 U7237 ( .B1(n6257), .B2(n6256), .A(n6255), .ZN(n6261) );
  AOI222_X1 U7238 ( .A1(n6261), .A2(n6260), .B1(REIP_REG_2__SCAN_IN), .B2(
        n6018), .C1(n6259), .C2(n6258), .ZN(n6266) );
  AOI22_X1 U7239 ( .A1(n6264), .A2(n6263), .B1(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .B2(n6262), .ZN(n6265) );
  OAI211_X1 U7240 ( .C1(INSTADDRPOINTER_REG_2__SCAN_IN), .C2(n6267), .A(n6266), 
        .B(n6265), .ZN(U3016) );
  NOR2_X1 U7241 ( .A1(n6412), .A2(n6268), .ZN(U3019) );
  AOI22_X1 U7242 ( .A1(n6286), .A2(n6269), .B1(n6296), .B2(n6283), .ZN(n6271)
         );
  AOI22_X1 U7243 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6288), .B1(n6318), 
        .B2(n6287), .ZN(n6270) );
  OAI211_X1 U7244 ( .C1(n6291), .C2(n6321), .A(n6271), .B(n6270), .ZN(U3045)
         );
  AOI22_X1 U7245 ( .A1(n6286), .A2(n6272), .B1(n6300), .B2(n6283), .ZN(n6274)
         );
  AOI22_X1 U7246 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6288), .B1(n6343), 
        .B2(n6287), .ZN(n6273) );
  OAI211_X1 U7247 ( .C1(n6291), .C2(n6346), .A(n6274), .B(n6273), .ZN(U3046)
         );
  AOI22_X1 U7248 ( .A1(n6286), .A2(n6276), .B1(n6275), .B2(n6283), .ZN(n6278)
         );
  AOI22_X1 U7249 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6288), .B1(n6357), 
        .B2(n6287), .ZN(n6277) );
  OAI211_X1 U7250 ( .C1(n6291), .C2(n6360), .A(n6278), .B(n6277), .ZN(U3048)
         );
  AOI22_X1 U7251 ( .A1(n6286), .A2(n6280), .B1(n6279), .B2(n6283), .ZN(n6282)
         );
  AOI22_X1 U7252 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6288), .B1(n6371), 
        .B2(n6287), .ZN(n6281) );
  OAI211_X1 U7253 ( .C1(n6291), .C2(n6374), .A(n6282), .B(n6281), .ZN(U3050)
         );
  AOI22_X1 U7254 ( .A1(n6286), .A2(n6285), .B1(n6284), .B2(n6283), .ZN(n6290)
         );
  AOI22_X1 U7255 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6288), .B1(n6381), 
        .B2(n6287), .ZN(n6289) );
  OAI211_X1 U7256 ( .C1(n6291), .C2(n6386), .A(n6290), .B(n6289), .ZN(U3051)
         );
  AOI22_X1 U7257 ( .A1(n6336), .A2(n6306), .B1(n6292), .B2(n6304), .ZN(n6295)
         );
  AOI22_X1 U7258 ( .A1(n6309), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6293), 
        .B2(n6307), .ZN(n6294) );
  OAI211_X1 U7259 ( .C1(n6334), .C2(n6332), .A(n6295), .B(n6294), .ZN(U3068)
         );
  AOI22_X1 U7260 ( .A1(n6318), .A2(n6306), .B1(n6296), .B2(n6304), .ZN(n6299)
         );
  AOI22_X1 U7261 ( .A1(n6309), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6297), 
        .B2(n6307), .ZN(n6298) );
  OAI211_X1 U7262 ( .C1(n6316), .C2(n6332), .A(n6299), .B(n6298), .ZN(U3069)
         );
  AOI22_X1 U7263 ( .A1(n6343), .A2(n6306), .B1(n6300), .B2(n6304), .ZN(n6303)
         );
  AOI22_X1 U7264 ( .A1(n6309), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6301), 
        .B2(n6307), .ZN(n6302) );
  OAI211_X1 U7265 ( .C1(n6341), .C2(n6332), .A(n6303), .B(n6302), .ZN(U3070)
         );
  AOI22_X1 U7266 ( .A1(n6350), .A2(n6306), .B1(n6305), .B2(n6304), .ZN(n6311)
         );
  AOI22_X1 U7267 ( .A1(n6309), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6308), 
        .B2(n6307), .ZN(n6310) );
  OAI211_X1 U7268 ( .C1(n6348), .C2(n6332), .A(n6311), .B(n6310), .ZN(U3071)
         );
  OAI22_X1 U7269 ( .A1(n6326), .A2(n6334), .B1(n6325), .B2(n6333), .ZN(n6312)
         );
  INV_X1 U7270 ( .A(n6312), .ZN(n6314) );
  AOI22_X1 U7271 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6329), .B1(n6336), 
        .B2(n6328), .ZN(n6313) );
  OAI211_X1 U7272 ( .C1(n6339), .C2(n6332), .A(n6314), .B(n6313), .ZN(U3076)
         );
  OAI22_X1 U7273 ( .A1(n6326), .A2(n6316), .B1(n6325), .B2(n6315), .ZN(n6317)
         );
  INV_X1 U7274 ( .A(n6317), .ZN(n6320) );
  AOI22_X1 U7275 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6329), .B1(n6318), 
        .B2(n6328), .ZN(n6319) );
  OAI211_X1 U7276 ( .C1(n6321), .C2(n6332), .A(n6320), .B(n6319), .ZN(U3077)
         );
  OAI22_X1 U7277 ( .A1(n6326), .A2(n6355), .B1(n6325), .B2(n6354), .ZN(n6322)
         );
  INV_X1 U7278 ( .A(n6322), .ZN(n6324) );
  AOI22_X1 U7279 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6329), .B1(n6357), 
        .B2(n6328), .ZN(n6323) );
  OAI211_X1 U7280 ( .C1(n6360), .C2(n6332), .A(n6324), .B(n6323), .ZN(U3080)
         );
  OAI22_X1 U7281 ( .A1(n6326), .A2(n6369), .B1(n6325), .B2(n6368), .ZN(n6327)
         );
  INV_X1 U7282 ( .A(n6327), .ZN(n6331) );
  AOI22_X1 U7283 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6329), .B1(n6371), 
        .B2(n6328), .ZN(n6330) );
  OAI211_X1 U7284 ( .C1(n6374), .C2(n6332), .A(n6331), .B(n6330), .ZN(U3082)
         );
  OAI22_X1 U7285 ( .A1(n6378), .A2(n6334), .B1(n6333), .B2(n6375), .ZN(n6335)
         );
  INV_X1 U7286 ( .A(n6335), .ZN(n6338) );
  AOI22_X1 U7287 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6382), .B1(n6336), 
        .B2(n6380), .ZN(n6337) );
  OAI211_X1 U7288 ( .C1(n6339), .C2(n6385), .A(n6338), .B(n6337), .ZN(U3108)
         );
  OAI22_X1 U7289 ( .A1(n6378), .A2(n6341), .B1(n6340), .B2(n6375), .ZN(n6342)
         );
  INV_X1 U7290 ( .A(n6342), .ZN(n6345) );
  AOI22_X1 U7291 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6382), .B1(n6343), 
        .B2(n6380), .ZN(n6344) );
  OAI211_X1 U7292 ( .C1(n6346), .C2(n6385), .A(n6345), .B(n6344), .ZN(U3110)
         );
  OAI22_X1 U7293 ( .A1(n6378), .A2(n6348), .B1(n6347), .B2(n6375), .ZN(n6349)
         );
  INV_X1 U7294 ( .A(n6349), .ZN(n6352) );
  AOI22_X1 U7295 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6382), .B1(n6350), 
        .B2(n6380), .ZN(n6351) );
  OAI211_X1 U7296 ( .C1(n6353), .C2(n6385), .A(n6352), .B(n6351), .ZN(U3111)
         );
  OAI22_X1 U7297 ( .A1(n6378), .A2(n6355), .B1(n6354), .B2(n6375), .ZN(n6356)
         );
  INV_X1 U7298 ( .A(n6356), .ZN(n6359) );
  AOI22_X1 U7299 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6382), .B1(n6357), 
        .B2(n6380), .ZN(n6358) );
  OAI211_X1 U7300 ( .C1(n6360), .C2(n6385), .A(n6359), .B(n6358), .ZN(U3112)
         );
  OAI22_X1 U7301 ( .A1(n6378), .A2(n6362), .B1(n6361), .B2(n6375), .ZN(n6363)
         );
  INV_X1 U7302 ( .A(n6363), .ZN(n6366) );
  AOI22_X1 U7303 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6382), .B1(n6364), 
        .B2(n6380), .ZN(n6365) );
  OAI211_X1 U7304 ( .C1(n6367), .C2(n6385), .A(n6366), .B(n6365), .ZN(U3113)
         );
  OAI22_X1 U7305 ( .A1(n6378), .A2(n6369), .B1(n6368), .B2(n6375), .ZN(n6370)
         );
  INV_X1 U7306 ( .A(n6370), .ZN(n6373) );
  AOI22_X1 U7307 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6382), .B1(n6371), 
        .B2(n6380), .ZN(n6372) );
  OAI211_X1 U7308 ( .C1(n6374), .C2(n6385), .A(n6373), .B(n6372), .ZN(U3114)
         );
  OAI22_X1 U7309 ( .A1(n6378), .A2(n6377), .B1(n6376), .B2(n6375), .ZN(n6379)
         );
  INV_X1 U7310 ( .A(n6379), .ZN(n6384) );
  AOI22_X1 U7311 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6382), .B1(n6381), 
        .B2(n6380), .ZN(n6383) );
  OAI211_X1 U7312 ( .C1(n6386), .C2(n6385), .A(n6384), .B(n6383), .ZN(U3115)
         );
  INV_X1 U7313 ( .A(n6387), .ZN(n6389) );
  NOR3_X1 U7314 ( .A1(n6389), .A2(n6388), .A3(n6691), .ZN(n6396) );
  INV_X1 U7315 ( .A(n6396), .ZN(n6394) );
  INV_X1 U7316 ( .A(n6390), .ZN(n6392) );
  OAI211_X1 U7317 ( .C1(n6394), .C2(n6393), .A(n6392), .B(n6391), .ZN(n6395)
         );
  OAI21_X1 U7318 ( .B1(n6396), .B2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n6395), 
        .ZN(n6397) );
  AOI222_X1 U7319 ( .A1(n6399), .A2(n6398), .B1(n6399), .B2(n6397), .C1(n6398), 
        .C2(n6397), .ZN(n6400) );
  AOI222_X1 U7320 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6401), .B1(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n6400), .C1(n6401), .C2(n6400), 
        .ZN(n6411) );
  INV_X1 U7321 ( .A(n6402), .ZN(n6403) );
  NOR2_X1 U7322 ( .A1(n6404), .A2(n6403), .ZN(n6407) );
  OAI21_X1 U7323 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6405), 
        .ZN(n6406) );
  NAND4_X1 U7324 ( .A1(n6409), .A2(n6408), .A3(n6407), .A4(n6406), .ZN(n6410)
         );
  AOI21_X1 U7325 ( .B1(n6412), .B2(n6411), .A(n6410), .ZN(n6422) );
  INV_X1 U7326 ( .A(n6422), .ZN(n6414) );
  OAI22_X1 U7327 ( .A1(n6414), .A2(n6424), .B1(n6413), .B2(n6441), .ZN(n6415)
         );
  OAI21_X1 U7328 ( .B1(n6417), .B2(n6416), .A(n6415), .ZN(n6511) );
  OAI21_X1 U7329 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6441), .A(n6511), .ZN(
        n6423) );
  AOI221_X1 U7330 ( .B1(n6419), .B2(STATE2_REG_0__SCAN_IN), .C1(n6423), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6418), .ZN(n6421) );
  OAI211_X1 U7331 ( .C1(n6431), .C2(n6550), .A(n6529), .B(n6511), .ZN(n6420)
         );
  OAI211_X1 U7332 ( .C1(n6422), .C2(n6424), .A(n6421), .B(n6420), .ZN(U3148)
         );
  NAND2_X1 U7333 ( .A1(n6423), .A2(STATE2_REG_1__SCAN_IN), .ZN(n6429) );
  OAI21_X1 U7334 ( .B1(READY_N), .B2(n6425), .A(n6424), .ZN(n6427) );
  AOI21_X1 U7335 ( .B1(n6511), .B2(n6427), .A(n6426), .ZN(n6428) );
  OAI21_X1 U7336 ( .B1(n6434), .B2(n6429), .A(n6428), .ZN(U3149) );
  INV_X1 U7337 ( .A(n6430), .ZN(n6510) );
  OAI211_X1 U7338 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6441), .A(n6510), .B(
        n6431), .ZN(n6433) );
  OAI21_X1 U7339 ( .B1(n6434), .B2(n6433), .A(n6432), .ZN(U3150) );
  INV_X1 U7340 ( .A(n6509), .ZN(n6435) );
  AND2_X1 U7341 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6435), .ZN(U3151) );
  INV_X1 U7342 ( .A(DATAWIDTH_REG_30__SCAN_IN), .ZN(n6612) );
  NOR2_X1 U7343 ( .A1(n6509), .A2(n6612), .ZN(U3152) );
  AND2_X1 U7344 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6435), .ZN(U3153) );
  AND2_X1 U7345 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6435), .ZN(U3154) );
  AND2_X1 U7346 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6435), .ZN(U3155) );
  AND2_X1 U7347 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6435), .ZN(U3156) );
  AND2_X1 U7348 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6435), .ZN(U3157) );
  AND2_X1 U7349 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6435), .ZN(U3158) );
  AND2_X1 U7350 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6435), .ZN(U3159) );
  AND2_X1 U7351 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6435), .ZN(U3160) );
  INV_X1 U7352 ( .A(DATAWIDTH_REG_21__SCAN_IN), .ZN(n6572) );
  NOR2_X1 U7353 ( .A1(n6509), .A2(n6572), .ZN(U3161) );
  AND2_X1 U7354 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6435), .ZN(U3162) );
  AND2_X1 U7355 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6435), .ZN(U3163) );
  AND2_X1 U7356 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6435), .ZN(U3164) );
  NOR2_X1 U7357 ( .A1(n6509), .A2(n6660), .ZN(U3165) );
  AND2_X1 U7358 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6435), .ZN(U3166) );
  AND2_X1 U7359 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6435), .ZN(U3167) );
  INV_X1 U7360 ( .A(DATAWIDTH_REG_14__SCAN_IN), .ZN(n6642) );
  NOR2_X1 U7361 ( .A1(n6509), .A2(n6642), .ZN(U3168) );
  AND2_X1 U7362 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6435), .ZN(U3169) );
  AND2_X1 U7363 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6435), .ZN(U3170) );
  AND2_X1 U7364 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6435), .ZN(U3171) );
  AND2_X1 U7365 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6435), .ZN(U3172) );
  AND2_X1 U7366 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6435), .ZN(U3173) );
  AND2_X1 U7367 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6435), .ZN(U3174) );
  AND2_X1 U7368 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6435), .ZN(U3175) );
  AND2_X1 U7369 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6435), .ZN(U3176) );
  NOR2_X1 U7370 ( .A1(n6509), .A2(n6646), .ZN(U3177) );
  AND2_X1 U7371 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6435), .ZN(U3178) );
  AND2_X1 U7372 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6435), .ZN(U3179) );
  AND2_X1 U7373 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6435), .ZN(U3180) );
  NOR2_X1 U7374 ( .A1(n6450), .A2(n6440), .ZN(n6444) );
  AOI22_X1 U7375 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6447) );
  AND2_X1 U7376 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6438) );
  INV_X1 U7377 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6539) );
  INV_X1 U7378 ( .A(NA_N), .ZN(n6591) );
  AOI211_X1 U7379 ( .C1(STATE_REG_2__SCAN_IN), .C2(n6591), .A(
        STATE_REG_0__SCAN_IN), .B(n6444), .ZN(n6449) );
  AOI221_X1 U7380 ( .B1(n6438), .B2(n6540), .C1(n6539), .C2(n6540), .A(n6449), 
        .ZN(n6436) );
  OAI21_X1 U7381 ( .B1(n6444), .B2(n6447), .A(n6436), .ZN(U3181) );
  NOR2_X1 U7382 ( .A1(n6442), .A2(n6539), .ZN(n6445) );
  NAND2_X1 U7383 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6437) );
  OAI21_X1 U7384 ( .B1(n6445), .B2(n6438), .A(n6437), .ZN(n6439) );
  OAI211_X1 U7385 ( .C1(n6440), .C2(n6441), .A(n6528), .B(n6439), .ZN(U3182)
         );
  AOI221_X1 U7386 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6441), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6443) );
  AOI221_X1 U7387 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6443), .C2(HOLD), .A(n6442), .ZN(n6448) );
  AOI21_X1 U7388 ( .B1(n6445), .B2(n6591), .A(n6444), .ZN(n6446) );
  OAI22_X1 U7389 ( .A1(n6449), .A2(n6448), .B1(n6447), .B2(n6446), .ZN(U3183)
         );
  NOR2_X1 U7390 ( .A1(n6450), .A2(n6540), .ZN(n6493) );
  INV_X1 U7391 ( .A(n6493), .ZN(n6504) );
  NAND2_X1 U7392 ( .A1(n6450), .A2(n6471), .ZN(n6495) );
  INV_X1 U7393 ( .A(n6495), .ZN(n6502) );
  AOI22_X1 U7394 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6502), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6540), .ZN(n6451) );
  OAI21_X1 U7395 ( .B1(n6513), .B2(n6504), .A(n6451), .ZN(U3184) );
  AOI22_X1 U7396 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6502), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6540), .ZN(n6452) );
  OAI21_X1 U7397 ( .B1(n5124), .B2(n6504), .A(n6452), .ZN(U3185) );
  AOI22_X1 U7398 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6502), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6540), .ZN(n6453) );
  OAI21_X1 U7399 ( .B1(n6454), .B2(n6504), .A(n6453), .ZN(U3186) );
  AOI22_X1 U7400 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6502), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6540), .ZN(n6455) );
  OAI21_X1 U7401 ( .B1(n6456), .B2(n6504), .A(n6455), .ZN(U3187) );
  INV_X1 U7402 ( .A(ADDRESS_REG_4__SCAN_IN), .ZN(n6577) );
  OAI222_X1 U7403 ( .A1(n6495), .A2(n6459), .B1(n6577), .B2(n6471), .C1(n6457), 
        .C2(n6504), .ZN(U3188) );
  AOI22_X1 U7404 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6502), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6540), .ZN(n6458) );
  OAI21_X1 U7405 ( .B1(n6459), .B2(n6504), .A(n6458), .ZN(U3189) );
  INV_X1 U7406 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n6559) );
  OAI222_X1 U7407 ( .A1(n6504), .A2(n6460), .B1(n6559), .B2(n6471), .C1(n6462), 
        .C2(n6495), .ZN(U3190) );
  AOI22_X1 U7408 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6502), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6540), .ZN(n6461) );
  OAI21_X1 U7409 ( .B1(n6462), .B2(n6504), .A(n6461), .ZN(U3191) );
  AOI22_X1 U7410 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6502), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6540), .ZN(n6463) );
  OAI21_X1 U7411 ( .B1(n6464), .B2(n6504), .A(n6463), .ZN(U3192) );
  AOI22_X1 U7412 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6493), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6540), .ZN(n6465) );
  OAI21_X1 U7413 ( .B1(n6466), .B2(n6495), .A(n6465), .ZN(U3193) );
  AOI22_X1 U7414 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6493), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6540), .ZN(n6467) );
  OAI21_X1 U7415 ( .B1(n6469), .B2(n6495), .A(n6467), .ZN(U3194) );
  AOI22_X1 U7416 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6502), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6540), .ZN(n6468) );
  OAI21_X1 U7417 ( .B1(n6469), .B2(n6504), .A(n6468), .ZN(U3195) );
  INV_X1 U7418 ( .A(ADDRESS_REG_12__SCAN_IN), .ZN(n6617) );
  OAI222_X1 U7419 ( .A1(n6504), .A2(n6472), .B1(n6617), .B2(n6471), .C1(n6470), 
        .C2(n6495), .ZN(U3196) );
  AOI22_X1 U7420 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6493), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6540), .ZN(n6473) );
  OAI21_X1 U7421 ( .B1(n6673), .B2(n6495), .A(n6473), .ZN(U3197) );
  AOI22_X1 U7422 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6502), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6540), .ZN(n6474) );
  OAI21_X1 U7423 ( .B1(n6673), .B2(n6504), .A(n6474), .ZN(U3198) );
  AOI22_X1 U7424 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6502), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6540), .ZN(n6475) );
  OAI21_X1 U7425 ( .B1(n6476), .B2(n6504), .A(n6475), .ZN(U3199) );
  AOI22_X1 U7426 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6502), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6540), .ZN(n6477) );
  OAI21_X1 U7427 ( .B1(n6478), .B2(n6504), .A(n6477), .ZN(U3200) );
  AOI22_X1 U7428 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6502), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6540), .ZN(n6479) );
  OAI21_X1 U7429 ( .B1(n6480), .B2(n6504), .A(n6479), .ZN(U3201) );
  INV_X1 U7430 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6482) );
  AOI22_X1 U7431 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6502), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6540), .ZN(n6481) );
  OAI21_X1 U7432 ( .B1(n6482), .B2(n6504), .A(n6481), .ZN(U3202) );
  AOI22_X1 U7433 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6493), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6540), .ZN(n6483) );
  OAI21_X1 U7434 ( .B1(n6484), .B2(n6495), .A(n6483), .ZN(U3203) );
  AOI22_X1 U7435 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6493), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6540), .ZN(n6485) );
  OAI21_X1 U7436 ( .B1(n6487), .B2(n6495), .A(n6485), .ZN(U3204) );
  AOI22_X1 U7437 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6502), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6540), .ZN(n6486) );
  OAI21_X1 U7438 ( .B1(n6487), .B2(n6504), .A(n6486), .ZN(U3205) );
  AOI22_X1 U7439 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6493), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6540), .ZN(n6488) );
  OAI21_X1 U7440 ( .B1(n6490), .B2(n6495), .A(n6488), .ZN(U3206) );
  AOI22_X1 U7441 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6502), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6540), .ZN(n6489) );
  OAI21_X1 U7442 ( .B1(n6490), .B2(n6504), .A(n6489), .ZN(U3207) );
  AOI22_X1 U7443 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6502), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6540), .ZN(n6491) );
  OAI21_X1 U7444 ( .B1(n6492), .B2(n6504), .A(n6491), .ZN(U3208) );
  AOI22_X1 U7445 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6493), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6540), .ZN(n6494) );
  OAI21_X1 U7446 ( .B1(n6497), .B2(n6495), .A(n6494), .ZN(U3209) );
  AOI22_X1 U7447 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6502), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6540), .ZN(n6496) );
  OAI21_X1 U7448 ( .B1(n6497), .B2(n6504), .A(n6496), .ZN(U3210) );
  AOI22_X1 U7449 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6502), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6540), .ZN(n6498) );
  OAI21_X1 U7450 ( .B1(n6499), .B2(n6504), .A(n6498), .ZN(U3211) );
  AOI22_X1 U7451 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6502), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6540), .ZN(n6500) );
  OAI21_X1 U7452 ( .B1(n6501), .B2(n6504), .A(n6500), .ZN(U3212) );
  AOI22_X1 U7453 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6502), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6540), .ZN(n6503) );
  OAI21_X1 U7454 ( .B1(n6505), .B2(n6504), .A(n6503), .ZN(U3213) );
  MUX2_X1 U7455 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(BE_N_REG_3__SCAN_IN), .S(
        n6540), .Z(U3445) );
  MUX2_X1 U7456 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6540), .Z(U3446) );
  MUX2_X1 U7457 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6540), .Z(U3447) );
  MUX2_X1 U7458 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6540), .Z(U3448) );
  OAI21_X1 U7459 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6509), .A(n6507), .ZN(
        n6506) );
  INV_X1 U7460 ( .A(n6506), .ZN(U3451) );
  OAI21_X1 U7461 ( .B1(n6509), .B2(n6508), .A(n6507), .ZN(U3452) );
  OAI221_X1 U7462 ( .B1(n6512), .B2(STATE2_REG_0__SCAN_IN), .C1(n6512), .C2(
        n6511), .A(n6510), .ZN(U3453) );
  AOI21_X1 U7463 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6514) );
  AOI22_X1 U7464 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6514), .B2(n6513), .ZN(n6515) );
  INV_X1 U7465 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6618) );
  AOI22_X1 U7466 ( .A1(n6516), .A2(n6515), .B1(n6618), .B2(n6519), .ZN(U3468)
         );
  INV_X1 U7467 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6520) );
  NOR2_X1 U7468 ( .A1(n6519), .A2(REIP_REG_1__SCAN_IN), .ZN(n6517) );
  AOI22_X1 U7469 ( .A1(n6520), .A2(n6519), .B1(n6518), .B2(n6517), .ZN(U3469)
         );
  NAND2_X1 U7470 ( .A1(n6540), .A2(W_R_N_REG_SCAN_IN), .ZN(n6521) );
  OAI21_X1 U7471 ( .B1(n6540), .B2(READREQUEST_REG_SCAN_IN), .A(n6521), .ZN(
        U3470) );
  NOR2_X1 U7472 ( .A1(READY_N), .A2(n6522), .ZN(n6530) );
  AOI211_X1 U7473 ( .C1(n6525), .C2(n6530), .A(n6524), .B(n6523), .ZN(n6538)
         );
  INV_X1 U7474 ( .A(n6526), .ZN(n6534) );
  OAI21_X1 U7475 ( .B1(n6528), .B2(n6527), .A(n3496), .ZN(n6531) );
  AOI21_X1 U7476 ( .B1(n6531), .B2(n6530), .A(n6529), .ZN(n6532) );
  AOI21_X1 U7477 ( .B1(n6534), .B2(n6533), .A(n6532), .ZN(n6537) );
  NOR2_X1 U7478 ( .A1(n6538), .A2(n6535), .ZN(n6536) );
  AOI22_X1 U7479 ( .A1(n6539), .A2(n6538), .B1(n6537), .B2(n6536), .ZN(U3472)
         );
  MUX2_X1 U7480 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(M_IO_N_REG_SCAN_IN), .S(
        n6540), .Z(U3473) );
  INV_X1 U7481 ( .A(n6541), .ZN(n6544) );
  INV_X1 U7482 ( .A(n6549), .ZN(n6542) );
  NOR3_X1 U7483 ( .A1(n6550), .A2(n6552), .A3(n6542), .ZN(n6543) );
  AOI21_X1 U7484 ( .B1(n6545), .B2(n6544), .A(n6543), .ZN(n6546) );
  OAI21_X1 U7485 ( .B1(n6548), .B2(n6547), .A(n6546), .ZN(n6554) );
  OAI21_X1 U7486 ( .B1(n6550), .B2(n6549), .A(n6553), .ZN(n6551) );
  AOI22_X1 U7487 ( .A1(n6554), .A2(n6553), .B1(n6552), .B2(n6551), .ZN(n6707)
         );
  AOI22_X1 U7488 ( .A1(n6557), .A2(keyinput42), .B1(n6556), .B2(keyinput27), 
        .ZN(n6555) );
  OAI221_X1 U7489 ( .B1(n6557), .B2(keyinput42), .C1(n6556), .C2(keyinput27), 
        .A(n6555), .ZN(n6567) );
  AOI22_X1 U7490 ( .A1(n6560), .A2(keyinput40), .B1(keyinput59), .B2(n6559), 
        .ZN(n6558) );
  OAI221_X1 U7491 ( .B1(n6560), .B2(keyinput40), .C1(n6559), .C2(keyinput59), 
        .A(n6558), .ZN(n6566) );
  INV_X1 U7492 ( .A(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n6681) );
  AOI22_X1 U7493 ( .A1(n6681), .A2(keyinput5), .B1(n4660), .B2(keyinput56), 
        .ZN(n6561) );
  OAI221_X1 U7494 ( .B1(n6681), .B2(keyinput5), .C1(n4660), .C2(keyinput56), 
        .A(n6561), .ZN(n6565) );
  XNOR2_X1 U7495 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .B(keyinput63), .ZN(
        n6563) );
  XNOR2_X1 U7496 ( .A(INSTQUEUE_REG_13__4__SCAN_IN), .B(keyinput29), .ZN(n6562) );
  NAND2_X1 U7497 ( .A1(n6563), .A2(n6562), .ZN(n6564) );
  NOR4_X1 U7498 ( .A1(n6567), .A2(n6566), .A3(n6565), .A4(n6564), .ZN(n6610)
         );
  INV_X1 U7499 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n6682) );
  AOI22_X1 U7500 ( .A1(n6569), .A2(keyinput4), .B1(n6682), .B2(keyinput32), 
        .ZN(n6568) );
  OAI221_X1 U7501 ( .B1(n6569), .B2(keyinput4), .C1(n6682), .C2(keyinput32), 
        .A(n6568), .ZN(n6582) );
  AOI22_X1 U7502 ( .A1(n6572), .A2(keyinput14), .B1(n6571), .B2(keyinput0), 
        .ZN(n6570) );
  OAI221_X1 U7503 ( .B1(n6572), .B2(keyinput14), .C1(n6571), .C2(keyinput0), 
        .A(n6570), .ZN(n6581) );
  INV_X1 U7504 ( .A(DATAI_19_), .ZN(n6575) );
  AOI22_X1 U7505 ( .A1(n6575), .A2(keyinput7), .B1(n6574), .B2(keyinput18), 
        .ZN(n6573) );
  OAI221_X1 U7506 ( .B1(n6575), .B2(keyinput7), .C1(n6574), .C2(keyinput18), 
        .A(n6573), .ZN(n6580) );
  AOI22_X1 U7507 ( .A1(n6578), .A2(keyinput38), .B1(keyinput23), .B2(n6577), 
        .ZN(n6576) );
  OAI221_X1 U7508 ( .B1(n6578), .B2(keyinput38), .C1(n6577), .C2(keyinput23), 
        .A(n6576), .ZN(n6579) );
  NOR4_X1 U7509 ( .A1(n6582), .A2(n6581), .A3(n6580), .A4(n6579), .ZN(n6609)
         );
  AOI22_X1 U7510 ( .A1(n6585), .A2(keyinput39), .B1(keyinput25), .B2(n6584), 
        .ZN(n6583) );
  OAI221_X1 U7511 ( .B1(n6585), .B2(keyinput39), .C1(n6584), .C2(keyinput25), 
        .A(n6583), .ZN(n6595) );
  INV_X1 U7512 ( .A(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n6587) );
  AOI22_X1 U7513 ( .A1(n6587), .A2(keyinput20), .B1(keyinput34), .B2(n4315), 
        .ZN(n6586) );
  OAI221_X1 U7514 ( .B1(n6587), .B2(keyinput20), .C1(n4315), .C2(keyinput34), 
        .A(n6586), .ZN(n6594) );
  XOR2_X1 U7515 ( .A(n4650), .B(keyinput26), .Z(n6590) );
  XNOR2_X1 U7516 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .B(keyinput15), .ZN(n6589)
         );
  XNOR2_X1 U7517 ( .A(INSTQUEUE_REG_11__6__SCAN_IN), .B(keyinput62), .ZN(n6588) );
  NAND3_X1 U7518 ( .A1(n6590), .A2(n6589), .A3(n6588), .ZN(n6593) );
  XNOR2_X1 U7519 ( .A(n6591), .B(keyinput46), .ZN(n6592) );
  NOR4_X1 U7520 ( .A1(n6595), .A2(n6594), .A3(n6593), .A4(n6592), .ZN(n6608)
         );
  AOI22_X1 U7521 ( .A1(n4330), .A2(keyinput48), .B1(n6597), .B2(keyinput8), 
        .ZN(n6596) );
  OAI221_X1 U7522 ( .B1(n4330), .B2(keyinput48), .C1(n6597), .C2(keyinput8), 
        .A(n6596), .ZN(n6606) );
  AOI22_X1 U7523 ( .A1(n3728), .A2(keyinput36), .B1(n6683), .B2(keyinput16), 
        .ZN(n6598) );
  OAI221_X1 U7524 ( .B1(n3728), .B2(keyinput36), .C1(n6683), .C2(keyinput16), 
        .A(n6598), .ZN(n6605) );
  AOI22_X1 U7525 ( .A1(n4574), .A2(keyinput19), .B1(keyinput52), .B2(n6600), 
        .ZN(n6599) );
  OAI221_X1 U7526 ( .B1(n4574), .B2(keyinput19), .C1(n6600), .C2(keyinput52), 
        .A(n6599), .ZN(n6604) );
  INV_X1 U7527 ( .A(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n6688) );
  AOI22_X1 U7528 ( .A1(n6602), .A2(keyinput10), .B1(n6688), .B2(keyinput24), 
        .ZN(n6601) );
  OAI221_X1 U7529 ( .B1(n6602), .B2(keyinput10), .C1(n6688), .C2(keyinput24), 
        .A(n6601), .ZN(n6603) );
  NOR4_X1 U7530 ( .A1(n6606), .A2(n6605), .A3(n6604), .A4(n6603), .ZN(n6607)
         );
  NAND4_X1 U7531 ( .A1(n6610), .A2(n6609), .A3(n6608), .A4(n6607), .ZN(n6672)
         );
  AOI22_X1 U7532 ( .A1(n5124), .A2(keyinput54), .B1(keyinput22), .B2(n6612), 
        .ZN(n6611) );
  OAI221_X1 U7533 ( .B1(n5124), .B2(keyinput54), .C1(n6612), .C2(keyinput22), 
        .A(n6611), .ZN(n6625) );
  INV_X1 U7534 ( .A(DATAI_18_), .ZN(n6614) );
  AOI22_X1 U7535 ( .A1(n6615), .A2(keyinput55), .B1(keyinput53), .B2(n6614), 
        .ZN(n6613) );
  OAI221_X1 U7536 ( .B1(n6615), .B2(keyinput55), .C1(n6614), .C2(keyinput53), 
        .A(n6613), .ZN(n6624) );
  AOI22_X1 U7537 ( .A1(n6618), .A2(keyinput49), .B1(n6617), .B2(keyinput1), 
        .ZN(n6616) );
  OAI221_X1 U7538 ( .B1(n6618), .B2(keyinput49), .C1(n6617), .C2(keyinput1), 
        .A(n6616), .ZN(n6623) );
  INV_X1 U7539 ( .A(LWORD_REG_4__SCAN_IN), .ZN(n6621) );
  INV_X1 U7540 ( .A(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n6620) );
  AOI22_X1 U7541 ( .A1(n6621), .A2(keyinput58), .B1(n6620), .B2(keyinput57), 
        .ZN(n6619) );
  OAI221_X1 U7542 ( .B1(n6621), .B2(keyinput58), .C1(n6620), .C2(keyinput57), 
        .A(n6619), .ZN(n6622) );
  NOR4_X1 U7543 ( .A1(n6625), .A2(n6624), .A3(n6623), .A4(n6622), .ZN(n6670)
         );
  AOI22_X1 U7544 ( .A1(n6691), .A2(keyinput9), .B1(keyinput61), .B2(n6627), 
        .ZN(n6626) );
  OAI221_X1 U7545 ( .B1(n6691), .B2(keyinput9), .C1(n6627), .C2(keyinput61), 
        .A(n6626), .ZN(n6639) );
  AOI22_X1 U7546 ( .A1(n6629), .A2(keyinput37), .B1(keyinput44), .B2(n3082), 
        .ZN(n6628) );
  OAI221_X1 U7547 ( .B1(n6629), .B2(keyinput37), .C1(n3082), .C2(keyinput44), 
        .A(n6628), .ZN(n6638) );
  AOI22_X1 U7548 ( .A1(n6632), .A2(keyinput13), .B1(keyinput47), .B2(n6631), 
        .ZN(n6630) );
  OAI221_X1 U7549 ( .B1(n6632), .B2(keyinput13), .C1(n6631), .C2(keyinput47), 
        .A(n6630), .ZN(n6637) );
  AOI22_X1 U7550 ( .A1(n6635), .A2(keyinput51), .B1(keyinput30), .B2(n6634), 
        .ZN(n6633) );
  OAI221_X1 U7551 ( .B1(n6635), .B2(keyinput51), .C1(n6634), .C2(keyinput30), 
        .A(n6633), .ZN(n6636) );
  NOR4_X1 U7552 ( .A1(n6639), .A2(n6638), .A3(n6637), .A4(n6636), .ZN(n6669)
         );
  INV_X1 U7553 ( .A(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n6684) );
  AOI22_X1 U7554 ( .A1(n4314), .A2(keyinput43), .B1(n6684), .B2(keyinput41), 
        .ZN(n6640) );
  OAI221_X1 U7555 ( .B1(n4314), .B2(keyinput43), .C1(n6684), .C2(keyinput41), 
        .A(n6640), .ZN(n6652) );
  AOI22_X1 U7556 ( .A1(n6643), .A2(keyinput28), .B1(keyinput6), .B2(n6642), 
        .ZN(n6641) );
  OAI221_X1 U7557 ( .B1(n6643), .B2(keyinput28), .C1(n6642), .C2(keyinput6), 
        .A(n6641), .ZN(n6651) );
  INV_X1 U7558 ( .A(D_C_N_REG_SCAN_IN), .ZN(n6645) );
  AOI22_X1 U7559 ( .A1(n6646), .A2(keyinput35), .B1(n6645), .B2(keyinput33), 
        .ZN(n6644) );
  OAI221_X1 U7560 ( .B1(n6646), .B2(keyinput35), .C1(n6645), .C2(keyinput33), 
        .A(n6644), .ZN(n6650) );
  XOR2_X1 U7561 ( .A(n6673), .B(keyinput60), .Z(n6648) );
  XNOR2_X1 U7562 ( .A(INSTQUEUE_REG_6__3__SCAN_IN), .B(keyinput12), .ZN(n6647)
         );
  NAND2_X1 U7563 ( .A1(n6648), .A2(n6647), .ZN(n6649) );
  NOR4_X1 U7564 ( .A1(n6652), .A2(n6651), .A3(n6650), .A4(n6649), .ZN(n6668)
         );
  INV_X1 U7565 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n6654) );
  AOI22_X1 U7566 ( .A1(n6655), .A2(keyinput45), .B1(n6654), .B2(keyinput2), 
        .ZN(n6653) );
  OAI221_X1 U7567 ( .B1(n6655), .B2(keyinput45), .C1(n6654), .C2(keyinput2), 
        .A(n6653), .ZN(n6666) );
  INV_X1 U7568 ( .A(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n6687) );
  INV_X1 U7569 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6657) );
  AOI22_X1 U7570 ( .A1(n6687), .A2(keyinput50), .B1(keyinput21), .B2(n6657), 
        .ZN(n6656) );
  OAI221_X1 U7571 ( .B1(n6687), .B2(keyinput50), .C1(n6657), .C2(keyinput21), 
        .A(n6656), .ZN(n6665) );
  AOI22_X1 U7572 ( .A1(n6660), .A2(keyinput31), .B1(n6659), .B2(keyinput11), 
        .ZN(n6658) );
  OAI221_X1 U7573 ( .B1(n6660), .B2(keyinput31), .C1(n6659), .C2(keyinput11), 
        .A(n6658), .ZN(n6664) );
  XOR2_X1 U7574 ( .A(n4968), .B(keyinput17), .Z(n6662) );
  XNOR2_X1 U7575 ( .A(INSTQUEUE_REG_1__5__SCAN_IN), .B(keyinput3), .ZN(n6661)
         );
  NAND2_X1 U7576 ( .A1(n6662), .A2(n6661), .ZN(n6663) );
  NOR4_X1 U7577 ( .A1(n6666), .A2(n6665), .A3(n6664), .A4(n6663), .ZN(n6667)
         );
  NAND4_X1 U7578 ( .A1(n6670), .A2(n6669), .A3(n6668), .A4(n6667), .ZN(n6671)
         );
  NOR2_X1 U7579 ( .A1(n6672), .A2(n6671), .ZN(n6705) );
  NOR4_X1 U7580 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(DATAI_6_), .A3(
        DATAI_4_), .A4(CODEFETCH_REG_SCAN_IN), .ZN(n6703) );
  NAND4_X1 U7581 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .A3(DATAO_REG_21__SCAN_IN), .A4(n6673), 
        .ZN(n6676) );
  NAND4_X1 U7582 ( .A1(DATAO_REG_20__SCAN_IN), .A2(DATAO_REG_17__SCAN_IN), 
        .A3(UWORD_REG_6__SCAN_IN), .A4(ADDRESS_REG_4__SCAN_IN), .ZN(n6675) );
  NAND4_X1 U7583 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        ADDRESS_REG_6__SCAN_IN), .A3(NA_N), .A4(DATAWIDTH_REG_14__SCAN_IN), 
        .ZN(n6674) );
  NOR3_X1 U7584 ( .A1(n6676), .A2(n6675), .A3(n6674), .ZN(n6702) );
  NAND4_X1 U7585 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(DATAI_2_), .A3(
        DATAO_REG_18__SCAN_IN), .A4(LWORD_REG_4__SCAN_IN), .ZN(n6680) );
  NAND4_X1 U7586 ( .A1(EBX_REG_13__SCAN_IN), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .A3(EAX_REG_18__SCAN_IN), .A4(DATAI_1_), .ZN(n6679) );
  NAND4_X1 U7587 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        EBX_REG_17__SCAN_IN), .A3(PHYADDRPOINTER_REG_30__SCAN_IN), .A4(
        DATAI_19_), .ZN(n6678) );
  NAND4_X1 U7588 ( .A1(EBX_REG_20__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_29__SCAN_IN), .A3(PHYADDRPOINTER_REG_25__SCAN_IN), 
        .A4(DATAI_10_), .ZN(n6677) );
  NOR4_X1 U7589 ( .A1(n6680), .A2(n6679), .A3(n6678), .A4(n6677), .ZN(n6701)
         );
  NOR4_X1 U7590 ( .A1(D_C_N_REG_SCAN_IN), .A2(INSTQUEUE_REG_4__3__SCAN_IN), 
        .A3(UWORD_REG_14__SCAN_IN), .A4(n6681), .ZN(n6699) );
  NOR4_X1 U7591 ( .A1(EBX_REG_3__SCAN_IN), .A2(ADDRESS_REG_12__SCAN_IN), .A3(
        DATAO_REG_11__SCAN_IN), .A4(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6698) );
  NOR4_X1 U7592 ( .A1(INSTQUEUE_REG_14__5__SCAN_IN), .A2(
        INSTQUEUE_REG_13__7__SCAN_IN), .A3(INSTQUEUE_REG_15__7__SCAN_IN), .A4(
        n6682), .ZN(n6685) );
  AND4_X1 U7593 ( .A1(n6686), .A2(n6685), .A3(n6684), .A4(n6683), .ZN(n6697)
         );
  NAND4_X1 U7594 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(
        INSTQUEUE_REG_5__1__SCAN_IN), .A3(INSTQUEUE_REG_4__2__SCAN_IN), .A4(
        n6687), .ZN(n6695) );
  AND4_X1 U7595 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(
        INSTQUEUE_REG_9__0__SCAN_IN), .A3(INSTQUEUE_REG_11__6__SCAN_IN), .A4(
        INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n6693) );
  NOR4_X1 U7596 ( .A1(EBX_REG_10__SCAN_IN), .A2(EAX_REG_6__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .A4(DATAI_18_), .ZN(n6689) );
  NAND3_X1 U7597 ( .A1(n6689), .A2(n4650), .A3(n6688), .ZN(n6690) );
  NOR2_X1 U7598 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n6690), .ZN(n6692) );
  NAND3_X1 U7599 ( .A1(n6693), .A2(n6692), .A3(n6691), .ZN(n6694) );
  NOR2_X1 U7600 ( .A1(n6695), .A2(n6694), .ZN(n6696) );
  AND4_X1 U7601 ( .A1(n6699), .A2(n6698), .A3(n6697), .A4(n6696), .ZN(n6700)
         );
  NAND4_X1 U7602 ( .A1(n6703), .A2(n6702), .A3(n6701), .A4(n6700), .ZN(n6704)
         );
  XNOR2_X1 U7603 ( .A(n6705), .B(n6704), .ZN(n6706) );
  XNOR2_X1 U7604 ( .A(n6707), .B(n6706), .ZN(U3459) );
  CLKBUF_X2 U4521 ( .A(n4010), .Z(n5835) );
  CLKBUF_X1 U3424 ( .A(n3491), .Z(n4450) );
  NOR2_X1 U3551 ( .A1(n4112), .A2(n3935), .ZN(n4116) );
  CLKBUF_X1 U3604 ( .A(n5097), .Z(n5109) );
  NAND2_X2 U4288 ( .A1(n4059), .A2(n3996), .ZN(n4079) );
  CLKBUF_X1 U4845 ( .A(n3376), .Z(n3769) );
endmodule

