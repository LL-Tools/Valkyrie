

module b20_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, 
        SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, 
        SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, 
        SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, 
        P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n5124, n5125, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11124;

  INV_X4 U5187 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  AOI21_X1 U5188 ( .B1(n8261), .B2(n8260), .A(n8259), .ZN(n11008) );
  INV_X2 U5189 ( .A(n7089), .ZN(n5129) );
  INV_X1 U5190 ( .A(n6928), .ZN(n7086) );
  CLKBUF_X2 U5192 ( .A(n6477), .Z(n5125) );
  CLKBUF_X2 U5193 ( .A(n8666), .Z(n5128) );
  CLKBUF_X1 U5194 ( .A(n5768), .Z(n5369) );
  INV_X1 U5195 ( .A(n9018), .ZN(n9007) );
  INV_X1 U5196 ( .A(n7130), .ZN(n6683) );
  NAND2_X1 U5197 ( .A1(n8888), .A2(n8896), .ZN(n8849) );
  INV_X1 U5198 ( .A(n9709), .ZN(n6153) );
  OAI21_X1 U5199 ( .B1(n6177), .B2(n5349), .A(n6180), .ZN(n6196) );
  NOR2_X2 U5200 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5962) );
  AND4_X1 U5201 ( .A1(n6503), .A2(n6502), .A3(n6501), .A4(n6500), .ZN(n7798)
         );
  INV_X1 U5202 ( .A(n8841), .ZN(n8837) );
  INV_X1 U5203 ( .A(n9151), .ZN(n5535) );
  AOI21_X1 U5204 ( .B1(n10140), .B2(n11107), .A(n5287), .ZN(n6914) );
  CLKBUF_X2 U5205 ( .A(n6916), .Z(n5130) );
  AND2_X1 U5206 ( .A1(n6431), .A2(n6434), .ZN(n6477) );
  XOR2_X1 U5207 ( .A(n9183), .B(n9182), .Z(n5124) );
  OAI211_X2 U5208 ( .C1(n8869), .C2(n8870), .A(n8999), .B(n9004), .ZN(n8871)
         );
  OAI22_X2 U5209 ( .A1(n7457), .A2(n7458), .B1(n6947), .B2(n6946), .ZN(n7754)
         );
  OAI222_X1 U5210 ( .A1(n9376), .A2(n7798), .B1(n9361), .B2(n7486), .C1(n9373), 
        .C2(n7449), .ZN(n7971) );
  NAND2_X2 U5211 ( .A1(n9731), .A2(n9842), .ZN(n9847) );
  AND2_X2 U5212 ( .A1(n6221), .A2(n6220), .ZN(n10445) );
  INV_X1 U5213 ( .A(n8032), .ZN(n7432) );
  NAND2_X2 U5214 ( .A1(n5242), .A2(n6474), .ZN(n8032) );
  BUF_X8 U5215 ( .A(n6475), .Z(n6839) );
  NAND2_X2 U5216 ( .A1(n9628), .A2(n7003), .ZN(n9522) );
  AOI22_X2 U5217 ( .A1(n7438), .A2(n7437), .B1(n6942), .B2(n6941), .ZN(n7457)
         );
  NAND2_X1 U5218 ( .A1(n7398), .A2(n7402), .ZN(n7438) );
  OAI22_X2 U5219 ( .A1(n10185), .A2(n6249), .B1(n7080), .B2(n10441), .ZN(
        n10170) );
  INV_X2 U5220 ( .A(n6324), .ZN(n6328) );
  NAND2_X2 U5221 ( .A1(n6442), .A2(n6441), .ZN(n6837) );
  XNOR2_X2 U5222 ( .A(n5262), .B(n6444), .ZN(n6838) );
  AOI21_X2 U5223 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n9081), .A(n9082), .ZN(
        n8582) );
  BUF_X2 U5224 ( .A(n7238), .Z(n5127) );
  AOI21_X2 U5225 ( .B1(n8183), .B2(n8173), .A(n8172), .ZN(n8261) );
  AND2_X1 U5226 ( .A1(n5405), .A2(n5404), .ZN(n10150) );
  XNOR2_X1 U5227 ( .A(n5380), .B(n6835), .ZN(n6846) );
  CLKBUF_X1 U5228 ( .A(n9530), .Z(n9612) );
  AND2_X1 U5229 ( .A1(n9619), .A2(n5194), .ZN(n9561) );
  INV_X1 U5230 ( .A(n10445), .ZN(n10201) );
  AOI22_X1 U5231 ( .A1(n5270), .A2(n5698), .B1(n7907), .B2(n6340), .ZN(n8099)
         );
  AND2_X1 U5232 ( .A1(n5646), .A2(n5645), .ZN(n8232) );
  OAI21_X1 U5233 ( .B1(n8897), .B2(n5375), .A(n8852), .ZN(n5374) );
  AND2_X1 U5234 ( .A1(n8909), .A2(n8905), .ZN(n8852) );
  NAND2_X1 U5235 ( .A1(n8127), .A2(n7806), .ZN(n8909) );
  INV_X2 U5236 ( .A(n7798), .ZN(n9048) );
  INV_X2 U5237 ( .A(n7839), .ZN(n9049) );
  INV_X2 U5238 ( .A(n8127), .ZN(n9047) );
  INV_X2 U5239 ( .A(n7940), .ZN(n10002) );
  INV_X1 U5240 ( .A(n7486), .ZN(n9050) );
  AND4_X1 U5241 ( .A1(n6490), .A2(n6489), .A3(n6488), .A4(n6487), .ZN(n7839)
         );
  NAND2_X1 U5242 ( .A1(n6921), .A2(n6920), .ZN(n6928) );
  INV_X1 U5243 ( .A(n7485), .ZN(n7976) );
  XNOR2_X1 U5244 ( .A(n6806), .B(P2_IR_REG_21__SCAN_IN), .ZN(n7476) );
  NAND2_X1 U5245 ( .A1(n6328), .A2(n7848), .ZN(n6917) );
  BUF_X2 U5246 ( .A(n5971), .Z(n5131) );
  CLKBUF_X2 U5247 ( .A(n5971), .Z(n5132) );
  AND2_X1 U5248 ( .A1(n7848), .A2(n6916), .ZN(n9758) );
  AND3_X2 U5249 ( .A1(n5967), .A2(n5966), .A3(n5965), .ZN(n11034) );
  AND2_X1 U5250 ( .A1(n8634), .A2(n5871), .ZN(n5971) );
  INV_X1 U5251 ( .A(n8541), .ZN(n5871) );
  XNOR2_X1 U5252 ( .A(n6802), .B(P2_IR_REG_19__SCAN_IN), .ZN(n9151) );
  NAND2_X2 U5253 ( .A1(n5857), .A2(n5856), .ZN(n5889) );
  NAND2_X1 U5254 ( .A1(n5275), .A2(n5271), .ZN(n8634) );
  OAI21_X1 U5255 ( .B1(n6113), .B2(n5652), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6129) );
  NAND2_X1 U5256 ( .A1(n6360), .A2(n5852), .ZN(n6370) );
  AND3_X2 U5257 ( .A1(n5846), .A2(n5845), .A3(n5710), .ZN(n6360) );
  NAND2_X1 U5258 ( .A1(n6457), .A2(n6456), .ZN(n8666) );
  INV_X1 U5259 ( .A(n5927), .ZN(n5845) );
  NAND2_X1 U5260 ( .A1(n10150), .A2(n5288), .ZN(n5287) );
  AND2_X1 U5261 ( .A1(n9025), .A2(n6897), .ZN(n5339) );
  OAI21_X1 U5262 ( .B1(n9674), .B2(n9673), .A(n9672), .ZN(n9677) );
  NAND2_X1 U5263 ( .A1(n8747), .A2(n8748), .ZN(n8810) );
  OAI21_X1 U5264 ( .B1(n6401), .B2(n9799), .A(n6400), .ZN(n8677) );
  NAND2_X1 U5265 ( .A1(n5606), .A2(n5610), .ZN(n9577) );
  NAND2_X1 U5266 ( .A1(n5614), .A2(n9610), .ZN(n9609) );
  OAI21_X1 U5267 ( .B1(n10199), .B2(n6230), .A(n6231), .ZN(n10185) );
  AND2_X1 U5268 ( .A1(n10144), .A2(n5212), .ZN(n5288) );
  NAND2_X1 U5269 ( .A1(n5284), .A2(n6215), .ZN(n10199) );
  AOI211_X1 U5270 ( .C1(n8673), .C2(n11065), .A(n8672), .B(n8671), .ZN(n8676)
         );
  NOR2_X1 U5271 ( .A1(n10134), .A2(n10135), .ZN(n5394) );
  NAND2_X1 U5272 ( .A1(n10235), .A2(n10234), .ZN(n5708) );
  AOI21_X1 U5273 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n9118), .A(n9119), .ZN(
        n8585) );
  OAI21_X1 U5274 ( .B1(n8507), .B2(n8467), .A(n8466), .ZN(n8517) );
  OAI21_X1 U5275 ( .B1(n8103), .B2(n5424), .A(n5422), .ZN(n6341) );
  OAI21_X1 U5276 ( .B1(n8089), .B2(n8088), .A(n8087), .ZN(n8091) );
  NAND2_X1 U5277 ( .A1(n7880), .A2(n9781), .ZN(n7879) );
  NAND2_X1 U5278 ( .A1(n5918), .A2(n5917), .ZN(n9527) );
  NAND2_X1 U5279 ( .A1(n6101), .A2(n6100), .ZN(n8207) );
  NOR2_X1 U5280 ( .A1(n7993), .A2(n5428), .ZN(n8166) );
  NAND2_X1 U5281 ( .A1(n5343), .A2(n5341), .ZN(n5809) );
  NAND2_X1 U5282 ( .A1(n5935), .A2(n5934), .ZN(n9547) );
  NAND2_X2 U5283 ( .A1(n7592), .A2(n9380), .ZN(n9377) );
  NAND2_X1 U5284 ( .A1(n7283), .A2(n7282), .ZN(n7625) );
  OR2_X1 U5285 ( .A1(n7281), .A2(n7280), .ZN(n7283) );
  INV_X8 U5286 ( .A(n8678), .ZN(n8694) );
  OR2_X1 U5287 ( .A1(n8851), .A2(n7429), .ZN(n7430) );
  NAND2_X1 U5288 ( .A1(n7432), .A2(n9051), .ZN(n8883) );
  NAND2_X1 U5289 ( .A1(n7240), .A2(n7271), .ZN(n7279) );
  CLKBUF_X3 U5290 ( .A(n6928), .Z(n8706) );
  OR2_X1 U5291 ( .A1(n10978), .A2(n7239), .ZN(n7240) );
  AND4_X1 U5292 ( .A1(n6000), .A2(n5999), .A3(n5998), .A4(n5997), .ZN(n7940)
         );
  AND2_X2 U5293 ( .A1(n7476), .A2(n9028), .ZN(n9018) );
  NAND2_X1 U5294 ( .A1(n6327), .A2(n5130), .ZN(n6921) );
  AND4_X1 U5295 ( .A1(n5975), .A2(n5974), .A3(n5973), .A4(n5972), .ZN(n7568)
         );
  INV_X2 U5297 ( .A(n6492), .ZN(n8838) );
  NAND2_X1 U5298 ( .A1(n6430), .A2(n6429), .ZN(n9515) );
  NAND2_X1 U5299 ( .A1(n6319), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6388) );
  NAND2_X1 U5300 ( .A1(n6386), .A2(n6385), .ZN(n7126) );
  AND2_X1 U5301 ( .A1(n5872), .A2(n5871), .ZN(n5980) );
  MUX2_X1 U5302 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6428), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n6430) );
  NOR2_X1 U5303 ( .A1(n8417), .A2(n8244), .ZN(n6385) );
  INV_X2 U5304 ( .A(n6013), .ZN(n9708) );
  NAND2_X1 U5305 ( .A1(n6365), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6320) );
  NAND2_X1 U5306 ( .A1(n5889), .A2(n8604), .ZN(n6013) );
  NAND2_X1 U5307 ( .A1(n10474), .A2(n5870), .ZN(n8541) );
  NAND2_X1 U5308 ( .A1(n6443), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5262) );
  NAND2_X1 U5309 ( .A1(n5869), .A2(n5868), .ZN(n5870) );
  NAND2_X1 U5310 ( .A1(n10474), .A2(n5274), .ZN(n5271) );
  AND2_X1 U5311 ( .A1(n5272), .A2(n5203), .ZN(n5275) );
  XNOR2_X1 U5312 ( .A(n6504), .B(P2_IR_REG_4__SCAN_IN), .ZN(n7238) );
  OR2_X1 U5313 ( .A1(n6362), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n6368) );
  INV_X2 U5314 ( .A(n8609), .ZN(n8667) );
  AND2_X1 U5315 ( .A1(n11124), .A2(n6424), .ZN(n6886) );
  XNOR2_X1 U5316 ( .A(n6491), .B(n6558), .ZN(n8623) );
  AND4_X1 U5317 ( .A1(n5167), .A2(n6666), .A3(n6667), .A4(n6423), .ZN(n6424)
         );
  CLKBUF_X1 U5318 ( .A(n6453), .Z(n7205) );
  NAND3_X1 U5319 ( .A1(n5683), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n5685) );
  NAND3_X1 U5320 ( .A1(n5679), .A2(n5678), .A3(n5677), .ZN(n5686) );
  AND2_X1 U5321 ( .A1(n6559), .A2(n5555), .ZN(n5554) );
  AND2_X1 U5322 ( .A1(n5556), .A2(n6537), .ZN(n6560) );
  AND2_X1 U5323 ( .A1(n6422), .A2(n6421), .ZN(n6666) );
  AND4_X1 U5324 ( .A1(n5844), .A2(n5843), .A3(n5842), .A4(n5841), .ZN(n5846)
         );
  NOR2_X1 U5325 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n5616) );
  NOR2_X1 U5326 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n6318) );
  INV_X1 U5327 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n10835) );
  INV_X4 U5328 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U5329 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6804) );
  INV_X1 U5330 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5679) );
  NOR2_X1 U5331 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5841) );
  NOR2_X1 U5332 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5842) );
  NOR2_X1 U5333 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5843) );
  INV_X1 U5334 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n10830) );
  NOR2_X1 U5335 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n5861) );
  INV_X1 U5336 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6387) );
  NOR2_X2 U5337 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6453) );
  INV_X1 U5338 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6592) );
  NOR2_X1 U5339 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n5556) );
  NOR2_X1 U5340 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n6559) );
  NOR2_X1 U5341 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n6422) );
  NOR2_X1 U5342 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n6421) );
  NAND2_X2 U5343 ( .A1(n5384), .A2(n6830), .ZN(n9245) );
  NAND4_X2 U5344 ( .A1(n5957), .A2(n5956), .A3(n5955), .A4(n5954), .ZN(n6332)
         );
  OAI211_X2 U5345 ( .C1(n5636), .C2(n5628), .A(n5627), .B(n5625), .ZN(n8021)
         );
  NOR2_X1 U5346 ( .A1(n5160), .A2(n5629), .ZN(n5628) );
  NOR2_X2 U5347 ( .A1(n8718), .A2(n10155), .ZN(n6403) );
  OAI22_X2 U5348 ( .A1(n10952), .A2(n10953), .B1(n10936), .B2(n7195), .ZN(
        n10973) );
  AOI211_X2 U5349 ( .C1(n8674), .C2(n10411), .A(n6404), .B(n8673), .ZN(n6405)
         );
  AOI21_X4 U5350 ( .B1(n8295), .B2(n8294), .A(n6975), .ZN(n9541) );
  OAI22_X2 U5351 ( .A1(n8232), .A2(n8231), .B1(n6968), .B2(n6967), .ZN(n8295)
         );
  XNOR2_X1 U5352 ( .A(n6151), .B(n6150), .ZN(n6916) );
  OAI22_X1 U5353 ( .A1(n5133), .A2(n9018), .B1(n5138), .B2(n9007), .ZN(n5320)
         );
  OR2_X1 U5354 ( .A1(n8845), .A2(n8844), .ZN(n8877) );
  AND2_X1 U5355 ( .A1(n5344), .A2(n5342), .ZN(n5341) );
  INV_X1 U5356 ( .A(n5914), .ZN(n5342) );
  OR2_X1 U5357 ( .A1(n6893), .A2(n9179), .ZN(n8875) );
  OR2_X1 U5358 ( .A1(n9196), .A2(n9204), .ZN(n9004) );
  AOI21_X1 U5359 ( .B1(n5136), .B2(n5722), .A(n5183), .ZN(n5718) );
  INV_X1 U5360 ( .A(n6642), .ZN(n5722) );
  INV_X1 U5361 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5259) );
  AOI21_X1 U5362 ( .B1(n5283), .B2(n9770), .A(n5282), .ZN(n5281) );
  INV_X1 U5363 ( .A(n10270), .ZN(n5282) );
  NAND2_X1 U5364 ( .A1(n5840), .A2(n5839), .ZN(n6177) );
  NOR2_X1 U5365 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5710) );
  NAND2_X1 U5366 ( .A1(n7625), .A2(n7624), .ZN(n7851) );
  AOI21_X1 U5367 ( .B1(n9178), .B2(n6794), .A(n5241), .ZN(n5240) );
  AND2_X1 U5368 ( .A1(n8698), .A2(n9033), .ZN(n5241) );
  INV_X1 U5369 ( .A(n5391), .ZN(n6439) );
  INV_X1 U5370 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6529) );
  NAND2_X1 U5371 ( .A1(n5620), .A2(n5185), .ZN(n5619) );
  INV_X1 U5372 ( .A(n5621), .ZN(n5620) );
  OR2_X1 U5373 ( .A1(n7627), .A2(n8212), .ZN(n5237) );
  AND2_X1 U5374 ( .A1(n5302), .A2(n5298), .ZN(n5297) );
  NAND2_X1 U5375 ( .A1(n8950), .A2(n9018), .ZN(n5298) );
  AND2_X1 U5376 ( .A1(n9295), .A2(n5313), .ZN(n5312) );
  AOI21_X1 U5377 ( .B1(n5320), .B2(n8965), .A(n5314), .ZN(n5313) );
  NAND2_X1 U5378 ( .A1(n5318), .A2(n5319), .ZN(n5314) );
  AND2_X1 U5379 ( .A1(n8973), .A2(n9280), .ZN(n5321) );
  OR2_X1 U5380 ( .A1(n6574), .A2(n6573), .ZN(n6576) );
  INV_X1 U5381 ( .A(SI_17_), .ZN(n10690) );
  AND2_X1 U5382 ( .A1(n5348), .A2(n5803), .ZN(n5347) );
  NAND2_X1 U5383 ( .A1(n5802), .A2(n5801), .ZN(n5348) );
  NOR2_X1 U5384 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(n6697), .ZN(n6708) );
  AND2_X1 U5385 ( .A1(n8519), .A2(n5161), .ZN(n5519) );
  CLKBUF_X1 U5386 ( .A(n5125), .Z(n6728) );
  INV_X1 U5387 ( .A(n9515), .ZN(n6434) );
  NAND2_X1 U5388 ( .A1(n10964), .A2(n7209), .ZN(n7229) );
  NOR2_X1 U5389 ( .A1(n7996), .A2(n5228), .ZN(n8182) );
  AND2_X1 U5390 ( .A1(n7997), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5228) );
  OR2_X1 U5391 ( .A1(n8685), .A2(n9225), .ZN(n8997) );
  OR2_X1 U5392 ( .A1(n9418), .A2(n9257), .ZN(n8979) );
  OR2_X1 U5393 ( .A1(n9433), .A2(n8765), .ZN(n8970) );
  OR2_X1 U5394 ( .A1(n9441), .A2(n9359), .ZN(n9308) );
  OR2_X1 U5395 ( .A1(n8321), .A2(n8390), .ZN(n8920) );
  NAND2_X1 U5396 ( .A1(n7466), .A2(n8032), .ZN(n8886) );
  NAND2_X1 U5397 ( .A1(n5135), .A2(n5170), .ZN(n5255) );
  NAND2_X1 U5398 ( .A1(n6803), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6807) );
  INV_X1 U5399 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6801) );
  AND2_X1 U5400 ( .A1(n9785), .A2(n9891), .ZN(n5425) );
  INV_X1 U5401 ( .A(n8199), .ZN(n5707) );
  XNOR2_X1 U5402 ( .A(n8597), .B(n8596), .ZN(n8599) );
  NAND2_X1 U5403 ( .A1(n5651), .A2(n6318), .ZN(n5650) );
  INV_X1 U5404 ( .A(n5652), .ZN(n5651) );
  AND2_X1 U5405 ( .A1(n5833), .A2(n5832), .ZN(n5834) );
  OR2_X1 U5406 ( .A1(n6147), .A2(n6145), .ZN(n5833) );
  AOI21_X1 U5407 ( .B1(n5675), .B2(n5813), .A(n5674), .ZN(n5672) );
  INV_X1 U5408 ( .A(n5818), .ZN(n5674) );
  INV_X1 U5409 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5890) );
  NAND2_X1 U5410 ( .A1(n5818), .A2(n5817), .ZN(n5887) );
  OAI21_X1 U5411 ( .B1(n6072), .B2(n6071), .A(n5799), .ZN(n6078) );
  AOI22_X1 U5412 ( .A1(n8755), .A2(n8754), .B1(n9325), .B2(n8639), .ZN(n8761)
         );
  AND2_X1 U5413 ( .A1(n8630), .A2(n9515), .ZN(n6476) );
  MUX2_X1 U5414 ( .A(n8881), .B(n8880), .S(n7476), .Z(n9025) );
  AND2_X1 U5415 ( .A1(n5735), .A2(n5230), .ZN(n5390) );
  AND2_X1 U5416 ( .A1(n6444), .A2(n6888), .ZN(n5230) );
  NAND2_X1 U5417 ( .A1(n5505), .A2(n7231), .ZN(n7233) );
  NAND2_X1 U5418 ( .A1(n5226), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5235) );
  INV_X1 U5419 ( .A(n7994), .ZN(n5226) );
  NAND2_X1 U5420 ( .A1(n5439), .A2(n5438), .ZN(n5437) );
  INV_X1 U5421 ( .A(n8169), .ZN(n5438) );
  NAND2_X1 U5422 ( .A1(n5239), .A2(n5238), .ZN(n5233) );
  NAND2_X1 U5423 ( .A1(n9118), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5238) );
  AND2_X1 U5424 ( .A1(n6834), .A2(n8872), .ZN(n9182) );
  NAND2_X1 U5425 ( .A1(n6771), .A2(n8686), .ZN(n9188) );
  AOI21_X1 U5426 ( .B1(n5267), .B2(n5165), .A(n5263), .ZN(n5711) );
  NAND2_X1 U5427 ( .A1(n5245), .A2(n5244), .ZN(n5723) );
  NOR2_X1 U5428 ( .A1(n5248), .A2(n5207), .ZN(n5244) );
  NAND2_X1 U5429 ( .A1(n9356), .A2(n5249), .ZN(n5245) );
  AND2_X1 U5430 ( .A1(n5136), .A2(n6823), .ZN(n5249) );
  OR2_X1 U5431 ( .A1(n6595), .A2(n5147), .ZN(n5731) );
  NAND2_X1 U5432 ( .A1(n5733), .A2(n5732), .ZN(n8367) );
  NOR2_X1 U5433 ( .A1(n8942), .A2(n5147), .ZN(n5732) );
  NAND2_X1 U5434 ( .A1(n6429), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5725) );
  NAND2_X1 U5435 ( .A1(n6439), .A2(n6426), .ZN(n6441) );
  AND2_X1 U5436 ( .A1(n9552), .A2(n5205), .ZN(n5617) );
  INV_X1 U5437 ( .A(n7848), .ZN(n9986) );
  AND2_X1 U5438 ( .A1(n9974), .A2(n9975), .ZN(n9972) );
  NAND2_X1 U5439 ( .A1(n6399), .A2(n6300), .ZN(n6400) );
  NAND2_X1 U5440 ( .A1(n5277), .A2(n5276), .ZN(n6176) );
  AOI21_X1 U5441 ( .B1(n5278), .B2(n5280), .A(n9936), .ZN(n5276) );
  OR2_X1 U5442 ( .A1(n8299), .A2(n9997), .ZN(n6062) );
  OR2_X1 U5443 ( .A1(n10300), .A2(n5130), .ZN(n7110) );
  NAND2_X1 U5444 ( .A1(n6351), .A2(n5854), .ZN(n5857) );
  AND2_X1 U5445 ( .A1(n5744), .A2(n5860), .ZN(n5866) );
  INV_X1 U5446 ( .A(n9478), .ZN(n8698) );
  XNOR2_X1 U5447 ( .A(n7851), .B(n7626), .ZN(n7627) );
  AND2_X1 U5448 ( .A1(n5430), .A2(n5429), .ZN(n7993) );
  INV_X1 U5449 ( .A(n7855), .ZN(n5429) );
  AOI21_X1 U5450 ( .B1(n6846), .B2(n8385), .A(n6844), .ZN(n5268) );
  OAI21_X1 U5451 ( .B1(n6959), .B2(n8134), .A(n5647), .ZN(n5646) );
  NAND2_X1 U5452 ( .A1(n6959), .A2(n8134), .ZN(n5645) );
  INV_X1 U5453 ( .A(n8135), .ZN(n5647) );
  XNOR2_X1 U5454 ( .A(n5394), .B(n10127), .ZN(n10310) );
  NAND2_X1 U5455 ( .A1(n10508), .A2(n10684), .ZN(n5590) );
  INV_X1 U5456 ( .A(SI_25_), .ZN(n10675) );
  NOR2_X1 U5457 ( .A1(n10689), .A2(n5445), .ZN(n5444) );
  AND2_X1 U5458 ( .A1(n10690), .A2(keyinput_143), .ZN(n5445) );
  NAND2_X1 U5459 ( .A1(n5332), .A2(n5331), .ZN(n8929) );
  OAI21_X1 U5460 ( .B1(n10719), .B2(n5483), .A(n5482), .ZN(n5481) );
  NAND2_X1 U5461 ( .A1(n5485), .A2(n5484), .ZN(n5483) );
  INV_X1 U5462 ( .A(n10721), .ZN(n5482) );
  NOR2_X1 U5463 ( .A1(n10718), .A2(n10717), .ZN(n10719) );
  XNOR2_X1 U5464 ( .A(n10722), .B(n5480), .ZN(n5479) );
  INV_X1 U5465 ( .A(keyinput_164), .ZN(n5480) );
  NAND2_X1 U5466 ( .A1(n5478), .A2(n5477), .ZN(n5476) );
  NAND2_X1 U5467 ( .A1(keyinput_165), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5477)
         );
  NAND2_X1 U5468 ( .A1(n10724), .A2(n10723), .ZN(n5478) );
  NAND2_X1 U5469 ( .A1(n8914), .A2(n9018), .ZN(n5329) );
  INV_X1 U5470 ( .A(n8937), .ZN(n5327) );
  AOI21_X1 U5471 ( .B1(n5568), .B2(n5567), .A(n5564), .ZN(n10572) );
  INV_X1 U5472 ( .A(n10557), .ZN(n5567) );
  NAND2_X1 U5473 ( .A1(n5566), .A2(n5565), .ZN(n5564) );
  NAND2_X1 U5474 ( .A1(n5569), .A2(n10558), .ZN(n5568) );
  OAI22_X1 U5475 ( .A1(n10760), .A2(n10574), .B1(P2_DATAO_REG_30__SCAN_IN), 
        .B2(keyinput_66), .ZN(n5563) );
  AOI21_X1 U5476 ( .B1(n5468), .B2(n10736), .A(n5465), .ZN(n5464) );
  INV_X1 U5477 ( .A(n10738), .ZN(n5465) );
  INV_X1 U5478 ( .A(keyinput_177), .ZN(n5467) );
  NAND2_X1 U5479 ( .A1(n10737), .A2(n5468), .ZN(n5466) );
  INV_X1 U5480 ( .A(n5297), .ZN(n5296) );
  NAND2_X1 U5481 ( .A1(n5297), .A2(n5294), .ZN(n5293) );
  INV_X1 U5482 ( .A(n8950), .ZN(n5294) );
  NAND2_X1 U5483 ( .A1(n5291), .A2(n5297), .ZN(n5300) );
  OR2_X1 U5484 ( .A1(n8944), .A2(n5301), .ZN(n5299) );
  NAND2_X1 U5485 ( .A1(n5302), .A2(n9018), .ZN(n5301) );
  NAND2_X1 U5486 ( .A1(n5312), .A2(n5164), .ZN(n5309) );
  INV_X1 U5487 ( .A(n5320), .ZN(n5317) );
  NAND2_X1 U5488 ( .A1(n5189), .A2(n9018), .ZN(n5315) );
  OR2_X1 U5489 ( .A1(n8969), .A2(n5311), .ZN(n5310) );
  INV_X1 U5490 ( .A(n5312), .ZN(n5311) );
  INV_X1 U5491 ( .A(n10778), .ZN(n5461) );
  NAND2_X1 U5492 ( .A1(n5602), .A2(n5600), .ZN(n10589) );
  NOR2_X1 U5493 ( .A1(n10588), .A2(n5601), .ZN(n5600) );
  XNOR2_X1 U5494 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput_81), .ZN(n5601)
         );
  AOI211_X1 U5495 ( .C1(n10772), .C2(n5459), .A(n5457), .B(n5218), .ZN(n10787)
         );
  NAND2_X1 U5496 ( .A1(n9280), .A2(n6703), .ZN(n5730) );
  NOR2_X1 U5497 ( .A1(n10192), .A2(n10201), .ZN(n5399) );
  INV_X1 U5498 ( .A(n5812), .ZN(n5676) );
  INV_X1 U5499 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5683) );
  INV_X1 U5500 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5678) );
  INV_X1 U5501 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5677) );
  INV_X1 U5502 ( .A(n8692), .ZN(n5530) );
  NAND2_X1 U5503 ( .A1(n7478), .A2(n7582), .ZN(n7484) );
  NAND2_X1 U5504 ( .A1(n8401), .A2(n8402), .ZN(n5549) );
  NAND2_X1 U5505 ( .A1(n8653), .A2(n9266), .ZN(n8654) );
  OAI22_X1 U5506 ( .A1(n5383), .A2(n5382), .B1(n9020), .B2(n8875), .ZN(n5381)
         );
  NAND2_X1 U5507 ( .A1(n9016), .A2(n8872), .ZN(n5382) );
  AOI21_X1 U5508 ( .B1(n9022), .B2(n9021), .A(n9020), .ZN(n9023) );
  NAND2_X1 U5509 ( .A1(n7233), .A2(n7232), .ZN(n7234) );
  AND2_X1 U5510 ( .A1(n7639), .A2(n7638), .ZN(n7866) );
  NAND2_X1 U5511 ( .A1(n5500), .A2(n5499), .ZN(n5498) );
  NAND2_X1 U5512 ( .A1(n8577), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5499) );
  NOR2_X1 U5513 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n6667) );
  INV_X1 U5514 ( .A(n8992), .ZN(n5663) );
  AOI21_X1 U5515 ( .B1(n5662), .B2(n9226), .A(n5660), .ZN(n5659) );
  INV_X1 U5516 ( .A(n8996), .ZN(n5660) );
  NAND2_X1 U5517 ( .A1(n9290), .A2(n5265), .ZN(n5267) );
  NOR2_X1 U5518 ( .A1(n5729), .A2(n5266), .ZN(n5265) );
  INV_X1 U5519 ( .A(n6693), .ZN(n5266) );
  NOR2_X1 U5520 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(n6716), .ZN(n6724) );
  NAND2_X1 U5521 ( .A1(n6687), .A2(n10729), .ZN(n6697) );
  NAND2_X1 U5522 ( .A1(n9311), .A2(n9330), .ZN(n5687) );
  OR2_X1 U5523 ( .A1(n9462), .A2(n9374), .ZN(n8946) );
  OR2_X1 U5524 ( .A1(n8344), .A2(n8402), .ZN(n8938) );
  AND2_X1 U5525 ( .A1(n5139), .A2(n6521), .ZN(n5251) );
  NAND2_X1 U5526 ( .A1(n6476), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n6463) );
  OR2_X1 U5527 ( .A1(n7144), .A2(n6872), .ZN(n6902) );
  OR2_X1 U5528 ( .A1(n7838), .A2(n8897), .ZN(n5734) );
  INV_X1 U5529 ( .A(n6614), .ZN(n5551) );
  AND2_X1 U5530 ( .A1(n6917), .A2(n7126), .ZN(n6920) );
  AOI21_X1 U5531 ( .B1(n6943), .B2(n11024), .A(n6924), .ZN(n6929) );
  AND2_X1 U5532 ( .A1(n7089), .A2(n10005), .ZN(n6924) );
  INV_X1 U5533 ( .A(n8704), .ZN(n7097) );
  NOR2_X1 U5534 ( .A1(n5452), .A2(n5448), .ZN(n5447) );
  OAI21_X1 U5535 ( .B1(n5449), .B2(n5448), .A(n5221), .ZN(n5446) );
  OR2_X1 U5536 ( .A1(n10253), .A2(n10273), .ZN(n9939) );
  NAND2_X1 U5537 ( .A1(n5875), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6187) );
  NOR2_X1 U5538 ( .A1(n8530), .A2(n10385), .ZN(n5402) );
  OR2_X1 U5539 ( .A1(n10398), .A2(n10389), .ZN(n9914) );
  NAND2_X1 U5540 ( .A1(n6104), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5908) );
  INV_X1 U5541 ( .A(n9869), .ZN(n5415) );
  OAI21_X1 U5542 ( .B1(n7884), .B2(n5415), .A(n9879), .ZN(n5414) );
  NAND2_X1 U5543 ( .A1(n5700), .A2(n9654), .ZN(n5699) );
  OR2_X1 U5544 ( .A1(n6055), .A2(n6054), .ZN(n6057) );
  NAND2_X1 U5545 ( .A1(n9836), .A2(n9834), .ZN(n7549) );
  NAND2_X1 U5546 ( .A1(n5360), .A2(n5358), .ZN(n6303) );
  AOI21_X1 U5547 ( .B1(n5362), .B2(n5364), .A(n5359), .ZN(n5358) );
  INV_X1 U5548 ( .A(n6290), .ZN(n5359) );
  AND2_X1 U5549 ( .A1(n6290), .A2(n6276), .ZN(n6288) );
  NAND2_X1 U5550 ( .A1(n6251), .A2(n6250), .ZN(n6255) );
  INV_X1 U5551 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5847) );
  INV_X1 U5552 ( .A(n6178), .ZN(n5349) );
  AND2_X1 U5553 ( .A1(n5839), .A2(n5838), .ZN(n6163) );
  OR2_X1 U5554 ( .A1(n5831), .A2(n5830), .ZN(n6145) );
  AND2_X1 U5555 ( .A1(n6123), .A2(n6125), .ZN(n5830) );
  INV_X1 U5556 ( .A(n6122), .ZN(n5670) );
  NOR2_X1 U5557 ( .A1(n5671), .A2(n5667), .ZN(n5666) );
  INV_X1 U5558 ( .A(n5808), .ZN(n5667) );
  INV_X1 U5559 ( .A(n5668), .ZN(n6144) );
  AOI21_X1 U5560 ( .B1(n5895), .B2(n5675), .A(n5671), .ZN(n5668) );
  XNOR2_X1 U5561 ( .A(n5800), .B(n10664), .ZN(n6077) );
  INV_X1 U5562 ( .A(n5353), .ZN(n5352) );
  NAND2_X1 U5563 ( .A1(n5369), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5367) );
  NAND2_X1 U5564 ( .A1(n8517), .A2(n8516), .ZN(n5520) );
  XNOR2_X1 U5565 ( .A(n8032), .B(n7484), .ZN(n7479) );
  NOR2_X1 U5566 ( .A1(n7542), .A2(n7593), .ZN(n7481) );
  OR2_X1 U5567 ( .A1(n5546), .A2(n5543), .ZN(n5542) );
  INV_X1 U5568 ( .A(n5549), .ZN(n5543) );
  AND2_X1 U5569 ( .A1(n8403), .A2(n5159), .ZN(n5546) );
  OR2_X1 U5570 ( .A1(n8656), .A2(n8655), .ZN(n8769) );
  NAND2_X1 U5571 ( .A1(n8732), .A2(n8731), .ZN(n5537) );
  OR2_X1 U5572 ( .A1(n8330), .A2(n9042), .ZN(n5548) );
  NAND2_X1 U5573 ( .A1(n8221), .A2(n5743), .ZN(n8331) );
  OR2_X1 U5574 ( .A1(n6754), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6765) );
  NAND2_X1 U5575 ( .A1(n5520), .A2(n5519), .ZN(n8822) );
  NAND2_X1 U5576 ( .A1(n6851), .A2(n5735), .ZN(n6443) );
  AND4_X1 U5577 ( .A1(n6438), .A2(n6437), .A3(n6436), .A4(n6435), .ZN(n8127)
         );
  OAI21_X1 U5578 ( .B1(n5128), .B2(n7475), .A(n5225), .ZN(n10959) );
  NAND2_X1 U5579 ( .A1(n5128), .A2(n7475), .ZN(n5225) );
  OAI21_X1 U5580 ( .B1(n5128), .B2(n7982), .A(n5494), .ZN(n10966) );
  NAND2_X1 U5581 ( .A1(n5128), .A2(n7982), .ZN(n5494) );
  NAND2_X1 U5582 ( .A1(n7200), .A2(n8623), .ZN(n5435) );
  NAND2_X1 U5583 ( .A1(n7228), .A2(n5175), .ZN(n5505) );
  XNOR2_X1 U5584 ( .A(n7866), .B(n7867), .ZN(n7640) );
  NOR2_X1 U5585 ( .A1(n7640), .A2(n7628), .ZN(n7868) );
  XNOR2_X1 U5586 ( .A(n8182), .B(n8183), .ZN(n7998) );
  XNOR2_X1 U5587 ( .A(n5234), .B(n8271), .ZN(n11003) );
  NAND2_X1 U5588 ( .A1(n5437), .A2(n5436), .ZN(n5234) );
  NAND2_X1 U5589 ( .A1(n8269), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5436) );
  NOR2_X1 U5590 ( .A1(n11004), .A2(n11003), .ZN(n11002) );
  NOR2_X1 U5591 ( .A1(n10999), .A2(n8272), .ZN(n8277) );
  OR2_X1 U5592 ( .A1(n8277), .A2(n8276), .ZN(n5500) );
  XNOR2_X1 U5593 ( .A(n5498), .B(n5497), .ZN(n9057) );
  NOR2_X1 U5594 ( .A1(n8558), .A2(n9455), .ZN(n5227) );
  AOI21_X1 U5595 ( .B1(n9188), .B2(n6782), .A(n6781), .ZN(n9178) );
  INV_X1 U5596 ( .A(n9214), .ZN(n5717) );
  AND2_X1 U5597 ( .A1(n5715), .A2(n6760), .ZN(n5714) );
  NAND2_X1 U5598 ( .A1(n9214), .A2(n5716), .ZN(n5715) );
  INV_X1 U5599 ( .A(n6750), .ZN(n5716) );
  INV_X1 U5600 ( .A(n9034), .ZN(n9204) );
  NAND2_X1 U5601 ( .A1(n9222), .A2(n9226), .ZN(n6751) );
  NAND2_X1 U5602 ( .A1(n5664), .A2(n9223), .ZN(n9229) );
  INV_X1 U5603 ( .A(n9227), .ZN(n5664) );
  NAND2_X1 U5604 ( .A1(n5267), .A2(n5726), .ZN(n9222) );
  INV_X1 U5605 ( .A(n9244), .ZN(n9239) );
  AND4_X1 U5606 ( .A1(n6713), .A2(n6712), .A3(n6711), .A4(n6710), .ZN(n9257)
         );
  AOI21_X1 U5607 ( .B1(n9280), .B2(n5378), .A(n5377), .ZN(n5376) );
  INV_X1 U5608 ( .A(n8975), .ZN(n5377) );
  INV_X1 U5609 ( .A(n6828), .ZN(n5378) );
  NAND2_X1 U5610 ( .A1(n9310), .A2(n8970), .ZN(n9296) );
  AND2_X1 U5611 ( .A1(n8970), .A2(n8967), .ZN(n9311) );
  OAI21_X1 U5612 ( .B1(n5718), .B2(n9330), .A(n5158), .ZN(n5248) );
  NAND2_X1 U5613 ( .A1(n5721), .A2(n6642), .ZN(n5720) );
  INV_X1 U5614 ( .A(n5718), .ZN(n5247) );
  AND4_X1 U5615 ( .A1(n6652), .A2(n6651), .A3(n6650), .A4(n6649), .ZN(n9359)
         );
  AND2_X1 U5616 ( .A1(n8955), .A2(n6630), .ZN(n9370) );
  OAI21_X1 U5617 ( .B1(n6617), .B2(n9039), .A(n9462), .ZN(n6618) );
  INV_X1 U5618 ( .A(n5389), .ZN(n8374) );
  OAI21_X1 U5619 ( .B1(n6819), .B2(n8326), .A(n6821), .ZN(n5389) );
  OR2_X1 U5620 ( .A1(n6579), .A2(n6578), .ZN(n6580) );
  INV_X1 U5621 ( .A(n9361), .ZN(n9339) );
  NOR2_X1 U5622 ( .A1(n8919), .A2(n5386), .ZN(n5385) );
  INV_X1 U5623 ( .A(n8910), .ZN(n5386) );
  AND2_X1 U5624 ( .A1(n8910), .A2(n8912), .ZN(n8853) );
  NAND2_X1 U5625 ( .A1(n7835), .A2(n8897), .ZN(n7834) );
  NAND2_X1 U5626 ( .A1(n7486), .A2(n7485), .ZN(n8888) );
  AND2_X1 U5627 ( .A1(n7595), .A2(n6836), .ZN(n8385) );
  NAND2_X1 U5628 ( .A1(n7590), .A2(n7589), .ZN(n7592) );
  AND2_X1 U5629 ( .A1(n7588), .A2(n7587), .ZN(n7590) );
  INV_X1 U5630 ( .A(n9376), .ZN(n9337) );
  AND2_X1 U5631 ( .A1(n6861), .A2(n7145), .ZN(n7582) );
  OR2_X1 U5632 ( .A1(n7144), .A2(P2_D_REG_0__SCAN_IN), .ZN(n6861) );
  AND2_X1 U5633 ( .A1(n9463), .A2(n7513), .ZN(n9466) );
  NAND2_X1 U5634 ( .A1(n6741), .A2(n6740), .ZN(n8991) );
  NAND2_X1 U5635 ( .A1(n6673), .A2(n6672), .ZN(n9433) );
  INV_X1 U5636 ( .A(n9450), .ZN(n9463) );
  NAND2_X1 U5637 ( .A1(n7477), .A2(n6874), .ZN(n9342) );
  AND2_X1 U5638 ( .A1(n7505), .A2(n7150), .ZN(n7513) );
  XNOR2_X1 U5639 ( .A(n6850), .B(P2_IR_REG_26__SCAN_IN), .ZN(n6885) );
  NAND2_X1 U5640 ( .A1(n6851), .A2(n5737), .ZN(n6849) );
  NAND2_X1 U5641 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n6454) );
  INV_X1 U5642 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6418) );
  NAND2_X1 U5643 ( .A1(n6472), .A2(n6471), .ZN(n7207) );
  INV_X1 U5644 ( .A(n7038), .ZN(n5623) );
  NOR2_X1 U5645 ( .A1(n5613), .A2(n9611), .ZN(n5609) );
  INV_X1 U5646 ( .A(n7079), .ZN(n5613) );
  NAND2_X1 U5647 ( .A1(n5612), .A2(n7079), .ZN(n5611) );
  INV_X1 U5648 ( .A(n9610), .ZN(n5612) );
  OR2_X1 U5649 ( .A1(n6979), .A2(n5644), .ZN(n9656) );
  NOR2_X1 U5650 ( .A1(n5622), .A2(n7038), .ZN(n5621) );
  INV_X1 U5651 ( .A(n7036), .ZN(n5622) );
  NAND2_X1 U5652 ( .A1(n7035), .A2(n9598), .ZN(n9601) );
  INV_X1 U5653 ( .A(n7984), .ZN(n5630) );
  AND2_X1 U5654 ( .A1(n5638), .A2(n6952), .ZN(n5629) );
  NAND2_X1 U5655 ( .A1(n6949), .A2(n6950), .ZN(n5638) );
  AND2_X1 U5656 ( .A1(n9969), .A2(n9968), .ZN(n9965) );
  AOI21_X1 U5657 ( .B1(n5420), .B2(n5419), .A(n5418), .ZN(n5417) );
  INV_X1 U5658 ( .A(n9947), .ZN(n5418) );
  INV_X1 U5659 ( .A(n6345), .ZN(n5419) );
  NAND2_X1 U5660 ( .A1(n5708), .A2(n5176), .ZN(n5284) );
  OR2_X1 U5661 ( .A1(n10237), .A2(n10248), .ZN(n10208) );
  AOI21_X1 U5662 ( .B1(n5281), .B2(n5279), .A(n5181), .ZN(n5278) );
  INV_X1 U5663 ( .A(n9770), .ZN(n5279) );
  INV_X1 U5664 ( .A(n5281), .ZN(n5280) );
  INV_X1 U5665 ( .A(n5173), .ZN(n5283) );
  NAND2_X1 U5666 ( .A1(n8535), .A2(n5179), .ZN(n5408) );
  OR2_X1 U5667 ( .A1(n8530), .A2(n10297), .ZN(n9920) );
  NAND2_X1 U5668 ( .A1(n10396), .A2(n5162), .ZN(n8526) );
  NAND2_X1 U5669 ( .A1(n8526), .A2(n9792), .ZN(n8525) );
  INV_X1 U5670 ( .A(n5423), .ZN(n5422) );
  AOI21_X1 U5671 ( .B1(n5137), .B2(n5705), .A(n5191), .ZN(n5704) );
  INV_X1 U5672 ( .A(n6109), .ZN(n5705) );
  NAND2_X1 U5673 ( .A1(n8103), .A2(n5425), .ZN(n8197) );
  NAND2_X1 U5674 ( .A1(n8099), .A2(n6093), .ZN(n6094) );
  OR2_X1 U5675 ( .A1(n8108), .A2(n11087), .ZN(n6093) );
  AND2_X1 U5676 ( .A1(n9879), .A2(n9881), .ZN(n9783) );
  NAND2_X1 U5677 ( .A1(n7711), .A2(n9779), .ZN(n6339) );
  NAND2_X1 U5678 ( .A1(n7883), .A2(n7884), .ZN(n7882) );
  NAND2_X1 U5679 ( .A1(n5693), .A2(n5696), .ZN(n5691) );
  NOR2_X1 U5680 ( .A1(n6031), .A2(n6030), .ZN(n6044) );
  AND2_X1 U5681 ( .A1(n5694), .A2(n9858), .ZN(n5693) );
  NAND2_X1 U5682 ( .A1(n5695), .A2(n6037), .ZN(n5694) );
  INV_X1 U5683 ( .A(n6037), .ZN(n5696) );
  NAND2_X1 U5684 ( .A1(n7713), .A2(n9852), .ZN(n7712) );
  NAND2_X1 U5685 ( .A1(n7550), .A2(n7549), .ZN(n7548) );
  NAND2_X1 U5686 ( .A1(n6350), .A2(n6349), .ZN(n10411) );
  OR2_X1 U5687 ( .A1(n9808), .A2(n8497), .ZN(n10388) );
  INV_X1 U5688 ( .A(n5889), .ZN(n6152) );
  INV_X1 U5689 ( .A(n10411), .ZN(n11022) );
  OAI21_X1 U5690 ( .B1(n8599), .B2(n10497), .A(n8598), .ZN(n8629) );
  OR2_X1 U5691 ( .A1(n8597), .A2(n8596), .ZN(n8598) );
  XNOR2_X1 U5692 ( .A(n6289), .B(n6288), .ZN(n8380) );
  NAND2_X1 U5693 ( .A1(n5361), .A2(n6271), .ZN(n6289) );
  NAND2_X1 U5694 ( .A1(n6255), .A2(n5365), .ZN(n5361) );
  NAND2_X1 U5695 ( .A1(n5649), .A2(n5648), .ZN(n6365) );
  NOR2_X1 U5696 ( .A1(n5650), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n5648) );
  INV_X1 U5697 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6150) );
  OAI21_X1 U5698 ( .B1(n5895), .B2(n5813), .A(n5812), .ZN(n5888) );
  NAND2_X1 U5699 ( .A1(n5343), .A2(n5344), .ZN(n5915) );
  INV_X1 U5700 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5709) );
  XNOR2_X1 U5701 ( .A(n5351), .B(n5338), .ZN(n7162) );
  INV_X1 U5702 ( .A(n5751), .ZN(n5338) );
  AOI21_X1 U5703 ( .B1(n5357), .B2(n5355), .A(n5354), .ZN(n5351) );
  NAND2_X1 U5704 ( .A1(n5357), .A2(n5780), .ZN(n6039) );
  NAND2_X1 U5705 ( .A1(n5774), .A2(n5773), .ZN(n6012) );
  NAND2_X1 U5706 ( .A1(n5290), .A2(n5767), .ZN(n6006) );
  NAND2_X1 U5707 ( .A1(n6685), .A2(n6684), .ZN(n9298) );
  AND4_X1 U5708 ( .A1(n6749), .A2(n6748), .A3(n6747), .A4(n6746), .ZN(n9242)
         );
  NAND2_X1 U5709 ( .A1(n5514), .A2(n5513), .ZN(n8755) );
  AOI21_X1 U5710 ( .B1(n5515), .B2(n5518), .A(n5168), .ZN(n5513) );
  AND4_X1 U5711 ( .A1(n6513), .A2(n6512), .A3(n6511), .A4(n6510), .ZN(n8150)
         );
  INV_X1 U5712 ( .A(n9324), .ZN(n8765) );
  NAND2_X1 U5713 ( .A1(n8091), .A2(n8090), .ZN(n8221) );
  NAND2_X1 U5714 ( .A1(n6475), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6469) );
  NAND2_X1 U5715 ( .A1(n6476), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6467) );
  INV_X1 U5716 ( .A(n9286), .ZN(n9422) );
  AOI21_X2 U5717 ( .B1(n7187), .B2(n8838), .A(n5229), .ZN(n8339) );
  INV_X1 U5718 ( .A(n6594), .ZN(n5229) );
  NAND2_X1 U5719 ( .A1(n9470), .A2(n9172), .ZN(n5340) );
  MUX2_X1 U5720 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6440), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n6442) );
  NAND2_X1 U5721 ( .A1(n5391), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6440) );
  AND4_X1 U5722 ( .A1(n7815), .A2(n6800), .A3(n6799), .A4(n6798), .ZN(n9179)
         );
  NAND2_X1 U5723 ( .A1(n5237), .A2(n5157), .ZN(n5430) );
  INV_X1 U5724 ( .A(n7851), .ZN(n7852) );
  NAND2_X1 U5725 ( .A1(n5235), .A2(n5154), .ZN(n5439) );
  INV_X1 U5726 ( .A(n5437), .ZN(n8254) );
  INV_X1 U5727 ( .A(n5233), .ZN(n8548) );
  INV_X1 U5728 ( .A(n8588), .ZN(n5503) );
  OAI21_X1 U5729 ( .B1(n9135), .B2(n8552), .A(n5502), .ZN(n5501) );
  NAND2_X1 U5730 ( .A1(n5654), .A2(n6834), .ZN(n5380) );
  NAND2_X1 U5731 ( .A1(n9183), .A2(n9182), .ZN(n5654) );
  INV_X1 U5732 ( .A(n6893), .ZN(n8616) );
  AND2_X1 U5733 ( .A1(n6426), .A2(n6427), .ZN(n5724) );
  XNOR2_X1 U5734 ( .A(n6536), .B(n6540), .ZN(n7997) );
  XNOR2_X1 U5735 ( .A(n6538), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7867) );
  AND4_X1 U5736 ( .A1(n5984), .A2(n5983), .A3(n5982), .A4(n5981), .ZN(n7439)
         );
  INV_X1 U5737 ( .A(n11073), .ZN(n8022) );
  AND2_X1 U5738 ( .A1(n6281), .A2(n6264), .ZN(n10171) );
  NAND2_X1 U5739 ( .A1(n7112), .A2(n7919), .ZN(n9694) );
  INV_X1 U5740 ( .A(n10174), .ZN(n10326) );
  XNOR2_X1 U5741 ( .A(n6317), .B(n9972), .ZN(n10140) );
  INV_X1 U5742 ( .A(n10317), .ZN(n10334) );
  NAND2_X1 U5743 ( .A1(n7553), .A2(n7919), .ZN(n10307) );
  AND2_X1 U5744 ( .A1(n9703), .A2(n9702), .ZN(n10426) );
  AOI21_X1 U5745 ( .B1(n10310), .B2(n10400), .A(n10312), .ZN(n10423) );
  NAND2_X1 U5746 ( .A1(n6310), .A2(n6309), .ZN(n10147) );
  OR2_X1 U5747 ( .A1(n10507), .A2(n5588), .ZN(n5587) );
  NAND2_X1 U5748 ( .A1(n5590), .A2(n5589), .ZN(n5588) );
  NAND2_X1 U5749 ( .A1(keyinput_11), .A2(SI_21_), .ZN(n5589) );
  AOI22_X1 U5750 ( .A1(n10509), .A2(n10685), .B1(keyinput_12), .B2(SI_20_), 
        .ZN(n5586) );
  AOI21_X1 U5751 ( .B1(n5585), .B2(n5584), .A(n5583), .ZN(n10513) );
  XNOR2_X1 U5752 ( .A(n10690), .B(keyinput_15), .ZN(n5583) );
  INV_X1 U5753 ( .A(n10511), .ZN(n5584) );
  NAND2_X1 U5754 ( .A1(n5587), .A2(n5586), .ZN(n5585) );
  OR2_X1 U5755 ( .A1(n10681), .A2(n10682), .ZN(n5493) );
  NOR4_X1 U5756 ( .A1(n10680), .A2(n10679), .A3(n10678), .A4(n10677), .ZN(
        n10681) );
  XNOR2_X1 U5757 ( .A(n5492), .B(keyinput_138), .ZN(n5491) );
  NAND2_X1 U5758 ( .A1(n10685), .A2(keyinput_140), .ZN(n5487) );
  NAND2_X1 U5759 ( .A1(n10686), .A2(SI_20_), .ZN(n5488) );
  AOI21_X1 U5760 ( .B1(n5490), .B2(n5489), .A(n5486), .ZN(n10687) );
  NAND2_X1 U5761 ( .A1(n5488), .A2(n5487), .ZN(n5486) );
  AOI22_X1 U5762 ( .A1(n10683), .A2(n10684), .B1(keyinput_139), .B2(SI_21_), 
        .ZN(n5489) );
  NAND2_X1 U5763 ( .A1(n5493), .A2(n5491), .ZN(n5490) );
  NAND2_X1 U5764 ( .A1(n5443), .A2(n10696), .ZN(n10701) );
  OAI21_X1 U5765 ( .B1(n5444), .B2(n10691), .A(n10693), .ZN(n5443) );
  INV_X1 U5766 ( .A(n10545), .ZN(n5596) );
  NAND2_X1 U5767 ( .A1(n5599), .A2(n5598), .ZN(n5597) );
  NAND2_X1 U5768 ( .A1(n10544), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5598) );
  NAND2_X1 U5769 ( .A1(n10724), .A2(keyinput_37), .ZN(n5599) );
  NAND2_X1 U5770 ( .A1(n10729), .A2(n10546), .ZN(n5593) );
  NAND2_X1 U5771 ( .A1(keyinput_41), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5592)
         );
  NAND2_X1 U5772 ( .A1(n8918), .A2(n9018), .ZN(n5331) );
  AOI21_X1 U5773 ( .B1(n5595), .B2(n5594), .A(n5591), .ZN(n10552) );
  XNOR2_X1 U5774 ( .A(n6486), .B(keyinput_40), .ZN(n5594) );
  NAND2_X1 U5775 ( .A1(n5593), .A2(n5592), .ZN(n5591) );
  OAI21_X1 U5776 ( .B1(n10543), .B2(n5597), .A(n5596), .ZN(n5595) );
  NAND2_X1 U5777 ( .A1(n11020), .A2(n10720), .ZN(n5485) );
  NAND2_X1 U5778 ( .A1(keyinput_161), .A2(P2_RD_REG_SCAN_IN), .ZN(n5484) );
  AND3_X1 U5779 ( .A1(n5328), .A2(n5329), .A3(n5324), .ZN(n8933) );
  AND2_X1 U5780 ( .A1(n5332), .A2(n5330), .ZN(n5324) );
  NAND2_X1 U5781 ( .A1(n5572), .A2(n5570), .ZN(n5569) );
  XNOR2_X1 U5782 ( .A(n5571), .B(P2_REG3_REG_5__SCAN_IN), .ZN(n5570) );
  NAND2_X1 U5783 ( .A1(n10553), .A2(n10554), .ZN(n5572) );
  INV_X1 U5784 ( .A(keyinput_49), .ZN(n5571) );
  INV_X1 U5785 ( .A(n10563), .ZN(n5566) );
  NOR2_X1 U5786 ( .A1(n10565), .A2(n10564), .ZN(n5565) );
  AOI21_X1 U5787 ( .B1(n5481), .B2(n5479), .A(n5476), .ZN(n10725) );
  AND2_X1 U5788 ( .A1(n10735), .A2(n10734), .ZN(n5468) );
  INV_X1 U5789 ( .A(n8949), .ZN(n5302) );
  OAI211_X1 U5790 ( .C1(n5333), .C2(n8937), .A(n5326), .B(n5325), .ZN(n8940)
         );
  NAND2_X1 U5791 ( .A1(n8934), .A2(n5327), .ZN(n5325) );
  NAND2_X1 U5792 ( .A1(n8936), .A2(n8935), .ZN(n5333) );
  NAND2_X1 U5793 ( .A1(n5323), .A2(n9018), .ZN(n5318) );
  NAND2_X1 U5794 ( .A1(n5322), .A2(n9007), .ZN(n5319) );
  INV_X1 U5795 ( .A(n8967), .ZN(n5322) );
  AOI21_X1 U5796 ( .B1(n10573), .B2(n5562), .A(n5561), .ZN(n5560) );
  OAI22_X1 U5797 ( .A1(n10763), .A2(keyinput_67), .B1(n10575), .B2(
        P2_DATAO_REG_29__SCAN_IN), .ZN(n5561) );
  INV_X1 U5798 ( .A(n5563), .ZN(n5562) );
  AOI211_X1 U5799 ( .C1(n5466), .C2(n5463), .A(n5462), .B(n10741), .ZN(n10750)
         );
  AND2_X1 U5800 ( .A1(n10742), .A2(n5219), .ZN(n5462) );
  AND2_X1 U5801 ( .A1(n5464), .A2(n10742), .ZN(n5463) );
  NAND2_X1 U5802 ( .A1(n5184), .A2(n9007), .ZN(n5316) );
  AND2_X1 U5803 ( .A1(n5295), .A2(n5204), .ZN(n5292) );
  AND2_X1 U5804 ( .A1(n5558), .A2(n5557), .ZN(n10578) );
  NAND2_X1 U5805 ( .A1(n8116), .A2(keyinput_73), .ZN(n5557) );
  OAI21_X1 U5806 ( .B1(n5560), .B2(n5559), .A(n10577), .ZN(n5558) );
  OAI22_X1 U5807 ( .A1(n10768), .A2(n10576), .B1(P2_DATAO_REG_28__SCAN_IN), 
        .B2(keyinput_68), .ZN(n5559) );
  XNOR2_X1 U5808 ( .A(n5604), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n5603) );
  INV_X1 U5809 ( .A(keyinput_76), .ZN(n5604) );
  NAND2_X1 U5810 ( .A1(n5310), .A2(n5308), .ZN(n8977) );
  AND2_X1 U5811 ( .A1(n5321), .A2(n5309), .ZN(n5308) );
  NOR2_X1 U5812 ( .A1(n5461), .A2(n5460), .ZN(n5459) );
  INV_X1 U5813 ( .A(n10771), .ZN(n5460) );
  NOR2_X1 U5814 ( .A1(n5461), .A2(n5458), .ZN(n5457) );
  NOR2_X1 U5815 ( .A1(n10779), .A2(n5217), .ZN(n5458) );
  INV_X1 U5816 ( .A(keyinput_211), .ZN(n5473) );
  OR2_X1 U5817 ( .A1(n10591), .A2(n5581), .ZN(n5580) );
  NAND2_X1 U5818 ( .A1(n10596), .A2(n5582), .ZN(n5581) );
  NAND2_X1 U5819 ( .A1(keyinput_85), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n5582)
         );
  NOR2_X1 U5820 ( .A1(n10594), .A2(n5579), .ZN(n5578) );
  AND2_X1 U5821 ( .A1(n10595), .A2(keyinput_87), .ZN(n5579) );
  INV_X1 U5822 ( .A(n10601), .ZN(n5575) );
  NOR2_X1 U5823 ( .A1(n10600), .A2(n10599), .ZN(n5574) );
  XNOR2_X1 U5824 ( .A(n5473), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n5472) );
  NAND2_X1 U5825 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n5475), .ZN(n5474) );
  INV_X1 U5826 ( .A(keyinput_207), .ZN(n5475) );
  AOI21_X1 U5827 ( .B1(n5577), .B2(n5576), .A(n5573), .ZN(n10604) );
  AOI22_X1 U5828 ( .A1(n10597), .A2(n10795), .B1(keyinput_88), .B2(
        P2_DATAO_REG_8__SCAN_IN), .ZN(n5576) );
  NAND2_X1 U5829 ( .A1(n5575), .A2(n5574), .ZN(n5573) );
  NAND2_X1 U5830 ( .A1(n5580), .A2(n5578), .ZN(n5577) );
  NOR2_X1 U5831 ( .A1(n5470), .A2(n5469), .ZN(n10801) );
  OR2_X1 U5832 ( .A1(n10793), .A2(n5224), .ZN(n5469) );
  AOI21_X1 U5833 ( .B1(n10788), .B2(n5474), .A(n5471), .ZN(n5470) );
  AOI21_X1 U5834 ( .B1(n5456), .B2(n5455), .A(n10822), .ZN(n5454) );
  INV_X1 U5835 ( .A(n10820), .ZN(n5455) );
  AOI21_X1 U5836 ( .B1(n5454), .B2(n10819), .A(n5223), .ZN(n5453) );
  INV_X1 U5837 ( .A(SI_20_), .ZN(n10685) );
  INV_X1 U5838 ( .A(SI_19_), .ZN(n10667) );
  INV_X1 U5839 ( .A(SI_14_), .ZN(n10695) );
  INV_X1 U5840 ( .A(SI_11_), .ZN(n10491) );
  INV_X1 U5841 ( .A(SI_8_), .ZN(n10518) );
  NAND2_X1 U5842 ( .A1(n5305), .A2(n5303), .ZN(n9017) );
  AOI21_X1 U5843 ( .B1(n8569), .B2(n9138), .A(n8568), .ZN(n8571) );
  AOI21_X1 U5844 ( .B1(n5453), .B2(n5451), .A(n5450), .ZN(n5449) );
  INV_X1 U5845 ( .A(n10828), .ZN(n5450) );
  INV_X1 U5846 ( .A(n5454), .ZN(n5451) );
  INV_X1 U5847 ( .A(n5453), .ZN(n5452) );
  INV_X1 U5848 ( .A(n10833), .ZN(n5448) );
  INV_X1 U5849 ( .A(n5363), .ZN(n5362) );
  OAI21_X1 U5850 ( .B1(n5365), .B2(n5364), .A(n6288), .ZN(n5363) );
  INV_X1 U5851 ( .A(n6271), .ZN(n5364) );
  INV_X1 U5852 ( .A(SI_26_), .ZN(n10673) );
  INV_X1 U5853 ( .A(SI_21_), .ZN(n10684) );
  AND2_X1 U5854 ( .A1(n6143), .A2(n5826), .ZN(n5827) );
  INV_X1 U5855 ( .A(n5672), .ZN(n5671) );
  NAND2_X1 U5856 ( .A1(n5815), .A2(n5814), .ZN(n5818) );
  INV_X1 U5857 ( .A(SI_12_), .ZN(n10664) );
  OAI21_X1 U5858 ( .B1(n5355), .B2(n5354), .A(n5751), .ZN(n5353) );
  NOR2_X1 U5859 ( .A1(n6659), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6675) );
  NAND2_X1 U5860 ( .A1(n8877), .A2(n8875), .ZN(n9019) );
  AND2_X1 U5861 ( .A1(n5737), .A2(n5736), .ZN(n5735) );
  INV_X1 U5862 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5736) );
  XNOR2_X1 U5863 ( .A(n7229), .B(n7223), .ZN(n7210) );
  NAND2_X1 U5864 ( .A1(n5712), .A2(n5264), .ZN(n5263) );
  NAND2_X1 U5865 ( .A1(n5714), .A2(n9223), .ZN(n5264) );
  INV_X1 U5866 ( .A(n8691), .ZN(n5713) );
  AOI21_X1 U5867 ( .B1(n5728), .B2(n5727), .A(n5190), .ZN(n5726) );
  INV_X1 U5868 ( .A(n6703), .ZN(n5727) );
  OR2_X1 U5869 ( .A1(n6572), .A2(n6571), .ZN(n6577) );
  AND2_X1 U5870 ( .A1(n6425), .A2(n6855), .ZN(n5737) );
  INV_X1 U5871 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6888) );
  NOR2_X1 U5872 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5555) );
  AND2_X1 U5873 ( .A1(n9568), .A2(n9659), .ZN(n6992) );
  OAI21_X1 U5874 ( .B1(n7024), .B2(n7023), .A(n9597), .ZN(n7025) );
  NAND2_X1 U5875 ( .A1(n5653), .A2(n6127), .ZN(n5652) );
  INV_X1 U5876 ( .A(n6112), .ZN(n5653) );
  OR2_X1 U5877 ( .A1(n10147), .A2(n8714), .ZN(n9974) );
  INV_X1 U5878 ( .A(n10325), .ZN(n7080) );
  NAND2_X1 U5879 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(n6133), .ZN(n6169) );
  OR2_X1 U5880 ( .A1(n5908), .A2(n5901), .ZN(n5903) );
  INV_X1 U5881 ( .A(n9892), .ZN(n5424) );
  OR2_X1 U5882 ( .A1(n9695), .A2(n9523), .ZN(n9909) );
  AND2_X1 U5883 ( .A1(n6102), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n6104) );
  INV_X1 U5884 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6063) );
  INV_X1 U5885 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5919) );
  INV_X1 U5886 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6054) );
  INV_X1 U5887 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6030) );
  NAND2_X1 U5888 ( .A1(n5269), .A2(n7946), .ZN(n9731) );
  NAND2_X1 U5889 ( .A1(n7567), .A2(n5178), .ZN(n9729) );
  NAND2_X1 U5890 ( .A1(n10200), .A2(n5399), .ZN(n10189) );
  OR2_X1 U5891 ( .A1(n8203), .A2(n8207), .ZN(n8360) );
  NAND2_X1 U5892 ( .A1(n7690), .A2(n5978), .ZN(n7550) );
  OR2_X1 U5893 ( .A1(n10466), .A2(n6384), .ZN(n7104) );
  NAND2_X1 U5894 ( .A1(n6308), .A2(n6307), .ZN(n8597) );
  NOR2_X1 U5895 ( .A1(n6272), .A2(n5366), .ZN(n5365) );
  INV_X1 U5896 ( .A(n6254), .ZN(n5366) );
  NAND2_X1 U5897 ( .A1(n6237), .A2(n6236), .ZN(n6251) );
  INV_X1 U5898 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6110) );
  AOI21_X1 U5899 ( .B1(n5347), .B2(n5345), .A(n5188), .ZN(n5344) );
  INV_X1 U5900 ( .A(n5801), .ZN(n5345) );
  INV_X1 U5901 ( .A(n5347), .ZN(n5346) );
  INV_X1 U5902 ( .A(n6077), .ZN(n5802) );
  OAI21_X2 U5903 ( .B1(n5926), .B2(n5792), .A(n5795), .ZN(n6072) );
  NOR2_X1 U5904 ( .A1(n6038), .A2(n5356), .ZN(n5355) );
  INV_X1 U5905 ( .A(n5780), .ZN(n5356) );
  INV_X1 U5906 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n10803) );
  OAI211_X1 U5907 ( .C1(n5686), .C2(n5684), .A(n5681), .B(n5680), .ZN(n5759)
         );
  NAND2_X1 U5908 ( .A1(n5682), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5681) );
  INV_X1 U5909 ( .A(n5685), .ZN(n5682) );
  OR2_X1 U5910 ( .A1(n7487), .A2(n9050), .ZN(n7488) );
  INV_X1 U5911 ( .A(n5148), .ZN(n5526) );
  AOI21_X1 U5912 ( .B1(n5528), .B2(n5530), .A(n5211), .ZN(n5527) );
  INV_X1 U5913 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10732) );
  NAND2_X1 U5914 ( .A1(n10658), .A2(n6648), .ZN(n6659) );
  AND2_X1 U5915 ( .A1(n8645), .A2(n8648), .ZN(n5536) );
  NAND2_X1 U5916 ( .A1(n6708), .A2(n6707), .ZN(n6716) );
  OR2_X1 U5917 ( .A1(n6566), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6582) );
  NOR2_X1 U5918 ( .A1(n6582), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6599) );
  NOR2_X1 U5919 ( .A1(n9051), .A2(n7479), .ZN(n7482) );
  NOR2_X1 U5920 ( .A1(n5533), .A2(n5532), .ZN(n5531) );
  INV_X1 U5921 ( .A(n8812), .ZN(n5532) );
  AND2_X1 U5922 ( .A1(n8637), .A2(n5516), .ZN(n5515) );
  NAND2_X1 U5923 ( .A1(n5519), .A2(n5517), .ZN(n5516) );
  INV_X1 U5924 ( .A(n8516), .ZN(n5517) );
  INV_X1 U5925 ( .A(n5519), .ZN(n5518) );
  NAND2_X1 U5926 ( .A1(n9015), .A2(n9014), .ZN(n9024) );
  NOR2_X1 U5927 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n6423) );
  INV_X1 U5928 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6420) );
  AND4_X1 U5929 ( .A1(n6481), .A2(n6480), .A3(n6479), .A4(n6478), .ZN(n7542)
         );
  NAND2_X1 U5930 ( .A1(n5232), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10946) );
  OR2_X1 U5931 ( .A1(n10938), .A2(n10937), .ZN(n10940) );
  INV_X1 U5932 ( .A(n5432), .ZN(n5431) );
  AND2_X1 U5933 ( .A1(n5432), .A2(n5435), .ZN(n10980) );
  NAND2_X1 U5934 ( .A1(n5495), .A2(n7244), .ZN(n5496) );
  NOR2_X1 U5935 ( .A1(n7632), .A2(n7631), .ZN(n7633) );
  NOR2_X1 U5936 ( .A1(n7868), .A2(n7869), .ZN(n7872) );
  NOR2_X1 U5937 ( .A1(n8002), .A2(n8001), .ZN(n8003) );
  AND2_X1 U5938 ( .A1(n7997), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5428) );
  NAND2_X1 U5939 ( .A1(n5508), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5507) );
  INV_X1 U5940 ( .A(n8187), .ZN(n5508) );
  NOR2_X1 U5941 ( .A1(n7998), .A2(n7999), .ZN(n8184) );
  NOR2_X1 U5942 ( .A1(n8273), .A2(n8502), .ZN(n5236) );
  NOR2_X1 U5943 ( .A1(n9066), .A2(n9067), .ZN(n9065) );
  INV_X1 U5944 ( .A(n5498), .ZN(n8578) );
  OAI21_X1 U5945 ( .B1(n9097), .B2(n5510), .A(n5509), .ZN(n9119) );
  NAND2_X1 U5946 ( .A1(n5511), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5510) );
  NOR2_X1 U5947 ( .A1(n9097), .A2(n8556), .ZN(n9096) );
  AND2_X1 U5948 ( .A1(n6670), .A2(n6592), .ZN(n5550) );
  AND2_X1 U5949 ( .A1(n9004), .A2(n9003), .ZN(n9195) );
  OAI21_X1 U5950 ( .B1(n9227), .B2(n5658), .A(n5656), .ZN(n9193) );
  INV_X1 U5951 ( .A(n5659), .ZN(n5658) );
  AOI21_X1 U5952 ( .B1(n5659), .B2(n5661), .A(n5657), .ZN(n5656) );
  NAND2_X1 U5953 ( .A1(n5655), .A2(n5659), .ZN(n8869) );
  NAND2_X1 U5954 ( .A1(n9227), .A2(n5662), .ZN(n5655) );
  NAND2_X1 U5955 ( .A1(n6743), .A2(n6742), .ZN(n6754) );
  OR2_X1 U5956 ( .A1(n6736), .A2(n6735), .ZN(n9237) );
  OR2_X1 U5957 ( .A1(n8986), .A2(n8848), .ZN(n9244) );
  NAND2_X1 U5958 ( .A1(n5206), .A2(n5379), .ZN(n9277) );
  NAND2_X1 U5959 ( .A1(n5723), .A2(n5177), .ZN(n9290) );
  NAND2_X1 U5960 ( .A1(n5193), .A2(n6827), .ZN(n5387) );
  INV_X1 U5961 ( .A(n5687), .ZN(n6824) );
  NOR2_X1 U5962 ( .A1(n6637), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6648) );
  INV_X1 U5963 ( .A(n9370), .ZN(n9368) );
  NAND2_X1 U5964 ( .A1(n8374), .A2(n8927), .ZN(n8504) );
  AND2_X1 U5965 ( .A1(n8503), .A2(n8946), .ZN(n8950) );
  OR2_X1 U5966 ( .A1(n6818), .A2(n8860), .ZN(n8372) );
  AND2_X1 U5967 ( .A1(n8938), .A2(n8925), .ZN(n8860) );
  INV_X1 U5968 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n10556) );
  AND2_X1 U5969 ( .A1(n6816), .A2(n8930), .ZN(n5754) );
  NAND2_X1 U5970 ( .A1(n5754), .A2(n6817), .ZN(n8312) );
  INV_X1 U5971 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6543) );
  INV_X1 U5972 ( .A(n5253), .ZN(n5252) );
  OAI21_X1 U5973 ( .B1(n5255), .B2(n5254), .A(n6522), .ZN(n5253) );
  OR2_X1 U5974 ( .A1(n6508), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6523) );
  NAND2_X1 U5975 ( .A1(n7467), .A2(n5260), .ZN(n7448) );
  NAND2_X1 U5976 ( .A1(n7486), .A2(n7976), .ZN(n5260) );
  OAI21_X1 U5977 ( .B1(n7469), .B2(n7468), .A(n8849), .ZN(n7467) );
  AND2_X1 U5978 ( .A1(n8851), .A2(n5261), .ZN(n7469) );
  INV_X1 U5979 ( .A(n7481), .ZN(n5261) );
  INV_X1 U5980 ( .A(n8851), .ZN(n7433) );
  OR2_X1 U5981 ( .A1(n9007), .A2(n6895), .ZN(n7500) );
  OR2_X1 U5982 ( .A1(n9007), .A2(n6896), .ZN(n7583) );
  NAND2_X1 U5983 ( .A1(n8843), .A2(n8842), .ZN(n8845) );
  NAND2_X1 U5984 ( .A1(n6796), .A2(n6795), .ZN(n6893) );
  NAND2_X1 U5985 ( .A1(n6762), .A2(n6761), .ZN(n6832) );
  NAND2_X1 U5986 ( .A1(n6753), .A2(n6752), .ZN(n8685) );
  NAND2_X1 U5987 ( .A1(n6715), .A2(n6714), .ZN(n8982) );
  NAND2_X1 U5988 ( .A1(n5256), .A2(n5255), .ZN(n8125) );
  NAND2_X1 U5989 ( .A1(n5734), .A2(n5139), .ZN(n5256) );
  AND3_X1 U5990 ( .A1(n6452), .A2(n6451), .A3(n6450), .ZN(n8012) );
  INV_X1 U5991 ( .A(n5734), .ZN(n7837) );
  NAND2_X1 U5992 ( .A1(n7892), .A2(n8060), .ZN(n9450) );
  NAND2_X1 U5993 ( .A1(n6885), .A2(n6858), .ZN(n7144) );
  INV_X1 U5994 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6855) );
  NAND2_X1 U5995 ( .A1(n6805), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6806) );
  NAND2_X1 U5996 ( .A1(n6590), .A2(n6589), .ZN(n6614) );
  NAND2_X1 U5997 ( .A1(n5551), .A2(n6592), .ZN(n6665) );
  INV_X1 U5998 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6537) );
  OR2_X1 U5999 ( .A1(n6445), .A2(n6446), .ZN(n6491) );
  INV_X1 U6000 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n6558) );
  NAND2_X1 U6001 ( .A1(n6186), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6209) );
  NAND2_X1 U6002 ( .A1(n7302), .A2(n6930), .ZN(n6935) );
  XNOR2_X1 U6003 ( .A(n6933), .B(n8706), .ZN(n6936) );
  NOR2_X1 U6004 ( .A1(n6064), .A2(n6063), .ZN(n6087) );
  INV_X1 U6005 ( .A(n10001), .ZN(n5269) );
  NOR2_X1 U6006 ( .A1(n5903), .A2(n5882), .ZN(n6117) );
  NAND2_X1 U6007 ( .A1(n5615), .A2(n7074), .ZN(n5614) );
  NAND2_X1 U6008 ( .A1(n9656), .A2(n9657), .ZN(n9655) );
  AOI21_X1 U6009 ( .B1(n5610), .B2(n5608), .A(n5180), .ZN(n5607) );
  INV_X1 U6010 ( .A(n5609), .ZN(n5608) );
  OR2_X1 U6011 ( .A1(n10856), .A2(n10855), .ZN(n10858) );
  INV_X1 U6012 ( .A(n10426), .ZN(n10127) );
  INV_X1 U6013 ( .A(n9965), .ZN(n9799) );
  NOR2_X1 U6014 ( .A1(n10157), .A2(n5397), .ZN(n5395) );
  AND2_X1 U6015 ( .A1(n9962), .A2(n9963), .ZN(n10153) );
  INV_X1 U6016 ( .A(n6346), .ZN(n10169) );
  NAND2_X1 U6017 ( .A1(n10209), .A2(n5420), .ZN(n10195) );
  NAND2_X1 U6018 ( .A1(n10227), .A2(n6345), .ZN(n10209) );
  AND2_X1 U6019 ( .A1(n5134), .A2(n10368), .ZN(n5400) );
  NAND2_X1 U6020 ( .A1(n8527), .A2(n5402), .ZN(n10298) );
  INV_X1 U6021 ( .A(n6156), .ZN(n6133) );
  NAND2_X1 U6022 ( .A1(n8527), .A2(n10390), .ZN(n10301) );
  AND2_X1 U6023 ( .A1(n8492), .A2(n8457), .ZN(n8527) );
  NOR2_X1 U6024 ( .A1(n8360), .A2(n9527), .ZN(n8458) );
  AND2_X1 U6025 ( .A1(n9901), .A2(n9892), .ZN(n9785) );
  NAND2_X1 U6026 ( .A1(n6085), .A2(n6084), .ZN(n8108) );
  NAND2_X1 U6027 ( .A1(n8106), .A2(n11104), .ZN(n8203) );
  NAND2_X1 U6028 ( .A1(n7879), .A2(n5141), .ZN(n5270) );
  NAND2_X1 U6029 ( .A1(n5413), .A2(n5415), .ZN(n5411) );
  INV_X1 U6030 ( .A(n5414), .ZN(n5413) );
  NAND2_X1 U6031 ( .A1(n7879), .A2(n5699), .ZN(n7907) );
  AND2_X1 U6032 ( .A1(n7910), .A2(n5698), .ZN(n8106) );
  AND4_X1 U6033 ( .A1(n6036), .A2(n6035), .A3(n6034), .A4(n6033), .ZN(n8235)
         );
  NOR2_X1 U6034 ( .A1(n7944), .A2(n8022), .ZN(n7714) );
  OR2_X1 U6035 ( .A1(n7943), .A2(n7946), .ZN(n7944) );
  NOR2_X1 U6036 ( .A1(n7555), .A2(n5994), .ZN(n7684) );
  NAND2_X1 U6037 ( .A1(n7684), .A2(n6009), .ZN(n7943) );
  NAND2_X1 U6038 ( .A1(n7567), .A2(n6333), .ZN(n9832) );
  NAND2_X1 U6039 ( .A1(n7571), .A2(n7572), .ZN(n7570) );
  INV_X1 U6040 ( .A(n5130), .ZN(n9987) );
  NAND2_X1 U6041 ( .A1(n9711), .A2(n9710), .ZN(n10135) );
  NAND2_X1 U6042 ( .A1(n5859), .A2(n5858), .ZN(n10253) );
  NAND2_X1 U6043 ( .A1(n5706), .A2(n5137), .ZN(n8355) );
  AND2_X1 U6044 ( .A1(n5706), .A2(n5156), .ZN(n8356) );
  NAND2_X1 U6045 ( .A1(n5707), .A2(n6109), .ZN(n5706) );
  OR2_X1 U6046 ( .A1(n5690), .A2(n5689), .ZN(n7694) );
  OAI21_X1 U6047 ( .B1(n5889), .B2(n7388), .A(n5688), .ZN(n5689) );
  NOR2_X1 U6048 ( .A1(n6458), .A2(n6013), .ZN(n5690) );
  NAND2_X1 U6049 ( .A1(n5889), .A2(n5142), .ZN(n5688) );
  AND2_X1 U6050 ( .A1(n7304), .A2(n7107), .ZN(n7551) );
  AND3_X1 U6051 ( .A1(n7105), .A2(n7104), .A3(n7110), .ZN(n6408) );
  INV_X1 U6052 ( .A(n10375), .ZN(n11088) );
  NOR2_X1 U6053 ( .A1(n10470), .A2(n6098), .ZN(n5274) );
  NOR2_X1 U6054 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n5273) );
  XNOR2_X1 U6055 ( .A(n8629), .B(n8628), .ZN(n8839) );
  AND2_X1 U6056 ( .A1(n6359), .A2(n5861), .ZN(n5852) );
  XNOR2_X1 U6057 ( .A(n6273), .B(n6272), .ZN(n8414) );
  NAND2_X1 U6058 ( .A1(n6255), .A2(n6254), .ZN(n6273) );
  OAI21_X1 U6059 ( .B1(n6365), .B2(n6364), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6366) );
  XNOR2_X1 U6060 ( .A(n6219), .B(n6218), .ZN(n8194) );
  OAI21_X1 U6061 ( .B1(n6196), .B2(n6195), .A(n6194), .ZN(n6203) );
  XNOR2_X1 U6062 ( .A(n6148), .B(n6147), .ZN(n7846) );
  AND2_X1 U6063 ( .A1(n6146), .A2(n6145), .ZN(n6148) );
  XNOR2_X1 U6064 ( .A(n6126), .B(n6125), .ZN(n7793) );
  NAND2_X1 U6065 ( .A1(n5665), .A2(n5669), .ZN(n6124) );
  AOI21_X1 U6066 ( .B1(n5672), .B2(n5673), .A(n5670), .ZN(n5669) );
  AND2_X1 U6067 ( .A1(n5933), .A2(n6073), .ZN(n7617) );
  OR2_X1 U6068 ( .A1(n6040), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5928) );
  OR3_X1 U6069 ( .A1(n6026), .A2(P1_IR_REG_6__SCAN_IN), .A3(
        P1_IR_REG_7__SCAN_IN), .ZN(n6040) );
  NAND2_X1 U6070 ( .A1(n5289), .A2(n5770), .ZN(n5942) );
  NAND2_X1 U6071 ( .A1(n5764), .A2(n5763), .ZN(n5991) );
  NAND2_X1 U6072 ( .A1(n7895), .A2(n5747), .ZN(n7898) );
  NAND2_X1 U6073 ( .A1(n8811), .A2(n8692), .ZN(n8725) );
  NAND2_X1 U6074 ( .A1(n6774), .A2(n6773), .ZN(n9196) );
  AND2_X1 U6075 ( .A1(n5520), .A2(n5161), .ZN(n8518) );
  INV_X1 U6076 ( .A(n5553), .ZN(n5552) );
  NAND2_X1 U6077 ( .A1(n8769), .A2(n8657), .ZN(n8658) );
  NAND2_X1 U6078 ( .A1(n6723), .A2(n6722), .ZN(n8663) );
  XNOR2_X1 U6079 ( .A(n8331), .B(n8330), .ZN(n8332) );
  AND2_X1 U6080 ( .A1(n7519), .A2(n7502), .ZN(n8827) );
  OAI21_X1 U6081 ( .B1(n5527), .B2(n5148), .A(n5523), .ZN(n5522) );
  NAND2_X1 U6082 ( .A1(n5527), .A2(n5524), .ZN(n5523) );
  NAND2_X1 U6083 ( .A1(n5526), .A2(n5529), .ZN(n5524) );
  NAND2_X1 U6084 ( .A1(n5527), .A2(n5526), .ZN(n5525) );
  AND4_X1 U6085 ( .A1(n6570), .A2(n6569), .A3(n6568), .A4(n6567), .ZN(n8390)
         );
  OAI21_X2 U6086 ( .B1(n8331), .B2(n5541), .A(n5539), .ZN(n8466) );
  INV_X1 U6087 ( .A(n5542), .ZN(n5541) );
  AOI21_X1 U6088 ( .B1(n5542), .B2(n5545), .A(n5540), .ZN(n5539) );
  INV_X1 U6089 ( .A(n8406), .ZN(n5540) );
  NAND2_X1 U6090 ( .A1(n5538), .A2(n5542), .ZN(n8407) );
  NAND2_X1 U6091 ( .A1(n8331), .A2(n5544), .ZN(n5538) );
  NAND2_X1 U6092 ( .A1(n5537), .A2(n8645), .ZN(n8782) );
  INV_X1 U6093 ( .A(n9038), .ZN(n9360) );
  NAND2_X1 U6094 ( .A1(n6616), .A2(n6615), .ZN(n9462) );
  NAND2_X1 U6095 ( .A1(n7517), .A2(n9380), .ZN(n8786) );
  AND2_X1 U6096 ( .A1(n8793), .A2(n8790), .ZN(n8652) );
  AND2_X1 U6097 ( .A1(n5547), .A2(n5159), .ZN(n8404) );
  NAND2_X1 U6098 ( .A1(n8331), .A2(n5548), .ZN(n5547) );
  AND2_X1 U6099 ( .A1(n8802), .A2(n8799), .ZN(n8642) );
  OAI21_X1 U6100 ( .B1(n8517), .B2(n5518), .A(n5515), .ZN(n8823) );
  INV_X1 U6101 ( .A(n8788), .ZN(n8824) );
  OR2_X1 U6102 ( .A1(n7500), .A2(n7499), .ZN(n9027) );
  AND4_X1 U6103 ( .A1(n7815), .A2(n6842), .A3(n6841), .A4(n6840), .ZN(n8844)
         );
  OR2_X1 U6104 ( .A1(n7505), .A2(n7132), .ZN(n9045) );
  NAND2_X1 U6105 ( .A1(n5433), .A2(n5435), .ZN(n7201) );
  INV_X1 U6106 ( .A(n5505), .ZN(n10990) );
  INV_X1 U6107 ( .A(n7233), .ZN(n10988) );
  INV_X1 U6108 ( .A(n5235), .ZN(n8167) );
  INV_X1 U6109 ( .A(n5234), .ZN(n8255) );
  INV_X1 U6110 ( .A(n5500), .ZN(n8576) );
  NOR2_X1 U6111 ( .A1(n9092), .A2(n9093), .ZN(n9091) );
  INV_X1 U6112 ( .A(n9164), .ZN(n11010) );
  OAI21_X1 U6113 ( .B1(n9092), .B2(n5441), .A(n5440), .ZN(n9111) );
  NAND2_X1 U6114 ( .A1(n5442), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5441) );
  INV_X1 U6115 ( .A(n9112), .ZN(n5442) );
  XNOR2_X1 U6116 ( .A(n5233), .B(n8553), .ZN(n9128) );
  AND2_X1 U6117 ( .A1(n5504), .A2(n9150), .ZN(n9153) );
  AND2_X1 U6118 ( .A1(n7203), .A2(n7193), .ZN(n10968) );
  AOI21_X1 U6119 ( .B1(n9181), .B2(n9342), .A(n9180), .ZN(n9392) );
  OAI21_X1 U6120 ( .B1(n6751), .B2(n5717), .A(n5714), .ZN(n9202) );
  NAND2_X1 U6121 ( .A1(n6751), .A2(n6750), .ZN(n9211) );
  NAND2_X1 U6122 ( .A1(n9229), .A2(n8992), .ZN(n9215) );
  NAND2_X1 U6123 ( .A1(n6705), .A2(n6704), .ZN(n9418) );
  NAND2_X1 U6124 ( .A1(n9281), .A2(n9280), .ZN(n9283) );
  NAND2_X1 U6125 ( .A1(n9428), .A2(n6828), .ZN(n9281) );
  AND2_X1 U6126 ( .A1(n6696), .A2(n6695), .ZN(n9286) );
  INV_X1 U6127 ( .A(n5248), .ZN(n5243) );
  NAND2_X1 U6128 ( .A1(n6658), .A2(n6657), .ZN(n9437) );
  INV_X1 U6129 ( .A(n5246), .ZN(n9323) );
  AOI21_X1 U6130 ( .B1(n9356), .B2(n5136), .A(n5247), .ZN(n5246) );
  NAND2_X1 U6131 ( .A1(n6647), .A2(n6646), .ZN(n9441) );
  NAND2_X1 U6132 ( .A1(n5719), .A2(n6642), .ZN(n9336) );
  NAND2_X1 U6133 ( .A1(n9356), .A2(n9357), .ZN(n5719) );
  NAND2_X1 U6134 ( .A1(n6636), .A2(n6635), .ZN(n9448) );
  NAND2_X1 U6135 ( .A1(n6623), .A2(n6622), .ZN(n9385) );
  NAND2_X1 U6136 ( .A1(n5731), .A2(n5146), .ZN(n6606) );
  NAND2_X1 U6137 ( .A1(n6552), .A2(n6551), .ZN(n8479) );
  NAND2_X1 U6138 ( .A1(n8124), .A2(n8910), .ZN(n8154) );
  INV_X1 U6139 ( .A(n8012), .ZN(n7806) );
  NAND2_X1 U6140 ( .A1(n7834), .A2(n8901), .ZN(n7795) );
  NAND2_X1 U6141 ( .A1(n8620), .A2(n7969), .ZN(n9320) );
  OR2_X1 U6142 ( .A1(n6493), .A2(n7133), .ZN(n6474) );
  INV_X1 U6143 ( .A(n6473), .ZN(n5242) );
  INV_X1 U6144 ( .A(n9317), .ZN(n9364) );
  INV_X1 U6145 ( .A(n9380), .ZN(n9314) );
  NAND2_X1 U6146 ( .A1(n9465), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5740) );
  NAND2_X1 U6147 ( .A1(n6563), .A2(n5337), .ZN(n8321) );
  NAND2_X1 U6148 ( .A1(n7162), .A2(n8838), .ZN(n5337) );
  INV_X1 U6149 ( .A(n8845), .ZN(n9474) );
  AND2_X1 U6150 ( .A1(n6785), .A2(n6784), .ZN(n9478) );
  NAND2_X1 U6151 ( .A1(n9392), .A2(n5742), .ZN(n9475) );
  NAND2_X1 U6152 ( .A1(n5124), .A2(n9414), .ZN(n5742) );
  INV_X1 U6153 ( .A(n6832), .ZN(n9486) );
  INV_X1 U6154 ( .A(n8685), .ZN(n9490) );
  INV_X1 U6155 ( .A(n8991), .ZN(n9494) );
  INV_X1 U6156 ( .A(n8663), .ZN(n9498) );
  AND2_X1 U6157 ( .A1(n6542), .A2(n6541), .ZN(n8290) );
  AND2_X1 U6158 ( .A1(n6533), .A2(n6532), .ZN(n8931) );
  INV_X1 U6159 ( .A(n6812), .ZN(n7970) );
  NAND2_X1 U6160 ( .A1(n7513), .A2(n7144), .ZN(n7157) );
  NAND2_X1 U6161 ( .A1(n6441), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6428) );
  NOR2_X1 U6162 ( .A1(n5369), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8609) );
  INV_X1 U6163 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8061) );
  INV_X1 U6164 ( .A(n9028), .ZN(n8060) );
  INV_X1 U6165 ( .A(n7476), .ZN(n7892) );
  INV_X1 U6166 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7847) );
  INV_X1 U6167 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7826) );
  INV_X1 U6168 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7609) );
  INV_X1 U6169 ( .A(n8554), .ZN(n9118) );
  INV_X1 U6170 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7397) );
  INV_X1 U6171 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n7188) );
  INV_X1 U6172 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n7167) );
  INV_X1 U6173 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n7159) );
  INV_X1 U6174 ( .A(n7287), .ZN(n7637) );
  INV_X1 U6175 ( .A(n6455), .ZN(n6457) );
  CLKBUF_X1 U6176 ( .A(n7207), .Z(n5231) );
  XNOR2_X1 U6177 ( .A(n6390), .B(n10835), .ZN(n8114) );
  INV_X1 U6178 ( .A(n6959), .ZN(n8137) );
  AND4_X1 U6179 ( .A1(n6061), .A2(n6060), .A3(n6059), .A4(n6058), .ZN(n9545)
         );
  AND2_X1 U6180 ( .A1(n6974), .A2(n6973), .ZN(n6975) );
  AND2_X1 U6181 ( .A1(n5618), .A2(n5205), .ZN(n9551) );
  INV_X1 U6182 ( .A(n8108), .ZN(n11104) );
  NAND2_X1 U6183 ( .A1(n9609), .A2(n7079), .ZN(n9578) );
  NAND2_X1 U6184 ( .A1(n5615), .A2(n5609), .ZN(n5606) );
  NAND2_X1 U6185 ( .A1(n5893), .A2(n5892), .ZN(n10398) );
  OAI22_X1 U6186 ( .A1(n11056), .A2(n5129), .B1(n5269), .B2(n8704), .ZN(n7984)
         );
  NAND2_X1 U6187 ( .A1(n5631), .A2(n5632), .ZN(n7983) );
  INV_X1 U6188 ( .A(n9697), .ZN(n9676) );
  AND4_X1 U6189 ( .A1(n5881), .A2(n5880), .A3(n5879), .A4(n5878), .ZN(n10273)
         );
  NAND2_X1 U6190 ( .A1(n6185), .A2(n6184), .ZN(n10237) );
  AND2_X1 U6191 ( .A1(n9601), .A2(n5621), .ZN(n9665) );
  NAND2_X1 U6192 ( .A1(n9601), .A2(n7036), .ZN(n5624) );
  NAND2_X1 U6193 ( .A1(n5626), .A2(n5629), .ZN(n5625) );
  INV_X1 U6194 ( .A(n9646), .ZN(n9689) );
  INV_X1 U6195 ( .A(n9644), .ZN(n9687) );
  INV_X1 U6196 ( .A(n9691), .ZN(n9678) );
  OR2_X1 U6197 ( .A1(n7120), .A2(n8497), .ZN(n9691) );
  OR3_X1 U6198 ( .A1(n7116), .A2(n9701), .A3(n7113), .ZN(n9697) );
  AND4_X1 U6199 ( .A1(n6299), .A2(n6298), .A3(n6297), .A4(n6296), .ZN(n10316)
         );
  NAND2_X1 U6200 ( .A1(n10130), .A2(n9994), .ZN(n5404) );
  NAND2_X1 U6201 ( .A1(n5406), .A2(n10411), .ZN(n5405) );
  XNOR2_X1 U6202 ( .A(n6348), .B(n9800), .ZN(n5406) );
  AND4_X1 U6203 ( .A1(n6286), .A2(n6285), .A3(n6284), .A4(n6283), .ZN(n10174)
         );
  AND4_X1 U6204 ( .A1(n6268), .A2(n6267), .A3(n6266), .A4(n6265), .ZN(n10317)
         );
  NAND2_X1 U6205 ( .A1(n6240), .A2(n6239), .ZN(n10192) );
  AND4_X1 U6206 ( .A1(n6229), .A2(n6228), .A3(n6227), .A4(n6226), .ZN(n10217)
         );
  NAND2_X1 U6207 ( .A1(n5708), .A2(n6193), .ZN(n10213) );
  NAND2_X1 U6208 ( .A1(n6206), .A2(n6205), .ZN(n10222) );
  OAI21_X1 U6209 ( .B1(n10280), .B2(n5280), .A(n5278), .ZN(n10250) );
  OAI21_X1 U6210 ( .B1(n10280), .B2(n5283), .A(n9770), .ZN(n10260) );
  INV_X1 U6211 ( .A(n9562), .ZN(n10376) );
  NOR2_X1 U6212 ( .A1(n5407), .A2(n5409), .ZN(n10278) );
  INV_X1 U6213 ( .A(n5408), .ZN(n5407) );
  NAND2_X1 U6214 ( .A1(n8535), .A2(n9920), .ZN(n10295) );
  NAND2_X1 U6215 ( .A1(n5285), .A2(n5166), .ZN(n10396) );
  AND2_X1 U6216 ( .A1(n5285), .A2(n5144), .ZN(n8489) );
  NAND2_X1 U6217 ( .A1(n8197), .A2(n9892), .ZN(n8353) );
  AND4_X1 U6218 ( .A1(n5913), .A2(n5912), .A3(n5911), .A4(n5910), .ZN(n9692)
         );
  NAND2_X1 U6219 ( .A1(n7882), .A2(n9869), .ZN(n7908) );
  OAI21_X1 U6220 ( .B1(n7713), .B2(n5696), .A(n5693), .ZN(n7722) );
  NAND2_X1 U6221 ( .A1(n7712), .A2(n6037), .ZN(n7723) );
  AND4_X1 U6222 ( .A1(n6049), .A2(n6048), .A3(n6047), .A4(n6046), .ZN(n7962)
         );
  NAND2_X1 U6223 ( .A1(n7548), .A2(n5995), .ZN(n7680) );
  INV_X1 U6224 ( .A(n10309), .ZN(n11075) );
  NAND2_X1 U6225 ( .A1(n7111), .A2(n10468), .ZN(n7919) );
  INV_X1 U6226 ( .A(n11072), .ZN(n10223) );
  INV_X1 U6227 ( .A(n10135), .ZN(n10430) );
  INV_X1 U6228 ( .A(n10192), .ZN(n10441) );
  INV_X1 U6229 ( .A(n10237), .ZN(n10453) );
  AND2_X1 U6230 ( .A1(n6016), .A2(n6015), .ZN(n11073) );
  INV_X1 U6231 ( .A(n7923), .ZN(n6009) );
  INV_X1 U6232 ( .A(n7694), .ZN(n8074) );
  XNOR2_X1 U6233 ( .A(n8608), .B(n8607), .ZN(n10477) );
  OAI21_X1 U6234 ( .B1(n8629), .B2(n8628), .A(n8603), .ZN(n8608) );
  NAND2_X1 U6235 ( .A1(n5867), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5868) );
  OAI21_X1 U6236 ( .B1(n5866), .B2(n6098), .A(P1_IR_REG_29__SCAN_IN), .ZN(
        n5869) );
  INV_X1 U6237 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n10775) );
  NAND2_X1 U6238 ( .A1(n6363), .A2(n6368), .ZN(n8244) );
  AND2_X1 U6239 ( .A1(n5369), .A2(P1_U3086), .ZN(n10476) );
  INV_X1 U6240 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7850) );
  NAND2_X1 U6241 ( .A1(n6365), .A2(n6323), .ZN(n7848) );
  INV_X1 U6242 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8723) );
  INV_X1 U6243 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7794) );
  INV_X1 U6244 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10593) );
  INV_X1 U6245 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n7169) );
  INV_X1 U6246 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10595) );
  INV_X1 U6247 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10795) );
  INV_X1 U6248 ( .A(n5237), .ZN(n7853) );
  INV_X1 U6249 ( .A(n5430), .ZN(n7856) );
  INV_X1 U6250 ( .A(n5439), .ZN(n8170) );
  AOI211_X1 U6251 ( .C1(n9157), .C2(n8592), .A(n8591), .B(n8590), .ZN(n8593)
         );
  INV_X1 U6252 ( .A(n6846), .ZN(n8621) );
  NAND2_X1 U6253 ( .A1(n5741), .A2(n5738), .ZN(P2_U3487) );
  INV_X1 U6254 ( .A(n5739), .ZN(n5738) );
  NAND2_X1 U6255 ( .A1(n9475), .A2(n9456), .ZN(n5741) );
  OAI21_X1 U6256 ( .B1(n9478), .B2(n9432), .A(n5740), .ZN(n5739) );
  INV_X1 U6257 ( .A(n5392), .ZN(n10311) );
  AOI21_X1 U6258 ( .B1(n10423), .B2(n11110), .A(n5393), .ZN(n5392) );
  NOR2_X1 U6259 ( .A1(n11110), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n5393) );
  NOR2_X1 U6260 ( .A1(n6396), .A2(n5753), .ZN(n6397) );
  XNOR2_X1 U6261 ( .A(n6388), .B(n6387), .ZN(n6918) );
  NAND2_X1 U6262 ( .A1(n8970), .A2(n9437), .ZN(n5133) );
  AND2_X1 U6263 ( .A1(n5402), .A2(n5401), .ZN(n5134) );
  NAND2_X1 U6264 ( .A1(n9047), .A2(n7806), .ZN(n5135) );
  AND2_X1 U6265 ( .A1(n9346), .A2(n5720), .ZN(n5136) );
  AND2_X1 U6266 ( .A1(n9787), .A2(n5156), .ZN(n5137) );
  INV_X1 U6267 ( .A(n6823), .ZN(n9330) );
  NAND2_X1 U6268 ( .A1(n8967), .A2(n9338), .ZN(n5138) );
  AND2_X1 U6269 ( .A1(n5135), .A2(n5152), .ZN(n5139) );
  AND2_X1 U6270 ( .A1(n7569), .A2(n11024), .ZN(n5140) );
  NAND2_X1 U6271 ( .A1(n6278), .A2(n6277), .ZN(n10157) );
  AOI22_X1 U6272 ( .A1(n10477), .A2(n8838), .B1(n8837), .B2(
        P1_DATAO_REG_31__SCAN_IN), .ZN(n9470) );
  AND2_X1 U6273 ( .A1(n5699), .A2(n9996), .ZN(n5141) );
  AND2_X1 U6274 ( .A1(n7134), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5142) );
  INV_X1 U6275 ( .A(n9695), .ZN(n10409) );
  NAND2_X1 U6276 ( .A1(n5900), .A2(n5899), .ZN(n9695) );
  NAND2_X1 U6277 ( .A1(n6846), .A2(n8016), .ZN(n5143) );
  OR2_X1 U6278 ( .A1(n9695), .A2(n5697), .ZN(n5144) );
  INV_X1 U6279 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5867) );
  AND2_X1 U6280 ( .A1(n5704), .A2(n5286), .ZN(n5145) );
  AND2_X1 U6281 ( .A1(n6166), .A2(n6165), .ZN(n10368) );
  INV_X1 U6282 ( .A(n10368), .ZN(n10263) );
  INV_X1 U6283 ( .A(n9280), .ZN(n5379) );
  OR2_X1 U6284 ( .A1(n8339), .A2(n8402), .ZN(n5146) );
  AND2_X1 U6285 ( .A1(n8339), .A2(n8402), .ZN(n5147) );
  INV_X1 U6286 ( .A(n10819), .ZN(n5456) );
  NOR2_X2 U6287 ( .A1(n8634), .A2(n5871), .ZN(n5970) );
  XOR2_X1 U6288 ( .A(n9182), .B(n8694), .Z(n5148) );
  INV_X2 U6289 ( .A(n6086), .ZN(n6167) );
  AND2_X1 U6290 ( .A1(n5552), .A2(n8769), .ZN(n5149) );
  NAND2_X1 U6291 ( .A1(n10200), .A2(n5396), .ZN(n5150) );
  NAND2_X1 U6292 ( .A1(n6851), .A2(n6425), .ZN(n5151) );
  NAND2_X1 U6293 ( .A1(n9048), .A2(n8040), .ZN(n5152) );
  AND2_X1 U6294 ( .A1(n10200), .A2(n10445), .ZN(n5153) );
  INV_X1 U6295 ( .A(n9357), .ZN(n5721) );
  OR2_X1 U6296 ( .A1(n8183), .A2(n8166), .ZN(n5154) );
  AND2_X1 U6297 ( .A1(n7009), .A2(n9519), .ZN(n5155) );
  INV_X1 U6298 ( .A(n9663), .ZN(n5698) );
  OR2_X1 U6299 ( .A1(n8207), .A2(n10415), .ZN(n5156) );
  INV_X1 U6300 ( .A(n6588), .ZN(n6590) );
  INV_X1 U6301 ( .A(n8919), .ZN(n6815) );
  INV_X1 U6302 ( .A(n7244), .ZN(n7271) );
  NAND2_X1 U6303 ( .A1(n9277), .A2(n6703), .ZN(n9235) );
  OR2_X1 U6304 ( .A1(n7867), .A2(n7852), .ZN(n5157) );
  INV_X1 U6305 ( .A(n8999), .ZN(n5657) );
  INV_X1 U6306 ( .A(n9919), .ZN(n5410) );
  XNOR2_X1 U6307 ( .A(n5725), .B(P2_IR_REG_30__SCAN_IN), .ZN(n6431) );
  OR2_X1 U6308 ( .A1(n8968), .A2(n8966), .ZN(n5158) );
  NAND2_X1 U6309 ( .A1(n8330), .A2(n9042), .ZN(n5159) );
  AND2_X1 U6310 ( .A1(n5632), .A2(n5630), .ZN(n5160) );
  NAND2_X1 U6311 ( .A1(n8515), .A2(n9039), .ZN(n5161) );
  INV_X1 U6312 ( .A(n6952), .ZN(n5637) );
  NAND2_X1 U6313 ( .A1(n6424), .A2(n6590), .ZN(n6808) );
  OR2_X1 U6314 ( .A1(n8492), .A2(n10389), .ZN(n5162) );
  AND2_X1 U6315 ( .A1(n5624), .A2(n7038), .ZN(n5163) );
  AND3_X1 U6316 ( .A1(n5317), .A2(n5316), .A3(n5315), .ZN(n5164) );
  INV_X1 U6317 ( .A(n5675), .ZN(n5673) );
  NOR2_X1 U6318 ( .A1(n5887), .A2(n5676), .ZN(n5675) );
  AND2_X1 U6319 ( .A1(n5714), .A2(n5726), .ZN(n5165) );
  AND2_X1 U6320 ( .A1(n9771), .A2(n5144), .ZN(n5166) );
  AND3_X1 U6321 ( .A1(n6519), .A2(n6518), .A3(n6517), .ZN(n8160) );
  AND4_X1 U6322 ( .A1(n6592), .A2(n6420), .A3(n6804), .A4(n6419), .ZN(n5167)
         );
  AND2_X1 U6323 ( .A1(n8638), .A2(n9340), .ZN(n5168) );
  NOR2_X1 U6324 ( .A1(n8546), .A2(n9091), .ZN(n5169) );
  AND2_X1 U6325 ( .A1(n8127), .A2(n8012), .ZN(n5170) );
  NOR2_X1 U6326 ( .A1(n9096), .A2(n8583), .ZN(n5171) );
  OR2_X1 U6327 ( .A1(n11104), .A2(n7914), .ZN(n5172) );
  INV_X1 U6328 ( .A(n8530), .ZN(n10390) );
  NAND2_X1 U6329 ( .A1(n6116), .A2(n6115), .ZN(n8530) );
  INV_X1 U6330 ( .A(n5662), .ZN(n5661) );
  NOR2_X1 U6331 ( .A1(n6831), .A2(n5663), .ZN(n5662) );
  INV_X1 U6332 ( .A(n5529), .ZN(n5528) );
  OAI21_X1 U6333 ( .B1(n5531), .B2(n5530), .A(n8724), .ZN(n5529) );
  NAND2_X1 U6334 ( .A1(n10379), .A2(n10265), .ZN(n5173) );
  INV_X1 U6335 ( .A(n5784), .ZN(n5354) );
  OR2_X1 U6336 ( .A1(n6113), .A2(n5650), .ZN(n5174) );
  NAND2_X1 U6337 ( .A1(n7229), .A2(n8623), .ZN(n5175) );
  INV_X1 U6338 ( .A(n5545), .ZN(n5544) );
  NAND2_X1 U6339 ( .A1(n5549), .A2(n5548), .ZN(n5545) );
  AND2_X1 U6340 ( .A1(n5752), .A2(n6193), .ZN(n5176) );
  AND2_X1 U6341 ( .A1(n9291), .A2(n6681), .ZN(n5177) );
  AND2_X1 U6342 ( .A1(n9833), .A2(n6333), .ZN(n5178) );
  AND2_X1 U6343 ( .A1(n5410), .A2(n9920), .ZN(n5179) );
  OR2_X1 U6344 ( .A1(n9672), .A2(n9673), .ZN(n5180) );
  NAND2_X1 U6345 ( .A1(n5501), .A2(n5503), .ZN(n5504) );
  AND2_X1 U6346 ( .A1(n10368), .A2(n10376), .ZN(n5181) );
  NOR2_X1 U6347 ( .A1(n9137), .A2(n8586), .ZN(n5182) );
  OR2_X1 U6348 ( .A1(n8698), .A2(n9189), .ZN(n6834) );
  AND2_X1 U6349 ( .A1(n9441), .A2(n9325), .ZN(n5183) );
  AND2_X1 U6350 ( .A1(n9311), .A2(n8966), .ZN(n5184) );
  INV_X1 U6351 ( .A(n5729), .ZN(n5728) );
  NAND2_X1 U6352 ( .A1(n6733), .A2(n5730), .ZN(n5729) );
  NAND2_X1 U6353 ( .A1(n7036), .A2(n9666), .ZN(n5185) );
  INV_X1 U6354 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5863) );
  AND3_X1 U6355 ( .A1(n5938), .A2(n5939), .A3(n5940), .ZN(n5186) );
  OR2_X1 U6356 ( .A1(n9470), .A2(n9172), .ZN(n5187) );
  AND2_X1 U6357 ( .A1(n5804), .A2(SI_13_), .ZN(n5188) );
  INV_X1 U6358 ( .A(n5397), .ZN(n5396) );
  NAND2_X1 U6359 ( .A1(n5399), .A2(n5398), .ZN(n5397) );
  AND2_X1 U6360 ( .A1(n9311), .A2(n8968), .ZN(n5189) );
  INV_X1 U6361 ( .A(n5421), .ZN(n5420) );
  NAND2_X1 U6362 ( .A1(n10198), .A2(n9943), .ZN(n5421) );
  INV_X1 U6363 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6321) );
  NAND2_X1 U6364 ( .A1(n6739), .A2(n6738), .ZN(n5190) );
  AND4_X1 U6365 ( .A1(n6464), .A2(n6463), .A3(n6462), .A4(n6461), .ZN(n7486)
         );
  NOR2_X1 U6366 ( .A1(n10418), .A2(n9692), .ZN(n5191) );
  AOI21_X1 U6367 ( .B1(n5714), .B2(n5717), .A(n5713), .ZN(n5712) );
  AND2_X1 U6368 ( .A1(n5721), .A2(n8956), .ZN(n5192) );
  AND2_X1 U6369 ( .A1(n6431), .A2(n9515), .ZN(n6465) );
  OR2_X1 U6370 ( .A1(n5687), .A2(n9308), .ZN(n5193) );
  INV_X1 U6371 ( .A(n9295), .ZN(n9291) );
  XNOR2_X1 U6372 ( .A(n9298), .B(n9304), .ZN(n9295) );
  AND2_X1 U6373 ( .A1(n9558), .A2(n9559), .ZN(n5194) );
  AND2_X1 U6374 ( .A1(n5245), .A2(n5243), .ZN(n5195) );
  INV_X1 U6375 ( .A(n8731), .ZN(n8646) );
  INV_X1 U6376 ( .A(n8901), .ZN(n5375) );
  AOI22_X1 U6377 ( .A1(n9013), .A2(n9189), .B1(n9018), .B2(n9478), .ZN(n9009)
         );
  AND2_X1 U6378 ( .A1(n10209), .A2(n9943), .ZN(n5196) );
  AND2_X1 U6379 ( .A1(n9928), .A2(n9921), .ZN(n5197) );
  INV_X1 U6380 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n6329) );
  AND2_X1 U6381 ( .A1(n5148), .A2(n5528), .ZN(n5198) );
  AND2_X1 U6382 ( .A1(n5330), .A2(n5327), .ZN(n5199) );
  AND2_X1 U6383 ( .A1(n5778), .A2(n5784), .ZN(n5200) );
  AND2_X1 U6384 ( .A1(n6287), .A2(n6269), .ZN(n5201) );
  AND2_X1 U6385 ( .A1(n7896), .A2(n5747), .ZN(n5202) );
  INV_X1 U6386 ( .A(n6521), .ZN(n5254) );
  NAND2_X1 U6387 ( .A1(n10470), .A2(n6098), .ZN(n5203) );
  AND2_X1 U6388 ( .A1(n5192), .A2(n5293), .ZN(n5204) );
  AND2_X1 U6389 ( .A1(n5611), .A2(n9579), .ZN(n5610) );
  INV_X1 U6390 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n10470) );
  NAND2_X1 U6391 ( .A1(n7439), .A2(n11044), .ZN(n5995) );
  INV_X1 U6392 ( .A(n9547), .ZN(n5700) );
  NAND2_X1 U6393 ( .A1(n6260), .A2(n6259), .ZN(n10178) );
  INV_X1 U6394 ( .A(n10178), .ZN(n5398) );
  NAND2_X1 U6395 ( .A1(n8312), .A2(n8920), .ZN(n8326) );
  NAND2_X1 U6396 ( .A1(n5388), .A2(n5721), .ZN(n9306) );
  INV_X1 U6397 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5684) );
  NAND2_X1 U6398 ( .A1(n6292), .A2(n6291), .ZN(n8718) );
  XNOR2_X1 U6399 ( .A(n6332), .B(n11034), .ZN(n7572) );
  INV_X1 U6400 ( .A(n7572), .ZN(n5416) );
  INV_X1 U6401 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5368) );
  NAND2_X1 U6402 ( .A1(n6132), .A2(n6131), .ZN(n10385) );
  INV_X1 U6403 ( .A(n10385), .ZN(n10305) );
  NAND2_X1 U6404 ( .A1(n5623), .A2(n9666), .ZN(n5205) );
  AND2_X1 U6405 ( .A1(n9290), .A2(n6693), .ZN(n5206) );
  NAND2_X1 U6406 ( .A1(n5846), .A2(n5845), .ZN(n6079) );
  AND2_X1 U6407 ( .A1(n9433), .A2(n9324), .ZN(n5207) );
  NAND2_X1 U6408 ( .A1(n8527), .A2(n5134), .ZN(n5403) );
  AND2_X1 U6409 ( .A1(n10813), .A2(n10812), .ZN(n5208) );
  AND2_X1 U6410 ( .A1(n5723), .A2(n6681), .ZN(n5209) );
  OR2_X1 U6411 ( .A1(n6113), .A2(n6112), .ZN(n5210) );
  AND2_X1 U6412 ( .A1(n8693), .A2(n9034), .ZN(n5211) );
  OR2_X1 U6413 ( .A1(n10316), .A2(n10388), .ZN(n5212) );
  AND2_X1 U6414 ( .A1(n8103), .A2(n9891), .ZN(n5213) );
  INV_X1 U6415 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6536) );
  INV_X1 U6416 ( .A(n8579), .ZN(n5497) );
  NAND2_X1 U6417 ( .A1(n6155), .A2(n6154), .ZN(n10379) );
  INV_X1 U6418 ( .A(n10379), .ZN(n5401) );
  INV_X1 U6419 ( .A(n9852), .ZN(n5695) );
  NAND2_X1 U6420 ( .A1(n5250), .A2(n5252), .ZN(n8148) );
  INV_X1 U6421 ( .A(n8558), .ZN(n9081) );
  NAND2_X1 U6422 ( .A1(n6581), .A2(n6580), .ZN(n6595) );
  XNOR2_X1 U6423 ( .A(n6366), .B(P1_IR_REG_24__SCAN_IN), .ZN(n6386) );
  NOR2_X1 U6424 ( .A1(n8184), .A2(n8185), .ZN(n5214) );
  INV_X1 U6425 ( .A(SI_22_), .ZN(n5492) );
  AND2_X1 U6426 ( .A1(n5639), .A2(n5629), .ZN(n5215) );
  AND2_X1 U6427 ( .A1(n5734), .A2(n5152), .ZN(n5216) );
  INV_X1 U6428 ( .A(n6838), .ZN(n7193) );
  AND4_X1 U6429 ( .A1(n5907), .A2(n5906), .A3(n5905), .A4(n5904), .ZN(n9523)
         );
  INV_X1 U6430 ( .A(n9523), .ZN(n5697) );
  XOR2_X1 U6431 ( .A(n10773), .B(keyinput_200), .Z(n5217) );
  AND2_X2 U6432 ( .A1(n6408), .A2(n6407), .ZN(n11110) );
  NAND2_X1 U6433 ( .A1(n6370), .A2(n5853), .ZN(n6351) );
  NAND2_X1 U6434 ( .A1(n10783), .A2(n10782), .ZN(n5218) );
  XOR2_X1 U6435 ( .A(n6432), .B(n5467), .Z(n5219) );
  AND2_X1 U6436 ( .A1(n5496), .A2(n7289), .ZN(n5220) );
  XNOR2_X1 U6437 ( .A(n6807), .B(P2_IR_REG_20__SCAN_IN), .ZN(n6897) );
  NOR2_X1 U6438 ( .A1(n10832), .A2(n10831), .ZN(n5221) );
  AND2_X1 U6439 ( .A1(n5431), .A2(n5435), .ZN(n5222) );
  NAND3_X1 U6440 ( .A1(n10826), .A2(n10825), .A3(n10824), .ZN(n5223) );
  INV_X1 U6441 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10789) );
  AND2_X1 U6442 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(keyinput_215), .ZN(n5224)
         );
  XNOR2_X1 U6443 ( .A(n8545), .B(n9103), .ZN(n9092) );
  XNOR2_X1 U6444 ( .A(n8582), .B(n9103), .ZN(n9097) );
  OAI21_X2 U6445 ( .B1(n8504), .B2(n8947), .A(n8946), .ZN(n9369) );
  NAND2_X1 U6446 ( .A1(n10957), .A2(n7199), .ZN(n7200) );
  NOR2_X1 U6447 ( .A1(n10980), .A2(n10979), .ZN(n10978) );
  OAI21_X1 U6448 ( .B1(n7240), .B2(n7271), .A(n7279), .ZN(n5427) );
  NOR2_X1 U6449 ( .A1(n9065), .A2(n8544), .ZN(n9075) );
  NOR2_X1 U6450 ( .A1(n9073), .A2(n5227), .ZN(n8545) );
  NOR2_X1 U6451 ( .A1(n8542), .A2(n5236), .ZN(n8543) );
  XNOR2_X1 U6452 ( .A(n8543), .B(n8579), .ZN(n9066) );
  NAND2_X1 U6453 ( .A1(n5433), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5432) );
  NOR2_X1 U6454 ( .A1(n5427), .A2(n8018), .ZN(n7281) );
  NOR2_X1 U6455 ( .A1(n9127), .A2(n8549), .ZN(n8551) );
  NOR2_X1 U6456 ( .A1(n11002), .A2(n8256), .ZN(n8258) );
  OAI22_X1 U6457 ( .A1(n6453), .A2(n6454), .B1(P2_IR_REG_2__SCAN_IN), .B2(
        P2_IR_REG_31__SCAN_IN), .ZN(n6455) );
  INV_X1 U6458 ( .A(n9111), .ZN(n5239) );
  NAND2_X1 U6459 ( .A1(n5182), .A2(n8588), .ZN(n8589) );
  NOR2_X1 U6460 ( .A1(n9135), .A2(n8552), .ZN(n9137) );
  NAND2_X1 U6461 ( .A1(n8583), .A2(n5511), .ZN(n5509) );
  NOR2_X1 U6462 ( .A1(n9058), .A2(n8580), .ZN(n9084) );
  XNOR2_X1 U6463 ( .A(n8270), .B(n10998), .ZN(n11000) );
  NOR2_X1 U6464 ( .A1(n11000), .A2(n11001), .ZN(n10999) );
  NAND2_X1 U6465 ( .A1(n9620), .A2(n9621), .ZN(n9619) );
  NAND2_X1 U6466 ( .A1(n5618), .A2(n5617), .ZN(n9550) );
  XNOR2_X1 U6467 ( .A(n6948), .B(n6950), .ZN(n5635) );
  NAND3_X1 U6468 ( .A1(n9193), .A2(n9003), .A3(n9192), .ZN(n6833) );
  NAND2_X2 U6469 ( .A1(n5777), .A2(n5776), .ZN(n6025) );
  NAND2_X2 U6470 ( .A1(n9296), .A2(n9295), .ZN(n9428) );
  NAND2_X1 U6471 ( .A1(n6845), .A2(n5268), .ZN(n8614) );
  INV_X1 U6472 ( .A(n8614), .ZN(n6848) );
  AND2_X2 U6473 ( .A1(n8901), .A2(n8906), .ZN(n8897) );
  INV_X1 U6474 ( .A(n9355), .ZN(n5388) );
  NAND2_X1 U6475 ( .A1(n9269), .A2(n9268), .ZN(n9271) );
  NAND2_X1 U6476 ( .A1(n9258), .A2(n6829), .ZN(n5384) );
  NAND2_X1 U6477 ( .A1(n8124), .A2(n5385), .ZN(n8152) );
  AOI21_X1 U6478 ( .B1(n5381), .B2(n8879), .A(n8878), .ZN(n8880) );
  OAI21_X1 U6479 ( .B1(n5374), .B2(n8901), .A(n8909), .ZN(n5371) );
  AOI21_X1 U6480 ( .B1(n8871), .B2(n9003), .A(n8873), .ZN(n5383) );
  NOR2_X1 U6481 ( .A1(n9128), .A2(n9129), .ZN(n9127) );
  NAND2_X1 U6482 ( .A1(n5434), .A2(n7223), .ZN(n5433) );
  INV_X1 U6483 ( .A(n10944), .ZN(n5232) );
  NOR2_X1 U6484 ( .A1(n8258), .A2(n8257), .ZN(n8542) );
  AOI22_X2 U6485 ( .A1(n7225), .A2(n7224), .B1(n7223), .B2(n7222), .ZN(n10987)
         );
  NAND2_X1 U6486 ( .A1(n8546), .A2(n5442), .ZN(n5440) );
  NAND2_X1 U6487 ( .A1(n10965), .A2(n10966), .ZN(n10964) );
  NAND2_X1 U6488 ( .A1(n8185), .A2(n5508), .ZN(n5506) );
  NOR2_X1 U6489 ( .A1(n9075), .A2(n9074), .ZN(n9073) );
  XNOR2_X1 U6490 ( .A(n5240), .B(n6835), .ZN(n6810) );
  NAND2_X1 U6491 ( .A1(n5734), .A2(n5251), .ZN(n5250) );
  NAND3_X1 U6494 ( .A1(n6445), .A2(n5554), .A3(n6560), .ZN(n6588) );
  NAND2_X2 U6495 ( .A1(n6837), .A2(n6838), .ZN(n7130) );
  NAND2_X2 U6496 ( .A1(n5186), .A2(n5937), .ZN(n10001) );
  NAND3_X1 U6497 ( .A1(n5744), .A2(n5860), .A3(n5867), .ZN(n10474) );
  NAND3_X1 U6498 ( .A1(n5860), .A2(n5744), .A3(n5273), .ZN(n5272) );
  AND2_X4 U6499 ( .A1(n8541), .A2(n8634), .ZN(n6066) );
  NAND2_X1 U6500 ( .A1(n10280), .A2(n5278), .ZN(n5277) );
  NAND2_X1 U6501 ( .A1(n5703), .A2(n5145), .ZN(n5285) );
  NAND2_X1 U6502 ( .A1(n5703), .A2(n5704), .ZN(n8455) );
  INV_X1 U6503 ( .A(n5285), .ZN(n8454) );
  INV_X1 U6504 ( .A(n9789), .ZN(n5286) );
  NAND2_X1 U6505 ( .A1(n6006), .A2(n6005), .ZN(n5289) );
  NAND2_X1 U6506 ( .A1(n5991), .A2(n5990), .ZN(n5290) );
  NAND2_X1 U6507 ( .A1(n8945), .A2(n8950), .ZN(n5291) );
  OR2_X1 U6508 ( .A1(n8945), .A2(n5296), .ZN(n5295) );
  NAND2_X1 U6509 ( .A1(n5299), .A2(n5292), .ZN(n8960) );
  NAND2_X1 U6510 ( .A1(n5299), .A2(n5300), .ZN(n8954) );
  NAND2_X1 U6511 ( .A1(n9017), .A2(n9016), .ZN(n9022) );
  NAND2_X1 U6512 ( .A1(n5304), .A2(n9009), .ZN(n5303) );
  INV_X1 U6513 ( .A(n5307), .ZN(n5304) );
  NAND2_X1 U6514 ( .A1(n5306), .A2(n9008), .ZN(n5305) );
  NAND2_X1 U6515 ( .A1(n5307), .A2(n9010), .ZN(n5306) );
  NAND2_X1 U6516 ( .A1(n9006), .A2(n9005), .ZN(n5307) );
  INV_X1 U6517 ( .A(n8970), .ZN(n5323) );
  NAND2_X1 U6518 ( .A1(n8915), .A2(n9007), .ZN(n5328) );
  NAND4_X1 U6519 ( .A1(n5329), .A2(n5328), .A3(n5332), .A4(n5199), .ZN(n5326)
         );
  NAND2_X1 U6520 ( .A1(n8917), .A2(n9007), .ZN(n5332) );
  AND2_X1 U6521 ( .A1(n5331), .A2(n6815), .ZN(n5330) );
  AOI21_X2 U6522 ( .B1(n5334), .B2(n6847), .A(n5339), .ZN(n9026) );
  NAND2_X1 U6523 ( .A1(n5335), .A2(n5340), .ZN(n5334) );
  NAND2_X1 U6524 ( .A1(n5336), .A2(n5187), .ZN(n5335) );
  NAND2_X1 U6525 ( .A1(n9024), .A2(n9023), .ZN(n5336) );
  INV_X2 U6526 ( .A(n5768), .ZN(n7134) );
  NAND2_X2 U6527 ( .A1(n5686), .A2(n5685), .ZN(n5768) );
  MUX2_X1 U6528 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n7134), .Z(n5766) );
  OR2_X2 U6529 ( .A1(n6078), .A2(n5346), .ZN(n5343) );
  OAI21_X1 U6530 ( .B1(n6078), .B2(n5802), .A(n5801), .ZN(n6096) );
  NAND3_X1 U6531 ( .A1(n8877), .A2(n8875), .A3(n9018), .ZN(n9013) );
  NAND2_X1 U6532 ( .A1(n6025), .A2(n5200), .ZN(n5350) );
  NAND2_X1 U6533 ( .A1(n6025), .A2(n5778), .ZN(n5357) );
  NAND2_X1 U6534 ( .A1(n5350), .A2(n5352), .ZN(n5791) );
  NAND2_X1 U6535 ( .A1(n6255), .A2(n5362), .ZN(n5360) );
  OAI21_X1 U6536 ( .B1(n5369), .B2(n5368), .A(n5367), .ZN(n5769) );
  MUX2_X1 U6537 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n5768), .Z(n5772) );
  MUX2_X1 U6538 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n5768), .Z(n5775) );
  MUX2_X1 U6539 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n5369), .Z(n5779) );
  MUX2_X1 U6540 ( .A(n7159), .B(n10795), .S(n5369), .Z(n5781) );
  MUX2_X1 U6541 ( .A(n5785), .B(n10595), .S(n5369), .Z(n5787) );
  MUX2_X1 U6542 ( .A(n7167), .B(n7169), .S(n5369), .Z(n5793) );
  MUX2_X1 U6543 ( .A(n7188), .B(n10792), .S(n5369), .Z(n5796) );
  OAI21_X1 U6544 ( .B1(n7835), .B2(n5375), .A(n5373), .ZN(n8122) );
  NAND2_X1 U6545 ( .A1(n5372), .A2(n5370), .ZN(n6814) );
  INV_X1 U6546 ( .A(n5371), .ZN(n5370) );
  NAND2_X1 U6547 ( .A1(n7835), .A2(n5373), .ZN(n5372) );
  INV_X1 U6548 ( .A(n5374), .ZN(n5373) );
  OAI21_X1 U6549 ( .B1(n9428), .B2(n5379), .A(n5376), .ZN(n9269) );
  OAI21_X2 U6550 ( .B1(n9245), .B2(n8986), .A(n8987), .ZN(n9227) );
  NAND2_X1 U6551 ( .A1(n8152), .A2(n8921), .ZN(n6816) );
  AOI21_X2 U6552 ( .B1(n9306), .B2(n6825), .A(n5387), .ZN(n9310) );
  AND2_X2 U6553 ( .A1(n6886), .A2(n6888), .ZN(n6851) );
  NAND2_X1 U6554 ( .A1(n6886), .A2(n5390), .ZN(n5391) );
  NAND2_X2 U6555 ( .A1(n8883), .A2(n8886), .ZN(n8851) );
  INV_X2 U6556 ( .A(n7466), .ZN(n9051) );
  NAND2_X1 U6557 ( .A1(n10200), .A2(n5395), .ZN(n10155) );
  NAND2_X1 U6558 ( .A1(n8527), .A2(n5400), .ZN(n10261) );
  INV_X1 U6559 ( .A(n5403), .ZN(n10281) );
  NAND2_X1 U6560 ( .A1(n5408), .A2(n5197), .ZN(n10271) );
  INV_X1 U6561 ( .A(n9921), .ZN(n5409) );
  NAND2_X1 U6562 ( .A1(n7883), .A2(n5413), .ZN(n5412) );
  NAND3_X1 U6563 ( .A1(n5412), .A2(n5411), .A3(n9881), .ZN(n8101) );
  NAND2_X1 U6564 ( .A1(n5140), .A2(n5416), .ZN(n7567) );
  OAI21_X2 U6565 ( .B1(n10227), .B2(n5421), .A(n5417), .ZN(n10183) );
  OAI21_X1 U6566 ( .B1(n5425), .B2(n5424), .A(n9896), .ZN(n5423) );
  OAI21_X1 U6567 ( .B1(n7658), .B2(n6336), .A(n9849), .ZN(n7711) );
  NAND2_X1 U6568 ( .A1(n6335), .A2(n9842), .ZN(n7658) );
  NOR2_X1 U6569 ( .A1(n7281), .A2(n5426), .ZN(n7241) );
  AND2_X1 U6570 ( .A1(n5427), .A2(n8018), .ZN(n5426) );
  INV_X1 U6571 ( .A(n7200), .ZN(n5434) );
  AOI21_X1 U6572 ( .B1(n5208), .B2(n5447), .A(n5446), .ZN(n10840) );
  NAND3_X1 U6573 ( .A1(n10790), .A2(n10794), .A3(n5472), .ZN(n5471) );
  AOI211_X1 U6574 ( .C1(n10789), .C2(keyinput_207), .A(n10787), .B(n10786), 
        .ZN(n10788) );
  NOR2_X1 U6575 ( .A1(n8551), .A2(n8550), .ZN(n9147) );
  NOR2_X1 U6576 ( .A1(n9147), .A2(n9146), .ZN(n9149) );
  AOI22_X1 U6577 ( .A1(n10676), .A2(keyinput_133), .B1(keyinput_135), .B2(
        n10675), .ZN(n10674) );
  INV_X1 U6578 ( .A(n6445), .ZN(n6456) );
  NAND3_X1 U6579 ( .A1(n5496), .A2(P2_REG2_REG_5__SCAN_IN), .A3(n7289), .ZN(
        n7290) );
  NAND2_X1 U6580 ( .A1(n7234), .A2(n7271), .ZN(n7289) );
  INV_X1 U6581 ( .A(n7234), .ZN(n5495) );
  INV_X1 U6582 ( .A(n8586), .ZN(n5502) );
  OAI21_X1 U6583 ( .B1(n7998), .B2(n5507), .A(n5506), .ZN(n8268) );
  INV_X1 U6584 ( .A(n9120), .ZN(n5511) );
  NAND4_X1 U6585 ( .A1(n6445), .A2(n6560), .A3(n6558), .A4(n6559), .ZN(n6561)
         );
  OAI21_X1 U6586 ( .B1(n7531), .B2(n5512), .A(n7532), .ZN(n7533) );
  NAND2_X1 U6587 ( .A1(n7531), .A2(n5512), .ZN(n7532) );
  XNOR2_X1 U6588 ( .A(n7487), .B(n7486), .ZN(n5512) );
  NAND2_X1 U6589 ( .A1(n8517), .A2(n5515), .ZN(n5514) );
  NAND2_X1 U6590 ( .A1(n8810), .A2(n5198), .ZN(n5521) );
  OAI211_X1 U6591 ( .C1(n8810), .C2(n5525), .A(n5522), .B(n5521), .ZN(n8700)
         );
  NAND2_X1 U6592 ( .A1(n8810), .A2(n5531), .ZN(n8811) );
  INV_X1 U6593 ( .A(n8809), .ZN(n5533) );
  INV_X1 U6594 ( .A(n6897), .ZN(n6847) );
  INV_X1 U6595 ( .A(n5534), .ZN(n7478) );
  OAI21_X1 U6596 ( .B1(n7476), .B2(n7515), .A(n7477), .ZN(n5534) );
  OR2_X1 U6597 ( .A1(n6897), .A2(n5535), .ZN(n7515) );
  NAND2_X1 U6598 ( .A1(n5537), .A2(n5536), .ZN(n8779) );
  NAND2_X1 U6599 ( .A1(n7895), .A2(n5202), .ZN(n8049) );
  NAND2_X2 U6600 ( .A1(n7780), .A2(n7779), .ZN(n7895) );
  NAND2_X1 U6601 ( .A1(n5551), .A2(n5550), .ZN(n6682) );
  NAND2_X1 U6602 ( .A1(n8657), .A2(n9256), .ZN(n5553) );
  NAND2_X1 U6603 ( .A1(n8769), .A2(n5553), .ZN(n8682) );
  AND2_X2 U6604 ( .A1(n6453), .A2(n6418), .ZN(n6445) );
  NAND3_X1 U6605 ( .A1(n10585), .A2(n10586), .A3(n5603), .ZN(n5602) );
  INV_X1 U6606 ( .A(n9530), .ZN(n5615) );
  NAND2_X1 U6607 ( .A1(n9530), .A2(n5610), .ZN(n5605) );
  NAND2_X2 U6608 ( .A1(n5605), .A2(n5607), .ZN(n9675) );
  NAND2_X1 U6609 ( .A1(n5962), .A2(n5616), .ZN(n5927) );
  NAND2_X1 U6610 ( .A1(n9601), .A2(n5619), .ZN(n5618) );
  NAND3_X1 U6611 ( .A1(n5637), .A2(n6950), .A3(n6949), .ZN(n5632) );
  NAND2_X1 U6612 ( .A1(n5633), .A2(n5636), .ZN(n5631) );
  NAND2_X1 U6613 ( .A1(n5636), .A2(n5635), .ZN(n5639) );
  INV_X1 U6614 ( .A(n5635), .ZN(n5626) );
  NAND2_X1 U6615 ( .A1(n5634), .A2(n5160), .ZN(n5627) );
  INV_X1 U6616 ( .A(n5634), .ZN(n5633) );
  NAND2_X1 U6617 ( .A1(n5635), .A2(n5637), .ZN(n5634) );
  INV_X1 U6618 ( .A(n5639), .ZN(n7753) );
  INV_X1 U6619 ( .A(n7754), .ZN(n5636) );
  NOR2_X2 U6620 ( .A1(n9561), .A2(n7059), .ZN(n7070) );
  NOR2_X1 U6621 ( .A1(n9541), .A2(n6978), .ZN(n5644) );
  NAND2_X1 U6622 ( .A1(n5643), .A2(n5640), .ZN(n9567) );
  INV_X1 U6623 ( .A(n5641), .ZN(n5640) );
  OAI21_X1 U6624 ( .B1(n9541), .B2(n5642), .A(n6992), .ZN(n5641) );
  NAND2_X1 U6625 ( .A1(n9657), .A2(n9538), .ZN(n5642) );
  NAND2_X1 U6626 ( .A1(n6979), .A2(n9657), .ZN(n5643) );
  INV_X1 U6627 ( .A(n6113), .ZN(n5649) );
  NAND2_X1 U6628 ( .A1(n5809), .A2(n5808), .ZN(n5895) );
  NAND2_X1 U6629 ( .A1(n5809), .A2(n5666), .ZN(n5665) );
  NAND3_X1 U6630 ( .A1(n5686), .A2(n5685), .A3(P1_DATAO_REG_1__SCAN_IN), .ZN(
        n5680) );
  NAND2_X2 U6631 ( .A1(n5889), .A2(n7134), .ZN(n9709) );
  NAND2_X1 U6632 ( .A1(n7713), .A2(n5693), .ZN(n5692) );
  NAND3_X1 U6633 ( .A1(n5692), .A2(n5691), .A3(n6050), .ZN(n7701) );
  NAND3_X1 U6634 ( .A1(n5995), .A2(n5978), .A3(n7690), .ZN(n5701) );
  NAND3_X1 U6635 ( .A1(n5701), .A2(n5702), .A3(n9775), .ZN(n7679) );
  NAND3_X1 U6636 ( .A1(n9836), .A2(n9834), .A3(n5995), .ZN(n5702) );
  NAND2_X1 U6637 ( .A1(n8199), .A2(n5137), .ZN(n5703) );
  NAND2_X1 U6638 ( .A1(n6270), .A2(n6269), .ZN(n10151) );
  NAND2_X1 U6639 ( .A1(n6270), .A2(n5201), .ZN(n6399) );
  AND3_X1 U6640 ( .A1(n5846), .A2(n5709), .A3(n5845), .ZN(n5860) );
  AND4_X2 U6641 ( .A1(n6469), .A2(n6466), .A3(n6468), .A4(n6467), .ZN(n7466)
         );
  INV_X1 U6642 ( .A(n5711), .ZN(n6771) );
  NAND2_X1 U6643 ( .A1(n6439), .A2(n5724), .ZN(n6429) );
  NAND2_X1 U6644 ( .A1(n6595), .A2(n5146), .ZN(n5733) );
  NAND2_X1 U6645 ( .A1(n6203), .A2(n6202), .ZN(n6235) );
  INV_X1 U6646 ( .A(n6203), .ZN(n6200) );
  XNOR2_X1 U6647 ( .A(n8599), .B(SI_29_), .ZN(n8540) );
  OR2_X1 U6648 ( .A1(n7601), .A2(n9758), .ZN(n11103) );
  OR2_X1 U6649 ( .A1(n9808), .A2(n9758), .ZN(n7117) );
  INV_X1 U6650 ( .A(n6935), .ZN(n6938) );
  XNOR2_X1 U6651 ( .A(n6320), .B(n10830), .ZN(n6324) );
  NAND2_X1 U6652 ( .A1(n8656), .A2(n8655), .ZN(n8657) );
  NAND2_X1 U6653 ( .A1(n7130), .A2(n8604), .ZN(n6493) );
  AND2_X1 U6654 ( .A1(n7479), .A2(n9051), .ZN(n7480) );
  AOI21_X1 U6655 ( .B1(n8678), .B2(n7593), .A(n7481), .ZN(n7540) );
  NAND2_X2 U6656 ( .A1(n8704), .A2(n6928), .ZN(n6943) );
  NAND2_X2 U6657 ( .A1(n6142), .A2(n5749), .ZN(n10280) );
  OAI21_X2 U6658 ( .B1(n8021), .B2(n6958), .A(n5755), .ZN(n6959) );
  OR2_X1 U6659 ( .A1(n6492), .A2(n6458), .ZN(n6460) );
  OR2_X1 U6660 ( .A1(n8220), .A2(n8390), .ZN(n5743) );
  INV_X1 U6661 ( .A(n8856), .ZN(n6817) );
  INV_X1 U6662 ( .A(n8718), .ZN(n8705) );
  AND4_X1 U6663 ( .A1(n6641), .A2(n6640), .A3(n6639), .A4(n6638), .ZN(n9375)
         );
  INV_X1 U6664 ( .A(n9266), .ZN(n9243) );
  AND2_X1 U6665 ( .A1(n6359), .A2(n5865), .ZN(n5744) );
  INV_X1 U6666 ( .A(n10366), .ZN(n6410) );
  OR2_X1 U6667 ( .A1(n8616), .A2(n9432), .ZN(n5745) );
  OR2_X1 U6668 ( .A1(n8616), .A2(n9508), .ZN(n5746) );
  OR2_X1 U6669 ( .A1(n7894), .A2(n8150), .ZN(n5747) );
  OR2_X1 U6670 ( .A1(n10390), .A2(n10297), .ZN(n5748) );
  OR2_X1 U6671 ( .A1(n10305), .A2(n6140), .ZN(n5749) );
  AND2_X1 U6672 ( .A1(n7490), .A2(n9049), .ZN(n5750) );
  INV_X2 U6673 ( .A(n11111), .ZN(n11114) );
  INV_X1 U6674 ( .A(n8659), .ZN(n9256) );
  INV_X1 U6675 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6432) );
  AND2_X1 U6676 ( .A1(n11114), .A2(n10399), .ZN(n6415) );
  INV_X1 U6677 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8116) );
  AND2_X1 U6678 ( .A1(n5790), .A2(n5789), .ZN(n5751) );
  OR2_X1 U6679 ( .A1(n10222), .A2(n10230), .ZN(n5752) );
  NAND2_X1 U6680 ( .A1(n7518), .A2(n9018), .ZN(n9376) );
  NAND2_X1 U6681 ( .A1(n7502), .A2(n9018), .ZN(n9361) );
  INV_X1 U6682 ( .A(n8150), .ZN(n6520) );
  INV_X1 U6683 ( .A(n5131), .ZN(n6086) );
  AND2_X1 U6684 ( .A1(n10147), .A2(n6415), .ZN(n5753) );
  INV_X1 U6685 ( .A(n10147), .ZN(n6910) );
  INV_X1 U6686 ( .A(n8207), .ZN(n9637) );
  AND2_X2 U6687 ( .A1(n9467), .A2(n7513), .ZN(n11121) );
  OR2_X1 U6688 ( .A1(n6957), .A2(n6956), .ZN(n5755) );
  INV_X1 U6689 ( .A(n7439), .ZN(n10003) );
  INV_X1 U6690 ( .A(n6332), .ZN(n5968) );
  INV_X1 U6691 ( .A(n8942), .ZN(n6605) );
  INV_X1 U6692 ( .A(keyinput_145), .ZN(n10692) );
  XNOR2_X1 U6693 ( .A(n10692), .B(SI_15_), .ZN(n10693) );
  NOR4_X1 U6694 ( .A1(n10750), .A2(n10749), .A3(n10748), .A4(n10747), .ZN(
        n10758) );
  OAI22_X1 U6695 ( .A1(n10763), .A2(keyinput_195), .B1(n10762), .B2(
        P2_DATAO_REG_29__SCAN_IN), .ZN(n10764) );
  INV_X1 U6696 ( .A(n10764), .ZN(n10765) );
  NAND2_X1 U6697 ( .A1(n10766), .A2(n10765), .ZN(n10767) );
  INV_X1 U6698 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n10773) );
  INV_X1 U6699 ( .A(keyinput_204), .ZN(n10781) );
  XNOR2_X1 U6700 ( .A(n10781), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n10782) );
  XNOR2_X1 U6701 ( .A(n10803), .B(keyinput_223), .ZN(n10804) );
  AOI21_X1 U6702 ( .B1(n10806), .B2(n10805), .A(n10804), .ZN(n10807) );
  INV_X1 U6703 ( .A(n10807), .ZN(n10810) );
  INV_X1 U6704 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6419) );
  INV_X1 U6705 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6111) );
  NAND2_X1 U6706 ( .A1(n7637), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7638) );
  INV_X1 U6707 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6425) );
  INV_X1 U6708 ( .A(n6134), .ZN(n5873) );
  INV_X1 U6709 ( .A(n10282), .ZN(n6140) );
  AND2_X1 U6710 ( .A1(n5864), .A2(n5863), .ZN(n5865) );
  INV_X1 U6711 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6694) );
  INV_X1 U6712 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6589) );
  AND2_X1 U6713 ( .A1(n7058), .A2(n7057), .ZN(n7059) );
  NAND2_X1 U6714 ( .A1(n5873), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6156) );
  NAND2_X1 U6715 ( .A1(n5874), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6171) );
  OR2_X1 U6716 ( .A1(n6057), .A2(n5919), .ZN(n6064) );
  AND2_X1 U6717 ( .A1(n6122), .A2(n5828), .ZN(n6143) );
  INV_X1 U6718 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6444) );
  INV_X1 U6719 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10724) );
  INV_X1 U6720 ( .A(n9046), .ZN(n8047) );
  INV_X1 U6721 ( .A(n8781), .ZN(n8648) );
  AND2_X1 U6722 ( .A1(n7781), .A2(n7782), .ZN(n7779) );
  OR2_X1 U6723 ( .A1(n6775), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6788) );
  NAND2_X1 U6724 ( .A1(n7637), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7624) );
  NOR2_X1 U6725 ( .A1(n6608), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6624) );
  NOR2_X1 U6726 ( .A1(n6523), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6544) );
  AND2_X1 U6727 ( .A1(n8975), .A2(n8974), .ZN(n9280) );
  OAI22_X1 U6728 ( .A1(n6497), .A2(n6812), .B1(n6496), .B2(n9049), .ZN(n7838)
         );
  INV_X1 U6729 ( .A(n7001), .ZN(n7002) );
  AND2_X1 U6730 ( .A1(n6087), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6102) );
  OR2_X1 U6731 ( .A1(n7077), .A2(n7076), .ZN(n7079) );
  OR2_X1 U6732 ( .A1(n7116), .A2(n7114), .ZN(n7120) );
  AND2_X1 U6733 ( .A1(n6294), .A2(n6282), .ZN(n10158) );
  AND2_X1 U6734 ( .A1(n10068), .A2(n8439), .ZN(n8440) );
  AND2_X1 U6735 ( .A1(n6311), .A2(n6295), .ZN(n8713) );
  OR2_X1 U6736 ( .A1(n7716), .A2(n9999), .ZN(n6037) );
  OR2_X1 U6737 ( .A1(n8239), .A2(n9998), .ZN(n6050) );
  NAND2_X1 U6738 ( .A1(n6009), .A2(n7940), .ZN(n6010) );
  NAND2_X1 U6739 ( .A1(n5968), .A2(n11034), .ZN(n5969) );
  AND2_X1 U6740 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n5853) );
  NAND2_X1 U6741 ( .A1(n5805), .A2(n10695), .ZN(n5808) );
  NAND2_X1 U6742 ( .A1(n10724), .A2(n6624), .ZN(n6637) );
  NAND2_X1 U6743 ( .A1(n8046), .A2(n8047), .ZN(n8048) );
  NAND2_X1 U6744 ( .A1(n10732), .A2(n6599), .ZN(n6608) );
  INV_X1 U6745 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n10658) );
  AND2_X1 U6746 ( .A1(n8683), .A2(n8681), .ZN(n8770) );
  INV_X1 U6747 ( .A(n9292), .ZN(n8742) );
  NOR2_X1 U6748 ( .A1(n6904), .A2(n6873), .ZN(n7514) );
  AND2_X1 U6749 ( .A1(n8825), .A2(n8821), .ZN(n8637) );
  AND2_X1 U6750 ( .A1(n6883), .A2(n6882), .ZN(n6884) );
  NAND2_X1 U6751 ( .A1(n6564), .A2(n10556), .ZN(n6566) );
  AND2_X1 U6752 ( .A1(n6544), .A2(n6543), .ZN(n6564) );
  NOR2_X1 U6753 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6498) );
  AND2_X1 U6754 ( .A1(n7500), .A2(n9450), .ZN(n7595) );
  INV_X1 U6755 ( .A(n11121), .ZN(n6890) );
  INV_X1 U6756 ( .A(n9039), .ZN(n9374) );
  INV_X1 U6757 ( .A(n9040), .ZN(n8507) );
  INV_X1 U6758 ( .A(n9342), .ZN(n9373) );
  INV_X1 U6759 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6427) );
  INV_X1 U6760 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6446) );
  INV_X2 U6761 ( .A(n7134), .ZN(n8604) );
  NAND2_X1 U6762 ( .A1(n7000), .A2(n7002), .ZN(n7003) );
  NAND2_X1 U6763 ( .A1(n9675), .A2(n7103), .ZN(n8702) );
  INV_X1 U6764 ( .A(n6936), .ZN(n6937) );
  AND3_X1 U6765 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n6017) );
  AND2_X1 U6766 ( .A1(n7079), .A2(n7078), .ZN(n9610) );
  OR2_X1 U6767 ( .A1(n7120), .A2(n7258), .ZN(n9644) );
  OR2_X1 U6768 ( .A1(n11079), .A2(n9987), .ZN(n10219) );
  NAND2_X1 U6769 ( .A1(n6327), .A2(n6328), .ZN(n9808) );
  INV_X1 U6770 ( .A(n10300), .ZN(n10400) );
  OR2_X1 U6771 ( .A1(n7601), .A2(n9986), .ZN(n10300) );
  AND2_X1 U6772 ( .A1(n6123), .A2(n5821), .ZN(n6122) );
  INV_X1 U6773 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6098) );
  INV_X1 U6774 ( .A(n8829), .ZN(n8815) );
  AND4_X1 U6775 ( .A1(n6793), .A2(n6792), .A3(n6791), .A4(n6790), .ZN(n9189)
         );
  AND4_X1 U6776 ( .A1(n6759), .A2(n6758), .A3(n6757), .A4(n6756), .ZN(n9225)
         );
  AND4_X1 U6777 ( .A1(n6664), .A2(n6663), .A3(n6662), .A4(n6661), .ZN(n8966)
         );
  AND4_X1 U6778 ( .A1(n6587), .A2(n6586), .A3(n6585), .A4(n6584), .ZN(n8402)
         );
  NAND2_X1 U6779 ( .A1(n6885), .A2(n6884), .ZN(n7505) );
  INV_X1 U6780 ( .A(n10968), .ZN(n11014) );
  INV_X1 U6781 ( .A(n10983), .ZN(n10997) );
  AOI21_X1 U6782 ( .B1(n5504), .B2(n8589), .A(n11014), .ZN(n8590) );
  INV_X1 U6783 ( .A(n8160), .ZN(n8130) );
  OR2_X1 U6784 ( .A1(n7516), .A2(n7515), .ZN(n9380) );
  OR2_X1 U6785 ( .A1(n9456), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6907) );
  AND2_X1 U6786 ( .A1(n6904), .A2(n6903), .ZN(n7589) );
  INV_X1 U6787 ( .A(n9414), .ZN(n9458) );
  OR2_X1 U6788 ( .A1(n8385), .A2(n8016), .ZN(n9414) );
  XNOR2_X1 U6789 ( .A(n6809), .B(P2_IR_REG_22__SCAN_IN), .ZN(n9028) );
  NAND2_X1 U6790 ( .A1(n7119), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9646) );
  INV_X1 U6791 ( .A(n5970), .ZN(n6358) );
  AND4_X1 U6792 ( .A1(n6192), .A2(n6191), .A3(n6190), .A4(n6189), .ZN(n10248)
         );
  AND4_X1 U6793 ( .A1(n5886), .A2(n5885), .A3(n5884), .A4(n5883), .ZN(n10389)
         );
  AND4_X1 U6794 ( .A1(n5924), .A2(n5923), .A3(n5922), .A4(n5921), .ZN(n9654)
         );
  OR2_X1 U6795 ( .A1(n7259), .A2(n9699), .ZN(n8444) );
  INV_X1 U6796 ( .A(n10119), .ZN(n10869) );
  INV_X1 U6797 ( .A(n10121), .ZN(n10866) );
  INV_X1 U6798 ( .A(n8444), .ZN(n10871) );
  AND2_X1 U6799 ( .A1(n9909), .A2(n9910), .ZN(n9789) );
  INV_X1 U6800 ( .A(n10219), .ZN(n11065) );
  INV_X1 U6801 ( .A(n10388), .ZN(n11089) );
  OR2_X1 U6802 ( .A1(n9808), .A2(n7258), .ZN(n10375) );
  INV_X1 U6803 ( .A(n11103), .ZN(n10399) );
  INV_X1 U6804 ( .A(n11107), .ZN(n11023) );
  NAND2_X1 U6805 ( .A1(n11084), .A2(n11085), .ZN(n11107) );
  NAND2_X1 U6806 ( .A1(n6373), .A2(n6372), .ZN(n10466) );
  XNOR2_X1 U6807 ( .A(n6303), .B(n6302), .ZN(n8482) );
  OR3_X1 U6808 ( .A1(n7498), .A2(n7497), .A3(n7499), .ZN(n8788) );
  INV_X1 U6809 ( .A(n8786), .ZN(n8835) );
  INV_X1 U6810 ( .A(n8402), .ZN(n9041) );
  OR2_X1 U6811 ( .A1(P2_U3150), .A2(n7175), .ZN(n9095) );
  OR2_X1 U6812 ( .A1(n7202), .A2(n7193), .ZN(n11005) );
  NAND2_X1 U6813 ( .A1(n7594), .A2(n9216), .ZN(n9317) );
  INV_X1 U6814 ( .A(n9377), .ZN(n9315) );
  INV_X1 U6815 ( .A(n9377), .ZN(n9353) );
  INV_X1 U6816 ( .A(n9320), .ZN(n9388) );
  NAND2_X1 U6817 ( .A1(n9456), .A2(n9463), .ZN(n9432) );
  INV_X1 U6818 ( .A(n9456), .ZN(n9465) );
  AND2_X2 U6819 ( .A1(n6905), .A2(n7589), .ZN(n9456) );
  AND2_X1 U6820 ( .A1(n8118), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7150) );
  INV_X1 U6821 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8120) );
  INV_X1 U6822 ( .A(n9694), .ZN(n9636) );
  AND4_X1 U6823 ( .A1(n6316), .A2(n6315), .A3(n6314), .A4(n6313), .ZN(n8714)
         );
  AND4_X1 U6824 ( .A1(n6121), .A2(n6120), .A3(n6119), .A4(n6118), .ZN(n10297)
         );
  OR2_X1 U6825 ( .A1(n7250), .A2(n7249), .ZN(n7259) );
  OR2_X1 U6826 ( .A1(n7259), .A2(n7258), .ZN(n10121) );
  OR2_X1 U6827 ( .A1(n7259), .A2(n7378), .ZN(n10125) );
  OR2_X1 U6828 ( .A1(n11079), .A2(n7554), .ZN(n11072) );
  OR2_X1 U6829 ( .A1(n11069), .A2(n7744), .ZN(n10309) );
  INV_X1 U6830 ( .A(n10307), .ZN(n11069) );
  AOI21_X1 U6831 ( .B1(n10147), .B2(n6410), .A(n6912), .ZN(n6913) );
  NAND2_X1 U6832 ( .A1(n11110), .A2(n10399), .ZN(n10366) );
  INV_X1 U6833 ( .A(n11110), .ZN(n11109) );
  INV_X1 U6834 ( .A(n10157), .ZN(n10434) );
  INV_X1 U6835 ( .A(n6415), .ZN(n10457) );
  NAND2_X1 U6836 ( .A1(n6408), .A2(n7551), .ZN(n11111) );
  INV_X1 U6837 ( .A(n10480), .ZN(n10481) );
  AND2_X1 U6838 ( .A1(n6391), .A2(n8114), .ZN(n10468) );
  INV_X1 U6839 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n10485) );
  INV_X1 U6840 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n10581) );
  INV_X1 U6841 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10785) );
  INV_X1 U6842 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10792) );
  INV_X1 U6843 ( .A(n9045), .ZN(P2_U3893) );
  AND2_X2 U6844 ( .A1(n7127), .A2(n8114), .ZN(P1_U3973) );
  OAI21_X1 U6845 ( .B1(n6914), .B2(n11111), .A(n6397), .ZN(P1_U3519) );
  AND2_X1 U6846 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5756) );
  NAND2_X1 U6847 ( .A1(n5768), .A2(n5756), .ZN(n5952) );
  AND2_X1 U6848 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5757) );
  NAND2_X1 U6849 ( .A1(n7134), .A2(n5757), .ZN(n6484) );
  NAND2_X1 U6850 ( .A1(n5952), .A2(n6484), .ZN(n5958) );
  INV_X1 U6851 ( .A(SI_1_), .ZN(n5758) );
  XNOR2_X1 U6852 ( .A(n5759), .B(n5758), .ZN(n5959) );
  NAND2_X1 U6853 ( .A1(n5958), .A2(n5959), .ZN(n5761) );
  NAND2_X1 U6854 ( .A1(n5759), .A2(SI_1_), .ZN(n5760) );
  NAND2_X1 U6855 ( .A1(n5761), .A2(n5760), .ZN(n5977) );
  MUX2_X1 U6856 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5768), .Z(n5762) );
  INV_X1 U6857 ( .A(SI_2_), .ZN(n10706) );
  XNOR2_X1 U6858 ( .A(n5762), .B(n10706), .ZN(n5976) );
  NAND2_X1 U6859 ( .A1(n5977), .A2(n5976), .ZN(n5764) );
  NAND2_X1 U6860 ( .A1(n5762), .A2(SI_2_), .ZN(n5763) );
  INV_X1 U6861 ( .A(SI_3_), .ZN(n5765) );
  XNOR2_X1 U6862 ( .A(n5766), .B(n5765), .ZN(n5990) );
  NAND2_X1 U6863 ( .A1(n5766), .A2(SI_3_), .ZN(n5767) );
  INV_X1 U6864 ( .A(SI_4_), .ZN(n10526) );
  XNOR2_X1 U6865 ( .A(n5769), .B(n10526), .ZN(n6005) );
  NAND2_X1 U6866 ( .A1(n5769), .A2(SI_4_), .ZN(n5770) );
  INV_X1 U6867 ( .A(SI_5_), .ZN(n5771) );
  XNOR2_X1 U6868 ( .A(n5772), .B(n5771), .ZN(n5941) );
  NAND2_X1 U6869 ( .A1(n5942), .A2(n5941), .ZN(n5774) );
  NAND2_X1 U6870 ( .A1(n5772), .A2(SI_5_), .ZN(n5773) );
  INV_X1 U6871 ( .A(SI_6_), .ZN(n10707) );
  XNOR2_X1 U6872 ( .A(n5775), .B(n10707), .ZN(n6011) );
  NAND2_X1 U6873 ( .A1(n6012), .A2(n6011), .ZN(n5777) );
  NAND2_X1 U6874 ( .A1(n5775), .A2(SI_6_), .ZN(n5776) );
  XNOR2_X1 U6875 ( .A(n5779), .B(SI_7_), .ZN(n6024) );
  INV_X1 U6876 ( .A(n6024), .ZN(n5778) );
  NAND2_X1 U6877 ( .A1(n5779), .A2(SI_7_), .ZN(n5780) );
  NAND2_X1 U6878 ( .A1(n5781), .A2(n10518), .ZN(n5784) );
  INV_X1 U6879 ( .A(n5781), .ZN(n5782) );
  NAND2_X1 U6880 ( .A1(n5782), .A2(SI_8_), .ZN(n5783) );
  NAND2_X1 U6881 ( .A1(n5784), .A2(n5783), .ZN(n6038) );
  INV_X1 U6882 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5785) );
  INV_X1 U6883 ( .A(SI_9_), .ZN(n5786) );
  NAND2_X1 U6884 ( .A1(n5787), .A2(n5786), .ZN(n5790) );
  INV_X1 U6885 ( .A(n5787), .ZN(n5788) );
  NAND2_X1 U6886 ( .A1(n5788), .A2(SI_9_), .ZN(n5789) );
  NAND2_X1 U6887 ( .A1(n5791), .A2(n5790), .ZN(n5926) );
  XNOR2_X1 U6888 ( .A(n5793), .B(SI_10_), .ZN(n5925) );
  INV_X1 U6889 ( .A(n5925), .ZN(n5792) );
  INV_X1 U6890 ( .A(n5793), .ZN(n5794) );
  NAND2_X1 U6891 ( .A1(n5794), .A2(SI_10_), .ZN(n5795) );
  NAND2_X1 U6892 ( .A1(n5796), .A2(n10491), .ZN(n5799) );
  INV_X1 U6893 ( .A(n5796), .ZN(n5797) );
  NAND2_X1 U6894 ( .A1(n5797), .A2(SI_11_), .ZN(n5798) );
  NAND2_X1 U6895 ( .A1(n5799), .A2(n5798), .ZN(n6071) );
  MUX2_X1 U6896 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n8604), .Z(n5800) );
  NAND2_X1 U6897 ( .A1(n5800), .A2(SI_12_), .ZN(n5801) );
  MUX2_X1 U6898 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n8604), .Z(n5804) );
  XNOR2_X1 U6899 ( .A(n5804), .B(SI_13_), .ZN(n6095) );
  INV_X1 U6900 ( .A(n6095), .ZN(n5803) );
  MUX2_X1 U6901 ( .A(n7397), .B(n10593), .S(n8604), .Z(n5805) );
  INV_X1 U6902 ( .A(n5805), .ZN(n5806) );
  NAND2_X1 U6903 ( .A1(n5806), .A2(SI_14_), .ZN(n5807) );
  NAND2_X1 U6904 ( .A1(n5808), .A2(n5807), .ZN(n5914) );
  MUX2_X1 U6905 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n8604), .Z(n5811) );
  INV_X1 U6906 ( .A(SI_15_), .ZN(n5810) );
  XNOR2_X1 U6907 ( .A(n5811), .B(n5810), .ZN(n5894) );
  INV_X1 U6908 ( .A(n5894), .ZN(n5813) );
  NAND2_X1 U6909 ( .A1(n5811), .A2(SI_15_), .ZN(n5812) );
  MUX2_X1 U6910 ( .A(n7609), .B(n10785), .S(n8604), .Z(n5815) );
  INV_X1 U6911 ( .A(SI_16_), .ZN(n5814) );
  INV_X1 U6912 ( .A(n5815), .ZN(n5816) );
  NAND2_X1 U6913 ( .A1(n5816), .A2(SI_16_), .ZN(n5817) );
  INV_X1 U6914 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7740) );
  MUX2_X1 U6915 ( .A(n7740), .B(n10789), .S(n8604), .Z(n5819) );
  NAND2_X1 U6916 ( .A1(n5819), .A2(n10690), .ZN(n6123) );
  INV_X1 U6917 ( .A(n5819), .ZN(n5820) );
  NAND2_X1 U6918 ( .A1(n5820), .A2(SI_17_), .ZN(n5821) );
  MUX2_X1 U6919 ( .A(n7826), .B(n7794), .S(n8604), .Z(n5829) );
  INV_X1 U6920 ( .A(n5829), .ZN(n5822) );
  NAND2_X1 U6921 ( .A1(n5822), .A2(SI_18_), .ZN(n5828) );
  MUX2_X1 U6922 ( .A(n7847), .B(n8723), .S(n8604), .Z(n5823) );
  NAND2_X1 U6923 ( .A1(n5823), .A2(n10667), .ZN(n5832) );
  INV_X1 U6924 ( .A(n5823), .ZN(n5824) );
  NAND2_X1 U6925 ( .A1(n5824), .A2(SI_19_), .ZN(n5825) );
  NAND2_X1 U6926 ( .A1(n5832), .A2(n5825), .ZN(n6147) );
  INV_X1 U6927 ( .A(n6147), .ZN(n5826) );
  NAND2_X1 U6928 ( .A1(n6144), .A2(n5827), .ZN(n5835) );
  INV_X1 U6929 ( .A(n5828), .ZN(n5831) );
  XNOR2_X1 U6930 ( .A(n5829), .B(SI_18_), .ZN(n6125) );
  NAND2_X1 U6931 ( .A1(n5835), .A2(n5834), .ZN(n6164) );
  MUX2_X1 U6932 ( .A(n6694), .B(n7850), .S(n8604), .Z(n5836) );
  NAND2_X1 U6933 ( .A1(n5836), .A2(n10685), .ZN(n5839) );
  INV_X1 U6934 ( .A(n5836), .ZN(n5837) );
  NAND2_X1 U6935 ( .A1(n5837), .A2(SI_20_), .ZN(n5838) );
  NAND2_X1 U6936 ( .A1(n6164), .A2(n6163), .ZN(n5840) );
  MUX2_X1 U6937 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n8604), .Z(n6179) );
  XNOR2_X1 U6938 ( .A(n6179), .B(n10684), .ZN(n6178) );
  XNOR2_X1 U6939 ( .A(n6177), .B(n6178), .ZN(n7890) );
  NOR2_X1 U6940 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5844) );
  NOR2_X1 U6941 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5849) );
  NOR2_X1 U6942 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5848) );
  NAND4_X1 U6943 ( .A1(n6318), .A2(n5849), .A3(n5848), .A4(n5847), .ZN(n5851)
         );
  NAND4_X1 U6944 ( .A1(n10830), .A2(n6387), .A3(n6321), .A4(n10835), .ZN(n5850) );
  NOR2_X2 U6945 ( .A1(n5851), .A2(n5850), .ZN(n6359) );
  NOR2_X1 U6946 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n5862) );
  INV_X1 U6947 ( .A(n5862), .ZN(n5854) );
  INV_X1 U6948 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5855) );
  NAND3_X1 U6949 ( .A1(n6370), .A2(P1_IR_REG_31__SCAN_IN), .A3(n5855), .ZN(
        n5856) );
  NAND2_X1 U6950 ( .A1(n7890), .A2(n9708), .ZN(n5859) );
  INV_X1 U6951 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n10777) );
  OR2_X1 U6952 ( .A1(n9709), .A2(n10777), .ZN(n5858) );
  AND2_X1 U6953 ( .A1(n5862), .A2(n5861), .ZN(n5864) );
  NAND2_X1 U6954 ( .A1(n5131), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5881) );
  INV_X2 U6955 ( .A(n6358), .ZN(n9704) );
  NAND2_X1 U6956 ( .A1(n9704), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5880) );
  INV_X1 U6957 ( .A(n8634), .ZN(n5872) );
  CLKBUF_X3 U6958 ( .A(n5980), .Z(n6312) );
  NAND2_X1 U6959 ( .A1(n6017), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U6960 ( .A1(n6044), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6055) );
  INV_X1 U6961 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5901) );
  INV_X1 U6962 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5882) );
  NAND2_X1 U6963 ( .A1(n6117), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6134) );
  INV_X1 U6964 ( .A(n6169), .ZN(n5874) );
  INV_X1 U6965 ( .A(n6171), .ZN(n5875) );
  INV_X1 U6966 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5876) );
  NAND2_X1 U6967 ( .A1(n6171), .A2(n5876), .ZN(n5877) );
  AND2_X1 U6968 ( .A1(n6187), .A2(n5877), .ZN(n10254) );
  NAND2_X1 U6969 ( .A1(n6312), .A2(n10254), .ZN(n5879) );
  NAND2_X1 U6970 ( .A1(n6066), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5878) );
  INV_X1 U6971 ( .A(n10273), .ZN(n10231) );
  NAND2_X1 U6972 ( .A1(n9704), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5886) );
  NAND2_X1 U6973 ( .A1(n5132), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5885) );
  AOI21_X1 U6974 ( .B1(n5903), .B2(n5882), .A(n6117), .ZN(n9591) );
  NAND2_X1 U6975 ( .A1(n6312), .A2(n9591), .ZN(n5884) );
  NAND2_X1 U6976 ( .A1(n6066), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5883) );
  XNOR2_X1 U6977 ( .A(n5888), .B(n5887), .ZN(n7607) );
  NAND2_X1 U6978 ( .A1(n7607), .A2(n9708), .ZN(n5893) );
  NAND2_X1 U6979 ( .A1(n6360), .A2(n5890), .ZN(n6113) );
  NAND2_X1 U6980 ( .A1(n6113), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5896) );
  NAND2_X1 U6981 ( .A1(n5896), .A2(n6110), .ZN(n5898) );
  NAND2_X1 U6982 ( .A1(n5898), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5891) );
  XNOR2_X1 U6983 ( .A(n5891), .B(P1_IR_REG_16__SCAN_IN), .ZN(n10080) );
  AOI22_X1 U6984 ( .A1(n6153), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6152), .B2(
        n10080), .ZN(n5892) );
  INV_X1 U6985 ( .A(n10398), .ZN(n8492) );
  XNOR2_X1 U6986 ( .A(n5895), .B(n5894), .ZN(n7408) );
  NAND2_X1 U6987 ( .A1(n7408), .A2(n9708), .ZN(n5900) );
  OR2_X1 U6988 ( .A1(n5896), .A2(n6110), .ZN(n5897) );
  AND2_X1 U6989 ( .A1(n5898), .A2(n5897), .ZN(n10865) );
  AOI22_X1 U6990 ( .A1(n6153), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6152), .B2(
        n10865), .ZN(n5899) );
  NAND2_X1 U6991 ( .A1(n5131), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5907) );
  NAND2_X1 U6992 ( .A1(n9704), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5906) );
  NAND2_X1 U6993 ( .A1(n5908), .A2(n5901), .ZN(n5902) );
  AND2_X1 U6994 ( .A1(n5903), .A2(n5902), .ZN(n9688) );
  NAND2_X1 U6995 ( .A1(n6312), .A2(n9688), .ZN(n5905) );
  NAND2_X1 U6996 ( .A1(n6066), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5904) );
  NAND2_X1 U6997 ( .A1(n9704), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5913) );
  NAND2_X1 U6998 ( .A1(n5132), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5912) );
  OR2_X1 U6999 ( .A1(n6104), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5909) );
  AND2_X1 U7000 ( .A1(n5909), .A2(n5908), .ZN(n9524) );
  NAND2_X1 U7001 ( .A1(n6312), .A2(n9524), .ZN(n5911) );
  NAND2_X1 U7002 ( .A1(n6066), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5910) );
  XNOR2_X1 U7003 ( .A(n5915), .B(n5914), .ZN(n7395) );
  NAND2_X1 U7004 ( .A1(n7395), .A2(n9708), .ZN(n5918) );
  OR2_X1 U7005 ( .A1(n6360), .A2(n6098), .ZN(n5916) );
  XNOR2_X1 U7006 ( .A(n5916), .B(P1_IR_REG_14__SCAN_IN), .ZN(n10063) );
  AOI22_X1 U7007 ( .A1(n6153), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6152), .B2(
        n10063), .ZN(n5917) );
  INV_X1 U7008 ( .A(n9527), .ZN(n10418) );
  NAND2_X1 U7009 ( .A1(n9704), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5924) );
  NAND2_X1 U7010 ( .A1(n6167), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5923) );
  NAND2_X1 U7011 ( .A1(n6057), .A2(n5919), .ZN(n5920) );
  AND2_X1 U7012 ( .A1(n6064), .A2(n5920), .ZN(n9542) );
  NAND2_X1 U7013 ( .A1(n6312), .A2(n9542), .ZN(n5922) );
  NAND2_X1 U7014 ( .A1(n6066), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5921) );
  INV_X1 U7015 ( .A(n9654), .ZN(n11090) );
  XNOR2_X1 U7016 ( .A(n5926), .B(n5925), .ZN(n7166) );
  NAND2_X1 U7017 ( .A1(n7166), .A2(n9708), .ZN(n5935) );
  NOR2_X1 U7018 ( .A1(n5927), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n6001) );
  NAND2_X1 U7019 ( .A1(n6001), .A2(n10803), .ZN(n6026) );
  NAND2_X1 U7020 ( .A1(n5928), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6051) );
  INV_X1 U7021 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5929) );
  NAND2_X1 U7022 ( .A1(n6051), .A2(n5929), .ZN(n5930) );
  NAND2_X1 U7023 ( .A1(n5930), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5932) );
  INV_X1 U7024 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5931) );
  OR2_X1 U7025 ( .A1(n5932), .A2(n5931), .ZN(n5933) );
  NAND2_X1 U7026 ( .A1(n5932), .A2(n5931), .ZN(n6073) );
  AOI22_X1 U7027 ( .A1(n6153), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6152), .B2(
        n7617), .ZN(n5934) );
  NAND2_X1 U7028 ( .A1(n5970), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5940) );
  NAND2_X1 U7029 ( .A1(n6167), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5939) );
  AOI21_X1 U7030 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5936) );
  NOR2_X1 U7031 ( .A1(n5936), .A2(n6017), .ZN(n7989) );
  NAND2_X1 U7032 ( .A1(n6312), .A2(n7989), .ZN(n5938) );
  NAND2_X1 U7033 ( .A1(n6066), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5937) );
  XNOR2_X1 U7034 ( .A(n5942), .B(n5941), .ZN(n7138) );
  OR2_X1 U7035 ( .A1(n7138), .A2(n6013), .ZN(n5945) );
  OR2_X1 U7036 ( .A1(n6001), .A2(n6098), .ZN(n5943) );
  XNOR2_X1 U7037 ( .A(n5943), .B(P1_IR_REG_5__SCAN_IN), .ZN(n7342) );
  AOI22_X1 U7038 ( .A1(n6153), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6152), .B2(
        n7342), .ZN(n5944) );
  NAND2_X1 U7039 ( .A1(n5945), .A2(n5944), .ZN(n7946) );
  NAND2_X1 U7040 ( .A1(n5970), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5949) );
  NAND2_X1 U7041 ( .A1(n5131), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5948) );
  NAND2_X1 U7042 ( .A1(n5980), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5947) );
  NAND2_X1 U7043 ( .A1(n6066), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5946) );
  NAND4_X1 U7044 ( .A1(n5949), .A2(n5948), .A3(n5947), .A4(n5946), .ZN(n10005)
         );
  NAND2_X1 U7045 ( .A1(n8604), .A2(SI_0_), .ZN(n5951) );
  INV_X1 U7046 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5950) );
  NAND2_X1 U7047 ( .A1(n5951), .A2(n5950), .ZN(n5953) );
  AND2_X1 U7048 ( .A1(n5953), .A2(n5952), .ZN(n10479) );
  MUX2_X1 U7049 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10479), .S(n5889), .Z(n11024)
         );
  NAND2_X1 U7050 ( .A1(n10005), .A2(n11024), .ZN(n7571) );
  NAND2_X1 U7051 ( .A1(n5971), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5957) );
  NAND2_X1 U7052 ( .A1(n5970), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5956) );
  NAND2_X1 U7053 ( .A1(n5980), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5955) );
  NAND2_X1 U7054 ( .A1(n6066), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5954) );
  XNOR2_X1 U7055 ( .A(n5959), .B(n5958), .ZN(n7136) );
  OR2_X1 U7056 ( .A1(n6013), .A2(n7136), .ZN(n5967) );
  OR2_X1 U7057 ( .A1(n9709), .A2(n5684), .ZN(n5966) );
  NAND2_X1 U7058 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5961) );
  INV_X1 U7059 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5960) );
  MUX2_X1 U7060 ( .A(n5961), .B(P1_IR_REG_31__SCAN_IN), .S(n5960), .Z(n5964)
         );
  INV_X1 U7061 ( .A(n5962), .ZN(n5963) );
  NAND2_X1 U7062 ( .A1(n5964), .A2(n5963), .ZN(n7310) );
  OR2_X1 U7063 ( .A1(n5889), .A2(n7310), .ZN(n5965) );
  INV_X1 U7064 ( .A(n11034), .ZN(n6934) );
  NAND2_X1 U7065 ( .A1(n7570), .A2(n5969), .ZN(n7691) );
  NAND2_X1 U7066 ( .A1(n5970), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5975) );
  NAND2_X1 U7067 ( .A1(n5132), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5974) );
  NAND2_X1 U7068 ( .A1(n5980), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5973) );
  NAND2_X1 U7069 ( .A1(n6066), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5972) );
  OR2_X1 U7070 ( .A1(n5962), .A2(n6098), .ZN(n5986) );
  INV_X1 U7071 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5985) );
  XNOR2_X1 U7072 ( .A(n5986), .B(n5985), .ZN(n7388) );
  XNOR2_X1 U7073 ( .A(n5977), .B(n5976), .ZN(n6458) );
  INV_X1 U7074 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n7135) );
  NAND2_X1 U7075 ( .A1(n7568), .A2(n7694), .ZN(n9833) );
  INV_X1 U7076 ( .A(n7568), .ZN(n10004) );
  NAND2_X1 U7077 ( .A1(n10004), .A2(n8074), .ZN(n9831) );
  NAND2_X1 U7078 ( .A1(n9833), .A2(n9831), .ZN(n7689) );
  NAND2_X1 U7079 ( .A1(n7691), .A2(n7689), .ZN(n7690) );
  OR2_X1 U7080 ( .A1(n10004), .A2(n7694), .ZN(n5978) );
  NAND2_X1 U7081 ( .A1(n5131), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5984) );
  NAND2_X1 U7082 ( .A1(n6066), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5983) );
  INV_X1 U7083 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5979) );
  NAND2_X1 U7084 ( .A1(n5980), .A2(n5979), .ZN(n5982) );
  NAND2_X1 U7085 ( .A1(n5970), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5981) );
  NAND2_X1 U7086 ( .A1(n5986), .A2(n5985), .ZN(n5987) );
  NAND2_X1 U7087 ( .A1(n5987), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5989) );
  INV_X1 U7088 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5988) );
  XNOR2_X1 U7089 ( .A(n5989), .B(n5988), .ZN(n10006) );
  XNOR2_X1 U7090 ( .A(n5991), .B(n5990), .ZN(n8624) );
  OR2_X1 U7091 ( .A1(n6013), .A2(n8624), .ZN(n5993) );
  INV_X1 U7092 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n8622) );
  OR2_X1 U7093 ( .A1(n9709), .A2(n8622), .ZN(n5992) );
  OAI211_X1 U7094 ( .C1(n5889), .C2(n10006), .A(n5993), .B(n5992), .ZN(n5994)
         );
  NAND2_X1 U7095 ( .A1(n7439), .A2(n5994), .ZN(n9834) );
  INV_X1 U7096 ( .A(n5994), .ZN(n11044) );
  NAND2_X1 U7097 ( .A1(n10003), .A2(n11044), .ZN(n9836) );
  NAND2_X1 U7098 ( .A1(n5970), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6000) );
  NAND2_X1 U7099 ( .A1(n6167), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5999) );
  INV_X1 U7100 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5996) );
  XNOR2_X1 U7101 ( .A(n5996), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n7755) );
  NAND2_X1 U7102 ( .A1(n6312), .A2(n7755), .ZN(n5998) );
  NAND2_X1 U7103 ( .A1(n6066), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5997) );
  INV_X1 U7104 ( .A(n6001), .ZN(n6004) );
  NAND2_X1 U7105 ( .A1(n5927), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6002) );
  MUX2_X1 U7106 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6002), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n6003) );
  NAND2_X1 U7107 ( .A1(n6004), .A2(n6003), .ZN(n10022) );
  XNOR2_X1 U7108 ( .A(n6006), .B(n6005), .ZN(n6505) );
  OR2_X1 U7109 ( .A1(n6505), .A2(n6013), .ZN(n6008) );
  INV_X1 U7110 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n7141) );
  OR2_X1 U7111 ( .A1(n9709), .A2(n7141), .ZN(n6007) );
  OAI211_X1 U7112 ( .C1(n5889), .C2(n10022), .A(n6008), .B(n6007), .ZN(n7923)
         );
  NAND2_X1 U7113 ( .A1(n7940), .A2(n7923), .ZN(n9827) );
  NAND2_X1 U7114 ( .A1(n10002), .A2(n6009), .ZN(n9837) );
  NAND2_X1 U7115 ( .A1(n9827), .A2(n9837), .ZN(n9775) );
  NAND2_X1 U7116 ( .A1(n7679), .A2(n6010), .ZN(n7942) );
  INV_X1 U7117 ( .A(n7946), .ZN(n11056) );
  NAND2_X1 U7118 ( .A1(n10001), .A2(n11056), .ZN(n9842) );
  NAND2_X1 U7119 ( .A1(n7942), .A2(n9847), .ZN(n7941) );
  OAI21_X1 U7120 ( .B1(n10001), .B2(n7946), .A(n7941), .ZN(n7657) );
  XNOR2_X1 U7121 ( .A(n6012), .B(n6011), .ZN(n7142) );
  OR2_X1 U7122 ( .A1(n7142), .A2(n6013), .ZN(n6016) );
  NAND2_X1 U7123 ( .A1(n6026), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6014) );
  XNOR2_X1 U7124 ( .A(n6014), .B(P1_IR_REG_6__SCAN_IN), .ZN(n7356) );
  AOI22_X1 U7125 ( .A1(n6153), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6152), .B2(
        n7356), .ZN(n6015) );
  NAND2_X1 U7126 ( .A1(n9704), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6022) );
  NAND2_X1 U7127 ( .A1(n6167), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6021) );
  OAI21_X1 U7128 ( .B1(n6017), .B2(P1_REG3_REG_6__SCAN_IN), .A(n6031), .ZN(
        n6018) );
  INV_X1 U7129 ( .A(n6018), .ZN(n11068) );
  NAND2_X1 U7130 ( .A1(n6312), .A2(n11068), .ZN(n6020) );
  NAND2_X1 U7131 ( .A1(n6066), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6019) );
  NAND4_X1 U7132 ( .A1(n6022), .A2(n6021), .A3(n6020), .A4(n6019), .ZN(n10000)
         );
  NAND2_X1 U7133 ( .A1(n11073), .A2(n10000), .ZN(n9850) );
  INV_X1 U7134 ( .A(n10000), .ZN(n8141) );
  NAND2_X1 U7135 ( .A1(n8141), .A2(n8022), .ZN(n9849) );
  NAND2_X1 U7136 ( .A1(n9850), .A2(n9849), .ZN(n9843) );
  NAND2_X1 U7137 ( .A1(n7657), .A2(n9843), .ZN(n7656) );
  NAND2_X1 U7138 ( .A1(n11073), .A2(n8141), .ZN(n6023) );
  NAND2_X1 U7139 ( .A1(n7656), .A2(n6023), .ZN(n7713) );
  XNOR2_X1 U7140 ( .A(n6025), .B(n6024), .ZN(n7152) );
  NAND2_X1 U7141 ( .A1(n7152), .A2(n9708), .ZN(n6029) );
  OAI21_X1 U7142 ( .B1(n6026), .B2(P1_IR_REG_6__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6027) );
  XNOR2_X1 U7143 ( .A(n6027), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7371) );
  AOI22_X1 U7144 ( .A1(n6153), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6152), .B2(
        n7371), .ZN(n6028) );
  NAND2_X1 U7145 ( .A1(n6029), .A2(n6028), .ZN(n7716) );
  NAND2_X1 U7146 ( .A1(n6167), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6036) );
  NAND2_X1 U7147 ( .A1(n9704), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6035) );
  AND2_X1 U7148 ( .A1(n6031), .A2(n6030), .ZN(n6032) );
  NOR2_X1 U7149 ( .A1(n6044), .A2(n6032), .ZN(n8140) );
  NAND2_X1 U7150 ( .A1(n6312), .A2(n8140), .ZN(n6034) );
  NAND2_X1 U7151 ( .A1(n6066), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6033) );
  OR2_X1 U7152 ( .A1(n7716), .A2(n8235), .ZN(n9856) );
  NAND2_X1 U7153 ( .A1(n7716), .A2(n8235), .ZN(n7724) );
  NAND2_X1 U7154 ( .A1(n9856), .A2(n7724), .ZN(n9852) );
  INV_X1 U7155 ( .A(n8235), .ZN(n9999) );
  XNOR2_X1 U7156 ( .A(n6039), .B(n6038), .ZN(n7158) );
  NAND2_X1 U7157 ( .A1(n7158), .A2(n9708), .ZN(n6043) );
  NAND2_X1 U7158 ( .A1(n6040), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6041) );
  XNOR2_X1 U7159 ( .A(n6041), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7421) );
  AOI22_X1 U7160 ( .A1(n6153), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6152), .B2(
        n7421), .ZN(n6042) );
  NAND2_X1 U7161 ( .A1(n6043), .A2(n6042), .ZN(n8239) );
  NAND2_X1 U7162 ( .A1(n9704), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6049) );
  NAND2_X1 U7163 ( .A1(n6167), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6048) );
  OR2_X1 U7164 ( .A1(n6044), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6045) );
  AND2_X1 U7165 ( .A1(n6055), .A2(n6045), .ZN(n8234) );
  NAND2_X1 U7166 ( .A1(n6312), .A2(n8234), .ZN(n6047) );
  NAND2_X1 U7167 ( .A1(n6066), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6046) );
  OR2_X1 U7168 ( .A1(n8239), .A2(n7962), .ZN(n9883) );
  NAND2_X1 U7169 ( .A1(n8239), .A2(n7962), .ZN(n9859) );
  NAND2_X1 U7170 ( .A1(n9883), .A2(n9859), .ZN(n9858) );
  INV_X1 U7171 ( .A(n7962), .ZN(n9998) );
  NAND2_X1 U7172 ( .A1(n7162), .A2(n9708), .ZN(n6053) );
  XNOR2_X1 U7173 ( .A(n6051), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10044) );
  AOI22_X1 U7174 ( .A1(n6153), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6152), .B2(
        n10044), .ZN(n6052) );
  NAND2_X1 U7175 ( .A1(n6053), .A2(n6052), .ZN(n8299) );
  NAND2_X1 U7176 ( .A1(n9704), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6061) );
  NAND2_X1 U7177 ( .A1(n5132), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6060) );
  NAND2_X1 U7178 ( .A1(n6055), .A2(n6054), .ZN(n6056) );
  AND2_X1 U7179 ( .A1(n6057), .A2(n6056), .ZN(n8296) );
  NAND2_X1 U7180 ( .A1(n6312), .A2(n8296), .ZN(n6059) );
  NAND2_X1 U7181 ( .A1(n6066), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6058) );
  OR2_X1 U7182 ( .A1(n8299), .A2(n9545), .ZN(n9867) );
  NAND2_X1 U7183 ( .A1(n8299), .A2(n9545), .ZN(n9872) );
  NAND2_X1 U7184 ( .A1(n9867), .A2(n9872), .ZN(n7703) );
  NAND2_X1 U7185 ( .A1(n7701), .A2(n7703), .ZN(n7700) );
  INV_X1 U7186 ( .A(n9545), .ZN(n9997) );
  NAND2_X1 U7187 ( .A1(n7700), .A2(n6062), .ZN(n7880) );
  OR2_X1 U7188 ( .A1(n9547), .A2(n9654), .ZN(n9874) );
  NAND2_X1 U7189 ( .A1(n9547), .A2(n9654), .ZN(n9869) );
  NAND2_X1 U7190 ( .A1(n9874), .A2(n9869), .ZN(n9781) );
  NAND2_X1 U7191 ( .A1(n9704), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6070) );
  NAND2_X1 U7192 ( .A1(n6167), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6069) );
  AND2_X1 U7193 ( .A1(n6064), .A2(n6063), .ZN(n6065) );
  NOR2_X1 U7194 ( .A1(n6087), .A2(n6065), .ZN(n9651) );
  NAND2_X1 U7195 ( .A1(n6312), .A2(n9651), .ZN(n6068) );
  NAND2_X1 U7196 ( .A1(n6066), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6067) );
  NAND4_X1 U7197 ( .A1(n6070), .A2(n6069), .A3(n6068), .A4(n6067), .ZN(n9996)
         );
  INV_X1 U7198 ( .A(n9996), .ZN(n6340) );
  XNOR2_X1 U7199 ( .A(n6072), .B(n6071), .ZN(n7187) );
  NAND2_X1 U7200 ( .A1(n7187), .A2(n9708), .ZN(n6076) );
  NAND2_X1 U7201 ( .A1(n6073), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6074) );
  XNOR2_X1 U7202 ( .A(n6074), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7819) );
  AOI22_X1 U7203 ( .A1(n6153), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6152), .B2(
        n7819), .ZN(n6075) );
  NAND2_X1 U7204 ( .A1(n6076), .A2(n6075), .ZN(n9663) );
  XNOR2_X1 U7205 ( .A(n6078), .B(n6077), .ZN(n7255) );
  NAND2_X1 U7206 ( .A1(n7255), .A2(n9708), .ZN(n6085) );
  NAND2_X1 U7207 ( .A1(n6079), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6080) );
  MUX2_X1 U7208 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6080), .S(
        P1_IR_REG_12__SCAN_IN), .Z(n6082) );
  INV_X1 U7209 ( .A(n5860), .ZN(n6081) );
  NAND2_X1 U7210 ( .A1(n6082), .A2(n6081), .ZN(n8434) );
  INV_X1 U7211 ( .A(n8434), .ZN(n6083) );
  AOI22_X1 U7212 ( .A1(n6153), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6152), .B2(
        n6083), .ZN(n6084) );
  NAND2_X1 U7213 ( .A1(n5131), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6092) );
  NAND2_X1 U7214 ( .A1(n9704), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6091) );
  NOR2_X1 U7215 ( .A1(n6087), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6088) );
  OR2_X1 U7216 ( .A1(n6102), .A2(n6088), .ZN(n9572) );
  INV_X1 U7217 ( .A(n9572), .ZN(n8107) );
  NAND2_X1 U7218 ( .A1(n6312), .A2(n8107), .ZN(n6090) );
  NAND2_X1 U7219 ( .A1(n6066), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6089) );
  NAND4_X1 U7220 ( .A1(n6092), .A2(n6091), .A3(n6090), .A4(n6089), .ZN(n11087)
         );
  INV_X1 U7221 ( .A(n11087), .ZN(n7914) );
  NAND2_X1 U7222 ( .A1(n6094), .A2(n5172), .ZN(n8199) );
  XNOR2_X1 U7223 ( .A(n6096), .B(n6095), .ZN(n7332) );
  NAND2_X1 U7224 ( .A1(n7332), .A2(n9708), .ZN(n6101) );
  NOR2_X1 U7225 ( .A1(n5860), .A2(n6098), .ZN(n6097) );
  MUX2_X1 U7226 ( .A(n6098), .B(n6097), .S(P1_IR_REG_13__SCAN_IN), .Z(n6099)
         );
  NOR2_X1 U7227 ( .A1(n6099), .A2(n6360), .ZN(n10049) );
  AOI22_X1 U7228 ( .A1(n6153), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6152), .B2(
        n10049), .ZN(n6100) );
  NAND2_X1 U7229 ( .A1(n6167), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6108) );
  NAND2_X1 U7230 ( .A1(n9704), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6107) );
  NOR2_X1 U7231 ( .A1(n6102), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n6103) );
  OR2_X1 U7232 ( .A1(n6104), .A2(n6103), .ZN(n9631) );
  INV_X1 U7233 ( .A(n9631), .ZN(n8200) );
  NAND2_X1 U7234 ( .A1(n6312), .A2(n8200), .ZN(n6106) );
  NAND2_X1 U7235 ( .A1(n6066), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6105) );
  NAND4_X1 U7236 ( .A1(n6108), .A2(n6107), .A3(n6106), .A4(n6105), .ZN(n10415)
         );
  NAND2_X1 U7237 ( .A1(n8207), .A2(n10415), .ZN(n6109) );
  INV_X1 U7238 ( .A(n10415), .ZN(n9571) );
  OR2_X1 U7239 ( .A1(n9527), .A2(n9692), .ZN(n9903) );
  NAND2_X1 U7240 ( .A1(n9527), .A2(n9692), .ZN(n9905) );
  NAND2_X1 U7241 ( .A1(n9903), .A2(n9905), .ZN(n9787) );
  NAND2_X1 U7242 ( .A1(n9695), .A2(n9523), .ZN(n9910) );
  NAND2_X1 U7243 ( .A1(n10398), .A2(n10389), .ZN(n9913) );
  NAND2_X1 U7244 ( .A1(n9914), .A2(n9913), .ZN(n9771) );
  XNOR2_X1 U7245 ( .A(n6144), .B(n6122), .ZN(n7739) );
  NAND2_X1 U7246 ( .A1(n7739), .A2(n9708), .ZN(n6116) );
  NAND2_X1 U7247 ( .A1(n6111), .A2(n6110), .ZN(n6112) );
  NAND2_X1 U7248 ( .A1(n5210), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6114) );
  XNOR2_X1 U7249 ( .A(n6114), .B(P1_IR_REG_17__SCAN_IN), .ZN(n10078) );
  AOI22_X1 U7250 ( .A1(n6153), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6152), .B2(
        n10078), .ZN(n6115) );
  NAND2_X1 U7251 ( .A1(n5131), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6121) );
  NAND2_X1 U7252 ( .A1(n6066), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6120) );
  OAI21_X1 U7253 ( .B1(n6117), .B2(P1_REG3_REG_17__SCAN_IN), .A(n6134), .ZN(
        n9605) );
  INV_X1 U7254 ( .A(n9605), .ZN(n8531) );
  NAND2_X1 U7255 ( .A1(n6312), .A2(n8531), .ZN(n6119) );
  NAND2_X1 U7256 ( .A1(n9704), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6118) );
  NAND2_X1 U7257 ( .A1(n8530), .A2(n10297), .ZN(n9724) );
  NAND2_X1 U7258 ( .A1(n9920), .A2(n9724), .ZN(n9792) );
  NAND2_X1 U7259 ( .A1(n8525), .A2(n5748), .ZN(n10293) );
  NAND2_X1 U7260 ( .A1(n6124), .A2(n6123), .ZN(n6126) );
  NAND2_X1 U7261 ( .A1(n7793), .A2(n9708), .ZN(n6132) );
  INV_X1 U7262 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6127) );
  INV_X1 U7263 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6128) );
  NAND2_X1 U7264 ( .A1(n6129), .A2(n6128), .ZN(n6149) );
  OR2_X1 U7265 ( .A1(n6129), .A2(n6128), .ZN(n6130) );
  AND2_X1 U7266 ( .A1(n6149), .A2(n6130), .ZN(n10096) );
  AOI22_X1 U7267 ( .A1(n6153), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6152), .B2(
        n10096), .ZN(n6131) );
  NAND2_X1 U7268 ( .A1(n5132), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6139) );
  NAND2_X1 U7269 ( .A1(n6066), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6138) );
  INV_X1 U7270 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6135) );
  AOI21_X1 U7271 ( .B1(n6135), .B2(n6134), .A(n6133), .ZN(n10302) );
  NAND2_X1 U7272 ( .A1(n6312), .A2(n10302), .ZN(n6137) );
  NAND2_X1 U7273 ( .A1(n9704), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6136) );
  NAND4_X1 U7274 ( .A1(n6139), .A2(n6138), .A3(n6137), .A4(n6136), .ZN(n10282)
         );
  NAND2_X1 U7275 ( .A1(n10305), .A2(n6140), .ZN(n6141) );
  NAND2_X1 U7276 ( .A1(n10293), .A2(n6141), .ZN(n6142) );
  NAND2_X1 U7277 ( .A1(n6144), .A2(n6143), .ZN(n6146) );
  NAND2_X1 U7278 ( .A1(n7846), .A2(n9708), .ZN(n6155) );
  NAND2_X1 U7279 ( .A1(n6149), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6151) );
  AOI22_X1 U7280 ( .A1(n6153), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9987), .B2(
        n6152), .ZN(n6154) );
  NAND2_X1 U7281 ( .A1(n9704), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6162) );
  NAND2_X1 U7282 ( .A1(n6167), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n6161) );
  INV_X1 U7283 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6157) );
  NAND2_X1 U7284 ( .A1(n6157), .A2(n6156), .ZN(n6158) );
  AND2_X1 U7285 ( .A1(n6158), .A2(n6169), .ZN(n10284) );
  NAND2_X1 U7286 ( .A1(n6312), .A2(n10284), .ZN(n6160) );
  NAND2_X1 U7287 ( .A1(n6066), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6159) );
  NAND4_X1 U7288 ( .A1(n6162), .A2(n6161), .A3(n6160), .A4(n6159), .ZN(n10265)
         );
  OR2_X1 U7289 ( .A1(n10379), .A2(n10265), .ZN(n9770) );
  XNOR2_X1 U7290 ( .A(n6164), .B(n6163), .ZN(n7845) );
  NAND2_X1 U7291 ( .A1(n7845), .A2(n9708), .ZN(n6166) );
  OR2_X1 U7292 ( .A1(n9709), .A2(n7850), .ZN(n6165) );
  NAND2_X1 U7293 ( .A1(n9704), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6175) );
  NAND2_X1 U7294 ( .A1(n6167), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6174) );
  INV_X1 U7295 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n6168) );
  NAND2_X1 U7296 ( .A1(n6169), .A2(n6168), .ZN(n6170) );
  AND2_X1 U7297 ( .A1(n6171), .A2(n6170), .ZN(n10264) );
  NAND2_X1 U7298 ( .A1(n6312), .A2(n10264), .ZN(n6173) );
  NAND2_X1 U7299 ( .A1(n6066), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6172) );
  NAND4_X1 U7300 ( .A1(n6175), .A2(n6174), .A3(n6173), .A4(n6172), .ZN(n9562)
         );
  NAND2_X1 U7301 ( .A1(n10368), .A2(n9562), .ZN(n10244) );
  NAND2_X1 U7302 ( .A1(n10263), .A2(n10376), .ZN(n9934) );
  NAND2_X1 U7303 ( .A1(n10244), .A2(n9934), .ZN(n10270) );
  NAND2_X1 U7304 ( .A1(n10253), .A2(n10273), .ZN(n9938) );
  NAND2_X1 U7305 ( .A1(n9939), .A2(n9938), .ZN(n10249) );
  OAI21_X1 U7306 ( .B1(n10253), .B2(n10231), .A(n6176), .ZN(n10235) );
  NAND2_X1 U7307 ( .A1(n6179), .A2(SI_21_), .ZN(n6180) );
  MUX2_X1 U7308 ( .A(n8061), .B(n10581), .S(n8604), .Z(n6181) );
  NAND2_X1 U7309 ( .A1(n6181), .A2(n5492), .ZN(n6194) );
  INV_X1 U7310 ( .A(n6181), .ZN(n6182) );
  NAND2_X1 U7311 ( .A1(n6182), .A2(SI_22_), .ZN(n6183) );
  NAND2_X1 U7312 ( .A1(n6194), .A2(n6183), .ZN(n6195) );
  XNOR2_X1 U7313 ( .A(n6196), .B(n6195), .ZN(n8059) );
  NAND2_X1 U7314 ( .A1(n8059), .A2(n9708), .ZN(n6185) );
  OR2_X1 U7315 ( .A1(n9709), .A2(n10581), .ZN(n6184) );
  NAND2_X1 U7316 ( .A1(n5132), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6192) );
  NAND2_X1 U7317 ( .A1(n6066), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6191) );
  INV_X1 U7318 ( .A(n6187), .ZN(n6186) );
  INV_X1 U7319 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9642) );
  NAND2_X1 U7320 ( .A1(n6187), .A2(n9642), .ZN(n6188) );
  AND2_X1 U7321 ( .A1(n6209), .A2(n6188), .ZN(n10238) );
  NAND2_X1 U7322 ( .A1(n6312), .A2(n10238), .ZN(n6190) );
  NAND2_X1 U7323 ( .A1(n9704), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6189) );
  NAND2_X1 U7324 ( .A1(n10237), .A2(n10248), .ZN(n9720) );
  NAND2_X1 U7325 ( .A1(n10208), .A2(n9720), .ZN(n10234) );
  NAND2_X1 U7326 ( .A1(n10453), .A2(n10248), .ZN(n6193) );
  MUX2_X1 U7327 ( .A(n8120), .B(n8116), .S(n8604), .Z(n6197) );
  INV_X1 U7328 ( .A(SI_23_), .ZN(n10669) );
  NAND2_X1 U7329 ( .A1(n6197), .A2(n10669), .ZN(n6233) );
  INV_X1 U7330 ( .A(n6197), .ZN(n6198) );
  NAND2_X1 U7331 ( .A1(n6198), .A2(SI_23_), .ZN(n6199) );
  NAND2_X1 U7332 ( .A1(n6233), .A2(n6199), .ZN(n6201) );
  NAND2_X1 U7333 ( .A1(n6200), .A2(n6201), .ZN(n6204) );
  INV_X1 U7334 ( .A(n6201), .ZN(n6202) );
  NAND2_X1 U7335 ( .A1(n6204), .A2(n6235), .ZN(n8117) );
  NAND2_X1 U7336 ( .A1(n8117), .A2(n9708), .ZN(n6206) );
  OR2_X1 U7337 ( .A1(n9709), .A2(n8116), .ZN(n6205) );
  NAND2_X1 U7338 ( .A1(n9704), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6214) );
  NAND2_X1 U7339 ( .A1(n5131), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6213) );
  INV_X1 U7340 ( .A(n6209), .ZN(n6207) );
  NAND2_X1 U7341 ( .A1(n6207), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6224) );
  INV_X1 U7342 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6208) );
  NAND2_X1 U7343 ( .A1(n6209), .A2(n6208), .ZN(n6210) );
  AND2_X1 U7344 ( .A1(n6224), .A2(n6210), .ZN(n10214) );
  NAND2_X1 U7345 ( .A1(n6312), .A2(n10214), .ZN(n6212) );
  NAND2_X1 U7346 ( .A1(n6066), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6211) );
  NAND4_X1 U7347 ( .A1(n6214), .A2(n6213), .A3(n6212), .A4(n6211), .ZN(n10230)
         );
  NAND2_X1 U7348 ( .A1(n10222), .A2(n10230), .ZN(n6215) );
  NAND2_X1 U7349 ( .A1(n6235), .A2(n6233), .ZN(n6219) );
  INV_X1 U7350 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8195) );
  MUX2_X1 U7351 ( .A(n8195), .B(n10773), .S(n8604), .Z(n6216) );
  INV_X1 U7352 ( .A(SI_24_), .ZN(n10493) );
  NAND2_X1 U7353 ( .A1(n6216), .A2(n10493), .ZN(n6232) );
  INV_X1 U7354 ( .A(n6216), .ZN(n6217) );
  NAND2_X1 U7355 ( .A1(n6217), .A2(SI_24_), .ZN(n6236) );
  AND2_X1 U7356 ( .A1(n6232), .A2(n6236), .ZN(n6218) );
  NAND2_X1 U7357 ( .A1(n8194), .A2(n9708), .ZN(n6221) );
  OR2_X1 U7358 ( .A1(n9709), .A2(n10773), .ZN(n6220) );
  NAND2_X1 U7359 ( .A1(n9704), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6229) );
  NAND2_X1 U7360 ( .A1(n5132), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6228) );
  INV_X1 U7361 ( .A(n6224), .ZN(n6222) );
  NAND2_X1 U7362 ( .A1(n6222), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6243) );
  INV_X1 U7363 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6223) );
  NAND2_X1 U7364 ( .A1(n6224), .A2(n6223), .ZN(n6225) );
  AND2_X1 U7365 ( .A1(n6243), .A2(n6225), .ZN(n10202) );
  NAND2_X1 U7366 ( .A1(n6312), .A2(n10202), .ZN(n6227) );
  NAND2_X1 U7367 ( .A1(n6066), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6226) );
  NOR2_X1 U7368 ( .A1(n10445), .A2(n10217), .ZN(n6230) );
  NAND2_X1 U7369 ( .A1(n10445), .A2(n10217), .ZN(n6231) );
  AND2_X1 U7370 ( .A1(n6233), .A2(n6232), .ZN(n6234) );
  NAND2_X1 U7371 ( .A1(n6235), .A2(n6234), .ZN(n6237) );
  INV_X1 U7372 ( .A(n6251), .ZN(n6238) );
  INV_X1 U7373 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8229) );
  MUX2_X1 U7374 ( .A(n8229), .B(n10775), .S(n8604), .Z(n6252) );
  XNOR2_X1 U7375 ( .A(n6252), .B(SI_25_), .ZN(n6250) );
  XNOR2_X1 U7376 ( .A(n6238), .B(n6250), .ZN(n8228) );
  NAND2_X1 U7377 ( .A1(n8228), .A2(n9708), .ZN(n6240) );
  OR2_X1 U7378 ( .A1(n9709), .A2(n10775), .ZN(n6239) );
  NAND2_X1 U7379 ( .A1(n6167), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6248) );
  NAND2_X1 U7380 ( .A1(n6066), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6247) );
  INV_X1 U7381 ( .A(n6243), .ZN(n6241) );
  NAND2_X1 U7382 ( .A1(n6241), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6263) );
  INV_X1 U7383 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6242) );
  NAND2_X1 U7384 ( .A1(n6243), .A2(n6242), .ZN(n6244) );
  AND2_X1 U7385 ( .A1(n6263), .A2(n6244), .ZN(n10186) );
  NAND2_X1 U7386 ( .A1(n6312), .A2(n10186), .ZN(n6246) );
  NAND2_X1 U7387 ( .A1(n9704), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6245) );
  NAND4_X1 U7388 ( .A1(n6248), .A2(n6247), .A3(n6246), .A4(n6245), .ZN(n10325)
         );
  NOR2_X1 U7389 ( .A1(n10192), .A2(n10325), .ZN(n6249) );
  INV_X1 U7390 ( .A(n6252), .ZN(n6253) );
  NAND2_X1 U7391 ( .A1(n6253), .A2(SI_25_), .ZN(n6254) );
  INV_X1 U7392 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8416) );
  MUX2_X1 U7393 ( .A(n8416), .B(n10485), .S(n8604), .Z(n6256) );
  NAND2_X1 U7394 ( .A1(n6256), .A2(n10673), .ZN(n6271) );
  INV_X1 U7395 ( .A(n6256), .ZN(n6257) );
  NAND2_X1 U7396 ( .A1(n6257), .A2(SI_26_), .ZN(n6258) );
  NAND2_X1 U7397 ( .A1(n6271), .A2(n6258), .ZN(n6272) );
  NAND2_X1 U7398 ( .A1(n8414), .A2(n9708), .ZN(n6260) );
  OR2_X1 U7399 ( .A1(n9709), .A2(n10485), .ZN(n6259) );
  NAND2_X1 U7400 ( .A1(n5131), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6268) );
  NAND2_X1 U7401 ( .A1(n6066), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6267) );
  INV_X1 U7402 ( .A(n6263), .ZN(n6261) );
  NAND2_X1 U7403 ( .A1(n6261), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6281) );
  INV_X1 U7404 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6262) );
  NAND2_X1 U7405 ( .A1(n6263), .A2(n6262), .ZN(n6264) );
  NAND2_X1 U7406 ( .A1(n6312), .A2(n10171), .ZN(n6266) );
  NAND2_X1 U7407 ( .A1(n9704), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6265) );
  OR2_X1 U7408 ( .A1(n10178), .A2(n10317), .ZN(n9961) );
  NAND2_X1 U7409 ( .A1(n10178), .A2(n10317), .ZN(n9959) );
  NAND2_X1 U7410 ( .A1(n9961), .A2(n9959), .ZN(n6346) );
  NAND2_X1 U7411 ( .A1(n10170), .A2(n6346), .ZN(n6270) );
  NAND2_X1 U7412 ( .A1(n10178), .A2(n10334), .ZN(n6269) );
  INV_X1 U7413 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n6772) );
  INV_X1 U7414 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8451) );
  MUX2_X1 U7415 ( .A(n6772), .B(n8451), .S(n8604), .Z(n6274) );
  INV_X1 U7416 ( .A(SI_27_), .ZN(n10676) );
  NAND2_X1 U7417 ( .A1(n6274), .A2(n10676), .ZN(n6290) );
  INV_X1 U7418 ( .A(n6274), .ZN(n6275) );
  NAND2_X1 U7419 ( .A1(n6275), .A2(SI_27_), .ZN(n6276) );
  NAND2_X1 U7420 ( .A1(n8380), .A2(n9708), .ZN(n6278) );
  OR2_X1 U7421 ( .A1(n9709), .A2(n8451), .ZN(n6277) );
  NAND2_X1 U7422 ( .A1(n5132), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6286) );
  NAND2_X1 U7423 ( .A1(n6066), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6285) );
  INV_X1 U7424 ( .A(n6281), .ZN(n6279) );
  NAND2_X1 U7425 ( .A1(n6279), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n6294) );
  INV_X1 U7426 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6280) );
  NAND2_X1 U7427 ( .A1(n6281), .A2(n6280), .ZN(n6282) );
  NAND2_X1 U7428 ( .A1(n6312), .A2(n10158), .ZN(n6284) );
  NAND2_X1 U7429 ( .A1(n9704), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6283) );
  OR2_X1 U7430 ( .A1(n10157), .A2(n10174), .ZN(n9962) );
  NAND2_X1 U7431 ( .A1(n10157), .A2(n10174), .ZN(n9963) );
  INV_X1 U7432 ( .A(n10153), .ZN(n6287) );
  NAND2_X1 U7433 ( .A1(n10434), .A2(n10174), .ZN(n6398) );
  MUX2_X1 U7434 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n8604), .Z(n6304) );
  INV_X1 U7435 ( .A(SI_28_), .ZN(n6305) );
  XNOR2_X1 U7436 ( .A(n6304), .B(n6305), .ZN(n6302) );
  NAND2_X1 U7437 ( .A1(n8482), .A2(n9708), .ZN(n6292) );
  INV_X1 U7438 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10768) );
  OR2_X1 U7439 ( .A1(n9709), .A2(n10768), .ZN(n6291) );
  NAND2_X1 U7440 ( .A1(n9704), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6299) );
  NAND2_X1 U7441 ( .A1(n5131), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6298) );
  INV_X1 U7442 ( .A(n6294), .ZN(n6293) );
  NAND2_X1 U7443 ( .A1(n6293), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n6311) );
  INV_X1 U7444 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8712) );
  NAND2_X1 U7445 ( .A1(n6294), .A2(n8712), .ZN(n6295) );
  NAND2_X1 U7446 ( .A1(n6312), .A2(n8713), .ZN(n6297) );
  NAND2_X1 U7447 ( .A1(n6066), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6296) );
  OR2_X1 U7448 ( .A1(n8718), .A2(n10316), .ZN(n9969) );
  NAND2_X1 U7449 ( .A1(n8718), .A2(n10316), .ZN(n9968) );
  AND2_X1 U7450 ( .A1(n6398), .A2(n9799), .ZN(n6300) );
  INV_X1 U7451 ( .A(n10316), .ZN(n9995) );
  NAND2_X1 U7452 ( .A1(n8718), .A2(n9995), .ZN(n6301) );
  NAND2_X1 U7453 ( .A1(n6400), .A2(n6301), .ZN(n6317) );
  NAND2_X1 U7454 ( .A1(n6303), .A2(n6302), .ZN(n6308) );
  INV_X1 U7455 ( .A(n6304), .ZN(n6306) );
  NAND2_X1 U7456 ( .A1(n6306), .A2(n6305), .ZN(n6307) );
  INV_X1 U7457 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9514) );
  INV_X1 U7458 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10763) );
  MUX2_X1 U7459 ( .A(n9514), .B(n10763), .S(n8604), .Z(n8596) );
  NAND2_X1 U7460 ( .A1(n8540), .A2(n9708), .ZN(n6310) );
  OR2_X1 U7461 ( .A1(n9709), .A2(n10763), .ZN(n6309) );
  NAND2_X1 U7462 ( .A1(n9704), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6316) );
  NAND2_X1 U7463 ( .A1(n5132), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6315) );
  INV_X1 U7464 ( .A(n6311), .ZN(n10141) );
  NAND2_X1 U7465 ( .A1(n6312), .A2(n10141), .ZN(n6314) );
  NAND2_X1 U7466 ( .A1(n6066), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6313) );
  NAND2_X1 U7467 ( .A1(n10147), .A2(n8714), .ZN(n9975) );
  NAND2_X1 U7468 ( .A1(n6320), .A2(n10830), .ZN(n6319) );
  INV_X1 U7469 ( .A(n6918), .ZN(n6327) );
  NAND2_X1 U7470 ( .A1(n5174), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6322) );
  MUX2_X1 U7471 ( .A(n6322), .B(P1_IR_REG_31__SCAN_IN), .S(n6321), .Z(n6323)
         );
  OR2_X1 U7472 ( .A1(n6921), .A2(n6917), .ZN(n9700) );
  NAND2_X1 U7473 ( .A1(n6918), .A2(n6324), .ZN(n7601) );
  INV_X1 U7474 ( .A(n9758), .ZN(n6325) );
  NAND2_X1 U7475 ( .A1(n6921), .A2(n6325), .ZN(n6326) );
  NAND3_X1 U7476 ( .A1(n9700), .A2(n7601), .A3(n6326), .ZN(n11084) );
  NAND2_X2 U7477 ( .A1(n6918), .A2(n9987), .ZN(n9973) );
  OR2_X1 U7478 ( .A1(n9973), .A2(n9986), .ZN(n11085) );
  NAND2_X1 U7479 ( .A1(n6370), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6330) );
  NAND2_X1 U7480 ( .A1(n6330), .A2(n6329), .ZN(n6352) );
  NAND2_X1 U7481 ( .A1(n6352), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6331) );
  XNOR2_X1 U7482 ( .A(n6331), .B(P1_IR_REG_28__SCAN_IN), .ZN(n7258) );
  INV_X1 U7483 ( .A(n7258), .ZN(n8497) );
  INV_X1 U7484 ( .A(n11024), .ZN(n9725) );
  NAND2_X1 U7485 ( .A1(n5968), .A2(n6934), .ZN(n6333) );
  AND2_X1 U7486 ( .A1(n9831), .A2(n9729), .ZN(n9826) );
  INV_X1 U7487 ( .A(n7549), .ZN(n9773) );
  NAND2_X1 U7488 ( .A1(n9826), .A2(n9773), .ZN(n7560) );
  NAND2_X1 U7489 ( .A1(n7560), .A2(n9834), .ZN(n7681) );
  INV_X1 U7490 ( .A(n9775), .ZN(n7682) );
  NAND2_X1 U7491 ( .A1(n7681), .A2(n7682), .ZN(n7937) );
  INV_X1 U7492 ( .A(n9827), .ZN(n6334) );
  NOR2_X1 U7493 ( .A1(n9847), .A2(n6334), .ZN(n9841) );
  NAND2_X1 U7494 ( .A1(n7937), .A2(n9841), .ZN(n6335) );
  INV_X1 U7495 ( .A(n9850), .ZN(n6336) );
  AND2_X1 U7496 ( .A1(n9883), .A2(n9856), .ZN(n6337) );
  AND2_X1 U7497 ( .A1(n9867), .A2(n6337), .ZN(n9779) );
  NAND2_X1 U7498 ( .A1(n9859), .A2(n7724), .ZN(n9772) );
  NAND3_X1 U7499 ( .A1(n9867), .A2(n9883), .A3(n9772), .ZN(n6338) );
  AND2_X1 U7500 ( .A1(n6338), .A2(n9872), .ZN(n9736) );
  NAND2_X1 U7501 ( .A1(n6339), .A2(n9736), .ZN(n7883) );
  INV_X1 U7502 ( .A(n9781), .ZN(n7884) );
  OR2_X1 U7503 ( .A1(n9663), .A2(n6340), .ZN(n9879) );
  NAND2_X1 U7504 ( .A1(n9663), .A2(n6340), .ZN(n9881) );
  OR2_X1 U7505 ( .A1(n8108), .A2(n7914), .ZN(n9891) );
  NAND2_X1 U7506 ( .A1(n8108), .A2(n7914), .ZN(n9882) );
  NAND2_X1 U7507 ( .A1(n9891), .A2(n9882), .ZN(n8100) );
  OR2_X1 U7508 ( .A1(n8101), .A2(n8100), .ZN(n8103) );
  OR2_X1 U7509 ( .A1(n8207), .A2(n9571), .ZN(n9901) );
  NAND2_X1 U7510 ( .A1(n8207), .A2(n9571), .ZN(n9892) );
  INV_X1 U7511 ( .A(n9787), .ZN(n9896) );
  NAND2_X1 U7512 ( .A1(n6341), .A2(n9905), .ZN(n8456) );
  NAND2_X1 U7513 ( .A1(n8456), .A2(n9909), .ZN(n6342) );
  NAND2_X1 U7514 ( .A1(n6342), .A2(n9910), .ZN(n8485) );
  OR2_X1 U7515 ( .A1(n8485), .A2(n9771), .ZN(n8487) );
  NAND2_X1 U7516 ( .A1(n8487), .A2(n9914), .ZN(n8536) );
  INV_X1 U7517 ( .A(n9792), .ZN(n9916) );
  NAND2_X1 U7518 ( .A1(n8536), .A2(n9916), .ZN(n8535) );
  AND2_X1 U7519 ( .A1(n10305), .A2(n10282), .ZN(n9919) );
  NAND2_X1 U7520 ( .A1(n10385), .A2(n6140), .ZN(n9921) );
  INV_X1 U7521 ( .A(n10265), .ZN(n10367) );
  NAND2_X1 U7522 ( .A1(n10379), .A2(n10367), .ZN(n9928) );
  OR2_X1 U7523 ( .A1(n10379), .A2(n10367), .ZN(n10269) );
  AND2_X1 U7524 ( .A1(n10244), .A2(n10269), .ZN(n9930) );
  AND2_X1 U7525 ( .A1(n9930), .A2(n9939), .ZN(n9746) );
  NAND2_X1 U7526 ( .A1(n10271), .A2(n9746), .ZN(n9763) );
  NAND2_X1 U7527 ( .A1(n9938), .A2(n9934), .ZN(n6343) );
  NAND2_X1 U7528 ( .A1(n6343), .A2(n9939), .ZN(n9721) );
  NAND2_X1 U7529 ( .A1(n9763), .A2(n9721), .ZN(n10226) );
  OR2_X1 U7530 ( .A1(n10226), .A2(n10234), .ZN(n10227) );
  INV_X1 U7531 ( .A(n10230), .ZN(n9643) );
  OR2_X1 U7532 ( .A1(n10222), .A2(n9643), .ZN(n9942) );
  NAND2_X1 U7533 ( .A1(n10222), .A2(n9643), .ZN(n9943) );
  NAND2_X1 U7534 ( .A1(n9942), .A2(n9943), .ZN(n10212) );
  INV_X1 U7535 ( .A(n10208), .ZN(n6344) );
  NOR2_X1 U7536 ( .A1(n10212), .A2(n6344), .ZN(n6345) );
  OR2_X2 U7537 ( .A1(n10201), .A2(n10217), .ZN(n9947) );
  NAND2_X1 U7538 ( .A1(n10201), .A2(n10217), .ZN(n9949) );
  AND2_X2 U7539 ( .A1(n9947), .A2(n9949), .ZN(n10198) );
  OR2_X1 U7540 ( .A1(n10192), .A2(n7080), .ZN(n9952) );
  NAND2_X1 U7541 ( .A1(n10192), .A2(n7080), .ZN(n9950) );
  NAND2_X1 U7542 ( .A1(n9952), .A2(n9950), .ZN(n10184) );
  OR2_X1 U7543 ( .A1(n10183), .A2(n10184), .ZN(n10181) );
  NAND2_X1 U7544 ( .A1(n10181), .A2(n9950), .ZN(n10167) );
  NAND2_X1 U7545 ( .A1(n10167), .A2(n10169), .ZN(n10166) );
  NAND2_X1 U7546 ( .A1(n10166), .A2(n9959), .ZN(n10154) );
  NAND2_X1 U7547 ( .A1(n10154), .A2(n10153), .ZN(n10152) );
  NAND2_X1 U7548 ( .A1(n10152), .A2(n9963), .ZN(n6402) );
  INV_X1 U7549 ( .A(n9968), .ZN(n6347) );
  AOI21_X1 U7550 ( .B1(n6402), .B2(n9965), .A(n6347), .ZN(n6348) );
  INV_X1 U7551 ( .A(n9972), .ZN(n9800) );
  NAND2_X1 U7552 ( .A1(n6327), .A2(n9987), .ZN(n6350) );
  NAND2_X1 U7553 ( .A1(n6328), .A2(n9986), .ZN(n6349) );
  NAND2_X1 U7554 ( .A1(n6351), .A2(n6352), .ZN(n8453) );
  INV_X1 U7555 ( .A(P1_B_REG_SCAN_IN), .ZN(n6353) );
  NOR2_X1 U7556 ( .A1(n8453), .A2(n6353), .ZN(n6354) );
  NOR2_X1 U7557 ( .A1(n10375), .A2(n6354), .ZN(n10130) );
  INV_X1 U7558 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n6357) );
  NAND2_X1 U7559 ( .A1(n6167), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6356) );
  NAND2_X1 U7560 ( .A1(n6066), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6355) );
  OAI211_X1 U7561 ( .C1(n6358), .C2(n6357), .A(n6356), .B(n6355), .ZN(n9994)
         );
  INV_X1 U7562 ( .A(n10222), .ZN(n10449) );
  NAND2_X1 U7563 ( .A1(n11034), .A2(n9725), .ZN(n7693) );
  OR2_X1 U7564 ( .A1(n7693), .A2(n7694), .ZN(n7555) );
  INV_X1 U7565 ( .A(n7716), .ZN(n8147) );
  AND2_X1 U7566 ( .A1(n7714), .A2(n8147), .ZN(n7733) );
  INV_X1 U7567 ( .A(n8239), .ZN(n8083) );
  NAND2_X1 U7568 ( .A1(n7733), .A2(n8083), .ZN(n7732) );
  OR2_X1 U7569 ( .A1(n7732), .A2(n8299), .ZN(n7881) );
  NOR2_X1 U7570 ( .A1(n7881), .A2(n9547), .ZN(n7910) );
  AND2_X1 U7571 ( .A1(n8458), .A2(n10409), .ZN(n8457) );
  OR2_X2 U7572 ( .A1(n10261), .A2(n10253), .ZN(n10251) );
  NOR2_X1 U7573 ( .A1(n10237), .A2(n10251), .ZN(n10236) );
  AND2_X1 U7574 ( .A1(n10449), .A2(n10236), .ZN(n10200) );
  NAND2_X1 U7575 ( .A1(n6910), .A2(n6403), .ZN(n10134) );
  OAI211_X1 U7576 ( .C1(n6910), .C2(n6403), .A(n10400), .B(n10134), .ZN(n10144) );
  NAND2_X1 U7577 ( .A1(n6360), .A2(n6359), .ZN(n6362) );
  NAND2_X1 U7578 ( .A1(n6362), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6361) );
  MUX2_X1 U7579 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6361), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n6363) );
  NAND2_X1 U7580 ( .A1(n8244), .A2(P1_B_REG_SCAN_IN), .ZN(n6367) );
  NAND3_X1 U7581 ( .A1(n10830), .A2(n6387), .A3(n10835), .ZN(n6364) );
  INV_X1 U7582 ( .A(n6386), .ZN(n6392) );
  MUX2_X1 U7583 ( .A(n6367), .B(P1_B_REG_SCAN_IN), .S(n6386), .Z(n6373) );
  NAND2_X1 U7584 ( .A1(n6368), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6369) );
  MUX2_X1 U7585 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6369), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n6371) );
  NAND2_X1 U7586 ( .A1(n6371), .A2(n6370), .ZN(n8417) );
  INV_X1 U7587 ( .A(n8417), .ZN(n6372) );
  OR2_X1 U7588 ( .A1(n10466), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6374) );
  NAND2_X1 U7589 ( .A1(n8417), .A2(n8244), .ZN(n10467) );
  NAND2_X1 U7590 ( .A1(n6374), .A2(n10467), .ZN(n7105) );
  NOR4_X1 U7591 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6383) );
  NOR4_X1 U7592 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6382) );
  OR4_X1 U7593 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .A3(
        P1_D_REG_30__SCAN_IN), .A4(P1_D_REG_29__SCAN_IN), .ZN(n6380) );
  NOR4_X1 U7594 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6378) );
  NOR4_X1 U7595 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6377) );
  NOR4_X1 U7596 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n6376) );
  NOR4_X1 U7597 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6375) );
  NAND4_X1 U7598 ( .A1(n6378), .A2(n6377), .A3(n6376), .A4(n6375), .ZN(n6379)
         );
  NOR4_X1 U7599 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        n6380), .A4(n6379), .ZN(n6381) );
  AND3_X1 U7600 ( .A1(n6383), .A2(n6382), .A3(n6381), .ZN(n6384) );
  AND2_X1 U7601 ( .A1(n7126), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6391) );
  NAND2_X1 U7602 ( .A1(n6388), .A2(n6387), .ZN(n6389) );
  NAND2_X1 U7603 ( .A1(n6389), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6390) );
  NAND2_X1 U7604 ( .A1(n10468), .A2(n7117), .ZN(n6406) );
  INV_X1 U7605 ( .A(n6406), .ZN(n7304) );
  OR2_X1 U7606 ( .A1(n10466), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6394) );
  NAND2_X1 U7607 ( .A1(n6392), .A2(n8417), .ZN(n6393) );
  NAND2_X1 U7608 ( .A1(n6394), .A2(n6393), .ZN(n7107) );
  INV_X1 U7609 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6395) );
  NOR2_X1 U7610 ( .A1(n11114), .A2(n6395), .ZN(n6396) );
  AND2_X1 U7611 ( .A1(n6399), .A2(n6398), .ZN(n6401) );
  XNOR2_X1 U7612 ( .A(n6402), .B(n9965), .ZN(n8674) );
  OAI22_X1 U7613 ( .A1(n10174), .A2(n10388), .B1(n8714), .B2(n10375), .ZN(
        n6404) );
  AOI211_X1 U7614 ( .C1(n8718), .C2(n10155), .A(n10300), .B(n6403), .ZN(n8673)
         );
  OAI21_X1 U7615 ( .B1(n8677), .B2(n11023), .A(n6405), .ZN(n6413) );
  NOR2_X1 U7616 ( .A1(n7107), .A2(n6406), .ZN(n6407) );
  MUX2_X1 U7617 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n6413), .S(n11110), .Z(n6409) );
  INV_X1 U7618 ( .A(n6409), .ZN(n6412) );
  NAND2_X1 U7619 ( .A1(n8718), .A2(n6410), .ZN(n6411) );
  NAND2_X1 U7620 ( .A1(n6412), .A2(n6411), .ZN(P1_U3550) );
  MUX2_X1 U7621 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n6413), .S(n11114), .Z(n6414) );
  INV_X1 U7622 ( .A(n6414), .ZN(n6417) );
  NAND2_X1 U7623 ( .A1(n8718), .A2(n6415), .ZN(n6416) );
  NAND2_X1 U7624 ( .A1(n6417), .A2(n6416), .ZN(P1_U3518) );
  INV_X1 U7625 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6426) );
  INV_X1 U7626 ( .A(n6431), .ZN(n8630) );
  BUF_X4 U7627 ( .A(n6476), .Z(n7810) );
  NAND2_X1 U7628 ( .A1(n7810), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6438) );
  BUF_X4 U7629 ( .A(n6465), .Z(n7811) );
  NAND2_X1 U7630 ( .A1(n7811), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6437) );
  NAND2_X1 U7631 ( .A1(n6498), .A2(n6432), .ZN(n6508) );
  OR2_X1 U7632 ( .A1(n6432), .A2(n6498), .ZN(n6433) );
  NAND2_X1 U7633 ( .A1(n6508), .A2(n6433), .ZN(n7802) );
  NAND2_X1 U7634 ( .A1(n5125), .A2(n7802), .ZN(n6436) );
  AND2_X2 U7635 ( .A1(n8630), .A2(n6434), .ZN(n6475) );
  NAND2_X1 U7636 ( .A1(n6839), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6435) );
  NAND2_X2 U7637 ( .A1(n7130), .A2(n7134), .ZN(n6492) );
  OR2_X1 U7638 ( .A1(n6492), .A2(n7138), .ZN(n6452) );
  INV_X1 U7639 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n7139) );
  OR2_X1 U7640 ( .A1(n8841), .A2(n7139), .ZN(n6451) );
  NAND2_X1 U7641 ( .A1(n6491), .A2(n6558), .ZN(n6447) );
  NAND2_X1 U7642 ( .A1(n6447), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6504) );
  INV_X1 U7643 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6448) );
  NAND2_X1 U7644 ( .A1(n6504), .A2(n6448), .ZN(n6449) );
  NAND2_X1 U7645 ( .A1(n6449), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6515) );
  XNOR2_X1 U7646 ( .A(n6515), .B(P2_IR_REG_5__SCAN_IN), .ZN(n7244) );
  NAND2_X1 U7647 ( .A1(n6683), .A2(n7244), .ZN(n6450) );
  INV_X1 U7648 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n8668) );
  OR2_X1 U7649 ( .A1(n6493), .A2(n8668), .ZN(n6459) );
  OAI211_X1 U7650 ( .C1(n7130), .C2(n5128), .A(n6460), .B(n6459), .ZN(n7485)
         );
  NAND2_X1 U7651 ( .A1(n6477), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6464) );
  NAND2_X1 U7652 ( .A1(n6475), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6462) );
  NAND2_X1 U7653 ( .A1(n6465), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6461) );
  NAND2_X1 U7654 ( .A1(n6477), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n6468) );
  NAND2_X1 U7655 ( .A1(n6465), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6466) );
  NAND2_X1 U7656 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6470) );
  MUX2_X1 U7657 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6470), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n6472) );
  INV_X1 U7658 ( .A(n7205), .ZN(n6471) );
  OAI22_X1 U7659 ( .A1(n6492), .A2(n7136), .B1(n7130), .B2(n5231), .ZN(n6473)
         );
  INV_X1 U7660 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n7133) );
  NAND2_X1 U7661 ( .A1(n6465), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6481) );
  NAND2_X1 U7662 ( .A1(n6475), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6480) );
  NAND2_X1 U7663 ( .A1(n6476), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6479) );
  NAND2_X1 U7664 ( .A1(n5125), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6478) );
  INV_X1 U7665 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7204) );
  NAND2_X1 U7666 ( .A1(n7134), .A2(SI_0_), .ZN(n6483) );
  INV_X1 U7667 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6482) );
  NAND2_X1 U7668 ( .A1(n6483), .A2(n6482), .ZN(n6485) );
  NAND2_X1 U7669 ( .A1(n6485), .A2(n6484), .ZN(n9517) );
  MUX2_X1 U7670 ( .A(n7204), .B(n9517), .S(n7130), .Z(n7593) );
  NOR2_X1 U7671 ( .A1(n9051), .A2(n8032), .ZN(n7468) );
  NAND2_X1 U7672 ( .A1(n9050), .A2(n7976), .ZN(n8896) );
  INV_X1 U7673 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6486) );
  NAND2_X1 U7674 ( .A1(n5125), .A2(n6486), .ZN(n6490) );
  NAND2_X1 U7675 ( .A1(n7811), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6489) );
  NAND2_X1 U7676 ( .A1(n6839), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6488) );
  NAND2_X1 U7677 ( .A1(n6476), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6487) );
  NOR2_X1 U7678 ( .A1(n7448), .A2(n7839), .ZN(n6497) );
  OR2_X1 U7679 ( .A1(n6492), .A2(n8624), .ZN(n6495) );
  INV_X1 U7680 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n8625) );
  OR2_X1 U7681 ( .A1(n8841), .A2(n8625), .ZN(n6494) );
  OAI211_X1 U7682 ( .C1(n7130), .C2(n8623), .A(n6495), .B(n6494), .ZN(n6812)
         );
  INV_X1 U7683 ( .A(n7448), .ZN(n6496) );
  NAND2_X1 U7684 ( .A1(n7810), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6503) );
  NAND2_X1 U7685 ( .A1(n7811), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6502) );
  AND2_X1 U7686 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6499) );
  OR2_X1 U7687 ( .A1(n6499), .A2(n6498), .ZN(n8039) );
  NAND2_X1 U7688 ( .A1(n5125), .A2(n8039), .ZN(n6501) );
  NAND2_X1 U7689 ( .A1(n6839), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6500) );
  INV_X1 U7690 ( .A(n5127), .ZN(n10982) );
  OR2_X1 U7691 ( .A1(n6492), .A2(n6505), .ZN(n6507) );
  OR2_X1 U7692 ( .A1(n6493), .A2(n5368), .ZN(n6506) );
  OAI211_X1 U7693 ( .C1(n7130), .C2(n10982), .A(n6507), .B(n6506), .ZN(n8040)
         );
  NAND2_X1 U7694 ( .A1(n7798), .A2(n8040), .ZN(n8901) );
  INV_X1 U7695 ( .A(n8040), .ZN(n7836) );
  NAND2_X1 U7696 ( .A1(n9048), .A2(n7836), .ZN(n8906) );
  NAND2_X1 U7697 ( .A1(n7810), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6513) );
  NAND2_X1 U7698 ( .A1(n7811), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6512) );
  NAND2_X1 U7699 ( .A1(n6508), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6509) );
  NAND2_X1 U7700 ( .A1(n6523), .A2(n6509), .ZN(n8129) );
  NAND2_X1 U7701 ( .A1(n5125), .A2(n8129), .ZN(n6511) );
  NAND2_X1 U7702 ( .A1(n6839), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6510) );
  OR2_X1 U7703 ( .A1(n7142), .A2(n6492), .ZN(n6519) );
  INV_X1 U7704 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6514) );
  NAND2_X1 U7705 ( .A1(n6515), .A2(n6514), .ZN(n6516) );
  NAND2_X1 U7706 ( .A1(n6516), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6530) );
  XNOR2_X1 U7707 ( .A(n6530), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7287) );
  NAND2_X1 U7708 ( .A1(n6683), .A2(n7287), .ZN(n6518) );
  INV_X1 U7709 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7143) );
  OR2_X1 U7710 ( .A1(n8841), .A2(n7143), .ZN(n6517) );
  NAND2_X1 U7711 ( .A1(n6520), .A2(n8130), .ZN(n6521) );
  NAND2_X1 U7712 ( .A1(n8150), .A2(n8160), .ZN(n6522) );
  NAND2_X1 U7713 ( .A1(n7811), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6528) );
  NAND2_X1 U7714 ( .A1(n6839), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6527) );
  AND2_X1 U7715 ( .A1(n6523), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6524) );
  OR2_X1 U7716 ( .A1(n6524), .A2(n6544), .ZN(n8155) );
  NAND2_X1 U7717 ( .A1(n5125), .A2(n8155), .ZN(n6526) );
  NAND2_X1 U7718 ( .A1(n7810), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6525) );
  NAND4_X1 U7719 ( .A1(n6528), .A2(n6527), .A3(n6526), .A4(n6525), .ZN(n9046)
         );
  NAND2_X1 U7720 ( .A1(n7152), .A2(n8838), .ZN(n6533) );
  NAND2_X1 U7721 ( .A1(n6530), .A2(n6529), .ZN(n6531) );
  NAND2_X1 U7722 ( .A1(n6531), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6538) );
  AOI22_X1 U7723 ( .A1(n8837), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6683), .B2(
        n7867), .ZN(n6532) );
  XNOR2_X1 U7724 ( .A(n9046), .B(n8931), .ZN(n8919) );
  NAND2_X1 U7725 ( .A1(n8148), .A2(n8919), .ZN(n6535) );
  NAND2_X1 U7726 ( .A1(n8047), .A2(n8931), .ZN(n6534) );
  NAND2_X1 U7727 ( .A1(n6535), .A2(n6534), .ZN(n8247) );
  NAND2_X1 U7728 ( .A1(n7158), .A2(n8838), .ZN(n6542) );
  NAND2_X1 U7729 ( .A1(n6538), .A2(n6537), .ZN(n6539) );
  NAND2_X1 U7730 ( .A1(n6539), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6540) );
  INV_X1 U7731 ( .A(n7997), .ZN(n7876) );
  AOI22_X1 U7732 ( .A1(n8837), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6683), .B2(
        n7876), .ZN(n6541) );
  NAND2_X1 U7733 ( .A1(n7810), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6549) );
  NAND2_X1 U7734 ( .A1(n7811), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6548) );
  NOR2_X1 U7735 ( .A1(n6544), .A2(n6543), .ZN(n6545) );
  OR2_X1 U7736 ( .A1(n6564), .A2(n6545), .ZN(n8250) );
  NAND2_X1 U7737 ( .A1(n6728), .A2(n8250), .ZN(n6547) );
  NAND2_X1 U7738 ( .A1(n6839), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6546) );
  NAND4_X1 U7739 ( .A1(n6549), .A2(n6548), .A3(n6547), .A4(n6546), .ZN(n9044)
         );
  NAND2_X1 U7740 ( .A1(n8290), .A2(n9044), .ZN(n8916) );
  INV_X1 U7741 ( .A(n9044), .ZN(n8151) );
  INV_X1 U7742 ( .A(n8290), .ZN(n8251) );
  NAND2_X1 U7743 ( .A1(n8151), .A2(n8251), .ZN(n8930) );
  NAND2_X1 U7744 ( .A1(n8916), .A2(n8930), .ZN(n8855) );
  NAND2_X1 U7745 ( .A1(n7166), .A2(n8838), .ZN(n6552) );
  NAND2_X1 U7746 ( .A1(n6588), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6550) );
  XNOR2_X1 U7747 ( .A(n6550), .B(n6589), .ZN(n8269) );
  INV_X1 U7748 ( .A(n8269), .ZN(n8191) );
  AOI22_X1 U7749 ( .A1(n8837), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6683), .B2(
        n8191), .ZN(n6551) );
  NAND2_X1 U7750 ( .A1(n7811), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6557) );
  NAND2_X1 U7751 ( .A1(n6839), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6556) );
  NAND2_X1 U7752 ( .A1(n6566), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6553) );
  NAND2_X1 U7753 ( .A1(n6582), .A2(n6553), .ZN(n8395) );
  NAND2_X1 U7754 ( .A1(n5125), .A2(n8395), .ZN(n6555) );
  NAND2_X1 U7755 ( .A1(n7810), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6554) );
  NAND4_X1 U7756 ( .A1(n6557), .A2(n6556), .A3(n6555), .A4(n6554), .ZN(n9042)
         );
  NAND2_X1 U7757 ( .A1(n8479), .A2(n9042), .ZN(n8383) );
  INV_X1 U7758 ( .A(n8383), .ZN(n6572) );
  NAND2_X1 U7759 ( .A1(n6561), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6562) );
  XNOR2_X1 U7760 ( .A(n6562), .B(P2_IR_REG_9__SCAN_IN), .ZN(n8183) );
  AOI22_X1 U7761 ( .A1(n8837), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6683), .B2(
        n8183), .ZN(n6563) );
  INV_X1 U7762 ( .A(n8321), .ZN(n8349) );
  NAND2_X1 U7763 ( .A1(n7810), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6570) );
  NAND2_X1 U7764 ( .A1(n7811), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6569) );
  OR2_X1 U7765 ( .A1(n6564), .A2(n10556), .ZN(n6565) );
  NAND2_X1 U7766 ( .A1(n6566), .A2(n6565), .ZN(n8320) );
  NAND2_X1 U7767 ( .A1(n5125), .A2(n8320), .ZN(n6568) );
  NAND2_X1 U7768 ( .A1(n6839), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6567) );
  NAND2_X1 U7769 ( .A1(n8349), .A2(n8390), .ZN(n8387) );
  OR2_X1 U7770 ( .A1(n8479), .A2(n9042), .ZN(n8384) );
  AND2_X1 U7771 ( .A1(n8387), .A2(n8384), .ZN(n6571) );
  INV_X1 U7772 ( .A(n6577), .ZN(n6574) );
  NAND2_X1 U7773 ( .A1(n8321), .A2(n8390), .ZN(n8932) );
  NAND2_X1 U7774 ( .A1(n8920), .A2(n8932), .ZN(n8856) );
  AND2_X1 U7775 ( .A1(n8856), .A2(n8383), .ZN(n6573) );
  AND2_X1 U7776 ( .A1(n8855), .A2(n6576), .ZN(n6575) );
  NAND2_X1 U7777 ( .A1(n8247), .A2(n6575), .ZN(n6581) );
  INV_X1 U7778 ( .A(n6576), .ZN(n6579) );
  NAND2_X1 U7779 ( .A1(n8290), .A2(n8151), .ZN(n8313) );
  AND2_X1 U7780 ( .A1(n8313), .A2(n6577), .ZN(n6578) );
  NAND2_X1 U7781 ( .A1(n7810), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6587) );
  NAND2_X1 U7782 ( .A1(n7811), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6586) );
  AND2_X1 U7783 ( .A1(n6582), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6583) );
  OR2_X1 U7784 ( .A1(n6599), .A2(n6583), .ZN(n8341) );
  NAND2_X1 U7785 ( .A1(n6728), .A2(n8341), .ZN(n6585) );
  NAND2_X1 U7786 ( .A1(n6839), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6584) );
  NAND2_X1 U7787 ( .A1(n6614), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6591) );
  MUX2_X1 U7788 ( .A(n6591), .B(P2_IR_REG_31__SCAN_IN), .S(n6592), .Z(n6593)
         );
  NAND2_X1 U7789 ( .A1(n6593), .A2(n6665), .ZN(n8271) );
  INV_X1 U7790 ( .A(n8271), .ZN(n10998) );
  AOI22_X1 U7791 ( .A1(n8837), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6683), .B2(
        n10998), .ZN(n6594) );
  NAND2_X1 U7792 ( .A1(n7255), .A2(n8838), .ZN(n6598) );
  NAND2_X1 U7793 ( .A1(n6665), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6596) );
  XNOR2_X1 U7794 ( .A(n6596), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8273) );
  AOI22_X1 U7795 ( .A1(n8837), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6683), .B2(
        n8273), .ZN(n6597) );
  NAND2_X1 U7796 ( .A1(n6598), .A2(n6597), .ZN(n8405) );
  NAND2_X1 U7797 ( .A1(n7810), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6604) );
  NAND2_X1 U7798 ( .A1(n7811), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6603) );
  OR2_X1 U7799 ( .A1(n6599), .A2(n10732), .ZN(n6600) );
  NAND2_X1 U7800 ( .A1(n6600), .A2(n6608), .ZN(n8411) );
  NAND2_X1 U7801 ( .A1(n6728), .A2(n8411), .ZN(n6602) );
  NAND2_X1 U7802 ( .A1(n6839), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6601) );
  NAND4_X1 U7803 ( .A1(n6604), .A2(n6603), .A3(n6602), .A4(n6601), .ZN(n9040)
         );
  XNOR2_X1 U7804 ( .A(n8405), .B(n9040), .ZN(n8942) );
  NAND2_X1 U7805 ( .A1(n8405), .A2(n9040), .ZN(n6607) );
  NAND2_X1 U7806 ( .A1(n8367), .A2(n6607), .ZN(n6617) );
  INV_X1 U7807 ( .A(n6617), .ZN(n8505) );
  NAND2_X1 U7808 ( .A1(n7811), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6612) );
  NAND2_X1 U7809 ( .A1(n6839), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6611) );
  NAND2_X1 U7810 ( .A1(n7810), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6610) );
  AOI21_X1 U7811 ( .B1(P2_REG3_REG_13__SCAN_IN), .B2(n6608), .A(n6624), .ZN(
        n8508) );
  INV_X1 U7812 ( .A(n8508), .ZN(n8469) );
  NAND2_X1 U7813 ( .A1(n6728), .A2(n8469), .ZN(n6609) );
  NAND4_X1 U7814 ( .A1(n6612), .A2(n6611), .A3(n6610), .A4(n6609), .ZN(n9039)
         );
  NAND2_X1 U7815 ( .A1(n7332), .A2(n8838), .ZN(n6616) );
  OR2_X1 U7816 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n6613) );
  OAI21_X1 U7817 ( .B1(n6614), .B2(n6613), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6620) );
  XNOR2_X1 U7818 ( .A(n6620), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8579) );
  AOI22_X1 U7819 ( .A1(n8837), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6683), .B2(
        n8579), .ZN(n6615) );
  OAI21_X1 U7820 ( .B1(n8505), .B2(n9374), .A(n6618), .ZN(n9371) );
  NAND2_X1 U7821 ( .A1(n7395), .A2(n8838), .ZN(n6623) );
  INV_X1 U7822 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6619) );
  NAND2_X1 U7823 ( .A1(n6620), .A2(n6619), .ZN(n6621) );
  NAND2_X1 U7824 ( .A1(n6621), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6633) );
  XNOR2_X1 U7825 ( .A(n6633), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8558) );
  AOI22_X1 U7826 ( .A1(n8837), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6683), .B2(
        n8558), .ZN(n6622) );
  NAND2_X1 U7827 ( .A1(n7810), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6629) );
  NAND2_X1 U7828 ( .A1(n7811), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6628) );
  OR2_X1 U7829 ( .A1(n6624), .A2(n10724), .ZN(n6625) );
  NAND2_X1 U7830 ( .A1(n6625), .A2(n6637), .ZN(n9379) );
  NAND2_X1 U7831 ( .A1(n6728), .A2(n9379), .ZN(n6627) );
  NAND2_X1 U7832 ( .A1(n6839), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6626) );
  NAND4_X1 U7833 ( .A1(n6629), .A2(n6628), .A3(n6627), .A4(n6626), .ZN(n9038)
         );
  NAND2_X1 U7834 ( .A1(n9385), .A2(n9038), .ZN(n8955) );
  OR2_X1 U7835 ( .A1(n9385), .A2(n9038), .ZN(n6630) );
  NAND2_X1 U7836 ( .A1(n9371), .A2(n9370), .ZN(n6631) );
  NAND2_X1 U7837 ( .A1(n6631), .A2(n8955), .ZN(n9356) );
  NAND2_X1 U7838 ( .A1(n7408), .A2(n8838), .ZN(n6636) );
  INV_X1 U7839 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6632) );
  NAND2_X1 U7840 ( .A1(n6633), .A2(n6632), .ZN(n6634) );
  NAND2_X1 U7841 ( .A1(n6634), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6644) );
  XNOR2_X1 U7842 ( .A(n6644), .B(P2_IR_REG_15__SCAN_IN), .ZN(n9103) );
  AOI22_X1 U7843 ( .A1(n8837), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6683), .B2(
        n9103), .ZN(n6635) );
  NAND2_X1 U7844 ( .A1(n7811), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6641) );
  NAND2_X1 U7845 ( .A1(n6839), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6640) );
  NAND2_X1 U7846 ( .A1(n7810), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6639) );
  AOI21_X1 U7847 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(n6637), .A(n6648), .ZN(
        n9362) );
  INV_X1 U7848 ( .A(n9362), .ZN(n8832) );
  NAND2_X1 U7849 ( .A1(n6728), .A2(n8832), .ZN(n6638) );
  OR2_X1 U7850 ( .A1(n9448), .A2(n9375), .ZN(n8958) );
  NAND2_X1 U7851 ( .A1(n9448), .A2(n9375), .ZN(n8957) );
  NAND2_X1 U7852 ( .A1(n8958), .A2(n8957), .ZN(n9357) );
  INV_X1 U7853 ( .A(n9375), .ZN(n9340) );
  NAND2_X1 U7854 ( .A1(n9448), .A2(n9340), .ZN(n6642) );
  NAND2_X1 U7855 ( .A1(n7607), .A2(n8838), .ZN(n6647) );
  INV_X1 U7856 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6643) );
  NAND2_X1 U7857 ( .A1(n6644), .A2(n6643), .ZN(n6645) );
  NAND2_X1 U7858 ( .A1(n6645), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6654) );
  XNOR2_X1 U7859 ( .A(n6654), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8554) );
  AOI22_X1 U7860 ( .A1(n8837), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6683), .B2(
        n8554), .ZN(n6646) );
  NAND2_X1 U7861 ( .A1(n7811), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6652) );
  NAND2_X1 U7862 ( .A1(n6839), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6651) );
  NAND2_X1 U7863 ( .A1(n7810), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6650) );
  OAI21_X1 U7864 ( .B1(n10658), .B2(n6648), .A(n6659), .ZN(n9343) );
  NAND2_X1 U7865 ( .A1(n6728), .A2(n9343), .ZN(n6649) );
  NAND2_X1 U7866 ( .A1(n9441), .A2(n9359), .ZN(n8961) );
  NAND2_X1 U7867 ( .A1(n9308), .A2(n8961), .ZN(n9346) );
  INV_X1 U7868 ( .A(n9359), .ZN(n9325) );
  NAND2_X1 U7869 ( .A1(n7739), .A2(n8838), .ZN(n6658) );
  INV_X1 U7870 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6653) );
  NAND2_X1 U7871 ( .A1(n6654), .A2(n6653), .ZN(n6655) );
  NAND2_X1 U7872 ( .A1(n6655), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6656) );
  XNOR2_X1 U7873 ( .A(n6656), .B(P2_IR_REG_17__SCAN_IN), .ZN(n9138) );
  AOI22_X1 U7874 ( .A1(n8837), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6683), .B2(
        n9138), .ZN(n6657) );
  NAND2_X1 U7875 ( .A1(n7810), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6664) );
  NAND2_X1 U7876 ( .A1(n7811), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6663) );
  NAND2_X1 U7877 ( .A1(n6659), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6660) );
  INV_X1 U7878 ( .A(n6675), .ZN(n6674) );
  NAND2_X1 U7879 ( .A1(n6660), .A2(n6674), .ZN(n9327) );
  NAND2_X1 U7880 ( .A1(n6728), .A2(n9327), .ZN(n6662) );
  NAND2_X1 U7881 ( .A1(n6839), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6661) );
  XNOR2_X1 U7882 ( .A(n9437), .B(n8966), .ZN(n6823) );
  INV_X1 U7883 ( .A(n9437), .ZN(n8968) );
  NAND2_X1 U7884 ( .A1(n7793), .A2(n8838), .ZN(n6673) );
  INV_X1 U7885 ( .A(n6666), .ZN(n6669) );
  INV_X1 U7886 ( .A(n6667), .ZN(n6668) );
  NOR2_X1 U7887 ( .A1(n6669), .A2(n6668), .ZN(n6670) );
  NAND2_X1 U7888 ( .A1(n6682), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6671) );
  XNOR2_X1 U7889 ( .A(n6671), .B(P2_IR_REG_18__SCAN_IN), .ZN(n9157) );
  AOI22_X1 U7890 ( .A1(n8837), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6683), .B2(
        n9157), .ZN(n6672) );
  NAND2_X1 U7891 ( .A1(n7810), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6680) );
  NAND2_X1 U7892 ( .A1(n7811), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6679) );
  NAND2_X1 U7893 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(n6674), .ZN(n6676) );
  INV_X1 U7894 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10752) );
  NAND2_X1 U7895 ( .A1(n10752), .A2(n6675), .ZN(n6686) );
  NAND2_X1 U7896 ( .A1(n6676), .A2(n6686), .ZN(n9313) );
  NAND2_X1 U7897 ( .A1(n6728), .A2(n9313), .ZN(n6678) );
  NAND2_X1 U7898 ( .A1(n6839), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6677) );
  NAND4_X1 U7899 ( .A1(n6680), .A2(n6679), .A3(n6678), .A4(n6677), .ZN(n9324)
         );
  INV_X1 U7900 ( .A(n9433), .ZN(n9318) );
  NAND2_X1 U7901 ( .A1(n9318), .A2(n8765), .ZN(n6681) );
  NAND2_X1 U7902 ( .A1(n7846), .A2(n8838), .ZN(n6685) );
  OAI21_X2 U7903 ( .B1(n6682), .B2(P2_IR_REG_18__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6802) );
  AOI22_X1 U7904 ( .A1(n8837), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9151), .B2(
        n6683), .ZN(n6684) );
  NAND2_X1 U7905 ( .A1(n7810), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6692) );
  NAND2_X1 U7906 ( .A1(n7811), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6691) );
  NAND2_X1 U7907 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(n6686), .ZN(n6688) );
  INV_X1 U7908 ( .A(n6686), .ZN(n6687) );
  INV_X1 U7909 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10729) );
  NAND2_X1 U7910 ( .A1(n6688), .A2(n6697), .ZN(n9299) );
  NAND2_X1 U7911 ( .A1(n6728), .A2(n9299), .ZN(n6690) );
  NAND2_X1 U7912 ( .A1(n6839), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6689) );
  NAND4_X1 U7913 ( .A1(n6692), .A2(n6691), .A3(n6690), .A4(n6689), .ZN(n9304)
         );
  NAND2_X1 U7914 ( .A1(n9298), .A2(n9304), .ZN(n6693) );
  NAND2_X1 U7915 ( .A1(n7845), .A2(n8838), .ZN(n6696) );
  OR2_X1 U7916 ( .A1(n8841), .A2(n6694), .ZN(n6695) );
  NAND2_X1 U7917 ( .A1(n7810), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6702) );
  NAND2_X1 U7918 ( .A1(n7811), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6701) );
  NAND2_X1 U7919 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(n6697), .ZN(n6698) );
  INV_X1 U7920 ( .A(n6708), .ZN(n6706) );
  NAND2_X1 U7921 ( .A1(n6698), .A2(n6706), .ZN(n9284) );
  NAND2_X1 U7922 ( .A1(n6728), .A2(n9284), .ZN(n6700) );
  NAND2_X1 U7923 ( .A1(n6839), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6699) );
  NAND4_X1 U7924 ( .A1(n6702), .A2(n6701), .A3(n6700), .A4(n6699), .ZN(n9292)
         );
  NAND2_X1 U7925 ( .A1(n9286), .A2(n9292), .ZN(n8975) );
  NAND2_X1 U7926 ( .A1(n9422), .A2(n8742), .ZN(n8974) );
  NAND2_X1 U7927 ( .A1(n9286), .A2(n8742), .ZN(n6703) );
  NAND2_X1 U7928 ( .A1(n7890), .A2(n8838), .ZN(n6705) );
  INV_X1 U7929 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7891) );
  OR2_X1 U7930 ( .A1(n8841), .A2(n7891), .ZN(n6704) );
  NAND2_X1 U7931 ( .A1(n7811), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6713) );
  NAND2_X1 U7932 ( .A1(n6839), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6712) );
  NAND2_X1 U7933 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(n6706), .ZN(n6709) );
  INV_X1 U7934 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n6707) );
  NAND2_X1 U7935 ( .A1(n6709), .A2(n6716), .ZN(n9272) );
  NAND2_X1 U7936 ( .A1(n6728), .A2(n9272), .ZN(n6711) );
  NAND2_X1 U7937 ( .A1(n7810), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6710) );
  NAND2_X1 U7938 ( .A1(n9418), .A2(n9257), .ZN(n8978) );
  NAND2_X1 U7939 ( .A1(n8979), .A2(n8978), .ZN(n9265) );
  NAND2_X1 U7940 ( .A1(n8059), .A2(n8838), .ZN(n6715) );
  OR2_X1 U7941 ( .A1(n8841), .A2(n8061), .ZN(n6714) );
  NAND2_X1 U7942 ( .A1(n7810), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6721) );
  NAND2_X1 U7943 ( .A1(n7811), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6720) );
  NAND2_X1 U7944 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(n6716), .ZN(n6717) );
  INV_X1 U7945 ( .A(n6724), .ZN(n6726) );
  NAND2_X1 U7946 ( .A1(n6717), .A2(n6726), .ZN(n9260) );
  NAND2_X1 U7947 ( .A1(n6728), .A2(n9260), .ZN(n6719) );
  NAND2_X1 U7948 ( .A1(n6839), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6718) );
  NAND4_X1 U7949 ( .A1(n6721), .A2(n6720), .A3(n6719), .A4(n6718), .ZN(n9266)
         );
  NAND2_X1 U7950 ( .A1(n8982), .A2(n9266), .ZN(n8846) );
  AND2_X1 U7951 ( .A1(n9265), .A2(n8846), .ZN(n9236) );
  NAND2_X1 U7952 ( .A1(n8117), .A2(n8838), .ZN(n6723) );
  OR2_X1 U7953 ( .A1(n8841), .A2(n8120), .ZN(n6722) );
  NAND2_X1 U7954 ( .A1(n7811), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6732) );
  NAND2_X1 U7955 ( .A1(n7810), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6731) );
  INV_X1 U7956 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n6725) );
  NAND2_X1 U7957 ( .A1(n6725), .A2(n6724), .ZN(n6744) );
  NAND2_X1 U7958 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(n6726), .ZN(n6727) );
  NAND2_X1 U7959 ( .A1(n6744), .A2(n6727), .ZN(n9246) );
  NAND2_X1 U7960 ( .A1(n6728), .A2(n9246), .ZN(n6730) );
  NAND2_X1 U7961 ( .A1(n6839), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6729) );
  NAND4_X1 U7962 ( .A1(n6732), .A2(n6731), .A3(n6730), .A4(n6729), .ZN(n8659)
         );
  NAND2_X1 U7963 ( .A1(n8663), .A2(n8659), .ZN(n6734) );
  AND2_X1 U7964 ( .A1(n9236), .A2(n6734), .ZN(n6733) );
  INV_X1 U7965 ( .A(n6734), .ZN(n6737) );
  INV_X1 U7966 ( .A(n8846), .ZN(n6736) );
  INV_X1 U7967 ( .A(n9418), .ZN(n8746) );
  NAND2_X1 U7968 ( .A1(n8746), .A2(n9257), .ZN(n9251) );
  OR2_X1 U7969 ( .A1(n8982), .A2(n9266), .ZN(n8847) );
  AND2_X1 U7970 ( .A1(n9251), .A2(n8847), .ZN(n6735) );
  OR2_X1 U7971 ( .A1(n6737), .A2(n9237), .ZN(n6739) );
  NAND2_X1 U7972 ( .A1(n9498), .A2(n9256), .ZN(n6738) );
  NAND2_X1 U7973 ( .A1(n8194), .A2(n8838), .ZN(n6741) );
  OR2_X1 U7974 ( .A1(n8841), .A2(n8195), .ZN(n6740) );
  NAND2_X1 U7975 ( .A1(n7811), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6749) );
  NAND2_X1 U7976 ( .A1(n6839), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6748) );
  INV_X1 U7977 ( .A(n6744), .ZN(n6743) );
  INV_X1 U7978 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n6742) );
  NAND2_X1 U7979 ( .A1(n6744), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6745) );
  NAND2_X1 U7980 ( .A1(n6754), .A2(n6745), .ZN(n9230) );
  NAND2_X1 U7981 ( .A1(n6728), .A2(n9230), .ZN(n6747) );
  NAND2_X1 U7982 ( .A1(n7810), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6746) );
  XNOR2_X1 U7983 ( .A(n8991), .B(n9242), .ZN(n9226) );
  NAND2_X1 U7984 ( .A1(n9494), .A2(n9242), .ZN(n6750) );
  NAND2_X1 U7985 ( .A1(n8228), .A2(n8838), .ZN(n6753) );
  OR2_X1 U7986 ( .A1(n8841), .A2(n8229), .ZN(n6752) );
  NAND2_X1 U7987 ( .A1(n7810), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6759) );
  NAND2_X1 U7988 ( .A1(n7811), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6758) );
  NAND2_X1 U7989 ( .A1(n6754), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6755) );
  NAND2_X1 U7990 ( .A1(n6765), .A2(n6755), .ZN(n9217) );
  NAND2_X1 U7991 ( .A1(n6728), .A2(n9217), .ZN(n6757) );
  NAND2_X1 U7992 ( .A1(n6839), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6756) );
  NAND2_X1 U7993 ( .A1(n8685), .A2(n9225), .ZN(n8996) );
  NAND2_X1 U7994 ( .A1(n8997), .A2(n8996), .ZN(n9214) );
  NAND2_X1 U7995 ( .A1(n9490), .A2(n9225), .ZN(n6760) );
  NAND2_X1 U7996 ( .A1(n8414), .A2(n8838), .ZN(n6762) );
  OR2_X1 U7997 ( .A1(n8841), .A2(n8416), .ZN(n6761) );
  NAND2_X1 U7998 ( .A1(n7811), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6770) );
  NAND2_X1 U7999 ( .A1(n6839), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6769) );
  INV_X1 U8000 ( .A(n6765), .ZN(n6764) );
  INV_X1 U8001 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n6763) );
  NAND2_X1 U8002 ( .A1(n6764), .A2(n6763), .ZN(n6775) );
  NAND2_X1 U8003 ( .A1(n6765), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6766) );
  NAND2_X1 U8004 ( .A1(n6775), .A2(n6766), .ZN(n9206) );
  NAND2_X1 U8005 ( .A1(n6728), .A2(n9206), .ZN(n6768) );
  NAND2_X1 U8006 ( .A1(n7810), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6767) );
  NAND4_X1 U8007 ( .A1(n6770), .A2(n6769), .A3(n6768), .A4(n6767), .ZN(n9035)
         );
  NAND2_X1 U8008 ( .A1(n6832), .A2(n9035), .ZN(n8691) );
  OR2_X1 U8009 ( .A1(n6832), .A2(n9035), .ZN(n8686) );
  NAND2_X1 U8010 ( .A1(n8380), .A2(n8838), .ZN(n6774) );
  OR2_X1 U8011 ( .A1(n8841), .A2(n6772), .ZN(n6773) );
  NAND2_X1 U8012 ( .A1(n7811), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6780) );
  NAND2_X1 U8013 ( .A1(n6839), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6779) );
  NAND2_X1 U8014 ( .A1(n6775), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6776) );
  NAND2_X1 U8015 ( .A1(n6788), .A2(n6776), .ZN(n9197) );
  NAND2_X1 U8016 ( .A1(n6728), .A2(n9197), .ZN(n6778) );
  NAND2_X1 U8017 ( .A1(n7810), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6777) );
  NAND4_X1 U8018 ( .A1(n6780), .A2(n6779), .A3(n6778), .A4(n6777), .ZN(n9034)
         );
  NAND2_X1 U8019 ( .A1(n9196), .A2(n9034), .ZN(n6782) );
  NOR2_X1 U8020 ( .A1(n9196), .A2(n9034), .ZN(n6781) );
  NAND2_X1 U8021 ( .A1(n8482), .A2(n8838), .ZN(n6785) );
  INV_X1 U8022 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n6783) );
  OR2_X1 U8023 ( .A1(n8841), .A2(n6783), .ZN(n6784) );
  NAND2_X1 U8024 ( .A1(n7811), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6793) );
  NAND2_X1 U8025 ( .A1(n7810), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6792) );
  INV_X1 U8026 ( .A(n6788), .ZN(n6787) );
  INV_X1 U8027 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6786) );
  NAND2_X1 U8028 ( .A1(n6787), .A2(n6786), .ZN(n8615) );
  NAND2_X1 U8029 ( .A1(n6788), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6789) );
  NAND2_X1 U8030 ( .A1(n8615), .A2(n6789), .ZN(n9184) );
  NAND2_X1 U8031 ( .A1(n6728), .A2(n9184), .ZN(n6791) );
  NAND2_X1 U8032 ( .A1(n6839), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6790) );
  NAND2_X1 U8033 ( .A1(n9478), .A2(n9189), .ZN(n6794) );
  INV_X1 U8034 ( .A(n9189), .ZN(n9033) );
  NAND2_X1 U8035 ( .A1(n8540), .A2(n8838), .ZN(n6796) );
  OR2_X1 U8036 ( .A1(n8841), .A2(n9514), .ZN(n6795) );
  INV_X1 U8037 ( .A(n8615), .ZN(n6797) );
  NAND2_X1 U8038 ( .A1(n6728), .A2(n6797), .ZN(n7815) );
  NAND2_X1 U8039 ( .A1(n7811), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6800) );
  NAND2_X1 U8040 ( .A1(n6839), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6799) );
  NAND2_X1 U8041 ( .A1(n7810), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6798) );
  NAND2_X1 U8042 ( .A1(n6893), .A2(n9179), .ZN(n9011) );
  NAND2_X1 U8043 ( .A1(n8875), .A2(n9011), .ZN(n6835) );
  NAND2_X1 U8044 ( .A1(n6802), .A2(n6801), .ZN(n6803) );
  NAND2_X1 U8045 ( .A1(n6807), .A2(n6804), .ZN(n6805) );
  NAND2_X1 U8046 ( .A1(n7476), .A2(n6897), .ZN(n7477) );
  NAND2_X1 U8047 ( .A1(n6808), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6809) );
  NAND2_X1 U8048 ( .A1(n9151), .A2(n9028), .ZN(n6874) );
  NAND2_X1 U8049 ( .A1(n6810), .A2(n9342), .ZN(n6845) );
  INV_X1 U8050 ( .A(n7593), .ZN(n6811) );
  NAND2_X1 U8051 ( .A1(n7542), .A2(n6811), .ZN(n7429) );
  NAND2_X1 U8052 ( .A1(n7430), .A2(n8886), .ZN(n7465) );
  INV_X1 U8053 ( .A(n8849), .ZN(n8892) );
  NAND2_X1 U8054 ( .A1(n7465), .A2(n8892), .ZN(n7464) );
  NAND2_X1 U8055 ( .A1(n7464), .A2(n8888), .ZN(n6813) );
  NAND2_X1 U8056 ( .A1(n7839), .A2(n6812), .ZN(n8889) );
  NAND2_X1 U8057 ( .A1(n9049), .A2(n7970), .ZN(n8900) );
  AND2_X1 U8058 ( .A1(n8889), .A2(n8900), .ZN(n7447) );
  NAND2_X1 U8059 ( .A1(n6813), .A2(n7447), .ZN(n7446) );
  NAND2_X1 U8060 ( .A1(n7446), .A2(n8889), .ZN(n7835) );
  NAND2_X1 U8061 ( .A1(n9047), .A2(n8012), .ZN(n8905) );
  NAND2_X1 U8062 ( .A1(n8150), .A2(n8130), .ZN(n8910) );
  NAND2_X1 U8063 ( .A1(n6520), .A2(n8160), .ZN(n8912) );
  NAND2_X1 U8064 ( .A1(n6814), .A2(n8853), .ZN(n8124) );
  NAND2_X1 U8065 ( .A1(n9046), .A2(n8931), .ZN(n8245) );
  AND2_X1 U8066 ( .A1(n8916), .A2(n8245), .ZN(n8921) );
  INV_X1 U8067 ( .A(n9042), .ZN(n8334) );
  NOR2_X1 U8068 ( .A1(n8479), .A2(n8334), .ZN(n8937) );
  INV_X1 U8069 ( .A(n8339), .ZN(n8344) );
  NAND2_X1 U8070 ( .A1(n8344), .A2(n8402), .ZN(n8925) );
  INV_X1 U8071 ( .A(n8925), .ZN(n6818) );
  NAND2_X1 U8072 ( .A1(n8942), .A2(n8372), .ZN(n6820) );
  OR2_X1 U8073 ( .A1(n8937), .A2(n6820), .ZN(n6819) );
  NAND2_X1 U8074 ( .A1(n8479), .A2(n8334), .ZN(n8924) );
  AND2_X1 U8075 ( .A1(n8924), .A2(n8925), .ZN(n8370) );
  OR2_X1 U8076 ( .A1(n6820), .A2(n8370), .ZN(n6821) );
  NAND2_X1 U8077 ( .A1(n8405), .A2(n8507), .ZN(n8927) );
  AND2_X1 U8078 ( .A1(n9462), .A2(n9374), .ZN(n8947) );
  NAND2_X1 U8079 ( .A1(n9369), .A2(n9368), .ZN(n9367) );
  OR2_X1 U8080 ( .A1(n9385), .A2(n9360), .ZN(n6822) );
  NAND2_X1 U8081 ( .A1(n9367), .A2(n6822), .ZN(n9355) );
  INV_X1 U8082 ( .A(n8957), .ZN(n9347) );
  NOR2_X1 U8083 ( .A1(n9346), .A2(n9347), .ZN(n9307) );
  NAND2_X1 U8084 ( .A1(n9433), .A2(n8765), .ZN(n8967) );
  AND2_X1 U8085 ( .A1(n9307), .A2(n6824), .ZN(n6825) );
  INV_X1 U8086 ( .A(n9311), .ZN(n6826) );
  OR2_X1 U8087 ( .A1(n9437), .A2(n8966), .ZN(n9309) );
  OR2_X1 U8088 ( .A1(n6826), .A2(n9309), .ZN(n6827) );
  INV_X1 U8089 ( .A(n9304), .ZN(n8971) );
  OR2_X1 U8090 ( .A1(n9298), .A2(n8971), .ZN(n6828) );
  INV_X1 U8091 ( .A(n9265), .ZN(n9268) );
  NAND2_X1 U8092 ( .A1(n9271), .A2(n8979), .ZN(n9258) );
  NAND2_X1 U8093 ( .A1(n8982), .A2(n9243), .ZN(n6829) );
  OR2_X1 U8094 ( .A1(n8982), .A2(n9243), .ZN(n6830) );
  AND2_X1 U8095 ( .A1(n9498), .A2(n8659), .ZN(n8986) );
  NAND2_X1 U8096 ( .A1(n8663), .A2(n9256), .ZN(n8987) );
  INV_X1 U8097 ( .A(n9242), .ZN(n9037) );
  NAND2_X1 U8098 ( .A1(n9494), .A2(n9037), .ZN(n8992) );
  INV_X1 U8099 ( .A(n8997), .ZN(n6831) );
  NAND2_X1 U8100 ( .A1(n9486), .A2(n9035), .ZN(n8999) );
  INV_X1 U8101 ( .A(n9035), .ZN(n9213) );
  NAND2_X1 U8102 ( .A1(n6832), .A2(n9213), .ZN(n9192) );
  NAND2_X1 U8103 ( .A1(n9196), .A2(n9204), .ZN(n9003) );
  NAND2_X1 U8104 ( .A1(n6833), .A2(n9004), .ZN(n9183) );
  NAND2_X1 U8105 ( .A1(n8698), .A2(n9189), .ZN(n8872) );
  INV_X1 U8106 ( .A(n6834), .ZN(n8873) );
  NAND2_X1 U8107 ( .A1(n6847), .A2(n5535), .ZN(n6895) );
  AOI21_X1 U8108 ( .B1(n6897), .B2(n8060), .A(n9151), .ZN(n6836) );
  XNOR2_X1 U8109 ( .A(n6837), .B(n8174), .ZN(n7518) );
  INV_X1 U8110 ( .A(n7518), .ZN(n7502) );
  NAND2_X1 U8111 ( .A1(n7810), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6842) );
  NAND2_X1 U8112 ( .A1(n7811), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6841) );
  NAND2_X1 U8113 ( .A1(n6839), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6840) );
  AND2_X1 U8114 ( .A1(n7130), .A2(P2_B_REG_SCAN_IN), .ZN(n6843) );
  OR2_X1 U8115 ( .A1(n9376), .A2(n6843), .ZN(n9170) );
  OAI22_X1 U8116 ( .A1(n9189), .A2(n9361), .B1(n8844), .B2(n9170), .ZN(n6844)
         );
  OR2_X1 U8117 ( .A1(n7515), .A2(n9028), .ZN(n8475) );
  NAND2_X1 U8118 ( .A1(n6848), .A2(n5143), .ZN(n6906) );
  NAND2_X1 U8119 ( .A1(n6849), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6850) );
  INV_X1 U8120 ( .A(n6851), .ZN(n6852) );
  NAND2_X1 U8121 ( .A1(n6852), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6853) );
  MUX2_X1 U8122 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6853), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n6854) );
  NAND2_X1 U8123 ( .A1(n6854), .A2(n5151), .ZN(n8196) );
  XNOR2_X1 U8124 ( .A(n8196), .B(P2_B_REG_SCAN_IN), .ZN(n6857) );
  NAND2_X1 U8125 ( .A1(n5151), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6856) );
  XNOR2_X1 U8126 ( .A(n6856), .B(n6855), .ZN(n8230) );
  NAND2_X1 U8127 ( .A1(n6857), .A2(n8230), .ZN(n6858) );
  INV_X1 U8128 ( .A(n7144), .ZN(n6859) );
  INV_X1 U8129 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n7151) );
  NAND2_X1 U8130 ( .A1(n6859), .A2(n7151), .ZN(n6860) );
  INV_X1 U8131 ( .A(n6885), .ZN(n8415) );
  NAND2_X1 U8132 ( .A1(n8415), .A2(n8230), .ZN(n7148) );
  NAND2_X1 U8133 ( .A1(n6860), .A2(n7148), .ZN(n6899) );
  INV_X1 U8134 ( .A(n6899), .ZN(n7586) );
  NAND2_X1 U8135 ( .A1(n8415), .A2(n8196), .ZN(n7145) );
  NAND2_X1 U8136 ( .A1(n7586), .A2(n7582), .ZN(n6904) );
  NOR2_X1 U8137 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6865) );
  NOR4_X1 U8138 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6864) );
  NOR4_X1 U8139 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6863) );
  NOR4_X1 U8140 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6862) );
  NAND4_X1 U8141 ( .A1(n6865), .A2(n6864), .A3(n6863), .A4(n6862), .ZN(n6871)
         );
  NOR4_X1 U8142 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6869) );
  NOR4_X1 U8143 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6868) );
  NOR4_X1 U8144 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6867) );
  NOR4_X1 U8145 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6866) );
  NAND4_X1 U8146 ( .A1(n6869), .A2(n6868), .A3(n6867), .A4(n6866), .ZN(n6870)
         );
  NOR2_X1 U8147 ( .A1(n6871), .A2(n6870), .ZN(n6872) );
  INV_X1 U8148 ( .A(n6902), .ZN(n6873) );
  INV_X1 U8149 ( .A(n6874), .ZN(n6875) );
  NAND2_X1 U8150 ( .A1(n6875), .A2(n6897), .ZN(n6876) );
  OR2_X1 U8151 ( .A1(n7476), .A2(n6876), .ZN(n7496) );
  NAND2_X1 U8152 ( .A1(n7500), .A2(n7496), .ZN(n6877) );
  NAND2_X1 U8153 ( .A1(n7514), .A2(n6877), .ZN(n6881) );
  NAND2_X1 U8154 ( .A1(n6899), .A2(n6902), .ZN(n6878) );
  NOR2_X1 U8155 ( .A1(n6878), .A2(n7582), .ZN(n7510) );
  NAND3_X1 U8156 ( .A1(n9007), .A2(n7496), .A3(n9450), .ZN(n6879) );
  INV_X1 U8157 ( .A(n7515), .ZN(n7796) );
  OR2_X1 U8158 ( .A1(n9450), .A2(n7796), .ZN(n8509) );
  NAND2_X1 U8159 ( .A1(n6879), .A2(n8509), .ZN(n7504) );
  NAND2_X1 U8160 ( .A1(n7510), .A2(n7504), .ZN(n6880) );
  NAND2_X1 U8161 ( .A1(n6881), .A2(n6880), .ZN(n9467) );
  INV_X1 U8162 ( .A(n8230), .ZN(n6883) );
  INV_X1 U8163 ( .A(n8196), .ZN(n6882) );
  INV_X1 U8164 ( .A(n6886), .ZN(n6887) );
  NAND2_X1 U8165 ( .A1(n6887), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6889) );
  XNOR2_X1 U8166 ( .A(n6889), .B(n6888), .ZN(n8118) );
  OR2_X1 U8167 ( .A1(n6906), .A2(n6890), .ZN(n6892) );
  OR2_X1 U8168 ( .A1(n11121), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6891) );
  NAND2_X1 U8169 ( .A1(n6892), .A2(n6891), .ZN(n6894) );
  NAND2_X1 U8170 ( .A1(n11121), .A2(n9463), .ZN(n9508) );
  NAND2_X1 U8171 ( .A1(n6894), .A2(n5746), .ZN(P2_U3456) );
  OAI21_X1 U8172 ( .B1(n7476), .B2(n8475), .A(n7582), .ZN(n6901) );
  INV_X1 U8173 ( .A(n6895), .ZN(n6896) );
  NAND3_X1 U8174 ( .A1(n6897), .A2(n9028), .A3(n5535), .ZN(n6898) );
  NAND2_X1 U8175 ( .A1(n9007), .A2(n6898), .ZN(n7585) );
  NAND2_X1 U8176 ( .A1(n7583), .A2(n7585), .ZN(n6900) );
  AOI22_X1 U8177 ( .A1(n6901), .A2(n6900), .B1(n6899), .B2(n7585), .ZN(n6905)
         );
  AND2_X1 U8178 ( .A1(n6902), .A2(n7513), .ZN(n6903) );
  OR2_X1 U8179 ( .A1(n6906), .A2(n9465), .ZN(n6908) );
  NAND2_X1 U8180 ( .A1(n6908), .A2(n6907), .ZN(n6909) );
  NAND2_X1 U8181 ( .A1(n6909), .A2(n5745), .ZN(P2_U3488) );
  INV_X1 U8182 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6911) );
  NOR2_X1 U8183 ( .A1(n11110), .A2(n6911), .ZN(n6912) );
  OAI21_X1 U8184 ( .B1(n6914), .B2(n11109), .A(n6913), .ZN(P1_U3551) );
  INV_X1 U8185 ( .A(n6917), .ZN(n6915) );
  AND2_X4 U8186 ( .A1(n6915), .A2(n7126), .ZN(n7089) );
  OR2_X2 U8187 ( .A1(n6917), .A2(n5130), .ZN(n7743) );
  NAND2_X1 U8188 ( .A1(n6918), .A2(n9758), .ZN(n6919) );
  NAND3_X4 U8189 ( .A1(n7743), .A2(n7126), .A3(n6919), .ZN(n8704) );
  OAI22_X1 U8190 ( .A1(n10305), .A2(n5129), .B1(n6140), .B2(n8704), .ZN(n9666)
         );
  AOI22_X1 U8191 ( .A1(n7716), .A2(n7089), .B1(n9999), .B2(n7097), .ZN(n6961)
         );
  INV_X1 U8192 ( .A(n6961), .ZN(n8134) );
  OAI22_X1 U8193 ( .A1(n7940), .A2(n8704), .B1(n6009), .B2(n5129), .ZN(n6950)
         );
  INV_X2 U8194 ( .A(n6943), .ZN(n6922) );
  INV_X4 U8195 ( .A(n6922), .ZN(n8703) );
  AOI22_X1 U8196 ( .A1(n10002), .A2(n7089), .B1(n6943), .B2(n7923), .ZN(n6923)
         );
  XNOR2_X1 U8197 ( .A(n6923), .B(n8706), .ZN(n6948) );
  INV_X1 U8198 ( .A(n6948), .ZN(n6949) );
  INV_X1 U8199 ( .A(n7126), .ZN(n7170) );
  NAND2_X1 U8200 ( .A1(n7170), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6925) );
  NAND2_X1 U8201 ( .A1(n6929), .A2(n6925), .ZN(n7303) );
  OR2_X1 U8202 ( .A1(n8704), .A2(n7569), .ZN(n6927) );
  AOI22_X1 U8203 ( .A1(n7089), .A2(n11024), .B1(n7170), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n6926) );
  NAND2_X1 U8204 ( .A1(n6927), .A2(n6926), .ZN(n7301) );
  NAND2_X1 U8205 ( .A1(n7303), .A2(n7301), .ZN(n7302) );
  NAND2_X1 U8206 ( .A1(n6929), .A2(n7086), .ZN(n6930) );
  NAND2_X1 U8207 ( .A1(n6943), .A2(n6934), .ZN(n6932) );
  NAND2_X1 U8208 ( .A1(n6332), .A2(n7089), .ZN(n6931) );
  NAND2_X1 U8209 ( .A1(n6932), .A2(n6931), .ZN(n6933) );
  NAND2_X1 U8210 ( .A1(n6935), .A2(n6936), .ZN(n7400) );
  AOI22_X1 U8211 ( .A1(n7097), .A2(n6332), .B1(n7089), .B2(n6934), .ZN(n7399)
         );
  NAND2_X1 U8212 ( .A1(n7400), .A2(n7399), .ZN(n7398) );
  NAND2_X1 U8213 ( .A1(n6938), .A2(n6937), .ZN(n7402) );
  AOI22_X1 U8214 ( .A1(n10004), .A2(n7089), .B1(n6943), .B2(n7694), .ZN(n6939)
         );
  XNOR2_X1 U8215 ( .A(n6939), .B(n8706), .ZN(n6942) );
  OAI22_X1 U8216 ( .A1(n7568), .A2(n8704), .B1(n8074), .B2(n5129), .ZN(n6940)
         );
  XNOR2_X1 U8217 ( .A(n6942), .B(n6940), .ZN(n7437) );
  INV_X1 U8218 ( .A(n6940), .ZN(n6941) );
  OAI22_X1 U8219 ( .A1(n7439), .A2(n8704), .B1(n11044), .B2(n5129), .ZN(n6946)
         );
  AOI22_X1 U8220 ( .A1(n10003), .A2(n7089), .B1(n6943), .B2(n5994), .ZN(n6944)
         );
  XNOR2_X1 U8221 ( .A(n6944), .B(n8706), .ZN(n6945) );
  XOR2_X1 U8222 ( .A(n6946), .B(n6945), .Z(n7458) );
  INV_X1 U8223 ( .A(n6945), .ZN(n6947) );
  AOI22_X1 U8224 ( .A1(n10001), .A2(n7089), .B1(n8703), .B2(n7946), .ZN(n6951)
         );
  XNOR2_X1 U8225 ( .A(n6951), .B(n8706), .ZN(n6952) );
  OAI22_X1 U8226 ( .A1(n6922), .A2(n11073), .B1(n8141), .B2(n5129), .ZN(n6953)
         );
  XNOR2_X1 U8227 ( .A(n6953), .B(n7086), .ZN(n6957) );
  OR2_X1 U8228 ( .A1(n11073), .A2(n5129), .ZN(n6955) );
  NAND2_X1 U8229 ( .A1(n7097), .A2(n10000), .ZN(n6954) );
  AND2_X1 U8230 ( .A1(n6955), .A2(n6954), .ZN(n6956) );
  NAND2_X1 U8231 ( .A1(n6957), .A2(n6956), .ZN(n8019) );
  INV_X1 U8232 ( .A(n8019), .ZN(n6958) );
  AOI22_X1 U8233 ( .A1(n7716), .A2(n8703), .B1(n9999), .B2(n7089), .ZN(n6960)
         );
  XNOR2_X1 U8234 ( .A(n6960), .B(n8706), .ZN(n8135) );
  NAND2_X1 U8235 ( .A1(n8239), .A2(n8703), .ZN(n6963) );
  OR2_X1 U8236 ( .A1(n7962), .A2(n5129), .ZN(n6962) );
  NAND2_X1 U8237 ( .A1(n6963), .A2(n6962), .ZN(n6964) );
  XNOR2_X1 U8238 ( .A(n6964), .B(n8706), .ZN(n6966) );
  OAI22_X1 U8239 ( .A1(n8083), .A2(n5129), .B1(n7962), .B2(n8704), .ZN(n6965)
         );
  XNOR2_X1 U8240 ( .A(n6966), .B(n6965), .ZN(n8231) );
  INV_X1 U8241 ( .A(n6965), .ZN(n6968) );
  INV_X1 U8242 ( .A(n6966), .ZN(n6967) );
  NAND2_X1 U8243 ( .A1(n8299), .A2(n8703), .ZN(n6970) );
  OR2_X1 U8244 ( .A1(n9545), .A2(n5129), .ZN(n6969) );
  NAND2_X1 U8245 ( .A1(n6970), .A2(n6969), .ZN(n6971) );
  XNOR2_X1 U8246 ( .A(n6971), .B(n8706), .ZN(n6974) );
  AOI22_X1 U8247 ( .A1(n8299), .A2(n7089), .B1(n7097), .B2(n9997), .ZN(n6972)
         );
  XNOR2_X1 U8248 ( .A(n6974), .B(n6972), .ZN(n8294) );
  INV_X1 U8249 ( .A(n6972), .ZN(n6973) );
  OAI22_X1 U8250 ( .A1(n5700), .A2(n5129), .B1(n9654), .B2(n8704), .ZN(n9538)
         );
  INV_X1 U8251 ( .A(n9538), .ZN(n6978) );
  AOI22_X1 U8252 ( .A1(n9547), .A2(n8703), .B1(n7089), .B2(n11090), .ZN(n6976)
         );
  XOR2_X1 U8253 ( .A(n8706), .B(n6976), .Z(n9539) );
  INV_X1 U8254 ( .A(n9539), .ZN(n6977) );
  AOI21_X1 U8255 ( .B1(n9541), .B2(n6978), .A(n6977), .ZN(n6979) );
  NAND2_X1 U8256 ( .A1(n9663), .A2(n8703), .ZN(n6981) );
  NAND2_X1 U8257 ( .A1(n9996), .A2(n7089), .ZN(n6980) );
  NAND2_X1 U8258 ( .A1(n6981), .A2(n6980), .ZN(n6982) );
  XNOR2_X1 U8259 ( .A(n6982), .B(n7086), .ZN(n6988) );
  AND2_X1 U8260 ( .A1(n7097), .A2(n9996), .ZN(n6983) );
  AOI21_X1 U8261 ( .B1(n9663), .B2(n7089), .A(n6983), .ZN(n6989) );
  NAND2_X1 U8262 ( .A1(n6988), .A2(n6989), .ZN(n9657) );
  NAND2_X1 U8263 ( .A1(n8108), .A2(n8703), .ZN(n6985) );
  NAND2_X1 U8264 ( .A1(n11087), .A2(n7089), .ZN(n6984) );
  NAND2_X1 U8265 ( .A1(n6985), .A2(n6984), .ZN(n6986) );
  XNOR2_X1 U8266 ( .A(n6986), .B(n8706), .ZN(n6997) );
  AND2_X1 U8267 ( .A1(n7097), .A2(n11087), .ZN(n6987) );
  AOI21_X1 U8268 ( .B1(n8108), .B2(n7089), .A(n6987), .ZN(n6998) );
  XNOR2_X1 U8269 ( .A(n6997), .B(n6998), .ZN(n9568) );
  INV_X1 U8270 ( .A(n6988), .ZN(n6991) );
  INV_X1 U8271 ( .A(n6989), .ZN(n6990) );
  NAND2_X1 U8272 ( .A1(n6991), .A2(n6990), .ZN(n9659) );
  NAND2_X1 U8273 ( .A1(n8207), .A2(n8703), .ZN(n6994) );
  NAND2_X1 U8274 ( .A1(n10415), .A2(n7089), .ZN(n6993) );
  NAND2_X1 U8275 ( .A1(n6994), .A2(n6993), .ZN(n6995) );
  XNOR2_X1 U8276 ( .A(n6995), .B(n8706), .ZN(n7000) );
  AND2_X1 U8277 ( .A1(n7097), .A2(n10415), .ZN(n6996) );
  AOI21_X1 U8278 ( .B1(n8207), .B2(n7089), .A(n6996), .ZN(n7001) );
  XNOR2_X1 U8279 ( .A(n7000), .B(n7001), .ZN(n9629) );
  INV_X1 U8280 ( .A(n6997), .ZN(n6999) );
  NAND2_X1 U8281 ( .A1(n6999), .A2(n6998), .ZN(n9627) );
  NAND3_X1 U8282 ( .A1(n9567), .A2(n9629), .A3(n9627), .ZN(n9628) );
  NAND2_X1 U8283 ( .A1(n9527), .A2(n8703), .ZN(n7005) );
  OR2_X1 U8284 ( .A1(n9692), .A2(n5129), .ZN(n7004) );
  NAND2_X1 U8285 ( .A1(n7005), .A2(n7004), .ZN(n7006) );
  XNOR2_X1 U8286 ( .A(n7006), .B(n7086), .ZN(n9520) );
  NOR2_X1 U8287 ( .A1(n9692), .A2(n8704), .ZN(n7007) );
  AOI21_X1 U8288 ( .B1(n9527), .B2(n7089), .A(n7007), .ZN(n7008) );
  NAND2_X1 U8289 ( .A1(n9520), .A2(n7008), .ZN(n7010) );
  INV_X1 U8290 ( .A(n9520), .ZN(n7009) );
  INV_X1 U8291 ( .A(n7008), .ZN(n9519) );
  AOI21_X2 U8292 ( .B1(n9522), .B2(n7010), .A(n5155), .ZN(n9686) );
  NAND2_X1 U8293 ( .A1(n10398), .A2(n8703), .ZN(n7012) );
  OR2_X1 U8294 ( .A1(n10389), .A2(n5129), .ZN(n7011) );
  NAND2_X1 U8295 ( .A1(n7012), .A2(n7011), .ZN(n7013) );
  XNOR2_X1 U8296 ( .A(n7013), .B(n7086), .ZN(n7022) );
  NOR2_X1 U8297 ( .A1(n10389), .A2(n8704), .ZN(n7014) );
  AOI21_X1 U8298 ( .B1(n10398), .B2(n7089), .A(n7014), .ZN(n7021) );
  OR2_X1 U8299 ( .A1(n7022), .A2(n7021), .ZN(n9585) );
  NAND2_X1 U8300 ( .A1(n9695), .A2(n8703), .ZN(n7016) );
  OR2_X1 U8301 ( .A1(n9523), .A2(n5129), .ZN(n7015) );
  NAND2_X1 U8302 ( .A1(n7016), .A2(n7015), .ZN(n7017) );
  XNOR2_X1 U8303 ( .A(n7017), .B(n7086), .ZN(n9684) );
  NOR2_X1 U8304 ( .A1(n9523), .A2(n8704), .ZN(n7018) );
  AOI21_X1 U8305 ( .B1(n9695), .B2(n7089), .A(n7018), .ZN(n9683) );
  OR2_X1 U8306 ( .A1(n9684), .A2(n9683), .ZN(n7019) );
  AND2_X1 U8307 ( .A1(n9585), .A2(n7019), .ZN(n7020) );
  NAND2_X1 U8308 ( .A1(n9686), .A2(n7020), .ZN(n7027) );
  INV_X1 U8309 ( .A(n9585), .ZN(n7024) );
  NAND2_X1 U8310 ( .A1(n9684), .A2(n9683), .ZN(n7023) );
  NAND2_X1 U8311 ( .A1(n7022), .A2(n7021), .ZN(n9597) );
  INV_X1 U8312 ( .A(n7025), .ZN(n7026) );
  NAND2_X1 U8313 ( .A1(n7027), .A2(n7026), .ZN(n7035) );
  NAND2_X1 U8314 ( .A1(n8530), .A2(n8703), .ZN(n7029) );
  OR2_X1 U8315 ( .A1(n10297), .A2(n5129), .ZN(n7028) );
  NAND2_X1 U8316 ( .A1(n7029), .A2(n7028), .ZN(n7030) );
  XNOR2_X1 U8317 ( .A(n7030), .B(n7086), .ZN(n7033) );
  NOR2_X1 U8318 ( .A1(n10297), .A2(n8704), .ZN(n7031) );
  AOI21_X1 U8319 ( .B1(n8530), .B2(n7089), .A(n7031), .ZN(n7032) );
  NAND2_X1 U8320 ( .A1(n7033), .A2(n7032), .ZN(n7036) );
  OR2_X1 U8321 ( .A1(n7033), .A2(n7032), .ZN(n7034) );
  AND2_X1 U8322 ( .A1(n7036), .A2(n7034), .ZN(n9598) );
  AOI22_X1 U8323 ( .A1(n10385), .A2(n8703), .B1(n7089), .B2(n10282), .ZN(n7037) );
  XNOR2_X1 U8324 ( .A(n7037), .B(n8706), .ZN(n7038) );
  NAND2_X1 U8325 ( .A1(n10379), .A2(n8703), .ZN(n7040) );
  NAND2_X1 U8326 ( .A1(n10265), .A2(n7089), .ZN(n7039) );
  NAND2_X1 U8327 ( .A1(n7040), .A2(n7039), .ZN(n7041) );
  XNOR2_X1 U8328 ( .A(n7041), .B(n8706), .ZN(n7045) );
  NAND2_X1 U8329 ( .A1(n10379), .A2(n7089), .ZN(n7043) );
  NAND2_X1 U8330 ( .A1(n7097), .A2(n10265), .ZN(n7042) );
  NAND2_X1 U8331 ( .A1(n7043), .A2(n7042), .ZN(n7044) );
  NOR2_X1 U8332 ( .A1(n7045), .A2(n7044), .ZN(n7046) );
  AOI21_X1 U8333 ( .B1(n7045), .B2(n7044), .A(n7046), .ZN(n9552) );
  INV_X1 U8334 ( .A(n7046), .ZN(n7047) );
  NAND2_X1 U8335 ( .A1(n9550), .A2(n7047), .ZN(n9620) );
  AOI22_X1 U8336 ( .A1(n10263), .A2(n8703), .B1(n7089), .B2(n9562), .ZN(n7048)
         );
  XNOR2_X1 U8337 ( .A(n7048), .B(n8706), .ZN(n7053) );
  OAI22_X1 U8338 ( .A1(n10368), .A2(n5129), .B1(n10376), .B2(n8704), .ZN(n7054) );
  XNOR2_X1 U8339 ( .A(n7053), .B(n7054), .ZN(n9621) );
  NAND2_X1 U8340 ( .A1(n10253), .A2(n8703), .ZN(n7050) );
  OR2_X1 U8341 ( .A1(n10273), .A2(n5129), .ZN(n7049) );
  NAND2_X1 U8342 ( .A1(n7050), .A2(n7049), .ZN(n7051) );
  XNOR2_X1 U8343 ( .A(n7051), .B(n8706), .ZN(n7058) );
  NOR2_X1 U8344 ( .A1(n10273), .A2(n8704), .ZN(n7052) );
  AOI21_X1 U8345 ( .B1(n10253), .B2(n7089), .A(n7052), .ZN(n7056) );
  XNOR2_X1 U8346 ( .A(n7058), .B(n7056), .ZN(n9558) );
  INV_X1 U8347 ( .A(n7053), .ZN(n7055) );
  OR2_X1 U8348 ( .A1(n7055), .A2(n7054), .ZN(n9559) );
  INV_X1 U8349 ( .A(n7056), .ZN(n7057) );
  OAI22_X1 U8350 ( .A1(n10453), .A2(n6922), .B1(n10248), .B2(n5129), .ZN(n7060) );
  XOR2_X1 U8351 ( .A(n8706), .B(n7060), .Z(n7071) );
  NAND2_X1 U8352 ( .A1(n7070), .A2(n7071), .ZN(n9639) );
  OAI22_X1 U8353 ( .A1(n10453), .A2(n5129), .B1(n10248), .B2(n8704), .ZN(n9641) );
  NAND2_X1 U8354 ( .A1(n9639), .A2(n9641), .ZN(n9532) );
  NAND2_X1 U8355 ( .A1(n10222), .A2(n8703), .ZN(n7062) );
  NAND2_X1 U8356 ( .A1(n10230), .A2(n7089), .ZN(n7061) );
  NAND2_X1 U8357 ( .A1(n7062), .A2(n7061), .ZN(n7063) );
  XNOR2_X1 U8358 ( .A(n7063), .B(n7086), .ZN(n7065) );
  AND2_X1 U8359 ( .A1(n7097), .A2(n10230), .ZN(n7064) );
  AOI21_X1 U8360 ( .B1(n10222), .B2(n7089), .A(n7064), .ZN(n7066) );
  NAND2_X1 U8361 ( .A1(n7065), .A2(n7066), .ZN(n7074) );
  INV_X1 U8362 ( .A(n7065), .ZN(n7068) );
  INV_X1 U8363 ( .A(n7066), .ZN(n7067) );
  NAND2_X1 U8364 ( .A1(n7068), .A2(n7067), .ZN(n7069) );
  AND2_X1 U8365 ( .A1(n7074), .A2(n7069), .ZN(n9531) );
  INV_X1 U8366 ( .A(n7070), .ZN(n7073) );
  INV_X1 U8367 ( .A(n7071), .ZN(n7072) );
  NAND2_X1 U8368 ( .A1(n7073), .A2(n7072), .ZN(n9638) );
  AND3_X2 U8369 ( .A1(n9532), .A2(n9531), .A3(n9638), .ZN(n9530) );
  INV_X1 U8370 ( .A(n7074), .ZN(n9611) );
  OAI22_X1 U8371 ( .A1(n10445), .A2(n6922), .B1(n10217), .B2(n5129), .ZN(n7075) );
  XNOR2_X1 U8372 ( .A(n7075), .B(n8706), .ZN(n7077) );
  OAI22_X1 U8373 ( .A1(n10445), .A2(n5129), .B1(n10217), .B2(n8704), .ZN(n7076) );
  NAND2_X1 U8374 ( .A1(n7077), .A2(n7076), .ZN(n7078) );
  OAI22_X1 U8375 ( .A1(n10441), .A2(n5129), .B1(n7080), .B2(n8704), .ZN(n7090)
         );
  NAND2_X1 U8376 ( .A1(n10192), .A2(n8703), .ZN(n7082) );
  NAND2_X1 U8377 ( .A1(n10325), .A2(n7089), .ZN(n7081) );
  NAND2_X1 U8378 ( .A1(n7082), .A2(n7081), .ZN(n7083) );
  XNOR2_X1 U8379 ( .A(n7083), .B(n8706), .ZN(n7091) );
  XOR2_X1 U8380 ( .A(n7090), .B(n7091), .Z(n9579) );
  NAND2_X1 U8381 ( .A1(n10178), .A2(n8703), .ZN(n7085) );
  OR2_X1 U8382 ( .A1(n10317), .A2(n5129), .ZN(n7084) );
  NAND2_X1 U8383 ( .A1(n7085), .A2(n7084), .ZN(n7087) );
  XNOR2_X1 U8384 ( .A(n7087), .B(n7086), .ZN(n7092) );
  NOR2_X1 U8385 ( .A1(n10317), .A2(n8704), .ZN(n7088) );
  AOI21_X1 U8386 ( .B1(n10178), .B2(n7089), .A(n7088), .ZN(n7093) );
  XNOR2_X1 U8387 ( .A(n7092), .B(n7093), .ZN(n9672) );
  NOR2_X1 U8388 ( .A1(n7091), .A2(n7090), .ZN(n9673) );
  INV_X1 U8389 ( .A(n9675), .ZN(n7100) );
  INV_X1 U8390 ( .A(n7092), .ZN(n7095) );
  INV_X1 U8391 ( .A(n7093), .ZN(n7094) );
  AND2_X1 U8392 ( .A1(n7095), .A2(n7094), .ZN(n7101) );
  AOI22_X1 U8393 ( .A1(n10157), .A2(n8703), .B1(n7089), .B2(n10326), .ZN(n7096) );
  XNOR2_X1 U8394 ( .A(n7096), .B(n8706), .ZN(n7099) );
  AOI22_X1 U8395 ( .A1(n10157), .A2(n7089), .B1(n7097), .B2(n10326), .ZN(n7098) );
  NAND2_X1 U8396 ( .A1(n7099), .A2(n7098), .ZN(n8701) );
  OAI21_X1 U8397 ( .B1(n7099), .B2(n7098), .A(n8701), .ZN(n7102) );
  OAI21_X2 U8398 ( .B1(n7100), .B2(n7101), .A(n7102), .ZN(n7108) );
  NOR2_X1 U8399 ( .A1(n7102), .A2(n7101), .ZN(n7103) );
  INV_X1 U8400 ( .A(n7104), .ZN(n7106) );
  NOR2_X1 U8401 ( .A1(n7106), .A2(n7105), .ZN(n7552) );
  INV_X1 U8402 ( .A(n7107), .ZN(n10469) );
  NAND2_X1 U8403 ( .A1(n7552), .A2(n10469), .ZN(n7116) );
  INV_X1 U8404 ( .A(n10468), .ZN(n9701) );
  NAND2_X1 U8405 ( .A1(n11103), .A2(n9808), .ZN(n7113) );
  AOI21_X1 U8406 ( .B1(n7108), .B2(n8702), .A(n9697), .ZN(n7109) );
  INV_X1 U8407 ( .A(n7109), .ZN(n7125) );
  OR2_X1 U8408 ( .A1(n7601), .A2(n7848), .ZN(n7554) );
  OR3_X1 U8409 ( .A1(n7116), .A2(n9701), .A3(n7554), .ZN(n7112) );
  INV_X1 U8410 ( .A(n7110), .ZN(n7111) );
  INV_X1 U8411 ( .A(n9700), .ZN(n7602) );
  NAND2_X1 U8412 ( .A1(n7602), .A2(n10468), .ZN(n7114) );
  AOI22_X1 U8413 ( .A1(n9678), .A2(n10334), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n7122) );
  NAND3_X1 U8414 ( .A1(n7114), .A2(n7554), .A3(n7113), .ZN(n7115) );
  NAND2_X1 U8415 ( .A1(n7116), .A2(n7115), .ZN(n7305) );
  AND3_X1 U8416 ( .A1(n7117), .A2(n8114), .A3(n7126), .ZN(n7118) );
  NAND2_X1 U8417 ( .A1(n7305), .A2(n7118), .ZN(n7119) );
  AOI22_X1 U8418 ( .A1(n9689), .A2(n10158), .B1(n9687), .B2(n9995), .ZN(n7121)
         );
  OAI211_X1 U8419 ( .C1(n10434), .C2(n9636), .A(n7122), .B(n7121), .ZN(n7123)
         );
  INV_X1 U8420 ( .A(n7123), .ZN(n7124) );
  NAND2_X1 U8421 ( .A1(n7125), .A2(n7124), .ZN(P1_U3214) );
  NOR2_X1 U8422 ( .A1(n7126), .A2(P1_U3086), .ZN(n7127) );
  INV_X1 U8423 ( .A(n7505), .ZN(n7128) );
  OR2_X1 U8424 ( .A1(n9018), .A2(n7128), .ZN(n7129) );
  NAND2_X1 U8425 ( .A1(n7129), .A2(n8118), .ZN(n7182) );
  NAND2_X1 U8426 ( .A1(n7182), .A2(n7130), .ZN(n7131) );
  NAND2_X1 U8427 ( .A1(n7131), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U8428 ( .A(n7150), .ZN(n7132) );
  AND2_X1 U8429 ( .A1(n8604), .A2(P2_U3151), .ZN(n8610) );
  INV_X1 U8430 ( .A(n8610), .ZN(n9513) );
  OAI222_X1 U8431 ( .A1(n9513), .A2(n7133), .B1(n8667), .B2(n7136), .C1(
        P2_U3151), .C2(n5231), .ZN(P2_U3294) );
  OAI222_X1 U8432 ( .A1(n9513), .A2(n5368), .B1(n8667), .B2(n6505), .C1(
        P2_U3151), .C2(n10982), .ZN(P2_U3291) );
  NAND2_X1 U8433 ( .A1(n7134), .A2(P1_U3086), .ZN(n8627) );
  INV_X2 U8434 ( .A(n10476), .ZN(n8633) );
  OAI222_X1 U8435 ( .A1(n8627), .A2(n7135), .B1(n8633), .B2(n6458), .C1(
        P1_U3086), .C2(n7388), .ZN(P1_U3353) );
  OAI222_X1 U8436 ( .A1(n8627), .A2(n5684), .B1(n8633), .B2(n7136), .C1(
        P1_U3086), .C2(n7310), .ZN(P1_U3354) );
  INV_X1 U8437 ( .A(n8627), .ZN(n7154) );
  AOI22_X1 U8438 ( .A1(n7342), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n7154), .ZN(n7137) );
  OAI21_X1 U8439 ( .B1(n7138), .B2(n8633), .A(n7137), .ZN(P1_U3350) );
  OAI222_X1 U8440 ( .A1(n9513), .A2(n7139), .B1(n8667), .B2(n7138), .C1(
        P2_U3151), .C2(n7271), .ZN(P2_U3290) );
  AOI22_X1 U8441 ( .A1(n7356), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n7154), .ZN(n7140) );
  OAI21_X1 U8442 ( .B1(n7142), .B2(n8633), .A(n7140), .ZN(P1_U3349) );
  INV_X1 U8443 ( .A(n7154), .ZN(n10471) );
  OAI222_X1 U8444 ( .A1(n10471), .A2(n7141), .B1(n8633), .B2(n6505), .C1(
        P1_U3086), .C2(n10022), .ZN(P1_U3351) );
  OAI222_X1 U8445 ( .A1(n9513), .A2(n7143), .B1(n8667), .B2(n7142), .C1(
        P2_U3151), .C2(n7637), .ZN(P2_U3289) );
  INV_X1 U8446 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n7147) );
  INV_X1 U8447 ( .A(n7145), .ZN(n7146) );
  AOI22_X1 U8448 ( .A1(n7157), .A2(n7147), .B1(n7150), .B2(n7146), .ZN(
        P2_U3376) );
  INV_X1 U8449 ( .A(n7148), .ZN(n7149) );
  AOI22_X1 U8450 ( .A1(n7157), .A2(n7151), .B1(n7150), .B2(n7149), .ZN(
        P2_U3377) );
  INV_X1 U8451 ( .A(n7152), .ZN(n7156) );
  AOI22_X1 U8452 ( .A1(n7867), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n8610), .ZN(n7153) );
  OAI21_X1 U8453 ( .B1(n7156), .B2(n8667), .A(n7153), .ZN(P2_U3288) );
  AOI22_X1 U8454 ( .A1(n7371), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n7154), .ZN(n7155) );
  OAI21_X1 U8455 ( .B1(n7156), .B2(n8633), .A(n7155), .ZN(P1_U3348) );
  AND2_X1 U8456 ( .A1(n7157), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8457 ( .A1(n7157), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8458 ( .A1(n7157), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8459 ( .A1(n7157), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8460 ( .A1(n7157), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8461 ( .A1(n7157), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8462 ( .A1(n7157), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8463 ( .A1(n7157), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8464 ( .A1(n7157), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8465 ( .A1(n7157), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8466 ( .A1(n7157), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8467 ( .A1(n7157), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8468 ( .A1(n7157), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8469 ( .A1(n7157), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8470 ( .A1(n7157), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8471 ( .A1(n7157), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8472 ( .A1(n7157), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8473 ( .A1(n7157), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8474 ( .A1(n7157), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8475 ( .A1(n7157), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8476 ( .A1(n7157), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8477 ( .A1(n7157), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8478 ( .A1(n7157), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8479 ( .A1(n7157), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8480 ( .A1(n7157), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8481 ( .A1(n7157), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8482 ( .A1(n7157), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8483 ( .A1(n7157), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8484 ( .A1(n7157), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8485 ( .A1(n7157), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  INV_X1 U8486 ( .A(n7158), .ZN(n7161) );
  OAI222_X1 U8487 ( .A1(n9513), .A2(n7159), .B1(n8667), .B2(n7161), .C1(
        P2_U3151), .C2(n7997), .ZN(P2_U3287) );
  INV_X1 U8488 ( .A(n7421), .ZN(n7160) );
  OAI222_X1 U8489 ( .A1(n8627), .A2(n10795), .B1(n8633), .B2(n7161), .C1(
        P1_U3086), .C2(n7160), .ZN(P1_U3347) );
  INV_X1 U8490 ( .A(n7162), .ZN(n7165) );
  AOI22_X1 U8491 ( .A1(n8183), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n8610), .ZN(n7163) );
  OAI21_X1 U8492 ( .B1(n7165), .B2(n8667), .A(n7163), .ZN(P2_U3286) );
  INV_X1 U8493 ( .A(n10044), .ZN(n7164) );
  OAI222_X1 U8494 ( .A1(n8627), .A2(n10595), .B1(n8633), .B2(n7165), .C1(n7164), .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U8495 ( .A(n7166), .ZN(n7168) );
  OAI222_X1 U8496 ( .A1(n8667), .A2(n7168), .B1(n8269), .B2(P2_U3151), .C1(
        n7167), .C2(n9513), .ZN(P2_U3285) );
  INV_X1 U8497 ( .A(n7617), .ZN(n7422) );
  OAI222_X1 U8498 ( .A1(n8627), .A2(n7169), .B1(n8633), .B2(n7168), .C1(n7422), 
        .C2(P1_U3086), .ZN(P1_U3345) );
  NAND2_X1 U8499 ( .A1(n8114), .A2(n7170), .ZN(n7171) );
  NAND2_X1 U8500 ( .A1(n7171), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7249) );
  INV_X1 U8501 ( .A(n7249), .ZN(n7173) );
  INV_X1 U8502 ( .A(n9808), .ZN(n9817) );
  NAND2_X1 U8503 ( .A1(n9817), .A2(n8114), .ZN(n7172) );
  NAND2_X1 U8504 ( .A1(n7172), .A2(n5889), .ZN(n7250) );
  AND2_X1 U8505 ( .A1(n7173), .A2(n7250), .ZN(n10119) );
  NOR2_X1 U8506 ( .A1(n10119), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8507 ( .A(n8118), .ZN(n7174) );
  NOR2_X1 U8508 ( .A1(n7505), .A2(n7174), .ZN(n7175) );
  INV_X1 U8509 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n7186) );
  NOR2_X1 U8510 ( .A1(n6837), .A2(P2_U3151), .ZN(n8483) );
  AND2_X1 U8511 ( .A1(n8483), .A2(n7182), .ZN(n7203) );
  INV_X1 U8512 ( .A(n7203), .ZN(n7202) );
  NAND2_X1 U8513 ( .A1(P2_U3893), .A2(n6837), .ZN(n9164) );
  MUX2_X1 U8514 ( .A(P2_REG2_REG_0__SCAN_IN), .B(P2_REG1_REG_0__SCAN_IN), .S(
        n8174), .Z(n7179) );
  INV_X1 U8515 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7177) );
  INV_X1 U8516 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n7176) );
  MUX2_X1 U8517 ( .A(n7177), .B(n7176), .S(n8174), .Z(n7178) );
  AND2_X1 U8518 ( .A1(n7178), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n10953) );
  AOI21_X1 U8519 ( .B1(n7204), .B2(n7179), .A(n10953), .ZN(n7180) );
  AOI21_X1 U8520 ( .B1(n7202), .B2(n9164), .A(n7180), .ZN(n7181) );
  AOI21_X1 U8521 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .A(n7181), .ZN(
        n7185) );
  NOR2_X1 U8522 ( .A1(n8174), .A2(P2_U3151), .ZN(n8381) );
  NAND2_X1 U8523 ( .A1(n7182), .A2(n8381), .ZN(n7183) );
  MUX2_X1 U8524 ( .A(n9045), .B(n7183), .S(n6837), .Z(n10983) );
  NAND2_X1 U8525 ( .A1(n10997), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n7184) );
  OAI211_X1 U8526 ( .C1(n9095), .C2(n7186), .A(n7185), .B(n7184), .ZN(P2_U3182) );
  INV_X1 U8527 ( .A(n7187), .ZN(n7190) );
  OAI222_X1 U8528 ( .A1(n9513), .A2(n7188), .B1(n8667), .B2(n7190), .C1(
        P2_U3151), .C2(n8271), .ZN(P2_U3284) );
  INV_X1 U8529 ( .A(n7819), .ZN(n7189) );
  OAI222_X1 U8530 ( .A1(n10471), .A2(n10792), .B1(n8633), .B2(n7190), .C1(
        P1_U3086), .C2(n7189), .ZN(P1_U3344) );
  NAND2_X1 U8531 ( .A1(P1_U3973), .A2(n9562), .ZN(n7191) );
  OAI21_X1 U8532 ( .B1(P1_U3973), .B2(n6694), .A(n7191), .ZN(P1_U3574) );
  INV_X1 U8533 ( .A(P1_U3973), .ZN(n7530) );
  NAND2_X1 U8534 ( .A1(n7530), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n7192) );
  OAI21_X1 U8535 ( .B1(n7530), .B2(n10297), .A(n7192), .ZN(P1_U3571) );
  INV_X4 U8536 ( .A(n7193), .ZN(n8174) );
  MUX2_X1 U8537 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8174), .Z(n7221) );
  XOR2_X1 U8538 ( .A(n8623), .B(n7221), .Z(n7224) );
  MUX2_X1 U8539 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n8174), .Z(n7194) );
  XNOR2_X1 U8540 ( .A(n7194), .B(n5231), .ZN(n10952) );
  INV_X1 U8541 ( .A(n5231), .ZN(n10936) );
  INV_X1 U8542 ( .A(n7194), .ZN(n7195) );
  MUX2_X1 U8543 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8174), .Z(n7196) );
  INV_X1 U8544 ( .A(n5128), .ZN(n10963) );
  XNOR2_X1 U8545 ( .A(n7196), .B(n10963), .ZN(n10974) );
  AOI22_X1 U8546 ( .A1(n10973), .A2(n10974), .B1(n7196), .B2(n5128), .ZN(n7225) );
  XOR2_X1 U8547 ( .A(n7224), .B(n7225), .Z(n7220) );
  INV_X1 U8548 ( .A(n9095), .ZN(n10996) );
  NOR2_X1 U8549 ( .A1(n10983), .A2(n8623), .ZN(n7218) );
  INV_X1 U8550 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7475) );
  AND2_X1 U8551 ( .A1(n7204), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7197) );
  NAND2_X1 U8552 ( .A1(n7205), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7198) );
  OAI21_X1 U8553 ( .B1(n7207), .B2(n7197), .A(n7198), .ZN(n10944) );
  INV_X1 U8554 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10943) );
  NAND2_X1 U8555 ( .A1(n10946), .A2(n7198), .ZN(n10958) );
  NAND2_X1 U8556 ( .A1(n10959), .A2(n10958), .ZN(n10957) );
  NAND2_X1 U8557 ( .A1(n5128), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7199) );
  INV_X1 U8558 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7453) );
  AOI21_X1 U8559 ( .B1(n7201), .B2(n7453), .A(n5222), .ZN(n7216) );
  INV_X1 U8560 ( .A(n8623), .ZN(n7223) );
  INV_X1 U8561 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7982) );
  AND2_X1 U8562 ( .A1(n7204), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7206) );
  NAND2_X1 U8563 ( .A1(n7205), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7208) );
  OAI21_X1 U8564 ( .B1(n7207), .B2(n7206), .A(n7208), .ZN(n10938) );
  INV_X1 U8565 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10937) );
  NAND2_X1 U8566 ( .A1(n10940), .A2(n7208), .ZN(n10965) );
  NAND2_X1 U8567 ( .A1(n5128), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7209) );
  NAND2_X1 U8568 ( .A1(n7210), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7228) );
  INV_X1 U8569 ( .A(n7210), .ZN(n7212) );
  INV_X1 U8570 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7211) );
  NAND2_X1 U8571 ( .A1(n7212), .A2(n7211), .ZN(n7213) );
  NAND2_X1 U8572 ( .A1(n7228), .A2(n7213), .ZN(n7214) );
  NAND2_X1 U8573 ( .A1(n10968), .A2(n7214), .ZN(n7215) );
  NAND2_X1 U8574 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7650) );
  OAI211_X1 U8575 ( .C1(n7216), .C2(n11005), .A(n7215), .B(n7650), .ZN(n7217)
         );
  AOI211_X1 U8576 ( .C1(n10996), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n7218), .B(
        n7217), .ZN(n7219) );
  OAI21_X1 U8577 ( .B1(n7220), .B2(n9164), .A(n7219), .ZN(P2_U3185) );
  MUX2_X1 U8578 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8174), .Z(n7226) );
  INV_X1 U8579 ( .A(n7226), .ZN(n7227) );
  INV_X1 U8580 ( .A(n7221), .ZN(n7222) );
  XNOR2_X1 U8581 ( .A(n7226), .B(n5127), .ZN(n10986) );
  NAND2_X1 U8582 ( .A1(n10987), .A2(n10986), .ZN(n10985) );
  OAI21_X1 U8583 ( .B1(n5127), .B2(n7227), .A(n10985), .ZN(n7274) );
  MUX2_X1 U8584 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8174), .Z(n7272) );
  XNOR2_X1 U8585 ( .A(n7272), .B(n7244), .ZN(n7273) );
  XNOR2_X1 U8586 ( .A(n7274), .B(n7273), .ZN(n7246) );
  INV_X1 U8587 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n7237) );
  INV_X1 U8588 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7230) );
  MUX2_X1 U8589 ( .A(n7230), .B(P2_REG2_REG_4__SCAN_IN), .S(n5127), .Z(n7231)
         );
  INV_X1 U8590 ( .A(n7231), .ZN(n10989) );
  OR2_X1 U8591 ( .A1(n5127), .A2(n7230), .ZN(n7232) );
  OAI21_X1 U8592 ( .B1(n5220), .B2(P2_REG2_REG_5__SCAN_IN), .A(n7290), .ZN(
        n7235) );
  NAND2_X1 U8593 ( .A1(n10968), .A2(n7235), .ZN(n7236) );
  NAND2_X1 U8594 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7670) );
  OAI211_X1 U8595 ( .C1(n9095), .C2(n7237), .A(n7236), .B(n7670), .ZN(n7243)
         );
  INV_X1 U8596 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7844) );
  AOI22_X1 U8597 ( .A1(n5127), .A2(P2_REG1_REG_4__SCAN_IN), .B1(n7844), .B2(
        n10982), .ZN(n10979) );
  NOR2_X1 U8598 ( .A1(n5127), .A2(n7844), .ZN(n7239) );
  INV_X1 U8599 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n8018) );
  NOR2_X1 U8600 ( .A1(n7241), .A2(n11005), .ZN(n7242) );
  AOI211_X1 U8601 ( .C1(n10997), .C2(n7244), .A(n7243), .B(n7242), .ZN(n7245)
         );
  OAI21_X1 U8602 ( .B1(n7246), .B2(n9164), .A(n7245), .ZN(P2_U3187) );
  INV_X1 U8603 ( .A(n8453), .ZN(n7378) );
  INV_X1 U8604 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n11028) );
  INV_X1 U8605 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7247) );
  AOI21_X1 U8606 ( .B1(n7378), .B2(n7247), .A(n8497), .ZN(n7380) );
  OAI21_X1 U8607 ( .B1(n7378), .B2(P1_REG1_REG_0__SCAN_IN), .A(n7380), .ZN(
        n7248) );
  MUX2_X1 U8608 ( .A(n7248), .B(n7380), .S(P1_IR_REG_0__SCAN_IN), .Z(n7254) );
  INV_X1 U8609 ( .A(n10125), .ZN(n10877) );
  NAND3_X1 U8610 ( .A1(n10877), .A2(P1_IR_REG_0__SCAN_IN), .A3(n11028), .ZN(
        n7253) );
  INV_X1 U8611 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7600) );
  NOR2_X1 U8612 ( .A1(n7600), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7251) );
  AOI21_X1 U8613 ( .B1(n10119), .B2(P1_ADDR_REG_0__SCAN_IN), .A(n7251), .ZN(
        n7252) );
  OAI211_X1 U8614 ( .C1(n7254), .C2(n7259), .A(n7253), .B(n7252), .ZN(P1_U3243) );
  INV_X1 U8615 ( .A(n7255), .ZN(n7257) );
  INV_X1 U8616 ( .A(n8273), .ZN(n8577) );
  INV_X1 U8617 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7256) );
  OAI222_X1 U8618 ( .A1(n8667), .A2(n7257), .B1(n8577), .B2(P2_U3151), .C1(
        n7256), .C2(n9513), .ZN(P2_U3283) );
  INV_X1 U8619 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10655) );
  OAI222_X1 U8620 ( .A1(n10471), .A2(n10655), .B1(n8633), .B2(n7257), .C1(
        n8434), .C2(P1_U3086), .ZN(P1_U3343) );
  NAND2_X1 U8621 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n7379) );
  XOR2_X1 U8622 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n7310), .Z(n7260) );
  NOR2_X1 U8623 ( .A1(n7260), .A2(n7379), .ZN(n7311) );
  NAND2_X1 U8624 ( .A1(n7258), .A2(n7378), .ZN(n9699) );
  AOI211_X1 U8625 ( .C1(n7379), .C2(n7260), .A(n7311), .B(n8444), .ZN(n7266)
         );
  NAND2_X1 U8626 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n7264) );
  INV_X1 U8627 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n7261) );
  XNOR2_X1 U8628 ( .A(n7310), .B(n7261), .ZN(n7263) );
  INV_X1 U8629 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7262) );
  NOR3_X1 U8630 ( .A1(n7263), .A2(n11028), .A3(n7262), .ZN(n7317) );
  AOI211_X1 U8631 ( .C1(n7264), .C2(n7263), .A(n7317), .B(n10125), .ZN(n7265)
         );
  NOR2_X1 U8632 ( .A1(n7266), .A2(n7265), .ZN(n7268) );
  AOI22_X1 U8633 ( .A1(n10119), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n7267) );
  OAI211_X1 U8634 ( .C1(n7310), .C2(n10121), .A(n7268), .B(n7267), .ZN(
        P1_U3244) );
  INV_X1 U8635 ( .A(n8475), .ZN(n8016) );
  INV_X1 U8636 ( .A(n7542), .ZN(n9052) );
  NAND2_X1 U8637 ( .A1(n9052), .A2(n7593), .ZN(n8884) );
  NAND2_X1 U8638 ( .A1(n8884), .A2(n7429), .ZN(n8885) );
  OAI21_X1 U8639 ( .B1(n9342), .B2(n9414), .A(n8885), .ZN(n7269) );
  NAND2_X1 U8640 ( .A1(n9051), .A2(n9337), .ZN(n7591) );
  OAI211_X1 U8641 ( .C1(n9450), .C2(n7593), .A(n7269), .B(n7591), .ZN(n7329)
         );
  NAND2_X1 U8642 ( .A1(n7329), .A2(n9456), .ZN(n7270) );
  OAI21_X1 U8643 ( .B1(n9456), .B2(n7176), .A(n7270), .ZN(P2_U3459) );
  AOI22_X1 U8644 ( .A1(n7274), .A2(n7273), .B1(n7272), .B2(n7271), .ZN(n7277)
         );
  MUX2_X1 U8645 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8174), .Z(n7275) );
  NOR2_X1 U8646 ( .A1(n7275), .A2(n7637), .ZN(n7632) );
  AOI21_X1 U8647 ( .B1(n7275), .B2(n7637), .A(n7632), .ZN(n7276) );
  AND2_X1 U8648 ( .A1(n7277), .A2(n7276), .ZN(n7631) );
  NOR2_X1 U8649 ( .A1(n7277), .A2(n7276), .ZN(n7278) );
  OAI21_X1 U8650 ( .B1(n7631), .B2(n7278), .A(n11010), .ZN(n7300) );
  INV_X1 U8651 ( .A(n7279), .ZN(n7280) );
  INV_X1 U8652 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n8165) );
  MUX2_X1 U8653 ( .A(n8165), .B(P2_REG1_REG_6__SCAN_IN), .S(n7287), .Z(n7282)
         );
  INV_X1 U8654 ( .A(n7282), .ZN(n7285) );
  INV_X1 U8655 ( .A(n7283), .ZN(n7284) );
  NAND2_X1 U8656 ( .A1(n7285), .A2(n7284), .ZN(n7286) );
  AND2_X1 U8657 ( .A1(n7625), .A2(n7286), .ZN(n7295) );
  INV_X1 U8658 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7288) );
  MUX2_X1 U8659 ( .A(n7288), .B(P2_REG2_REG_6__SCAN_IN), .S(n7287), .Z(n7292)
         );
  NAND2_X1 U8660 ( .A1(n7290), .A2(n7289), .ZN(n7291) );
  NAND2_X1 U8661 ( .A1(n7291), .A2(n7292), .ZN(n7639) );
  OAI21_X1 U8662 ( .B1(n7292), .B2(n7291), .A(n7639), .ZN(n7293) );
  NAND2_X1 U8663 ( .A1(n10968), .A2(n7293), .ZN(n7294) );
  NAND2_X1 U8664 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7785) );
  OAI211_X1 U8665 ( .C1(n7295), .C2(n11005), .A(n7294), .B(n7785), .ZN(n7298)
         );
  INV_X1 U8666 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7296) );
  NOR2_X1 U8667 ( .A1(n9095), .A2(n7296), .ZN(n7297) );
  NOR2_X1 U8668 ( .A1(n7298), .A2(n7297), .ZN(n7299) );
  OAI211_X1 U8669 ( .C1(n10983), .C2(n7637), .A(n7300), .B(n7299), .ZN(
        P2_U3188) );
  OAI21_X1 U8670 ( .B1(n7303), .B2(n7301), .A(n7302), .ZN(n7383) );
  NAND2_X1 U8671 ( .A1(n7305), .A2(n7304), .ZN(n7442) );
  AOI22_X1 U8672 ( .A1(n9687), .A2(n6332), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n7442), .ZN(n7307) );
  NAND2_X1 U8673 ( .A1(n9694), .A2(n11024), .ZN(n7306) );
  OAI211_X1 U8674 ( .C1(n9697), .C2(n7383), .A(n7307), .B(n7306), .ZN(P1_U3232) );
  INV_X1 U8675 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n7309) );
  NAND2_X1 U8676 ( .A1(n10866), .A2(n7342), .ZN(n7308) );
  NAND2_X1 U8677 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7986) );
  OAI211_X1 U8678 ( .C1(n7309), .C2(n10869), .A(n7308), .B(n7986), .ZN(n7328)
         );
  INV_X1 U8679 ( .A(n10022), .ZN(n7323) );
  INV_X1 U8680 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7557) );
  INV_X1 U8681 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7313) );
  INV_X1 U8682 ( .A(n7310), .ZN(n7318) );
  AOI21_X1 U8683 ( .B1(P1_REG2_REG_1__SCAN_IN), .B2(n7318), .A(n7311), .ZN(
        n7386) );
  XOR2_X1 U8684 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n7388), .Z(n7385) );
  NOR2_X1 U8685 ( .A1(n7386), .A2(n7385), .ZN(n7384) );
  INV_X1 U8686 ( .A(n7384), .ZN(n7312) );
  OAI21_X1 U8687 ( .B1(n7313), .B2(n7388), .A(n7312), .ZN(n10013) );
  XNOR2_X1 U8688 ( .A(n10006), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n10014) );
  NAND2_X1 U8689 ( .A1(n10013), .A2(n10014), .ZN(n10012) );
  OAI21_X1 U8690 ( .B1(n10006), .B2(n7557), .A(n10012), .ZN(n10029) );
  INV_X1 U8691 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7921) );
  MUX2_X1 U8692 ( .A(n7921), .B(P1_REG2_REG_4__SCAN_IN), .S(n10022), .Z(n10030) );
  NAND2_X1 U8693 ( .A1(n10029), .A2(n10030), .ZN(n10028) );
  INV_X1 U8694 ( .A(n10028), .ZN(n7314) );
  AOI21_X1 U8695 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n7323), .A(n7314), .ZN(
        n7316) );
  XNOR2_X1 U8696 ( .A(n7342), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n7315) );
  NOR2_X1 U8697 ( .A1(n7316), .A2(n7315), .ZN(n7336) );
  AOI211_X1 U8698 ( .C1(n7316), .C2(n7315), .A(n8444), .B(n7336), .ZN(n7327)
         );
  INV_X1 U8699 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7321) );
  INV_X1 U8700 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n7320) );
  AOI21_X1 U8701 ( .B1(P1_REG1_REG_1__SCAN_IN), .B2(n7318), .A(n7317), .ZN(
        n7391) );
  XOR2_X1 U8702 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n7388), .Z(n7390) );
  NOR2_X1 U8703 ( .A1(n7391), .A2(n7390), .ZN(n7389) );
  INV_X1 U8704 ( .A(n7389), .ZN(n7319) );
  OAI21_X1 U8705 ( .B1(n7320), .B2(n7388), .A(n7319), .ZN(n10016) );
  XNOR2_X1 U8706 ( .A(n10006), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n10017) );
  NAND2_X1 U8707 ( .A1(n10016), .A2(n10017), .ZN(n10015) );
  OAI21_X1 U8708 ( .B1(n10006), .B2(n7321), .A(n10015), .ZN(n10026) );
  INV_X1 U8709 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n8070) );
  MUX2_X1 U8710 ( .A(n8070), .B(P1_REG1_REG_4__SCAN_IN), .S(n10022), .Z(n10027) );
  NAND2_X1 U8711 ( .A1(n10026), .A2(n10027), .ZN(n10025) );
  INV_X1 U8712 ( .A(n10025), .ZN(n7322) );
  AOI21_X1 U8713 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n7323), .A(n7322), .ZN(
        n7325) );
  XNOR2_X1 U8714 ( .A(n7342), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n7324) );
  NOR2_X1 U8715 ( .A1(n7325), .A2(n7324), .ZN(n7341) );
  AOI211_X1 U8716 ( .C1(n7325), .C2(n7324), .A(n10125), .B(n7341), .ZN(n7326)
         );
  OR3_X1 U8717 ( .A1(n7328), .A2(n7327), .A3(n7326), .ZN(P1_U3248) );
  INV_X1 U8718 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7331) );
  NAND2_X1 U8719 ( .A1(n7329), .A2(n11121), .ZN(n7330) );
  OAI21_X1 U8720 ( .B1(n11121), .B2(n7331), .A(n7330), .ZN(P2_U3390) );
  INV_X1 U8721 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n7333) );
  INV_X1 U8722 ( .A(n7332), .ZN(n7334) );
  INV_X1 U8723 ( .A(n10049), .ZN(n8422) );
  OAI222_X1 U8724 ( .A1(n8627), .A2(n7333), .B1(n8633), .B2(n7334), .C1(
        P1_U3086), .C2(n8422), .ZN(P1_U3342) );
  INV_X1 U8725 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7335) );
  OAI222_X1 U8726 ( .A1(n9513), .A2(n7335), .B1(n8667), .B2(n7334), .C1(
        P2_U3151), .C2(n5497), .ZN(P2_U3282) );
  AOI21_X1 U8727 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n7342), .A(n7336), .ZN(
        n7340) );
  INV_X1 U8728 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7337) );
  MUX2_X1 U8729 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n7337), .S(n7356), .Z(n7338)
         );
  INV_X1 U8730 ( .A(n7338), .ZN(n7339) );
  NOR2_X1 U8731 ( .A1(n7340), .A2(n7339), .ZN(n7355) );
  AOI211_X1 U8732 ( .C1(n7340), .C2(n7339), .A(n8444), .B(n7355), .ZN(n7350)
         );
  AOI21_X1 U8733 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n7342), .A(n7341), .ZN(
        n7345) );
  INV_X1 U8734 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7343) );
  MUX2_X1 U8735 ( .A(n7343), .B(P1_REG1_REG_6__SCAN_IN), .S(n7356), .Z(n7344)
         );
  NOR2_X1 U8736 ( .A1(n7345), .A2(n7344), .ZN(n7351) );
  AOI211_X1 U8737 ( .C1(n7345), .C2(n7344), .A(n10125), .B(n7351), .ZN(n7349)
         );
  INV_X1 U8738 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n7347) );
  NAND2_X1 U8739 ( .A1(n10866), .A2(n7356), .ZN(n7346) );
  NAND2_X1 U8740 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8023) );
  OAI211_X1 U8741 ( .C1(n7347), .C2(n10869), .A(n7346), .B(n8023), .ZN(n7348)
         );
  OR3_X1 U8742 ( .A1(n7350), .A2(n7349), .A3(n7348), .ZN(P1_U3249) );
  AOI21_X1 U8743 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n7356), .A(n7351), .ZN(
        n7367) );
  NAND2_X1 U8744 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n7371), .ZN(n7352) );
  OAI21_X1 U8745 ( .B1(n7371), .B2(P1_REG1_REG_7__SCAN_IN), .A(n7352), .ZN(
        n7366) );
  NOR2_X1 U8746 ( .A1(n7367), .A2(n7366), .ZN(n7365) );
  AOI21_X1 U8747 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n7371), .A(n7365), .ZN(
        n7354) );
  XNOR2_X1 U8748 ( .A(n7421), .B(P1_REG1_REG_8__SCAN_IN), .ZN(n7353) );
  NOR2_X1 U8749 ( .A1(n7354), .A2(n7353), .ZN(n7415) );
  AOI211_X1 U8750 ( .C1(n7354), .C2(n7353), .A(n10125), .B(n7415), .ZN(n7364)
         );
  AOI21_X1 U8751 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n7356), .A(n7355), .ZN(
        n7370) );
  NAND2_X1 U8752 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n7371), .ZN(n7357) );
  OAI21_X1 U8753 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n7371), .A(n7357), .ZN(
        n7369) );
  NOR2_X1 U8754 ( .A1(n7370), .A2(n7369), .ZN(n7368) );
  AOI21_X1 U8755 ( .B1(n7371), .B2(P1_REG2_REG_7__SCAN_IN), .A(n7368), .ZN(
        n7359) );
  XNOR2_X1 U8756 ( .A(n7421), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n7358) );
  NOR2_X1 U8757 ( .A1(n7358), .A2(n7359), .ZN(n7420) );
  AOI211_X1 U8758 ( .C1(n7359), .C2(n7358), .A(n7420), .B(n8444), .ZN(n7363)
         );
  INV_X1 U8759 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n7361) );
  NAND2_X1 U8760 ( .A1(n10866), .A2(n7421), .ZN(n7360) );
  NAND2_X1 U8761 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n8233) );
  OAI211_X1 U8762 ( .C1(n7361), .C2(n10869), .A(n7360), .B(n8233), .ZN(n7362)
         );
  OR3_X1 U8763 ( .A1(n7364), .A2(n7363), .A3(n7362), .ZN(P1_U3251) );
  AOI211_X1 U8764 ( .C1(n7367), .C2(n7366), .A(n10125), .B(n7365), .ZN(n7376)
         );
  AOI211_X1 U8765 ( .C1(n7370), .C2(n7369), .A(n7368), .B(n8444), .ZN(n7375)
         );
  INV_X1 U8766 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n7373) );
  NAND2_X1 U8767 ( .A1(n10866), .A2(n7371), .ZN(n7372) );
  NAND2_X1 U8768 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n8139) );
  OAI211_X1 U8769 ( .C1(n7373), .C2(n10869), .A(n7372), .B(n8139), .ZN(n7374)
         );
  OR3_X1 U8770 ( .A1(n7376), .A2(n7375), .A3(n7374), .ZN(P1_U3250) );
  NAND2_X1 U8771 ( .A1(n8659), .A2(P2_U3893), .ZN(n7377) );
  OAI21_X1 U8772 ( .B1(P2_U3893), .B2(n8116), .A(n7377), .ZN(P2_U3514) );
  NOR2_X1 U8773 ( .A1(n8497), .A2(n7378), .ZN(n7382) );
  OAI22_X1 U8774 ( .A1(n7380), .A2(P1_IR_REG_0__SCAN_IN), .B1(n7379), .B2(
        n9699), .ZN(n7381) );
  AOI211_X1 U8775 ( .C1(n7383), .C2(n7382), .A(n7530), .B(n7381), .ZN(n10021)
         );
  AOI211_X1 U8776 ( .C1(n7386), .C2(n7385), .A(n7384), .B(n8444), .ZN(n7394)
         );
  AOI22_X1 U8777 ( .A1(n10119), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n7387) );
  OAI21_X1 U8778 ( .B1(n7388), .B2(n10121), .A(n7387), .ZN(n7393) );
  AOI211_X1 U8779 ( .C1(n7391), .C2(n7390), .A(n7389), .B(n10125), .ZN(n7392)
         );
  OR4_X1 U8780 ( .A1(n10021), .A2(n7394), .A3(n7393), .A4(n7392), .ZN(P1_U3245) );
  INV_X1 U8781 ( .A(n7395), .ZN(n7396) );
  INV_X1 U8782 ( .A(n10063), .ZN(n8425) );
  OAI222_X1 U8783 ( .A1(n8627), .A2(n10593), .B1(n8633), .B2(n7396), .C1(
        P1_U3086), .C2(n8425), .ZN(P1_U3341) );
  OAI222_X1 U8784 ( .A1(n9513), .A2(n7397), .B1(n8667), .B2(n7396), .C1(
        P2_U3151), .C2(n9081), .ZN(P2_U3281) );
  INV_X1 U8785 ( .A(n7398), .ZN(n7403) );
  AOI21_X1 U8786 ( .B1(n7402), .B2(n7400), .A(n7399), .ZN(n7401) );
  AOI21_X1 U8787 ( .B1(n7403), .B2(n7402), .A(n7401), .ZN(n7407) );
  NOR2_X1 U8788 ( .A1(n9636), .A2(n11034), .ZN(n7405) );
  INV_X1 U8789 ( .A(n10005), .ZN(n7569) );
  OAI22_X1 U8790 ( .A1(n7569), .A2(n9691), .B1(n9644), .B2(n7568), .ZN(n7404)
         );
  AOI211_X1 U8791 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(n7442), .A(n7405), .B(
        n7404), .ZN(n7406) );
  OAI21_X1 U8792 ( .B1(n7407), .B2(n9697), .A(n7406), .ZN(P1_U3222) );
  INV_X1 U8793 ( .A(n7408), .ZN(n7410) );
  AOI22_X1 U8794 ( .A1(n9103), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n8610), .ZN(n7409) );
  OAI21_X1 U8795 ( .B1(n7410), .B2(n8667), .A(n7409), .ZN(P2_U3280) );
  INV_X1 U8796 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7411) );
  INV_X1 U8797 ( .A(n10865), .ZN(n8441) );
  OAI222_X1 U8798 ( .A1(n8627), .A2(n7411), .B1(n8633), .B2(n7410), .C1(n8441), 
        .C2(P1_U3086), .ZN(P1_U3340) );
  INV_X1 U8799 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7413) );
  NAND2_X1 U8800 ( .A1(n10866), .A2(n7617), .ZN(n7412) );
  NAND2_X1 U8801 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n9543) );
  OAI211_X1 U8802 ( .C1(n7413), .C2(n10869), .A(n7412), .B(n9543), .ZN(n7428)
         );
  NOR2_X1 U8803 ( .A1(n10044), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7414) );
  AOI21_X1 U8804 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n10044), .A(n7414), .ZN(
        n10036) );
  AOI21_X1 U8805 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n7421), .A(n7415), .ZN(
        n10037) );
  NAND2_X1 U8806 ( .A1(n10036), .A2(n10037), .ZN(n10035) );
  OAI21_X1 U8807 ( .B1(n10044), .B2(P1_REG1_REG_9__SCAN_IN), .A(n10035), .ZN(
        n7418) );
  INV_X1 U8808 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7416) );
  MUX2_X1 U8809 ( .A(n7416), .B(P1_REG1_REG_10__SCAN_IN), .S(n7617), .Z(n7417)
         );
  NOR2_X1 U8810 ( .A1(n7417), .A2(n7418), .ZN(n7612) );
  AOI211_X1 U8811 ( .C1(n7418), .C2(n7417), .A(n7612), .B(n10125), .ZN(n7427)
         );
  NOR2_X1 U8812 ( .A1(n10044), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7419) );
  AOI21_X1 U8813 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n10044), .A(n7419), .ZN(
        n10042) );
  AOI21_X1 U8814 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n7421), .A(n7420), .ZN(
        n10041) );
  NAND2_X1 U8815 ( .A1(n10042), .A2(n10041), .ZN(n10040) );
  OAI21_X1 U8816 ( .B1(n10044), .B2(P1_REG2_REG_9__SCAN_IN), .A(n10040), .ZN(
        n7425) );
  INV_X1 U8817 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7423) );
  AOI22_X1 U8818 ( .A1(n7617), .A2(n7423), .B1(P1_REG2_REG_10__SCAN_IN), .B2(
        n7422), .ZN(n7424) );
  NOR2_X1 U8819 ( .A1(n7425), .A2(n7424), .ZN(n7616) );
  AOI211_X1 U8820 ( .C1(n7425), .C2(n7424), .A(n7616), .B(n8444), .ZN(n7426)
         );
  OR3_X1 U8821 ( .A1(n7428), .A2(n7427), .A3(n7426), .ZN(P1_U3253) );
  INV_X1 U8822 ( .A(n7429), .ZN(n7431) );
  OAI21_X1 U8823 ( .B1(n7433), .B2(n7431), .A(n7430), .ZN(n8029) );
  NOR2_X1 U8824 ( .A1(n7432), .A2(n9450), .ZN(n7435) );
  AOI21_X1 U8825 ( .B1(n7481), .B2(n7433), .A(n7469), .ZN(n7434) );
  OAI222_X1 U8826 ( .A1(n9376), .A2(n7486), .B1(n9361), .B2(n7542), .C1(n9373), 
        .C2(n7434), .ZN(n8030) );
  AOI211_X1 U8827 ( .C1(n9414), .C2(n8029), .A(n7435), .B(n8030), .ZN(n11032)
         );
  OR2_X1 U8828 ( .A1(n11032), .A2(n9465), .ZN(n7436) );
  OAI21_X1 U8829 ( .B1(n9456), .B2(n10943), .A(n7436), .ZN(P2_U3460) );
  XOR2_X1 U8830 ( .A(n7438), .B(n7437), .Z(n7444) );
  NOR2_X1 U8831 ( .A1(n9636), .A2(n8074), .ZN(n7441) );
  OAI22_X1 U8832 ( .A1(n5968), .A2(n9691), .B1(n9644), .B2(n7439), .ZN(n7440)
         );
  AOI211_X1 U8833 ( .C1(P1_REG3_REG_2__SCAN_IN), .C2(n7442), .A(n7441), .B(
        n7440), .ZN(n7443) );
  OAI21_X1 U8834 ( .B1(n9697), .B2(n7444), .A(n7443), .ZN(P1_U3237) );
  INV_X1 U8835 ( .A(n7447), .ZN(n8850) );
  NAND3_X1 U8836 ( .A1(n7464), .A2(n8888), .A3(n8850), .ZN(n7445) );
  NAND2_X1 U8837 ( .A1(n7446), .A2(n7445), .ZN(n7974) );
  XNOR2_X1 U8838 ( .A(n7448), .B(n7447), .ZN(n7449) );
  AOI21_X1 U8839 ( .B1(n9414), .B2(n7974), .A(n7971), .ZN(n7456) );
  INV_X1 U8840 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7450) );
  OAI22_X1 U8841 ( .A1(n9508), .A2(n7970), .B1(n11121), .B2(n7450), .ZN(n7451)
         );
  INV_X1 U8842 ( .A(n7451), .ZN(n7452) );
  OAI21_X1 U8843 ( .B1(n7456), .B2(n6890), .A(n7452), .ZN(P2_U3399) );
  OAI22_X1 U8844 ( .A1(n9432), .A2(n7970), .B1(n9456), .B2(n7453), .ZN(n7454)
         );
  INV_X1 U8845 ( .A(n7454), .ZN(n7455) );
  OAI21_X1 U8846 ( .B1(n7456), .B2(n9465), .A(n7455), .ZN(P2_U3462) );
  XOR2_X1 U8847 ( .A(n7458), .B(n7457), .Z(n7463) );
  AOI22_X1 U8848 ( .A1(n9678), .A2(n10004), .B1(n9687), .B2(n10002), .ZN(n7462) );
  NAND2_X1 U8849 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n10008) );
  INV_X1 U8850 ( .A(n10008), .ZN(n7460) );
  NOR2_X1 U8851 ( .A1(n9646), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n7459) );
  AOI211_X1 U8852 ( .C1(n5994), .C2(n9694), .A(n7460), .B(n7459), .ZN(n7461)
         );
  OAI211_X1 U8853 ( .C1(n7463), .C2(n9697), .A(n7462), .B(n7461), .ZN(P1_U3218) );
  OAI21_X1 U8854 ( .B1(n7465), .B2(n8892), .A(n7464), .ZN(n7979) );
  NOR2_X1 U8855 ( .A1(n7976), .A2(n9450), .ZN(n7473) );
  INV_X1 U8856 ( .A(n7467), .ZN(n7471) );
  NOR3_X1 U8857 ( .A1(n7469), .A2(n7468), .A3(n8849), .ZN(n7470) );
  NOR2_X1 U8858 ( .A1(n7471), .A2(n7470), .ZN(n7472) );
  OAI222_X1 U8859 ( .A1(n9376), .A2(n7839), .B1(n9361), .B2(n7466), .C1(n9373), 
        .C2(n7472), .ZN(n7978) );
  AOI211_X1 U8860 ( .C1(n9414), .C2(n7979), .A(n7473), .B(n7978), .ZN(n11042)
         );
  OR2_X1 U8861 ( .A1(n11042), .A2(n9465), .ZN(n7474) );
  OAI21_X1 U8862 ( .B1(n9456), .B2(n7475), .A(n7474), .ZN(P2_U3461) );
  NOR2_X1 U8863 ( .A1(n7480), .A2(n7482), .ZN(n7539) );
  NAND2_X1 U8864 ( .A1(n7539), .A2(n7540), .ZN(n7538) );
  INV_X1 U8865 ( .A(n7482), .ZN(n7483) );
  NAND2_X1 U8866 ( .A1(n7538), .A2(n7483), .ZN(n7531) );
  INV_X2 U8867 ( .A(n7484), .ZN(n8678) );
  INV_X1 U8868 ( .A(n8678), .ZN(n8684) );
  XNOR2_X1 U8869 ( .A(n7485), .B(n8684), .ZN(n7487) );
  NAND2_X1 U8870 ( .A1(n7532), .A2(n7488), .ZN(n7647) );
  XNOR2_X1 U8871 ( .A(n7970), .B(n8694), .ZN(n7489) );
  XNOR2_X1 U8872 ( .A(n7489), .B(n7839), .ZN(n7648) );
  NOR2_X1 U8873 ( .A1(n7647), .A2(n7648), .ZN(n7646) );
  INV_X1 U8874 ( .A(n7489), .ZN(n7490) );
  NOR2_X1 U8875 ( .A1(n7646), .A2(n5750), .ZN(n7493) );
  XNOR2_X1 U8876 ( .A(n8040), .B(n8694), .ZN(n7491) );
  NOR2_X1 U8877 ( .A1(n9048), .A2(n7491), .ZN(n7665) );
  AOI21_X1 U8878 ( .B1(n9048), .B2(n7491), .A(n7665), .ZN(n7492) );
  NAND2_X1 U8879 ( .A1(n7493), .A2(n7492), .ZN(n7667) );
  OAI21_X1 U8880 ( .B1(n7493), .B2(n7492), .A(n7667), .ZN(n7525) );
  NOR2_X1 U8881 ( .A1(n9463), .A2(n9018), .ZN(n7495) );
  INV_X1 U8882 ( .A(n7496), .ZN(n7494) );
  AOI21_X1 U8883 ( .B1(n7514), .B2(n7495), .A(n7494), .ZN(n7498) );
  OR2_X1 U8884 ( .A1(n7510), .A2(n7496), .ZN(n7506) );
  INV_X1 U8885 ( .A(n7506), .ZN(n7497) );
  INV_X1 U8886 ( .A(n7513), .ZN(n7499) );
  INV_X1 U8887 ( .A(n9027), .ZN(n7501) );
  AND2_X1 U8888 ( .A1(n7510), .A2(n7501), .ZN(n7519) );
  NAND2_X1 U8889 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n10994) );
  INV_X1 U8890 ( .A(n10994), .ZN(n7503) );
  AOI21_X1 U8891 ( .B1(n9049), .B2(n8827), .A(n7503), .ZN(n7523) );
  INV_X1 U8892 ( .A(n7504), .ZN(n7508) );
  AND3_X1 U8893 ( .A1(n7583), .A2(n7505), .A3(n8118), .ZN(n7507) );
  OAI211_X1 U8894 ( .C1(n7514), .C2(n7508), .A(n7507), .B(n7506), .ZN(n7509)
         );
  NAND2_X1 U8895 ( .A1(n7509), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7512) );
  OR2_X1 U8896 ( .A1(n9027), .A2(n7510), .ZN(n7511) );
  NAND2_X2 U8897 ( .A1(n7512), .A2(n7511), .ZN(n8831) );
  NAND2_X1 U8898 ( .A1(n8831), .A2(n8039), .ZN(n7522) );
  NAND2_X1 U8899 ( .A1(n7514), .A2(n9466), .ZN(n7517) );
  INV_X1 U8900 ( .A(n9466), .ZN(n7516) );
  NAND2_X1 U8901 ( .A1(n8786), .A2(n8040), .ZN(n7521) );
  NAND2_X1 U8902 ( .A1(n7519), .A2(n7518), .ZN(n8829) );
  OR2_X1 U8903 ( .A1(n8127), .A2(n8829), .ZN(n7520) );
  NAND4_X1 U8904 ( .A1(n7523), .A2(n7522), .A3(n7521), .A4(n7520), .ZN(n7524)
         );
  AOI21_X1 U8905 ( .B1(n7525), .B2(n8824), .A(n7524), .ZN(n7526) );
  INV_X1 U8906 ( .A(n7526), .ZN(P2_U3170) );
  NOR2_X1 U8907 ( .A1(n8831), .A2(P2_U3151), .ZN(n7547) );
  INV_X1 U8908 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10562) );
  OAI22_X1 U8909 ( .A1(n7466), .A2(n8829), .B1(n8835), .B2(n7593), .ZN(n7527)
         );
  AOI21_X1 U8910 ( .B1(n8885), .B2(n8824), .A(n7527), .ZN(n7528) );
  OAI21_X1 U8911 ( .B1(n7547), .B2(n10562), .A(n7528), .ZN(P2_U3172) );
  NAND2_X1 U8912 ( .A1(n7530), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7529) );
  OAI21_X1 U8913 ( .B1(n7530), .B2(n8714), .A(n7529), .ZN(P1_U3583) );
  INV_X1 U8914 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7537) );
  NAND2_X1 U8915 ( .A1(n7533), .A2(n8824), .ZN(n7536) );
  INV_X1 U8916 ( .A(n8827), .ZN(n8817) );
  OAI22_X1 U8917 ( .A1(n7466), .A2(n8817), .B1(n7976), .B2(n8835), .ZN(n7534)
         );
  AOI21_X1 U8918 ( .B1(n8815), .B2(n9049), .A(n7534), .ZN(n7535) );
  OAI211_X1 U8919 ( .C1(n7547), .C2(n7537), .A(n7536), .B(n7535), .ZN(P2_U3177) );
  INV_X1 U8920 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7546) );
  OAI21_X1 U8921 ( .B1(n7540), .B2(n7539), .A(n7538), .ZN(n7541) );
  NAND2_X1 U8922 ( .A1(n7541), .A2(n8824), .ZN(n7545) );
  OAI22_X1 U8923 ( .A1(n7542), .A2(n8817), .B1(n7432), .B2(n8835), .ZN(n7543)
         );
  AOI21_X1 U8924 ( .B1(n8815), .B2(n9050), .A(n7543), .ZN(n7544) );
  OAI211_X1 U8925 ( .C1(n7547), .C2(n7546), .A(n7545), .B(n7544), .ZN(P2_U3162) );
  OAI21_X1 U8926 ( .B1(n7550), .B2(n7549), .A(n7548), .ZN(n11047) );
  INV_X1 U8927 ( .A(n11047), .ZN(n7566) );
  NAND2_X1 U8928 ( .A1(n7552), .A2(n7551), .ZN(n7553) );
  INV_X2 U8929 ( .A(n10307), .ZN(n11079) );
  OR2_X1 U8930 ( .A1(n11079), .A2(n7743), .ZN(n7577) );
  INV_X1 U8931 ( .A(n7555), .ZN(n7692) );
  INV_X1 U8932 ( .A(n7684), .ZN(n7556) );
  OAI211_X1 U8933 ( .C1(n11044), .C2(n7692), .A(n7556), .B(n10400), .ZN(n11043) );
  NOR2_X1 U8934 ( .A1(n10219), .A2(n11043), .ZN(n7559) );
  OAI22_X1 U8935 ( .A1(n10307), .A2(n7557), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n7919), .ZN(n7558) );
  AOI211_X1 U8936 ( .C1(n10223), .C2(n5994), .A(n7559), .B(n7558), .ZN(n7565)
         );
  OAI21_X1 U8937 ( .B1(n9773), .B2(n9826), .A(n7560), .ZN(n7562) );
  OAI22_X1 U8938 ( .A1(n7568), .A2(n10388), .B1(n7940), .B2(n10375), .ZN(n7561) );
  AOI21_X1 U8939 ( .B1(n7562), .B2(n10411), .A(n7561), .ZN(n7563) );
  OAI21_X1 U8940 ( .B1(n7566), .B2(n11084), .A(n7563), .ZN(n11045) );
  NAND2_X1 U8941 ( .A1(n11045), .A2(n10307), .ZN(n7564) );
  OAI211_X1 U8942 ( .C1(n7566), .C2(n7577), .A(n7565), .B(n7564), .ZN(P1_U3290) );
  OAI21_X1 U8943 ( .B1(n5416), .B2(n5140), .A(n7567), .ZN(n7576) );
  OAI22_X1 U8944 ( .A1(n7569), .A2(n10388), .B1(n7568), .B2(n10375), .ZN(n7575) );
  OAI21_X1 U8945 ( .B1(n7572), .B2(n7571), .A(n7570), .ZN(n11038) );
  INV_X1 U8946 ( .A(n11038), .ZN(n7573) );
  NOR2_X1 U8947 ( .A1(n7573), .A2(n11084), .ZN(n7574) );
  AOI211_X1 U8948 ( .C1(n10411), .C2(n7576), .A(n7575), .B(n7574), .ZN(n11035)
         );
  INV_X1 U8949 ( .A(n7577), .ZN(n7737) );
  OAI211_X1 U8950 ( .C1(n11034), .C2(n9725), .A(n10400), .B(n7693), .ZN(n11033) );
  NOR2_X1 U8951 ( .A1(n10219), .A2(n11033), .ZN(n7580) );
  INV_X2 U8952 ( .A(n7919), .ZN(n11067) );
  AOI22_X1 U8953 ( .A1(n11079), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n11067), .ZN(n7578) );
  OAI21_X1 U8954 ( .B1(n11072), .B2(n11034), .A(n7578), .ZN(n7579) );
  AOI211_X1 U8955 ( .C1(n7737), .C2(n11038), .A(n7580), .B(n7579), .ZN(n7581)
         );
  OAI21_X1 U8956 ( .B1(n11079), .B2(n11035), .A(n7581), .ZN(P1_U3292) );
  NAND2_X1 U8957 ( .A1(n7583), .A2(n7582), .ZN(n7584) );
  NAND2_X1 U8958 ( .A1(n7584), .A2(n7585), .ZN(n7588) );
  OR2_X1 U8959 ( .A1(n7586), .A2(n7585), .ZN(n7587) );
  OAI21_X1 U8960 ( .B1(n9380), .B2(n10562), .A(n7591), .ZN(n7598) );
  INV_X1 U8961 ( .A(n7592), .ZN(n7594) );
  INV_X1 U8962 ( .A(n8509), .ZN(n9216) );
  OAI22_X1 U8963 ( .A1(n9317), .A2(n7593), .B1(n9377), .B2(n7177), .ZN(n7597)
         );
  AND3_X1 U8964 ( .A1(n8885), .A2(n7595), .A3(n7594), .ZN(n7596) );
  AOI211_X1 U8965 ( .C1(n9377), .C2(n7598), .A(n7597), .B(n7596), .ZN(n7599)
         );
  INV_X1 U8966 ( .A(n7599), .ZN(P2_U3233) );
  OR2_X1 U8967 ( .A1(n11079), .A2(n10375), .ZN(n10287) );
  NOR2_X1 U8968 ( .A1(n7919), .A2(n7600), .ZN(n7604) );
  INV_X1 U8969 ( .A(n7601), .ZN(n11025) );
  XNOR2_X1 U8970 ( .A(n10005), .B(n11024), .ZN(n11021) );
  NOR4_X1 U8971 ( .A1(n11069), .A2(n7602), .A3(n11025), .A4(n11021), .ZN(n7603) );
  AOI211_X1 U8972 ( .C1(n11079), .C2(P1_REG2_REG_0__SCAN_IN), .A(n7604), .B(
        n7603), .ZN(n7606) );
  NOR2_X1 U8973 ( .A1(n10219), .A2(n10300), .ZN(n10128) );
  OAI21_X1 U8974 ( .B1(n10128), .B2(n10223), .A(n11024), .ZN(n7605) );
  OAI211_X1 U8975 ( .C1(n5968), .C2(n10287), .A(n7606), .B(n7605), .ZN(
        P1_U3293) );
  INV_X1 U8976 ( .A(n7607), .ZN(n7608) );
  INV_X1 U8977 ( .A(n10080), .ZN(n8431) );
  OAI222_X1 U8978 ( .A1(n8627), .A2(n10785), .B1(n8633), .B2(n7608), .C1(
        P1_U3086), .C2(n8431), .ZN(P1_U3339) );
  OAI222_X1 U8979 ( .A1(n9513), .A2(n7609), .B1(n8667), .B2(n7608), .C1(
        P2_U3151), .C2(n9118), .ZN(P2_U3279) );
  INV_X1 U8980 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7611) );
  NAND2_X1 U8981 ( .A1(n10866), .A2(n7819), .ZN(n7610) );
  NAND2_X1 U8982 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9652) );
  OAI211_X1 U8983 ( .C1(n7611), .C2(n10869), .A(n7610), .B(n9652), .ZN(n7623)
         );
  AOI21_X1 U8984 ( .B1(n7617), .B2(P1_REG1_REG_10__SCAN_IN), .A(n7612), .ZN(
        n7615) );
  NAND2_X1 U8985 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n7819), .ZN(n7613) );
  OAI21_X1 U8986 ( .B1(n7819), .B2(P1_REG1_REG_11__SCAN_IN), .A(n7613), .ZN(
        n7614) );
  NOR2_X1 U8987 ( .A1(n7615), .A2(n7614), .ZN(n7818) );
  AOI211_X1 U8988 ( .C1(n7615), .C2(n7614), .A(n7818), .B(n10125), .ZN(n7622)
         );
  AOI21_X1 U8989 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n7617), .A(n7616), .ZN(
        n7620) );
  NAND2_X1 U8990 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n7819), .ZN(n7618) );
  OAI21_X1 U8991 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n7819), .A(n7618), .ZN(
        n7619) );
  NOR2_X1 U8992 ( .A1(n7620), .A2(n7619), .ZN(n7817) );
  AOI211_X1 U8993 ( .C1(n7620), .C2(n7619), .A(n7817), .B(n8444), .ZN(n7621)
         );
  OR3_X1 U8994 ( .A1(n7623), .A2(n7622), .A3(n7621), .ZN(P1_U3254) );
  INV_X1 U8995 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n8212) );
  INV_X1 U8996 ( .A(n7867), .ZN(n7626) );
  AOI21_X1 U8997 ( .B1(n8212), .B2(n7627), .A(n7853), .ZN(n7645) );
  INV_X1 U8998 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7628) );
  MUX2_X1 U8999 ( .A(n7628), .B(n8212), .S(n8174), .Z(n7630) );
  AND2_X1 U9000 ( .A1(n7630), .A2(n7867), .ZN(n7861) );
  INV_X1 U9001 ( .A(n7861), .ZN(n7629) );
  OAI21_X1 U9002 ( .B1(n7867), .B2(n7630), .A(n7629), .ZN(n7634) );
  NOR2_X1 U9003 ( .A1(n7633), .A2(n7634), .ZN(n7860) );
  AOI21_X1 U9004 ( .B1(n7634), .B2(n7633), .A(n7860), .ZN(n7636) );
  AND2_X1 U9005 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7900) );
  AOI21_X1 U9006 ( .B1(n10996), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n7900), .ZN(
        n7635) );
  OAI21_X1 U9007 ( .B1(n7636), .B2(n9164), .A(n7635), .ZN(n7643) );
  AOI21_X1 U9008 ( .B1(n7628), .B2(n7640), .A(n7868), .ZN(n7641) );
  NOR2_X1 U9009 ( .A1(n7641), .A2(n11014), .ZN(n7642) );
  AOI211_X1 U9010 ( .C1(n10997), .C2(n7867), .A(n7643), .B(n7642), .ZN(n7644)
         );
  OAI21_X1 U9011 ( .B1(n7645), .B2(n11005), .A(n7644), .ZN(P2_U3189) );
  INV_X1 U9012 ( .A(n8831), .ZN(n7655) );
  AOI211_X1 U9013 ( .C1(n7648), .C2(n7647), .A(n8788), .B(n7646), .ZN(n7649)
         );
  INV_X1 U9014 ( .A(n7649), .ZN(n7654) );
  INV_X1 U9015 ( .A(n7650), .ZN(n7652) );
  OAI22_X1 U9016 ( .A1(n7798), .A2(n8829), .B1(n7970), .B2(n8835), .ZN(n7651)
         );
  AOI211_X1 U9017 ( .C1(n8827), .C2(n9050), .A(n7652), .B(n7651), .ZN(n7653)
         );
  OAI211_X1 U9018 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n7655), .A(n7654), .B(
        n7653), .ZN(P2_U3158) );
  OAI21_X1 U9019 ( .B1(n7657), .B2(n9843), .A(n7656), .ZN(n11076) );
  AOI211_X1 U9020 ( .C1(n8022), .C2(n7944), .A(n10300), .B(n7714), .ZN(n11066)
         );
  XNOR2_X1 U9021 ( .A(n7658), .B(n9843), .ZN(n7659) );
  AOI222_X1 U9022 ( .A1(n10411), .A2(n7659), .B1(n9999), .B2(n11088), .C1(
        n10001), .C2(n11089), .ZN(n11078) );
  INV_X1 U9023 ( .A(n11078), .ZN(n7660) );
  AOI211_X1 U9024 ( .C1(n11107), .C2(n11076), .A(n11066), .B(n7660), .ZN(n8069) );
  INV_X1 U9025 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7661) );
  OAI22_X1 U9026 ( .A1(n10457), .A2(n11073), .B1(n11114), .B2(n7661), .ZN(
        n7662) );
  INV_X1 U9027 ( .A(n7662), .ZN(n7663) );
  OAI21_X1 U9028 ( .B1(n8069), .B2(n11111), .A(n7663), .ZN(P1_U3471) );
  NAND2_X1 U9029 ( .A1(n9045), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7664) );
  OAI21_X1 U9030 ( .B1(n8844), .B2(n9045), .A(n7664), .ZN(P2_U3521) );
  XNOR2_X1 U9031 ( .A(n8012), .B(n8694), .ZN(n7778) );
  XNOR2_X1 U9032 ( .A(n9047), .B(n7778), .ZN(n7669) );
  INV_X1 U9033 ( .A(n7665), .ZN(n7666) );
  NAND2_X1 U9034 ( .A1(n7667), .A2(n7666), .ZN(n7668) );
  NAND2_X1 U9035 ( .A1(n7668), .A2(n7669), .ZN(n7780) );
  OAI21_X1 U9036 ( .B1(n7669), .B2(n7668), .A(n7780), .ZN(n7676) );
  AND2_X1 U9037 ( .A1(n7806), .A2(n8786), .ZN(n7675) );
  INV_X1 U9038 ( .A(n7670), .ZN(n7671) );
  AOI21_X1 U9039 ( .B1(n9048), .B2(n8827), .A(n7671), .ZN(n7673) );
  NAND2_X1 U9040 ( .A1(n8831), .A2(n7802), .ZN(n7672) );
  OAI211_X1 U9041 ( .C1(n8150), .C2(n8829), .A(n7673), .B(n7672), .ZN(n7674)
         );
  AOI211_X1 U9042 ( .C1(n7676), .C2(n8824), .A(n7675), .B(n7674), .ZN(n7677)
         );
  INV_X1 U9043 ( .A(n7677), .ZN(P2_U3167) );
  NAND2_X1 U9044 ( .A1(n9045), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7678) );
  OAI21_X1 U9045 ( .B1(n9179), .B2(n9045), .A(n7678), .ZN(P2_U3520) );
  OAI21_X1 U9046 ( .B1(n7680), .B2(n9775), .A(n7679), .ZN(n7927) );
  INV_X1 U9047 ( .A(n7927), .ZN(n7685) );
  OAI21_X1 U9048 ( .B1(n7682), .B2(n7681), .A(n7937), .ZN(n7683) );
  AOI222_X1 U9049 ( .A1(n10411), .A2(n7683), .B1(n10001), .B2(n11088), .C1(
        n10003), .C2(n11089), .ZN(n7929) );
  OAI211_X1 U9050 ( .C1(n7684), .C2(n6009), .A(n7943), .B(n10400), .ZN(n7925)
         );
  OAI211_X1 U9051 ( .C1(n11023), .C2(n7685), .A(n7929), .B(n7925), .ZN(n8072)
         );
  INV_X1 U9052 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7686) );
  OAI22_X1 U9053 ( .A1(n10457), .A2(n6009), .B1(n11114), .B2(n7686), .ZN(n7687) );
  AOI21_X1 U9054 ( .B1(n8072), .B2(n11114), .A(n7687), .ZN(n7688) );
  INV_X1 U9055 ( .A(n7688), .ZN(P1_U3465) );
  OAI21_X1 U9056 ( .B1(n7691), .B2(n7689), .A(n7690), .ZN(n7934) );
  AOI211_X1 U9057 ( .C1(n7694), .C2(n7693), .A(n10300), .B(n7692), .ZN(n7930)
         );
  XOR2_X1 U9058 ( .A(n7689), .B(n9832), .Z(n7695) );
  AOI222_X1 U9059 ( .A1(n10411), .A2(n7695), .B1(n10003), .B2(n11088), .C1(
        n6332), .C2(n11089), .ZN(n7936) );
  INV_X1 U9060 ( .A(n7936), .ZN(n7696) );
  AOI211_X1 U9061 ( .C1(n11107), .C2(n7934), .A(n7930), .B(n7696), .ZN(n8077)
         );
  INV_X1 U9062 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n7697) );
  OAI22_X1 U9063 ( .A1(n10457), .A2(n8074), .B1(n11114), .B2(n7697), .ZN(n7698) );
  INV_X1 U9064 ( .A(n7698), .ZN(n7699) );
  OAI21_X1 U9065 ( .B1(n8077), .B2(n11111), .A(n7699), .ZN(P1_U3459) );
  OAI21_X1 U9066 ( .B1(n7701), .B2(n7703), .A(n7700), .ZN(n7742) );
  NAND2_X1 U9067 ( .A1(n7711), .A2(n5695), .ZN(n7725) );
  INV_X1 U9068 ( .A(n7724), .ZN(n7702) );
  NOR2_X1 U9069 ( .A1(n9858), .A2(n7702), .ZN(n9862) );
  NAND2_X1 U9070 ( .A1(n7725), .A2(n9862), .ZN(n7726) );
  NAND2_X1 U9071 ( .A1(n7726), .A2(n9883), .ZN(n7704) );
  XNOR2_X1 U9072 ( .A(n7704), .B(n7703), .ZN(n7750) );
  NAND2_X1 U9073 ( .A1(n7750), .A2(n10411), .ZN(n7706) );
  AOI21_X1 U9074 ( .B1(n7732), .B2(n8299), .A(n10300), .ZN(n7705) );
  AOI22_X1 U9075 ( .A1(n7705), .A2(n7881), .B1(n11088), .B2(n11090), .ZN(n7748) );
  OAI211_X1 U9076 ( .C1(n7962), .C2(n10388), .A(n7706), .B(n7748), .ZN(n7707)
         );
  AOI21_X1 U9077 ( .B1(n7742), .B2(n11107), .A(n7707), .ZN(n8066) );
  INV_X1 U9078 ( .A(n8299), .ZN(n8063) );
  INV_X1 U9079 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n7708) );
  OAI22_X1 U9080 ( .A1(n10457), .A2(n8063), .B1(n11114), .B2(n7708), .ZN(n7709) );
  INV_X1 U9081 ( .A(n7709), .ZN(n7710) );
  OAI21_X1 U9082 ( .B1(n8066), .B2(n11111), .A(n7710), .ZN(P1_U3480) );
  XNOR2_X1 U9083 ( .A(n7711), .B(n9852), .ZN(n7968) );
  OAI21_X1 U9084 ( .B1(n7713), .B2(n9852), .A(n7712), .ZN(n7959) );
  INV_X1 U9085 ( .A(n7714), .ZN(n7715) );
  AOI211_X1 U9086 ( .C1(n7716), .C2(n7715), .A(n10300), .B(n7733), .ZN(n7965)
         );
  OAI22_X1 U9087 ( .A1(n8141), .A2(n10388), .B1(n7962), .B2(n10375), .ZN(n7717) );
  AOI211_X1 U9088 ( .C1(n7959), .C2(n11107), .A(n7965), .B(n7717), .ZN(n7718)
         );
  OAI21_X1 U9089 ( .B1(n11022), .B2(n7968), .A(n7718), .ZN(n8080) );
  INV_X1 U9090 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7719) );
  OAI22_X1 U9091 ( .A1(n10457), .A2(n8147), .B1(n11114), .B2(n7719), .ZN(n7720) );
  AOI21_X1 U9092 ( .B1(n8080), .B2(n11114), .A(n7720), .ZN(n7721) );
  INV_X1 U9093 ( .A(n7721), .ZN(P1_U3474) );
  INV_X1 U9094 ( .A(n11084), .ZN(n7731) );
  OAI21_X1 U9095 ( .B1(n7723), .B2(n9858), .A(n7722), .ZN(n7827) );
  OAI22_X1 U9096 ( .A1(n8235), .A2(n10388), .B1(n9545), .B2(n10375), .ZN(n7730) );
  NAND2_X1 U9097 ( .A1(n7725), .A2(n7724), .ZN(n7728) );
  INV_X1 U9098 ( .A(n7726), .ZN(n7727) );
  AOI211_X1 U9099 ( .C1(n9858), .C2(n7728), .A(n11022), .B(n7727), .ZN(n7729)
         );
  AOI211_X1 U9100 ( .C1(n7731), .C2(n7827), .A(n7730), .B(n7729), .ZN(n7829)
         );
  OAI211_X1 U9101 ( .C1(n7733), .C2(n8083), .A(n10400), .B(n7732), .ZN(n7828)
         );
  AOI22_X1 U9102 ( .A1(n11069), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n8234), .B2(
        n11067), .ZN(n7735) );
  NAND2_X1 U9103 ( .A1(n10223), .A2(n8239), .ZN(n7734) );
  OAI211_X1 U9104 ( .C1(n7828), .C2(n10219), .A(n7735), .B(n7734), .ZN(n7736)
         );
  AOI21_X1 U9105 ( .B1(n7827), .B2(n7737), .A(n7736), .ZN(n7738) );
  OAI21_X1 U9106 ( .B1(n7829), .B2(n11069), .A(n7738), .ZN(P1_U3285) );
  INV_X1 U9107 ( .A(n7739), .ZN(n7741) );
  INV_X1 U9108 ( .A(n9138), .ZN(n8553) );
  OAI222_X1 U9109 ( .A1(n8667), .A2(n7741), .B1(n8553), .B2(P2_U3151), .C1(
        n7740), .C2(n9513), .ZN(P2_U3278) );
  INV_X1 U9110 ( .A(n10078), .ZN(n10099) );
  OAI222_X1 U9111 ( .A1(P1_U3086), .A2(n10099), .B1(n8633), .B2(n7741), .C1(
        n10789), .C2(n10471), .ZN(P1_U3338) );
  INV_X1 U9112 ( .A(n7742), .ZN(n7752) );
  AND2_X1 U9113 ( .A1(n7743), .A2(n11084), .ZN(n7744) );
  OR2_X1 U9114 ( .A1(n11079), .A2(n11022), .ZN(n10292) );
  INV_X1 U9115 ( .A(n10292), .ZN(n10164) );
  OR2_X1 U9116 ( .A1(n11079), .A2(n10388), .ZN(n10143) );
  AOI22_X1 U9117 ( .A1(n11069), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n8296), .B2(
        n11067), .ZN(n7745) );
  OAI21_X1 U9118 ( .B1(n10143), .B2(n7962), .A(n7745), .ZN(n7746) );
  AOI21_X1 U9119 ( .B1(n10223), .B2(n8299), .A(n7746), .ZN(n7747) );
  OAI21_X1 U9120 ( .B1(n7748), .B2(n10219), .A(n7747), .ZN(n7749) );
  AOI21_X1 U9121 ( .B1(n7750), .B2(n10164), .A(n7749), .ZN(n7751) );
  OAI21_X1 U9122 ( .B1(n7752), .B2(n10309), .A(n7751), .ZN(P1_U3284) );
  AOI211_X1 U9123 ( .C1(n5626), .C2(n7754), .A(n9697), .B(n7753), .ZN(n7759)
         );
  INV_X1 U9124 ( .A(n7755), .ZN(n7920) );
  AOI22_X1 U9125 ( .A1(n9678), .A2(n10003), .B1(n9687), .B2(n10001), .ZN(n7757) );
  AND2_X1 U9126 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n10024) );
  AOI21_X1 U9127 ( .B1(n9694), .B2(n7923), .A(n10024), .ZN(n7756) );
  OAI211_X1 U9128 ( .C1(n7920), .C2(n9646), .A(n7757), .B(n7756), .ZN(n7758)
         );
  OR2_X1 U9129 ( .A1(n7759), .A2(n7758), .ZN(P1_U3230) );
  INV_X1 U9130 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10094) );
  INV_X1 U9131 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8575) );
  AOI22_X1 U9132 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(P1_ADDR_REG_18__SCAN_IN), 
        .B1(n10094), .B2(n8575), .ZN(n10935) );
  NOR2_X1 U9133 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7760) );
  AOI21_X1 U9134 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7760), .ZN(n10932) );
  NOR2_X1 U9135 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7761) );
  AOI21_X1 U9136 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7761), .ZN(n10929) );
  INV_X1 U9137 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n9094) );
  INV_X1 U9138 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10870) );
  AOI22_X1 U9139 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(P2_ADDR_REG_15__SCAN_IN), 
        .B1(n9094), .B2(n10870), .ZN(n10926) );
  NOR2_X1 U9140 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7762) );
  AOI21_X1 U9141 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7762), .ZN(n10923) );
  NOR2_X1 U9142 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7763) );
  AOI21_X1 U9143 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7763), .ZN(n10920) );
  NOR2_X1 U9144 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7764) );
  AOI21_X1 U9145 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7764), .ZN(n10917) );
  NOR2_X1 U9146 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7765) );
  AOI21_X1 U9147 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7765), .ZN(n10914) );
  NOR2_X1 U9148 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7766) );
  AOI21_X1 U9149 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7766), .ZN(n10911) );
  NOR2_X1 U9150 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7767) );
  AOI21_X1 U9151 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7767), .ZN(n10908) );
  NOR2_X1 U9152 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7768) );
  AOI21_X1 U9153 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7768), .ZN(n10905) );
  NOR2_X1 U9154 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7769) );
  AOI21_X1 U9155 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7769), .ZN(n10902) );
  NOR2_X1 U9156 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7770) );
  AOI21_X1 U9157 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n7770), .ZN(n10899) );
  NOR2_X1 U9158 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7771) );
  AOI21_X1 U9159 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n7771), .ZN(n10896) );
  AND2_X1 U9160 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .ZN(n7772) );
  NOR2_X1 U9161 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7772), .ZN(n10881) );
  INV_X1 U9162 ( .A(n10881), .ZN(n10882) );
  INV_X1 U9163 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10884) );
  NAND3_X1 U9164 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_0__SCAN_IN), .ZN(n10883) );
  NAND2_X1 U9165 ( .A1(n10884), .A2(n10883), .ZN(n10880) );
  NAND2_X1 U9166 ( .A1(n10882), .A2(n10880), .ZN(n10887) );
  NAND2_X1 U9167 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7773) );
  OAI21_X1 U9168 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7773), .ZN(n10886) );
  NOR2_X1 U9169 ( .A1(n10887), .A2(n10886), .ZN(n10885) );
  AOI21_X1 U9170 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10885), .ZN(n10890) );
  NAND2_X1 U9171 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n7774) );
  OAI21_X1 U9172 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n7774), .ZN(n10889) );
  NOR2_X1 U9173 ( .A1(n10890), .A2(n10889), .ZN(n10888) );
  AOI21_X1 U9174 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n10888), .ZN(n10893) );
  NOR2_X1 U9175 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7775) );
  AOI21_X1 U9176 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7775), .ZN(n10892) );
  NAND2_X1 U9177 ( .A1(n10893), .A2(n10892), .ZN(n10891) );
  OAI21_X1 U9178 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10891), .ZN(n10895) );
  NAND2_X1 U9179 ( .A1(n10896), .A2(n10895), .ZN(n10894) );
  OAI21_X1 U9180 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10894), .ZN(n10898) );
  NAND2_X1 U9181 ( .A1(n10899), .A2(n10898), .ZN(n10897) );
  OAI21_X1 U9182 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10897), .ZN(n10901) );
  NAND2_X1 U9183 ( .A1(n10902), .A2(n10901), .ZN(n10900) );
  OAI21_X1 U9184 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10900), .ZN(n10904) );
  NAND2_X1 U9185 ( .A1(n10905), .A2(n10904), .ZN(n10903) );
  OAI21_X1 U9186 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10903), .ZN(n10907) );
  NAND2_X1 U9187 ( .A1(n10908), .A2(n10907), .ZN(n10906) );
  OAI21_X1 U9188 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10906), .ZN(n10910) );
  NAND2_X1 U9189 ( .A1(n10911), .A2(n10910), .ZN(n10909) );
  OAI21_X1 U9190 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10909), .ZN(n10913) );
  NAND2_X1 U9191 ( .A1(n10914), .A2(n10913), .ZN(n10912) );
  OAI21_X1 U9192 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10912), .ZN(n10916) );
  NAND2_X1 U9193 ( .A1(n10917), .A2(n10916), .ZN(n10915) );
  OAI21_X1 U9194 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10915), .ZN(n10919) );
  NAND2_X1 U9195 ( .A1(n10920), .A2(n10919), .ZN(n10918) );
  OAI21_X1 U9196 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10918), .ZN(n10922) );
  NAND2_X1 U9197 ( .A1(n10923), .A2(n10922), .ZN(n10921) );
  OAI21_X1 U9198 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10921), .ZN(n10925) );
  NAND2_X1 U9199 ( .A1(n10926), .A2(n10925), .ZN(n10924) );
  OAI21_X1 U9200 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n10924), .ZN(n10928) );
  NAND2_X1 U9201 ( .A1(n10929), .A2(n10928), .ZN(n10927) );
  OAI21_X1 U9202 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10927), .ZN(n10931) );
  NAND2_X1 U9203 ( .A1(n10932), .A2(n10931), .ZN(n10930) );
  OAI21_X1 U9204 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10930), .ZN(n10934) );
  NAND2_X1 U9205 ( .A1(n10935), .A2(n10934), .ZN(n10933) );
  OAI21_X1 U9206 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(P1_ADDR_REG_18__SCAN_IN), 
        .A(n10933), .ZN(n7777) );
  XNOR2_X1 U9207 ( .A(n5679), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n7776) );
  XNOR2_X1 U9208 ( .A(n7777), .B(n7776), .ZN(ADD_1068_U4) );
  XNOR2_X1 U9209 ( .A(n8160), .B(n8678), .ZN(n7893) );
  XNOR2_X1 U9210 ( .A(n7893), .B(n8150), .ZN(n7781) );
  NAND2_X1 U9211 ( .A1(n8127), .A2(n7778), .ZN(n7782) );
  INV_X1 U9212 ( .A(n7895), .ZN(n7784) );
  AOI21_X1 U9213 ( .B1(n7780), .B2(n7782), .A(n7781), .ZN(n7783) );
  NOR3_X1 U9214 ( .A1(n7784), .A2(n7783), .A3(n8788), .ZN(n7792) );
  INV_X1 U9215 ( .A(n7785), .ZN(n7786) );
  AOI21_X1 U9216 ( .B1(n9047), .B2(n8827), .A(n7786), .ZN(n7790) );
  NAND2_X1 U9217 ( .A1(n8130), .A2(n8786), .ZN(n7789) );
  NAND2_X1 U9218 ( .A1(n8831), .A2(n8129), .ZN(n7788) );
  NAND2_X1 U9219 ( .A1(n9046), .A2(n8815), .ZN(n7787) );
  NAND4_X1 U9220 ( .A1(n7790), .A2(n7789), .A3(n7788), .A4(n7787), .ZN(n7791)
         );
  OR2_X1 U9221 ( .A1(n7792), .A2(n7791), .ZN(P2_U3179) );
  INV_X1 U9222 ( .A(n10096), .ZN(n10098) );
  INV_X1 U9223 ( .A(n7793), .ZN(n7825) );
  OAI222_X1 U9224 ( .A1(P1_U3086), .A2(n10098), .B1(n8633), .B2(n7825), .C1(
        n7794), .C2(n10471), .ZN(P1_U3337) );
  OAI21_X1 U9225 ( .B1(n7795), .B2(n8852), .A(n8122), .ZN(n8015) );
  INV_X1 U9226 ( .A(n8015), .ZN(n7809) );
  AND2_X1 U9227 ( .A1(n7796), .A2(n7476), .ZN(n7797) );
  NAND2_X1 U9228 ( .A1(n9377), .A2(n7797), .ZN(n8620) );
  XNOR2_X1 U9229 ( .A(n5216), .B(n8852), .ZN(n7801) );
  OAI22_X1 U9230 ( .A1(n7798), .A2(n9361), .B1(n8150), .B2(n9376), .ZN(n7799)
         );
  AOI21_X1 U9231 ( .B1(n8015), .B2(n8385), .A(n7799), .ZN(n7800) );
  OAI21_X1 U9232 ( .B1(n7801), .B2(n9373), .A(n7800), .ZN(n8013) );
  NAND2_X1 U9233 ( .A1(n8013), .A2(n9377), .ZN(n7808) );
  INV_X1 U9234 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7804) );
  INV_X1 U9235 ( .A(n7802), .ZN(n7803) );
  OAI22_X1 U9236 ( .A1(n9377), .A2(n7804), .B1(n7803), .B2(n9380), .ZN(n7805)
         );
  AOI21_X1 U9237 ( .B1(n9364), .B2(n7806), .A(n7805), .ZN(n7807) );
  OAI211_X1 U9238 ( .C1(n7809), .C2(n8620), .A(n7808), .B(n7807), .ZN(P2_U3228) );
  NAND2_X1 U9239 ( .A1(n7810), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7814) );
  NAND2_X1 U9240 ( .A1(n7811), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n7813) );
  NAND2_X1 U9241 ( .A1(n6839), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n7812) );
  NAND4_X1 U9242 ( .A1(n7815), .A2(n7814), .A3(n7813), .A4(n7812), .ZN(n9172)
         );
  NAND2_X1 U9243 ( .A1(n9172), .A2(P2_U3893), .ZN(n7816) );
  OAI21_X1 U9244 ( .B1(P2_U3893), .B2(n10472), .A(n7816), .ZN(P2_U3522) );
  XNOR2_X1 U9245 ( .A(n8434), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n8436) );
  AOI21_X1 U9246 ( .B1(n7819), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7817), .ZN(
        n8435) );
  XNOR2_X1 U9247 ( .A(n8436), .B(n8435), .ZN(n7821) );
  XNOR2_X1 U9248 ( .A(n8434), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n8421) );
  AOI21_X1 U9249 ( .B1(n7819), .B2(P1_REG1_REG_11__SCAN_IN), .A(n7818), .ZN(
        n8420) );
  XNOR2_X1 U9250 ( .A(n8421), .B(n8420), .ZN(n7820) );
  AOI22_X1 U9251 ( .A1(n10871), .A2(n7821), .B1(n10877), .B2(n7820), .ZN(n7824) );
  INV_X1 U9252 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7822) );
  NOR2_X1 U9253 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7822), .ZN(n9574) );
  AOI21_X1 U9254 ( .B1(n10119), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n9574), .ZN(
        n7823) );
  OAI211_X1 U9255 ( .C1(n8434), .C2(n10121), .A(n7824), .B(n7823), .ZN(
        P1_U3255) );
  INV_X1 U9256 ( .A(n9157), .ZN(n8587) );
  OAI222_X1 U9257 ( .A1(n9513), .A2(n7826), .B1(n8587), .B2(P2_U3151), .C1(
        n8667), .C2(n7825), .ZN(P2_U3277) );
  INV_X1 U9258 ( .A(n7827), .ZN(n7830) );
  OAI211_X1 U9259 ( .C1(n7830), .C2(n11085), .A(n7829), .B(n7828), .ZN(n8085)
         );
  INV_X1 U9260 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7831) );
  OAI22_X1 U9261 ( .A1(n10457), .A2(n8083), .B1(n11114), .B2(n7831), .ZN(n7832) );
  AOI21_X1 U9262 ( .B1(n8085), .B2(n11114), .A(n7832), .ZN(n7833) );
  INV_X1 U9263 ( .A(n7833), .ZN(P1_U3477) );
  OAI21_X1 U9264 ( .B1(n7835), .B2(n8897), .A(n7834), .ZN(n8036) );
  NOR2_X1 U9265 ( .A1(n7836), .A2(n9450), .ZN(n7842) );
  AOI211_X1 U9266 ( .C1(n8897), .C2(n7838), .A(n9373), .B(n7837), .ZN(n7841)
         );
  OAI22_X1 U9267 ( .A1(n8127), .A2(n9376), .B1(n7839), .B2(n9361), .ZN(n7840)
         );
  OR2_X1 U9268 ( .A1(n7841), .A2(n7840), .ZN(n8037) );
  AOI211_X1 U9269 ( .C1(n9414), .C2(n8036), .A(n7842), .B(n8037), .ZN(n11052)
         );
  OR2_X1 U9270 ( .A1(n11052), .A2(n9465), .ZN(n7843) );
  OAI21_X1 U9271 ( .B1(n9456), .B2(n7844), .A(n7843), .ZN(P2_U3463) );
  INV_X1 U9272 ( .A(n7845), .ZN(n7849) );
  OAI222_X1 U9273 ( .A1(n8667), .A2(n7849), .B1(n9513), .B2(n6694), .C1(
        P2_U3151), .C2(n6847), .ZN(P2_U3275) );
  INV_X1 U9274 ( .A(n7846), .ZN(n8722) );
  OAI222_X1 U9275 ( .A1(n9513), .A2(n7847), .B1(n8667), .B2(n8722), .C1(
        P2_U3151), .C2(n5535), .ZN(P2_U3276) );
  OAI222_X1 U9276 ( .A1(n8627), .A2(n7850), .B1(n8633), .B2(n7849), .C1(n7848), 
        .C2(P1_U3086), .ZN(P1_U3335) );
  NAND2_X1 U9277 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n7997), .ZN(n7854) );
  OAI21_X1 U9278 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n7997), .A(n7854), .ZN(
        n7855) );
  AOI21_X1 U9279 ( .B1(n7856), .B2(n7855), .A(n7993), .ZN(n7878) );
  INV_X1 U9280 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n8249) );
  INV_X1 U9281 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7857) );
  MUX2_X1 U9282 ( .A(n8249), .B(n7857), .S(n8174), .Z(n7859) );
  AND2_X1 U9283 ( .A1(n7859), .A2(n7876), .ZN(n8002) );
  INV_X1 U9284 ( .A(n8002), .ZN(n7858) );
  OAI21_X1 U9285 ( .B1(n7876), .B2(n7859), .A(n7858), .ZN(n7863) );
  NOR2_X1 U9286 ( .A1(n7861), .A2(n7860), .ZN(n7862) );
  NOR2_X1 U9287 ( .A1(n7862), .A2(n7863), .ZN(n8001) );
  AOI21_X1 U9288 ( .B1(n7863), .B2(n7862), .A(n8001), .ZN(n7865) );
  AND2_X1 U9289 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3151), .ZN(n8053) );
  AOI21_X1 U9290 ( .B1(n10996), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n8053), .ZN(
        n7864) );
  OAI21_X1 U9291 ( .B1(n7865), .B2(n9164), .A(n7864), .ZN(n7875) );
  NOR2_X1 U9292 ( .A1(n7867), .A2(n7866), .ZN(n7869) );
  NAND2_X1 U9293 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n7997), .ZN(n7870) );
  OAI21_X1 U9294 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n7997), .A(n7870), .ZN(
        n7871) );
  NOR2_X1 U9295 ( .A1(n7872), .A2(n7871), .ZN(n7996) );
  AOI21_X1 U9296 ( .B1(n7872), .B2(n7871), .A(n7996), .ZN(n7873) );
  NOR2_X1 U9297 ( .A1(n7873), .A2(n11014), .ZN(n7874) );
  AOI211_X1 U9298 ( .C1(n10997), .C2(n7876), .A(n7875), .B(n7874), .ZN(n7877)
         );
  OAI21_X1 U9299 ( .B1(n7878), .B2(n11005), .A(n7877), .ZN(P2_U3190) );
  OAI21_X1 U9300 ( .B1(n7880), .B2(n9781), .A(n7879), .ZN(n7952) );
  AOI211_X1 U9301 ( .C1(n9547), .C2(n7881), .A(n10300), .B(n7910), .ZN(n7955)
         );
  OAI21_X1 U9302 ( .B1(n7884), .B2(n7883), .A(n7882), .ZN(n7885) );
  AOI222_X1 U9303 ( .A1(n10411), .A2(n7885), .B1(n9996), .B2(n11088), .C1(
        n9997), .C2(n11089), .ZN(n7958) );
  INV_X1 U9304 ( .A(n7958), .ZN(n7886) );
  AOI211_X1 U9305 ( .C1(n7952), .C2(n11107), .A(n7955), .B(n7886), .ZN(n8045)
         );
  INV_X1 U9306 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7887) );
  OAI22_X1 U9307 ( .A1(n10457), .A2(n5700), .B1(n11114), .B2(n7887), .ZN(n7888) );
  INV_X1 U9308 ( .A(n7888), .ZN(n7889) );
  OAI21_X1 U9309 ( .B1(n8045), .B2(n11111), .A(n7889), .ZN(P1_U3483) );
  INV_X1 U9310 ( .A(n7890), .ZN(n8626) );
  OAI222_X1 U9311 ( .A1(n8667), .A2(n8626), .B1(n7892), .B2(P2_U3151), .C1(
        n7891), .C2(n9513), .ZN(P2_U3274) );
  XNOR2_X1 U9312 ( .A(n8931), .B(n8694), .ZN(n8046) );
  XNOR2_X1 U9313 ( .A(n8046), .B(n8047), .ZN(n7899) );
  INV_X1 U9314 ( .A(n7893), .ZN(n7894) );
  INV_X1 U9315 ( .A(n7899), .ZN(n7896) );
  INV_X1 U9316 ( .A(n8049), .ZN(n7897) );
  AOI21_X1 U9317 ( .B1(n7899), .B2(n7898), .A(n7897), .ZN(n7906) );
  INV_X1 U9318 ( .A(n8931), .ZN(n7904) );
  AOI21_X1 U9319 ( .B1(n6520), .B2(n8827), .A(n7900), .ZN(n7902) );
  NAND2_X1 U9320 ( .A1(n8831), .A2(n8155), .ZN(n7901) );
  OAI211_X1 U9321 ( .C1(n8151), .C2(n8829), .A(n7902), .B(n7901), .ZN(n7903)
         );
  AOI21_X1 U9322 ( .B1(n7904), .B2(n8786), .A(n7903), .ZN(n7905) );
  OAI21_X1 U9323 ( .B1(n7906), .B2(n8788), .A(n7905), .ZN(P2_U3153) );
  XNOR2_X1 U9324 ( .A(n7907), .B(n9783), .ZN(n11086) );
  XOR2_X1 U9325 ( .A(n9783), .B(n7908), .Z(n7909) );
  NOR2_X1 U9326 ( .A1(n7909), .A2(n11022), .ZN(n11094) );
  OAI21_X1 U9327 ( .B1(n7910), .B2(n5698), .A(n10400), .ZN(n7911) );
  OR2_X1 U9328 ( .A1(n7911), .A2(n8106), .ZN(n11092) );
  INV_X1 U9329 ( .A(n10143), .ZN(n10283) );
  NAND2_X1 U9330 ( .A1(n10283), .A2(n11090), .ZN(n7913) );
  AOI22_X1 U9331 ( .A1(n11069), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n9651), .B2(
        n11067), .ZN(n7912) );
  OAI211_X1 U9332 ( .C1(n7914), .C2(n10287), .A(n7913), .B(n7912), .ZN(n7915)
         );
  AOI21_X1 U9333 ( .B1(n10223), .B2(n9663), .A(n7915), .ZN(n7916) );
  OAI21_X1 U9334 ( .B1(n11092), .B2(n10219), .A(n7916), .ZN(n7917) );
  AOI21_X1 U9335 ( .B1(n11094), .B2(n10307), .A(n7917), .ZN(n7918) );
  OAI21_X1 U9336 ( .B1(n11086), .B2(n10309), .A(n7918), .ZN(P1_U3282) );
  OAI22_X1 U9337 ( .A1(n10307), .A2(n7921), .B1(n7920), .B2(n7919), .ZN(n7922)
         );
  AOI21_X1 U9338 ( .B1(n10223), .B2(n7923), .A(n7922), .ZN(n7924) );
  OAI21_X1 U9339 ( .B1(n10219), .B2(n7925), .A(n7924), .ZN(n7926) );
  AOI21_X1 U9340 ( .B1(n11075), .B2(n7927), .A(n7926), .ZN(n7928) );
  OAI21_X1 U9341 ( .B1(n7929), .B2(n11079), .A(n7928), .ZN(P1_U3289) );
  NAND2_X1 U9342 ( .A1(n11065), .A2(n7930), .ZN(n7932) );
  AOI22_X1 U9343 ( .A1(n11069), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n11067), .ZN(n7931) );
  OAI211_X1 U9344 ( .C1(n8074), .C2(n11072), .A(n7932), .B(n7931), .ZN(n7933)
         );
  AOI21_X1 U9345 ( .B1(n11075), .B2(n7934), .A(n7933), .ZN(n7935) );
  OAI21_X1 U9346 ( .B1(n7936), .B2(n11069), .A(n7935), .ZN(P1_U3291) );
  NAND2_X1 U9347 ( .A1(n7937), .A2(n9827), .ZN(n7938) );
  XNOR2_X1 U9348 ( .A(n7938), .B(n9847), .ZN(n7939) );
  OAI222_X1 U9349 ( .A1(n10375), .A2(n8141), .B1(n10388), .B2(n7940), .C1(
        n7939), .C2(n11022), .ZN(n11057) );
  INV_X1 U9350 ( .A(n11057), .ZN(n7951) );
  OAI21_X1 U9351 ( .B1(n7942), .B2(n9847), .A(n7941), .ZN(n11059) );
  INV_X1 U9352 ( .A(n7943), .ZN(n7945) );
  OAI211_X1 U9353 ( .C1(n7945), .C2(n11056), .A(n10400), .B(n7944), .ZN(n11055) );
  NAND2_X1 U9354 ( .A1(n10223), .A2(n7946), .ZN(n7948) );
  AOI22_X1 U9355 ( .A1(n11069), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7989), .B2(
        n11067), .ZN(n7947) );
  OAI211_X1 U9356 ( .C1(n11055), .C2(n10219), .A(n7948), .B(n7947), .ZN(n7949)
         );
  AOI21_X1 U9357 ( .B1(n11059), .B2(n11075), .A(n7949), .ZN(n7950) );
  OAI21_X1 U9358 ( .B1(n7951), .B2(n11079), .A(n7950), .ZN(P1_U3288) );
  NAND2_X1 U9359 ( .A1(n7952), .A2(n11075), .ZN(n7957) );
  AOI22_X1 U9360 ( .A1(n11069), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n9542), .B2(
        n11067), .ZN(n7953) );
  OAI21_X1 U9361 ( .B1(n5700), .B2(n11072), .A(n7953), .ZN(n7954) );
  AOI21_X1 U9362 ( .B1(n7955), .B2(n11065), .A(n7954), .ZN(n7956) );
  OAI211_X1 U9363 ( .C1(n11079), .C2(n7958), .A(n7957), .B(n7956), .ZN(
        P1_U3283) );
  NAND2_X1 U9364 ( .A1(n7959), .A2(n11075), .ZN(n7967) );
  NOR2_X1 U9365 ( .A1(n11072), .A2(n8147), .ZN(n7964) );
  NAND2_X1 U9366 ( .A1(n10283), .A2(n10000), .ZN(n7961) );
  AOI22_X1 U9367 ( .A1(n11069), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n8140), .B2(
        n11067), .ZN(n7960) );
  OAI211_X1 U9368 ( .C1(n7962), .C2(n10287), .A(n7961), .B(n7960), .ZN(n7963)
         );
  AOI211_X1 U9369 ( .C1(n7965), .C2(n11065), .A(n7964), .B(n7963), .ZN(n7966)
         );
  OAI211_X1 U9370 ( .C1(n7968), .C2(n10292), .A(n7967), .B(n7966), .ZN(
        P1_U3286) );
  NAND2_X1 U9371 ( .A1(n9377), .A2(n8385), .ZN(n7969) );
  OAI22_X1 U9372 ( .A1(n9317), .A2(n7970), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n9380), .ZN(n7973) );
  MUX2_X1 U9373 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n7971), .S(n9377), .Z(n7972)
         );
  AOI211_X1 U9374 ( .C1(n9320), .C2(n7974), .A(n7973), .B(n7972), .ZN(n7975)
         );
  INV_X1 U9375 ( .A(n7975), .ZN(P2_U3230) );
  OAI22_X1 U9376 ( .A1(n7976), .A2(n8509), .B1(n7537), .B2(n9380), .ZN(n7977)
         );
  OAI21_X1 U9377 ( .B1(n7978), .B2(n7977), .A(n9377), .ZN(n7981) );
  NAND2_X1 U9378 ( .A1(n7979), .A2(n9320), .ZN(n7980) );
  OAI211_X1 U9379 ( .C1(n7982), .C2(n9377), .A(n7981), .B(n7980), .ZN(P2_U3231) );
  NOR2_X1 U9380 ( .A1(n7983), .A2(n5215), .ZN(n7985) );
  XNOR2_X1 U9381 ( .A(n7985), .B(n7984), .ZN(n7992) );
  AOI22_X1 U9382 ( .A1(n9678), .A2(n10002), .B1(n9687), .B2(n10000), .ZN(n7991) );
  INV_X1 U9383 ( .A(n7986), .ZN(n7988) );
  NOR2_X1 U9384 ( .A1(n9636), .A2(n11056), .ZN(n7987) );
  AOI211_X1 U9385 ( .C1(n9689), .C2(n7989), .A(n7988), .B(n7987), .ZN(n7990)
         );
  OAI211_X1 U9386 ( .C1(n7992), .C2(n9697), .A(n7991), .B(n7990), .ZN(P1_U3227) );
  INV_X1 U9387 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7995) );
  XNOR2_X1 U9388 ( .A(n8166), .B(n8183), .ZN(n7994) );
  AOI21_X1 U9389 ( .B1(n7995), .B2(n7994), .A(n8167), .ZN(n8011) );
  INV_X1 U9390 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7999) );
  AOI21_X1 U9391 ( .B1(n7999), .B2(n7998), .A(n8184), .ZN(n8000) );
  NOR2_X1 U9392 ( .A1(n8000), .A2(n11014), .ZN(n8009) );
  MUX2_X1 U9393 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8174), .Z(n8171) );
  XOR2_X1 U9394 ( .A(n8183), .B(n8171), .Z(n8004) );
  NOR2_X1 U9395 ( .A1(n8003), .A2(n8004), .ZN(n8172) );
  AOI21_X1 U9396 ( .B1(n8004), .B2(n8003), .A(n8172), .ZN(n8007) );
  NOR2_X1 U9397 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10556), .ZN(n8092) );
  AOI21_X1 U9398 ( .B1(n10996), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n8092), .ZN(
        n8006) );
  NAND2_X1 U9399 ( .A1(n10997), .A2(n8183), .ZN(n8005) );
  OAI211_X1 U9400 ( .C1(n8007), .C2(n9164), .A(n8006), .B(n8005), .ZN(n8008)
         );
  NOR2_X1 U9401 ( .A1(n8009), .A2(n8008), .ZN(n8010) );
  OAI21_X1 U9402 ( .B1(n8011), .B2(n11005), .A(n8010), .ZN(P2_U3191) );
  NOR2_X1 U9403 ( .A1(n8012), .A2(n9450), .ZN(n8014) );
  AOI211_X1 U9404 ( .C1(n8016), .C2(n8015), .A(n8014), .B(n8013), .ZN(n11054)
         );
  OR2_X1 U9405 ( .A1(n11054), .A2(n9465), .ZN(n8017) );
  OAI21_X1 U9406 ( .B1(n9456), .B2(n8018), .A(n8017), .ZN(P2_U3464) );
  NAND2_X1 U9407 ( .A1(n5755), .A2(n8019), .ZN(n8020) );
  XNOR2_X1 U9408 ( .A(n8021), .B(n8020), .ZN(n8028) );
  AOI22_X1 U9409 ( .A1(n9678), .A2(n10001), .B1(n8022), .B2(n9694), .ZN(n8027)
         );
  INV_X1 U9410 ( .A(n8023), .ZN(n8025) );
  NOR2_X1 U9411 ( .A1(n9644), .A2(n8235), .ZN(n8024) );
  AOI211_X1 U9412 ( .C1(n9689), .C2(n11068), .A(n8025), .B(n8024), .ZN(n8026)
         );
  OAI211_X1 U9413 ( .C1(n8028), .C2(n9697), .A(n8027), .B(n8026), .ZN(P1_U3239) );
  INV_X1 U9414 ( .A(n8029), .ZN(n8035) );
  INV_X1 U9415 ( .A(n8030), .ZN(n8031) );
  MUX2_X1 U9416 ( .A(n10937), .B(n8031), .S(n9377), .Z(n8034) );
  AOI22_X1 U9417 ( .A1(n9364), .A2(n8032), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n9314), .ZN(n8033) );
  OAI211_X1 U9418 ( .C1(n9388), .C2(n8035), .A(n8034), .B(n8033), .ZN(P2_U3232) );
  INV_X1 U9419 ( .A(n8036), .ZN(n8043) );
  INV_X1 U9420 ( .A(n8037), .ZN(n8038) );
  MUX2_X1 U9421 ( .A(n7230), .B(n8038), .S(n9377), .Z(n8042) );
  AOI22_X1 U9422 ( .A1(n9364), .A2(n8040), .B1(n9314), .B2(n8039), .ZN(n8041)
         );
  OAI211_X1 U9423 ( .C1(n9388), .C2(n8043), .A(n8042), .B(n8041), .ZN(P2_U3229) );
  AOI22_X1 U9424 ( .A1(n6410), .A2(n9547), .B1(n11109), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n8044) );
  OAI21_X1 U9425 ( .B1(n8045), .B2(n11109), .A(n8044), .ZN(P1_U3532) );
  NAND2_X1 U9426 ( .A1(n8049), .A2(n8048), .ZN(n8089) );
  XNOR2_X1 U9427 ( .A(n8290), .B(n8678), .ZN(n8050) );
  NOR2_X1 U9428 ( .A1(n8050), .A2(n9044), .ZN(n8088) );
  INV_X1 U9429 ( .A(n8088), .ZN(n8051) );
  NAND2_X1 U9430 ( .A1(n8050), .A2(n9044), .ZN(n8087) );
  NAND2_X1 U9431 ( .A1(n8051), .A2(n8087), .ZN(n8052) );
  XNOR2_X1 U9432 ( .A(n8089), .B(n8052), .ZN(n8058) );
  AOI21_X1 U9433 ( .B1(n9046), .B2(n8827), .A(n8053), .ZN(n8055) );
  NAND2_X1 U9434 ( .A1(n8831), .A2(n8250), .ZN(n8054) );
  OAI211_X1 U9435 ( .C1(n8390), .C2(n8829), .A(n8055), .B(n8054), .ZN(n8056)
         );
  AOI21_X1 U9436 ( .B1(n8251), .B2(n8786), .A(n8056), .ZN(n8057) );
  OAI21_X1 U9437 ( .B1(n8058), .B2(n8788), .A(n8057), .ZN(P2_U3161) );
  INV_X1 U9438 ( .A(n8059), .ZN(n8631) );
  OAI222_X1 U9439 ( .A1(n9513), .A2(n8061), .B1(n8667), .B2(n8631), .C1(
        P2_U3151), .C2(n8060), .ZN(P2_U3273) );
  INV_X1 U9440 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n8062) );
  OAI22_X1 U9441 ( .A1(n10366), .A2(n8063), .B1(n11110), .B2(n8062), .ZN(n8064) );
  INV_X1 U9442 ( .A(n8064), .ZN(n8065) );
  OAI21_X1 U9443 ( .B1(n8066), .B2(n11109), .A(n8065), .ZN(P1_U3531) );
  OAI22_X1 U9444 ( .A1(n10366), .A2(n11073), .B1(n11110), .B2(n7343), .ZN(
        n8067) );
  INV_X1 U9445 ( .A(n8067), .ZN(n8068) );
  OAI21_X1 U9446 ( .B1(n8069), .B2(n11109), .A(n8068), .ZN(P1_U3528) );
  OAI22_X1 U9447 ( .A1(n10366), .A2(n6009), .B1(n11110), .B2(n8070), .ZN(n8071) );
  AOI21_X1 U9448 ( .B1(n8072), .B2(n11110), .A(n8071), .ZN(n8073) );
  INV_X1 U9449 ( .A(n8073), .ZN(P1_U3526) );
  OAI22_X1 U9450 ( .A1(n10366), .A2(n8074), .B1(n11110), .B2(n7320), .ZN(n8075) );
  INV_X1 U9451 ( .A(n8075), .ZN(n8076) );
  OAI21_X1 U9452 ( .B1(n8077), .B2(n11109), .A(n8076), .ZN(P1_U3524) );
  INV_X1 U9453 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n8078) );
  OAI22_X1 U9454 ( .A1(n10366), .A2(n8147), .B1(n11110), .B2(n8078), .ZN(n8079) );
  AOI21_X1 U9455 ( .B1(n8080), .B2(n11110), .A(n8079), .ZN(n8081) );
  INV_X1 U9456 ( .A(n8081), .ZN(P1_U3529) );
  INV_X1 U9457 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n8082) );
  OAI22_X1 U9458 ( .A1(n10366), .A2(n8083), .B1(n11110), .B2(n8082), .ZN(n8084) );
  AOI21_X1 U9459 ( .B1(n8085), .B2(n11110), .A(n8084), .ZN(n8086) );
  INV_X1 U9460 ( .A(n8086), .ZN(P1_U3530) );
  XNOR2_X1 U9461 ( .A(n8321), .B(n8694), .ZN(n8219) );
  XNOR2_X1 U9462 ( .A(n8219), .B(n8390), .ZN(n8090) );
  OAI211_X1 U9463 ( .C1(n8091), .C2(n8090), .A(n8221), .B(n8824), .ZN(n8098)
         );
  AOI21_X1 U9464 ( .B1(n9044), .B2(n8827), .A(n8092), .ZN(n8095) );
  NAND2_X1 U9465 ( .A1(n8831), .A2(n8320), .ZN(n8094) );
  NAND2_X1 U9466 ( .A1(n9042), .A2(n8815), .ZN(n8093) );
  NAND3_X1 U9467 ( .A1(n8095), .A2(n8094), .A3(n8093), .ZN(n8096) );
  AOI21_X1 U9468 ( .B1(n8321), .B2(n8786), .A(n8096), .ZN(n8097) );
  NAND2_X1 U9469 ( .A1(n8098), .A2(n8097), .ZN(P2_U3171) );
  INV_X1 U9470 ( .A(n8100), .ZN(n9784) );
  XNOR2_X1 U9471 ( .A(n8099), .B(n9784), .ZN(n11108) );
  INV_X1 U9472 ( .A(n11108), .ZN(n8113) );
  NAND2_X1 U9473 ( .A1(n8101), .A2(n8100), .ZN(n8102) );
  NAND3_X1 U9474 ( .A1(n8103), .A2(n10411), .A3(n8102), .ZN(n8105) );
  AOI22_X1 U9475 ( .A1(n11089), .A2(n9996), .B1(n11088), .B2(n10415), .ZN(
        n8104) );
  NAND2_X1 U9476 ( .A1(n8105), .A2(n8104), .ZN(n11106) );
  OAI211_X1 U9477 ( .C1(n8106), .C2(n11104), .A(n10400), .B(n8203), .ZN(n11102) );
  AOI22_X1 U9478 ( .A1(n11069), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n8107), .B2(
        n11067), .ZN(n8110) );
  NAND2_X1 U9479 ( .A1(n8108), .A2(n10223), .ZN(n8109) );
  OAI211_X1 U9480 ( .C1(n11102), .C2(n10219), .A(n8110), .B(n8109), .ZN(n8111)
         );
  AOI21_X1 U9481 ( .B1(n11106), .B2(n10307), .A(n8111), .ZN(n8112) );
  OAI21_X1 U9482 ( .B1(n8113), .B2(n10309), .A(n8112), .ZN(P1_U3281) );
  NAND2_X1 U9483 ( .A1(n8117), .A2(n10476), .ZN(n8115) );
  OR2_X1 U9484 ( .A1(n8114), .A2(P1_U3086), .ZN(n9756) );
  OAI211_X1 U9485 ( .C1(n8116), .C2(n8627), .A(n8115), .B(n9756), .ZN(P1_U3332) );
  NAND2_X1 U9486 ( .A1(n8117), .A2(n8609), .ZN(n8119) );
  OR2_X1 U9487 ( .A1(n8118), .A2(P2_U3151), .ZN(n9031) );
  OAI211_X1 U9488 ( .C1(n8120), .C2(n9513), .A(n8119), .B(n9031), .ZN(P2_U3272) );
  INV_X1 U9489 ( .A(n8853), .ZN(n8121) );
  NAND3_X1 U9490 ( .A1(n8122), .A2(n8909), .A3(n8121), .ZN(n8123) );
  NAND2_X1 U9491 ( .A1(n8124), .A2(n8123), .ZN(n8163) );
  INV_X1 U9492 ( .A(n8163), .ZN(n8133) );
  XNOR2_X1 U9493 ( .A(n8125), .B(n8853), .ZN(n8126) );
  OAI222_X1 U9494 ( .A1(n9376), .A2(n8047), .B1(n9361), .B2(n8127), .C1(n8126), 
        .C2(n9373), .ZN(n8161) );
  INV_X1 U9495 ( .A(n8161), .ZN(n8128) );
  MUX2_X1 U9496 ( .A(n7288), .B(n8128), .S(n9377), .Z(n8132) );
  AOI22_X1 U9497 ( .A1(n9364), .A2(n8130), .B1(n9314), .B2(n8129), .ZN(n8131)
         );
  OAI211_X1 U9498 ( .C1(n9388), .C2(n8133), .A(n8132), .B(n8131), .ZN(P2_U3227) );
  XNOR2_X1 U9499 ( .A(n8135), .B(n8134), .ZN(n8136) );
  XNOR2_X1 U9500 ( .A(n8137), .B(n8136), .ZN(n8138) );
  NAND2_X1 U9501 ( .A1(n8138), .A2(n9676), .ZN(n8146) );
  INV_X1 U9502 ( .A(n8139), .ZN(n8144) );
  INV_X1 U9503 ( .A(n8140), .ZN(n8142) );
  OAI22_X1 U9504 ( .A1(n9646), .A2(n8142), .B1(n9691), .B2(n8141), .ZN(n8143)
         );
  AOI211_X1 U9505 ( .C1(n9687), .C2(n9998), .A(n8144), .B(n8143), .ZN(n8145)
         );
  OAI211_X1 U9506 ( .C1(n8147), .C2(n9636), .A(n8146), .B(n8145), .ZN(P1_U3213) );
  XOR2_X1 U9507 ( .A(n8148), .B(n8919), .Z(n8149) );
  OAI222_X1 U9508 ( .A1(n9376), .A2(n8151), .B1(n9361), .B2(n8150), .C1(n8149), 
        .C2(n9373), .ZN(n8210) );
  INV_X1 U9509 ( .A(n8210), .ZN(n8159) );
  INV_X1 U9510 ( .A(n8152), .ZN(n8153) );
  AOI21_X1 U9511 ( .B1(n8919), .B2(n8154), .A(n8153), .ZN(n8211) );
  AOI22_X1 U9512 ( .A1(n9315), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n9314), .B2(
        n8155), .ZN(n8156) );
  OAI21_X1 U9513 ( .B1(n8931), .B2(n9317), .A(n8156), .ZN(n8157) );
  AOI21_X1 U9514 ( .B1(n8211), .B2(n9320), .A(n8157), .ZN(n8158) );
  OAI21_X1 U9515 ( .B1(n8159), .B2(n9353), .A(n8158), .ZN(P2_U3226) );
  NOR2_X1 U9516 ( .A1(n8160), .A2(n9450), .ZN(n8162) );
  AOI211_X1 U9517 ( .C1(n9414), .C2(n8163), .A(n8162), .B(n8161), .ZN(n11064)
         );
  OR2_X1 U9518 ( .A1(n11064), .A2(n9465), .ZN(n8164) );
  OAI21_X1 U9519 ( .B1(n9456), .B2(n8165), .A(n8164), .ZN(P2_U3465) );
  NAND2_X1 U9520 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n8269), .ZN(n8168) );
  OAI21_X1 U9521 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n8269), .A(n8168), .ZN(
        n8169) );
  AOI21_X1 U9522 ( .B1(n8170), .B2(n8169), .A(n8254), .ZN(n8193) );
  INV_X1 U9523 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n8181) );
  INV_X1 U9524 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10661) );
  NOR2_X1 U9525 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10661), .ZN(n8222) );
  INV_X1 U9526 ( .A(n8171), .ZN(n8173) );
  MUX2_X1 U9527 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8174), .Z(n8175) );
  AND2_X1 U9528 ( .A1(n8175), .A2(n8269), .ZN(n8259) );
  OR2_X1 U9529 ( .A1(n8175), .A2(n8269), .ZN(n8260) );
  INV_X1 U9530 ( .A(n8260), .ZN(n8176) );
  NOR2_X1 U9531 ( .A1(n8259), .A2(n8176), .ZN(n8178) );
  OAI21_X1 U9532 ( .B1(n8261), .B2(n8178), .A(n11010), .ZN(n8177) );
  AOI21_X1 U9533 ( .B1(n8261), .B2(n8178), .A(n8177), .ZN(n8179) );
  NOR2_X1 U9534 ( .A1(n8222), .A2(n8179), .ZN(n8180) );
  OAI21_X1 U9535 ( .B1(n9095), .B2(n8181), .A(n8180), .ZN(n8190) );
  NOR2_X1 U9536 ( .A1(n8182), .A2(n8183), .ZN(n8185) );
  NAND2_X1 U9537 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n8269), .ZN(n8186) );
  OAI21_X1 U9538 ( .B1(n8269), .B2(P2_REG2_REG_10__SCAN_IN), .A(n8186), .ZN(
        n8187) );
  AOI21_X1 U9539 ( .B1(n5214), .B2(n8187), .A(n8268), .ZN(n8188) );
  NOR2_X1 U9540 ( .A1(n8188), .A2(n11014), .ZN(n8189) );
  AOI211_X1 U9541 ( .C1(n10997), .C2(n8191), .A(n8190), .B(n8189), .ZN(n8192)
         );
  OAI21_X1 U9542 ( .B1(n8193), .B2(n11005), .A(n8192), .ZN(P2_U3192) );
  INV_X1 U9543 ( .A(n8194), .ZN(n8284) );
  OAI222_X1 U9544 ( .A1(n8667), .A2(n8284), .B1(P2_U3151), .B2(n8196), .C1(
        n8195), .C2(n9513), .ZN(P2_U3271) );
  OAI21_X1 U9545 ( .B1(n5213), .B2(n9785), .A(n8197), .ZN(n8198) );
  INV_X1 U9546 ( .A(n8198), .ZN(n8305) );
  XNOR2_X1 U9547 ( .A(n8199), .B(n9785), .ZN(n8307) );
  NAND2_X1 U9548 ( .A1(n8307), .A2(n11075), .ZN(n8209) );
  NAND2_X1 U9549 ( .A1(n10283), .A2(n11087), .ZN(n8202) );
  AOI22_X1 U9550 ( .A1(n11069), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n8200), .B2(
        n11067), .ZN(n8201) );
  OAI211_X1 U9551 ( .C1(n9692), .C2(n10287), .A(n8202), .B(n8201), .ZN(n8206)
         );
  INV_X1 U9552 ( .A(n8203), .ZN(n8204) );
  OAI211_X1 U9553 ( .C1(n8204), .C2(n9637), .A(n10400), .B(n8360), .ZN(n8303)
         );
  NOR2_X1 U9554 ( .A1(n8303), .A2(n10219), .ZN(n8205) );
  AOI211_X1 U9555 ( .C1(n10223), .C2(n8207), .A(n8206), .B(n8205), .ZN(n8208)
         );
  OAI211_X1 U9556 ( .C1(n8305), .C2(n10292), .A(n8209), .B(n8208), .ZN(
        P1_U3280) );
  AOI21_X1 U9557 ( .B1(n8211), .B2(n9414), .A(n8210), .ZN(n8218) );
  OAI22_X1 U9558 ( .A1(n8931), .A2(n9432), .B1(n9456), .B2(n8212), .ZN(n8213)
         );
  INV_X1 U9559 ( .A(n8213), .ZN(n8214) );
  OAI21_X1 U9560 ( .B1(n8218), .B2(n9465), .A(n8214), .ZN(P2_U3466) );
  INV_X1 U9561 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n8215) );
  OAI22_X1 U9562 ( .A1(n9508), .A2(n8931), .B1(n11121), .B2(n8215), .ZN(n8216)
         );
  INV_X1 U9563 ( .A(n8216), .ZN(n8217) );
  OAI21_X1 U9564 ( .B1(n8218), .B2(n6890), .A(n8217), .ZN(P2_U3411) );
  INV_X1 U9565 ( .A(n8219), .ZN(n8220) );
  XNOR2_X1 U9566 ( .A(n8479), .B(n8694), .ZN(n8330) );
  XNOR2_X1 U9567 ( .A(n8332), .B(n8334), .ZN(n8227) );
  INV_X1 U9568 ( .A(n8390), .ZN(n9043) );
  AOI21_X1 U9569 ( .B1(n9043), .B2(n8827), .A(n8222), .ZN(n8224) );
  NAND2_X1 U9570 ( .A1(n8831), .A2(n8395), .ZN(n8223) );
  OAI211_X1 U9571 ( .C1(n8402), .C2(n8829), .A(n8224), .B(n8223), .ZN(n8225)
         );
  AOI21_X1 U9572 ( .B1(n8479), .B2(n8786), .A(n8225), .ZN(n8226) );
  OAI21_X1 U9573 ( .B1(n8227), .B2(n8788), .A(n8226), .ZN(P2_U3157) );
  INV_X1 U9574 ( .A(n8228), .ZN(n8243) );
  OAI222_X1 U9575 ( .A1(n8667), .A2(n8243), .B1(P2_U3151), .B2(n8230), .C1(
        n8229), .C2(n9513), .ZN(P2_U3270) );
  XNOR2_X1 U9576 ( .A(n8232), .B(n8231), .ZN(n8242) );
  INV_X1 U9577 ( .A(n8233), .ZN(n8238) );
  INV_X1 U9578 ( .A(n8234), .ZN(n8236) );
  OAI22_X1 U9579 ( .A1(n9646), .A2(n8236), .B1(n9691), .B2(n8235), .ZN(n8237)
         );
  AOI211_X1 U9580 ( .C1(n9687), .C2(n9997), .A(n8238), .B(n8237), .ZN(n8241)
         );
  NAND2_X1 U9581 ( .A1(n9694), .A2(n8239), .ZN(n8240) );
  OAI211_X1 U9582 ( .C1(n8242), .C2(n9697), .A(n8241), .B(n8240), .ZN(P1_U3221) );
  OAI222_X1 U9583 ( .A1(P1_U3086), .A2(n8244), .B1(n8633), .B2(n8243), .C1(
        n10775), .C2(n10471), .ZN(P1_U3330) );
  NAND2_X1 U9584 ( .A1(n8152), .A2(n8245), .ZN(n8246) );
  XOR2_X1 U9585 ( .A(n8855), .B(n8246), .Z(n8286) );
  XNOR2_X1 U9586 ( .A(n8247), .B(n8855), .ZN(n8248) );
  AOI222_X1 U9587 ( .A1(n9342), .A2(n8248), .B1(n9043), .B2(n9337), .C1(n9046), 
        .C2(n9339), .ZN(n8285) );
  MUX2_X1 U9588 ( .A(n8249), .B(n8285), .S(n9377), .Z(n8253) );
  AOI22_X1 U9589 ( .A1(n8251), .A2(n9364), .B1(n9314), .B2(n8250), .ZN(n8252)
         );
  OAI211_X1 U9590 ( .C1(n9388), .C2(n8286), .A(n8253), .B(n8252), .ZN(P2_U3225) );
  NOR2_X1 U9591 ( .A1(n10998), .A2(n8255), .ZN(n8256) );
  INV_X1 U9592 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n11004) );
  INV_X1 U9593 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8502) );
  AOI22_X1 U9594 ( .A1(n8273), .A2(P2_REG1_REG_12__SCAN_IN), .B1(n8502), .B2(
        n8577), .ZN(n8257) );
  AOI21_X1 U9595 ( .B1(n8258), .B2(n8257), .A(n8542), .ZN(n8283) );
  MUX2_X1 U9596 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8174), .Z(n8561) );
  XNOR2_X1 U9597 ( .A(n8561), .B(n8273), .ZN(n8265) );
  MUX2_X1 U9598 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8174), .Z(n8262) );
  OR2_X1 U9599 ( .A1(n8262), .A2(n8271), .ZN(n8263) );
  XNOR2_X1 U9600 ( .A(n8262), .B(n10998), .ZN(n11009) );
  NAND2_X1 U9601 ( .A1(n11008), .A2(n11009), .ZN(n11007) );
  NAND2_X1 U9602 ( .A1(n8263), .A2(n11007), .ZN(n8264) );
  NAND2_X1 U9603 ( .A1(n8265), .A2(n8264), .ZN(n8562) );
  OAI21_X1 U9604 ( .B1(n8265), .B2(n8264), .A(n8562), .ZN(n8281) );
  NAND2_X1 U9605 ( .A1(n10996), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n8267) );
  NOR2_X1 U9606 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10732), .ZN(n8408) );
  INV_X1 U9607 ( .A(n8408), .ZN(n8266) );
  OAI211_X1 U9608 ( .C1(n10983), .C2(n8577), .A(n8267), .B(n8266), .ZN(n8280)
         );
  AOI21_X1 U9609 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n8269), .A(n8268), .ZN(
        n8270) );
  NOR2_X1 U9610 ( .A1(n10998), .A2(n8270), .ZN(n8272) );
  INV_X1 U9611 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11001) );
  INV_X1 U9612 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8274) );
  MUX2_X1 U9613 ( .A(n8274), .B(P2_REG2_REG_12__SCAN_IN), .S(n8273), .Z(n8275)
         );
  INV_X1 U9614 ( .A(n8275), .ZN(n8276) );
  AOI21_X1 U9615 ( .B1(n8277), .B2(n8276), .A(n8576), .ZN(n8278) );
  NOR2_X1 U9616 ( .A1(n8278), .A2(n11014), .ZN(n8279) );
  AOI211_X1 U9617 ( .C1(n11010), .C2(n8281), .A(n8280), .B(n8279), .ZN(n8282)
         );
  OAI21_X1 U9618 ( .B1(n8283), .B2(n11005), .A(n8282), .ZN(P2_U3194) );
  OAI222_X1 U9619 ( .A1(P1_U3086), .A2(n6392), .B1(n8633), .B2(n8284), .C1(
        n10773), .C2(n10471), .ZN(P1_U3331) );
  OAI21_X1 U9620 ( .B1(n9458), .B2(n8286), .A(n8285), .ZN(n8292) );
  OAI22_X1 U9621 ( .A1(n8290), .A2(n9432), .B1(n9456), .B2(n7857), .ZN(n8287)
         );
  AOI21_X1 U9622 ( .B1(n8292), .B2(n9456), .A(n8287), .ZN(n8288) );
  INV_X1 U9623 ( .A(n8288), .ZN(P2_U3467) );
  INV_X1 U9624 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n8289) );
  OAI22_X1 U9625 ( .A1(n9508), .A2(n8290), .B1(n11121), .B2(n8289), .ZN(n8291)
         );
  AOI21_X1 U9626 ( .B1(n8292), .B2(n11121), .A(n8291), .ZN(n8293) );
  INV_X1 U9627 ( .A(n8293), .ZN(P2_U3414) );
  XNOR2_X1 U9628 ( .A(n8295), .B(n8294), .ZN(n8302) );
  AND2_X1 U9629 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n10039) );
  INV_X1 U9630 ( .A(n8296), .ZN(n8297) );
  OAI22_X1 U9631 ( .A1(n9646), .A2(n8297), .B1(n9644), .B2(n9654), .ZN(n8298)
         );
  AOI211_X1 U9632 ( .C1(n9678), .C2(n9998), .A(n10039), .B(n8298), .ZN(n8301)
         );
  NAND2_X1 U9633 ( .A1(n9694), .A2(n8299), .ZN(n8300) );
  OAI211_X1 U9634 ( .C1(n8302), .C2(n9697), .A(n8301), .B(n8300), .ZN(P1_U3231) );
  INV_X1 U9635 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n8423) );
  INV_X1 U9636 ( .A(n9692), .ZN(n10406) );
  AOI22_X1 U9637 ( .A1(n10406), .A2(n11088), .B1(n11089), .B2(n11087), .ZN(
        n8304) );
  OAI211_X1 U9638 ( .C1(n8305), .C2(n11022), .A(n8304), .B(n8303), .ZN(n8306)
         );
  AOI21_X1 U9639 ( .B1(n8307), .B2(n11107), .A(n8306), .ZN(n8309) );
  MUX2_X1 U9640 ( .A(n8423), .B(n8309), .S(n11110), .Z(n8308) );
  OAI21_X1 U9641 ( .B1(n9637), .B2(n10366), .A(n8308), .ZN(P1_U3535) );
  INV_X1 U9642 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n8310) );
  MUX2_X1 U9643 ( .A(n8310), .B(n8309), .S(n11114), .Z(n8311) );
  OAI21_X1 U9644 ( .B1(n9637), .B2(n10457), .A(n8311), .ZN(P1_U3492) );
  OAI21_X1 U9645 ( .B1(n5754), .B2(n6817), .A(n8312), .ZN(n8324) );
  NAND2_X1 U9646 ( .A1(n8247), .A2(n8855), .ZN(n8314) );
  NAND2_X1 U9647 ( .A1(n8314), .A2(n8313), .ZN(n8386) );
  XNOR2_X1 U9648 ( .A(n8386), .B(n8856), .ZN(n8315) );
  AOI222_X1 U9649 ( .A1(n9342), .A2(n8315), .B1(n9044), .B2(n9339), .C1(n9042), 
        .C2(n9337), .ZN(n8319) );
  OAI21_X1 U9650 ( .B1(n9458), .B2(n8324), .A(n8319), .ZN(n8351) );
  INV_X1 U9651 ( .A(n8351), .ZN(n8318) );
  INV_X1 U9652 ( .A(n9432), .ZN(n8316) );
  AOI22_X1 U9653 ( .A1(n8321), .A2(n8316), .B1(n9465), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n8317) );
  OAI21_X1 U9654 ( .B1(n8318), .B2(n9465), .A(n8317), .ZN(P2_U3468) );
  MUX2_X1 U9655 ( .A(n7999), .B(n8319), .S(n9377), .Z(n8323) );
  AOI22_X1 U9656 ( .A1(n8321), .A2(n9364), .B1(n9314), .B2(n8320), .ZN(n8322)
         );
  OAI211_X1 U9657 ( .C1(n9388), .C2(n8324), .A(n8323), .B(n8322), .ZN(P2_U3224) );
  XNOR2_X1 U9658 ( .A(n6595), .B(n8860), .ZN(n8325) );
  OAI222_X1 U9659 ( .A1(n9376), .A2(n8507), .B1(n9361), .B2(n8334), .C1(n9373), 
        .C2(n8325), .ZN(n8340) );
  OR2_X1 U9660 ( .A1(n8326), .A2(n8937), .ZN(n8371) );
  NAND2_X1 U9661 ( .A1(n8371), .A2(n8924), .ZN(n8327) );
  XOR2_X1 U9662 ( .A(n8860), .B(n8327), .Z(n8347) );
  OAI22_X1 U9663 ( .A1(n8347), .A2(n9458), .B1(n8339), .B2(n9450), .ZN(n8328)
         );
  NOR2_X1 U9664 ( .A1(n8340), .A2(n8328), .ZN(n11083) );
  NAND2_X1 U9665 ( .A1(n9465), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8329) );
  OAI21_X1 U9666 ( .B1(n11083), .B2(n9465), .A(n8329), .ZN(P2_U3470) );
  XNOR2_X1 U9667 ( .A(n8339), .B(n8694), .ZN(n8401) );
  XNOR2_X1 U9668 ( .A(n8401), .B(n9041), .ZN(n8403) );
  XNOR2_X1 U9669 ( .A(n8404), .B(n8403), .ZN(n8333) );
  NAND2_X1 U9670 ( .A1(n8333), .A2(n8824), .ZN(n8338) );
  NOR2_X1 U9671 ( .A1(n8507), .A2(n8829), .ZN(n8336) );
  INV_X1 U9672 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n11019) );
  OAI22_X1 U9673 ( .A1(n8334), .A2(n8817), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11019), .ZN(n8335) );
  AOI211_X1 U9674 ( .C1(n8341), .C2(n8831), .A(n8336), .B(n8335), .ZN(n8337)
         );
  OAI211_X1 U9675 ( .C1(n8339), .C2(n8835), .A(n8338), .B(n8337), .ZN(P2_U3176) );
  NAND2_X1 U9676 ( .A1(n8340), .A2(n9377), .ZN(n8346) );
  INV_X1 U9677 ( .A(n8341), .ZN(n8342) );
  OAI22_X1 U9678 ( .A1(n9377), .A2(n11001), .B1(n8342), .B2(n9380), .ZN(n8343)
         );
  AOI21_X1 U9679 ( .B1(n8344), .B2(n9364), .A(n8343), .ZN(n8345) );
  OAI211_X1 U9680 ( .C1(n9388), .C2(n8347), .A(n8346), .B(n8345), .ZN(P2_U3222) );
  INV_X1 U9681 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n8348) );
  OAI22_X1 U9682 ( .A1(n8349), .A2(n9508), .B1(n11121), .B2(n8348), .ZN(n8350)
         );
  AOI21_X1 U9683 ( .B1(n8351), .B2(n11121), .A(n8350), .ZN(n8352) );
  INV_X1 U9684 ( .A(n8352), .ZN(P2_U3417) );
  XNOR2_X1 U9685 ( .A(n8353), .B(n9896), .ZN(n8354) );
  NAND2_X1 U9686 ( .A1(n8354), .A2(n10411), .ZN(n10420) );
  OAI21_X1 U9687 ( .B1(n8356), .B2(n9787), .A(n8355), .ZN(n10422) );
  INV_X1 U9688 ( .A(n10422), .ZN(n8357) );
  NAND2_X1 U9689 ( .A1(n8357), .A2(n11075), .ZN(n8366) );
  NAND2_X1 U9690 ( .A1(n10283), .A2(n10415), .ZN(n8359) );
  AOI22_X1 U9691 ( .A1(n11079), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9524), .B2(
        n11067), .ZN(n8358) );
  OAI211_X1 U9692 ( .C1(n9523), .C2(n10287), .A(n8359), .B(n8358), .ZN(n8364)
         );
  NAND2_X1 U9693 ( .A1(n8360), .A2(n9527), .ZN(n8361) );
  NAND2_X1 U9694 ( .A1(n8361), .A2(n10400), .ZN(n8362) );
  OR2_X1 U9695 ( .A1(n8458), .A2(n8362), .ZN(n10417) );
  NOR2_X1 U9696 ( .A1(n10417), .A2(n10219), .ZN(n8363) );
  AOI211_X1 U9697 ( .C1(n10223), .C2(n9527), .A(n8364), .B(n8363), .ZN(n8365)
         );
  OAI211_X1 U9698 ( .C1(n11069), .C2(n10420), .A(n8366), .B(n8365), .ZN(
        P1_U3279) );
  OAI211_X1 U9699 ( .C1(n6606), .C2(n6605), .A(n8367), .B(n9342), .ZN(n8369)
         );
  AOI22_X1 U9700 ( .A1(n9041), .A2(n9339), .B1(n9337), .B2(n9039), .ZN(n8368)
         );
  NAND2_X1 U9701 ( .A1(n8369), .A2(n8368), .ZN(n8498) );
  INV_X1 U9702 ( .A(n8498), .ZN(n8379) );
  NAND2_X1 U9703 ( .A1(n8371), .A2(n8370), .ZN(n8373) );
  AND2_X1 U9704 ( .A1(n8373), .A2(n8372), .ZN(n8375) );
  OAI21_X1 U9705 ( .B1(n8375), .B2(n8942), .A(n8374), .ZN(n8500) );
  INV_X1 U9706 ( .A(n8405), .ZN(n8941) );
  AOI22_X1 U9707 ( .A1(n9315), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n9314), .B2(
        n8411), .ZN(n8376) );
  OAI21_X1 U9708 ( .B1(n8941), .B2(n9317), .A(n8376), .ZN(n8377) );
  AOI21_X1 U9709 ( .B1(n8500), .B2(n9320), .A(n8377), .ZN(n8378) );
  OAI21_X1 U9710 ( .B1(n8379), .B2(n9353), .A(n8378), .ZN(P2_U3221) );
  INV_X1 U9711 ( .A(n8380), .ZN(n8452) );
  AOI21_X1 U9712 ( .B1(P1_DATAO_REG_27__SCAN_IN), .B2(n8610), .A(n8381), .ZN(
        n8382) );
  OAI21_X1 U9713 ( .B1(n8452), .B2(n8667), .A(n8382), .ZN(P2_U3268) );
  NAND2_X1 U9714 ( .A1(n8384), .A2(n8383), .ZN(n8858) );
  XNOR2_X1 U9715 ( .A(n8326), .B(n8858), .ZN(n8476) );
  INV_X1 U9716 ( .A(n8385), .ZN(n8394) );
  NAND2_X1 U9717 ( .A1(n8386), .A2(n8856), .ZN(n8388) );
  NAND2_X1 U9718 ( .A1(n8388), .A2(n8387), .ZN(n8389) );
  XOR2_X1 U9719 ( .A(n8858), .B(n8389), .Z(n8392) );
  OAI22_X1 U9720 ( .A1(n8402), .A2(n9376), .B1(n8390), .B2(n9361), .ZN(n8391)
         );
  AOI21_X1 U9721 ( .B1(n8392), .B2(n9342), .A(n8391), .ZN(n8393) );
  OAI21_X1 U9722 ( .B1(n8394), .B2(n8476), .A(n8393), .ZN(n8477) );
  NAND2_X1 U9723 ( .A1(n8477), .A2(n9377), .ZN(n8400) );
  INV_X1 U9724 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8397) );
  INV_X1 U9725 ( .A(n8395), .ZN(n8396) );
  OAI22_X1 U9726 ( .A1(n9377), .A2(n8397), .B1(n8396), .B2(n9380), .ZN(n8398)
         );
  AOI21_X1 U9727 ( .B1(n8479), .B2(n9364), .A(n8398), .ZN(n8399) );
  OAI211_X1 U9728 ( .C1(n8476), .C2(n8620), .A(n8400), .B(n8399), .ZN(P2_U3223) );
  XNOR2_X1 U9729 ( .A(n8405), .B(n8694), .ZN(n8465) );
  XNOR2_X1 U9730 ( .A(n8465), .B(n8507), .ZN(n8406) );
  OAI211_X1 U9731 ( .C1(n8407), .C2(n8406), .A(n8466), .B(n8824), .ZN(n8413)
         );
  AOI21_X1 U9732 ( .B1(n9041), .B2(n8827), .A(n8408), .ZN(n8409) );
  OAI21_X1 U9733 ( .B1(n9374), .B2(n8829), .A(n8409), .ZN(n8410) );
  AOI21_X1 U9734 ( .B1(n8411), .B2(n8831), .A(n8410), .ZN(n8412) );
  OAI211_X1 U9735 ( .C1(n8941), .C2(n8835), .A(n8413), .B(n8412), .ZN(P2_U3164) );
  INV_X1 U9736 ( .A(n8414), .ZN(n8418) );
  OAI222_X1 U9737 ( .A1(n9513), .A2(n8416), .B1(n8667), .B2(n8418), .C1(n8415), 
        .C2(P2_U3151), .ZN(P2_U3269) );
  OAI222_X1 U9738 ( .A1(n10471), .A2(n10485), .B1(n8633), .B2(n8418), .C1(
        P1_U3086), .C2(n8417), .ZN(P1_U3329) );
  INV_X1 U9739 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n8424) );
  XNOR2_X1 U9740 ( .A(n10049), .B(n8423), .ZN(n10059) );
  INV_X1 U9741 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n8419) );
  AOI22_X1 U9742 ( .A1(n8421), .A2(n8420), .B1(n8434), .B2(n8419), .ZN(n10058)
         );
  NAND2_X1 U9743 ( .A1(n10059), .A2(n10058), .ZN(n10057) );
  OAI21_X1 U9744 ( .B1(n8423), .B2(n8422), .A(n10057), .ZN(n10072) );
  XOR2_X1 U9745 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10063), .Z(n10073) );
  NAND2_X1 U9746 ( .A1(n10072), .A2(n10073), .ZN(n10071) );
  OAI21_X1 U9747 ( .B1(n8425), .B2(n8424), .A(n10071), .ZN(n8426) );
  XNOR2_X1 U9748 ( .A(n8426), .B(n8441), .ZN(n10864) );
  AOI22_X1 U9749 ( .A1(n10865), .A2(n8426), .B1(P1_REG1_REG_15__SCAN_IN), .B2(
        n10864), .ZN(n8429) );
  INV_X1 U9750 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n8427) );
  AOI22_X1 U9751 ( .A1(n10080), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n8427), .B2(
        n8431), .ZN(n8428) );
  NAND2_X1 U9752 ( .A1(n8428), .A2(n8429), .ZN(n10077) );
  OAI21_X1 U9753 ( .B1(n8429), .B2(n8428), .A(n10077), .ZN(n8449) );
  NAND2_X1 U9754 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9592) );
  NAND2_X1 U9755 ( .A1(n10119), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n8430) );
  OAI211_X1 U9756 ( .C1(n10121), .C2(n8431), .A(n9592), .B(n8430), .ZN(n8448)
         );
  INV_X1 U9757 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n8432) );
  XNOR2_X1 U9758 ( .A(n10049), .B(n8432), .ZN(n10056) );
  INV_X1 U9759 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n8433) );
  AOI22_X1 U9760 ( .A1(n8436), .A2(n8435), .B1(n8434), .B2(n8433), .ZN(n10055)
         );
  NAND2_X1 U9761 ( .A1(n10056), .A2(n10055), .ZN(n10054) );
  NAND2_X1 U9762 ( .A1(n10049), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n8437) );
  NAND2_X1 U9763 ( .A1(n10054), .A2(n8437), .ZN(n10069) );
  INV_X1 U9764 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n8438) );
  XNOR2_X1 U9765 ( .A(n10063), .B(n8438), .ZN(n10070) );
  NAND2_X1 U9766 ( .A1(n10069), .A2(n10070), .ZN(n10068) );
  NAND2_X1 U9767 ( .A1(n10063), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n8439) );
  INV_X1 U9768 ( .A(n8440), .ZN(n8442) );
  XOR2_X1 U9769 ( .A(n8441), .B(n8440), .Z(n10873) );
  AOI22_X1 U9770 ( .A1(n10865), .A2(n8442), .B1(P1_REG2_REG_15__SCAN_IN), .B2(
        n10873), .ZN(n8446) );
  NAND2_X1 U9771 ( .A1(n10080), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8443) );
  OAI21_X1 U9772 ( .B1(n10080), .B2(P1_REG2_REG_16__SCAN_IN), .A(n8443), .ZN(
        n8445) );
  NOR2_X1 U9773 ( .A1(n8446), .A2(n8445), .ZN(n10079) );
  AOI211_X1 U9774 ( .C1(n8446), .C2(n8445), .A(n10079), .B(n8444), .ZN(n8447)
         );
  AOI211_X1 U9775 ( .C1(n10877), .C2(n8449), .A(n8448), .B(n8447), .ZN(n8450)
         );
  INV_X1 U9776 ( .A(n8450), .ZN(P1_U3259) );
  OAI222_X1 U9777 ( .A1(P1_U3086), .A2(n8453), .B1(n8633), .B2(n8452), .C1(
        n8451), .C2(n10471), .ZN(P1_U3328) );
  AOI21_X1 U9778 ( .B1(n9789), .B2(n8455), .A(n8454), .ZN(n10414) );
  XNOR2_X1 U9779 ( .A(n8456), .B(n9789), .ZN(n10412) );
  INV_X1 U9780 ( .A(n8457), .ZN(n8490) );
  OAI211_X1 U9781 ( .C1(n10409), .C2(n8458), .A(n8490), .B(n10400), .ZN(n10408) );
  NAND2_X1 U9782 ( .A1(n10283), .A2(n10406), .ZN(n8460) );
  AOI22_X1 U9783 ( .A1(n11069), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9688), .B2(
        n11067), .ZN(n8459) );
  OAI211_X1 U9784 ( .C1(n10389), .C2(n10287), .A(n8460), .B(n8459), .ZN(n8461)
         );
  AOI21_X1 U9785 ( .B1(n9695), .B2(n10223), .A(n8461), .ZN(n8462) );
  OAI21_X1 U9786 ( .B1(n10408), .B2(n10219), .A(n8462), .ZN(n8463) );
  AOI21_X1 U9787 ( .B1(n10412), .B2(n10164), .A(n8463), .ZN(n8464) );
  OAI21_X1 U9788 ( .B1(n10414), .B2(n10309), .A(n8464), .ZN(P1_U3278) );
  INV_X1 U9789 ( .A(n8465), .ZN(n8467) );
  XNOR2_X1 U9790 ( .A(n9462), .B(n8678), .ZN(n8514) );
  XNOR2_X1 U9791 ( .A(n8514), .B(n9039), .ZN(n8468) );
  XNOR2_X1 U9792 ( .A(n8517), .B(n8468), .ZN(n8474) );
  INV_X1 U9793 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n10746) );
  NOR2_X1 U9794 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10746), .ZN(n9061) );
  AOI21_X1 U9795 ( .B1(n9040), .B2(n8827), .A(n9061), .ZN(n8471) );
  NAND2_X1 U9796 ( .A1(n8831), .A2(n8469), .ZN(n8470) );
  OAI211_X1 U9797 ( .C1(n9360), .C2(n8829), .A(n8471), .B(n8470), .ZN(n8472)
         );
  AOI21_X1 U9798 ( .B1(n9462), .B2(n8786), .A(n8472), .ZN(n8473) );
  OAI21_X1 U9799 ( .B1(n8474), .B2(n8788), .A(n8473), .ZN(P2_U3174) );
  INV_X1 U9800 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8481) );
  NOR2_X1 U9801 ( .A1(n8476), .A2(n8475), .ZN(n8478) );
  AOI211_X1 U9802 ( .C1(n9463), .C2(n8479), .A(n8478), .B(n8477), .ZN(n11081)
         );
  OR2_X1 U9803 ( .A1(n11081), .A2(n9465), .ZN(n8480) );
  OAI21_X1 U9804 ( .B1(n9456), .B2(n8481), .A(n8480), .ZN(P2_U3469) );
  INV_X1 U9805 ( .A(n8482), .ZN(n8496) );
  AOI21_X1 U9806 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(n8610), .A(n8483), .ZN(
        n8484) );
  OAI21_X1 U9807 ( .B1(n8496), .B2(n8667), .A(n8484), .ZN(P2_U3267) );
  AOI21_X1 U9808 ( .B1(n8485), .B2(n9771), .A(n11022), .ZN(n8488) );
  OAI22_X1 U9809 ( .A1(n9523), .A2(n10388), .B1(n10297), .B2(n10375), .ZN(
        n8486) );
  AOI21_X1 U9810 ( .B1(n8488), .B2(n8487), .A(n8486), .ZN(n10403) );
  OR2_X1 U9811 ( .A1(n8489), .A2(n9771), .ZN(n10397) );
  NAND3_X1 U9812 ( .A1(n10397), .A2(n10396), .A3(n11075), .ZN(n8495) );
  AOI21_X1 U9813 ( .B1(n10398), .B2(n8490), .A(n8527), .ZN(n10401) );
  AOI22_X1 U9814 ( .A1(n11079), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9591), .B2(
        n11067), .ZN(n8491) );
  OAI21_X1 U9815 ( .B1(n8492), .B2(n11072), .A(n8491), .ZN(n8493) );
  AOI21_X1 U9816 ( .B1(n10401), .B2(n10128), .A(n8493), .ZN(n8494) );
  OAI211_X1 U9817 ( .C1(n11079), .C2(n10403), .A(n8495), .B(n8494), .ZN(
        P1_U3277) );
  OAI222_X1 U9818 ( .A1(P1_U3086), .A2(n8497), .B1(n8633), .B2(n8496), .C1(
        n10768), .C2(n10471), .ZN(P1_U3327) );
  NOR2_X1 U9819 ( .A1(n8941), .A2(n9450), .ZN(n8499) );
  AOI211_X1 U9820 ( .C1(n9414), .C2(n8500), .A(n8499), .B(n8498), .ZN(n11101)
         );
  OR2_X1 U9821 ( .A1(n11101), .A2(n9465), .ZN(n8501) );
  OAI21_X1 U9822 ( .B1(n9456), .B2(n8502), .A(n8501), .ZN(P2_U3471) );
  INV_X1 U9823 ( .A(n8947), .ZN(n8503) );
  XOR2_X1 U9824 ( .A(n8950), .B(n8504), .Z(n9459) );
  XNOR2_X1 U9825 ( .A(n8505), .B(n8950), .ZN(n8506) );
  OAI222_X1 U9826 ( .A1(n9376), .A2(n9360), .B1(n9361), .B2(n8507), .C1(n8506), 
        .C2(n9373), .ZN(n9460) );
  INV_X1 U9827 ( .A(n9462), .ZN(n8510) );
  OAI22_X1 U9828 ( .A1(n8510), .A2(n8509), .B1(n8508), .B2(n9380), .ZN(n8511)
         );
  OAI21_X1 U9829 ( .B1(n9460), .B2(n8511), .A(n9377), .ZN(n8513) );
  NAND2_X1 U9830 ( .A1(n9315), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8512) );
  OAI211_X1 U9831 ( .C1(n9388), .C2(n9459), .A(n8513), .B(n8512), .ZN(P2_U3220) );
  INV_X1 U9832 ( .A(n9385), .ZN(n9451) );
  XNOR2_X1 U9833 ( .A(n9385), .B(n8694), .ZN(n8635) );
  XNOR2_X1 U9834 ( .A(n8635), .B(n9360), .ZN(n8519) );
  NAND2_X1 U9835 ( .A1(n8514), .A2(n9374), .ZN(n8516) );
  INV_X1 U9836 ( .A(n8514), .ZN(n8515) );
  OAI21_X1 U9837 ( .B1(n8519), .B2(n8518), .A(n8822), .ZN(n8520) );
  NAND2_X1 U9838 ( .A1(n8520), .A2(n8824), .ZN(n8524) );
  NOR2_X1 U9839 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10724), .ZN(n9079) );
  AOI21_X1 U9840 ( .B1(n9039), .B2(n8827), .A(n9079), .ZN(n8521) );
  OAI21_X1 U9841 ( .B1(n9375), .B2(n8829), .A(n8521), .ZN(n8522) );
  AOI21_X1 U9842 ( .B1(n9379), .B2(n8831), .A(n8522), .ZN(n8523) );
  OAI211_X1 U9843 ( .C1(n9451), .C2(n8835), .A(n8524), .B(n8523), .ZN(P2_U3155) );
  OAI21_X1 U9844 ( .B1(n8526), .B2(n9792), .A(n8525), .ZN(n10395) );
  INV_X1 U9845 ( .A(n8527), .ZN(n8529) );
  INV_X1 U9846 ( .A(n10301), .ZN(n8528) );
  AOI211_X1 U9847 ( .C1(n8530), .C2(n8529), .A(n10300), .B(n8528), .ZN(n10392)
         );
  NAND2_X1 U9848 ( .A1(n8530), .A2(n10223), .ZN(n8533) );
  AOI22_X1 U9849 ( .A1(n11079), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n11067), 
        .B2(n8531), .ZN(n8532) );
  OAI211_X1 U9850 ( .C1(n10389), .C2(n10143), .A(n8533), .B(n8532), .ZN(n8534)
         );
  AOI21_X1 U9851 ( .B1(n10392), .B2(n11065), .A(n8534), .ZN(n8539) );
  OAI211_X1 U9852 ( .C1(n8536), .C2(n9916), .A(n8535), .B(n10411), .ZN(n8537)
         );
  OAI21_X1 U9853 ( .B1(n6140), .B2(n10375), .A(n8537), .ZN(n10393) );
  NAND2_X1 U9854 ( .A1(n10393), .A2(n10307), .ZN(n8538) );
  OAI211_X1 U9855 ( .C1(n10395), .C2(n10309), .A(n8539), .B(n8538), .ZN(
        P1_U3276) );
  INV_X1 U9856 ( .A(n8540), .ZN(n9516) );
  OAI222_X1 U9857 ( .A1(n10471), .A2(n10763), .B1(n8633), .B2(n9516), .C1(
        n8541), .C2(P1_U3086), .ZN(P1_U3326) );
  NOR2_X1 U9858 ( .A1(n8579), .A2(n8543), .ZN(n8544) );
  INV_X1 U9859 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9067) );
  INV_X1 U9860 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9455) );
  AOI22_X1 U9861 ( .A1(n8558), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n9455), .B2(
        n9081), .ZN(n9074) );
  NOR2_X1 U9862 ( .A1(n9103), .A2(n8545), .ZN(n8546) );
  INV_X1 U9863 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9093) );
  INV_X1 U9864 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8547) );
  AOI22_X1 U9865 ( .A1(n8554), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n8547), .B2(
        n9118), .ZN(n9112) );
  NOR2_X1 U9866 ( .A1(n9138), .A2(n8548), .ZN(n8549) );
  INV_X1 U9867 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9129) );
  NAND2_X1 U9868 ( .A1(n8587), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n9145) );
  OAI21_X1 U9869 ( .B1(n8587), .B2(P2_REG1_REG_18__SCAN_IN), .A(n9145), .ZN(
        n8550) );
  AOI21_X1 U9870 ( .B1(n8551), .B2(n8550), .A(n9147), .ZN(n8594) );
  INV_X1 U9871 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8552) );
  MUX2_X1 U9872 ( .A(n8552), .B(n9129), .S(n8174), .Z(n8569) );
  XNOR2_X1 U9873 ( .A(n8569), .B(n8553), .ZN(n9133) );
  MUX2_X1 U9874 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8174), .Z(n8555) );
  OR2_X1 U9875 ( .A1(n8555), .A2(n9118), .ZN(n8567) );
  XNOR2_X1 U9876 ( .A(n8555), .B(n8554), .ZN(n9114) );
  INV_X1 U9877 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8556) );
  MUX2_X1 U9878 ( .A(n8556), .B(n9093), .S(n8174), .Z(n8557) );
  NAND2_X1 U9879 ( .A1(n8557), .A2(n9103), .ZN(n8566) );
  XOR2_X1 U9880 ( .A(n9103), .B(n8557), .Z(n9106) );
  MUX2_X1 U9881 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8174), .Z(n8559) );
  OR2_X1 U9882 ( .A1(n8559), .A2(n9081), .ZN(n8565) );
  XNOR2_X1 U9883 ( .A(n8559), .B(n8558), .ZN(n9078) );
  MUX2_X1 U9884 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8174), .Z(n8560) );
  OR2_X1 U9885 ( .A1(n8560), .A2(n5497), .ZN(n8564) );
  XNOR2_X1 U9886 ( .A(n8560), .B(n8579), .ZN(n9055) );
  OR2_X1 U9887 ( .A1(n8561), .A2(n8577), .ZN(n8563) );
  NAND2_X1 U9888 ( .A1(n8563), .A2(n8562), .ZN(n9054) );
  NAND2_X1 U9889 ( .A1(n9055), .A2(n9054), .ZN(n9053) );
  NAND2_X1 U9890 ( .A1(n8564), .A2(n9053), .ZN(n9077) );
  NAND2_X1 U9891 ( .A1(n9078), .A2(n9077), .ZN(n9076) );
  NAND2_X1 U9892 ( .A1(n8565), .A2(n9076), .ZN(n9105) );
  NAND2_X1 U9893 ( .A1(n9106), .A2(n9105), .ZN(n9104) );
  NAND2_X1 U9894 ( .A1(n8566), .A2(n9104), .ZN(n9115) );
  NAND2_X1 U9895 ( .A1(n9114), .A2(n9115), .ZN(n9113) );
  NAND2_X1 U9896 ( .A1(n8567), .A2(n9113), .ZN(n9132) );
  NAND2_X1 U9897 ( .A1(n9133), .A2(n9132), .ZN(n9131) );
  INV_X1 U9898 ( .A(n9131), .ZN(n8568) );
  MUX2_X1 U9899 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8174), .Z(n8570) );
  NOR2_X1 U9900 ( .A1(n8571), .A2(n8570), .ZN(n9158) );
  INV_X1 U9901 ( .A(n9158), .ZN(n8572) );
  NAND2_X1 U9902 ( .A1(n8571), .A2(n8570), .ZN(n9156) );
  NAND2_X1 U9903 ( .A1(n8572), .A2(n9156), .ZN(n8573) );
  OAI21_X1 U9904 ( .B1(n8573), .B2(n9045), .A(n10983), .ZN(n8592) );
  NAND3_X1 U9905 ( .A1(n8573), .A2(n11010), .A3(n8587), .ZN(n8574) );
  NAND2_X1 U9906 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_U3151), .ZN(n8805) );
  OAI211_X1 U9907 ( .C1(n8575), .C2(n9095), .A(n8574), .B(n8805), .ZN(n8591)
         );
  NOR2_X1 U9908 ( .A1(n8579), .A2(n8578), .ZN(n8580) );
  INV_X1 U9909 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n9056) );
  NOR2_X1 U9910 ( .A1(n9056), .A2(n9057), .ZN(n9058) );
  INV_X1 U9911 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n9382) );
  NOR2_X1 U9912 ( .A1(n9081), .A2(n9382), .ZN(n8581) );
  AOI21_X1 U9913 ( .B1(n9382), .B2(n9081), .A(n8581), .ZN(n9083) );
  NOR2_X1 U9914 ( .A1(n9084), .A2(n9083), .ZN(n9082) );
  NOR2_X1 U9915 ( .A1(n9103), .A2(n8582), .ZN(n8583) );
  NAND2_X1 U9916 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n9118), .ZN(n8584) );
  OAI21_X1 U9917 ( .B1(n9118), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8584), .ZN(
        n9120) );
  XNOR2_X1 U9918 ( .A(n9138), .B(n8585), .ZN(n9135) );
  NOR2_X1 U9919 ( .A1(n9138), .A2(n8585), .ZN(n8586) );
  NAND2_X1 U9920 ( .A1(n8587), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n9150) );
  OAI21_X1 U9921 ( .B1(n8587), .B2(P2_REG2_REG_18__SCAN_IN), .A(n9150), .ZN(
        n8588) );
  OAI21_X1 U9922 ( .B1(n8594), .B2(n11005), .A(n8593), .ZN(P2_U3200) );
  INV_X1 U9923 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8595) );
  NAND3_X1 U9924 ( .A1(n8595), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n8613) );
  INV_X1 U9925 ( .A(SI_29_), .ZN(n10497) );
  INV_X1 U9926 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8840) );
  INV_X1 U9927 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10760) );
  MUX2_X1 U9928 ( .A(n8840), .B(n10760), .S(n8604), .Z(n8600) );
  NAND2_X1 U9929 ( .A1(n8600), .A2(n10499), .ZN(n8603) );
  INV_X1 U9930 ( .A(n8600), .ZN(n8601) );
  NAND2_X1 U9931 ( .A1(n8601), .A2(SI_30_), .ZN(n8602) );
  NAND2_X1 U9932 ( .A1(n8603), .A2(n8602), .ZN(n8628) );
  MUX2_X1 U9933 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n8604), .Z(n8606) );
  INV_X1 U9934 ( .A(SI_31_), .ZN(n8605) );
  XNOR2_X1 U9935 ( .A(n8606), .B(n8605), .ZN(n8607) );
  NAND2_X1 U9936 ( .A1(n10477), .A2(n8609), .ZN(n8612) );
  NAND2_X1 U9937 ( .A1(n8610), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8611) );
  OAI211_X1 U9938 ( .C1(n6429), .C2(n8613), .A(n8612), .B(n8611), .ZN(P2_U3264) );
  NAND2_X1 U9939 ( .A1(n8614), .A2(n9377), .ZN(n8619) );
  NOR2_X1 U9940 ( .A1(n9380), .A2(n8615), .ZN(n9173) );
  NOR2_X1 U9941 ( .A1(n8616), .A2(n9317), .ZN(n8617) );
  AOI211_X1 U9942 ( .C1(n9315), .C2(P2_REG2_REG_29__SCAN_IN), .A(n9173), .B(
        n8617), .ZN(n8618) );
  OAI211_X1 U9943 ( .C1(n8621), .C2(n8620), .A(n8619), .B(n8618), .ZN(P2_U3204) );
  OAI222_X1 U9944 ( .A1(n8627), .A2(n8622), .B1(n8633), .B2(n8624), .C1(
        P1_U3086), .C2(n10006), .ZN(P1_U3352) );
  OAI222_X1 U9945 ( .A1(n9513), .A2(n8625), .B1(n8667), .B2(n8624), .C1(
        P2_U3151), .C2(n8623), .ZN(P2_U3292) );
  OAI222_X1 U9946 ( .A1(n8627), .A2(n10777), .B1(n8633), .B2(n8626), .C1(n6324), .C2(P1_U3086), .ZN(P1_U3334) );
  INV_X1 U9947 ( .A(n8839), .ZN(n8632) );
  OAI222_X1 U9948 ( .A1(n9513), .A2(n8840), .B1(n8667), .B2(n8632), .C1(
        P2_U3151), .C2(n8630), .ZN(P2_U3265) );
  OAI222_X1 U9949 ( .A1(n10471), .A2(n10581), .B1(n8633), .B2(n8631), .C1(
        P1_U3086), .C2(n6918), .ZN(P1_U3333) );
  OAI222_X1 U9950 ( .A1(P1_U3086), .A2(n8634), .B1(n8633), .B2(n8632), .C1(
        n10760), .C2(n10471), .ZN(P1_U3325) );
  XNOR2_X1 U9951 ( .A(n9448), .B(n8694), .ZN(n8638) );
  XNOR2_X1 U9952 ( .A(n8638), .B(n9375), .ZN(n8825) );
  INV_X1 U9953 ( .A(n8635), .ZN(n8636) );
  NAND2_X1 U9954 ( .A1(n8636), .A2(n9360), .ZN(n8821) );
  XNOR2_X1 U9955 ( .A(n9441), .B(n8694), .ZN(n8639) );
  XNOR2_X1 U9956 ( .A(n8639), .B(n9359), .ZN(n8754) );
  XNOR2_X1 U9957 ( .A(n9437), .B(n8694), .ZN(n8640) );
  XNOR2_X1 U9958 ( .A(n8640), .B(n8966), .ZN(n8762) );
  NAND2_X1 U9959 ( .A1(n8761), .A2(n8762), .ZN(n8800) );
  XNOR2_X1 U9960 ( .A(n9433), .B(n8694), .ZN(n8643) );
  XNOR2_X1 U9961 ( .A(n8643), .B(n8765), .ZN(n8802) );
  INV_X1 U9962 ( .A(n8640), .ZN(n8641) );
  NAND2_X1 U9963 ( .A1(n8641), .A2(n8966), .ZN(n8799) );
  NAND2_X1 U9964 ( .A1(n8800), .A2(n8642), .ZN(n8801) );
  NAND2_X1 U9965 ( .A1(n8643), .A2(n9324), .ZN(n8644) );
  NAND2_X1 U9966 ( .A1(n8801), .A2(n8644), .ZN(n8732) );
  XNOR2_X1 U9967 ( .A(n9291), .B(n8694), .ZN(n8731) );
  NAND2_X1 U9968 ( .A1(n8646), .A2(n9304), .ZN(n8645) );
  XNOR2_X1 U9969 ( .A(n9286), .B(n8694), .ZN(n8647) );
  NAND2_X1 U9970 ( .A1(n8647), .A2(n8742), .ZN(n8649) );
  OAI21_X1 U9971 ( .B1(n8647), .B2(n8742), .A(n8649), .ZN(n8781) );
  NAND2_X1 U9972 ( .A1(n8779), .A2(n8649), .ZN(n8738) );
  XNOR2_X1 U9973 ( .A(n9418), .B(n8694), .ZN(n8650) );
  XNOR2_X1 U9974 ( .A(n8650), .B(n9257), .ZN(n8739) );
  NAND2_X1 U9975 ( .A1(n8738), .A2(n8739), .ZN(n8791) );
  XNOR2_X1 U9976 ( .A(n8982), .B(n8694), .ZN(n8653) );
  XNOR2_X1 U9977 ( .A(n8653), .B(n9243), .ZN(n8793) );
  INV_X1 U9978 ( .A(n8650), .ZN(n8651) );
  NAND2_X1 U9979 ( .A1(n8651), .A2(n9257), .ZN(n8790) );
  NAND2_X1 U9980 ( .A1(n8791), .A2(n8652), .ZN(n8792) );
  NAND2_X1 U9981 ( .A1(n8792), .A2(n8654), .ZN(n8656) );
  XNOR2_X1 U9982 ( .A(n8663), .B(n8694), .ZN(n8655) );
  AOI21_X1 U9983 ( .B1(n8659), .B2(n8658), .A(n5149), .ZN(n8665) );
  AOI22_X1 U9984 ( .A1(n9037), .A2(n8815), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8661) );
  NAND2_X1 U9985 ( .A1(n8831), .A2(n9246), .ZN(n8660) );
  OAI211_X1 U9986 ( .C1(n9243), .C2(n8817), .A(n8661), .B(n8660), .ZN(n8662)
         );
  AOI21_X1 U9987 ( .B1(n8663), .B2(n8786), .A(n8662), .ZN(n8664) );
  OAI21_X1 U9988 ( .B1(n8665), .B2(n8788), .A(n8664), .ZN(P2_U3156) );
  OAI222_X1 U9989 ( .A1(n9513), .A2(n8668), .B1(n8667), .B2(n6458), .C1(
        P2_U3151), .C2(n5128), .ZN(P2_U3293) );
  NOR2_X1 U9990 ( .A1(n8705), .A2(n11072), .ZN(n8672) );
  NAND2_X1 U9991 ( .A1(n10283), .A2(n10326), .ZN(n8670) );
  AOI22_X1 U9992 ( .A1(n11079), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n8713), .B2(
        n11067), .ZN(n8669) );
  OAI211_X1 U9993 ( .C1(n8714), .C2(n10287), .A(n8670), .B(n8669), .ZN(n8671)
         );
  NAND2_X1 U9994 ( .A1(n8674), .A2(n10164), .ZN(n8675) );
  OAI211_X1 U9995 ( .C1(n8677), .C2(n10309), .A(n8676), .B(n8675), .ZN(
        P1_U3265) );
  XNOR2_X1 U9996 ( .A(n8991), .B(n8678), .ZN(n8679) );
  NAND2_X1 U9997 ( .A1(n8679), .A2(n9242), .ZN(n8683) );
  INV_X1 U9998 ( .A(n8679), .ZN(n8680) );
  NAND2_X1 U9999 ( .A1(n8680), .A2(n9037), .ZN(n8681) );
  NAND2_X1 U10000 ( .A1(n8682), .A2(n8770), .ZN(n8772) );
  NAND2_X1 U10001 ( .A1(n8772), .A2(n8683), .ZN(n8747) );
  XNOR2_X1 U10002 ( .A(n8685), .B(n8684), .ZN(n8689) );
  XNOR2_X1 U10003 ( .A(n8689), .B(n9225), .ZN(n8748) );
  INV_X1 U10004 ( .A(n9192), .ZN(n8870) );
  NOR2_X1 U10005 ( .A1(n5657), .A2(n8870), .ZN(n8688) );
  NAND2_X1 U10006 ( .A1(n8686), .A2(n8691), .ZN(n9205) );
  INV_X1 U10007 ( .A(n9205), .ZN(n8687) );
  MUX2_X1 U10008 ( .A(n8688), .B(n8687), .S(n8694), .Z(n8812) );
  INV_X1 U10009 ( .A(n8689), .ZN(n8690) );
  NAND2_X1 U10010 ( .A1(n8690), .A2(n9225), .ZN(n8809) );
  MUX2_X1 U10011 ( .A(n8999), .B(n8691), .S(n8694), .Z(n8692) );
  XNOR2_X1 U10012 ( .A(n9196), .B(n8694), .ZN(n8693) );
  XNOR2_X1 U10013 ( .A(n8693), .B(n9204), .ZN(n8724) );
  AOI22_X1 U10014 ( .A1(n9034), .A2(n8827), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8696) );
  NAND2_X1 U10015 ( .A1(n8831), .A2(n9184), .ZN(n8695) );
  OAI211_X1 U10016 ( .C1(n9179), .C2(n8829), .A(n8696), .B(n8695), .ZN(n8697)
         );
  AOI21_X1 U10017 ( .B1(n8698), .B2(n8786), .A(n8697), .ZN(n8699) );
  OAI21_X1 U10018 ( .B1(n8700), .B2(n8788), .A(n8699), .ZN(P2_U3160) );
  NAND2_X1 U10019 ( .A1(n8702), .A2(n8701), .ZN(n8711) );
  AOI22_X1 U10020 ( .A1(n8718), .A2(n8703), .B1(n7089), .B2(n9995), .ZN(n8709)
         );
  OAI22_X1 U10021 ( .A1(n8705), .A2(n5129), .B1(n10316), .B2(n8704), .ZN(n8707) );
  XNOR2_X1 U10022 ( .A(n8707), .B(n8706), .ZN(n8708) );
  XOR2_X1 U10023 ( .A(n8709), .B(n8708), .Z(n8710) );
  XNOR2_X1 U10024 ( .A(n8711), .B(n8710), .ZN(n8720) );
  OAI22_X1 U10025 ( .A1(n9691), .A2(n10174), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8712), .ZN(n8717) );
  INV_X1 U10026 ( .A(n8713), .ZN(n8715) );
  OAI22_X1 U10027 ( .A1(n9646), .A2(n8715), .B1(n9644), .B2(n8714), .ZN(n8716)
         );
  AOI211_X1 U10028 ( .C1(n8718), .C2(n9694), .A(n8717), .B(n8716), .ZN(n8719)
         );
  OAI21_X1 U10029 ( .B1(n8720), .B2(n9697), .A(n8719), .ZN(P1_U3220) );
  OAI222_X1 U10030 ( .A1(n10471), .A2(n8723), .B1(n8633), .B2(n8722), .C1(
        P1_U3086), .C2(n5130), .ZN(P1_U3336) );
  XNOR2_X1 U10031 ( .A(n8725), .B(n8724), .ZN(n8730) );
  AOI22_X1 U10032 ( .A1(n9035), .A2(n8827), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8727) );
  NAND2_X1 U10033 ( .A1(n8831), .A2(n9197), .ZN(n8726) );
  OAI211_X1 U10034 ( .C1(n9189), .C2(n8829), .A(n8727), .B(n8726), .ZN(n8728)
         );
  AOI21_X1 U10035 ( .B1(n9196), .B2(n8786), .A(n8728), .ZN(n8729) );
  OAI21_X1 U10036 ( .B1(n8730), .B2(n8788), .A(n8729), .ZN(P2_U3154) );
  XNOR2_X1 U10037 ( .A(n8732), .B(n8731), .ZN(n8737) );
  NOR2_X1 U10038 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10729), .ZN(n9162) );
  AOI21_X1 U10039 ( .B1(n9292), .B2(n8815), .A(n9162), .ZN(n8734) );
  NAND2_X1 U10040 ( .A1(n8831), .A2(n9299), .ZN(n8733) );
  OAI211_X1 U10041 ( .C1(n8765), .C2(n8817), .A(n8734), .B(n8733), .ZN(n8735)
         );
  AOI21_X1 U10042 ( .B1(n9298), .B2(n8786), .A(n8735), .ZN(n8736) );
  OAI21_X1 U10043 ( .B1(n8737), .B2(n8788), .A(n8736), .ZN(P2_U3159) );
  OAI21_X1 U10044 ( .B1(n8739), .B2(n8738), .A(n8791), .ZN(n8740) );
  NAND2_X1 U10045 ( .A1(n8740), .A2(n8824), .ZN(n8745) );
  AOI22_X1 U10046 ( .A1(n9266), .A2(n8815), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8741) );
  OAI21_X1 U10047 ( .B1(n8742), .B2(n8817), .A(n8741), .ZN(n8743) );
  AOI21_X1 U10048 ( .B1(n9272), .B2(n8831), .A(n8743), .ZN(n8744) );
  OAI211_X1 U10049 ( .C1(n8746), .C2(n8835), .A(n8745), .B(n8744), .ZN(
        P2_U3163) );
  OAI21_X1 U10050 ( .B1(n8748), .B2(n8747), .A(n8810), .ZN(n8749) );
  NAND2_X1 U10051 ( .A1(n8749), .A2(n8824), .ZN(n8753) );
  AOI22_X1 U10052 ( .A1(n9035), .A2(n8815), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8750) );
  OAI21_X1 U10053 ( .B1(n9242), .B2(n8817), .A(n8750), .ZN(n8751) );
  AOI21_X1 U10054 ( .B1(n9217), .B2(n8831), .A(n8751), .ZN(n8752) );
  OAI211_X1 U10055 ( .C1(n9490), .C2(n8835), .A(n8753), .B(n8752), .ZN(
        P2_U3165) );
  XNOR2_X1 U10056 ( .A(n8755), .B(n8754), .ZN(n8760) );
  INV_X1 U10057 ( .A(n8966), .ZN(n9338) );
  NAND2_X1 U10058 ( .A1(n9338), .A2(n8815), .ZN(n8756) );
  NAND2_X1 U10059 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3151), .ZN(n9116) );
  OAI211_X1 U10060 ( .C1(n9375), .C2(n8817), .A(n8756), .B(n9116), .ZN(n8757)
         );
  AOI21_X1 U10061 ( .B1(n9343), .B2(n8831), .A(n8757), .ZN(n8759) );
  NAND2_X1 U10062 ( .A1(n9441), .A2(n8786), .ZN(n8758) );
  OAI211_X1 U10063 ( .C1(n8760), .C2(n8788), .A(n8759), .B(n8758), .ZN(
        P2_U3166) );
  OAI21_X1 U10064 ( .B1(n8762), .B2(n8761), .A(n8800), .ZN(n8763) );
  NAND2_X1 U10065 ( .A1(n8763), .A2(n8824), .ZN(n8768) );
  AND2_X1 U10066 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9130) );
  AOI21_X1 U10067 ( .B1(n9325), .B2(n8827), .A(n9130), .ZN(n8764) );
  OAI21_X1 U10068 ( .B1(n8765), .B2(n8829), .A(n8764), .ZN(n8766) );
  AOI21_X1 U10069 ( .B1(n9327), .B2(n8831), .A(n8766), .ZN(n8767) );
  OAI211_X1 U10070 ( .C1(n8968), .C2(n8835), .A(n8768), .B(n8767), .ZN(
        P2_U3168) );
  INV_X1 U10071 ( .A(n8769), .ZN(n8771) );
  NOR3_X1 U10072 ( .A1(n5149), .A2(n8771), .A3(n8770), .ZN(n8774) );
  INV_X1 U10073 ( .A(n8772), .ZN(n8773) );
  OAI21_X1 U10074 ( .B1(n8774), .B2(n8773), .A(n8824), .ZN(n8778) );
  INV_X1 U10075 ( .A(n9225), .ZN(n9036) );
  AOI22_X1 U10076 ( .A1(n9036), .A2(n8815), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8775) );
  OAI21_X1 U10077 ( .B1(n9256), .B2(n8817), .A(n8775), .ZN(n8776) );
  AOI21_X1 U10078 ( .B1(n9230), .B2(n8831), .A(n8776), .ZN(n8777) );
  OAI211_X1 U10079 ( .C1(n9494), .C2(n8835), .A(n8778), .B(n8777), .ZN(
        P2_U3169) );
  INV_X1 U10080 ( .A(n8779), .ZN(n8780) );
  AOI21_X1 U10081 ( .B1(n8782), .B2(n8781), .A(n8780), .ZN(n8789) );
  INV_X1 U10082 ( .A(n9257), .ZN(n9278) );
  AOI22_X1 U10083 ( .A1(n9278), .A2(n8815), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8784) );
  NAND2_X1 U10084 ( .A1(n8831), .A2(n9284), .ZN(n8783) );
  OAI211_X1 U10085 ( .C1(n8971), .C2(n8817), .A(n8784), .B(n8783), .ZN(n8785)
         );
  AOI21_X1 U10086 ( .B1(n9422), .B2(n8786), .A(n8785), .ZN(n8787) );
  OAI21_X1 U10087 ( .B1(n8789), .B2(n8788), .A(n8787), .ZN(P2_U3173) );
  INV_X1 U10088 ( .A(n8982), .ZN(n9502) );
  AND2_X1 U10089 ( .A1(n8791), .A2(n8790), .ZN(n8794) );
  OAI211_X1 U10090 ( .C1(n8794), .C2(n8793), .A(n8824), .B(n8792), .ZN(n8798)
         );
  AOI22_X1 U10091 ( .A1(n9278), .A2(n8827), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8795) );
  OAI21_X1 U10092 ( .B1(n9256), .B2(n8829), .A(n8795), .ZN(n8796) );
  AOI21_X1 U10093 ( .B1(n9260), .B2(n8831), .A(n8796), .ZN(n8797) );
  OAI211_X1 U10094 ( .C1(n9502), .C2(n8835), .A(n8798), .B(n8797), .ZN(
        P2_U3175) );
  AND2_X1 U10095 ( .A1(n8800), .A2(n8799), .ZN(n8803) );
  OAI211_X1 U10096 ( .C1(n8803), .C2(n8802), .A(n8824), .B(n8801), .ZN(n8808)
         );
  NAND2_X1 U10097 ( .A1(n9304), .A2(n8815), .ZN(n8804) );
  OAI211_X1 U10098 ( .C1(n8966), .C2(n8817), .A(n8805), .B(n8804), .ZN(n8806)
         );
  AOI21_X1 U10099 ( .B1(n9313), .B2(n8831), .A(n8806), .ZN(n8807) );
  OAI211_X1 U10100 ( .C1(n9318), .C2(n8835), .A(n8808), .B(n8807), .ZN(
        P2_U3178) );
  AND2_X1 U10101 ( .A1(n8810), .A2(n8809), .ZN(n8813) );
  OAI211_X1 U10102 ( .C1(n8813), .C2(n8812), .A(n8824), .B(n8811), .ZN(n8820)
         );
  AOI22_X1 U10103 ( .A1(n9034), .A2(n8815), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8816) );
  OAI21_X1 U10104 ( .B1(n9225), .B2(n8817), .A(n8816), .ZN(n8818) );
  AOI21_X1 U10105 ( .B1(n9206), .B2(n8831), .A(n8818), .ZN(n8819) );
  OAI211_X1 U10106 ( .C1(n9486), .C2(n8835), .A(n8820), .B(n8819), .ZN(
        P2_U3180) );
  INV_X1 U10107 ( .A(n9448), .ZN(n8836) );
  AND2_X1 U10108 ( .A1(n8822), .A2(n8821), .ZN(n8826) );
  OAI211_X1 U10109 ( .C1(n8826), .C2(n8825), .A(n8824), .B(n8823), .ZN(n8834)
         );
  AND2_X1 U10110 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9098) );
  AOI21_X1 U10111 ( .B1(n9038), .B2(n8827), .A(n9098), .ZN(n8828) );
  OAI21_X1 U10112 ( .B1(n9359), .B2(n8829), .A(n8828), .ZN(n8830) );
  AOI21_X1 U10113 ( .B1(n8832), .B2(n8831), .A(n8830), .ZN(n8833) );
  OAI211_X1 U10114 ( .C1(n8836), .C2(n8835), .A(n8834), .B(n8833), .ZN(
        P2_U3181) );
  XNOR2_X1 U10115 ( .A(n9470), .B(n9172), .ZN(n8868) );
  NAND2_X1 U10116 ( .A1(n8839), .A2(n8838), .ZN(n8843) );
  OR2_X1 U10117 ( .A1(n8841), .A2(n8840), .ZN(n8842) );
  NAND2_X1 U10118 ( .A1(n8845), .A2(n8844), .ZN(n8874) );
  AND2_X1 U10119 ( .A1(n8874), .A2(n9011), .ZN(n9016) );
  INV_X1 U10120 ( .A(n9016), .ZN(n8876) );
  NAND2_X1 U10121 ( .A1(n8847), .A2(n8846), .ZN(n9253) );
  INV_X1 U10122 ( .A(n9253), .ZN(n9259) );
  INV_X1 U10123 ( .A(n8987), .ZN(n8848) );
  INV_X1 U10124 ( .A(n9346), .ZN(n9335) );
  NOR4_X1 U10125 ( .A1(n8851), .A2(n8850), .A3(n8885), .A4(n8849), .ZN(n8854)
         );
  NAND4_X1 U10126 ( .A1(n8854), .A2(n8897), .A3(n8853), .A4(n8852), .ZN(n8857)
         );
  NOR4_X1 U10127 ( .A1(n8857), .A2(n8919), .A3(n8856), .A4(n8855), .ZN(n8859)
         );
  NAND4_X1 U10128 ( .A1(n8950), .A2(n8860), .A3(n8859), .A4(n8858), .ZN(n8861)
         );
  NOR4_X1 U10129 ( .A1(n9357), .A2(n9370), .A3(n6605), .A4(n8861), .ZN(n8862)
         );
  NAND4_X1 U10130 ( .A1(n9311), .A2(n9335), .A3(n8862), .A4(n9330), .ZN(n8863)
         );
  NOR2_X1 U10131 ( .A1(n5379), .A2(n8863), .ZN(n8864) );
  NAND4_X1 U10132 ( .A1(n9239), .A2(n9268), .A3(n8864), .A4(n9295), .ZN(n8865)
         );
  NOR4_X1 U10133 ( .A1(n9226), .A2(n9259), .A3(n8865), .A4(n9214), .ZN(n8866)
         );
  NAND4_X1 U10134 ( .A1(n9182), .A2(n9195), .A3(n8866), .A4(n9205), .ZN(n8867)
         );
  NOR4_X1 U10135 ( .A1(n8868), .A2(n8876), .A3(n9019), .A4(n8867), .ZN(n8881)
         );
  INV_X1 U10136 ( .A(n8874), .ZN(n9020) );
  OAI21_X1 U10137 ( .B1(n8845), .B2(n9172), .A(n9470), .ZN(n8879) );
  AOI21_X1 U10138 ( .B1(n8877), .B2(n9172), .A(n9470), .ZN(n8878) );
  INV_X1 U10139 ( .A(n8886), .ZN(n8882) );
  AOI21_X1 U10140 ( .B1(n8884), .B2(n8883), .A(n8882), .ZN(n8893) );
  NOR2_X1 U10141 ( .A1(n8885), .A2(n7476), .ZN(n8887) );
  OAI211_X1 U10142 ( .C1(n8893), .C2(n8887), .A(n9007), .B(n8886), .ZN(n8891)
         );
  INV_X1 U10143 ( .A(n8888), .ZN(n8890) );
  INV_X1 U10144 ( .A(n8889), .ZN(n8907) );
  AOI211_X1 U10145 ( .C1(n8891), .C2(n8892), .A(n8890), .B(n8907), .ZN(n8895)
         );
  AOI21_X1 U10146 ( .B1(n8893), .B2(n8892), .A(n9007), .ZN(n8894) );
  NOR2_X1 U10147 ( .A1(n8895), .A2(n8894), .ZN(n8899) );
  AOI21_X1 U10148 ( .B1(n8900), .B2(n8896), .A(n9007), .ZN(n8898) );
  OAI21_X1 U10149 ( .B1(n8899), .B2(n8898), .A(n8897), .ZN(n8908) );
  INV_X1 U10150 ( .A(n8900), .ZN(n8902) );
  OAI211_X1 U10151 ( .C1(n8908), .C2(n8902), .A(n8909), .B(n8901), .ZN(n8903)
         );
  NAND3_X1 U10152 ( .A1(n8903), .A2(n8905), .A3(n8912), .ZN(n8904) );
  NAND2_X1 U10153 ( .A1(n8904), .A2(n8910), .ZN(n8915) );
  OAI211_X1 U10154 ( .C1(n8908), .C2(n8907), .A(n8906), .B(n8905), .ZN(n8911)
         );
  NAND3_X1 U10155 ( .A1(n8911), .A2(n8910), .A3(n8909), .ZN(n8913) );
  NAND2_X1 U10156 ( .A1(n8913), .A2(n8912), .ZN(n8914) );
  NAND2_X1 U10157 ( .A1(n8920), .A2(n8916), .ZN(n8918) );
  NAND2_X1 U10158 ( .A1(n6817), .A2(n8930), .ZN(n8917) );
  INV_X1 U10159 ( .A(n8920), .ZN(n8923) );
  NOR2_X1 U10160 ( .A1(n8929), .A2(n8921), .ZN(n8922) );
  NOR4_X1 U10161 ( .A1(n8933), .A2(n8923), .A3(n8922), .A4(n8937), .ZN(n8926)
         );
  NAND2_X1 U10162 ( .A1(n8925), .A2(n8924), .ZN(n8939) );
  OAI211_X1 U10163 ( .C1(n8926), .C2(n8939), .A(n8942), .B(n8938), .ZN(n8928)
         );
  AND2_X1 U10164 ( .A1(n8928), .A2(n8927), .ZN(n8945) );
  INV_X1 U10165 ( .A(n8929), .ZN(n8936) );
  OAI21_X1 U10166 ( .B1(n8931), .B2(n9046), .A(n8930), .ZN(n8935) );
  INV_X1 U10167 ( .A(n8932), .ZN(n8934) );
  OAI21_X1 U10168 ( .B1(n8940), .B2(n8939), .A(n8938), .ZN(n8943) );
  AOI22_X1 U10169 ( .A1(n8943), .A2(n8942), .B1(n8941), .B2(n9040), .ZN(n8944)
         );
  INV_X1 U10170 ( .A(n8946), .ZN(n8948) );
  MUX2_X1 U10171 ( .A(n8948), .B(n8947), .S(n9018), .Z(n8949) );
  NAND2_X1 U10172 ( .A1(n8957), .A2(n9451), .ZN(n8952) );
  NAND2_X1 U10173 ( .A1(n8958), .A2(n9360), .ZN(n8951) );
  MUX2_X1 U10174 ( .A(n8952), .B(n8951), .S(n9018), .Z(n8953) );
  AOI21_X1 U10175 ( .B1(n8954), .B2(n9368), .A(n8953), .ZN(n8964) );
  INV_X1 U10176 ( .A(n8955), .ZN(n8956) );
  MUX2_X1 U10177 ( .A(n8958), .B(n8957), .S(n9018), .Z(n8959) );
  NAND3_X1 U10178 ( .A1(n8960), .A2(n9335), .A3(n8959), .ZN(n8963) );
  MUX2_X1 U10179 ( .A(n8961), .B(n9308), .S(n9018), .Z(n8962) );
  OAI21_X1 U10180 ( .B1(n8964), .B2(n8963), .A(n8962), .ZN(n8969) );
  MUX2_X1 U10181 ( .A(n8968), .B(n8966), .S(n9007), .Z(n8965) );
  MUX2_X1 U10182 ( .A(n9007), .B(n8971), .S(n9298), .Z(n8972) );
  OAI21_X1 U10183 ( .B1(n9018), .B2(n9304), .A(n8972), .ZN(n8973) );
  MUX2_X1 U10184 ( .A(n8975), .B(n8974), .S(n9007), .Z(n8976) );
  NAND3_X1 U10185 ( .A1(n8977), .A2(n9268), .A3(n8976), .ZN(n8981) );
  MUX2_X1 U10186 ( .A(n8979), .B(n8978), .S(n9018), .Z(n8980) );
  NAND3_X1 U10187 ( .A1(n8981), .A2(n8980), .A3(n9253), .ZN(n8985) );
  MUX2_X1 U10188 ( .A(n9018), .B(n9243), .S(n8982), .Z(n8983) );
  OAI21_X1 U10189 ( .B1(n9266), .B2(n9007), .A(n8983), .ZN(n8984) );
  NAND3_X1 U10190 ( .A1(n8985), .A2(n9239), .A3(n8984), .ZN(n8990) );
  INV_X1 U10191 ( .A(n9226), .ZN(n9223) );
  INV_X1 U10192 ( .A(n8986), .ZN(n8988) );
  MUX2_X1 U10193 ( .A(n8988), .B(n8987), .S(n9018), .Z(n8989) );
  NAND3_X1 U10194 ( .A1(n8990), .A2(n9223), .A3(n8989), .ZN(n8995) );
  NAND2_X1 U10195 ( .A1(n8991), .A2(n9242), .ZN(n8993) );
  MUX2_X1 U10196 ( .A(n8993), .B(n8992), .S(n9018), .Z(n8994) );
  AOI21_X1 U10197 ( .B1(n8995), .B2(n8994), .A(n9214), .ZN(n9002) );
  MUX2_X1 U10198 ( .A(n8997), .B(n8996), .S(n9007), .Z(n8998) );
  NAND2_X1 U10199 ( .A1(n9205), .A2(n8998), .ZN(n9001) );
  MUX2_X1 U10200 ( .A(n8999), .B(n9192), .S(n9018), .Z(n9000) );
  OAI211_X1 U10201 ( .C1(n9002), .C2(n9001), .A(n9195), .B(n9000), .ZN(n9006)
         );
  MUX2_X1 U10202 ( .A(n9004), .B(n9003), .S(n9007), .Z(n9005) );
  INV_X1 U10203 ( .A(n9009), .ZN(n9010) );
  MUX2_X1 U10204 ( .A(n9189), .B(n9478), .S(n9007), .Z(n9008) );
  INV_X1 U10205 ( .A(n9017), .ZN(n9012) );
  NAND2_X1 U10206 ( .A1(n9012), .A2(n9011), .ZN(n9015) );
  INV_X1 U10207 ( .A(n9013), .ZN(n9014) );
  NOR2_X1 U10208 ( .A1(n9019), .A2(n9018), .ZN(n9021) );
  XNOR2_X1 U10209 ( .A(n9026), .B(n5535), .ZN(n9032) );
  NOR3_X1 U10210 ( .A1(n9027), .A2(n6837), .A3(n7193), .ZN(n9030) );
  OAI21_X1 U10211 ( .B1(n9031), .B2(n9028), .A(P2_B_REG_SCAN_IN), .ZN(n9029)
         );
  OAI22_X1 U10212 ( .A1(n9032), .A2(n9031), .B1(n9030), .B2(n9029), .ZN(
        P2_U3296) );
  MUX2_X1 U10213 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n9033), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U10214 ( .A(n9034), .B(P2_DATAO_REG_27__SCAN_IN), .S(n9045), .Z(
        P2_U3518) );
  MUX2_X1 U10215 ( .A(n9035), .B(P2_DATAO_REG_26__SCAN_IN), .S(n9045), .Z(
        P2_U3517) );
  MUX2_X1 U10216 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n9036), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10217 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n9037), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10218 ( .A(n9266), .B(P2_DATAO_REG_22__SCAN_IN), .S(n9045), .Z(
        P2_U3513) );
  MUX2_X1 U10219 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n9278), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10220 ( .A(n9292), .B(P2_DATAO_REG_20__SCAN_IN), .S(n9045), .Z(
        P2_U3511) );
  MUX2_X1 U10221 ( .A(n9304), .B(P2_DATAO_REG_19__SCAN_IN), .S(n9045), .Z(
        P2_U3510) );
  MUX2_X1 U10222 ( .A(n9324), .B(P2_DATAO_REG_18__SCAN_IN), .S(n9045), .Z(
        P2_U3509) );
  MUX2_X1 U10223 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n9338), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10224 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n9325), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U10225 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n9340), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U10226 ( .A(n9038), .B(P2_DATAO_REG_14__SCAN_IN), .S(n9045), .Z(
        P2_U3505) );
  MUX2_X1 U10227 ( .A(n9039), .B(P2_DATAO_REG_13__SCAN_IN), .S(n9045), .Z(
        P2_U3504) );
  MUX2_X1 U10228 ( .A(n9040), .B(P2_DATAO_REG_12__SCAN_IN), .S(n9045), .Z(
        P2_U3503) );
  MUX2_X1 U10229 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n9041), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U10230 ( .A(n9042), .B(P2_DATAO_REG_10__SCAN_IN), .S(n9045), .Z(
        P2_U3501) );
  MUX2_X1 U10231 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n9043), .S(P2_U3893), .Z(
        P2_U3500) );
  MUX2_X1 U10232 ( .A(n9044), .B(P2_DATAO_REG_8__SCAN_IN), .S(n9045), .Z(
        P2_U3499) );
  MUX2_X1 U10233 ( .A(n9046), .B(P2_DATAO_REG_7__SCAN_IN), .S(n9045), .Z(
        P2_U3498) );
  MUX2_X1 U10234 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n6520), .S(P2_U3893), .Z(
        P2_U3497) );
  MUX2_X1 U10235 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n9047), .S(P2_U3893), .Z(
        P2_U3496) );
  MUX2_X1 U10236 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n9048), .S(P2_U3893), .Z(
        P2_U3495) );
  MUX2_X1 U10237 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n9049), .S(P2_U3893), .Z(
        P2_U3494) );
  MUX2_X1 U10238 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n9050), .S(P2_U3893), .Z(
        P2_U3493) );
  MUX2_X1 U10239 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n9051), .S(P2_U3893), .Z(
        P2_U3492) );
  MUX2_X1 U10240 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n9052), .S(P2_U3893), .Z(
        P2_U3491) );
  OAI21_X1 U10241 ( .B1(n9055), .B2(n9054), .A(n9053), .ZN(n9071) );
  NAND2_X1 U10242 ( .A1(n9057), .A2(n9056), .ZN(n9060) );
  INV_X1 U10243 ( .A(n9058), .ZN(n9059) );
  NAND2_X1 U10244 ( .A1(n9060), .A2(n9059), .ZN(n9062) );
  AOI21_X1 U10245 ( .B1(n10968), .B2(n9062), .A(n9061), .ZN(n9064) );
  NAND2_X1 U10246 ( .A1(n10996), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n9063) );
  OAI211_X1 U10247 ( .C1(n10983), .C2(n5497), .A(n9064), .B(n9063), .ZN(n9070)
         );
  AOI21_X1 U10248 ( .B1(n9067), .B2(n9066), .A(n9065), .ZN(n9068) );
  NOR2_X1 U10249 ( .A1(n9068), .A2(n11005), .ZN(n9069) );
  AOI211_X1 U10250 ( .C1(n11010), .C2(n9071), .A(n9070), .B(n9069), .ZN(n9072)
         );
  INV_X1 U10251 ( .A(n9072), .ZN(P2_U3195) );
  AOI21_X1 U10252 ( .B1(n9075), .B2(n9074), .A(n9073), .ZN(n9090) );
  OAI21_X1 U10253 ( .B1(n9078), .B2(n9077), .A(n9076), .ZN(n9088) );
  AOI21_X1 U10254 ( .B1(n10996), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n9079), .ZN(
        n9080) );
  OAI21_X1 U10255 ( .B1(n9081), .B2(n10983), .A(n9080), .ZN(n9087) );
  AOI21_X1 U10256 ( .B1(n9084), .B2(n9083), .A(n9082), .ZN(n9085) );
  NOR2_X1 U10257 ( .A1(n9085), .A2(n11014), .ZN(n9086) );
  AOI211_X1 U10258 ( .C1(n11010), .C2(n9088), .A(n9087), .B(n9086), .ZN(n9089)
         );
  OAI21_X1 U10259 ( .B1(n9090), .B2(n11005), .A(n9089), .ZN(P2_U3196) );
  AOI21_X1 U10260 ( .B1(n9093), .B2(n9092), .A(n9091), .ZN(n9110) );
  NOR2_X1 U10261 ( .A1(n9095), .A2(n9094), .ZN(n9102) );
  AOI21_X1 U10262 ( .B1(n9097), .B2(n8556), .A(n9096), .ZN(n9100) );
  INV_X1 U10263 ( .A(n9098), .ZN(n9099) );
  OAI21_X1 U10264 ( .B1(n11014), .B2(n9100), .A(n9099), .ZN(n9101) );
  AOI211_X1 U10265 ( .C1(n10997), .C2(n9103), .A(n9102), .B(n9101), .ZN(n9109)
         );
  OAI21_X1 U10266 ( .B1(n9106), .B2(n9105), .A(n9104), .ZN(n9107) );
  NAND2_X1 U10267 ( .A1(n9107), .A2(n11010), .ZN(n9108) );
  OAI211_X1 U10268 ( .C1(n9110), .C2(n11005), .A(n9109), .B(n9108), .ZN(
        P2_U3197) );
  AOI21_X1 U10269 ( .B1(n5169), .B2(n9112), .A(n9111), .ZN(n9126) );
  OAI21_X1 U10270 ( .B1(n9115), .B2(n9114), .A(n9113), .ZN(n9124) );
  NAND2_X1 U10271 ( .A1(n10996), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n9117) );
  OAI211_X1 U10272 ( .C1(n10983), .C2(n9118), .A(n9117), .B(n9116), .ZN(n9123)
         );
  AOI21_X1 U10273 ( .B1(n5171), .B2(n9120), .A(n9119), .ZN(n9121) );
  NOR2_X1 U10274 ( .A1(n9121), .A2(n11014), .ZN(n9122) );
  AOI211_X1 U10275 ( .C1(n11010), .C2(n9124), .A(n9123), .B(n9122), .ZN(n9125)
         );
  OAI21_X1 U10276 ( .B1(n9126), .B2(n11005), .A(n9125), .ZN(P2_U3198) );
  AOI21_X1 U10277 ( .B1(n9129), .B2(n9128), .A(n9127), .ZN(n9144) );
  AOI21_X1 U10278 ( .B1(n10996), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n9130), .ZN(
        n9142) );
  OAI21_X1 U10279 ( .B1(n9133), .B2(n9132), .A(n9131), .ZN(n9134) );
  NAND2_X1 U10280 ( .A1(n9134), .A2(n11010), .ZN(n9141) );
  AND2_X1 U10281 ( .A1(n9135), .A2(n8552), .ZN(n9136) );
  OAI21_X1 U10282 ( .B1(n9137), .B2(n9136), .A(n10968), .ZN(n9140) );
  NAND2_X1 U10283 ( .A1(n10997), .A2(n9138), .ZN(n9139) );
  AND4_X1 U10284 ( .A1(n9142), .A2(n9141), .A3(n9140), .A4(n9139), .ZN(n9143)
         );
  OAI21_X1 U10285 ( .B1(n9144), .B2(n11005), .A(n9143), .ZN(P2_U3199) );
  INV_X1 U10286 ( .A(n9145), .ZN(n9146) );
  INV_X1 U10287 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9430) );
  XNOR2_X1 U10288 ( .A(n9151), .B(n9430), .ZN(n9154) );
  INV_X1 U10289 ( .A(n9154), .ZN(n9148) );
  XNOR2_X1 U10290 ( .A(n9149), .B(n9148), .ZN(n9169) );
  INV_X1 U10291 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n9152) );
  MUX2_X1 U10292 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n9152), .S(n9151), .Z(n9155) );
  XNOR2_X1 U10293 ( .A(n9153), .B(n9155), .ZN(n9167) );
  MUX2_X1 U10294 ( .A(n9155), .B(n9154), .S(n8174), .Z(n9160) );
  OAI21_X1 U10295 ( .B1(n9158), .B2(n9157), .A(n9156), .ZN(n9159) );
  XOR2_X1 U10296 ( .A(n9160), .B(n9159), .Z(n9165) );
  NOR2_X1 U10297 ( .A1(n10983), .A2(n5535), .ZN(n9161) );
  AOI211_X1 U10298 ( .C1(P2_ADDR_REG_19__SCAN_IN), .C2(n10996), .A(n9162), .B(
        n9161), .ZN(n9163) );
  OAI21_X1 U10299 ( .B1(n9165), .B2(n9164), .A(n9163), .ZN(n9166) );
  AOI21_X1 U10300 ( .B1(n9167), .B2(n10968), .A(n9166), .ZN(n9168) );
  OAI21_X1 U10301 ( .B1(n9169), .B2(n11005), .A(n9168), .ZN(P2_U3201) );
  INV_X1 U10302 ( .A(n9170), .ZN(n9171) );
  NAND2_X1 U10303 ( .A1(n9172), .A2(n9171), .ZN(n9468) );
  INV_X1 U10304 ( .A(n9468), .ZN(n9174) );
  NOR3_X1 U10305 ( .A1(n9174), .A2(n9315), .A3(n9173), .ZN(n9177) );
  NOR2_X1 U10306 ( .A1(n9377), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9175) );
  OAI22_X1 U10307 ( .A1(n9470), .A2(n9317), .B1(n9177), .B2(n9175), .ZN(
        P2_U3202) );
  NOR2_X1 U10308 ( .A1(n9377), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n9176) );
  OAI22_X1 U10309 ( .A1(n9474), .A2(n9317), .B1(n9177), .B2(n9176), .ZN(
        P2_U3203) );
  XNOR2_X1 U10310 ( .A(n9178), .B(n9182), .ZN(n9181) );
  OAI22_X1 U10311 ( .A1(n9204), .A2(n9361), .B1(n9179), .B2(n9376), .ZN(n9180)
         );
  AOI22_X1 U10312 ( .A1(n9315), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n9314), .B2(
        n9184), .ZN(n9185) );
  OAI21_X1 U10313 ( .B1(n9478), .B2(n9317), .A(n9185), .ZN(n9186) );
  AOI21_X1 U10314 ( .B1(n5124), .B2(n9320), .A(n9186), .ZN(n9187) );
  OAI21_X1 U10315 ( .B1(n9392), .B2(n9353), .A(n9187), .ZN(P2_U3205) );
  XOR2_X1 U10316 ( .A(n9195), .B(n9188), .Z(n9191) );
  OAI22_X1 U10317 ( .A1(n9213), .A2(n9361), .B1(n9189), .B2(n9376), .ZN(n9190)
         );
  AOI21_X1 U10318 ( .B1(n9191), .B2(n9342), .A(n9190), .ZN(n9393) );
  NAND2_X1 U10319 ( .A1(n9193), .A2(n9192), .ZN(n9194) );
  XOR2_X1 U10320 ( .A(n9195), .B(n9194), .Z(n9394) );
  INV_X1 U10321 ( .A(n9394), .ZN(n9200) );
  INV_X1 U10322 ( .A(n9196), .ZN(n9482) );
  AOI22_X1 U10323 ( .A1(n9315), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n9314), .B2(
        n9197), .ZN(n9198) );
  OAI21_X1 U10324 ( .B1(n9482), .B2(n9317), .A(n9198), .ZN(n9199) );
  AOI21_X1 U10325 ( .B1(n9200), .B2(n9320), .A(n9199), .ZN(n9201) );
  OAI21_X1 U10326 ( .B1(n9393), .B2(n9353), .A(n9201), .ZN(P2_U3206) );
  XNOR2_X1 U10327 ( .A(n9202), .B(n9205), .ZN(n9203) );
  OAI222_X1 U10328 ( .A1(n9361), .A2(n9225), .B1(n9376), .B2(n9204), .C1(n9203), .C2(n9373), .ZN(n9397) );
  INV_X1 U10329 ( .A(n9397), .ZN(n9210) );
  XNOR2_X1 U10330 ( .A(n8869), .B(n9205), .ZN(n9398) );
  AOI22_X1 U10331 ( .A1(n9315), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n9314), .B2(
        n9206), .ZN(n9207) );
  OAI21_X1 U10332 ( .B1(n9486), .B2(n9317), .A(n9207), .ZN(n9208) );
  AOI21_X1 U10333 ( .B1(n9398), .B2(n9320), .A(n9208), .ZN(n9209) );
  OAI21_X1 U10334 ( .B1(n9210), .B2(n9353), .A(n9209), .ZN(P2_U3207) );
  XOR2_X1 U10335 ( .A(n9214), .B(n9211), .Z(n9212) );
  OAI222_X1 U10336 ( .A1(n9376), .A2(n9213), .B1(n9361), .B2(n9242), .C1(n9373), .C2(n9212), .ZN(n9401) );
  INV_X1 U10337 ( .A(n9401), .ZN(n9221) );
  XNOR2_X1 U10338 ( .A(n9215), .B(n9214), .ZN(n9402) );
  NAND2_X1 U10339 ( .A1(n9377), .A2(n9216), .ZN(n9378) );
  AOI22_X1 U10340 ( .A1(n9315), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n9314), .B2(
        n9217), .ZN(n9218) );
  OAI21_X1 U10341 ( .B1(n9490), .B2(n9378), .A(n9218), .ZN(n9219) );
  AOI21_X1 U10342 ( .B1(n9402), .B2(n9320), .A(n9219), .ZN(n9220) );
  OAI21_X1 U10343 ( .B1(n9221), .B2(n9353), .A(n9220), .ZN(P2_U3208) );
  XNOR2_X1 U10344 ( .A(n9222), .B(n9223), .ZN(n9224) );
  OAI222_X1 U10345 ( .A1(n9376), .A2(n9225), .B1(n9361), .B2(n9256), .C1(n9224), .C2(n9373), .ZN(n9405) );
  NAND2_X1 U10346 ( .A1(n9227), .A2(n9226), .ZN(n9228) );
  AND2_X1 U10347 ( .A1(n9229), .A2(n9228), .ZN(n9406) );
  NAND2_X1 U10348 ( .A1(n9406), .A2(n9320), .ZN(n9232) );
  AOI22_X1 U10349 ( .A1(n9315), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n9314), .B2(
        n9230), .ZN(n9231) );
  OAI211_X1 U10350 ( .C1(n9494), .C2(n9378), .A(n9232), .B(n9231), .ZN(n9233)
         );
  AOI21_X1 U10351 ( .B1(n9405), .B2(n9377), .A(n9233), .ZN(n9234) );
  INV_X1 U10352 ( .A(n9234), .ZN(P2_U3209) );
  NAND2_X1 U10353 ( .A1(n9235), .A2(n9236), .ZN(n9238) );
  NAND2_X1 U10354 ( .A1(n9238), .A2(n9237), .ZN(n9240) );
  XNOR2_X1 U10355 ( .A(n9240), .B(n9239), .ZN(n9241) );
  OAI222_X1 U10356 ( .A1(n9361), .A2(n9243), .B1(n9376), .B2(n9242), .C1(n9373), .C2(n9241), .ZN(n9409) );
  INV_X1 U10357 ( .A(n9409), .ZN(n9250) );
  XNOR2_X1 U10358 ( .A(n9245), .B(n9244), .ZN(n9410) );
  AOI22_X1 U10359 ( .A1(n9315), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n9314), .B2(
        n9246), .ZN(n9247) );
  OAI21_X1 U10360 ( .B1(n9498), .B2(n9317), .A(n9247), .ZN(n9248) );
  AOI21_X1 U10361 ( .B1(n9410), .B2(n9320), .A(n9248), .ZN(n9249) );
  OAI21_X1 U10362 ( .B1(n9250), .B2(n9315), .A(n9249), .ZN(P2_U3210) );
  NAND2_X1 U10363 ( .A1(n9235), .A2(n9265), .ZN(n9252) );
  NAND2_X1 U10364 ( .A1(n9252), .A2(n9251), .ZN(n9254) );
  XNOR2_X1 U10365 ( .A(n9254), .B(n9253), .ZN(n9255) );
  OAI222_X1 U10366 ( .A1(n9361), .A2(n9257), .B1(n9376), .B2(n9256), .C1(n9255), .C2(n9373), .ZN(n9413) );
  INV_X1 U10367 ( .A(n9413), .ZN(n9264) );
  XNOR2_X1 U10368 ( .A(n9258), .B(n9259), .ZN(n9415) );
  AOI22_X1 U10369 ( .A1(n9315), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9314), .B2(
        n9260), .ZN(n9261) );
  OAI21_X1 U10370 ( .B1(n9502), .B2(n9317), .A(n9261), .ZN(n9262) );
  AOI21_X1 U10371 ( .B1(n9415), .B2(n9320), .A(n9262), .ZN(n9263) );
  OAI21_X1 U10372 ( .B1(n9264), .B2(n9353), .A(n9263), .ZN(P2_U3211) );
  XNOR2_X1 U10373 ( .A(n9235), .B(n9265), .ZN(n9267) );
  AOI222_X1 U10374 ( .A1(n9342), .A2(n9267), .B1(n9292), .B2(n9339), .C1(n9266), .C2(n9337), .ZN(n9420) );
  OR2_X1 U10375 ( .A1(n9269), .A2(n9268), .ZN(n9270) );
  NAND2_X1 U10376 ( .A1(n9271), .A2(n9270), .ZN(n9421) );
  AOI22_X1 U10377 ( .A1(n9315), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n9314), .B2(
        n9272), .ZN(n9274) );
  NAND2_X1 U10378 ( .A1(n9418), .A2(n9364), .ZN(n9273) );
  OAI211_X1 U10379 ( .C1(n9421), .C2(n9388), .A(n9274), .B(n9273), .ZN(n9275)
         );
  INV_X1 U10380 ( .A(n9275), .ZN(n9276) );
  OAI21_X1 U10381 ( .B1(n9420), .B2(n9353), .A(n9276), .ZN(P2_U3212) );
  OAI21_X1 U10382 ( .B1(n5206), .B2(n5379), .A(n9277), .ZN(n9279) );
  AOI222_X1 U10383 ( .A1(n9342), .A2(n9279), .B1(n9304), .B2(n9339), .C1(n9278), .C2(n9337), .ZN(n9424) );
  OR2_X1 U10384 ( .A1(n9281), .A2(n9280), .ZN(n9282) );
  NAND2_X1 U10385 ( .A1(n9283), .A2(n9282), .ZN(n9425) );
  INV_X1 U10386 ( .A(n9425), .ZN(n9288) );
  AOI22_X1 U10387 ( .A1(n9315), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9314), .B2(
        n9284), .ZN(n9285) );
  OAI21_X1 U10388 ( .B1(n9286), .B2(n9317), .A(n9285), .ZN(n9287) );
  AOI21_X1 U10389 ( .B1(n9288), .B2(n9320), .A(n9287), .ZN(n9289) );
  OAI21_X1 U10390 ( .B1(n9424), .B2(n9353), .A(n9289), .ZN(P2_U3213) );
  OAI211_X1 U10391 ( .C1(n5209), .C2(n9291), .A(n9290), .B(n9342), .ZN(n9294)
         );
  AOI22_X1 U10392 ( .A1(n9337), .A2(n9292), .B1(n9324), .B2(n9339), .ZN(n9293)
         );
  NAND2_X1 U10393 ( .A1(n9294), .A2(n9293), .ZN(n9427) );
  NOR2_X1 U10394 ( .A1(n9296), .A2(n9295), .ZN(n9426) );
  INV_X1 U10395 ( .A(n9428), .ZN(n9297) );
  NOR3_X1 U10396 ( .A1(n9426), .A2(n9297), .A3(n9388), .ZN(n9302) );
  INV_X1 U10397 ( .A(n9298), .ZN(n9509) );
  AOI22_X1 U10398 ( .A1(n9315), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n9314), .B2(
        n9299), .ZN(n9300) );
  OAI21_X1 U10399 ( .B1(n9509), .B2(n9317), .A(n9300), .ZN(n9301) );
  AOI211_X1 U10400 ( .C1(n9427), .C2(n9377), .A(n9302), .B(n9301), .ZN(n9303)
         );
  INV_X1 U10401 ( .A(n9303), .ZN(P2_U3214) );
  XOR2_X1 U10402 ( .A(n5195), .B(n9311), .Z(n9305) );
  AOI222_X1 U10403 ( .A1(n9342), .A2(n9305), .B1(n9304), .B2(n9337), .C1(n9338), .C2(n9339), .ZN(n9435) );
  NAND2_X1 U10404 ( .A1(n9306), .A2(n9307), .ZN(n9348) );
  NAND2_X1 U10405 ( .A1(n9348), .A2(n9308), .ZN(n9331) );
  NAND2_X1 U10406 ( .A1(n9331), .A2(n9330), .ZN(n9329) );
  NAND2_X1 U10407 ( .A1(n9329), .A2(n9309), .ZN(n9312) );
  OAI21_X1 U10408 ( .B1(n9312), .B2(n9311), .A(n9310), .ZN(n9436) );
  INV_X1 U10409 ( .A(n9436), .ZN(n9321) );
  AOI22_X1 U10410 ( .A1(n9315), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9314), .B2(
        n9313), .ZN(n9316) );
  OAI21_X1 U10411 ( .B1(n9318), .B2(n9317), .A(n9316), .ZN(n9319) );
  AOI21_X1 U10412 ( .B1(n9321), .B2(n9320), .A(n9319), .ZN(n9322) );
  OAI21_X1 U10413 ( .B1(n9435), .B2(n9353), .A(n9322), .ZN(P2_U3215) );
  XNOR2_X1 U10414 ( .A(n9323), .B(n9330), .ZN(n9326) );
  AOI222_X1 U10415 ( .A1(n9342), .A2(n9326), .B1(n9325), .B2(n9339), .C1(n9324), .C2(n9337), .ZN(n9439) );
  INV_X1 U10416 ( .A(n9327), .ZN(n9328) );
  OAI22_X1 U10417 ( .A1(n9377), .A2(n8552), .B1(n9328), .B2(n9380), .ZN(n9333)
         );
  OAI21_X1 U10418 ( .B1(n9331), .B2(n9330), .A(n9329), .ZN(n9440) );
  NOR2_X1 U10419 ( .A1(n9440), .A2(n9388), .ZN(n9332) );
  AOI211_X1 U10420 ( .C1(n9364), .C2(n9437), .A(n9333), .B(n9332), .ZN(n9334)
         );
  OAI21_X1 U10421 ( .B1(n9439), .B2(n9353), .A(n9334), .ZN(P2_U3216) );
  XNOR2_X1 U10422 ( .A(n9336), .B(n9335), .ZN(n9341) );
  AOI222_X1 U10423 ( .A1(n9342), .A2(n9341), .B1(n9340), .B2(n9339), .C1(n9338), .C2(n9337), .ZN(n9443) );
  INV_X1 U10424 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n9345) );
  INV_X1 U10425 ( .A(n9343), .ZN(n9344) );
  OAI22_X1 U10426 ( .A1(n9377), .A2(n9345), .B1(n9344), .B2(n9380), .ZN(n9351)
         );
  INV_X1 U10427 ( .A(n9306), .ZN(n9354) );
  OAI21_X1 U10428 ( .B1(n9354), .B2(n9347), .A(n9346), .ZN(n9349) );
  NAND2_X1 U10429 ( .A1(n9349), .A2(n9348), .ZN(n9444) );
  NOR2_X1 U10430 ( .A1(n9444), .A2(n9388), .ZN(n9350) );
  AOI211_X1 U10431 ( .C1(n9364), .C2(n9441), .A(n9351), .B(n9350), .ZN(n9352)
         );
  OAI21_X1 U10432 ( .B1(n9443), .B2(n9353), .A(n9352), .ZN(P2_U3217) );
  AOI21_X1 U10433 ( .B1(n9357), .B2(n9355), .A(n9354), .ZN(n9445) );
  XNOR2_X1 U10434 ( .A(n9356), .B(n9357), .ZN(n9358) );
  OAI222_X1 U10435 ( .A1(n9361), .A2(n9360), .B1(n9376), .B2(n9359), .C1(n9358), .C2(n9373), .ZN(n9446) );
  NAND2_X1 U10436 ( .A1(n9446), .A2(n9377), .ZN(n9366) );
  OAI22_X1 U10437 ( .A1(n9377), .A2(n8556), .B1(n9362), .B2(n9380), .ZN(n9363)
         );
  AOI21_X1 U10438 ( .B1(n9448), .B2(n9364), .A(n9363), .ZN(n9365) );
  OAI211_X1 U10439 ( .C1(n9388), .C2(n9445), .A(n9366), .B(n9365), .ZN(
        P2_U3218) );
  OAI21_X1 U10440 ( .B1(n9369), .B2(n9368), .A(n9367), .ZN(n9452) );
  XNOR2_X1 U10441 ( .A(n9371), .B(n9370), .ZN(n9372) );
  OAI222_X1 U10442 ( .A1(n9376), .A2(n9375), .B1(n9361), .B2(n9374), .C1(n9373), .C2(n9372), .ZN(n9454) );
  NAND2_X1 U10443 ( .A1(n9454), .A2(n9377), .ZN(n9387) );
  INV_X1 U10444 ( .A(n9378), .ZN(n9384) );
  INV_X1 U10445 ( .A(n9379), .ZN(n9381) );
  OAI22_X1 U10446 ( .A1(n9377), .A2(n9382), .B1(n9381), .B2(n9380), .ZN(n9383)
         );
  AOI21_X1 U10447 ( .B1(n9385), .B2(n9384), .A(n9383), .ZN(n9386) );
  OAI211_X1 U10448 ( .C1(n9388), .C2(n9452), .A(n9387), .B(n9386), .ZN(
        P2_U3219) );
  NOR2_X1 U10449 ( .A1(n9468), .A2(n9465), .ZN(n9390) );
  AOI21_X1 U10450 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n9465), .A(n9390), .ZN(
        n9389) );
  OAI21_X1 U10451 ( .B1(n9470), .B2(n9432), .A(n9389), .ZN(P2_U3490) );
  AOI21_X1 U10452 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(n9465), .A(n9390), .ZN(
        n9391) );
  OAI21_X1 U10453 ( .B1(n9474), .B2(n9432), .A(n9391), .ZN(P2_U3489) );
  OAI21_X1 U10454 ( .B1(n9458), .B2(n9394), .A(n9393), .ZN(n9479) );
  MUX2_X1 U10455 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9479), .S(n9456), .Z(n9395) );
  INV_X1 U10456 ( .A(n9395), .ZN(n9396) );
  OAI21_X1 U10457 ( .B1(n9482), .B2(n9432), .A(n9396), .ZN(P2_U3486) );
  INV_X1 U10458 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9399) );
  AOI21_X1 U10459 ( .B1(n9414), .B2(n9398), .A(n9397), .ZN(n9483) );
  MUX2_X1 U10460 ( .A(n9399), .B(n9483), .S(n9456), .Z(n9400) );
  OAI21_X1 U10461 ( .B1(n9486), .B2(n9432), .A(n9400), .ZN(P2_U3485) );
  INV_X1 U10462 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9403) );
  AOI21_X1 U10463 ( .B1(n9414), .B2(n9402), .A(n9401), .ZN(n9487) );
  MUX2_X1 U10464 ( .A(n9403), .B(n9487), .S(n9456), .Z(n9404) );
  OAI21_X1 U10465 ( .B1(n9490), .B2(n9432), .A(n9404), .ZN(P2_U3484) );
  INV_X1 U10466 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9407) );
  AOI21_X1 U10467 ( .B1(n9406), .B2(n9414), .A(n9405), .ZN(n9491) );
  MUX2_X1 U10468 ( .A(n9407), .B(n9491), .S(n9456), .Z(n9408) );
  OAI21_X1 U10469 ( .B1(n9494), .B2(n9432), .A(n9408), .ZN(P2_U3483) );
  INV_X1 U10470 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9411) );
  AOI21_X1 U10471 ( .B1(n9414), .B2(n9410), .A(n9409), .ZN(n9495) );
  MUX2_X1 U10472 ( .A(n9411), .B(n9495), .S(n9456), .Z(n9412) );
  OAI21_X1 U10473 ( .B1(n9498), .B2(n9432), .A(n9412), .ZN(P2_U3482) );
  INV_X1 U10474 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9416) );
  AOI21_X1 U10475 ( .B1(n9415), .B2(n9414), .A(n9413), .ZN(n9499) );
  MUX2_X1 U10476 ( .A(n9416), .B(n9499), .S(n9456), .Z(n9417) );
  OAI21_X1 U10477 ( .B1(n9502), .B2(n9432), .A(n9417), .ZN(P2_U3481) );
  NAND2_X1 U10478 ( .A1(n9418), .A2(n9463), .ZN(n9419) );
  OAI211_X1 U10479 ( .C1(n9458), .C2(n9421), .A(n9420), .B(n9419), .ZN(n9503)
         );
  MUX2_X1 U10480 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9503), .S(n9456), .Z(
        P2_U3480) );
  NAND2_X1 U10481 ( .A1(n9422), .A2(n9463), .ZN(n9423) );
  OAI211_X1 U10482 ( .C1(n9458), .C2(n9425), .A(n9424), .B(n9423), .ZN(n9504)
         );
  MUX2_X1 U10483 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9504), .S(n9456), .Z(
        P2_U3479) );
  NOR2_X1 U10484 ( .A1(n9426), .A2(n9458), .ZN(n9429) );
  AOI21_X1 U10485 ( .B1(n9429), .B2(n9428), .A(n9427), .ZN(n9505) );
  MUX2_X1 U10486 ( .A(n9430), .B(n9505), .S(n9456), .Z(n9431) );
  OAI21_X1 U10487 ( .B1(n9509), .B2(n9432), .A(n9431), .ZN(P2_U3478) );
  NAND2_X1 U10488 ( .A1(n9433), .A2(n9463), .ZN(n9434) );
  OAI211_X1 U10489 ( .C1(n9458), .C2(n9436), .A(n9435), .B(n9434), .ZN(n9510)
         );
  MUX2_X1 U10490 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9510), .S(n9456), .Z(
        P2_U3477) );
  NAND2_X1 U10491 ( .A1(n9437), .A2(n9463), .ZN(n9438) );
  OAI211_X1 U10492 ( .C1(n9458), .C2(n9440), .A(n9439), .B(n9438), .ZN(n9511)
         );
  MUX2_X1 U10493 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9511), .S(n9456), .Z(
        P2_U3476) );
  NAND2_X1 U10494 ( .A1(n9441), .A2(n9463), .ZN(n9442) );
  OAI211_X1 U10495 ( .C1(n9458), .C2(n9444), .A(n9443), .B(n9442), .ZN(n9512)
         );
  MUX2_X1 U10496 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9512), .S(n9456), .Z(
        P2_U3475) );
  NOR2_X1 U10497 ( .A1(n9445), .A2(n9458), .ZN(n9447) );
  AOI211_X1 U10498 ( .C1(n9463), .C2(n9448), .A(n9447), .B(n9446), .ZN(n11120)
         );
  NAND2_X1 U10499 ( .A1(n9465), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n9449) );
  OAI21_X1 U10500 ( .B1(n11120), .B2(n9465), .A(n9449), .ZN(P2_U3474) );
  OAI22_X1 U10501 ( .A1(n9452), .A2(n9458), .B1(n9451), .B2(n9450), .ZN(n9453)
         );
  NOR2_X1 U10502 ( .A1(n9454), .A2(n9453), .ZN(n11118) );
  OR2_X1 U10503 ( .A1(n9456), .A2(n9455), .ZN(n9457) );
  OAI21_X1 U10504 ( .B1(n11118), .B2(n9465), .A(n9457), .ZN(P2_U3473) );
  NOR2_X1 U10505 ( .A1(n9459), .A2(n9458), .ZN(n9461) );
  AOI211_X1 U10506 ( .C1(n9463), .C2(n9462), .A(n9461), .B(n9460), .ZN(n11116)
         );
  NAND2_X1 U10507 ( .A1(n9465), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n9464) );
  OAI21_X1 U10508 ( .B1(n11116), .B2(n9465), .A(n9464), .ZN(P2_U3472) );
  NAND2_X1 U10509 ( .A1(n9467), .A2(n9466), .ZN(n9473) );
  NOR2_X1 U10510 ( .A1(n6890), .A2(n9468), .ZN(n9471) );
  AOI21_X1 U10511 ( .B1(P2_REG0_REG_31__SCAN_IN), .B2(n6890), .A(n9471), .ZN(
        n9469) );
  OAI21_X1 U10512 ( .B1(n9470), .B2(n9473), .A(n9469), .ZN(P2_U3458) );
  AOI21_X1 U10513 ( .B1(P2_REG0_REG_30__SCAN_IN), .B2(n6890), .A(n9471), .ZN(
        n9472) );
  OAI21_X1 U10514 ( .B1(n9474), .B2(n9473), .A(n9472), .ZN(P2_U3457) );
  MUX2_X1 U10515 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9475), .S(n11121), .Z(
        n9476) );
  INV_X1 U10516 ( .A(n9476), .ZN(n9477) );
  OAI21_X1 U10517 ( .B1(n9478), .B2(n9508), .A(n9477), .ZN(P2_U3455) );
  MUX2_X1 U10518 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9479), .S(n11121), .Z(
        n9480) );
  INV_X1 U10519 ( .A(n9480), .ZN(n9481) );
  OAI21_X1 U10520 ( .B1(n9482), .B2(n9508), .A(n9481), .ZN(P2_U3454) );
  INV_X1 U10521 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9484) );
  MUX2_X1 U10522 ( .A(n9484), .B(n9483), .S(n11121), .Z(n9485) );
  OAI21_X1 U10523 ( .B1(n9486), .B2(n9508), .A(n9485), .ZN(P2_U3453) );
  INV_X1 U10524 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9488) );
  MUX2_X1 U10525 ( .A(n9488), .B(n9487), .S(n11121), .Z(n9489) );
  OAI21_X1 U10526 ( .B1(n9490), .B2(n9508), .A(n9489), .ZN(P2_U3452) );
  INV_X1 U10527 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9492) );
  MUX2_X1 U10528 ( .A(n9492), .B(n9491), .S(n11121), .Z(n9493) );
  OAI21_X1 U10529 ( .B1(n9494), .B2(n9508), .A(n9493), .ZN(P2_U3451) );
  INV_X1 U10530 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9496) );
  MUX2_X1 U10531 ( .A(n9496), .B(n9495), .S(n11121), .Z(n9497) );
  OAI21_X1 U10532 ( .B1(n9498), .B2(n9508), .A(n9497), .ZN(P2_U3450) );
  INV_X1 U10533 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9500) );
  MUX2_X1 U10534 ( .A(n9500), .B(n9499), .S(n11121), .Z(n9501) );
  OAI21_X1 U10535 ( .B1(n9502), .B2(n9508), .A(n9501), .ZN(P2_U3449) );
  MUX2_X1 U10536 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9503), .S(n11121), .Z(
        P2_U3448) );
  MUX2_X1 U10537 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9504), .S(n11121), .Z(
        P2_U3447) );
  INV_X1 U10538 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9506) );
  MUX2_X1 U10539 ( .A(n9506), .B(n9505), .S(n11121), .Z(n9507) );
  OAI21_X1 U10540 ( .B1(n9509), .B2(n9508), .A(n9507), .ZN(P2_U3446) );
  MUX2_X1 U10541 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9510), .S(n11121), .Z(
        P2_U3444) );
  MUX2_X1 U10542 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9511), .S(n11121), .Z(
        P2_U3441) );
  MUX2_X1 U10543 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9512), .S(n11121), .Z(
        P2_U3438) );
  OAI222_X1 U10544 ( .A1(n8667), .A2(n9516), .B1(n9515), .B2(P2_U3151), .C1(
        n9514), .C2(n9513), .ZN(P2_U3266) );
  INV_X1 U10545 ( .A(n9517), .ZN(n9518) );
  MUX2_X1 U10546 ( .A(n9518), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  XNOR2_X1 U10547 ( .A(n9520), .B(n9519), .ZN(n9521) );
  XNOR2_X1 U10548 ( .A(n9522), .B(n9521), .ZN(n9529) );
  AOI22_X1 U10549 ( .A1(n9689), .A2(n9524), .B1(n9687), .B2(n5697), .ZN(n9525)
         );
  NAND2_X1 U10550 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n10064)
         );
  OAI211_X1 U10551 ( .C1(n9571), .C2(n9691), .A(n9525), .B(n10064), .ZN(n9526)
         );
  AOI21_X1 U10552 ( .B1(n9527), .B2(n9694), .A(n9526), .ZN(n9528) );
  OAI21_X1 U10553 ( .B1(n9529), .B2(n9697), .A(n9528), .ZN(P1_U3215) );
  AOI21_X1 U10554 ( .B1(n9532), .B2(n9638), .A(n9531), .ZN(n9533) );
  OAI21_X1 U10555 ( .B1(n9612), .B2(n9533), .A(n9676), .ZN(n9537) );
  INV_X1 U10556 ( .A(n10217), .ZN(n10347) );
  AOI22_X1 U10557 ( .A1(n9687), .A2(n10347), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9536) );
  INV_X1 U10558 ( .A(n10248), .ZN(n10348) );
  AOI22_X1 U10559 ( .A1(n9689), .A2(n10214), .B1(n9678), .B2(n10348), .ZN(
        n9535) );
  NAND2_X1 U10560 ( .A1(n10222), .A2(n9694), .ZN(n9534) );
  NAND4_X1 U10561 ( .A1(n9537), .A2(n9536), .A3(n9535), .A4(n9534), .ZN(
        P1_U3216) );
  XNOR2_X1 U10562 ( .A(n9539), .B(n9538), .ZN(n9540) );
  XNOR2_X1 U10563 ( .A(n9541), .B(n9540), .ZN(n9549) );
  AOI22_X1 U10564 ( .A1(n9689), .A2(n9542), .B1(n9687), .B2(n9996), .ZN(n9544)
         );
  OAI211_X1 U10565 ( .C1(n9545), .C2(n9691), .A(n9544), .B(n9543), .ZN(n9546)
         );
  AOI21_X1 U10566 ( .B1(n9547), .B2(n9694), .A(n9546), .ZN(n9548) );
  OAI21_X1 U10567 ( .B1(n9549), .B2(n9697), .A(n9548), .ZN(P1_U3217) );
  OAI21_X1 U10568 ( .B1(n9552), .B2(n9551), .A(n9550), .ZN(n9553) );
  NAND2_X1 U10569 ( .A1(n9553), .A2(n9676), .ZN(n9557) );
  AND2_X1 U10570 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n10118) );
  INV_X1 U10571 ( .A(n10284), .ZN(n9554) );
  OAI22_X1 U10572 ( .A1(n9691), .A2(n6140), .B1(n9554), .B2(n9646), .ZN(n9555)
         );
  AOI211_X1 U10573 ( .C1(n9687), .C2(n9562), .A(n10118), .B(n9555), .ZN(n9556)
         );
  OAI211_X1 U10574 ( .C1(n5401), .C2(n9636), .A(n9557), .B(n9556), .ZN(
        P1_U3219) );
  AOI21_X1 U10575 ( .B1(n9619), .B2(n9559), .A(n9558), .ZN(n9560) );
  NOR3_X1 U10576 ( .A1(n9561), .A2(n9560), .A3(n9697), .ZN(n9566) );
  INV_X1 U10577 ( .A(n10253), .ZN(n10458) );
  AOI22_X1 U10578 ( .A1(n9678), .A2(n9562), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n9564) );
  AOI22_X1 U10579 ( .A1(n9689), .A2(n10254), .B1(n9687), .B2(n10348), .ZN(
        n9563) );
  OAI211_X1 U10580 ( .C1(n10458), .C2(n9636), .A(n9564), .B(n9563), .ZN(n9565)
         );
  OR2_X1 U10581 ( .A1(n9566), .A2(n9565), .ZN(P1_U3223) );
  INV_X1 U10582 ( .A(n9567), .ZN(n9570) );
  AOI21_X1 U10583 ( .B1(n9655), .B2(n9659), .A(n9568), .ZN(n9569) );
  OAI21_X1 U10584 ( .B1(n9570), .B2(n9569), .A(n9676), .ZN(n9576) );
  OAI22_X1 U10585 ( .A1(n9646), .A2(n9572), .B1(n9644), .B2(n9571), .ZN(n9573)
         );
  AOI211_X1 U10586 ( .C1(n9678), .C2(n9996), .A(n9574), .B(n9573), .ZN(n9575)
         );
  OAI211_X1 U10587 ( .C1(n11104), .C2(n9636), .A(n9576), .B(n9575), .ZN(
        P1_U3224) );
  OAI21_X1 U10588 ( .B1(n9579), .B2(n9578), .A(n9577), .ZN(n9583) );
  AOI22_X1 U10589 ( .A1(n9687), .A2(n10334), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9581) );
  AOI22_X1 U10590 ( .A1(n9689), .A2(n10186), .B1(n9678), .B2(n10347), .ZN(
        n9580) );
  OAI211_X1 U10591 ( .C1(n10441), .C2(n9636), .A(n9581), .B(n9580), .ZN(n9582)
         );
  AOI21_X1 U10592 ( .B1(n9583), .B2(n9676), .A(n9582), .ZN(n9584) );
  INV_X1 U10593 ( .A(n9584), .ZN(P1_U3225) );
  NAND2_X1 U10594 ( .A1(n9585), .A2(n9597), .ZN(n9590) );
  INV_X1 U10595 ( .A(n9686), .ZN(n9587) );
  INV_X1 U10596 ( .A(n9684), .ZN(n9586) );
  NOR2_X1 U10597 ( .A1(n9587), .A2(n9586), .ZN(n9588) );
  OAI22_X1 U10598 ( .A1(n9588), .A2(n9683), .B1(n9686), .B2(n9684), .ZN(n9589)
         );
  NOR2_X1 U10599 ( .A1(n9589), .A2(n9590), .ZN(n9600) );
  AOI21_X1 U10600 ( .B1(n9590), .B2(n9589), .A(n9600), .ZN(n9596) );
  AOI22_X1 U10601 ( .A1(n9591), .A2(n9689), .B1(n9678), .B2(n5697), .ZN(n9593)
         );
  OAI211_X1 U10602 ( .C1(n10297), .C2(n9644), .A(n9593), .B(n9592), .ZN(n9594)
         );
  AOI21_X1 U10603 ( .B1(n10398), .B2(n9694), .A(n9594), .ZN(n9595) );
  OAI21_X1 U10604 ( .B1(n9596), .B2(n9697), .A(n9595), .ZN(P1_U3226) );
  INV_X1 U10605 ( .A(n9597), .ZN(n9599) );
  NOR3_X1 U10606 ( .A1(n9600), .A2(n9599), .A3(n9598), .ZN(n9603) );
  INV_X1 U10607 ( .A(n9601), .ZN(n9602) );
  OAI21_X1 U10608 ( .B1(n9603), .B2(n9602), .A(n9676), .ZN(n9608) );
  INV_X1 U10609 ( .A(n10389), .ZN(n10405) );
  INV_X1 U10610 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9604) );
  NOR2_X1 U10611 ( .A1(n9604), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10081) );
  OAI22_X1 U10612 ( .A1(n9644), .A2(n6140), .B1(n9605), .B2(n9646), .ZN(n9606)
         );
  AOI211_X1 U10613 ( .C1(n9678), .C2(n10405), .A(n10081), .B(n9606), .ZN(n9607) );
  OAI211_X1 U10614 ( .C1(n10390), .C2(n9636), .A(n9608), .B(n9607), .ZN(
        P1_U3228) );
  INV_X1 U10615 ( .A(n9609), .ZN(n9614) );
  NOR3_X1 U10616 ( .A1(n9612), .A2(n9611), .A3(n9610), .ZN(n9613) );
  OAI21_X1 U10617 ( .B1(n9614), .B2(n9613), .A(n9676), .ZN(n9618) );
  AOI22_X1 U10618 ( .A1(n9687), .A2(n10325), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9617) );
  AOI22_X1 U10619 ( .A1(n10202), .A2(n9689), .B1(n9678), .B2(n10230), .ZN(
        n9616) );
  NAND2_X1 U10620 ( .A1(n10201), .A2(n9694), .ZN(n9615) );
  NAND4_X1 U10621 ( .A1(n9618), .A2(n9617), .A3(n9616), .A4(n9615), .ZN(
        P1_U3229) );
  OAI21_X1 U10622 ( .B1(n9621), .B2(n9620), .A(n9619), .ZN(n9625) );
  AOI22_X1 U10623 ( .A1(n9687), .A2(n10231), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9623) );
  AOI22_X1 U10624 ( .A1(n9689), .A2(n10264), .B1(n9678), .B2(n10265), .ZN(
        n9622) );
  OAI211_X1 U10625 ( .C1(n10368), .C2(n9636), .A(n9623), .B(n9622), .ZN(n9624)
         );
  AOI21_X1 U10626 ( .B1(n9625), .B2(n9676), .A(n9624), .ZN(n9626) );
  INV_X1 U10627 ( .A(n9626), .ZN(P1_U3233) );
  AND2_X1 U10628 ( .A1(n9567), .A2(n9627), .ZN(n9630) );
  OAI211_X1 U10629 ( .C1(n9630), .C2(n9629), .A(n9676), .B(n9628), .ZN(n9635)
         );
  NAND2_X1 U10630 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n10050)
         );
  INV_X1 U10631 ( .A(n10050), .ZN(n9633) );
  OAI22_X1 U10632 ( .A1(n9646), .A2(n9631), .B1(n9644), .B2(n9692), .ZN(n9632)
         );
  AOI211_X1 U10633 ( .C1(n9678), .C2(n11087), .A(n9633), .B(n9632), .ZN(n9634)
         );
  OAI211_X1 U10634 ( .C1(n9637), .C2(n9636), .A(n9635), .B(n9634), .ZN(
        P1_U3234) );
  NAND2_X1 U10635 ( .A1(n9639), .A2(n9638), .ZN(n9640) );
  XOR2_X1 U10636 ( .A(n9641), .B(n9640), .Z(n9650) );
  OAI22_X1 U10637 ( .A1(n9691), .A2(n10273), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9642), .ZN(n9648) );
  INV_X1 U10638 ( .A(n10238), .ZN(n9645) );
  OAI22_X1 U10639 ( .A1(n9646), .A2(n9645), .B1(n9644), .B2(n9643), .ZN(n9647)
         );
  AOI211_X1 U10640 ( .C1(n10237), .C2(n9694), .A(n9648), .B(n9647), .ZN(n9649)
         );
  OAI21_X1 U10641 ( .B1(n9650), .B2(n9697), .A(n9649), .ZN(P1_U3235) );
  AOI22_X1 U10642 ( .A1(n9689), .A2(n9651), .B1(n9687), .B2(n11087), .ZN(n9653) );
  OAI211_X1 U10643 ( .C1(n9654), .C2(n9691), .A(n9653), .B(n9652), .ZN(n9662)
         );
  INV_X1 U10644 ( .A(n9655), .ZN(n9660) );
  AOI21_X1 U10645 ( .B1(n9657), .B2(n9659), .A(n9656), .ZN(n9658) );
  AOI211_X1 U10646 ( .C1(n9660), .C2(n9659), .A(n9697), .B(n9658), .ZN(n9661)
         );
  AOI211_X1 U10647 ( .C1(n9663), .C2(n9694), .A(n9662), .B(n9661), .ZN(n9664)
         );
  INV_X1 U10648 ( .A(n9664), .ZN(P1_U3236) );
  NOR2_X1 U10649 ( .A1(n9665), .A2(n5163), .ZN(n9667) );
  XNOR2_X1 U10650 ( .A(n9667), .B(n9666), .ZN(n9671) );
  AOI22_X1 U10651 ( .A1(n9689), .A2(n10302), .B1(n9687), .B2(n10265), .ZN(
        n9668) );
  NAND2_X1 U10652 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10093)
         );
  OAI211_X1 U10653 ( .C1(n10297), .C2(n9691), .A(n9668), .B(n10093), .ZN(n9669) );
  AOI21_X1 U10654 ( .B1(n10385), .B2(n9694), .A(n9669), .ZN(n9670) );
  OAI21_X1 U10655 ( .B1(n9671), .B2(n9697), .A(n9670), .ZN(P1_U3238) );
  INV_X1 U10656 ( .A(n9577), .ZN(n9674) );
  NAND3_X1 U10657 ( .A1(n9677), .A2(n9676), .A3(n9675), .ZN(n9682) );
  AOI22_X1 U10658 ( .A1(n9678), .A2(n10325), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9681) );
  AOI22_X1 U10659 ( .A1(n9689), .A2(n10171), .B1(n9687), .B2(n10326), .ZN(
        n9680) );
  NAND2_X1 U10660 ( .A1(n10178), .A2(n9694), .ZN(n9679) );
  NAND4_X1 U10661 ( .A1(n9682), .A2(n9681), .A3(n9680), .A4(n9679), .ZN(
        P1_U3240) );
  XNOR2_X1 U10662 ( .A(n9684), .B(n9683), .ZN(n9685) );
  XNOR2_X1 U10663 ( .A(n9686), .B(n9685), .ZN(n9698) );
  AOI22_X1 U10664 ( .A1(n9689), .A2(n9688), .B1(n9687), .B2(n10405), .ZN(n9690) );
  NAND2_X1 U10665 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10867)
         );
  OAI211_X1 U10666 ( .C1(n9692), .C2(n9691), .A(n9690), .B(n10867), .ZN(n9693)
         );
  AOI21_X1 U10667 ( .B1(n9695), .B2(n9694), .A(n9693), .ZN(n9696) );
  OAI21_X1 U10668 ( .B1(n9698), .B2(n9697), .A(n9696), .ZN(P1_U3241) );
  NOR3_X1 U10669 ( .A1(n9701), .A2(n9700), .A3(n9699), .ZN(n9993) );
  OAI21_X1 U10670 ( .B1(n9756), .B2(n6327), .A(P1_B_REG_SCAN_IN), .ZN(n9992)
         );
  NAND2_X1 U10671 ( .A1(n10477), .A2(n9708), .ZN(n9703) );
  INV_X1 U10672 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10472) );
  OR2_X1 U10673 ( .A1(n9709), .A2(n10472), .ZN(n9702) );
  NAND2_X1 U10674 ( .A1(n5131), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n9707) );
  NAND2_X1 U10675 ( .A1(n9704), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n9706) );
  NAND2_X1 U10676 ( .A1(n6066), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n9705) );
  NAND3_X1 U10677 ( .A1(n9707), .A2(n9706), .A3(n9705), .ZN(n10129) );
  NOR2_X1 U10678 ( .A1(n10426), .A2(n10129), .ZN(n9816) );
  NAND2_X1 U10679 ( .A1(n8839), .A2(n9708), .ZN(n9711) );
  OR2_X1 U10680 ( .A1(n9709), .A2(n10760), .ZN(n9710) );
  INV_X1 U10681 ( .A(n9994), .ZN(n9752) );
  NOR2_X1 U10682 ( .A1(n10135), .A2(n9752), .ZN(n9812) );
  NOR2_X1 U10683 ( .A1(n9816), .A2(n9812), .ZN(n9804) );
  AND2_X1 U10684 ( .A1(n9968), .A2(n9963), .ZN(n9715) );
  NAND2_X1 U10685 ( .A1(n9962), .A2(n9961), .ZN(n9713) );
  INV_X1 U10686 ( .A(n9969), .ZN(n9712) );
  AOI21_X1 U10687 ( .B1(n9715), .B2(n9713), .A(n9712), .ZN(n9714) );
  NAND2_X1 U10688 ( .A1(n9974), .A2(n9714), .ZN(n9769) );
  INV_X1 U10689 ( .A(n9715), .ZN(n9716) );
  NAND2_X1 U10690 ( .A1(n9959), .A2(n9950), .ZN(n9957) );
  OR2_X1 U10691 ( .A1(n9716), .A2(n9957), .ZN(n9766) );
  NAND2_X1 U10692 ( .A1(n9942), .A2(n10208), .ZN(n9825) );
  NAND2_X1 U10693 ( .A1(n9825), .A2(n9943), .ZN(n9717) );
  NAND2_X1 U10694 ( .A1(n9947), .A2(n9717), .ZN(n9718) );
  NAND2_X1 U10695 ( .A1(n9718), .A2(n9949), .ZN(n9719) );
  NAND2_X1 U10696 ( .A1(n9952), .A2(n9719), .ZN(n9762) );
  NAND2_X1 U10697 ( .A1(n9943), .A2(n9720), .ZN(n9824) );
  INV_X1 U10698 ( .A(n9721), .ZN(n9722) );
  NOR2_X1 U10699 ( .A1(n9824), .A2(n9722), .ZN(n9723) );
  NAND2_X1 U10700 ( .A1(n9723), .A2(n9949), .ZN(n9761) );
  INV_X1 U10701 ( .A(n9928), .ZN(n9933) );
  AND2_X1 U10702 ( .A1(n9921), .A2(n9724), .ZN(n9923) );
  AND2_X1 U10703 ( .A1(n9910), .A2(n9905), .ZN(n9894) );
  NAND2_X1 U10704 ( .A1(n6332), .A2(n11034), .ZN(n9727) );
  NAND2_X1 U10705 ( .A1(n10005), .A2(n9725), .ZN(n9726) );
  AND3_X1 U10706 ( .A1(n9727), .A2(n9726), .A3(n6328), .ZN(n9728) );
  OAI211_X1 U10707 ( .C1(n9729), .C2(n9728), .A(n9836), .B(n9831), .ZN(n9730)
         );
  INV_X1 U10708 ( .A(n9837), .ZN(n9828) );
  AOI21_X1 U10709 ( .B1(n9730), .B2(n9834), .A(n9828), .ZN(n9733) );
  NAND2_X1 U10710 ( .A1(n9827), .A2(n9731), .ZN(n9732) );
  OAI21_X1 U10711 ( .B1(n9733), .B2(n9732), .A(n9842), .ZN(n9734) );
  NAND2_X1 U10712 ( .A1(n9734), .A2(n9849), .ZN(n9735) );
  NAND3_X1 U10713 ( .A1(n9735), .A2(n9779), .A3(n9850), .ZN(n9737) );
  NAND2_X1 U10714 ( .A1(n9737), .A2(n9736), .ZN(n9738) );
  NAND2_X1 U10715 ( .A1(n9738), .A2(n9874), .ZN(n9739) );
  AND2_X1 U10716 ( .A1(n9881), .A2(n9869), .ZN(n9871) );
  NAND2_X1 U10717 ( .A1(n9891), .A2(n9879), .ZN(n9884) );
  AOI21_X1 U10718 ( .B1(n9739), .B2(n9871), .A(n9884), .ZN(n9740) );
  NAND2_X1 U10719 ( .A1(n9892), .A2(n9882), .ZN(n9898) );
  OAI211_X1 U10720 ( .C1(n9740), .C2(n9898), .A(n9903), .B(n9901), .ZN(n9742)
         );
  INV_X1 U10721 ( .A(n9909), .ZN(n9741) );
  AOI21_X1 U10722 ( .B1(n9894), .B2(n9742), .A(n9741), .ZN(n9744) );
  INV_X1 U10723 ( .A(n9913), .ZN(n9743) );
  OAI211_X1 U10724 ( .C1(n9744), .C2(n9743), .A(n9920), .B(n9914), .ZN(n9745)
         );
  AOI21_X1 U10725 ( .B1(n9923), .B2(n9745), .A(n9919), .ZN(n9747) );
  OAI21_X1 U10726 ( .B1(n9933), .B2(n9747), .A(n9746), .ZN(n9748) );
  INV_X1 U10727 ( .A(n9748), .ZN(n9749) );
  NOR2_X1 U10728 ( .A1(n9761), .A2(n9749), .ZN(n9750) );
  NOR2_X1 U10729 ( .A1(n9762), .A2(n9750), .ZN(n9751) );
  NOR2_X1 U10730 ( .A1(n9766), .A2(n9751), .ZN(n9753) );
  NAND2_X1 U10731 ( .A1(n10135), .A2(n9752), .ZN(n9802) );
  OAI211_X1 U10732 ( .C1(n9769), .C2(n9753), .A(n9975), .B(n9802), .ZN(n9754)
         );
  AND2_X1 U10733 ( .A1(n10426), .A2(n10129), .ZN(n9818) );
  AOI21_X1 U10734 ( .B1(n9804), .B2(n9754), .A(n9818), .ZN(n9757) );
  NOR3_X1 U10735 ( .A1(n9757), .A2(n9986), .A3(n5130), .ZN(n9755) );
  AOI211_X1 U10736 ( .C1(n9758), .C2(n9757), .A(n9756), .B(n9755), .ZN(n9990)
         );
  INV_X1 U10737 ( .A(n9812), .ZN(n9759) );
  NAND2_X1 U10738 ( .A1(n9759), .A2(n10129), .ZN(n9760) );
  AOI21_X1 U10739 ( .B1(n9760), .B2(n10127), .A(n9808), .ZN(n9807) );
  INV_X1 U10740 ( .A(n9761), .ZN(n9764) );
  AOI21_X1 U10741 ( .B1(n9764), .B2(n9763), .A(n9762), .ZN(n9765) );
  NOR2_X1 U10742 ( .A1(n9766), .A2(n9765), .ZN(n9768) );
  NAND2_X1 U10743 ( .A1(n10129), .A2(n9994), .ZN(n9767) );
  NAND2_X1 U10744 ( .A1(n10135), .A2(n9767), .ZN(n9977) );
  OAI211_X1 U10745 ( .C1(n9769), .C2(n9768), .A(n9975), .B(n9977), .ZN(n9806)
         );
  INV_X1 U10746 ( .A(n10184), .ZN(n9948) );
  INV_X1 U10747 ( .A(n10249), .ZN(n9936) );
  NAND2_X1 U10748 ( .A1(n5173), .A2(n9770), .ZN(n10279) );
  INV_X1 U10749 ( .A(n9771), .ZN(n9790) );
  INV_X1 U10750 ( .A(n9772), .ZN(n9778) );
  NOR2_X1 U10751 ( .A1(n7689), .A2(n6328), .ZN(n9774) );
  NAND4_X1 U10752 ( .A1(n9774), .A2(n9773), .A3(n11021), .A4(n5416), .ZN(n9776) );
  NOR4_X1 U10753 ( .A1(n9776), .A2(n9843), .A3(n9775), .A4(n9847), .ZN(n9777)
         );
  NAND4_X1 U10754 ( .A1(n9779), .A2(n9778), .A3(n9777), .A4(n9872), .ZN(n9780)
         );
  NOR2_X1 U10755 ( .A1(n9781), .A2(n9780), .ZN(n9782) );
  NAND4_X1 U10756 ( .A1(n9785), .A2(n9784), .A3(n9783), .A4(n9782), .ZN(n9786)
         );
  NOR2_X1 U10757 ( .A1(n9787), .A2(n9786), .ZN(n9788) );
  NAND3_X1 U10758 ( .A1(n9790), .A2(n9789), .A3(n9788), .ZN(n9791) );
  NOR2_X1 U10759 ( .A1(n9792), .A2(n9791), .ZN(n9793) );
  XNOR2_X1 U10760 ( .A(n10385), .B(n10282), .ZN(n10294) );
  NAND3_X1 U10761 ( .A1(n10279), .A2(n9793), .A3(n10294), .ZN(n9794) );
  NOR2_X1 U10762 ( .A1(n10270), .A2(n9794), .ZN(n9795) );
  NAND2_X1 U10763 ( .A1(n9936), .A2(n9795), .ZN(n9796) );
  NOR3_X1 U10764 ( .A1(n10212), .A2(n10234), .A3(n9796), .ZN(n9797) );
  NAND4_X1 U10765 ( .A1(n10169), .A2(n10198), .A3(n9948), .A4(n9797), .ZN(
        n9798) );
  NOR4_X1 U10766 ( .A1(n9800), .A2(n9799), .A3(n6287), .A4(n9798), .ZN(n9803)
         );
  INV_X1 U10767 ( .A(n9818), .ZN(n9801) );
  NAND4_X1 U10768 ( .A1(n9804), .A2(n9803), .A3(n9802), .A4(n9801), .ZN(n9982)
         );
  INV_X1 U10769 ( .A(n9982), .ZN(n9805) );
  AOI21_X1 U10770 ( .B1(n9807), .B2(n9806), .A(n9805), .ZN(n9988) );
  NOR2_X1 U10771 ( .A1(n6324), .A2(n5130), .ZN(n9815) );
  OR3_X1 U10772 ( .A1(n10127), .A2(n9808), .A3(n9977), .ZN(n9811) );
  INV_X1 U10773 ( .A(n10129), .ZN(n9809) );
  OR3_X1 U10774 ( .A1(n9977), .A2(n9809), .A3(n9808), .ZN(n9810) );
  OAI211_X1 U10775 ( .C1(n6328), .C2(n9987), .A(n9811), .B(n9810), .ZN(n9814)
         );
  NAND2_X1 U10776 ( .A1(n9812), .A2(n10129), .ZN(n9821) );
  AOI211_X1 U10777 ( .C1(n10129), .C2(n9821), .A(n9987), .B(n10426), .ZN(n9813) );
  AOI211_X1 U10778 ( .C1(n9818), .C2(n9815), .A(n9814), .B(n9813), .ZN(n9984)
         );
  INV_X1 U10779 ( .A(n9816), .ZN(n9822) );
  NAND3_X1 U10780 ( .A1(n9821), .A2(n9817), .A3(n9822), .ZN(n9981) );
  INV_X1 U10781 ( .A(n9977), .ZN(n9820) );
  AOI21_X1 U10782 ( .B1(n6918), .B2(n6328), .A(n5130), .ZN(n9819) );
  AOI211_X1 U10783 ( .C1(n9820), .C2(n5130), .A(n9819), .B(n9818), .ZN(n9823)
         );
  NAND3_X1 U10784 ( .A1(n9823), .A2(n9822), .A3(n9821), .ZN(n9980) );
  MUX2_X1 U10785 ( .A(n9825), .B(n9824), .S(n9973), .Z(n9946) );
  NAND2_X1 U10786 ( .A1(n9826), .A2(n9836), .ZN(n9830) );
  AND2_X1 U10787 ( .A1(n9827), .A2(n9834), .ZN(n9829) );
  AOI21_X1 U10788 ( .B1(n9830), .B2(n9829), .A(n9828), .ZN(n9840) );
  NAND2_X1 U10789 ( .A1(n9832), .A2(n9831), .ZN(n9835) );
  NAND3_X1 U10790 ( .A1(n9835), .A2(n9834), .A3(n9833), .ZN(n9838) );
  NAND3_X1 U10791 ( .A1(n9838), .A2(n9837), .A3(n9836), .ZN(n9839) );
  MUX2_X1 U10792 ( .A(n9840), .B(n9839), .S(n9973), .Z(n9848) );
  INV_X1 U10793 ( .A(n9841), .ZN(n9845) );
  XNOR2_X1 U10794 ( .A(n9842), .B(n9973), .ZN(n9844) );
  AOI21_X1 U10795 ( .B1(n9845), .B2(n9844), .A(n9843), .ZN(n9846) );
  OAI21_X1 U10796 ( .B1(n9848), .B2(n9847), .A(n9846), .ZN(n9855) );
  INV_X1 U10797 ( .A(n9973), .ZN(n9958) );
  MUX2_X1 U10798 ( .A(n9850), .B(n9849), .S(n9958), .Z(n9851) );
  INV_X1 U10799 ( .A(n9851), .ZN(n9853) );
  NOR2_X1 U10800 ( .A1(n9853), .A2(n9852), .ZN(n9854) );
  NAND2_X1 U10801 ( .A1(n9855), .A2(n9854), .ZN(n9863) );
  INV_X1 U10802 ( .A(n9856), .ZN(n9857) );
  NOR2_X1 U10803 ( .A1(n9858), .A2(n9857), .ZN(n9861) );
  NAND3_X1 U10804 ( .A1(n9869), .A2(n9872), .A3(n9859), .ZN(n9860) );
  AOI21_X1 U10805 ( .B1(n9863), .B2(n9861), .A(n9860), .ZN(n9865) );
  NAND2_X1 U10806 ( .A1(n9863), .A2(n9862), .ZN(n9864) );
  MUX2_X1 U10807 ( .A(n9865), .B(n9864), .S(n9973), .Z(n9866) );
  NAND3_X1 U10808 ( .A1(n9866), .A2(n9874), .A3(n9867), .ZN(n9880) );
  INV_X1 U10809 ( .A(n9867), .ZN(n9868) );
  NAND2_X1 U10810 ( .A1(n9869), .A2(n9868), .ZN(n9870) );
  AND2_X1 U10811 ( .A1(n9870), .A2(n9874), .ZN(n9878) );
  INV_X1 U10812 ( .A(n9871), .ZN(n9876) );
  INV_X1 U10813 ( .A(n9872), .ZN(n9873) );
  AND2_X1 U10814 ( .A1(n9874), .A2(n9873), .ZN(n9875) );
  NOR2_X1 U10815 ( .A1(n9876), .A2(n9875), .ZN(n9877) );
  MUX2_X1 U10816 ( .A(n9878), .B(n9877), .S(n9973), .Z(n9886) );
  NAND3_X1 U10817 ( .A1(n9880), .A2(n9886), .A3(n9879), .ZN(n9890) );
  AND2_X1 U10818 ( .A1(n9882), .A2(n9881), .ZN(n9888) );
  INV_X1 U10819 ( .A(n9883), .ZN(n9885) );
  AOI21_X1 U10820 ( .B1(n9886), .B2(n9885), .A(n9884), .ZN(n9887) );
  MUX2_X1 U10821 ( .A(n9888), .B(n9887), .S(n9973), .Z(n9889) );
  NAND2_X1 U10822 ( .A1(n9890), .A2(n9889), .ZN(n9900) );
  NAND3_X1 U10823 ( .A1(n9900), .A2(n9901), .A3(n9891), .ZN(n9893) );
  NAND2_X1 U10824 ( .A1(n9893), .A2(n9892), .ZN(n9897) );
  INV_X1 U10825 ( .A(n9894), .ZN(n9895) );
  AOI21_X1 U10826 ( .B1(n9897), .B2(n9896), .A(n9895), .ZN(n9908) );
  INV_X1 U10827 ( .A(n9898), .ZN(n9899) );
  NAND2_X1 U10828 ( .A1(n9900), .A2(n9899), .ZN(n9902) );
  NAND2_X1 U10829 ( .A1(n9902), .A2(n9901), .ZN(n9906) );
  NAND2_X1 U10830 ( .A1(n9909), .A2(n9903), .ZN(n9904) );
  AOI21_X1 U10831 ( .B1(n9906), .B2(n9905), .A(n9904), .ZN(n9907) );
  MUX2_X1 U10832 ( .A(n9908), .B(n9907), .S(n9973), .Z(n9918) );
  NAND2_X1 U10833 ( .A1(n9914), .A2(n9909), .ZN(n9912) );
  NAND2_X1 U10834 ( .A1(n9913), .A2(n9910), .ZN(n9911) );
  MUX2_X1 U10835 ( .A(n9912), .B(n9911), .S(n9973), .Z(n9917) );
  MUX2_X1 U10836 ( .A(n9914), .B(n9913), .S(n9958), .Z(n9915) );
  OAI211_X1 U10837 ( .C1(n9918), .C2(n9917), .A(n9916), .B(n9915), .ZN(n9924)
         );
  NAND3_X1 U10838 ( .A1(n9924), .A2(n9920), .A3(n5410), .ZN(n9922) );
  NAND2_X1 U10839 ( .A1(n9922), .A2(n9921), .ZN(n9927) );
  NAND2_X1 U10840 ( .A1(n9924), .A2(n9923), .ZN(n9925) );
  NAND3_X1 U10841 ( .A1(n9925), .A2(n5410), .A3(n10269), .ZN(n9926) );
  MUX2_X1 U10842 ( .A(n9927), .B(n9926), .S(n9973), .Z(n9932) );
  AND2_X1 U10843 ( .A1(n9934), .A2(n9928), .ZN(n9929) );
  MUX2_X1 U10844 ( .A(n9930), .B(n9929), .S(n9973), .Z(n9931) );
  OAI21_X1 U10845 ( .B1(n9933), .B2(n9932), .A(n9931), .ZN(n9937) );
  MUX2_X1 U10846 ( .A(n9934), .B(n10244), .S(n9973), .Z(n9935) );
  NAND3_X1 U10847 ( .A1(n9937), .A2(n9936), .A3(n9935), .ZN(n9941) );
  MUX2_X1 U10848 ( .A(n9939), .B(n9938), .S(n9973), .Z(n9940) );
  AOI21_X1 U10849 ( .B1(n9941), .B2(n9940), .A(n10234), .ZN(n9945) );
  MUX2_X1 U10850 ( .A(n9943), .B(n9942), .S(n9973), .Z(n9944) );
  OAI211_X1 U10851 ( .C1(n9946), .C2(n9945), .A(n10198), .B(n9944), .ZN(n9951)
         );
  NAND3_X1 U10852 ( .A1(n9948), .A2(n9947), .A3(n9951), .ZN(n9955) );
  NAND3_X1 U10853 ( .A1(n9951), .A2(n9950), .A3(n9949), .ZN(n9953) );
  AND2_X1 U10854 ( .A1(n9953), .A2(n9952), .ZN(n9954) );
  MUX2_X1 U10855 ( .A(n9955), .B(n9954), .S(n9973), .Z(n9956) );
  NAND2_X1 U10856 ( .A1(n9956), .A2(n9961), .ZN(n9960) );
  AOI22_X1 U10857 ( .A1(n9960), .A2(n9959), .B1(n9958), .B2(n9957), .ZN(n9967)
         );
  OAI21_X1 U10858 ( .B1(n9973), .B2(n9961), .A(n10153), .ZN(n9966) );
  MUX2_X1 U10859 ( .A(n9963), .B(n9962), .S(n9973), .Z(n9964) );
  OAI211_X1 U10860 ( .C1(n9967), .C2(n9966), .A(n9965), .B(n9964), .ZN(n9971)
         );
  MUX2_X1 U10861 ( .A(n9969), .B(n9968), .S(n9973), .Z(n9970) );
  NAND3_X1 U10862 ( .A1(n9972), .A2(n9971), .A3(n9970), .ZN(n9978) );
  MUX2_X1 U10863 ( .A(n9975), .B(n9974), .S(n9973), .Z(n9976) );
  NAND3_X1 U10864 ( .A1(n9978), .A2(n9977), .A3(n9976), .ZN(n9979) );
  MUX2_X1 U10865 ( .A(n9981), .B(n9980), .S(n9979), .Z(n9983) );
  NAND3_X1 U10866 ( .A1(n9984), .A2(n9983), .A3(n9982), .ZN(n9985) );
  OAI211_X1 U10867 ( .C1(n9988), .C2(n9987), .A(n9986), .B(n9985), .ZN(n9989)
         );
  NAND2_X1 U10868 ( .A1(n9990), .A2(n9989), .ZN(n9991) );
  OAI21_X1 U10869 ( .B1(n9993), .B2(n9992), .A(n9991), .ZN(P1_U3242) );
  MUX2_X1 U10870 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n10129), .S(P1_U3973), .Z(
        P1_U3585) );
  MUX2_X1 U10871 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9994), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10872 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9995), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10873 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n10326), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10874 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n10334), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10875 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n10325), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10876 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n10347), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10877 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n10230), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10878 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n10348), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10879 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n10231), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10880 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n10265), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10881 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n10282), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10882 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n10405), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10883 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n5697), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10884 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n10406), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10885 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n10415), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10886 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n11087), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10887 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9996), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10888 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n11090), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10889 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9997), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10890 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9998), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10891 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9999), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10892 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n10000), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10893 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n10001), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10894 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n10002), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10895 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n10003), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10896 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n10004), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10897 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6332), .S(P1_U3973), .Z(
        P1_U3555) );
  MUX2_X1 U10898 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n10005), .S(P1_U3973), .Z(
        P1_U3554) );
  INV_X1 U10899 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n10010) );
  INV_X1 U10900 ( .A(n10006), .ZN(n10007) );
  NAND2_X1 U10901 ( .A1(n10866), .A2(n10007), .ZN(n10009) );
  OAI211_X1 U10902 ( .C1(n10010), .C2(n10869), .A(n10009), .B(n10008), .ZN(
        n10011) );
  INV_X1 U10903 ( .A(n10011), .ZN(n10020) );
  OAI211_X1 U10904 ( .C1(n10014), .C2(n10013), .A(n10871), .B(n10012), .ZN(
        n10019) );
  OAI211_X1 U10905 ( .C1(n10017), .C2(n10016), .A(n10877), .B(n10015), .ZN(
        n10018) );
  NAND3_X1 U10906 ( .A1(n10020), .A2(n10019), .A3(n10018), .ZN(P1_U3246) );
  INV_X1 U10907 ( .A(n10021), .ZN(n10034) );
  NOR2_X1 U10908 ( .A1(n10121), .A2(n10022), .ZN(n10023) );
  AOI211_X1 U10909 ( .C1(n10119), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n10024), .B(
        n10023), .ZN(n10033) );
  OAI211_X1 U10910 ( .C1(n10027), .C2(n10026), .A(n10877), .B(n10025), .ZN(
        n10032) );
  OAI211_X1 U10911 ( .C1(n10030), .C2(n10029), .A(n10871), .B(n10028), .ZN(
        n10031) );
  NAND4_X1 U10912 ( .A1(n10034), .A2(n10033), .A3(n10032), .A4(n10031), .ZN(
        P1_U3247) );
  OAI21_X1 U10913 ( .B1(n10037), .B2(n10036), .A(n10035), .ZN(n10038) );
  NAND2_X1 U10914 ( .A1(n10038), .A2(n10877), .ZN(n10048) );
  AOI21_X1 U10915 ( .B1(n10119), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n10039), .ZN(
        n10047) );
  OAI21_X1 U10916 ( .B1(n10042), .B2(n10041), .A(n10040), .ZN(n10043) );
  NAND2_X1 U10917 ( .A1(n10871), .A2(n10043), .ZN(n10046) );
  NAND2_X1 U10918 ( .A1(n10866), .A2(n10044), .ZN(n10045) );
  NAND4_X1 U10919 ( .A1(n10048), .A2(n10047), .A3(n10046), .A4(n10045), .ZN(
        P1_U3252) );
  INV_X1 U10920 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10052) );
  NAND2_X1 U10921 ( .A1(n10866), .A2(n10049), .ZN(n10051) );
  OAI211_X1 U10922 ( .C1(n10052), .C2(n10869), .A(n10051), .B(n10050), .ZN(
        n10053) );
  INV_X1 U10923 ( .A(n10053), .ZN(n10062) );
  OAI211_X1 U10924 ( .C1(n10056), .C2(n10055), .A(n10871), .B(n10054), .ZN(
        n10061) );
  OAI211_X1 U10925 ( .C1(n10059), .C2(n10058), .A(n10877), .B(n10057), .ZN(
        n10060) );
  NAND3_X1 U10926 ( .A1(n10062), .A2(n10061), .A3(n10060), .ZN(P1_U3256) );
  INV_X1 U10927 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10066) );
  NAND2_X1 U10928 ( .A1(n10866), .A2(n10063), .ZN(n10065) );
  OAI211_X1 U10929 ( .C1(n10066), .C2(n10869), .A(n10065), .B(n10064), .ZN(
        n10067) );
  INV_X1 U10930 ( .A(n10067), .ZN(n10076) );
  OAI211_X1 U10931 ( .C1(n10070), .C2(n10069), .A(n10871), .B(n10068), .ZN(
        n10075) );
  OAI211_X1 U10932 ( .C1(n10073), .C2(n10072), .A(n10877), .B(n10071), .ZN(
        n10074) );
  NAND3_X1 U10933 ( .A1(n10076), .A2(n10075), .A3(n10074), .ZN(P1_U3257) );
  XOR2_X1 U10934 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10078), .Z(n10088) );
  OAI21_X1 U10935 ( .B1(n10080), .B2(P1_REG1_REG_16__SCAN_IN), .A(n10077), 
        .ZN(n10089) );
  XOR2_X1 U10936 ( .A(n10088), .B(n10089), .Z(n10086) );
  XOR2_X1 U10937 ( .A(P1_REG2_REG_17__SCAN_IN), .B(n10078), .Z(n10102) );
  AOI21_X1 U10938 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n10080), .A(n10079), 
        .ZN(n10101) );
  XNOR2_X1 U10939 ( .A(n10102), .B(n10101), .ZN(n10084) );
  AOI21_X1 U10940 ( .B1(n10119), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n10081), 
        .ZN(n10082) );
  OAI21_X1 U10941 ( .B1(n10099), .B2(n10121), .A(n10082), .ZN(n10083) );
  AOI21_X1 U10942 ( .B1(n10871), .B2(n10084), .A(n10083), .ZN(n10085) );
  OAI21_X1 U10943 ( .B1(n10086), .B2(n10125), .A(n10085), .ZN(P1_U3260) );
  INV_X1 U10944 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n10087) );
  AOI22_X1 U10945 ( .A1(n10089), .A2(n10088), .B1(n10087), .B2(n10099), .ZN(
        n10092) );
  NAND2_X1 U10946 ( .A1(n10096), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n10108) );
  OAI21_X1 U10947 ( .B1(n10096), .B2(P1_REG1_REG_18__SCAN_IN), .A(n10108), 
        .ZN(n10090) );
  INV_X1 U10948 ( .A(n10090), .ZN(n10091) );
  NAND2_X1 U10949 ( .A1(n10092), .A2(n10091), .ZN(n10109) );
  OAI211_X1 U10950 ( .C1(n10092), .C2(n10091), .A(n10109), .B(n10877), .ZN(
        n10107) );
  OAI21_X1 U10951 ( .B1(n10869), .B2(n10094), .A(n10093), .ZN(n10095) );
  AOI21_X1 U10952 ( .B1(n10096), .B2(n10866), .A(n10095), .ZN(n10106) );
  INV_X1 U10953 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n10097) );
  AND2_X1 U10954 ( .A1(n10096), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n10112) );
  AOI21_X1 U10955 ( .B1(n10098), .B2(n10097), .A(n10112), .ZN(n10104) );
  INV_X1 U10956 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n10100) );
  AOI22_X1 U10957 ( .A1(n10102), .A2(n10101), .B1(n10100), .B2(n10099), .ZN(
        n10103) );
  NAND2_X1 U10958 ( .A1(n10103), .A2(n10104), .ZN(n10114) );
  OAI211_X1 U10959 ( .C1(n10104), .C2(n10103), .A(n10871), .B(n10114), .ZN(
        n10105) );
  NAND3_X1 U10960 ( .A1(n10107), .A2(n10106), .A3(n10105), .ZN(P1_U3261) );
  NAND2_X1 U10961 ( .A1(n10109), .A2(n10108), .ZN(n10111) );
  XNOR2_X1 U10962 ( .A(n5130), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n10110) );
  XNOR2_X1 U10963 ( .A(n10111), .B(n10110), .ZN(n10126) );
  INV_X1 U10964 ( .A(n10112), .ZN(n10113) );
  NAND2_X1 U10965 ( .A1(n10114), .A2(n10113), .ZN(n10117) );
  INV_X1 U10966 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n10115) );
  MUX2_X1 U10967 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n10115), .S(n5130), .Z(
        n10116) );
  XNOR2_X1 U10968 ( .A(n10117), .B(n10116), .ZN(n10123) );
  AOI21_X1 U10969 ( .B1(n10119), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n10118), 
        .ZN(n10120) );
  OAI21_X1 U10970 ( .B1(n5130), .B2(n10121), .A(n10120), .ZN(n10122) );
  AOI21_X1 U10971 ( .B1(n10871), .B2(n10123), .A(n10122), .ZN(n10124) );
  OAI21_X1 U10972 ( .B1(n10126), .B2(n10125), .A(n10124), .ZN(P1_U3262) );
  NAND2_X1 U10973 ( .A1(n10310), .A2(n10128), .ZN(n10133) );
  AND2_X1 U10974 ( .A1(n10130), .A2(n10129), .ZN(n10312) );
  INV_X1 U10975 ( .A(n10312), .ZN(n10131) );
  NOR2_X1 U10976 ( .A1(n11079), .A2(n10131), .ZN(n10137) );
  AOI21_X1 U10977 ( .B1(n11069), .B2(P1_REG2_REG_31__SCAN_IN), .A(n10137), 
        .ZN(n10132) );
  OAI211_X1 U10978 ( .C1(n10426), .C2(n11072), .A(n10133), .B(n10132), .ZN(
        P1_U3263) );
  XNOR2_X1 U10979 ( .A(n10135), .B(n10134), .ZN(n10136) );
  NOR2_X1 U10980 ( .A1(n10136), .A2(n10300), .ZN(n10313) );
  NAND2_X1 U10981 ( .A1(n10313), .A2(n11065), .ZN(n10139) );
  AOI21_X1 U10982 ( .B1(n11079), .B2(P1_REG2_REG_30__SCAN_IN), .A(n10137), 
        .ZN(n10138) );
  OAI211_X1 U10983 ( .C1(n10430), .C2(n11072), .A(n10139), .B(n10138), .ZN(
        P1_U3264) );
  NAND2_X1 U10984 ( .A1(n10140), .A2(n11075), .ZN(n10149) );
  AOI22_X1 U10985 ( .A1(n11069), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n10141), 
        .B2(n11067), .ZN(n10142) );
  OAI21_X1 U10986 ( .B1(n10143), .B2(n10316), .A(n10142), .ZN(n10146) );
  NOR2_X1 U10987 ( .A1(n10144), .A2(n10219), .ZN(n10145) );
  AOI211_X1 U10988 ( .C1(n10223), .C2(n10147), .A(n10146), .B(n10145), .ZN(
        n10148) );
  OAI211_X1 U10989 ( .C1(n10150), .C2(n11079), .A(n10149), .B(n10148), .ZN(
        P1_U3356) );
  XOR2_X1 U10990 ( .A(n10153), .B(n10151), .Z(n10322) );
  OAI21_X1 U10991 ( .B1(n10154), .B2(n10153), .A(n10152), .ZN(n10320) );
  INV_X1 U10992 ( .A(n10155), .ZN(n10156) );
  AOI211_X1 U10993 ( .C1(n10157), .C2(n5150), .A(n10300), .B(n10156), .ZN(
        n10318) );
  NAND2_X1 U10994 ( .A1(n10318), .A2(n11065), .ZN(n10162) );
  AOI22_X1 U10995 ( .A1(n11069), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n10158), 
        .B2(n11067), .ZN(n10159) );
  OAI21_X1 U10996 ( .B1(n10287), .B2(n10316), .A(n10159), .ZN(n10160) );
  AOI21_X1 U10997 ( .B1(n10283), .B2(n10334), .A(n10160), .ZN(n10161) );
  OAI211_X1 U10998 ( .C1(n10434), .C2(n11072), .A(n10162), .B(n10161), .ZN(
        n10163) );
  AOI21_X1 U10999 ( .B1(n10164), .B2(n10320), .A(n10163), .ZN(n10165) );
  OAI21_X1 U11000 ( .B1(n10322), .B2(n10309), .A(n10165), .ZN(P1_U3266) );
  OAI21_X1 U11001 ( .B1(n10167), .B2(n10169), .A(n10166), .ZN(n10168) );
  INV_X1 U11002 ( .A(n10168), .ZN(n10329) );
  XNOR2_X1 U11003 ( .A(n10170), .B(n10169), .ZN(n10331) );
  NAND2_X1 U11004 ( .A1(n10331), .A2(n11075), .ZN(n10180) );
  NAND2_X1 U11005 ( .A1(n10283), .A2(n10325), .ZN(n10173) );
  AOI22_X1 U11006 ( .A1(n11069), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n10171), 
        .B2(n11067), .ZN(n10172) );
  OAI211_X1 U11007 ( .C1(n10174), .C2(n10287), .A(n10173), .B(n10172), .ZN(
        n10177) );
  INV_X1 U11008 ( .A(n10189), .ZN(n10175) );
  OAI211_X1 U11009 ( .C1(n5398), .C2(n10175), .A(n5150), .B(n10400), .ZN(
        n10327) );
  NOR2_X1 U11010 ( .A1(n10327), .A2(n10219), .ZN(n10176) );
  AOI211_X1 U11011 ( .C1(n10223), .C2(n10178), .A(n10177), .B(n10176), .ZN(
        n10179) );
  OAI211_X1 U11012 ( .C1(n10329), .C2(n10292), .A(n10180), .B(n10179), .ZN(
        P1_U3267) );
  INV_X1 U11013 ( .A(n10181), .ZN(n10182) );
  AOI21_X1 U11014 ( .B1(n10183), .B2(n10184), .A(n10182), .ZN(n10337) );
  XNOR2_X1 U11015 ( .A(n10185), .B(n10184), .ZN(n10339) );
  NAND2_X1 U11016 ( .A1(n10339), .A2(n11075), .ZN(n10194) );
  NAND2_X1 U11017 ( .A1(n10283), .A2(n10347), .ZN(n10188) );
  AOI22_X1 U11018 ( .A1(n11069), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n10186), 
        .B2(n11067), .ZN(n10187) );
  OAI211_X1 U11019 ( .C1(n10317), .C2(n10287), .A(n10188), .B(n10187), .ZN(
        n10191) );
  OAI211_X1 U11020 ( .C1(n10441), .C2(n5153), .A(n10400), .B(n10189), .ZN(
        n10335) );
  NOR2_X1 U11021 ( .A1(n10335), .A2(n10219), .ZN(n10190) );
  AOI211_X1 U11022 ( .C1(n10223), .C2(n10192), .A(n10191), .B(n10190), .ZN(
        n10193) );
  OAI211_X1 U11023 ( .C1(n10337), .C2(n10292), .A(n10194), .B(n10193), .ZN(
        P1_U3268) );
  OAI211_X1 U11024 ( .C1(n5196), .C2(n10198), .A(n10195), .B(n10411), .ZN(
        n10197) );
  AOI22_X1 U11025 ( .A1(n11089), .A2(n10230), .B1(n11088), .B2(n10325), .ZN(
        n10196) );
  NAND2_X1 U11026 ( .A1(n10197), .A2(n10196), .ZN(n10342) );
  INV_X1 U11027 ( .A(n10342), .ZN(n10207) );
  XNOR2_X1 U11028 ( .A(n10199), .B(n10198), .ZN(n10344) );
  NAND2_X1 U11029 ( .A1(n10344), .A2(n11075), .ZN(n10206) );
  INV_X1 U11030 ( .A(n10200), .ZN(n10218) );
  AOI211_X1 U11031 ( .C1(n10201), .C2(n10218), .A(n10300), .B(n5153), .ZN(
        n10343) );
  AOI22_X1 U11032 ( .A1(n11069), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n10202), 
        .B2(n11067), .ZN(n10203) );
  OAI21_X1 U11033 ( .B1(n10445), .B2(n11072), .A(n10203), .ZN(n10204) );
  AOI21_X1 U11034 ( .B1(n10343), .B2(n11065), .A(n10204), .ZN(n10205) );
  OAI211_X1 U11035 ( .C1(n11069), .C2(n10207), .A(n10206), .B(n10205), .ZN(
        P1_U3269) );
  NAND2_X1 U11036 ( .A1(n10227), .A2(n10208), .ZN(n10211) );
  INV_X1 U11037 ( .A(n10209), .ZN(n10210) );
  AOI21_X1 U11038 ( .B1(n10212), .B2(n10211), .A(n10210), .ZN(n10351) );
  XNOR2_X1 U11039 ( .A(n10213), .B(n10212), .ZN(n10353) );
  NAND2_X1 U11040 ( .A1(n10353), .A2(n11075), .ZN(n10225) );
  NAND2_X1 U11041 ( .A1(n10283), .A2(n10348), .ZN(n10216) );
  AOI22_X1 U11042 ( .A1(n11079), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n10214), 
        .B2(n11067), .ZN(n10215) );
  OAI211_X1 U11043 ( .C1(n10217), .C2(n10287), .A(n10216), .B(n10215), .ZN(
        n10221) );
  OAI211_X1 U11044 ( .C1(n10449), .C2(n10236), .A(n10218), .B(n10400), .ZN(
        n10349) );
  NOR2_X1 U11045 ( .A1(n10349), .A2(n10219), .ZN(n10220) );
  AOI211_X1 U11046 ( .C1(n10223), .C2(n10222), .A(n10221), .B(n10220), .ZN(
        n10224) );
  OAI211_X1 U11047 ( .C1(n10351), .C2(n10292), .A(n10225), .B(n10224), .ZN(
        P1_U3270) );
  INV_X1 U11048 ( .A(n10234), .ZN(n10229) );
  INV_X1 U11049 ( .A(n10226), .ZN(n10228) );
  OAI211_X1 U11050 ( .C1(n10229), .C2(n10228), .A(n10227), .B(n10411), .ZN(
        n10233) );
  AOI22_X1 U11051 ( .A1(n10231), .A2(n11089), .B1(n11088), .B2(n10230), .ZN(
        n10232) );
  NAND2_X1 U11052 ( .A1(n10233), .A2(n10232), .ZN(n10356) );
  INV_X1 U11053 ( .A(n10356), .ZN(n10243) );
  XNOR2_X1 U11054 ( .A(n10235), .B(n10234), .ZN(n10358) );
  NAND2_X1 U11055 ( .A1(n10358), .A2(n11075), .ZN(n10242) );
  AOI211_X1 U11056 ( .C1(n10237), .C2(n10251), .A(n10300), .B(n10236), .ZN(
        n10357) );
  AOI22_X1 U11057 ( .A1(n11079), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n10238), 
        .B2(n11067), .ZN(n10239) );
  OAI21_X1 U11058 ( .B1(n10453), .B2(n11072), .A(n10239), .ZN(n10240) );
  AOI21_X1 U11059 ( .B1(n10357), .B2(n11065), .A(n10240), .ZN(n10241) );
  OAI211_X1 U11060 ( .C1(n11069), .C2(n10243), .A(n10242), .B(n10241), .ZN(
        P1_U3271) );
  AOI21_X1 U11061 ( .B1(n10271), .B2(n10269), .A(n10270), .ZN(n10275) );
  INV_X1 U11062 ( .A(n10244), .ZN(n10245) );
  NOR2_X1 U11063 ( .A1(n10275), .A2(n10245), .ZN(n10246) );
  XNOR2_X1 U11064 ( .A(n10246), .B(n10249), .ZN(n10247) );
  OAI222_X1 U11065 ( .A1(n10375), .A2(n10248), .B1(n10388), .B2(n10376), .C1(
        n11022), .C2(n10247), .ZN(n10361) );
  INV_X1 U11066 ( .A(n10361), .ZN(n10259) );
  XNOR2_X1 U11067 ( .A(n10250), .B(n10249), .ZN(n10363) );
  NAND2_X1 U11068 ( .A1(n10363), .A2(n11075), .ZN(n10258) );
  INV_X1 U11069 ( .A(n10251), .ZN(n10252) );
  AOI211_X1 U11070 ( .C1(n10253), .C2(n10261), .A(n10300), .B(n10252), .ZN(
        n10362) );
  AOI22_X1 U11071 ( .A1(n11079), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n10254), 
        .B2(n11067), .ZN(n10255) );
  OAI21_X1 U11072 ( .B1(n10458), .B2(n11072), .A(n10255), .ZN(n10256) );
  AOI21_X1 U11073 ( .B1(n10362), .B2(n11065), .A(n10256), .ZN(n10257) );
  OAI211_X1 U11074 ( .C1(n11069), .C2(n10259), .A(n10258), .B(n10257), .ZN(
        P1_U3272) );
  XOR2_X1 U11075 ( .A(n10260), .B(n10270), .Z(n10373) );
  INV_X1 U11076 ( .A(n10261), .ZN(n10262) );
  AOI211_X1 U11077 ( .C1(n10263), .C2(n5403), .A(n10300), .B(n10262), .ZN(
        n10370) );
  AOI22_X1 U11078 ( .A1(n11079), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n10264), 
        .B2(n11067), .ZN(n10267) );
  NAND2_X1 U11079 ( .A1(n10283), .A2(n10265), .ZN(n10266) );
  OAI211_X1 U11080 ( .C1(n10368), .C2(n11072), .A(n10267), .B(n10266), .ZN(
        n10268) );
  AOI21_X1 U11081 ( .B1(n10370), .B2(n11065), .A(n10268), .ZN(n10277) );
  NAND3_X1 U11082 ( .A1(n10271), .A2(n10270), .A3(n10269), .ZN(n10272) );
  NAND2_X1 U11083 ( .A1(n10272), .A2(n10411), .ZN(n10274) );
  OAI22_X1 U11084 ( .A1(n10275), .A2(n10274), .B1(n10273), .B2(n10375), .ZN(
        n10371) );
  NAND2_X1 U11085 ( .A1(n10371), .A2(n10307), .ZN(n10276) );
  OAI211_X1 U11086 ( .C1(n10373), .C2(n10309), .A(n10277), .B(n10276), .ZN(
        P1_U3273) );
  XNOR2_X1 U11087 ( .A(n10278), .B(n10279), .ZN(n10382) );
  XNOR2_X1 U11088 ( .A(n10280), .B(n10279), .ZN(n10374) );
  NAND2_X1 U11089 ( .A1(n10374), .A2(n11075), .ZN(n10291) );
  AOI211_X1 U11090 ( .C1(n10379), .C2(n10298), .A(n10300), .B(n10281), .ZN(
        n10377) );
  NOR2_X1 U11091 ( .A1(n5401), .A2(n11072), .ZN(n10289) );
  NAND2_X1 U11092 ( .A1(n10283), .A2(n10282), .ZN(n10286) );
  AOI22_X1 U11093 ( .A1(n11079), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n10284), 
        .B2(n11067), .ZN(n10285) );
  OAI211_X1 U11094 ( .C1(n10376), .C2(n10287), .A(n10286), .B(n10285), .ZN(
        n10288) );
  AOI211_X1 U11095 ( .C1(n10377), .C2(n11065), .A(n10289), .B(n10288), .ZN(
        n10290) );
  OAI211_X1 U11096 ( .C1(n10382), .C2(n10292), .A(n10291), .B(n10290), .ZN(
        P1_U3274) );
  XOR2_X1 U11097 ( .A(n10293), .B(n10294), .Z(n10387) );
  XNOR2_X1 U11098 ( .A(n10295), .B(n10294), .ZN(n10296) );
  OAI222_X1 U11099 ( .A1(n10375), .A2(n10367), .B1(n10388), .B2(n10297), .C1(
        n10296), .C2(n11022), .ZN(n10383) );
  INV_X1 U11100 ( .A(n10298), .ZN(n10299) );
  AOI211_X1 U11101 ( .C1(n10385), .C2(n10301), .A(n10300), .B(n10299), .ZN(
        n10384) );
  NAND2_X1 U11102 ( .A1(n10384), .A2(n11065), .ZN(n10304) );
  AOI22_X1 U11103 ( .A1(n11079), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n10302), 
        .B2(n11067), .ZN(n10303) );
  OAI211_X1 U11104 ( .C1(n10305), .C2(n11072), .A(n10304), .B(n10303), .ZN(
        n10306) );
  AOI21_X1 U11105 ( .B1(n10383), .B2(n10307), .A(n10306), .ZN(n10308) );
  OAI21_X1 U11106 ( .B1(n10387), .B2(n10309), .A(n10308), .ZN(P1_U3275) );
  OAI21_X1 U11107 ( .B1(n10426), .B2(n10366), .A(n10311), .ZN(P1_U3553) );
  INV_X1 U11108 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n10314) );
  NOR2_X1 U11109 ( .A1(n10313), .A2(n10312), .ZN(n10427) );
  MUX2_X1 U11110 ( .A(n10314), .B(n10427), .S(n11110), .Z(n10315) );
  OAI21_X1 U11111 ( .B1(n10430), .B2(n10366), .A(n10315), .ZN(P1_U3552) );
  OAI22_X1 U11112 ( .A1(n10317), .A2(n10388), .B1(n10316), .B2(n10375), .ZN(
        n10319) );
  AOI211_X1 U11113 ( .C1(n10411), .C2(n10320), .A(n10319), .B(n10318), .ZN(
        n10321) );
  OAI21_X1 U11114 ( .B1(n10322), .B2(n11023), .A(n10321), .ZN(n10431) );
  MUX2_X1 U11115 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10431), .S(n11110), .Z(
        n10323) );
  INV_X1 U11116 ( .A(n10323), .ZN(n10324) );
  OAI21_X1 U11117 ( .B1(n10434), .B2(n10366), .A(n10324), .ZN(P1_U3549) );
  INV_X1 U11118 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n10332) );
  AOI22_X1 U11119 ( .A1(n10326), .A2(n11088), .B1(n11089), .B2(n10325), .ZN(
        n10328) );
  OAI211_X1 U11120 ( .C1(n10329), .C2(n11022), .A(n10328), .B(n10327), .ZN(
        n10330) );
  AOI21_X1 U11121 ( .B1(n10331), .B2(n11107), .A(n10330), .ZN(n10435) );
  MUX2_X1 U11122 ( .A(n10332), .B(n10435), .S(n11110), .Z(n10333) );
  OAI21_X1 U11123 ( .B1(n5398), .B2(n10366), .A(n10333), .ZN(P1_U3548) );
  INV_X1 U11124 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n10340) );
  AOI22_X1 U11125 ( .A1(n11089), .A2(n10347), .B1(n10334), .B2(n11088), .ZN(
        n10336) );
  OAI211_X1 U11126 ( .C1(n10337), .C2(n11022), .A(n10336), .B(n10335), .ZN(
        n10338) );
  AOI21_X1 U11127 ( .B1(n10339), .B2(n11107), .A(n10338), .ZN(n10438) );
  MUX2_X1 U11128 ( .A(n10340), .B(n10438), .S(n11110), .Z(n10341) );
  OAI21_X1 U11129 ( .B1(n10441), .B2(n10366), .A(n10341), .ZN(P1_U3547) );
  INV_X1 U11130 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n10345) );
  AOI211_X1 U11131 ( .C1(n10344), .C2(n11107), .A(n10343), .B(n10342), .ZN(
        n10442) );
  MUX2_X1 U11132 ( .A(n10345), .B(n10442), .S(n11110), .Z(n10346) );
  OAI21_X1 U11133 ( .B1(n10445), .B2(n10366), .A(n10346), .ZN(P1_U3546) );
  INV_X1 U11134 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n10354) );
  AOI22_X1 U11135 ( .A1(n11089), .A2(n10348), .B1(n10347), .B2(n11088), .ZN(
        n10350) );
  OAI211_X1 U11136 ( .C1(n10351), .C2(n11022), .A(n10350), .B(n10349), .ZN(
        n10352) );
  AOI21_X1 U11137 ( .B1(n10353), .B2(n11107), .A(n10352), .ZN(n10446) );
  MUX2_X1 U11138 ( .A(n10354), .B(n10446), .S(n11110), .Z(n10355) );
  OAI21_X1 U11139 ( .B1(n10449), .B2(n10366), .A(n10355), .ZN(P1_U3545) );
  INV_X1 U11140 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n10359) );
  AOI211_X1 U11141 ( .C1(n10358), .C2(n11107), .A(n10357), .B(n10356), .ZN(
        n10450) );
  MUX2_X1 U11142 ( .A(n10359), .B(n10450), .S(n11110), .Z(n10360) );
  OAI21_X1 U11143 ( .B1(n10453), .B2(n10366), .A(n10360), .ZN(P1_U3544) );
  INV_X1 U11144 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n10364) );
  AOI211_X1 U11145 ( .C1(n10363), .C2(n11107), .A(n10362), .B(n10361), .ZN(
        n10454) );
  MUX2_X1 U11146 ( .A(n10364), .B(n10454), .S(n11110), .Z(n10365) );
  OAI21_X1 U11147 ( .B1(n10458), .B2(n10366), .A(n10365), .ZN(P1_U3543) );
  OAI22_X1 U11148 ( .A1(n10368), .A2(n11103), .B1(n10367), .B2(n10388), .ZN(
        n10369) );
  NOR3_X1 U11149 ( .A1(n10371), .A2(n10370), .A3(n10369), .ZN(n10372) );
  OAI21_X1 U11150 ( .B1(n10373), .B2(n11023), .A(n10372), .ZN(n10459) );
  MUX2_X1 U11151 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10459), .S(n11110), .Z(
        P1_U3542) );
  NAND2_X1 U11152 ( .A1(n10374), .A2(n11107), .ZN(n10381) );
  OAI22_X1 U11153 ( .A1(n6140), .A2(n10388), .B1(n10376), .B2(n10375), .ZN(
        n10378) );
  AOI211_X1 U11154 ( .C1(n10399), .C2(n10379), .A(n10378), .B(n10377), .ZN(
        n10380) );
  OAI211_X1 U11155 ( .C1(n11022), .C2(n10382), .A(n10381), .B(n10380), .ZN(
        n10460) );
  MUX2_X1 U11156 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10460), .S(n11110), .Z(
        P1_U3541) );
  AOI211_X1 U11157 ( .C1(n10399), .C2(n10385), .A(n10384), .B(n10383), .ZN(
        n10386) );
  OAI21_X1 U11158 ( .B1(n10387), .B2(n11023), .A(n10386), .ZN(n10461) );
  MUX2_X1 U11159 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10461), .S(n11110), .Z(
        P1_U3540) );
  OAI22_X1 U11160 ( .A1(n10390), .A2(n11103), .B1(n10389), .B2(n10388), .ZN(
        n10391) );
  NOR3_X1 U11161 ( .A1(n10393), .A2(n10392), .A3(n10391), .ZN(n10394) );
  OAI21_X1 U11162 ( .B1(n10395), .B2(n11023), .A(n10394), .ZN(n10462) );
  MUX2_X1 U11163 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10462), .S(n11110), .Z(
        P1_U3539) );
  NAND3_X1 U11164 ( .A1(n10397), .A2(n10396), .A3(n11107), .ZN(n10404) );
  AOI22_X1 U11165 ( .A1(n10401), .A2(n10400), .B1(n10399), .B2(n10398), .ZN(
        n10402) );
  NAND3_X1 U11166 ( .A1(n10404), .A2(n10403), .A3(n10402), .ZN(n10463) );
  MUX2_X1 U11167 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10463), .S(n11110), .Z(
        P1_U3538) );
  AOI22_X1 U11168 ( .A1(n11089), .A2(n10406), .B1(n10405), .B2(n11088), .ZN(
        n10407) );
  OAI211_X1 U11169 ( .C1(n10409), .C2(n11103), .A(n10408), .B(n10407), .ZN(
        n10410) );
  AOI21_X1 U11170 ( .B1(n10412), .B2(n10411), .A(n10410), .ZN(n10413) );
  OAI21_X1 U11171 ( .B1(n10414), .B2(n11023), .A(n10413), .ZN(n10464) );
  MUX2_X1 U11172 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n10464), .S(n11110), .Z(
        P1_U3537) );
  AOI22_X1 U11173 ( .A1(n5697), .A2(n11088), .B1(n11089), .B2(n10415), .ZN(
        n10416) );
  OAI211_X1 U11174 ( .C1(n10418), .C2(n11103), .A(n10417), .B(n10416), .ZN(
        n10419) );
  INV_X1 U11175 ( .A(n10419), .ZN(n10421) );
  OAI211_X1 U11176 ( .C1(n10422), .C2(n11023), .A(n10421), .B(n10420), .ZN(
        n10465) );
  MUX2_X1 U11177 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10465), .S(n11110), .Z(
        P1_U3536) );
  INV_X1 U11178 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n10424) );
  MUX2_X1 U11179 ( .A(n10424), .B(n10423), .S(n11114), .Z(n10425) );
  OAI21_X1 U11180 ( .B1(n10426), .B2(n10457), .A(n10425), .ZN(P1_U3521) );
  INV_X1 U11181 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10428) );
  MUX2_X1 U11182 ( .A(n10428), .B(n10427), .S(n11114), .Z(n10429) );
  OAI21_X1 U11183 ( .B1(n10430), .B2(n10457), .A(n10429), .ZN(P1_U3520) );
  MUX2_X1 U11184 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10431), .S(n11114), .Z(
        n10432) );
  INV_X1 U11185 ( .A(n10432), .ZN(n10433) );
  OAI21_X1 U11186 ( .B1(n10434), .B2(n10457), .A(n10433), .ZN(P1_U3517) );
  INV_X1 U11187 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n10436) );
  MUX2_X1 U11188 ( .A(n10436), .B(n10435), .S(n11114), .Z(n10437) );
  OAI21_X1 U11189 ( .B1(n5398), .B2(n10457), .A(n10437), .ZN(P1_U3516) );
  INV_X1 U11190 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n10439) );
  MUX2_X1 U11191 ( .A(n10439), .B(n10438), .S(n11114), .Z(n10440) );
  OAI21_X1 U11192 ( .B1(n10441), .B2(n10457), .A(n10440), .ZN(P1_U3515) );
  INV_X1 U11193 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n10443) );
  MUX2_X1 U11194 ( .A(n10443), .B(n10442), .S(n11114), .Z(n10444) );
  OAI21_X1 U11195 ( .B1(n10445), .B2(n10457), .A(n10444), .ZN(P1_U3514) );
  INV_X1 U11196 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n10447) );
  MUX2_X1 U11197 ( .A(n10447), .B(n10446), .S(n11114), .Z(n10448) );
  OAI21_X1 U11198 ( .B1(n10449), .B2(n10457), .A(n10448), .ZN(P1_U3513) );
  INV_X1 U11199 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n10451) );
  MUX2_X1 U11200 ( .A(n10451), .B(n10450), .S(n11114), .Z(n10452) );
  OAI21_X1 U11201 ( .B1(n10453), .B2(n10457), .A(n10452), .ZN(P1_U3512) );
  INV_X1 U11202 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n10455) );
  MUX2_X1 U11203 ( .A(n10455), .B(n10454), .S(n11114), .Z(n10456) );
  OAI21_X1 U11204 ( .B1(n10458), .B2(n10457), .A(n10456), .ZN(P1_U3511) );
  MUX2_X1 U11205 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10459), .S(n11114), .Z(
        P1_U3510) );
  MUX2_X1 U11206 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10460), .S(n11114), .Z(
        P1_U3509) );
  MUX2_X1 U11207 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10461), .S(n11114), .Z(
        P1_U3507) );
  MUX2_X1 U11208 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10462), .S(n11114), .Z(
        P1_U3504) );
  MUX2_X1 U11209 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10463), .S(n11114), .Z(
        P1_U3501) );
  MUX2_X1 U11210 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n10464), .S(n11114), .Z(
        P1_U3498) );
  MUX2_X1 U11211 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10465), .S(n11114), .Z(
        P1_U3495) );
  AND2_X1 U11212 ( .A1(n10468), .A2(n10466), .ZN(n10480) );
  MUX2_X1 U11213 ( .A(P1_D_REG_1__SCAN_IN), .B(n10467), .S(n10480), .Z(
        P1_U3440) );
  MUX2_X1 U11214 ( .A(P1_D_REG_0__SCAN_IN), .B(n10469), .S(n10468), .Z(
        P1_U3439) );
  NAND3_X1 U11215 ( .A1(n10470), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n10473) );
  OAI22_X1 U11216 ( .A1(n10474), .A2(n10473), .B1(n10472), .B2(n10471), .ZN(
        n10475) );
  AOI21_X1 U11217 ( .B1(n10477), .B2(n10476), .A(n10475), .ZN(n10478) );
  INV_X1 U11218 ( .A(n10478), .ZN(P1_U3324) );
  MUX2_X1 U11219 ( .A(n10479), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AND2_X1 U11220 ( .A1(n10481), .A2(P1_D_REG_2__SCAN_IN), .ZN(P1_U3323) );
  AND2_X1 U11221 ( .A1(n10481), .A2(P1_D_REG_3__SCAN_IN), .ZN(P1_U3322) );
  INV_X1 U11222 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10842) );
  NOR2_X1 U11223 ( .A1(n10480), .A2(n10842), .ZN(P1_U3321) );
  AND2_X1 U11224 ( .A1(n10481), .A2(P1_D_REG_5__SCAN_IN), .ZN(P1_U3320) );
  AND2_X1 U11225 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10481), .ZN(P1_U3319) );
  AND2_X1 U11226 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10481), .ZN(P1_U3318) );
  AND2_X1 U11227 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10481), .ZN(P1_U3317) );
  AND2_X1 U11228 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10481), .ZN(P1_U3316) );
  AND2_X1 U11229 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10481), .ZN(P1_U3315) );
  AND2_X1 U11230 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10481), .ZN(P1_U3314) );
  AND2_X1 U11231 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10481), .ZN(P1_U3313) );
  AND2_X1 U11232 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10481), .ZN(P1_U3312) );
  AND2_X1 U11233 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10481), .ZN(P1_U3311) );
  AND2_X1 U11234 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10481), .ZN(P1_U3310) );
  AND2_X1 U11235 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10481), .ZN(P1_U3309) );
  AND2_X1 U11236 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10481), .ZN(P1_U3308) );
  AND2_X1 U11237 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10481), .ZN(P1_U3307) );
  AND2_X1 U11238 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10481), .ZN(P1_U3306) );
  AND2_X1 U11239 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10481), .ZN(P1_U3305) );
  AND2_X1 U11240 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10481), .ZN(P1_U3304) );
  AND2_X1 U11241 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10481), .ZN(P1_U3303) );
  AND2_X1 U11242 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10481), .ZN(P1_U3302) );
  AND2_X1 U11243 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10481), .ZN(P1_U3301) );
  AND2_X1 U11244 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10481), .ZN(P1_U3300) );
  AND2_X1 U11245 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10481), .ZN(P1_U3299) );
  AND2_X1 U11246 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10481), .ZN(P1_U3298) );
  AND2_X1 U11247 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10481), .ZN(P1_U3297) );
  AND2_X1 U11248 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10481), .ZN(P1_U3296) );
  AND2_X1 U11249 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10481), .ZN(P1_U3295) );
  AND2_X1 U11250 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10481), .ZN(P1_U3294) );
  INV_X1 U11251 ( .A(keyinput_88), .ZN(n10597) );
  OAI22_X1 U11252 ( .A1(n10655), .A2(keyinput_84), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(keyinput_83), .ZN(n10482) );
  AOI221_X1 U11253 ( .B1(n10655), .B2(keyinput_84), .C1(keyinput_83), .C2(
        P2_DATAO_REG_13__SCAN_IN), .A(n10482), .ZN(n10590) );
  OAI22_X1 U11254 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(keyinput_77), .B1(
        keyinput_78), .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n10483) );
  AOI221_X1 U11255 ( .B1(P2_DATAO_REG_19__SCAN_IN), .B2(keyinput_77), .C1(
        P2_DATAO_REG_18__SCAN_IN), .C2(keyinput_78), .A(n10483), .ZN(n10586)
         );
  OAI22_X1 U11256 ( .A1(n10485), .A2(keyinput_70), .B1(keyinput_69), .B2(
        P2_DATAO_REG_27__SCAN_IN), .ZN(n10484) );
  AOI221_X1 U11257 ( .B1(n10485), .B2(keyinput_70), .C1(
        P2_DATAO_REG_27__SCAN_IN), .C2(keyinput_69), .A(n10484), .ZN(n10577)
         );
  INV_X1 U11258 ( .A(keyinput_68), .ZN(n10576) );
  INV_X1 U11259 ( .A(keyinput_67), .ZN(n10575) );
  INV_X1 U11260 ( .A(keyinput_66), .ZN(n10574) );
  OAI22_X1 U11261 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(keyinput_51), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(keyinput_50), .ZN(n10486) );
  AOI221_X1 U11262 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_51), .C1(
        keyinput_50), .C2(P2_REG3_REG_17__SCAN_IN), .A(n10486), .ZN(n10558) );
  INV_X1 U11263 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n10659) );
  OAI22_X1 U11264 ( .A1(n10659), .A2(keyinput_47), .B1(keyinput_48), .B2(
        P2_REG3_REG_16__SCAN_IN), .ZN(n10487) );
  AOI221_X1 U11265 ( .B1(n10659), .B2(keyinput_47), .C1(
        P2_REG3_REG_16__SCAN_IN), .C2(keyinput_48), .A(n10487), .ZN(n10554) );
  INV_X1 U11266 ( .A(keyinput_41), .ZN(n10546) );
  AOI22_X1 U11267 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(keyinput_38), .B1(n10661), .B2(keyinput_39), .ZN(n10488) );
  OAI221_X1 U11268 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(keyinput_38), .C1(
        n10661), .C2(keyinput_39), .A(n10488), .ZN(n10545) );
  INV_X1 U11269 ( .A(keyinput_37), .ZN(n10544) );
  INV_X1 U11270 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n10722) );
  AOI22_X1 U11271 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(keyinput_35), .B1(
        P2_STATE_REG_SCAN_IN), .B2(keyinput_34), .ZN(n10489) );
  OAI221_X1 U11272 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(keyinput_35), .C1(
        P2_STATE_REG_SCAN_IN), .C2(keyinput_34), .A(n10489), .ZN(n10541) );
  INV_X1 U11273 ( .A(keyinput_33), .ZN(n10539) );
  INV_X1 U11274 ( .A(P2_RD_REG_SCAN_IN), .ZN(n11020) );
  OAI22_X1 U11275 ( .A1(n10491), .A2(keyinput_21), .B1(SI_12_), .B2(
        keyinput_20), .ZN(n10490) );
  AOI221_X1 U11276 ( .B1(n10491), .B2(keyinput_21), .C1(keyinput_20), .C2(
        SI_12_), .A(n10490), .ZN(n10522) );
  INV_X1 U11277 ( .A(keyinput_12), .ZN(n10509) );
  INV_X1 U11278 ( .A(keyinput_11), .ZN(n10508) );
  AOI22_X1 U11279 ( .A1(SI_23_), .A2(keyinput_9), .B1(n10493), .B2(keyinput_8), 
        .ZN(n10492) );
  OAI221_X1 U11280 ( .B1(SI_23_), .B2(keyinput_9), .C1(n10493), .C2(keyinput_8), .A(n10492), .ZN(n10505) );
  AOI22_X1 U11281 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_0), .B1(SI_31_), .B2(
        keyinput_1), .ZN(n10494) );
  OAI221_X1 U11282 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_0), .C1(SI_31_), 
        .C2(keyinput_1), .A(n10494), .ZN(n10503) );
  AOI22_X1 U11283 ( .A1(SI_28_), .A2(keyinput_4), .B1(n10675), .B2(keyinput_7), 
        .ZN(n10495) );
  OAI221_X1 U11284 ( .B1(SI_28_), .B2(keyinput_4), .C1(n10675), .C2(keyinput_7), .A(n10495), .ZN(n10502) );
  AOI22_X1 U11285 ( .A1(n10497), .A2(keyinput_3), .B1(n10673), .B2(keyinput_6), 
        .ZN(n10496) );
  OAI221_X1 U11286 ( .B1(n10497), .B2(keyinput_3), .C1(n10673), .C2(keyinput_6), .A(n10496), .ZN(n10501) );
  INV_X1 U11287 ( .A(SI_30_), .ZN(n10499) );
  AOI22_X1 U11288 ( .A1(n10676), .A2(keyinput_5), .B1(keyinput_2), .B2(n10499), 
        .ZN(n10498) );
  OAI221_X1 U11289 ( .B1(n10676), .B2(keyinput_5), .C1(n10499), .C2(keyinput_2), .A(n10498), .ZN(n10500) );
  NOR4_X1 U11290 ( .A1(n10503), .A2(n10502), .A3(n10501), .A4(n10500), .ZN(
        n10504) );
  OAI22_X1 U11291 ( .A1(n10505), .A2(n10504), .B1(keyinput_10), .B2(SI_22_), 
        .ZN(n10506) );
  AOI21_X1 U11292 ( .B1(keyinput_10), .B2(SI_22_), .A(n10506), .ZN(n10507) );
  AOI22_X1 U11293 ( .A1(SI_18_), .A2(keyinput_14), .B1(SI_19_), .B2(
        keyinput_13), .ZN(n10510) );
  OAI221_X1 U11294 ( .B1(SI_18_), .B2(keyinput_14), .C1(SI_19_), .C2(
        keyinput_13), .A(n10510), .ZN(n10511) );
  XOR2_X1 U11295 ( .A(SI_16_), .B(keyinput_16), .Z(n10512) );
  OAI22_X1 U11296 ( .A1(n10513), .A2(n10512), .B1(SI_15_), .B2(keyinput_17), 
        .ZN(n10516) );
  OAI22_X1 U11297 ( .A1(SI_14_), .A2(keyinput_18), .B1(SI_13_), .B2(
        keyinput_19), .ZN(n10514) );
  AOI221_X1 U11298 ( .B1(SI_14_), .B2(keyinput_18), .C1(keyinput_19), .C2(
        SI_13_), .A(n10514), .ZN(n10515) );
  OAI221_X1 U11299 ( .B1(n10516), .B2(keyinput_17), .C1(n10516), .C2(SI_15_), 
        .A(n10515), .ZN(n10521) );
  INV_X1 U11300 ( .A(SI_10_), .ZN(n10698) );
  XNOR2_X1 U11301 ( .A(n10698), .B(keyinput_22), .ZN(n10520) );
  AOI22_X1 U11302 ( .A1(SI_9_), .A2(keyinput_23), .B1(n10518), .B2(keyinput_24), .ZN(n10517) );
  OAI221_X1 U11303 ( .B1(SI_9_), .B2(keyinput_23), .C1(n10518), .C2(
        keyinput_24), .A(n10517), .ZN(n10519) );
  AOI211_X1 U11304 ( .C1(n10522), .C2(n10521), .A(n10520), .B(n10519), .ZN(
        n10523) );
  INV_X1 U11305 ( .A(n10523), .ZN(n10534) );
  AOI22_X1 U11306 ( .A1(SI_2_), .A2(keyinput_30), .B1(SI_5_), .B2(keyinput_27), 
        .ZN(n10524) );
  OAI221_X1 U11307 ( .B1(SI_2_), .B2(keyinput_30), .C1(SI_5_), .C2(keyinput_27), .A(n10524), .ZN(n10530) );
  AOI22_X1 U11308 ( .A1(SI_3_), .A2(keyinput_29), .B1(SI_6_), .B2(keyinput_26), 
        .ZN(n10525) );
  OAI221_X1 U11309 ( .B1(SI_3_), .B2(keyinput_29), .C1(SI_6_), .C2(keyinput_26), .A(n10525), .ZN(n10529) );
  XNOR2_X1 U11310 ( .A(n10526), .B(keyinput_28), .ZN(n10528) );
  XOR2_X1 U11311 ( .A(SI_7_), .B(keyinput_25), .Z(n10527) );
  NOR4_X1 U11312 ( .A1(n10530), .A2(n10529), .A3(n10528), .A4(n10527), .ZN(
        n10533) );
  INV_X1 U11313 ( .A(keyinput_31), .ZN(n10531) );
  MUX2_X1 U11314 ( .A(n10531), .B(keyinput_31), .S(SI_1_), .Z(n10532) );
  AOI21_X1 U11315 ( .B1(n10534), .B2(n10533), .A(n10532), .ZN(n10537) );
  INV_X1 U11316 ( .A(keyinput_32), .ZN(n10535) );
  MUX2_X1 U11317 ( .A(n10535), .B(keyinput_32), .S(SI_0_), .Z(n10536) );
  NOR2_X1 U11318 ( .A1(n10537), .A2(n10536), .ZN(n10538) );
  AOI221_X1 U11319 ( .B1(P2_RD_REG_SCAN_IN), .B2(n10539), .C1(n11020), .C2(
        keyinput_33), .A(n10538), .ZN(n10540) );
  OAI22_X1 U11320 ( .A1(keyinput_36), .A2(n10722), .B1(n10541), .B2(n10540), 
        .ZN(n10542) );
  AOI21_X1 U11321 ( .B1(keyinput_36), .B2(n10722), .A(n10542), .ZN(n10543) );
  XNOR2_X1 U11322 ( .A(P2_REG3_REG_28__SCAN_IN), .B(keyinput_42), .ZN(n10551)
         );
  OAI22_X1 U11323 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(keyinput_45), .B1(
        keyinput_46), .B2(P2_REG3_REG_12__SCAN_IN), .ZN(n10547) );
  AOI221_X1 U11324 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_45), .C1(
        P2_REG3_REG_12__SCAN_IN), .C2(keyinput_46), .A(n10547), .ZN(n10550) );
  OAI22_X1 U11325 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_43), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(keyinput_44), .ZN(n10548) );
  AOI221_X1 U11326 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_43), .C1(
        keyinput_44), .C2(P2_REG3_REG_1__SCAN_IN), .A(n10548), .ZN(n10549) );
  OAI211_X1 U11327 ( .C1(n10552), .C2(n10551), .A(n10550), .B(n10549), .ZN(
        n10553) );
  AOI22_X1 U11328 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(keyinput_52), .B1(n10556), 
        .B2(keyinput_53), .ZN(n10555) );
  OAI221_X1 U11329 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput_52), .C1(n10556), .C2(keyinput_53), .A(n10555), .ZN(n10557) );
  AOI22_X1 U11330 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(keyinput_58), .B1(
        P2_REG3_REG_22__SCAN_IN), .B2(keyinput_57), .ZN(n10559) );
  OAI221_X1 U11331 ( .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput_58), .C1(
        P2_REG3_REG_22__SCAN_IN), .C2(keyinput_57), .A(n10559), .ZN(n10565) );
  AOI22_X1 U11332 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(keyinput_56), .B1(
        P2_REG3_REG_20__SCAN_IN), .B2(keyinput_55), .ZN(n10560) );
  OAI221_X1 U11333 ( .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput_56), .C1(
        P2_REG3_REG_20__SCAN_IN), .C2(keyinput_55), .A(n10560), .ZN(n10564) );
  AOI22_X1 U11334 ( .A1(n10562), .A2(keyinput_54), .B1(n7537), .B2(keyinput_59), .ZN(n10561) );
  OAI221_X1 U11335 ( .B1(n10562), .B2(keyinput_54), .C1(n7537), .C2(
        keyinput_59), .A(n10561), .ZN(n10563) );
  AOI22_X1 U11336 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput_61), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(keyinput_60), .ZN(n10566) );
  OAI221_X1 U11337 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_61), .C1(
        P2_REG3_REG_18__SCAN_IN), .C2(keyinput_60), .A(n10566), .ZN(n10571) );
  OAI22_X1 U11338 ( .A1(n10472), .A2(keyinput_65), .B1(keyinput_64), .B2(
        P2_B_REG_SCAN_IN), .ZN(n10567) );
  AOI221_X1 U11339 ( .B1(n10472), .B2(keyinput_65), .C1(P2_B_REG_SCAN_IN), 
        .C2(keyinput_64), .A(n10567), .ZN(n10570) );
  OAI22_X1 U11340 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(keyinput_62), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(keyinput_63), .ZN(n10568) );
  AOI221_X1 U11341 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_62), .C1(
        keyinput_63), .C2(P2_REG3_REG_15__SCAN_IN), .A(n10568), .ZN(n10569) );
  OAI211_X1 U11342 ( .C1(n10572), .C2(n10571), .A(n10570), .B(n10569), .ZN(
        n10573) );
  OAI21_X1 U11343 ( .B1(keyinput_73), .B2(n8116), .A(n10578), .ZN(n10584) );
  AOI22_X1 U11344 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(keyinput_72), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(keyinput_71), .ZN(n10579) );
  OAI221_X1 U11345 ( .B1(P2_DATAO_REG_24__SCAN_IN), .B2(keyinput_72), .C1(
        P2_DATAO_REG_25__SCAN_IN), .C2(keyinput_71), .A(n10579), .ZN(n10583)
         );
  OAI22_X1 U11346 ( .A1(n10581), .A2(keyinput_74), .B1(keyinput_75), .B2(
        P2_DATAO_REG_21__SCAN_IN), .ZN(n10580) );
  AOI221_X1 U11347 ( .B1(n10581), .B2(keyinput_74), .C1(
        P2_DATAO_REG_21__SCAN_IN), .C2(keyinput_75), .A(n10580), .ZN(n10582)
         );
  OAI21_X1 U11348 ( .B1(n10584), .B2(n10583), .A(n10582), .ZN(n10585) );
  AOI22_X1 U11349 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(keyinput_80), .B1(
        n10789), .B2(keyinput_79), .ZN(n10587) );
  OAI221_X1 U11350 ( .B1(P2_DATAO_REG_16__SCAN_IN), .B2(keyinput_80), .C1(
        n10789), .C2(keyinput_79), .A(n10587), .ZN(n10588) );
  OAI211_X1 U11351 ( .C1(P2_DATAO_REG_11__SCAN_IN), .C2(keyinput_85), .A(
        n10590), .B(n10589), .ZN(n10591) );
  OAI22_X1 U11352 ( .A1(n10593), .A2(keyinput_82), .B1(keyinput_86), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n10592) );
  AOI221_X1 U11353 ( .B1(n10593), .B2(keyinput_82), .C1(
        P2_DATAO_REG_10__SCAN_IN), .C2(keyinput_86), .A(n10592), .ZN(n10596)
         );
  NOR2_X1 U11354 ( .A1(n10595), .A2(keyinput_87), .ZN(n10594) );
  AOI22_X1 U11355 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(keyinput_91), .B1(
        P1_IR_REG_0__SCAN_IN), .B2(keyinput_90), .ZN(n10598) );
  OAI221_X1 U11356 ( .B1(P1_IR_REG_1__SCAN_IN), .B2(keyinput_91), .C1(
        P1_IR_REG_0__SCAN_IN), .C2(keyinput_90), .A(n10598), .ZN(n10601) );
  XOR2_X1 U11357 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_89), .Z(n10600) );
  XOR2_X1 U11358 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_92), .Z(n10599) );
  XOR2_X1 U11359 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_94), .Z(n10603) );
  XNOR2_X1 U11360 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_93), .ZN(n10602) );
  NOR3_X1 U11361 ( .A1(n10604), .A2(n10603), .A3(n10602), .ZN(n10609) );
  NAND2_X1 U11362 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(keyinput_95), .ZN(n10605)
         );
  OAI21_X1 U11363 ( .B1(P1_IR_REG_5__SCAN_IN), .B2(keyinput_95), .A(n10605), 
        .ZN(n10608) );
  INV_X1 U11364 ( .A(keyinput_96), .ZN(n10606) );
  MUX2_X1 U11365 ( .A(n10606), .B(keyinput_96), .S(P1_IR_REG_6__SCAN_IN), .Z(
        n10607) );
  OAI21_X1 U11366 ( .B1(n10609), .B2(n10608), .A(n10607), .ZN(n10614) );
  INV_X1 U11367 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n10610) );
  XNOR2_X1 U11368 ( .A(keyinput_97), .B(n10610), .ZN(n10613) );
  XOR2_X1 U11369 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_99), .Z(n10612) );
  XOR2_X1 U11370 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_98), .Z(n10611) );
  AOI211_X1 U11371 ( .C1(n10614), .C2(n10613), .A(n10612), .B(n10611), .ZN(
        n10622) );
  XOR2_X1 U11372 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_101), .Z(n10618) );
  XNOR2_X1 U11373 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_102), .ZN(n10617)
         );
  XNOR2_X1 U11374 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_103), .ZN(n10616)
         );
  XNOR2_X1 U11375 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_100), .ZN(n10615)
         );
  NAND4_X1 U11376 ( .A1(n10618), .A2(n10617), .A3(n10616), .A4(n10615), .ZN(
        n10621) );
  XNOR2_X1 U11377 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_105), .ZN(n10620)
         );
  XNOR2_X1 U11378 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_104), .ZN(n10619)
         );
  OAI211_X1 U11379 ( .C1(n10622), .C2(n10621), .A(n10620), .B(n10619), .ZN(
        n10626) );
  XNOR2_X1 U11380 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_106), .ZN(n10625)
         );
  OAI22_X1 U11381 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(keyinput_107), .B1(
        keyinput_108), .B2(P1_IR_REG_18__SCAN_IN), .ZN(n10623) );
  AOI221_X1 U11382 ( .B1(P1_IR_REG_17__SCAN_IN), .B2(keyinput_107), .C1(
        P1_IR_REG_18__SCAN_IN), .C2(keyinput_108), .A(n10623), .ZN(n10624) );
  NAND3_X1 U11383 ( .A1(n10626), .A2(n10625), .A3(n10624), .ZN(n10629) );
  INV_X1 U11384 ( .A(keyinput_109), .ZN(n10627) );
  MUX2_X1 U11385 ( .A(n10627), .B(keyinput_109), .S(P1_IR_REG_19__SCAN_IN), 
        .Z(n10628) );
  NAND2_X1 U11386 ( .A1(n10629), .A2(n10628), .ZN(n10632) );
  INV_X1 U11387 ( .A(keyinput_110), .ZN(n10630) );
  MUX2_X1 U11388 ( .A(n10630), .B(keyinput_110), .S(P1_IR_REG_20__SCAN_IN), 
        .Z(n10631) );
  NAND2_X1 U11389 ( .A1(n10632), .A2(n10631), .ZN(n10640) );
  OAI22_X1 U11390 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(keyinput_112), .B1(
        keyinput_111), .B2(P1_IR_REG_21__SCAN_IN), .ZN(n10633) );
  AOI221_X1 U11391 ( .B1(P1_IR_REG_22__SCAN_IN), .B2(keyinput_112), .C1(
        P1_IR_REG_21__SCAN_IN), .C2(keyinput_111), .A(n10633), .ZN(n10639) );
  XNOR2_X1 U11392 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_115), .ZN(n10637)
         );
  XNOR2_X1 U11393 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_116), .ZN(n10636)
         );
  XNOR2_X1 U11394 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_114), .ZN(n10635)
         );
  XNOR2_X1 U11395 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput_113), .ZN(n10634)
         );
  NAND4_X1 U11396 ( .A1(n10637), .A2(n10636), .A3(n10635), .A4(n10634), .ZN(
        n10638) );
  AOI21_X1 U11397 ( .B1(n10640), .B2(n10639), .A(n10638), .ZN(n10643) );
  XOR2_X1 U11398 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput_119), .Z(n10642) );
  XNOR2_X1 U11399 ( .A(n10842), .B(keyinput_126), .ZN(n10641) );
  NOR3_X1 U11400 ( .A1(n10643), .A2(n10642), .A3(n10641), .ZN(n10863) );
  INV_X1 U11401 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10645) );
  INV_X1 U11402 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10843) );
  AOI22_X1 U11403 ( .A1(n10645), .A2(keyinput_123), .B1(n10843), .B2(
        keyinput_122), .ZN(n10644) );
  OAI221_X1 U11404 ( .B1(n10645), .B2(keyinput_123), .C1(n10843), .C2(
        keyinput_122), .A(n10644), .ZN(n10653) );
  AOI22_X1 U11405 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(keyinput_117), .B1(
        P1_IR_REG_31__SCAN_IN), .B2(keyinput_121), .ZN(n10646) );
  OAI221_X1 U11406 ( .B1(P1_IR_REG_27__SCAN_IN), .B2(keyinput_117), .C1(
        P1_IR_REG_31__SCAN_IN), .C2(keyinput_121), .A(n10646), .ZN(n10652) );
  AOI22_X1 U11407 ( .A1(P1_D_REG_2__SCAN_IN), .A2(keyinput_124), .B1(
        P1_IR_REG_28__SCAN_IN), .B2(keyinput_118), .ZN(n10647) );
  OAI221_X1 U11408 ( .B1(P1_D_REG_2__SCAN_IN), .B2(keyinput_124), .C1(
        P1_IR_REG_28__SCAN_IN), .C2(keyinput_118), .A(n10647), .ZN(n10651) );
  XOR2_X1 U11409 ( .A(P1_D_REG_3__SCAN_IN), .B(keyinput_125), .Z(n10649) );
  XNOR2_X1 U11410 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_120), .ZN(n10648)
         );
  NAND2_X1 U11411 ( .A1(n10649), .A2(n10648), .ZN(n10650) );
  NOR4_X1 U11412 ( .A1(n10653), .A2(n10652), .A3(n10651), .A4(n10650), .ZN(
        n10862) );
  OAI22_X1 U11413 ( .A1(n10655), .A2(keyinput_212), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(keyinput_214), .ZN(n10654) );
  AOI221_X1 U11414 ( .B1(n10655), .B2(keyinput_212), .C1(keyinput_214), .C2(
        P2_DATAO_REG_10__SCAN_IN), .A(n10654), .ZN(n10790) );
  INV_X1 U11415 ( .A(keyinput_196), .ZN(n10769) );
  INV_X1 U11416 ( .A(keyinput_194), .ZN(n10761) );
  OAI22_X1 U11417 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(keyinput_179), .B1(
        keyinput_178), .B2(P2_REG3_REG_17__SCAN_IN), .ZN(n10656) );
  AOI221_X1 U11418 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_179), .C1(
        P2_REG3_REG_17__SCAN_IN), .C2(keyinput_178), .A(n10656), .ZN(n10742)
         );
  OAI22_X1 U11419 ( .A1(n10659), .A2(keyinput_175), .B1(n10658), .B2(
        keyinput_176), .ZN(n10657) );
  AOI221_X1 U11420 ( .B1(n10659), .B2(keyinput_175), .C1(keyinput_176), .C2(
        n10658), .A(n10657), .ZN(n10738) );
  INV_X1 U11421 ( .A(keyinput_169), .ZN(n10730) );
  AOI22_X1 U11422 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(keyinput_166), .B1(
        n10661), .B2(keyinput_167), .ZN(n10660) );
  OAI221_X1 U11423 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(keyinput_166), .C1(
        n10661), .C2(keyinput_167), .A(n10660), .ZN(n10726) );
  INV_X1 U11424 ( .A(keyinput_165), .ZN(n10723) );
  AOI22_X1 U11425 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(keyinput_163), .B1(
        P2_STATE_REG_SCAN_IN), .B2(keyinput_162), .ZN(n10662) );
  OAI221_X1 U11426 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(keyinput_163), .C1(
        P2_STATE_REG_SCAN_IN), .C2(keyinput_162), .A(n10662), .ZN(n10721) );
  INV_X1 U11427 ( .A(keyinput_161), .ZN(n10720) );
  OAI22_X1 U11428 ( .A1(n10664), .A2(keyinput_148), .B1(SI_11_), .B2(
        keyinput_149), .ZN(n10663) );
  AOI221_X1 U11429 ( .B1(n10664), .B2(keyinput_148), .C1(keyinput_149), .C2(
        SI_11_), .A(n10663), .ZN(n10702) );
  INV_X1 U11430 ( .A(SI_18_), .ZN(n10666) );
  AOI22_X1 U11431 ( .A1(n10667), .A2(keyinput_141), .B1(keyinput_142), .B2(
        n10666), .ZN(n10665) );
  OAI221_X1 U11432 ( .B1(n10667), .B2(keyinput_141), .C1(n10666), .C2(
        keyinput_142), .A(n10665), .ZN(n10688) );
  INV_X1 U11433 ( .A(keyinput_140), .ZN(n10686) );
  INV_X1 U11434 ( .A(keyinput_139), .ZN(n10683) );
  AOI22_X1 U11435 ( .A1(SI_24_), .A2(keyinput_136), .B1(n10669), .B2(
        keyinput_137), .ZN(n10668) );
  OAI221_X1 U11436 ( .B1(SI_24_), .B2(keyinput_136), .C1(n10669), .C2(
        keyinput_137), .A(n10668), .ZN(n10682) );
  AOI22_X1 U11437 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_128), .B1(SI_31_), 
        .B2(keyinput_129), .ZN(n10670) );
  OAI221_X1 U11438 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_128), .C1(SI_31_), 
        .C2(keyinput_129), .A(n10670), .ZN(n10680) );
  AOI22_X1 U11439 ( .A1(SI_30_), .A2(keyinput_130), .B1(SI_28_), .B2(
        keyinput_132), .ZN(n10671) );
  OAI221_X1 U11440 ( .B1(SI_30_), .B2(keyinput_130), .C1(SI_28_), .C2(
        keyinput_132), .A(n10671), .ZN(n10679) );
  AOI22_X1 U11441 ( .A1(SI_29_), .A2(keyinput_131), .B1(n10673), .B2(
        keyinput_134), .ZN(n10672) );
  OAI221_X1 U11442 ( .B1(SI_29_), .B2(keyinput_131), .C1(n10673), .C2(
        keyinput_134), .A(n10672), .ZN(n10678) );
  OAI221_X1 U11443 ( .B1(n10676), .B2(keyinput_133), .C1(n10675), .C2(
        keyinput_135), .A(n10674), .ZN(n10677) );
  OAI22_X1 U11444 ( .A1(keyinput_143), .A2(n10690), .B1(n10688), .B2(n10687), 
        .ZN(n10689) );
  XOR2_X1 U11445 ( .A(SI_16_), .B(keyinput_144), .Z(n10691) );
  OAI22_X1 U11446 ( .A1(n10695), .A2(keyinput_146), .B1(SI_13_), .B2(
        keyinput_147), .ZN(n10694) );
  AOI221_X1 U11447 ( .B1(n10695), .B2(keyinput_146), .C1(keyinput_147), .C2(
        SI_13_), .A(n10694), .ZN(n10696) );
  XOR2_X1 U11448 ( .A(SI_9_), .B(keyinput_151), .Z(n10700) );
  AOI22_X1 U11449 ( .A1(SI_8_), .A2(keyinput_152), .B1(n10698), .B2(
        keyinput_150), .ZN(n10697) );
  OAI221_X1 U11450 ( .B1(SI_8_), .B2(keyinput_152), .C1(n10698), .C2(
        keyinput_150), .A(n10697), .ZN(n10699) );
  AOI211_X1 U11451 ( .C1(n10702), .C2(n10701), .A(n10700), .B(n10699), .ZN(
        n10703) );
  INV_X1 U11452 ( .A(n10703), .ZN(n10715) );
  AOI22_X1 U11453 ( .A1(SI_4_), .A2(keyinput_156), .B1(SI_7_), .B2(
        keyinput_153), .ZN(n10704) );
  OAI221_X1 U11454 ( .B1(SI_4_), .B2(keyinput_156), .C1(SI_7_), .C2(
        keyinput_153), .A(n10704), .ZN(n10711) );
  AOI22_X1 U11455 ( .A1(SI_3_), .A2(keyinput_157), .B1(SI_5_), .B2(
        keyinput_155), .ZN(n10705) );
  OAI221_X1 U11456 ( .B1(SI_3_), .B2(keyinput_157), .C1(SI_5_), .C2(
        keyinput_155), .A(n10705), .ZN(n10710) );
  XNOR2_X1 U11457 ( .A(n10706), .B(keyinput_158), .ZN(n10709) );
  XNOR2_X1 U11458 ( .A(n10707), .B(keyinput_154), .ZN(n10708) );
  NOR4_X1 U11459 ( .A1(n10711), .A2(n10710), .A3(n10709), .A4(n10708), .ZN(
        n10714) );
  INV_X1 U11460 ( .A(keyinput_159), .ZN(n10712) );
  MUX2_X1 U11461 ( .A(keyinput_159), .B(n10712), .S(SI_1_), .Z(n10713) );
  AOI21_X1 U11462 ( .B1(n10715), .B2(n10714), .A(n10713), .ZN(n10718) );
  INV_X1 U11463 ( .A(keyinput_160), .ZN(n10716) );
  MUX2_X1 U11464 ( .A(keyinput_160), .B(n10716), .S(SI_0_), .Z(n10717) );
  OAI22_X1 U11465 ( .A1(n10726), .A2(n10725), .B1(keyinput_168), .B2(
        P2_REG3_REG_3__SCAN_IN), .ZN(n10727) );
  AOI21_X1 U11466 ( .B1(keyinput_168), .B2(P2_REG3_REG_3__SCAN_IN), .A(n10727), 
        .ZN(n10728) );
  AOI221_X1 U11467 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(n10730), .C1(n10729), 
        .C2(keyinput_169), .A(n10728), .ZN(n10737) );
  XNOR2_X1 U11468 ( .A(P2_REG3_REG_28__SCAN_IN), .B(keyinput_170), .ZN(n10736)
         );
  OAI22_X1 U11469 ( .A1(n10732), .A2(keyinput_174), .B1(n7546), .B2(
        keyinput_172), .ZN(n10731) );
  AOI221_X1 U11470 ( .B1(n10732), .B2(keyinput_174), .C1(keyinput_172), .C2(
        n7546), .A(n10731), .ZN(n10735) );
  OAI22_X1 U11471 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(keyinput_173), .B1(
        P2_REG3_REG_8__SCAN_IN), .B2(keyinput_171), .ZN(n10733) );
  AOI221_X1 U11472 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_173), .C1(
        keyinput_171), .C2(P2_REG3_REG_8__SCAN_IN), .A(n10733), .ZN(n10734) );
  INV_X1 U11473 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n10740) );
  AOI22_X1 U11474 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput_181), .B1(n10740), .B2(keyinput_180), .ZN(n10739) );
  OAI221_X1 U11475 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput_181), .C1(
        n10740), .C2(keyinput_180), .A(n10739), .ZN(n10741) );
  AOI22_X1 U11476 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(keyinput_183), .B1(
        P2_REG3_REG_22__SCAN_IN), .B2(keyinput_185), .ZN(n10743) );
  OAI221_X1 U11477 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput_183), .C1(
        P2_REG3_REG_22__SCAN_IN), .C2(keyinput_185), .A(n10743), .ZN(n10749)
         );
  AOI22_X1 U11478 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_182), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(keyinput_187), .ZN(n10744) );
  OAI221_X1 U11479 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_182), .C1(
        P2_REG3_REG_2__SCAN_IN), .C2(keyinput_187), .A(n10744), .ZN(n10748) );
  AOI22_X1 U11480 ( .A1(n11019), .A2(keyinput_186), .B1(n10746), .B2(
        keyinput_184), .ZN(n10745) );
  OAI221_X1 U11481 ( .B1(n11019), .B2(keyinput_186), .C1(n10746), .C2(
        keyinput_184), .A(n10745), .ZN(n10747) );
  AOI22_X1 U11482 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput_189), .B1(n10752), .B2(keyinput_188), .ZN(n10751) );
  OAI221_X1 U11483 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_189), .C1(
        n10752), .C2(keyinput_188), .A(n10751), .ZN(n10757) );
  OAI22_X1 U11484 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(keyinput_190), .B1(
        keyinput_193), .B2(P2_DATAO_REG_31__SCAN_IN), .ZN(n10753) );
  AOI221_X1 U11485 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_190), .C1(
        P2_DATAO_REG_31__SCAN_IN), .C2(keyinput_193), .A(n10753), .ZN(n10756)
         );
  OAI22_X1 U11486 ( .A1(P2_B_REG_SCAN_IN), .A2(keyinput_192), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(keyinput_191), .ZN(n10754) );
  AOI221_X1 U11487 ( .B1(P2_B_REG_SCAN_IN), .B2(keyinput_192), .C1(
        keyinput_191), .C2(P2_REG3_REG_15__SCAN_IN), .A(n10754), .ZN(n10755)
         );
  OAI211_X1 U11488 ( .C1(n10758), .C2(n10757), .A(n10756), .B(n10755), .ZN(
        n10759) );
  OAI221_X1 U11489 ( .B1(P2_DATAO_REG_30__SCAN_IN), .B2(n10761), .C1(n10760), 
        .C2(keyinput_194), .A(n10759), .ZN(n10766) );
  INV_X1 U11490 ( .A(keyinput_195), .ZN(n10762) );
  OAI221_X1 U11491 ( .B1(P2_DATAO_REG_28__SCAN_IN), .B2(n10769), .C1(n10768), 
        .C2(keyinput_196), .A(n10767), .ZN(n10772) );
  OAI22_X1 U11492 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(keyinput_197), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(keyinput_198), .ZN(n10770) );
  AOI221_X1 U11493 ( .B1(P2_DATAO_REG_27__SCAN_IN), .B2(keyinput_197), .C1(
        keyinput_198), .C2(P2_DATAO_REG_26__SCAN_IN), .A(n10770), .ZN(n10771)
         );
  AOI22_X1 U11494 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(keyinput_201), .B1(
        n10775), .B2(keyinput_199), .ZN(n10774) );
  OAI221_X1 U11495 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(keyinput_201), .C1(
        n10775), .C2(keyinput_199), .A(n10774), .ZN(n10779) );
  OAI22_X1 U11496 ( .A1(n10777), .A2(keyinput_203), .B1(keyinput_202), .B2(
        P2_DATAO_REG_22__SCAN_IN), .ZN(n10776) );
  AOI221_X1 U11497 ( .B1(n10777), .B2(keyinput_203), .C1(
        P2_DATAO_REG_22__SCAN_IN), .C2(keyinput_202), .A(n10776), .ZN(n10778)
         );
  OAI22_X1 U11498 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(keyinput_205), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(keyinput_206), .ZN(n10780) );
  AOI221_X1 U11499 ( .B1(P2_DATAO_REG_19__SCAN_IN), .B2(keyinput_205), .C1(
        keyinput_206), .C2(P2_DATAO_REG_18__SCAN_IN), .A(n10780), .ZN(n10783)
         );
  AOI22_X1 U11500 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(keyinput_209), .B1(
        n10785), .B2(keyinput_208), .ZN(n10784) );
  OAI221_X1 U11501 ( .B1(P2_DATAO_REG_15__SCAN_IN), .B2(keyinput_209), .C1(
        n10785), .C2(keyinput_208), .A(n10784), .ZN(n10786) );
  OAI22_X1 U11502 ( .A1(n10792), .A2(keyinput_213), .B1(keyinput_210), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n10791) );
  AOI221_X1 U11503 ( .B1(n10792), .B2(keyinput_213), .C1(
        P2_DATAO_REG_14__SCAN_IN), .C2(keyinput_210), .A(n10791), .ZN(n10794)
         );
  NOR2_X1 U11504 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(keyinput_215), .ZN(n10793) );
  XOR2_X1 U11505 ( .A(n10795), .B(keyinput_216), .Z(n10800) );
  OAI22_X1 U11506 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(keyinput_218), .B1(
        P1_IR_REG_2__SCAN_IN), .B2(keyinput_220), .ZN(n10796) );
  AOI221_X1 U11507 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(keyinput_218), .C1(
        keyinput_220), .C2(P1_IR_REG_2__SCAN_IN), .A(n10796), .ZN(n10799) );
  OAI22_X1 U11508 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(keyinput_217), .B1(
        P1_IR_REG_1__SCAN_IN), .B2(keyinput_219), .ZN(n10797) );
  AOI221_X1 U11509 ( .B1(P2_DATAO_REG_7__SCAN_IN), .B2(keyinput_217), .C1(
        keyinput_219), .C2(P1_IR_REG_1__SCAN_IN), .A(n10797), .ZN(n10798) );
  OAI211_X1 U11510 ( .C1(n10801), .C2(n10800), .A(n10799), .B(n10798), .ZN(
        n10806) );
  OAI22_X1 U11511 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(keyinput_222), .B1(
        keyinput_221), .B2(P1_IR_REG_3__SCAN_IN), .ZN(n10802) );
  AOI221_X1 U11512 ( .B1(P1_IR_REG_4__SCAN_IN), .B2(keyinput_222), .C1(
        P1_IR_REG_3__SCAN_IN), .C2(keyinput_221), .A(n10802), .ZN(n10805) );
  INV_X1 U11513 ( .A(keyinput_224), .ZN(n10808) );
  MUX2_X1 U11514 ( .A(keyinput_224), .B(n10808), .S(P1_IR_REG_6__SCAN_IN), .Z(
        n10809) );
  NAND2_X1 U11515 ( .A1(n10810), .A2(n10809), .ZN(n10813) );
  INV_X1 U11516 ( .A(keyinput_225), .ZN(n10811) );
  MUX2_X1 U11517 ( .A(n10811), .B(keyinput_225), .S(P1_IR_REG_7__SCAN_IN), .Z(
        n10812) );
  OAI22_X1 U11518 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(keyinput_226), .B1(
        keyinput_227), .B2(P1_IR_REG_9__SCAN_IN), .ZN(n10814) );
  AOI221_X1 U11519 ( .B1(P1_IR_REG_8__SCAN_IN), .B2(keyinput_226), .C1(
        P1_IR_REG_9__SCAN_IN), .C2(keyinput_227), .A(n10814), .ZN(n10820) );
  XNOR2_X1 U11520 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_230), .ZN(n10818)
         );
  XNOR2_X1 U11521 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_231), .ZN(n10817)
         );
  XNOR2_X1 U11522 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_229), .ZN(n10816)
         );
  XNOR2_X1 U11523 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_228), .ZN(n10815)
         );
  NAND4_X1 U11524 ( .A1(n10818), .A2(n10817), .A3(n10816), .A4(n10815), .ZN(
        n10819) );
  AOI22_X1 U11525 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(keyinput_233), .B1(
        P1_IR_REG_14__SCAN_IN), .B2(keyinput_232), .ZN(n10821) );
  OAI221_X1 U11526 ( .B1(P1_IR_REG_15__SCAN_IN), .B2(keyinput_233), .C1(
        P1_IR_REG_14__SCAN_IN), .C2(keyinput_232), .A(n10821), .ZN(n10822) );
  XOR2_X1 U11527 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_236), .Z(n10826) );
  INV_X1 U11528 ( .A(keyinput_234), .ZN(n10823) );
  XNOR2_X1 U11529 ( .A(n10823), .B(P1_IR_REG_16__SCAN_IN), .ZN(n10825) );
  XNOR2_X1 U11530 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_235), .ZN(n10824)
         );
  INV_X1 U11531 ( .A(keyinput_237), .ZN(n10827) );
  MUX2_X1 U11532 ( .A(n10827), .B(keyinput_237), .S(P1_IR_REG_19__SCAN_IN), 
        .Z(n10828) );
  INV_X1 U11533 ( .A(keyinput_238), .ZN(n10829) );
  MUX2_X1 U11534 ( .A(keyinput_238), .B(n10829), .S(P1_IR_REG_20__SCAN_IN), 
        .Z(n10833) );
  XNOR2_X1 U11535 ( .A(n10830), .B(keyinput_239), .ZN(n10832) );
  XNOR2_X1 U11536 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput_240), .ZN(n10831)
         );
  AOI22_X1 U11537 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(keyinput_242), .B1(
        P1_IR_REG_25__SCAN_IN), .B2(keyinput_243), .ZN(n10834) );
  OAI221_X1 U11538 ( .B1(P1_IR_REG_24__SCAN_IN), .B2(keyinput_242), .C1(
        P1_IR_REG_25__SCAN_IN), .C2(keyinput_243), .A(n10834), .ZN(n10839) );
  XNOR2_X1 U11539 ( .A(n10835), .B(keyinput_241), .ZN(n10838) );
  INV_X1 U11540 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n10836) );
  XNOR2_X1 U11541 ( .A(n10836), .B(keyinput_244), .ZN(n10837) );
  NOR4_X1 U11542 ( .A1(n10840), .A2(n10839), .A3(n10838), .A4(n10837), .ZN(
        n10856) );
  AOI22_X1 U11543 ( .A1(n10843), .A2(keyinput_250), .B1(keyinput_254), .B2(
        n10842), .ZN(n10841) );
  OAI221_X1 U11544 ( .B1(n10843), .B2(keyinput_250), .C1(n10842), .C2(
        keyinput_254), .A(n10841), .ZN(n10849) );
  XOR2_X1 U11545 ( .A(P1_D_REG_3__SCAN_IN), .B(keyinput_253), .Z(n10847) );
  XNOR2_X1 U11546 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_249), .ZN(n10846)
         );
  XNOR2_X1 U11547 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput_245), .ZN(n10845)
         );
  XNOR2_X1 U11548 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput_247), .ZN(n10844)
         );
  NAND4_X1 U11549 ( .A1(n10847), .A2(n10846), .A3(n10845), .A4(n10844), .ZN(
        n10848) );
  NOR2_X1 U11550 ( .A1(n10849), .A2(n10848), .ZN(n10854) );
  OAI22_X1 U11551 ( .A1(P1_D_REG_1__SCAN_IN), .A2(keyinput_251), .B1(
        keyinput_248), .B2(P1_IR_REG_30__SCAN_IN), .ZN(n10850) );
  AOI221_X1 U11552 ( .B1(P1_D_REG_1__SCAN_IN), .B2(keyinput_251), .C1(
        P1_IR_REG_30__SCAN_IN), .C2(keyinput_248), .A(n10850), .ZN(n10853) );
  OAI22_X1 U11553 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(keyinput_246), .B1(
        keyinput_252), .B2(P1_D_REG_2__SCAN_IN), .ZN(n10851) );
  AOI221_X1 U11554 ( .B1(P1_IR_REG_28__SCAN_IN), .B2(keyinput_246), .C1(
        P1_D_REG_2__SCAN_IN), .C2(keyinput_252), .A(n10851), .ZN(n10852) );
  NAND3_X1 U11555 ( .A1(n10854), .A2(n10853), .A3(n10852), .ZN(n10855) );
  AOI21_X1 U11556 ( .B1(keyinput_255), .B2(n10858), .A(keyinput_127), .ZN(
        n10860) );
  INV_X1 U11557 ( .A(keyinput_255), .ZN(n10857) );
  AOI21_X1 U11558 ( .B1(n10858), .B2(n10857), .A(P1_D_REG_5__SCAN_IN), .ZN(
        n10859) );
  AOI22_X1 U11559 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10860), .B1(keyinput_127), 
        .B2(n10859), .ZN(n10861) );
  AOI21_X1 U11560 ( .B1(n10863), .B2(n10862), .A(n10861), .ZN(n10879) );
  XOR2_X1 U11561 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n10864), .Z(n10876) );
  NAND2_X1 U11562 ( .A1(n10866), .A2(n10865), .ZN(n10868) );
  OAI211_X1 U11563 ( .C1(n10870), .C2(n10869), .A(n10868), .B(n10867), .ZN(
        n10875) );
  OAI21_X1 U11564 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n10873), .A(n10871), 
        .ZN(n10872) );
  AOI21_X1 U11565 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n10873), .A(n10872), 
        .ZN(n10874) );
  AOI211_X1 U11566 ( .C1(n10877), .C2(n10876), .A(n10875), .B(n10874), .ZN(
        n10878) );
  XNOR2_X1 U11567 ( .A(n10879), .B(n10878), .ZN(P1_U3258) );
  XOR2_X1 U11568 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  OAI222_X1 U11569 ( .A1(n10884), .A2(n10883), .B1(n10884), .B2(n10882), .C1(
        n10881), .C2(n10880), .ZN(ADD_1068_U5) );
  AOI21_X1 U11570 ( .B1(n10887), .B2(n10886), .A(n10885), .ZN(ADD_1068_U54) );
  AOI21_X1 U11571 ( .B1(n10890), .B2(n10889), .A(n10888), .ZN(ADD_1068_U53) );
  OAI21_X1 U11572 ( .B1(n10893), .B2(n10892), .A(n10891), .ZN(ADD_1068_U52) );
  OAI21_X1 U11573 ( .B1(n10896), .B2(n10895), .A(n10894), .ZN(ADD_1068_U51) );
  OAI21_X1 U11574 ( .B1(n10899), .B2(n10898), .A(n10897), .ZN(ADD_1068_U50) );
  OAI21_X1 U11575 ( .B1(n10902), .B2(n10901), .A(n10900), .ZN(ADD_1068_U49) );
  OAI21_X1 U11576 ( .B1(n10905), .B2(n10904), .A(n10903), .ZN(ADD_1068_U48) );
  OAI21_X1 U11577 ( .B1(n10908), .B2(n10907), .A(n10906), .ZN(ADD_1068_U47) );
  OAI21_X1 U11578 ( .B1(n10911), .B2(n10910), .A(n10909), .ZN(ADD_1068_U63) );
  OAI21_X1 U11579 ( .B1(n10914), .B2(n10913), .A(n10912), .ZN(ADD_1068_U62) );
  OAI21_X1 U11580 ( .B1(n10917), .B2(n10916), .A(n10915), .ZN(ADD_1068_U61) );
  OAI21_X1 U11581 ( .B1(n10920), .B2(n10919), .A(n10918), .ZN(ADD_1068_U60) );
  OAI21_X1 U11582 ( .B1(n10923), .B2(n10922), .A(n10921), .ZN(ADD_1068_U59) );
  OAI21_X1 U11583 ( .B1(n10926), .B2(n10925), .A(n10924), .ZN(ADD_1068_U58) );
  OAI21_X1 U11584 ( .B1(n10929), .B2(n10928), .A(n10927), .ZN(ADD_1068_U57) );
  OAI21_X1 U11585 ( .B1(n10932), .B2(n10931), .A(n10930), .ZN(ADD_1068_U56) );
  OAI21_X1 U11586 ( .B1(n10935), .B2(n10934), .A(n10933), .ZN(ADD_1068_U55) );
  NAND2_X1 U11587 ( .A1(n10997), .A2(n10936), .ZN(n10951) );
  NAND2_X1 U11588 ( .A1(n10996), .A2(P2_ADDR_REG_1__SCAN_IN), .ZN(n10950) );
  NAND2_X1 U11589 ( .A1(n10938), .A2(n10937), .ZN(n10939) );
  NAND2_X1 U11590 ( .A1(n10940), .A2(n10939), .ZN(n10942) );
  NOR2_X1 U11591 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7546), .ZN(n10941) );
  AOI21_X1 U11592 ( .B1(n10968), .B2(n10942), .A(n10941), .ZN(n10949) );
  INV_X1 U11593 ( .A(n11005), .ZN(n10962) );
  NAND2_X1 U11594 ( .A1(n10944), .A2(n10943), .ZN(n10945) );
  NAND2_X1 U11595 ( .A1(n10946), .A2(n10945), .ZN(n10947) );
  NAND2_X1 U11596 ( .A1(n10962), .A2(n10947), .ZN(n10948) );
  AND4_X1 U11597 ( .A1(n10951), .A2(n10950), .A3(n10949), .A4(n10948), .ZN(
        n10956) );
  XOR2_X1 U11598 ( .A(n10953), .B(n10952), .Z(n10954) );
  NAND2_X1 U11599 ( .A1(n10954), .A2(n11010), .ZN(n10955) );
  NAND2_X1 U11600 ( .A1(n10956), .A2(n10955), .ZN(P2_U3183) );
  OAI21_X1 U11601 ( .B1(n10959), .B2(n10958), .A(n10957), .ZN(n10961) );
  NOR2_X1 U11602 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7537), .ZN(n10960) );
  AOI21_X1 U11603 ( .B1(n10962), .B2(n10961), .A(n10960), .ZN(n10972) );
  NAND2_X1 U11604 ( .A1(n10997), .A2(n10963), .ZN(n10971) );
  NAND2_X1 U11605 ( .A1(n10996), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n10970) );
  OAI21_X1 U11606 ( .B1(n10966), .B2(n10965), .A(n10964), .ZN(n10967) );
  NAND2_X1 U11607 ( .A1(n10968), .A2(n10967), .ZN(n10969) );
  AND4_X1 U11608 ( .A1(n10972), .A2(n10971), .A3(n10970), .A4(n10969), .ZN(
        n10977) );
  XOR2_X1 U11609 ( .A(n10974), .B(n10973), .Z(n10975) );
  NAND2_X1 U11610 ( .A1(n10975), .A2(n11010), .ZN(n10976) );
  NAND2_X1 U11611 ( .A1(n10977), .A2(n10976), .ZN(P2_U3184) );
  AOI21_X1 U11612 ( .B1(n10980), .B2(n10979), .A(n10978), .ZN(n10981) );
  OAI22_X1 U11613 ( .A1(n10983), .A2(n10982), .B1(n11005), .B2(n10981), .ZN(
        n10984) );
  AOI21_X1 U11614 ( .B1(n10996), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n10984), .ZN(
        n10995) );
  OAI211_X1 U11615 ( .C1(n10987), .C2(n10986), .A(n10985), .B(n11010), .ZN(
        n10993) );
  AOI21_X1 U11616 ( .B1(n10990), .B2(n10989), .A(n10988), .ZN(n10991) );
  OR2_X1 U11617 ( .A1(n11014), .A2(n10991), .ZN(n10992) );
  NAND4_X1 U11618 ( .A1(n10995), .A2(n10994), .A3(n10993), .A4(n10992), .ZN(
        P2_U3186) );
  AOI22_X1 U11619 ( .A1(n10998), .A2(n10997), .B1(n10996), .B2(
        P2_ADDR_REG_11__SCAN_IN), .ZN(n11018) );
  AOI21_X1 U11620 ( .B1(n11001), .B2(n11000), .A(n10999), .ZN(n11015) );
  AOI21_X1 U11621 ( .B1(n11004), .B2(n11003), .A(n11002), .ZN(n11006) );
  OR2_X1 U11622 ( .A1(n11006), .A2(n11005), .ZN(n11013) );
  OAI21_X1 U11623 ( .B1(n11009), .B2(n11008), .A(n11007), .ZN(n11011) );
  NAND2_X1 U11624 ( .A1(n11011), .A2(n11010), .ZN(n11012) );
  OAI211_X1 U11625 ( .C1(n11015), .C2(n11014), .A(n11013), .B(n11012), .ZN(
        n11016) );
  INV_X1 U11626 ( .A(n11016), .ZN(n11017) );
  OAI211_X1 U11627 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n11019), .A(n11018), .B(
        n11017), .ZN(P2_U3193) );
  XOR2_X1 U11628 ( .A(n11020), .B(P1_RD_REG_SCAN_IN), .Z(U126) );
  INV_X1 U11629 ( .A(n11021), .ZN(n11027) );
  NAND2_X1 U11630 ( .A1(n11023), .A2(n11022), .ZN(n11026) );
  AOI222_X1 U11631 ( .A1(n11027), .A2(n11026), .B1(n11025), .B2(n11024), .C1(
        n6332), .C2(n11088), .ZN(n11030) );
  AOI22_X1 U11632 ( .A1(n11110), .A2(n11030), .B1(n11028), .B2(n11109), .ZN(
        P1_U3522) );
  INV_X1 U11633 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n11029) );
  AOI22_X1 U11634 ( .A1(n11114), .A2(n11030), .B1(n11029), .B2(n11111), .ZN(
        P1_U3453) );
  INV_X1 U11635 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n11031) );
  AOI22_X1 U11636 ( .A1(n11121), .A2(n11032), .B1(n11031), .B2(n6890), .ZN(
        P2_U3393) );
  INV_X1 U11637 ( .A(n11085), .ZN(n11048) );
  OAI21_X1 U11638 ( .B1(n11034), .B2(n11103), .A(n11033), .ZN(n11037) );
  INV_X1 U11639 ( .A(n11035), .ZN(n11036) );
  AOI211_X1 U11640 ( .C1(n11048), .C2(n11038), .A(n11037), .B(n11036), .ZN(
        n11040) );
  AOI22_X1 U11641 ( .A1(n11110), .A2(n11040), .B1(n7261), .B2(n11109), .ZN(
        P1_U3523) );
  INV_X1 U11642 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n11039) );
  AOI22_X1 U11643 ( .A1(n11114), .A2(n11040), .B1(n11039), .B2(n11111), .ZN(
        P1_U3456) );
  INV_X1 U11644 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n11041) );
  AOI22_X1 U11645 ( .A1(n11121), .A2(n11042), .B1(n11041), .B2(n6890), .ZN(
        P2_U3396) );
  OAI21_X1 U11646 ( .B1(n11044), .B2(n11103), .A(n11043), .ZN(n11046) );
  AOI211_X1 U11647 ( .C1(n11048), .C2(n11047), .A(n11046), .B(n11045), .ZN(
        n11050) );
  AOI22_X1 U11648 ( .A1(n11110), .A2(n11050), .B1(n7321), .B2(n11109), .ZN(
        P1_U3525) );
  INV_X1 U11649 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n11049) );
  AOI22_X1 U11650 ( .A1(n11114), .A2(n11050), .B1(n11049), .B2(n11111), .ZN(
        P1_U3462) );
  INV_X1 U11651 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n11051) );
  AOI22_X1 U11652 ( .A1(n11121), .A2(n11052), .B1(n11051), .B2(n6890), .ZN(
        P2_U3402) );
  INV_X1 U11653 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n11053) );
  AOI22_X1 U11654 ( .A1(n11121), .A2(n11054), .B1(n11053), .B2(n6890), .ZN(
        P2_U3405) );
  OAI21_X1 U11655 ( .B1(n11056), .B2(n11103), .A(n11055), .ZN(n11058) );
  AOI211_X1 U11656 ( .C1(n11107), .C2(n11059), .A(n11058), .B(n11057), .ZN(
        n11062) );
  INV_X1 U11657 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n11060) );
  AOI22_X1 U11658 ( .A1(n11110), .A2(n11062), .B1(n11060), .B2(n11109), .ZN(
        P1_U3527) );
  INV_X1 U11659 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n11061) );
  AOI22_X1 U11660 ( .A1(n11114), .A2(n11062), .B1(n11061), .B2(n11111), .ZN(
        P1_U3468) );
  INV_X1 U11661 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n11063) );
  AOI22_X1 U11662 ( .A1(n11121), .A2(n11064), .B1(n11063), .B2(n6890), .ZN(
        P2_U3408) );
  NAND2_X1 U11663 ( .A1(n11066), .A2(n11065), .ZN(n11071) );
  AOI22_X1 U11664 ( .A1(n11069), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n11068), 
        .B2(n11067), .ZN(n11070) );
  OAI211_X1 U11665 ( .C1(n11073), .C2(n11072), .A(n11071), .B(n11070), .ZN(
        n11074) );
  AOI21_X1 U11666 ( .B1(n11076), .B2(n11075), .A(n11074), .ZN(n11077) );
  OAI21_X1 U11667 ( .B1(n11079), .B2(n11078), .A(n11077), .ZN(P1_U3287) );
  INV_X1 U11668 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n11080) );
  AOI22_X1 U11669 ( .A1(n11121), .A2(n11081), .B1(n11080), .B2(n6890), .ZN(
        P2_U3420) );
  INV_X1 U11670 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n11082) );
  AOI22_X1 U11671 ( .A1(n11121), .A2(n11083), .B1(n11082), .B2(n6890), .ZN(
        P2_U3423) );
  NOR2_X1 U11672 ( .A1(n11086), .A2(n11084), .ZN(n11096) );
  NOR2_X1 U11673 ( .A1(n11086), .A2(n11085), .ZN(n11095) );
  AOI22_X1 U11674 ( .A1(n11090), .A2(n11089), .B1(n11088), .B2(n11087), .ZN(
        n11091) );
  OAI211_X1 U11675 ( .C1(n5698), .C2(n11103), .A(n11092), .B(n11091), .ZN(
        n11093) );
  NOR4_X1 U11676 ( .A1(n11096), .A2(n11095), .A3(n11094), .A4(n11093), .ZN(
        n11099) );
  INV_X1 U11677 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n11097) );
  AOI22_X1 U11678 ( .A1(n11110), .A2(n11099), .B1(n11097), .B2(n11109), .ZN(
        P1_U3533) );
  INV_X1 U11679 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n11098) );
  AOI22_X1 U11680 ( .A1(n11114), .A2(n11099), .B1(n11098), .B2(n11111), .ZN(
        P1_U3486) );
  INV_X1 U11681 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n11100) );
  AOI22_X1 U11682 ( .A1(n11121), .A2(n11101), .B1(n11100), .B2(n6890), .ZN(
        P2_U3426) );
  OAI21_X1 U11683 ( .B1(n11104), .B2(n11103), .A(n11102), .ZN(n11105) );
  AOI211_X1 U11684 ( .C1(n11108), .C2(n11107), .A(n11106), .B(n11105), .ZN(
        n11113) );
  AOI22_X1 U11685 ( .A1(n11110), .A2(n11113), .B1(n8419), .B2(n11109), .ZN(
        P1_U3534) );
  INV_X1 U11686 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n11112) );
  AOI22_X1 U11687 ( .A1(n11114), .A2(n11113), .B1(n11112), .B2(n11111), .ZN(
        P1_U3489) );
  INV_X1 U11688 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n11115) );
  AOI22_X1 U11689 ( .A1(n11121), .A2(n11116), .B1(n11115), .B2(n6890), .ZN(
        P2_U3429) );
  INV_X1 U11690 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n11117) );
  AOI22_X1 U11691 ( .A1(n11121), .A2(n11118), .B1(n11117), .B2(n6890), .ZN(
        P2_U3432) );
  INV_X1 U11692 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n11119) );
  AOI22_X1 U11693 ( .A1(n11121), .A2(n11120), .B1(n11119), .B2(n6890), .ZN(
        P2_U3435) );
  XNOR2_X1 U11694 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  AND4_X1 U5191 ( .A1(n6445), .A2(n5554), .A3(n5259), .A4(n6560), .ZN(n11124)
         );
  CLKBUF_X3 U5296 ( .A(n6493), .Z(n8841) );
endmodule

