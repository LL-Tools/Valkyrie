

module b14_C_AntiSAT_k_128_7 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3352, 
        U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343, U3342, 
        U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333, U3332, 
        U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323, U3322, 
        U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315, U3314, 
        U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305, U3304, 
        U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295, U3294, 
        U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477, U3479, 
        U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497, U3499, 
        U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511, U3512, 
        U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521, U3522, 
        U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531, U3532, 
        U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541, U3542, 
        U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289, U3288, 
        U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279, U3278, 
        U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269, U3268, 
        U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260, U3259, 
        U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250, U3249, 
        U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240, U3550, 
        U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559, U3560, 
        U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569, U3570, 
        U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579, U3580, 
        U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232, U3231, 
        U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222, U3221, 
        U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212, U3211, 
        U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2041, n2042, n2043, n2044, n2045, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735;

  AOI21_X1 U2283 ( .B1(n4282), .B2(n4715), .A(n2202), .ZN(n2201) );
  CLKBUF_X2 U2285 ( .A(n2814), .Z(n2042) );
  OAI22_X1 U2286 ( .A1(n4447), .A2(n3255), .B1(n3254), .B2(n3253), .ZN(n4457)
         );
  CLKBUF_X2 U2287 ( .A(n2401), .Z(n2853) );
  CLKBUF_X2 U2288 ( .A(n2390), .Z(n2043) );
  INV_X1 U2289 ( .A(n4622), .ZN(n4612) );
  AND2_X1 U2290 ( .A1(n2376), .A2(n2114), .ZN(n4622) );
  XNOR2_X1 U2291 ( .A(n2196), .B(IR_REG_30__SCAN_IN), .ZN(n4389) );
  OAI21_X1 U2292 ( .B1(n3724), .B2(n2163), .A(n2160), .ZN(n2159) );
  NAND2_X1 U2293 ( .A1(n2084), .A2(n3818), .ZN(n3452) );
  INV_X1 U2294 ( .A(n2814), .ZN(n2788) );
  INV_X1 U2295 ( .A(n2401), .ZN(n2048) );
  XNOR2_X1 U2296 ( .A(n3252), .B(n4444), .ZN(n4447) );
  NOR2_X1 U2297 ( .A1(n4280), .A2(n4337), .ZN(n2202) );
  OAI21_X1 U2298 ( .B1(n2348), .B2(n3241), .A(n2347), .ZN(n2350) );
  INV_X1 U2299 ( .A(n4389), .ZN(n2092) );
  NAND2_X2 U2300 ( .A1(n2350), .A2(n2349), .ZN(n3787) );
  AND2_X1 U2301 ( .A1(n4605), .A2(n3051), .ZN(n3447) );
  NAND2_X1 U2302 ( .A1(n2547), .A2(n2295), .ZN(n2549) );
  NAND2_X1 U2303 ( .A1(n3194), .A2(IR_REG_31__SCAN_IN), .ZN(n2196) );
  NAND2_X1 U2304 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2395)
         );
  NAND2_X1 U2305 ( .A1(n2350), .A2(n2349), .ZN(n2041) );
  AOI211_X2 U2306 ( .C1(n4581), .C2(n4036), .A(n4035), .B(n4034), .ZN(n4284)
         );
  NAND2_X1 U2307 ( .A1(n3092), .A2(n2852), .ZN(n2814) );
  OAI22_X2 U2308 ( .A1(n4480), .A2(n2289), .B1(REG1_REG_7__SCAN_IN), .B2(n4478), .ZN(n3258) );
  XNOR2_X2 U2309 ( .A(n2108), .B(n2414), .ZN(n3971) );
  AND2_X1 U2310 ( .A1(n2148), .A2(n2067), .ZN(n3609) );
  OR2_X1 U2311 ( .A1(n3137), .A2(n4720), .ZN(n2099) );
  NAND2_X1 U2312 ( .A1(n4212), .A2(n4211), .ZN(n4210) );
  AOI22_X1 U2313 ( .A1(n3581), .A2(n3572), .B1(n4418), .B2(n4224), .ZN(n4228)
         );
  NAND2_X1 U2314 ( .A1(n2278), .A2(n2275), .ZN(n3581) );
  NAND2_X1 U2315 ( .A1(n2198), .A2(n3884), .ZN(n3503) );
  OR2_X1 U2316 ( .A1(n2493), .A2(n3345), .ZN(n3329) );
  AOI21_X1 U2317 ( .B1(n2251), .B2(n2252), .A(n2071), .ZN(n2250) );
  AND2_X2 U2318 ( .A1(n2857), .A2(n4255), .ZN(n3762) );
  NAND2_X1 U2319 ( .A1(n2178), .A2(n2177), .ZN(n3395) );
  NAND2_X2 U2320 ( .A1(n3312), .A2(n4255), .ZN(n3379) );
  INV_X2 U2321 ( .A(n2401), .ZN(n2047) );
  AND2_X2 U2322 ( .A1(n2816), .A2(n4701), .ZN(n2472) );
  INV_X4 U2323 ( .A(n2397), .ZN(n2816) );
  CLKBUF_X1 U2324 ( .A(n3095), .Z(n4607) );
  AND2_X1 U2325 ( .A1(n3050), .A2(n4612), .ZN(n4606) );
  NAND2_X1 U2326 ( .A1(n2231), .A2(n2230), .ZN(n3854) );
  INV_X1 U2327 ( .A(n3948), .ZN(n3859) );
  NAND2_X1 U2328 ( .A1(n4470), .A2(REG1_REG_6__SCAN_IN), .ZN(n4469) );
  NOR2_X1 U2329 ( .A1(n3050), .A2(n4622), .ZN(n4600) );
  XNOR2_X1 U2330 ( .A(n3256), .B(n4659), .ZN(n4470) );
  AND3_X1 U2331 ( .A1(n2393), .A2(n2392), .A3(n2093), .ZN(n2394) );
  OR2_X1 U2332 ( .A1(n2336), .A2(n2335), .ZN(n2339) );
  CLKBUF_X2 U2333 ( .A(n2389), .Z(n2780) );
  NAND2_X1 U2334 ( .A1(n2331), .A2(IR_REG_31__SCAN_IN), .ZN(n2835) );
  NAND2_X4 U2335 ( .A1(n2092), .A2(n4390), .ZN(n3786) );
  INV_X1 U2336 ( .A(n2310), .ZN(n4390) );
  NAND2_X1 U2337 ( .A1(n2325), .A2(n2340), .ZN(n2331) );
  XNOR2_X1 U2338 ( .A(n2358), .B(IR_REG_22__SCAN_IN), .ZN(n4394) );
  NAND2_X1 U2339 ( .A1(n2175), .A2(n2174), .ZN(n2691) );
  XNOR2_X1 U2340 ( .A(n2307), .B(n2306), .ZN(n2310) );
  XNOR2_X1 U2341 ( .A(n2323), .B(IR_REG_21__SCAN_IN), .ZN(n4395) );
  OR2_X1 U2342 ( .A1(n2305), .A2(n3193), .ZN(n2307) );
  OR2_X1 U2343 ( .A1(n2346), .A2(n3193), .ZN(n3241) );
  INV_X1 U2344 ( .A(n2634), .ZN(n2175) );
  NOR2_X2 U2345 ( .A1(n2342), .A2(n2124), .ZN(n2346) );
  XNOR2_X1 U2346 ( .A(n3250), .B(n2180), .ZN(n4403) );
  NAND2_X1 U2347 ( .A1(n2097), .A2(n2273), .ZN(n2342) );
  AND2_X1 U2348 ( .A1(n2097), .A2(n2274), .ZN(n2632) );
  NOR2_X1 U2349 ( .A1(n2328), .A2(IR_REG_26__SCAN_IN), .ZN(n2228) );
  NOR2_X1 U2350 ( .A1(n2292), .A2(IR_REG_5__SCAN_IN), .ZN(n2259) );
  NOR2_X1 U2351 ( .A1(n2298), .A2(IR_REG_10__SCAN_IN), .ZN(n2274) );
  AND4_X1 U2352 ( .A1(n2316), .A2(n2301), .A3(n2300), .A4(n2299), .ZN(n2302)
         );
  AND3_X1 U2353 ( .A1(n2293), .A2(n2507), .A3(n2509), .ZN(n2294) );
  INV_X1 U2354 ( .A(IR_REG_28__SCAN_IN), .ZN(n2348) );
  NOR2_X1 U2355 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2316)
         );
  INV_X1 U2356 ( .A(IR_REG_3__SCAN_IN), .ZN(n2433) );
  INV_X1 U2357 ( .A(IR_REG_6__SCAN_IN), .ZN(n2507) );
  INV_X1 U2358 ( .A(IR_REG_7__SCAN_IN), .ZN(n2509) );
  INV_X1 U2359 ( .A(IR_REG_2__SCAN_IN), .ZN(n2414) );
  INV_X1 U2360 ( .A(IR_REG_11__SCAN_IN), .ZN(n2585) );
  NAND2_X1 U2361 ( .A1(n2265), .A2(n2262), .ZN(n3421) );
  OR2_X1 U2362 ( .A1(n3786), .A2(n4723), .ZN(n2382) );
  OAI21_X1 U2363 ( .B1(n3667), .B2(n2142), .A(n2139), .ZN(n2873) );
  AOI21_X2 U2364 ( .B1(n4183), .B2(n3078), .A(n2288), .ZN(n4158) );
  NAND2_X2 U2365 ( .A1(n2360), .A2(n4395), .ZN(n3092) );
  XNOR2_X2 U2366 ( .A(n2322), .B(n2321), .ZN(n2360) );
  AND2_X1 U2367 ( .A1(n2816), .A2(n4701), .ZN(n2044) );
  AND2_X1 U2368 ( .A1(n2816), .A2(n4701), .ZN(n2045) );
  NOR2_X1 U2370 ( .A1(n4490), .A2(n2524), .ZN(n4489) );
  AOI21_X1 U2371 ( .B1(n2168), .B2(n2166), .A(n2165), .ZN(n2164) );
  INV_X1 U2372 ( .A(n3651), .ZN(n2165) );
  INV_X1 U2373 ( .A(n2172), .ZN(n2166) );
  AND2_X1 U2374 ( .A1(n3395), .A2(n3394), .ZN(n3397) );
  AND2_X1 U2375 ( .A1(n3906), .A2(n2224), .ZN(n2223) );
  NAND2_X1 U2376 ( .A1(n2225), .A2(n3572), .ZN(n2224) );
  AND2_X1 U2377 ( .A1(n4052), .A2(n4603), .ZN(n2102) );
  OR2_X1 U2378 ( .A1(n4249), .A2(n4248), .ZN(n4246) );
  OR2_X1 U2379 ( .A1(IR_REG_25__SCAN_IN), .A2(n2326), .ZN(n2328) );
  INV_X1 U2380 ( .A(IR_REG_23__SCAN_IN), .ZN(n2112) );
  INV_X1 U2381 ( .A(IR_REG_21__SCAN_IN), .ZN(n2341) );
  INV_X1 U2382 ( .A(IR_REG_9__SCAN_IN), .ZN(n2295) );
  OR2_X1 U2383 ( .A1(n2778), .A2(n3746), .ZN(n2793) );
  INV_X1 U2384 ( .A(n2780), .ZN(n2811) );
  NAND2_X1 U2385 ( .A1(n4460), .A2(n4461), .ZN(n4459) );
  OR2_X1 U2386 ( .A1(n4489), .A2(n3260), .ZN(n2178) );
  INV_X1 U2387 ( .A(IR_REG_13__SCAN_IN), .ZN(n2315) );
  AND2_X1 U2388 ( .A1(n2804), .A2(REG3_REG_28__SCAN_IN), .ZN(n3594) );
  OR2_X1 U2389 ( .A1(n4037), .A2(n3584), .ZN(n3588) );
  AND2_X1 U2390 ( .A1(n4090), .A2(n4072), .ZN(n4074) );
  NAND2_X1 U2391 ( .A1(n2360), .A2(n2836), .ZN(n4701) );
  XNOR2_X1 U2392 ( .A(n3987), .B(n2110), .ZN(n4557) );
  INV_X1 U2393 ( .A(n4645), .ZN(n2110) );
  OAI21_X1 U2394 ( .B1(n2164), .B2(n2162), .A(n2072), .ZN(n2161) );
  INV_X1 U2395 ( .A(n2648), .ZN(n2162) );
  INV_X1 U2396 ( .A(n3781), .ZN(n2214) );
  AND2_X1 U2397 ( .A1(n3608), .A2(n2067), .ZN(n2147) );
  OR2_X1 U2398 ( .A1(n3721), .A2(n3722), .ZN(n2172) );
  INV_X1 U2399 ( .A(n2130), .ZN(n2129) );
  INV_X1 U2400 ( .A(n2171), .ZN(n2169) );
  NAND2_X1 U2401 ( .A1(n2345), .A2(n3163), .ZN(n2401) );
  NOR2_X1 U2402 ( .A1(n2682), .A2(n3675), .ZN(n2135) );
  INV_X1 U2403 ( .A(n2213), .ZN(n2212) );
  OAI21_X1 U2404 ( .B1(n2215), .B2(n2214), .A(n3794), .ZN(n2213) );
  AOI21_X1 U2405 ( .B1(n2212), .B2(n2214), .A(n2211), .ZN(n2210) );
  INV_X1 U2406 ( .A(n3782), .ZN(n2211) );
  NAND2_X1 U2407 ( .A1(n2212), .A2(n3916), .ZN(n2208) );
  NOR2_X1 U2408 ( .A1(n3772), .A2(n2068), .ZN(n2225) );
  INV_X1 U2409 ( .A(n3769), .ZN(n2226) );
  NOR2_X1 U2410 ( .A1(n3074), .A2(n3534), .ZN(n2279) );
  NAND2_X1 U2411 ( .A1(n2280), .A2(n3075), .ZN(n2277) );
  AND2_X1 U2412 ( .A1(n2283), .A2(n2281), .ZN(n2280) );
  OAI21_X1 U2413 ( .B1(n3503), .B2(n3878), .A(n3875), .ZN(n3472) );
  AND2_X1 U2414 ( .A1(n3428), .A2(n2117), .ZN(n2116) );
  NOR2_X1 U2415 ( .A1(n2268), .A2(n2267), .ZN(n2266) );
  INV_X1 U2416 ( .A(n3813), .ZN(n2268) );
  NAND2_X1 U2417 ( .A1(n2271), .A2(n2272), .ZN(n2267) );
  INV_X1 U2418 ( .A(n3061), .ZN(n2271) );
  AOI21_X1 U2419 ( .B1(n2089), .B2(n2091), .A(n2087), .ZN(n2086) );
  INV_X1 U2420 ( .A(n3767), .ZN(n2087) );
  AOI21_X1 U2421 ( .B1(n2290), .B2(n2284), .A(n2079), .ZN(n2283) );
  NAND2_X1 U2422 ( .A1(n3072), .A2(n2284), .ZN(n2282) );
  NAND2_X1 U2423 ( .A1(n2585), .A2(n2297), .ZN(n2298) );
  INV_X1 U2424 ( .A(IR_REG_12__SCAN_IN), .ZN(n2297) );
  NAND2_X1 U2425 ( .A1(n2228), .A2(n2056), .ZN(n2124) );
  INV_X1 U2426 ( .A(IR_REG_24__SCAN_IN), .ZN(n2333) );
  NOR2_X1 U2427 ( .A1(n2145), .A2(n3665), .ZN(n2144) );
  INV_X1 U2428 ( .A(n3744), .ZN(n2145) );
  INV_X1 U2429 ( .A(n3632), .ZN(n2752) );
  INV_X1 U2430 ( .A(n2157), .ZN(n2150) );
  NAND2_X1 U2431 ( .A1(n3437), .A2(n3436), .ZN(n2173) );
  AOI21_X1 U2432 ( .B1(n2134), .B2(n2683), .A(n2131), .ZN(n2130) );
  INV_X1 U2433 ( .A(n3733), .ZN(n2131) );
  NAND2_X1 U2434 ( .A1(n3787), .A2(n2396), .ZN(n2229) );
  NOR2_X1 U2435 ( .A1(n3141), .A2(n3144), .ZN(n3155) );
  NAND2_X1 U2436 ( .A1(n3721), .A2(n3722), .ZN(n2171) );
  NAND2_X1 U2437 ( .A1(n3724), .A2(n2172), .ZN(n2170) );
  NOR2_X2 U2438 ( .A1(n3142), .A2(n3143), .ZN(n3141) );
  NOR2_X1 U2439 ( .A1(n3713), .A2(n2153), .ZN(n2152) );
  INV_X1 U2440 ( .A(n2156), .ZN(n2153) );
  NAND2_X1 U2441 ( .A1(n2138), .A2(n2137), .ZN(n2136) );
  INV_X1 U2442 ( .A(n3674), .ZN(n2138) );
  INV_X1 U2443 ( .A(n2135), .ZN(n2133) );
  OR2_X1 U2444 ( .A1(n2794), .A2(n2804), .ZN(n3610) );
  NAND4_X1 U2445 ( .A1(n2412), .A2(n2411), .A3(n2410), .A4(n2409), .ZN(n3054)
         );
  NAND2_X1 U2446 ( .A1(n2390), .A2(REG0_REG_1__SCAN_IN), .ZN(n2093) );
  NAND2_X1 U2447 ( .A1(n3976), .A2(n3229), .ZN(n3230) );
  NAND2_X1 U2448 ( .A1(n4459), .A2(n2070), .ZN(n3235) );
  NAND2_X1 U2449 ( .A1(n4456), .A2(n2053), .ZN(n3256) );
  INV_X1 U2450 ( .A(n3263), .ZN(n2177) );
  XNOR2_X1 U2451 ( .A(n3397), .B(n4654), .ZN(n4498) );
  NOR2_X1 U2452 ( .A1(n4498), .A2(n2562), .ZN(n4497) );
  NAND2_X1 U2453 ( .A1(n2182), .A2(n2181), .ZN(n3994) );
  INV_X1 U2454 ( .A(n3401), .ZN(n2181) );
  NAND2_X1 U2455 ( .A1(n3982), .A2(n2106), .ZN(n3983) );
  NAND2_X1 U2456 ( .A1(n2107), .A2(REG2_REG_11__SCAN_IN), .ZN(n2106) );
  INV_X1 U2457 ( .A(n4391), .ZN(n3225) );
  INV_X1 U2458 ( .A(n3587), .ZN(n3791) );
  NOR2_X1 U2459 ( .A1(n2793), .A2(n3611), .ZN(n2804) );
  OR2_X1 U2460 ( .A1(n2253), .A2(n2062), .ZN(n2251) );
  AND2_X1 U2461 ( .A1(n2065), .A2(n3084), .ZN(n2253) );
  OR2_X1 U2462 ( .A1(n3085), .A2(n2062), .ZN(n2252) );
  INV_X1 U2463 ( .A(n4110), .ZN(n4067) );
  AND2_X1 U2464 ( .A1(n4105), .A2(n4104), .ZN(n4125) );
  NAND2_X1 U2465 ( .A1(n2075), .A2(n2049), .ZN(n2242) );
  AOI21_X1 U2466 ( .B1(n2242), .B2(n2244), .A(n2240), .ZN(n2239) );
  INV_X1 U2467 ( .A(n4124), .ZN(n2240) );
  INV_X1 U2468 ( .A(n2242), .ZN(n2241) );
  NAND2_X1 U2469 ( .A1(n4210), .A2(n3077), .ZN(n4183) );
  NAND2_X1 U2470 ( .A1(n4213), .A2(n3076), .ZN(n3077) );
  AOI21_X1 U2471 ( .B1(n2257), .B2(n2256), .A(n2255), .ZN(n4212) );
  AND2_X1 U2472 ( .A1(n3939), .A2(n4229), .ZN(n2255) );
  NAND2_X1 U2473 ( .A1(n4412), .A2(n4222), .ZN(n2256) );
  INV_X1 U2474 ( .A(n4228), .ZN(n2257) );
  AND2_X1 U2475 ( .A1(n2282), .A2(n2280), .ZN(n4240) );
  AND2_X1 U2476 ( .A1(n2116), .A2(n3476), .ZN(n2115) );
  NAND2_X1 U2477 ( .A1(n2098), .A2(n3867), .ZN(n3370) );
  NAND2_X1 U2478 ( .A1(n3357), .A2(n3883), .ZN(n2098) );
  INV_X1 U2479 ( .A(n2267), .ZN(n2264) );
  NAND2_X1 U2480 ( .A1(n3059), .A2(n2272), .ZN(n2261) );
  OR2_X1 U2481 ( .A1(n3946), .A2(n3488), .ZN(n2272) );
  OAI21_X1 U2482 ( .B1(n3487), .B2(n3486), .A(n3881), .ZN(n3357) );
  NAND2_X1 U2483 ( .A1(n3093), .A2(n2707), .ZN(n4608) );
  INV_X1 U2484 ( .A(n4585), .ZN(n4624) );
  NOR2_X1 U2485 ( .A1(n3118), .A2(n2101), .ZN(n3602) );
  OR2_X1 U2486 ( .A1(n3119), .A2(n2102), .ZN(n2101) );
  AND2_X1 U2487 ( .A1(n4175), .A2(n2081), .ZN(n4090) );
  AND2_X1 U2488 ( .A1(n4194), .A2(n4177), .ZN(n4175) );
  INV_X1 U2489 ( .A(IR_REG_29__SCAN_IN), .ZN(n2306) );
  NOR2_X1 U2490 ( .A1(n2303), .A2(IR_REG_22__SCAN_IN), .ZN(n2227) );
  OR2_X1 U2491 ( .A1(IR_REG_27__SCAN_IN), .A2(IR_REG_28__SCAN_IN), .ZN(n2303)
         );
  INV_X1 U2492 ( .A(IR_REG_27__SCAN_IN), .ZN(n2861) );
  NAND2_X1 U2493 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_26__SCAN_IN), .ZN(n2335) );
  INV_X1 U2494 ( .A(IR_REG_26__SCAN_IN), .ZN(n2337) );
  NAND2_X1 U2495 ( .A1(n2112), .A2(n2333), .ZN(n2326) );
  NAND2_X1 U2496 ( .A1(n2175), .A2(n2318), .ZN(n2673) );
  INV_X1 U2497 ( .A(IR_REG_8__SCAN_IN), .ZN(n2293) );
  INV_X1 U2498 ( .A(n2432), .ZN(n2176) );
  NAND2_X1 U2499 ( .A1(n2109), .A2(IR_REG_31__SCAN_IN), .ZN(n2108) );
  INV_X1 U2500 ( .A(n2413), .ZN(n2109) );
  INV_X1 U2501 ( .A(IR_REG_1__SCAN_IN), .ZN(n2183) );
  OAI21_X1 U2502 ( .B1(n3686), .B2(n3690), .A(n3688), .ZN(n3667) );
  AND2_X1 U2503 ( .A1(n2854), .A2(n3285), .ZN(n4429) );
  NAND2_X1 U2504 ( .A1(n2785), .A2(n2784), .ZN(n4069) );
  INV_X1 U2505 ( .A(n4660), .ZN(n4464) );
  XNOR2_X1 U2506 ( .A(n3235), .B(n4659), .ZN(n4472) );
  XNOR2_X1 U2507 ( .A(n3983), .B(n2105), .ZN(n4512) );
  NAND2_X1 U2508 ( .A1(n4512), .A2(REG2_REG_12__SCAN_IN), .ZN(n4511) );
  NAND2_X1 U2509 ( .A1(n4556), .A2(n3988), .ZN(n4568) );
  AOI21_X1 U2510 ( .B1(n4008), .B2(n4007), .A(n4540), .ZN(n4011) );
  AND2_X1 U2511 ( .A1(n4440), .A2(n3931), .ZN(n4571) );
  NAND2_X1 U2512 ( .A1(n2197), .A2(n3853), .ZN(n4665) );
  INV_X1 U2513 ( .A(n4600), .ZN(n2197) );
  NAND2_X1 U2514 ( .A1(n3602), .A2(n2100), .ZN(n3137) );
  OR2_X1 U2515 ( .A1(n3607), .A2(n4337), .ZN(n2100) );
  NAND2_X1 U2516 ( .A1(n2203), .A2(n2201), .ZN(n4351) );
  INV_X1 U2517 ( .A(n4281), .ZN(n2203) );
  AND2_X1 U2518 ( .A1(n2216), .A2(n3115), .ZN(n2215) );
  INV_X1 U2519 ( .A(n4031), .ZN(n2216) );
  OAI21_X1 U2520 ( .B1(n2223), .B2(n2222), .A(n2221), .ZN(n2220) );
  INV_X1 U2521 ( .A(n3908), .ZN(n2221) );
  NAND2_X1 U2522 ( .A1(n2218), .A2(n2215), .ZN(n2217) );
  AOI21_X1 U2523 ( .B1(n3850), .B2(n2090), .A(n2281), .ZN(n2089) );
  INV_X1 U2524 ( .A(n3850), .ZN(n2091) );
  NAND2_X1 U2525 ( .A1(n2729), .A2(n2158), .ZN(n2157) );
  INV_X1 U2526 ( .A(n2159), .ZN(n2663) );
  NAND2_X1 U2527 ( .A1(n2168), .A2(n2648), .ZN(n2163) );
  INV_X1 U2528 ( .A(n2161), .ZN(n2160) );
  OR2_X1 U2529 ( .A1(n3786), .A2(n3245), .ZN(n2411) );
  AND2_X1 U2530 ( .A1(n3994), .A2(n3993), .ZN(n3995) );
  AOI21_X1 U2531 ( .B1(n3999), .B2(REG1_REG_13__SCAN_IN), .A(n4515), .ZN(n4000) );
  AND2_X1 U2532 ( .A1(n4184), .A2(n3828), .ZN(n4164) );
  NAND2_X1 U2533 ( .A1(n3053), .A2(n3052), .ZN(n3855) );
  INV_X1 U2534 ( .A(n3094), .ZN(n3209) );
  XNOR2_X1 U2535 ( .A(n2103), .B(n3807), .ZN(n3117) );
  NAND2_X1 U2536 ( .A1(n2217), .A2(n3781), .ZN(n2103) );
  INV_X1 U2537 ( .A(n2217), .ZN(n4030) );
  NOR2_X1 U2538 ( .A1(n4136), .A2(n3081), .ZN(n2120) );
  NAND2_X1 U2539 ( .A1(n4175), .A2(n4151), .ZN(n4150) );
  AND2_X1 U2540 ( .A1(n2856), .A2(n3123), .ZN(n2836) );
  NOR2_X2 U2541 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2413)
         );
  INV_X1 U2542 ( .A(n2144), .ZN(n2142) );
  AND2_X1 U2543 ( .A1(n2147), .A2(n2140), .ZN(n2139) );
  NAND2_X1 U2544 ( .A1(n2144), .A2(n2141), .ZN(n2140) );
  INV_X1 U2545 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2594) );
  INV_X1 U2546 ( .A(n4069), .ZN(n4029) );
  NOR2_X1 U2547 ( .A1(n2701), .A2(n2700), .ZN(n2715) );
  AND2_X1 U2548 ( .A1(n2715), .A2(REG3_REG_20__SCAN_IN), .ZN(n2717) );
  AND2_X1 U2549 ( .A1(n2128), .A2(n3642), .ZN(n2127) );
  NAND2_X1 U2550 ( .A1(n2130), .A2(n2132), .ZN(n2128) );
  OAI21_X1 U2551 ( .B1(n3724), .B2(n2167), .A(n2164), .ZN(n3701) );
  NOR2_X1 U2552 ( .A1(n2595), .A2(n2594), .ZN(n2625) );
  NAND2_X1 U2553 ( .A1(n3153), .A2(n2728), .ZN(n2156) );
  NAND2_X1 U2554 ( .A1(n3155), .A2(n2157), .ZN(n2154) );
  OR2_X1 U2555 ( .A1(n2731), .A2(n3714), .ZN(n2739) );
  XNOR2_X1 U2556 ( .A(n2400), .B(n2814), .ZN(n2403) );
  NAND2_X1 U2557 ( .A1(n2399), .A2(n2398), .ZN(n2400) );
  AOI21_X1 U2558 ( .B1(n3049), .B2(n2044), .A(n2402), .ZN(n2404) );
  NAND2_X1 U2559 ( .A1(n2667), .A2(REG3_REG_17__SCAN_IN), .ZN(n2685) );
  OR2_X1 U2560 ( .A1(n2685), .A2(n2684), .ZN(n2701) );
  OR3_X1 U2561 ( .A1(n2853), .A2(n2852), .A3(n3204), .ZN(n2859) );
  NAND2_X1 U2562 ( .A1(n4402), .A2(n3251), .ZN(n3252) );
  OAI22_X1 U2563 ( .A1(n4445), .A2(n3234), .B1(n3233), .B2(n3253), .ZN(n4460)
         );
  XNOR2_X1 U2564 ( .A(n3258), .B(n2179), .ZN(n4490) );
  NAND2_X1 U2565 ( .A1(n4484), .A2(n2104), .ZN(n3237) );
  NAND2_X1 U2566 ( .A1(n4478), .A2(REG2_REG_7__SCAN_IN), .ZN(n2104) );
  OR2_X1 U2567 ( .A1(n4497), .A2(n3398), .ZN(n2182) );
  XNOR2_X1 U2568 ( .A(n4000), .B(n4649), .ZN(n4528) );
  OAI21_X1 U2569 ( .B1(n4528), .B2(n2185), .A(n2184), .ZN(n4541) );
  NAND2_X1 U2570 ( .A1(n2186), .A2(REG1_REG_14__SCAN_IN), .ZN(n2185) );
  NAND2_X1 U2571 ( .A1(n4001), .A2(n2186), .ZN(n2184) );
  INV_X1 U2572 ( .A(n4542), .ZN(n2186) );
  NOR2_X1 U2573 ( .A1(n4528), .A2(n4529), .ZN(n4527) );
  NOR2_X1 U2574 ( .A1(n4545), .A2(n2111), .ZN(n3987) );
  AND2_X1 U2575 ( .A1(n4646), .A2(REG2_REG_15__SCAN_IN), .ZN(n2111) );
  AND2_X1 U2576 ( .A1(n2318), .A2(n2319), .ZN(n2174) );
  INV_X1 U2577 ( .A(IR_REG_17__SCAN_IN), .ZN(n2319) );
  NAND2_X1 U2578 ( .A1(n4643), .A2(n4326), .ZN(n2195) );
  NOR2_X1 U2579 ( .A1(n2193), .A2(n4007), .ZN(n2192) );
  INV_X1 U2580 ( .A(n2195), .ZN(n2193) );
  NOR3_X1 U2581 ( .A1(n4037), .A2(n3584), .A3(n3791), .ZN(n4271) );
  AND2_X1 U2582 ( .A1(n2210), .A2(n2208), .ZN(n2207) );
  AOI21_X1 U2583 ( .B1(n2239), .B2(n2241), .A(n2074), .ZN(n2236) );
  NAND2_X1 U2584 ( .A1(n2219), .A2(n2223), .ZN(n4103) );
  NAND2_X1 U2585 ( .A1(n4246), .A2(n2225), .ZN(n2219) );
  OR2_X1 U2586 ( .A1(n4160), .A2(n4159), .ZN(n4221) );
  NOR2_X1 U2587 ( .A1(n2649), .A2(n3760), .ZN(n2651) );
  NAND2_X1 U2588 ( .A1(n2277), .A2(n2276), .ZN(n2275) );
  INV_X1 U2589 ( .A(n3074), .ZN(n2276) );
  NAND2_X1 U2590 ( .A1(n4246), .A2(n3769), .ZN(n3571) );
  AND2_X1 U2591 ( .A1(n3571), .A2(n3819), .ZN(n4160) );
  NOR2_X1 U2592 ( .A1(n4340), .A2(n4254), .ZN(n4253) );
  NOR2_X1 U2593 ( .A1(n3545), .A2(n3544), .ZN(n2119) );
  NAND2_X1 U2594 ( .A1(n2088), .A2(n3850), .ZN(n3771) );
  NAND2_X1 U2595 ( .A1(n3537), .A2(n3847), .ZN(n2088) );
  OR2_X1 U2596 ( .A1(n2560), .A2(n2559), .ZN(n2578) );
  INV_X1 U2597 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3393) );
  NAND2_X1 U2598 ( .A1(n3427), .A2(n3874), .ZN(n2198) );
  NAND2_X1 U2599 ( .A1(n3422), .A2(n2116), .ZN(n3512) );
  AOI21_X1 U2600 ( .B1(n2260), .B2(n3813), .A(n2052), .ZN(n2262) );
  AND3_X1 U2601 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2474) );
  NAND2_X1 U2602 ( .A1(n2474), .A2(REG3_REG_6__SCAN_IN), .ZN(n2520) );
  OAI21_X1 U2603 ( .B1(n3302), .B2(n3097), .A(n3865), .ZN(n3487) );
  NAND2_X1 U2604 ( .A1(n3410), .A2(n3861), .ZN(n3302) );
  NAND2_X1 U2605 ( .A1(n3446), .A2(n3055), .ZN(n3406) );
  AND2_X1 U2606 ( .A1(n3804), .A2(n3116), .ZN(n4585) );
  NAND2_X1 U2607 ( .A1(n3855), .A2(n3857), .ZN(n3450) );
  NOR2_X1 U2608 ( .A1(n3207), .A2(n3120), .ZN(n3310) );
  NAND2_X1 U2609 ( .A1(n4622), .A2(n3128), .ZN(n4614) );
  NOR2_X1 U2610 ( .A1(n2122), .A2(n3089), .ZN(n2121) );
  NAND2_X1 U2611 ( .A1(n3131), .A2(n2123), .ZN(n2122) );
  NOR2_X1 U2612 ( .A1(n4277), .A2(n3791), .ZN(n2123) );
  AND2_X1 U2613 ( .A1(n4396), .A2(n2836), .ZN(n4602) );
  AND2_X1 U2614 ( .A1(n4074), .A2(n4058), .ZN(n4056) );
  NAND2_X1 U2615 ( .A1(n4175), .A2(n2051), .ZN(n4114) );
  NAND2_X1 U2616 ( .A1(n4175), .A2(n2120), .ZN(n4304) );
  NOR2_X1 U2617 ( .A1(n4232), .A2(n3130), .ZN(n4194) );
  NAND2_X1 U2618 ( .A1(n4253), .A2(n3576), .ZN(n4230) );
  OR2_X1 U2619 ( .A1(n4230), .A2(n4229), .ZN(n4232) );
  AND2_X1 U2620 ( .A1(n4608), .A2(n4679), .ZN(n4337) );
  NAND2_X1 U2621 ( .A1(n2282), .A2(n2283), .ZN(n3552) );
  INV_X1 U2622 ( .A(n2119), .ZN(n3557) );
  AND2_X1 U2623 ( .A1(n3422), .A2(n2077), .ZN(n4589) );
  NAND2_X1 U2624 ( .A1(n4589), .A2(n3658), .ZN(n3545) );
  AND2_X1 U2625 ( .A1(n3377), .A2(n3869), .ZN(n3422) );
  NAND2_X1 U2626 ( .A1(n3422), .A2(n3428), .ZN(n3510) );
  OR2_X1 U2627 ( .A1(n3494), .A2(n3488), .ZN(n3495) );
  NOR2_X1 U2628 ( .A1(n3495), .A2(n3364), .ZN(n3377) );
  NAND2_X1 U2629 ( .A1(n2113), .A2(n3455), .ZN(n4674) );
  INV_X1 U2630 ( .A(n4614), .ZN(n2113) );
  INV_X1 U2631 ( .A(n4701), .ZN(n4715) );
  INV_X1 U2632 ( .A(IR_REG_20__SCAN_IN), .ZN(n2321) );
  NAND2_X1 U2633 ( .A1(n2355), .A2(IR_REG_31__SCAN_IN), .ZN(n2322) );
  NAND2_X1 U2634 ( .A1(n2146), .A2(n2144), .ZN(n2148) );
  INV_X1 U2635 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3635) );
  INV_X1 U2636 ( .A(n2152), .ZN(n2151) );
  NOR2_X1 U2637 ( .A1(n2753), .A2(n2069), .ZN(n2149) );
  NAND2_X1 U2638 ( .A1(n2752), .A2(n2751), .ZN(n2753) );
  NAND2_X1 U2639 ( .A1(n2173), .A2(n2558), .ZN(n3186) );
  NAND2_X1 U2640 ( .A1(n2126), .A2(n2130), .ZN(n3643) );
  NAND2_X1 U2641 ( .A1(n3674), .A2(n2134), .ZN(n2126) );
  INV_X1 U2642 ( .A(n3100), .ZN(n3428) );
  XNOR2_X1 U2643 ( .A(n2403), .B(n2404), .ZN(n2125) );
  NAND2_X1 U2644 ( .A1(n2170), .A2(n2171), .ZN(n3654) );
  INV_X1 U2645 ( .A(n4205), .ZN(n3738) );
  AND2_X1 U2646 ( .A1(n2154), .A2(n2152), .ZN(n3711) );
  NAND2_X1 U2647 ( .A1(n2154), .A2(n2156), .ZN(n3712) );
  NAND2_X1 U2648 ( .A1(n2136), .A2(n2133), .ZN(n3736) );
  INV_X1 U2649 ( .A(n3665), .ZN(n2143) );
  AND2_X1 U2650 ( .A1(n2793), .A2(n2779), .ZN(n4059) );
  OAI21_X1 U2651 ( .B1(n3610), .B2(n2811), .A(n2799), .ZN(n4052) );
  OAI211_X1 U2652 ( .C1(n3668), .C2(n2811), .A(n2772), .B(n2771), .ZN(n4086)
         );
  OAI211_X1 U2653 ( .C1(n4094), .C2(n2811), .A(n2758), .B(n2757), .ZN(n4110)
         );
  NAND4_X1 U2654 ( .A1(n2744), .A2(n2743), .A3(n2742), .A4(n2741), .ZN(n4126)
         );
  AND2_X1 U2655 ( .A1(n3224), .A2(n3223), .ZN(n4440) );
  NAND2_X1 U2656 ( .A1(n3950), .A2(n3951), .ZN(n3965) );
  NAND2_X1 U2657 ( .A1(n3228), .A2(n3227), .ZN(n3976) );
  XNOR2_X1 U2658 ( .A(n3230), .B(n2180), .ZN(n4405) );
  NAND2_X1 U2659 ( .A1(n4405), .A2(REG2_REG_3__SCAN_IN), .ZN(n4404) );
  NAND2_X1 U2660 ( .A1(n4403), .A2(REG1_REG_3__SCAN_IN), .ZN(n4402) );
  NAND2_X1 U2661 ( .A1(n4471), .A2(n3236), .ZN(n4485) );
  NAND2_X1 U2662 ( .A1(n4485), .A2(n4486), .ZN(n4484) );
  NAND2_X1 U2663 ( .A1(n4469), .A2(n3257), .ZN(n4480) );
  XNOR2_X1 U2664 ( .A(n3237), .B(n2179), .ZN(n4494) );
  INV_X1 U2665 ( .A(n2178), .ZN(n3264) );
  INV_X1 U2666 ( .A(n2182), .ZN(n3402) );
  NAND2_X1 U2667 ( .A1(n3984), .A2(n4511), .ZN(n4523) );
  NAND2_X1 U2668 ( .A1(n4557), .A2(n3578), .ZN(n4556) );
  AND2_X1 U2669 ( .A1(n4440), .A2(n3960), .ZN(n4573) );
  INV_X1 U2670 ( .A(n4573), .ZN(n4540) );
  OAI21_X1 U2671 ( .B1(n2194), .B2(n2190), .A(n2189), .ZN(n2188) );
  NAND2_X1 U2672 ( .A1(n2194), .A2(n4015), .ZN(n2189) );
  NOR2_X1 U2673 ( .A1(n2192), .A2(n4016), .ZN(n2190) );
  NAND2_X1 U2674 ( .A1(n4017), .A2(n4015), .ZN(n2191) );
  NAND2_X1 U2675 ( .A1(n2206), .A2(n2204), .ZN(n4281) );
  NOR2_X1 U2676 ( .A1(n2061), .A2(n2205), .ZN(n2204) );
  OR2_X1 U2677 ( .A1(n3593), .A2(n4585), .ZN(n2206) );
  INV_X1 U2678 ( .A(n3592), .ZN(n2205) );
  OR2_X1 U2679 ( .A1(n3594), .A2(n2805), .ZN(n3601) );
  NAND2_X1 U2680 ( .A1(n2249), .A2(n2251), .ZN(n4045) );
  OR2_X1 U2681 ( .A1(n4080), .A2(n2252), .ZN(n2249) );
  OR2_X1 U2682 ( .A1(n4080), .A2(n3085), .ZN(n2254) );
  NAND2_X1 U2683 ( .A1(n2238), .A2(n2242), .ZN(n4123) );
  NAND2_X1 U2684 ( .A1(n4158), .A2(n2243), .ZN(n2238) );
  NAND2_X1 U2685 ( .A1(n4158), .A2(n3080), .ZN(n2245) );
  NAND2_X1 U2686 ( .A1(n2119), .A2(n3625), .ZN(n4340) );
  NAND2_X1 U2687 ( .A1(n3379), .A2(n3376), .ZN(n4262) );
  INV_X1 U2688 ( .A(n2260), .ZN(n2270) );
  NAND2_X1 U2689 ( .A1(n2269), .A2(n2272), .ZN(n3356) );
  OR2_X1 U2690 ( .A1(n3493), .A2(n3059), .ZN(n2269) );
  INV_X1 U2691 ( .A(n4262), .ZN(n4237) );
  AND2_X1 U2692 ( .A1(n3379), .A2(n3314), .ZN(n4630) );
  INV_X1 U2693 ( .A(n3049), .ZN(n3048) );
  INV_X2 U2694 ( .A(n3379), .ZN(n4634) );
  OR2_X1 U2695 ( .A1(n4074), .A2(n4073), .ZN(n4360) );
  INV_X1 U2696 ( .A(n4720), .ZN(n4722) );
  INV_X1 U2697 ( .A(n4640), .ZN(n3204) );
  AND2_X1 U2698 ( .A1(n2060), .A2(n2097), .ZN(n2095) );
  XNOR2_X1 U2699 ( .A(n2863), .B(IR_REG_28__SCAN_IN), .ZN(n4391) );
  NOR2_X1 U2700 ( .A1(n2343), .A2(n2346), .ZN(n4392) );
  NAND2_X1 U2701 ( .A1(n2339), .A2(n2338), .ZN(n2343) );
  NAND2_X1 U2702 ( .A1(n3193), .A2(n2337), .ZN(n2338) );
  OAI21_X1 U2703 ( .B1(n2331), .B2(n2326), .A(IR_REG_31__SCAN_IN), .ZN(n2327)
         );
  AND2_X1 U2704 ( .A1(n3208), .A2(STATE_REG_SCAN_IN), .ZN(n4640) );
  XNOR2_X1 U2705 ( .A(n2372), .B(n2371), .ZN(n4645) );
  NOR2_X1 U2706 ( .A1(n2550), .A2(n2097), .ZN(n4399) );
  INV_X1 U2707 ( .A(n2292), .ZN(n2258) );
  OR4_X1 U2708 ( .A1(n3162), .A2(n3161), .A3(n3160), .A4(n3159), .ZN(U3220) );
  AOI21_X1 U2709 ( .B1(n4011), .B2(n2055), .A(n4010), .ZN(n4012) );
  NAND2_X1 U2710 ( .A1(n2235), .A2(n2234), .ZN(U3547) );
  NAND2_X1 U2711 ( .A1(n4733), .A2(REG1_REG_29__SCAN_IN), .ZN(n2234) );
  NAND2_X1 U2712 ( .A1(n4351), .A2(n4735), .ZN(n2235) );
  OR2_X1 U2713 ( .A1(n3599), .A2(n4328), .ZN(n3133) );
  NAND2_X1 U2714 ( .A1(n2200), .A2(n2082), .ZN(U3515) );
  INV_X1 U2715 ( .A(REG0_REG_29__SCAN_IN), .ZN(n2199) );
  NAND2_X1 U2716 ( .A1(n2099), .A2(n2078), .ZN(n3139) );
  INV_X1 U2717 ( .A(n2728), .ZN(n2158) );
  NAND2_X2 U2718 ( .A1(n3163), .A2(n3092), .ZN(n2397) );
  AND2_X1 U2719 ( .A1(n2245), .A2(n2247), .ZN(n4148) );
  OR2_X1 U2720 ( .A1(n4171), .A2(n3081), .ZN(n2049) );
  AND2_X1 U2721 ( .A1(n2714), .A2(n2713), .ZN(n2050) );
  AND2_X1 U2722 ( .A1(n2529), .A2(n2511), .ZN(n4478) );
  AND2_X1 U2723 ( .A1(n3535), .A2(n3104), .ZN(n3847) );
  INV_X1 U2724 ( .A(n3847), .ZN(n2090) );
  INV_X1 U2725 ( .A(n2707), .ZN(n4397) );
  AND2_X1 U2726 ( .A1(n2120), .A2(n4115), .ZN(n2051) );
  INV_X1 U2727 ( .A(n3992), .ZN(n2107) );
  AND2_X1 U2728 ( .A1(n4389), .A2(n4390), .ZN(n2389) );
  INV_X2 U2729 ( .A(n2408), .ZN(n2730) );
  AND2_X1 U2730 ( .A1(n2302), .A2(n2274), .ZN(n2273) );
  NAND2_X1 U2731 ( .A1(n2254), .A2(n3084), .ZN(n4064) );
  NAND2_X1 U2732 ( .A1(n2237), .A2(n2236), .ZN(n4100) );
  AND2_X1 U2733 ( .A1(n2445), .A2(n2435), .ZN(n4406) );
  INV_X1 U2734 ( .A(n4406), .ZN(n2180) );
  AND2_X1 U2735 ( .A1(n3944), .A2(n3062), .ZN(n2052) );
  XNOR2_X1 U2736 ( .A(n3586), .B(n3839), .ZN(n4280) );
  OR2_X1 U2737 ( .A1(n4464), .A2(n2461), .ZN(n2053) );
  NOR2_X1 U2738 ( .A1(n4527), .A2(n4001), .ZN(n2054) );
  NAND2_X1 U2739 ( .A1(n4564), .A2(n2192), .ZN(n2055) );
  AND2_X1 U2740 ( .A1(n2341), .A2(n2340), .ZN(n2056) );
  INV_X1 U2741 ( .A(n2155), .ZN(n3631) );
  OAI21_X1 U2742 ( .B1(n3155), .B2(n2151), .A(n2149), .ZN(n2155) );
  AND2_X1 U2743 ( .A1(n2146), .A2(n2143), .ZN(n2057) );
  AND2_X1 U2744 ( .A1(n2228), .A2(n2227), .ZN(n2058) );
  AND2_X1 U2745 ( .A1(n2572), .A2(n2558), .ZN(n2059) );
  AND2_X1 U2746 ( .A1(n2273), .A2(n2306), .ZN(n2060) );
  INV_X1 U2747 ( .A(n3259), .ZN(n2179) );
  INV_X1 U2748 ( .A(n2472), .ZN(n2487) );
  INV_X1 U2749 ( .A(IR_REG_22__SCAN_IN), .ZN(n2340) );
  AND2_X1 U2750 ( .A1(n4036), .A2(n4603), .ZN(n2061) );
  INV_X1 U2751 ( .A(n4102), .ZN(n2222) );
  OAI21_X1 U2752 ( .B1(n2666), .B2(n2665), .A(n2664), .ZN(n3674) );
  AND2_X1 U2753 ( .A1(n4086), .A2(n3086), .ZN(n2062) );
  INV_X1 U2754 ( .A(n3509), .ZN(n2117) );
  NOR2_X1 U2755 ( .A1(n3072), .A2(n2290), .ZN(n2063) );
  AND2_X1 U2756 ( .A1(n4171), .A2(n3081), .ZN(n2064) );
  INV_X1 U2757 ( .A(n3664), .ZN(n2141) );
  OR2_X1 U2758 ( .A1(n4086), .A2(n3086), .ZN(n2065) );
  AND3_X1 U2759 ( .A1(n2259), .A2(n2294), .A3(n2176), .ZN(n2547) );
  OR2_X1 U2760 ( .A1(n4126), .A2(n3806), .ZN(n2066) );
  INV_X1 U2761 ( .A(n2683), .ZN(n2137) );
  NAND2_X1 U2762 ( .A1(n2097), .A2(n2296), .ZN(n2584) );
  NAND2_X1 U2763 ( .A1(n2792), .A2(n2791), .ZN(n2067) );
  INV_X1 U2764 ( .A(n3534), .ZN(n2284) );
  AND2_X1 U2765 ( .A1(n3819), .A2(n2226), .ZN(n2068) );
  AND2_X1 U2766 ( .A1(n2152), .A2(n2150), .ZN(n2069) );
  INV_X1 U2767 ( .A(n2244), .ZN(n2243) );
  NAND2_X1 U2768 ( .A1(n2049), .A2(n3080), .ZN(n2244) );
  OR2_X1 U2769 ( .A1(n4464), .A2(n3499), .ZN(n2070) );
  AND2_X1 U2770 ( .A1(n4069), .A2(n4051), .ZN(n2071) );
  AND2_X1 U2771 ( .A1(n2647), .A2(n3620), .ZN(n2072) );
  OR2_X1 U2772 ( .A1(n2129), .A2(n2050), .ZN(n2073) );
  NOR2_X1 U2773 ( .A1(n3636), .A2(n4129), .ZN(n2074) );
  INV_X1 U2774 ( .A(n2168), .ZN(n2167) );
  NOR2_X1 U2775 ( .A1(n3650), .A2(n2169), .ZN(n2168) );
  INV_X1 U2776 ( .A(IR_REG_31__SCAN_IN), .ZN(n3193) );
  OR2_X1 U2777 ( .A1(n2064), .A2(n2246), .ZN(n2075) );
  AND2_X1 U2778 ( .A1(n2225), .A2(n4102), .ZN(n2076) );
  AND2_X1 U2779 ( .A1(n2115), .A2(n3129), .ZN(n2077) );
  INV_X1 U2780 ( .A(n3996), .ZN(n2105) );
  OR2_X1 U2781 ( .A1(n4375), .A2(REG0_REG_28__SCAN_IN), .ZN(n2078) );
  NAND2_X1 U2782 ( .A1(n3422), .A2(n2115), .ZN(n2118) );
  NAND2_X1 U2783 ( .A1(n2263), .A2(n2270), .ZN(n3374) );
  INV_X1 U2784 ( .A(n4115), .ZN(n3806) );
  AND2_X1 U2785 ( .A1(n3767), .A2(n3768), .ZN(n3808) );
  INV_X1 U2786 ( .A(n3808), .ZN(n2281) );
  AND2_X1 U2787 ( .A1(n3941), .A2(n3544), .ZN(n2079) );
  NOR2_X1 U2788 ( .A1(n3176), .A2(n3177), .ZN(n2080) );
  INV_X1 U2789 ( .A(n2134), .ZN(n2132) );
  NOR2_X1 U2790 ( .A1(n3732), .A2(n2135), .ZN(n2134) );
  INV_X1 U2791 ( .A(n2247), .ZN(n2246) );
  NAND2_X1 U2792 ( .A1(n4142), .A2(n3079), .ZN(n2247) );
  AND2_X1 U2793 ( .A1(n2051), .A2(n4092), .ZN(n2081) );
  INV_X2 U2794 ( .A(n3938), .ZN(U4043) );
  INV_X1 U2795 ( .A(n3054), .ZN(n3053) );
  AND2_X1 U2796 ( .A1(n2360), .A2(n4395), .ZN(n2345) );
  OR2_X1 U2797 ( .A1(n4375), .A2(n2199), .ZN(n2082) );
  INV_X1 U2798 ( .A(n4005), .ZN(n4643) );
  INV_X2 U2799 ( .A(n4733), .ZN(n4735) );
  OR2_X1 U2800 ( .A1(n3136), .A2(n3309), .ZN(n4733) );
  INV_X1 U2801 ( .A(n4017), .ZN(n2194) );
  AND2_X1 U2802 ( .A1(n2194), .A2(n2192), .ZN(n2083) );
  INV_X1 U2803 ( .A(IR_REG_10__SCAN_IN), .ZN(n2296) );
  INV_X1 U2804 ( .A(n3952), .ZN(n2233) );
  NAND2_X1 U2805 ( .A1(n4351), .A2(n4375), .ZN(n2200) );
  NAND2_X1 U2806 ( .A1(n3452), .A2(n3855), .ZN(n3096) );
  NAND2_X1 U2807 ( .A1(n4599), .A2(n3854), .ZN(n2084) );
  NAND2_X1 U2808 ( .A1(n4601), .A2(n4600), .ZN(n4599) );
  NAND2_X1 U2809 ( .A1(n3537), .A2(n2089), .ZN(n2085) );
  NAND2_X1 U2810 ( .A1(n2085), .A2(n2086), .ZN(n4249) );
  NAND3_X1 U2811 ( .A1(n2092), .A2(n4390), .A3(REG1_REG_1__SCAN_IN), .ZN(n2232) );
  AND2_X1 U2812 ( .A1(n2394), .A2(n2232), .ZN(n2231) );
  NOR2_X2 U2813 ( .A1(n4389), .A2(n4390), .ZN(n2390) );
  NOR2_X1 U2815 ( .A1(n2304), .A2(n2342), .ZN(n2305) );
  INV_X2 U2816 ( .A(n2549), .ZN(n2097) );
  INV_X1 U2817 ( .A(n2304), .ZN(n2096) );
  NAND2_X1 U2818 ( .A1(n2096), .A2(n2095), .ZN(n3194) );
  OAI21_X2 U2819 ( .B1(n3370), .B2(n3099), .A(n3880), .ZN(n3427) );
  NAND2_X1 U2820 ( .A1(n2835), .A2(n2112), .ZN(n2332) );
  XNOR2_X1 U2821 ( .A(n2835), .B(n2112), .ZN(n3208) );
  INV_X1 U2822 ( .A(n3455), .ZN(n3052) );
  MUX2_X1 U2823 ( .A(n3971), .B(n2415), .S(n3787), .Z(n3455) );
  OR2_X1 U2824 ( .A1(n2041), .A2(n2377), .ZN(n2114) );
  INV_X1 U2825 ( .A(n2118), .ZN(n4708) );
  NAND2_X1 U2826 ( .A1(n4056), .A2(n2121), .ZN(n4272) );
  NAND2_X1 U2827 ( .A1(n4056), .A2(n4038), .ZN(n4037) );
  NAND2_X1 U2828 ( .A1(n2125), .A2(n3289), .ZN(n2407) );
  XNOR2_X1 U2829 ( .A(n2125), .B(n3289), .ZN(n3293) );
  OAI22_X2 U2830 ( .A1(n3674), .A2(n2073), .B1(n2127), .B2(n2050), .ZN(n3142)
         );
  NAND2_X1 U2831 ( .A1(n3667), .A2(n3664), .ZN(n2146) );
  INV_X1 U2832 ( .A(n2873), .ZN(n2840) );
  NAND2_X1 U2833 ( .A1(n2173), .A2(n2059), .ZN(n3184) );
  NAND2_X1 U2834 ( .A1(n2176), .A2(n2258), .ZN(n2466) );
  AND2_X1 U2835 ( .A1(n2259), .A2(n2176), .ZN(n2482) );
  NAND2_X1 U2836 ( .A1(n2422), .A2(n2425), .ZN(n3282) );
  NAND2_X2 U2837 ( .A1(n2232), .A2(n2394), .ZN(n3049) );
  MUX2_X1 U2838 ( .A(n3246), .B(REG1_REG_1__SCAN_IN), .S(n3952), .Z(n3950) );
  XNOR2_X2 U2839 ( .A(n2183), .B(n2395), .ZN(n3952) );
  NAND2_X1 U2840 ( .A1(n4564), .A2(n2083), .ZN(n2187) );
  OAI211_X1 U2841 ( .C1(n4564), .C2(n2191), .A(n2188), .B(n2187), .ZN(n4027)
         );
  NAND2_X1 U2842 ( .A1(n4564), .A2(n2195), .ZN(n4008) );
  OR2_X1 U2843 ( .A1(n4048), .A2(n3916), .ZN(n2218) );
  NAND2_X1 U2844 ( .A1(n2209), .A2(n2207), .ZN(n3589) );
  NAND2_X1 U2845 ( .A1(n4048), .A2(n2212), .ZN(n2209) );
  NAND2_X1 U2846 ( .A1(n2218), .A2(n3115), .ZN(n4032) );
  AOI21_X1 U2847 ( .B1(n4246), .B2(n2076), .A(n2220), .ZN(n3113) );
  INV_X1 U2848 ( .A(n3128), .ZN(n2230) );
  OAI21_X2 U2849 ( .B1(n3787), .B2(n2233), .A(n2229), .ZN(n3128) );
  NAND2_X1 U2850 ( .A1(n3852), .A2(n3854), .ZN(n3095) );
  NAND2_X1 U2851 ( .A1(n4158), .A2(n2239), .ZN(n2237) );
  OAI21_X1 U2852 ( .B1(n4158), .B2(n2241), .A(n2239), .ZN(n4122) );
  NAND2_X1 U2853 ( .A1(n2248), .A2(n2250), .ZN(n3088) );
  NAND2_X1 U2854 ( .A1(n4080), .A2(n2251), .ZN(n2248) );
  OAI21_X1 U2855 ( .B1(n2261), .B2(n3061), .A(n3060), .ZN(n2260) );
  NAND2_X1 U2856 ( .A1(n3493), .A2(n2264), .ZN(n2263) );
  NAND2_X1 U2857 ( .A1(n3493), .A2(n2266), .ZN(n2265) );
  NAND2_X1 U2858 ( .A1(n3072), .A2(n2279), .ZN(n2278) );
  XNOR2_X1 U2859 ( .A(n2334), .B(n2333), .ZN(n2819) );
  NAND2_X1 U2860 ( .A1(n2332), .A2(IR_REG_31__SCAN_IN), .ZN(n2334) );
  OR2_X1 U2861 ( .A1(n2421), .A2(n2420), .ZN(n2422) );
  NAND2_X1 U2862 ( .A1(n3163), .A2(n4640), .ZN(n3207) );
  NOR2_X1 U2863 ( .A1(n3631), .A2(n2766), .ZN(n3686) );
  NAND2_X1 U2864 ( .A1(n2632), .A2(n2315), .ZN(n2634) );
  OR2_X1 U2865 ( .A1(n3128), .A2(n2397), .ZN(n2398) );
  OAI21_X2 U2866 ( .B1(n4028), .B2(n3091), .A(n3090), .ZN(n3585) );
  NAND2_X1 U2867 ( .A1(n3787), .A2(DATAI_0_), .ZN(n2376) );
  NAND2_X1 U2868 ( .A1(n2872), .A2(n2871), .ZN(n2285) );
  AND3_X1 U2869 ( .A1(n2844), .A2(n2845), .A3(n4424), .ZN(n2286) );
  NAND2_X1 U2870 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n2287) );
  AND2_X1 U2871 ( .A1(n3738), .A2(n4188), .ZN(n2288) );
  AND2_X1 U2872 ( .A1(n4478), .A2(REG1_REG_7__SCAN_IN), .ZN(n2289) );
  AND2_X1 U2873 ( .A1(n4582), .A2(n3103), .ZN(n2290) );
  NOR2_X1 U2874 ( .A1(n2517), .A2(n2516), .ZN(n2291) );
  INV_X1 U2875 ( .A(n4191), .ZN(n3076) );
  INV_X1 U2876 ( .A(IR_REG_0__SCAN_IN), .ZN(n2377) );
  NAND2_X1 U2877 ( .A1(n2765), .A2(n2764), .ZN(n2766) );
  INV_X1 U2878 ( .A(n3633), .ZN(n2751) );
  INV_X1 U2879 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2559) );
  NAND2_X1 U2880 ( .A1(n3241), .A2(n2861), .ZN(n2347) );
  NOR2_X1 U2881 ( .A1(n3329), .A2(n2494), .ZN(n2495) );
  INV_X1 U2882 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2613) );
  OR2_X1 U2883 ( .A1(n2459), .A2(n2458), .ZN(n3346) );
  NAND2_X1 U2884 ( .A1(n2717), .A2(REG3_REG_21__SCAN_IN), .ZN(n2731) );
  INV_X1 U2885 ( .A(n3282), .ZN(n2423) );
  OR2_X1 U2886 ( .A1(n4602), .A2(n2837), .ZN(n2848) );
  AOI21_X1 U2887 ( .B1(n4646), .B2(REG1_REG_15__SCAN_IN), .A(n4541), .ZN(n4003) );
  OR2_X1 U2888 ( .A1(n3508), .A2(n3064), .ZN(n3066) );
  INV_X1 U2889 ( .A(n3625), .ZN(n3556) );
  OAI22_X1 U2890 ( .A1(n3406), .A2(n3056), .B1(n3859), .B2(n3407), .ZN(n3301)
         );
  OR2_X1 U2891 ( .A1(n2626), .A2(n2613), .ZN(n2649) );
  INV_X1 U2892 ( .A(n4195), .ZN(n4188) );
  NOR2_X1 U2893 ( .A1(n2520), .A2(n2308), .ZN(n2540) );
  OR2_X1 U2894 ( .A1(n2739), .A2(n3635), .ZN(n2754) );
  NAND2_X1 U2895 ( .A1(n2540), .A2(REG3_REG_9__SCAN_IN), .ZN(n2560) );
  NAND2_X1 U2896 ( .A1(n2424), .A2(n2423), .ZN(n3280) );
  NOR2_X1 U2897 ( .A1(n3997), .A2(n4506), .ZN(n4517) );
  INV_X1 U2898 ( .A(REG3_REG_15__SCAN_IN), .ZN(n3760) );
  AND2_X1 U2899 ( .A1(n3835), .A2(n4046), .ZN(n4065) );
  OR2_X1 U2900 ( .A1(n2578), .A2(n3393), .ZN(n2595) );
  INV_X1 U2901 ( .A(n4617), .ZN(n4235) );
  OR3_X1 U2902 ( .A1(n4679), .A2(n3207), .A3(n4395), .ZN(n4255) );
  INV_X1 U2903 ( .A(n4602), .ZN(n4267) );
  INV_X1 U2904 ( .A(n4627), .ZN(n4581) );
  INV_X1 U2905 ( .A(n4222), .ZN(n4229) );
  INV_X1 U2906 ( .A(n3103), .ZN(n3658) );
  AND2_X1 U2907 ( .A1(n2360), .A2(n4397), .ZN(n4623) );
  INV_X1 U2908 ( .A(IR_REG_4__SCAN_IN), .ZN(n2446) );
  INV_X1 U2909 ( .A(n4143), .ZN(n3636) );
  AND2_X1 U2910 ( .A1(n2651), .A2(REG3_REG_16__SCAN_IN), .ZN(n2667) );
  NOR2_X1 U2911 ( .A1(n2754), .A2(n3692), .ZN(n2769) );
  INV_X1 U2912 ( .A(n4429), .ZN(n3751) );
  AND2_X1 U2913 ( .A1(n2839), .A2(n2838), .ZN(n4424) );
  NAND2_X1 U2914 ( .A1(n4009), .A2(n2287), .ZN(n4010) );
  AND2_X1 U2915 ( .A1(n4440), .A2(n3225), .ZN(n4536) );
  AND2_X1 U2916 ( .A1(n4391), .A2(n3209), .ZN(n4603) );
  AND2_X1 U2917 ( .A1(n3379), .A2(n2707), .ZN(n4215) );
  AND2_X1 U2918 ( .A1(n4215), .A2(n4715), .ZN(n4617) );
  INV_X1 U2919 ( .A(n4255), .ZN(n4629) );
  OAI21_X1 U2920 ( .B1(n3199), .B2(D_REG_0__SCAN_IN), .A(n3205), .ZN(n3309) );
  INV_X1 U2921 ( .A(n3309), .ZN(n3135) );
  INV_X1 U2922 ( .A(n4716), .ZN(n4679) );
  INV_X1 U2923 ( .A(n4337), .ZN(n4704) );
  AND2_X1 U2924 ( .A1(n4623), .A2(n2856), .ZN(n4716) );
  NAND2_X1 U2925 ( .A1(n2821), .A2(n4392), .ZN(n3199) );
  AND2_X1 U2926 ( .A1(n2675), .A2(n2691), .ZN(n4005) );
  AND2_X1 U2927 ( .A1(n3224), .A2(n3211), .ZN(n4563) );
  INV_X1 U2928 ( .A(n4424), .ZN(n3753) );
  OAI21_X1 U2929 ( .B1(n3601), .B2(n2811), .A(n2810), .ZN(n4036) );
  OR2_X1 U2930 ( .A1(n3163), .A2(n3204), .ZN(n3938) );
  AND2_X1 U2931 ( .A1(n3480), .A2(n3479), .ZN(n4712) );
  NAND2_X1 U2932 ( .A1(n4735), .A2(n4715), .ZN(n4328) );
  OR2_X1 U2933 ( .A1(n3599), .A2(n4384), .ZN(n3138) );
  NOR2_X2 U2934 ( .A1(n3136), .A2(n3135), .ZN(n4375) );
  AND2_X1 U2935 ( .A1(n4712), .A2(n4711), .ZN(n4732) );
  INV_X1 U2936 ( .A(n4375), .ZN(n4720) );
  NAND2_X1 U2937 ( .A1(n3200), .A2(n3199), .ZN(n4639) );
  INV_X1 U2938 ( .A(n4535), .ZN(n4649) );
  INV_X1 U2939 ( .A(n4478), .ZN(n4657) );
  OR4_X1 U2940 ( .A1(n3152), .A2(n3151), .A3(n3150), .A4(n3149), .ZN(U3230) );
  NAND2_X1 U2941 ( .A1(n2413), .A2(n2414), .ZN(n2432) );
  NAND2_X1 U2942 ( .A1(n2433), .A2(n2446), .ZN(n2292) );
  NOR2_X1 U2943 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2301)
         );
  NOR2_X1 U2944 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2300)
         );
  NOR2_X1 U2945 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_13__SCAN_IN), .ZN(n2299)
         );
  NAND2_X1 U2946 ( .A1(n2341), .A2(n2058), .ZN(n2304) );
  AND2_X2 U2947 ( .A1(n4389), .A2(n2310), .ZN(n2391) );
  INV_X1 U2948 ( .A(n2391), .ZN(n2408) );
  NAND2_X1 U2949 ( .A1(n2730), .A2(REG2_REG_21__SCAN_IN), .ZN(n2314) );
  NAND2_X1 U2950 ( .A1(REG3_REG_7__SCAN_IN), .A2(REG3_REG_8__SCAN_IN), .ZN(
        n2308) );
  NAND2_X1 U2951 ( .A1(n2625), .A2(REG3_REG_13__SCAN_IN), .ZN(n2626) );
  INV_X1 U2952 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2684) );
  INV_X1 U2953 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2700) );
  OR2_X1 U2954 ( .A1(n2717), .A2(REG3_REG_21__SCAN_IN), .ZN(n2309) );
  AND2_X1 U2955 ( .A1(n2731), .A2(n2309), .ZN(n3157) );
  NAND2_X1 U2956 ( .A1(n2389), .A2(n3157), .ZN(n2313) );
  NAND2_X1 U2957 ( .A1(n2043), .A2(REG0_REG_21__SCAN_IN), .ZN(n2312) );
  INV_X1 U2958 ( .A(REG1_REG_21__SCAN_IN), .ZN(n2877) );
  OR2_X1 U2959 ( .A1(n3786), .A2(n2877), .ZN(n2311) );
  NAND4_X1 U2960 ( .A1(n2314), .A2(n2313), .A3(n2312), .A4(n2311), .ZN(n4171)
         );
  INV_X1 U2961 ( .A(n2316), .ZN(n2317) );
  NOR2_X1 U2962 ( .A1(n2317), .A2(IR_REG_16__SCAN_IN), .ZN(n2318) );
  OAI21_X2 U2963 ( .B1(n2691), .B2(IR_REG_18__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2353) );
  INV_X1 U2964 ( .A(IR_REG_19__SCAN_IN), .ZN(n2320) );
  NAND2_X1 U2965 ( .A1(n2353), .A2(n2320), .ZN(n2355) );
  NAND2_X1 U2966 ( .A1(n2342), .A2(IR_REG_31__SCAN_IN), .ZN(n2323) );
  INV_X1 U2967 ( .A(n2342), .ZN(n2324) );
  NAND2_X1 U2968 ( .A1(n2324), .A2(n2341), .ZN(n2357) );
  INV_X1 U2969 ( .A(n2357), .ZN(n2325) );
  MUX2_X1 U2970 ( .A(IR_REG_31__SCAN_IN), .B(n2327), .S(IR_REG_25__SCAN_IN), 
        .Z(n2330) );
  NOR2_X2 U2971 ( .A1(n2331), .A2(n2328), .ZN(n2336) );
  INV_X1 U2972 ( .A(n2336), .ZN(n2329) );
  NAND2_X1 U2973 ( .A1(n2330), .A2(n2329), .ZN(n3198) );
  NOR2_X1 U2974 ( .A1(n3198), .A2(n2819), .ZN(n2344) );
  NAND2_X2 U2975 ( .A1(n2344), .A2(n4392), .ZN(n3163) );
  NAND2_X1 U2976 ( .A1(n4171), .A2(n2047), .ZN(n2352) );
  NAND2_X1 U2977 ( .A1(n2861), .A2(IR_REG_28__SCAN_IN), .ZN(n2349) );
  NAND2_X1 U2978 ( .A1(n3787), .A2(DATAI_21_), .ZN(n4151) );
  OR2_X1 U2979 ( .A1(n2397), .A2(n4151), .ZN(n2351) );
  NAND2_X1 U2980 ( .A1(n2352), .A2(n2351), .ZN(n2359) );
  INV_X1 U2981 ( .A(n2353), .ZN(n2354) );
  NAND2_X1 U2982 ( .A1(n2354), .A2(IR_REG_19__SCAN_IN), .ZN(n2356) );
  NAND2_X1 U2983 ( .A1(n2356), .A2(n2355), .ZN(n2707) );
  NAND2_X1 U2984 ( .A1(n2357), .A2(IR_REG_31__SCAN_IN), .ZN(n2358) );
  NAND2_X1 U2985 ( .A1(n2707), .A2(n4394), .ZN(n2852) );
  XNOR2_X1 U2986 ( .A(n2359), .B(n2814), .ZN(n3153) );
  INV_X1 U2987 ( .A(n3153), .ZN(n2729) );
  INV_X1 U2988 ( .A(n4394), .ZN(n2856) );
  INV_X1 U2989 ( .A(n4395), .ZN(n3123) );
  NAND2_X1 U2990 ( .A1(n4171), .A2(n2045), .ZN(n2362) );
  OR2_X1 U2991 ( .A1(n2853), .A2(n4151), .ZN(n2361) );
  NAND2_X1 U2992 ( .A1(n2362), .A2(n2361), .ZN(n2728) );
  NOR2_X1 U2993 ( .A1(n2651), .A2(REG3_REG_16__SCAN_IN), .ZN(n2363) );
  OR2_X1 U2994 ( .A1(n2667), .A2(n2363), .ZN(n4428) );
  INV_X1 U2995 ( .A(n4428), .ZN(n2364) );
  NAND2_X1 U2996 ( .A1(n2780), .A2(n2364), .ZN(n2368) );
  NAND2_X1 U2997 ( .A1(n2391), .A2(REG2_REG_16__SCAN_IN), .ZN(n2367) );
  NAND2_X1 U2998 ( .A1(n2043), .A2(REG0_REG_16__SCAN_IN), .ZN(n2366) );
  INV_X1 U2999 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4554) );
  OR2_X1 U3000 ( .A1(n3786), .A2(n4554), .ZN(n2365) );
  NAND4_X1 U3001 ( .A1(n2368), .A2(n2367), .A3(n2366), .A4(n2365), .ZN(n4224)
         );
  NAND2_X1 U3002 ( .A1(n4224), .A2(n2047), .ZN(n2374) );
  OAI21_X1 U3003 ( .B1(n2634), .B2(IR_REG_14__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2656) );
  INV_X1 U3004 ( .A(IR_REG_15__SCAN_IN), .ZN(n2369) );
  NAND2_X1 U3005 ( .A1(n2656), .A2(n2369), .ZN(n2370) );
  NAND2_X1 U3006 ( .A1(n2370), .A2(IR_REG_31__SCAN_IN), .ZN(n2372) );
  INV_X1 U3007 ( .A(IR_REG_16__SCAN_IN), .ZN(n2371) );
  INV_X1 U3008 ( .A(DATAI_16_), .ZN(n4644) );
  MUX2_X1 U3009 ( .A(n4645), .B(n4644), .S(n3787), .Z(n3576) );
  OR2_X1 U3010 ( .A1(n3576), .A2(n2397), .ZN(n2373) );
  NAND2_X1 U3011 ( .A1(n2374), .A2(n2373), .ZN(n2375) );
  XNOR2_X1 U3012 ( .A(n2375), .B(n2042), .ZN(n2666) );
  INV_X1 U3013 ( .A(n3576), .ZN(n4418) );
  AOI22_X1 U3014 ( .A1(n4224), .A2(n2472), .B1(n2048), .B2(n4418), .ZN(n2661)
         );
  INV_X1 U3015 ( .A(n2661), .ZN(n2665) );
  NOR2_X1 U3016 ( .A1(n3163), .A2(n2377), .ZN(n2378) );
  AOI21_X1 U3017 ( .B1(n4612), .B2(n2047), .A(n2378), .ZN(n2384) );
  INV_X1 U3018 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4723) );
  NAND2_X1 U3019 ( .A1(n2390), .A2(REG0_REG_0__SCAN_IN), .ZN(n2381) );
  NAND2_X1 U3020 ( .A1(n2391), .A2(REG2_REG_0__SCAN_IN), .ZN(n2380) );
  NAND2_X1 U3021 ( .A1(n2389), .A2(REG3_REG_0__SCAN_IN), .ZN(n2379) );
  NAND4_X1 U3022 ( .A1(n2382), .A2(n2381), .A3(n2380), .A4(n2379), .ZN(n3050)
         );
  NAND2_X1 U3023 ( .A1(n3050), .A2(n2045), .ZN(n2383) );
  NAND2_X1 U3024 ( .A1(n2384), .A2(n2383), .ZN(n3295) );
  NAND2_X1 U3025 ( .A1(n3050), .A2(n2048), .ZN(n2385) );
  NAND2_X1 U3026 ( .A1(n4612), .A2(n2816), .ZN(n2386) );
  OAI211_X1 U3027 ( .C1(n3163), .C2(n4723), .A(n2385), .B(n2386), .ZN(n3294)
         );
  NAND2_X1 U3028 ( .A1(n3295), .A2(n3294), .ZN(n2388) );
  NAND2_X1 U3029 ( .A1(n2386), .A2(n2788), .ZN(n2387) );
  NAND2_X1 U3030 ( .A1(n2388), .A2(n2387), .ZN(n3289) );
  INV_X1 U3031 ( .A(REG1_REG_1__SCAN_IN), .ZN(n3246) );
  NAND2_X1 U3032 ( .A1(n2389), .A2(REG3_REG_1__SCAN_IN), .ZN(n2393) );
  NAND2_X1 U3033 ( .A1(n2391), .A2(REG2_REG_1__SCAN_IN), .ZN(n2392) );
  NAND2_X1 U3034 ( .A1(n3049), .A2(n2047), .ZN(n2399) );
  INV_X1 U3035 ( .A(DATAI_1_), .ZN(n2396) );
  NOR2_X1 U3036 ( .A1(n3128), .A2(n2401), .ZN(n2402) );
  INV_X1 U3037 ( .A(n2403), .ZN(n2405) );
  OR2_X1 U3038 ( .A1(n2405), .A2(n2404), .ZN(n2406) );
  NAND2_X1 U3039 ( .A1(n2407), .A2(n2406), .ZN(n3283) );
  INV_X1 U3040 ( .A(n3283), .ZN(n2424) );
  NAND2_X1 U3041 ( .A1(n2389), .A2(REG3_REG_2__SCAN_IN), .ZN(n2412) );
  INV_X1 U3042 ( .A(REG1_REG_2__SCAN_IN), .ZN(n3245) );
  NAND2_X1 U3043 ( .A1(n2390), .A2(REG0_REG_2__SCAN_IN), .ZN(n2410) );
  NAND2_X1 U3044 ( .A1(n2391), .A2(REG2_REG_2__SCAN_IN), .ZN(n2409) );
  NAND2_X1 U3045 ( .A1(n3054), .A2(n2047), .ZN(n2417) );
  INV_X1 U3046 ( .A(DATAI_2_), .ZN(n2415) );
  OR2_X1 U3047 ( .A1(n3455), .A2(n2397), .ZN(n2416) );
  NAND2_X1 U3048 ( .A1(n2417), .A2(n2416), .ZN(n2418) );
  XNOR2_X1 U3049 ( .A(n2418), .B(n2788), .ZN(n2421) );
  NOR2_X1 U3050 ( .A1(n3455), .A2(n2853), .ZN(n2419) );
  AOI21_X1 U3051 ( .B1(n3054), .B2(n2472), .A(n2419), .ZN(n2420) );
  NAND2_X1 U3052 ( .A1(n2421), .A2(n2420), .ZN(n2425) );
  NAND2_X1 U3053 ( .A1(n3280), .A2(n2425), .ZN(n3272) );
  INV_X1 U3054 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2426) );
  NAND2_X1 U3055 ( .A1(n2780), .A2(n2426), .ZN(n2431) );
  NAND2_X1 U3056 ( .A1(n2730), .A2(REG2_REG_3__SCAN_IN), .ZN(n2430) );
  NAND2_X1 U3057 ( .A1(n2390), .A2(REG0_REG_3__SCAN_IN), .ZN(n2429) );
  INV_X1 U3058 ( .A(REG1_REG_3__SCAN_IN), .ZN(n2427) );
  OR2_X1 U3059 ( .A1(n3786), .A2(n2427), .ZN(n2428) );
  NAND4_X1 U3060 ( .A1(n2431), .A2(n2430), .A3(n2429), .A4(n2428), .ZN(n3948)
         );
  NAND2_X1 U3061 ( .A1(n3948), .A2(n2048), .ZN(n2437) );
  NAND2_X1 U3062 ( .A1(n2432), .A2(IR_REG_31__SCAN_IN), .ZN(n2434) );
  NAND2_X1 U3063 ( .A1(n2434), .A2(n2433), .ZN(n2445) );
  OR2_X1 U3064 ( .A1(n2434), .A2(n2433), .ZN(n2435) );
  MUX2_X1 U3065 ( .A(n4406), .B(DATAI_3_), .S(n3787), .Z(n3860) );
  NAND2_X1 U3066 ( .A1(n3860), .A2(n2816), .ZN(n2436) );
  NAND2_X1 U3067 ( .A1(n2437), .A2(n2436), .ZN(n2438) );
  XNOR2_X1 U3068 ( .A(n2438), .B(n2042), .ZN(n2453) );
  AND2_X1 U3069 ( .A1(n3860), .A2(n2047), .ZN(n2439) );
  AOI21_X1 U3070 ( .B1(n3948), .B2(n2472), .A(n2439), .ZN(n2454) );
  XNOR2_X1 U3071 ( .A(n2453), .B(n2454), .ZN(n3273) );
  NAND2_X1 U3072 ( .A1(n3272), .A2(n3273), .ZN(n3271) );
  NAND2_X1 U3073 ( .A1(n2730), .A2(REG2_REG_4__SCAN_IN), .ZN(n2444) );
  INV_X1 U3074 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2440) );
  XNOR2_X1 U3075 ( .A(n2440), .B(REG3_REG_3__SCAN_IN), .ZN(n3317) );
  NAND2_X1 U3076 ( .A1(n2780), .A2(n3317), .ZN(n2443) );
  NAND2_X1 U3077 ( .A1(n2043), .A2(REG0_REG_4__SCAN_IN), .ZN(n2442) );
  INV_X1 U3078 ( .A(REG1_REG_4__SCAN_IN), .ZN(n3255) );
  OR2_X1 U3079 ( .A1(n3786), .A2(n3255), .ZN(n2441) );
  NAND4_X1 U3080 ( .A1(n2444), .A2(n2443), .A3(n2442), .A4(n2441), .ZN(n3947)
         );
  NAND2_X1 U3081 ( .A1(n3947), .A2(n2047), .ZN(n2450) );
  NAND2_X1 U3082 ( .A1(n2445), .A2(IR_REG_31__SCAN_IN), .ZN(n2447) );
  XNOR2_X1 U3083 ( .A(n2447), .B(n2446), .ZN(n3253) );
  INV_X1 U3084 ( .A(DATAI_4_), .ZN(n2448) );
  MUX2_X1 U3085 ( .A(n3253), .B(n2448), .S(n3787), .Z(n3322) );
  OR2_X1 U3086 ( .A1(n3322), .A2(n2397), .ZN(n2449) );
  NAND2_X1 U3087 ( .A1(n2450), .A2(n2449), .ZN(n2451) );
  XNOR2_X1 U3088 ( .A(n2451), .B(n2042), .ZN(n2457) );
  NOR2_X1 U3089 ( .A1(n3322), .A2(n2853), .ZN(n2452) );
  AOI21_X1 U3090 ( .B1(n3947), .B2(n2472), .A(n2452), .ZN(n2458) );
  XNOR2_X1 U3091 ( .A(n2457), .B(n2458), .ZN(n3319) );
  INV_X1 U3092 ( .A(n2453), .ZN(n2455) );
  NAND2_X1 U3093 ( .A1(n2455), .A2(n2454), .ZN(n3318) );
  AND2_X1 U3094 ( .A1(n3319), .A2(n3318), .ZN(n2456) );
  NAND2_X2 U3095 ( .A1(n3271), .A2(n2456), .ZN(n3347) );
  INV_X1 U3096 ( .A(n2457), .ZN(n2459) );
  NAND2_X1 U3097 ( .A1(n2730), .A2(REG2_REG_5__SCAN_IN), .ZN(n2465) );
  AOI21_X1 U3098 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        REG3_REG_5__SCAN_IN), .ZN(n2460) );
  NOR2_X1 U3099 ( .A1(n2460), .A2(n2474), .ZN(n3344) );
  NAND2_X1 U3100 ( .A1(n2780), .A2(n3344), .ZN(n2464) );
  NAND2_X1 U3101 ( .A1(n2390), .A2(REG0_REG_5__SCAN_IN), .ZN(n2463) );
  INV_X1 U3102 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2461) );
  OR2_X1 U3103 ( .A1(n3786), .A2(n2461), .ZN(n2462) );
  NAND4_X1 U3104 ( .A1(n2465), .A2(n2464), .A3(n2463), .A4(n2462), .ZN(n3946)
         );
  NAND2_X1 U3105 ( .A1(n3946), .A2(n2047), .ZN(n2469) );
  NAND2_X1 U3106 ( .A1(n2466), .A2(IR_REG_31__SCAN_IN), .ZN(n2467) );
  XNOR2_X1 U3107 ( .A(n2467), .B(IR_REG_5__SCAN_IN), .ZN(n4660) );
  MUX2_X1 U3108 ( .A(n4660), .B(DATAI_5_), .S(n3787), .Z(n3488) );
  NAND2_X1 U3109 ( .A1(n3488), .A2(n2816), .ZN(n2468) );
  NAND2_X1 U3110 ( .A1(n2469), .A2(n2468), .ZN(n2470) );
  XNOR2_X1 U3111 ( .A(n2470), .B(n2042), .ZN(n2492) );
  AND2_X1 U3112 ( .A1(n3488), .A2(n2047), .ZN(n2471) );
  AOI21_X1 U3113 ( .B1(n3946), .B2(n2472), .A(n2471), .ZN(n2491) );
  INV_X1 U3114 ( .A(n2491), .ZN(n2473) );
  NAND2_X1 U3115 ( .A1(n2492), .A2(n2473), .ZN(n2490) );
  AND2_X1 U3116 ( .A1(n3346), .A2(n2490), .ZN(n3328) );
  INV_X1 U3117 ( .A(n2474), .ZN(n2475) );
  INV_X1 U3118 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3337) );
  NAND2_X1 U3119 ( .A1(n2475), .A2(n3337), .ZN(n2476) );
  AND2_X1 U3120 ( .A1(n2476), .A2(n2520), .ZN(n4593) );
  NAND2_X1 U3121 ( .A1(n2780), .A2(n4593), .ZN(n2481) );
  NAND2_X1 U3122 ( .A1(n2730), .A2(REG2_REG_6__SCAN_IN), .ZN(n2480) );
  NAND2_X1 U3123 ( .A1(n2043), .A2(REG0_REG_6__SCAN_IN), .ZN(n2479) );
  INV_X1 U3124 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2477) );
  OR2_X1 U3125 ( .A1(n3786), .A2(n2477), .ZN(n2478) );
  NAND4_X1 U3126 ( .A1(n2481), .A2(n2480), .A3(n2479), .A4(n2478), .ZN(n3945)
         );
  NAND2_X1 U3127 ( .A1(n3945), .A2(n2048), .ZN(n2485) );
  OR2_X1 U3128 ( .A1(n2482), .A2(n3193), .ZN(n2483) );
  XNOR2_X1 U3129 ( .A(n2483), .B(IR_REG_6__SCAN_IN), .ZN(n4473) );
  MUX2_X1 U3130 ( .A(n4473), .B(DATAI_6_), .S(n3787), .Z(n3364) );
  NAND2_X1 U3131 ( .A1(n3364), .A2(n2816), .ZN(n2484) );
  NAND2_X1 U3132 ( .A1(n2485), .A2(n2484), .ZN(n2486) );
  XNOR2_X1 U3133 ( .A(n2486), .B(n2042), .ZN(n2497) );
  NAND2_X1 U3134 ( .A1(n3945), .A2(n2472), .ZN(n2489) );
  NAND2_X1 U3135 ( .A1(n3364), .A2(n2047), .ZN(n2488) );
  NAND2_X1 U3136 ( .A1(n2489), .A2(n2488), .ZN(n2498) );
  AND2_X1 U3137 ( .A1(n2497), .A2(n2498), .ZN(n2494) );
  INV_X1 U3138 ( .A(n2494), .ZN(n3332) );
  AND2_X1 U3139 ( .A1(n3328), .A2(n3332), .ZN(n2496) );
  INV_X1 U3140 ( .A(n2490), .ZN(n2493) );
  XNOR2_X1 U3141 ( .A(n2492), .B(n2491), .ZN(n3345) );
  AOI21_X1 U3142 ( .B1(n3347), .B2(n2496), .A(n2495), .ZN(n2501) );
  INV_X1 U3143 ( .A(n2497), .ZN(n2500) );
  INV_X1 U3144 ( .A(n2498), .ZN(n2499) );
  NAND2_X1 U3145 ( .A1(n2500), .A2(n2499), .ZN(n3331) );
  NAND2_X1 U3146 ( .A1(n2501), .A2(n3331), .ZN(n3176) );
  INV_X1 U3147 ( .A(n3176), .ZN(n2519) );
  NAND2_X1 U31480 ( .A1(n2730), .A2(REG2_REG_7__SCAN_IN), .ZN(n2506) );
  XNOR2_X1 U31490 ( .A(n2520), .B(REG3_REG_7__SCAN_IN), .ZN(n3178) );
  NAND2_X1 U3150 ( .A1(n2780), .A2(n3178), .ZN(n2505) );
  NAND2_X1 U3151 ( .A1(n2043), .A2(REG0_REG_7__SCAN_IN), .ZN(n2504) );
  INV_X1 U3152 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2502) );
  OR2_X1 U3153 ( .A1(n3786), .A2(n2502), .ZN(n2503) );
  NAND4_X1 U3154 ( .A1(n2506), .A2(n2505), .A3(n2504), .A4(n2503), .ZN(n3944)
         );
  NAND2_X1 U3155 ( .A1(n3944), .A2(n2048), .ZN(n2513) );
  NAND2_X1 U3156 ( .A1(n2482), .A2(n2507), .ZN(n2508) );
  NAND2_X1 U3157 ( .A1(n2508), .A2(IR_REG_31__SCAN_IN), .ZN(n2510) );
  NAND2_X1 U3158 ( .A1(n2510), .A2(n2509), .ZN(n2529) );
  OR2_X1 U3159 ( .A1(n2510), .A2(n2509), .ZN(n2511) );
  INV_X1 U3160 ( .A(DATAI_7_), .ZN(n4656) );
  MUX2_X1 U3161 ( .A(n4657), .B(n4656), .S(n3787), .Z(n3869) );
  OR2_X1 U3162 ( .A1(n3869), .A2(n2397), .ZN(n2512) );
  NAND2_X1 U3163 ( .A1(n2513), .A2(n2512), .ZN(n2514) );
  XNOR2_X1 U3164 ( .A(n2514), .B(n2788), .ZN(n2517) );
  NOR2_X1 U3165 ( .A1(n3869), .A2(n2853), .ZN(n2515) );
  AOI21_X1 U3166 ( .B1(n3944), .B2(n2472), .A(n2515), .ZN(n2516) );
  XNOR2_X1 U3167 ( .A(n2517), .B(n2516), .ZN(n3177) );
  INV_X1 U3168 ( .A(n3177), .ZN(n2518) );
  AOI21_X1 U3169 ( .B1(n2519), .B2(n2518), .A(n2291), .ZN(n3165) );
  NAND2_X1 U3170 ( .A1(n2730), .A2(REG2_REG_8__SCAN_IN), .ZN(n2528) );
  INV_X1 U3171 ( .A(n2520), .ZN(n2521) );
  AOI21_X1 U3172 ( .B1(n2521), .B2(REG3_REG_7__SCAN_IN), .A(
        REG3_REG_8__SCAN_IN), .ZN(n2522) );
  OR2_X1 U3173 ( .A1(n2522), .A2(n2540), .ZN(n3423) );
  INV_X1 U3174 ( .A(n3423), .ZN(n2523) );
  NAND2_X1 U3175 ( .A1(n2780), .A2(n2523), .ZN(n2527) );
  NAND2_X1 U3176 ( .A1(n2043), .A2(REG0_REG_8__SCAN_IN), .ZN(n2526) );
  INV_X1 U3177 ( .A(REG1_REG_8__SCAN_IN), .ZN(n2524) );
  OR2_X1 U3178 ( .A1(n3786), .A2(n2524), .ZN(n2525) );
  NAND4_X1 U3179 ( .A1(n2528), .A2(n2527), .A3(n2526), .A4(n2525), .ZN(n3943)
         );
  NAND2_X1 U3180 ( .A1(n3943), .A2(n2047), .ZN(n2532) );
  NAND2_X1 U3181 ( .A1(n2529), .A2(IR_REG_31__SCAN_IN), .ZN(n2530) );
  XNOR2_X1 U3182 ( .A(n2530), .B(IR_REG_8__SCAN_IN), .ZN(n3259) );
  MUX2_X1 U3183 ( .A(n3259), .B(DATAI_8_), .S(n3787), .Z(n3100) );
  NAND2_X1 U3184 ( .A1(n3100), .A2(n2816), .ZN(n2531) );
  NAND2_X1 U3185 ( .A1(n2532), .A2(n2531), .ZN(n2533) );
  XNOR2_X1 U3186 ( .A(n2533), .B(n2042), .ZN(n2536) );
  NAND2_X1 U3187 ( .A1(n3943), .A2(n2472), .ZN(n2535) );
  NAND2_X1 U3188 ( .A1(n3100), .A2(n2048), .ZN(n2534) );
  NAND2_X1 U3189 ( .A1(n2535), .A2(n2534), .ZN(n2537) );
  NAND2_X1 U3190 ( .A1(n2536), .A2(n2537), .ZN(n3166) );
  NAND2_X1 U3191 ( .A1(n3165), .A2(n3166), .ZN(n3164) );
  INV_X1 U3192 ( .A(n2536), .ZN(n2539) );
  INV_X1 U3193 ( .A(n2537), .ZN(n2538) );
  NAND2_X1 U3194 ( .A1(n2539), .A2(n2538), .ZN(n3168) );
  NAND2_X1 U3195 ( .A1(n3164), .A2(n3168), .ZN(n3437) );
  NAND2_X1 U3196 ( .A1(n2730), .A2(REG2_REG_9__SCAN_IN), .ZN(n2546) );
  OR2_X1 U3197 ( .A1(n2540), .A2(REG3_REG_9__SCAN_IN), .ZN(n2541) );
  AND2_X1 U3198 ( .A1(n2560), .A2(n2541), .ZN(n3513) );
  NAND2_X1 U3199 ( .A1(n2780), .A2(n3513), .ZN(n2545) );
  NAND2_X1 U3200 ( .A1(n2043), .A2(REG0_REG_9__SCAN_IN), .ZN(n2544) );
  INV_X1 U3201 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2542) );
  OR2_X1 U3202 ( .A1(n3786), .A2(n2542), .ZN(n2543) );
  NAND4_X1 U3203 ( .A1(n2546), .A2(n2545), .A3(n2544), .A4(n2543), .ZN(n3473)
         );
  NAND2_X1 U3204 ( .A1(n3473), .A2(n2047), .ZN(n2552) );
  NOR2_X1 U3205 ( .A1(n2547), .A2(n3193), .ZN(n2548) );
  MUX2_X1 U3206 ( .A(n3193), .B(n2548), .S(IR_REG_9__SCAN_IN), .Z(n2550) );
  MUX2_X1 U3207 ( .A(n4399), .B(DATAI_9_), .S(n3787), .Z(n3509) );
  NAND2_X1 U3208 ( .A1(n3509), .A2(n2816), .ZN(n2551) );
  NAND2_X1 U3209 ( .A1(n2552), .A2(n2551), .ZN(n2553) );
  XNOR2_X1 U32100 ( .A(n2553), .B(n2042), .ZN(n2555) );
  AND2_X1 U32110 ( .A1(n3509), .A2(n2048), .ZN(n2554) );
  AOI21_X1 U32120 ( .B1(n3473), .B2(n2472), .A(n2554), .ZN(n2556) );
  XNOR2_X1 U32130 ( .A(n2555), .B(n2556), .ZN(n3436) );
  INV_X1 U32140 ( .A(n2555), .ZN(n2557) );
  NAND2_X1 U32150 ( .A1(n2557), .A2(n2556), .ZN(n2558) );
  NAND2_X1 U32160 ( .A1(n2391), .A2(REG2_REG_10__SCAN_IN), .ZN(n2566) );
  NAND2_X1 U32170 ( .A1(n2560), .A2(n2559), .ZN(n2561) );
  AND2_X1 U32180 ( .A1(n2578), .A2(n2561), .ZN(n3188) );
  NAND2_X1 U32190 ( .A1(n2780), .A2(n3188), .ZN(n2565) );
  NAND2_X1 U32200 ( .A1(n2043), .A2(REG0_REG_10__SCAN_IN), .ZN(n2564) );
  INV_X1 U32210 ( .A(REG1_REG_10__SCAN_IN), .ZN(n2562) );
  OR2_X1 U32220 ( .A1(n3786), .A2(n2562), .ZN(n2563) );
  NAND4_X1 U32230 ( .A1(n2566), .A2(n2565), .A3(n2564), .A4(n2563), .ZN(n4580)
         );
  NAND2_X1 U32240 ( .A1(n4580), .A2(n2048), .ZN(n2569) );
  NAND2_X1 U32250 ( .A1(n2549), .A2(IR_REG_31__SCAN_IN), .ZN(n2567) );
  XNOR2_X1 U32260 ( .A(n2567), .B(IR_REG_10__SCAN_IN), .ZN(n3396) );
  MUX2_X1 U32270 ( .A(n3396), .B(DATAI_10_), .S(n3787), .Z(n3481) );
  NAND2_X1 U32280 ( .A1(n3481), .A2(n2816), .ZN(n2568) );
  NAND2_X1 U32290 ( .A1(n2569), .A2(n2568), .ZN(n2570) );
  XNOR2_X1 U32300 ( .A(n2570), .B(n2788), .ZN(n2573) );
  AND2_X1 U32310 ( .A1(n3481), .A2(n2047), .ZN(n2571) );
  AOI21_X1 U32320 ( .B1(n4580), .B2(n2472), .A(n2571), .ZN(n2574) );
  XNOR2_X1 U32330 ( .A(n2573), .B(n2574), .ZN(n3187) );
  INV_X1 U32340 ( .A(n3187), .ZN(n2572) );
  INV_X1 U32350 ( .A(n2573), .ZN(n2576) );
  INV_X1 U32360 ( .A(n2574), .ZN(n2575) );
  NAND2_X1 U32370 ( .A1(n2576), .A2(n2575), .ZN(n2577) );
  NAND2_X2 U32380 ( .A1(n3184), .A2(n2577), .ZN(n3724) );
  NAND2_X1 U32390 ( .A1(n2578), .A2(n3393), .ZN(n2579) );
  AND2_X1 U32400 ( .A1(n2595), .A2(n2579), .ZN(n4588) );
  NAND2_X1 U32410 ( .A1(n2780), .A2(n4588), .ZN(n2583) );
  NAND2_X1 U32420 ( .A1(n2391), .A2(REG2_REG_11__SCAN_IN), .ZN(n2582) );
  NAND2_X1 U32430 ( .A1(n2043), .A2(REG0_REG_11__SCAN_IN), .ZN(n2581) );
  INV_X1 U32440 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3399) );
  OR2_X1 U32450 ( .A1(n3786), .A2(n3399), .ZN(n2580) );
  NAND4_X1 U32460 ( .A1(n2583), .A2(n2582), .A3(n2581), .A4(n2580), .ZN(n3942)
         );
  NAND2_X1 U32470 ( .A1(n3942), .A2(n2048), .ZN(n2590) );
  NAND2_X1 U32480 ( .A1(n2584), .A2(IR_REG_31__SCAN_IN), .ZN(n2586) );
  NAND2_X1 U32490 ( .A1(n2586), .A2(n2585), .ZN(n2602) );
  OR2_X1 U32500 ( .A1(n2586), .A2(n2585), .ZN(n2587) );
  NAND2_X1 U32510 ( .A1(n2602), .A2(n2587), .ZN(n3992) );
  INV_X1 U32520 ( .A(DATAI_11_), .ZN(n2588) );
  MUX2_X1 U32530 ( .A(n3992), .B(n2588), .S(n3787), .Z(n3129) );
  OR2_X1 U32540 ( .A1(n3129), .A2(n2397), .ZN(n2589) );
  NAND2_X1 U32550 ( .A1(n2590), .A2(n2589), .ZN(n2591) );
  XNOR2_X1 U32560 ( .A(n2591), .B(n2042), .ZN(n3721) );
  NAND2_X1 U32570 ( .A1(n3942), .A2(n2472), .ZN(n2593) );
  OR2_X1 U32580 ( .A1(n3129), .A2(n2853), .ZN(n2592) );
  NAND2_X1 U32590 ( .A1(n2593), .A2(n2592), .ZN(n3722) );
  NAND2_X1 U32600 ( .A1(n2391), .A2(REG2_REG_12__SCAN_IN), .ZN(n2601) );
  AND2_X1 U32610 ( .A1(n2595), .A2(n2594), .ZN(n2596) );
  NOR2_X1 U32620 ( .A1(n2625), .A2(n2596), .ZN(n3649) );
  NAND2_X1 U32630 ( .A1(n2780), .A2(n3649), .ZN(n2600) );
  NAND2_X1 U32640 ( .A1(n2043), .A2(REG0_REG_12__SCAN_IN), .ZN(n2599) );
  INV_X1 U32650 ( .A(REG1_REG_12__SCAN_IN), .ZN(n2597) );
  OR2_X1 U32660 ( .A1(n3786), .A2(n2597), .ZN(n2598) );
  NAND4_X1 U32670 ( .A1(n2601), .A2(n2600), .A3(n2599), .A4(n2598), .ZN(n4582)
         );
  NAND2_X1 U32680 ( .A1(n4582), .A2(n2047), .ZN(n2605) );
  NAND2_X1 U32690 ( .A1(n2602), .A2(IR_REG_31__SCAN_IN), .ZN(n2603) );
  XNOR2_X1 U32700 ( .A(n2603), .B(IR_REG_12__SCAN_IN), .ZN(n3996) );
  MUX2_X1 U32710 ( .A(n3996), .B(DATAI_12_), .S(n2041), .Z(n3103) );
  NAND2_X1 U32720 ( .A1(n3103), .A2(n2816), .ZN(n2604) );
  NAND2_X1 U32730 ( .A1(n2605), .A2(n2604), .ZN(n2606) );
  XNOR2_X1 U32740 ( .A(n2606), .B(n2042), .ZN(n2609) );
  NAND2_X1 U32750 ( .A1(n4582), .A2(n2472), .ZN(n2608) );
  NAND2_X1 U32760 ( .A1(n3103), .A2(n2048), .ZN(n2607) );
  NAND2_X1 U32770 ( .A1(n2608), .A2(n2607), .ZN(n2610) );
  AND2_X1 U32780 ( .A1(n2609), .A2(n2610), .ZN(n3650) );
  INV_X1 U32790 ( .A(n2609), .ZN(n2612) );
  INV_X1 U32800 ( .A(n2610), .ZN(n2611) );
  NAND2_X1 U32810 ( .A1(n2612), .A2(n2611), .ZN(n3651) );
  NAND2_X1 U32820 ( .A1(n2730), .A2(REG2_REG_14__SCAN_IN), .ZN(n2618) );
  NAND2_X1 U32830 ( .A1(n2626), .A2(n2613), .ZN(n2614) );
  AND2_X1 U32840 ( .A1(n2649), .A2(n2614), .ZN(n3558) );
  NAND2_X1 U32850 ( .A1(n2780), .A2(n3558), .ZN(n2617) );
  NAND2_X1 U32860 ( .A1(n2043), .A2(REG0_REG_14__SCAN_IN), .ZN(n2616) );
  INV_X1 U32870 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4529) );
  OR2_X1 U32880 ( .A1(n3786), .A2(n4529), .ZN(n2615) );
  NAND4_X1 U32890 ( .A1(n2618), .A2(n2617), .A3(n2616), .A4(n2615), .ZN(n4252)
         );
  NAND2_X1 U32900 ( .A1(n4252), .A2(n2047), .ZN(n2621) );
  NAND2_X1 U32910 ( .A1(n2634), .A2(IR_REG_31__SCAN_IN), .ZN(n2619) );
  XNOR2_X1 U32920 ( .A(n2619), .B(IR_REG_14__SCAN_IN), .ZN(n4535) );
  INV_X1 U32930 ( .A(DATAI_14_), .ZN(n4648) );
  MUX2_X1 U32940 ( .A(n4649), .B(n4648), .S(n3787), .Z(n3625) );
  OR2_X1 U32950 ( .A1(n3625), .A2(n2397), .ZN(n2620) );
  NAND2_X1 U32960 ( .A1(n2621), .A2(n2620), .ZN(n2622) );
  XNOR2_X1 U32970 ( .A(n2622), .B(n2042), .ZN(n2643) );
  NAND2_X1 U32980 ( .A1(n4252), .A2(n2472), .ZN(n2624) );
  OR2_X1 U32990 ( .A1(n3625), .A2(n2853), .ZN(n2623) );
  NAND2_X1 U33000 ( .A1(n2624), .A2(n2623), .ZN(n2644) );
  NAND2_X1 U33010 ( .A1(n2643), .A2(n2644), .ZN(n3621) );
  NAND2_X1 U33020 ( .A1(n2391), .A2(REG2_REG_13__SCAN_IN), .ZN(n2631) );
  OR2_X1 U33030 ( .A1(n2625), .A2(REG3_REG_13__SCAN_IN), .ZN(n2627) );
  AND2_X1 U33040 ( .A1(n2627), .A2(n2626), .ZN(n3697) );
  NAND2_X1 U33050 ( .A1(n2780), .A2(n3697), .ZN(n2630) );
  NAND2_X1 U33060 ( .A1(n2043), .A2(REG0_REG_13__SCAN_IN), .ZN(n2629) );
  INV_X1 U33070 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3998) );
  OR2_X1 U33080 ( .A1(n3786), .A2(n3998), .ZN(n2628) );
  NAND4_X1 U33090 ( .A1(n2631), .A2(n2630), .A3(n2629), .A4(n2628), .ZN(n3941)
         );
  NAND2_X1 U33100 ( .A1(n3941), .A2(n2047), .ZN(n2637) );
  OR2_X1 U33110 ( .A1(n2632), .A2(n3193), .ZN(n2633) );
  MUX2_X1 U33120 ( .A(IR_REG_31__SCAN_IN), .B(n2633), .S(IR_REG_13__SCAN_IN), 
        .Z(n2635) );
  AND2_X1 U33130 ( .A1(n2635), .A2(n2634), .ZN(n3999) );
  MUX2_X1 U33140 ( .A(n3999), .B(DATAI_13_), .S(n3787), .Z(n3544) );
  NAND2_X1 U33150 ( .A1(n3544), .A2(n2816), .ZN(n2636) );
  NAND2_X1 U33160 ( .A1(n2637), .A2(n2636), .ZN(n2638) );
  XNOR2_X1 U33170 ( .A(n2638), .B(n2788), .ZN(n3699) );
  INV_X1 U33180 ( .A(n3699), .ZN(n3617) );
  NAND2_X1 U33190 ( .A1(n3941), .A2(n2472), .ZN(n2640) );
  NAND2_X1 U33200 ( .A1(n3544), .A2(n2048), .ZN(n2639) );
  AND2_X1 U33210 ( .A1(n2640), .A2(n2639), .ZN(n2642) );
  INV_X1 U33220 ( .A(n2642), .ZN(n3698) );
  NAND2_X1 U33230 ( .A1(n3617), .A2(n3698), .ZN(n2641) );
  AND2_X1 U33240 ( .A1(n3621), .A2(n2641), .ZN(n2648) );
  NAND3_X1 U33250 ( .A1(n3621), .A2(n2642), .A3(n3699), .ZN(n2647) );
  INV_X1 U33260 ( .A(n2643), .ZN(n2646) );
  INV_X1 U33270 ( .A(n2644), .ZN(n2645) );
  NAND2_X1 U33280 ( .A1(n2646), .A2(n2645), .ZN(n3620) );
  NAND2_X1 U33290 ( .A1(n2391), .A2(REG2_REG_15__SCAN_IN), .ZN(n2655) );
  AND2_X1 U33300 ( .A1(n2649), .A2(n3760), .ZN(n2650) );
  NOR2_X1 U33310 ( .A1(n2651), .A2(n2650), .ZN(n3755) );
  NAND2_X1 U33320 ( .A1(n2780), .A2(n3755), .ZN(n2654) );
  NAND2_X1 U33330 ( .A1(n2043), .A2(REG0_REG_15__SCAN_IN), .ZN(n2653) );
  INV_X1 U33340 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4002) );
  OR2_X1 U33350 ( .A1(n3786), .A2(n4002), .ZN(n2652) );
  NAND4_X1 U33360 ( .A1(n2655), .A2(n2654), .A3(n2653), .A4(n2652), .ZN(n3940)
         );
  NAND2_X1 U33370 ( .A1(n3940), .A2(n2047), .ZN(n2658) );
  XNOR2_X1 U33380 ( .A(n2656), .B(IR_REG_15__SCAN_IN), .ZN(n4646) );
  MUX2_X1 U33390 ( .A(n4646), .B(DATAI_15_), .S(n2041), .Z(n4254) );
  NAND2_X1 U33400 ( .A1(n4254), .A2(n2816), .ZN(n2657) );
  NAND2_X1 U33410 ( .A1(n2658), .A2(n2657), .ZN(n2659) );
  XNOR2_X1 U33420 ( .A(n2659), .B(n2042), .ZN(n2662) );
  NOR2_X2 U33430 ( .A1(n2663), .A2(n2662), .ZN(n4419) );
  AND2_X1 U33440 ( .A1(n4254), .A2(n2048), .ZN(n2660) );
  AOI21_X1 U33450 ( .B1(n3940), .B2(n2472), .A(n2660), .ZN(n4421) );
  XNOR2_X1 U33460 ( .A(n2666), .B(n2661), .ZN(n4423) );
  NAND2_X1 U33470 ( .A1(n2663), .A2(n2662), .ZN(n4420) );
  OAI211_X1 U33480 ( .C1(n4419), .C2(n4421), .A(n4423), .B(n4420), .ZN(n2664)
         );
  OR2_X1 U33490 ( .A1(n2667), .A2(REG3_REG_17__SCAN_IN), .ZN(n2668) );
  AND2_X1 U33500 ( .A1(n2685), .A2(n2668), .ZN(n4233) );
  NAND2_X1 U33510 ( .A1(n2780), .A2(n4233), .ZN(n2672) );
  NAND2_X1 U33520 ( .A1(n2391), .A2(REG2_REG_17__SCAN_IN), .ZN(n2671) );
  NAND2_X1 U3353 ( .A1(n2043), .A2(REG0_REG_17__SCAN_IN), .ZN(n2670) );
  INV_X1 U33540 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4326) );
  OR2_X1 U3355 ( .A1(n3786), .A2(n4326), .ZN(n2669) );
  NAND4_X1 U3356 ( .A1(n2672), .A2(n2671), .A3(n2670), .A4(n2669), .ZN(n3939)
         );
  NAND2_X1 U3357 ( .A1(n3939), .A2(n2047), .ZN(n2677) );
  NAND2_X1 U3358 ( .A1(n2673), .A2(IR_REG_31__SCAN_IN), .ZN(n2674) );
  MUX2_X1 U3359 ( .A(IR_REG_31__SCAN_IN), .B(n2674), .S(IR_REG_17__SCAN_IN), 
        .Z(n2675) );
  INV_X1 U3360 ( .A(DATAI_17_), .ZN(n4642) );
  MUX2_X1 U3361 ( .A(n4643), .B(n4642), .S(n3787), .Z(n4222) );
  OR2_X1 U3362 ( .A1(n4222), .A2(n2397), .ZN(n2676) );
  NAND2_X1 U3363 ( .A1(n2677), .A2(n2676), .ZN(n2678) );
  XNOR2_X1 U3364 ( .A(n2678), .B(n2042), .ZN(n3676) );
  NAND2_X1 U3365 ( .A1(n3939), .A2(n2472), .ZN(n2680) );
  OR2_X1 U3366 ( .A1(n4222), .A2(n2853), .ZN(n2679) );
  NAND2_X1 U3367 ( .A1(n2680), .A2(n2679), .ZN(n2681) );
  NOR2_X1 U3368 ( .A1(n3676), .A2(n2681), .ZN(n2683) );
  INV_X1 U3369 ( .A(n3676), .ZN(n2682) );
  INV_X1 U3370 ( .A(n2681), .ZN(n3675) );
  NAND2_X1 U3371 ( .A1(n2730), .A2(REG2_REG_18__SCAN_IN), .ZN(n2690) );
  NAND2_X1 U3372 ( .A1(n2685), .A2(n2684), .ZN(n2686) );
  AND2_X1 U3373 ( .A1(n2701), .A2(n2686), .ZN(n4216) );
  NAND2_X1 U3374 ( .A1(n2780), .A2(n4216), .ZN(n2689) );
  NAND2_X1 U3375 ( .A1(n2043), .A2(REG0_REG_18__SCAN_IN), .ZN(n2688) );
  INV_X1 U3376 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4006) );
  OR2_X1 U3377 ( .A1(n3786), .A2(n4006), .ZN(n2687) );
  NAND4_X1 U3378 ( .A1(n2690), .A2(n2689), .A3(n2688), .A4(n2687), .ZN(n4191)
         );
  NAND2_X1 U3379 ( .A1(n4191), .A2(n2048), .ZN(n2695) );
  NAND2_X1 U3380 ( .A1(n2691), .A2(IR_REG_31__SCAN_IN), .ZN(n2692) );
  INV_X1 U3381 ( .A(IR_REG_18__SCAN_IN), .ZN(n2996) );
  XNOR2_X1 U3382 ( .A(n2692), .B(n2996), .ZN(n4014) );
  INV_X1 U3383 ( .A(DATAI_18_), .ZN(n2693) );
  MUX2_X1 U3384 ( .A(n4014), .B(n2693), .S(n2041), .Z(n4213) );
  OR2_X1 U3385 ( .A1(n4213), .A2(n2397), .ZN(n2694) );
  NAND2_X1 U3386 ( .A1(n2695), .A2(n2694), .ZN(n2696) );
  XNOR2_X1 U3387 ( .A(n2696), .B(n2788), .ZN(n2699) );
  NOR2_X1 U3388 ( .A1(n4213), .A2(n2853), .ZN(n2697) );
  AOI21_X1 U3389 ( .B1(n4191), .B2(n2472), .A(n2697), .ZN(n2698) );
  NOR2_X1 U3390 ( .A1(n2699), .A2(n2698), .ZN(n3732) );
  NAND2_X1 U3391 ( .A1(n2699), .A2(n2698), .ZN(n3733) );
  NAND2_X1 U3392 ( .A1(n2391), .A2(REG2_REG_19__SCAN_IN), .ZN(n2706) );
  AND2_X1 U3393 ( .A1(n2701), .A2(n2700), .ZN(n2702) );
  NOR2_X1 U3394 ( .A1(n2715), .A2(n2702), .ZN(n3641) );
  NAND2_X1 U3395 ( .A1(n2780), .A2(n3641), .ZN(n2705) );
  NAND2_X1 U3396 ( .A1(n2043), .A2(REG0_REG_19__SCAN_IN), .ZN(n2704) );
  INV_X1 U3397 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4318) );
  OR2_X1 U3398 ( .A1(n3786), .A2(n4318), .ZN(n2703) );
  NAND4_X1 U3399 ( .A1(n2706), .A2(n2705), .A3(n2704), .A4(n2703), .ZN(n4205)
         );
  MUX2_X1 U3400 ( .A(n4397), .B(DATAI_19_), .S(n3787), .Z(n4195) );
  OAI22_X1 U3401 ( .A1(n3738), .A2(n2487), .B1(n2853), .B2(n4188), .ZN(n2712)
         );
  NAND2_X1 U3402 ( .A1(n4205), .A2(n2048), .ZN(n2709) );
  NAND2_X1 U3403 ( .A1(n4195), .A2(n2816), .ZN(n2708) );
  NAND2_X1 U3404 ( .A1(n2709), .A2(n2708), .ZN(n2710) );
  XNOR2_X1 U3405 ( .A(n2710), .B(n2042), .ZN(n2711) );
  XOR2_X1 U3406 ( .A(n2712), .B(n2711), .Z(n3642) );
  INV_X1 U3407 ( .A(n2711), .ZN(n2714) );
  INV_X1 U3408 ( .A(n2712), .ZN(n2713) );
  NAND2_X1 U3409 ( .A1(n2730), .A2(REG2_REG_20__SCAN_IN), .ZN(n2721) );
  NOR2_X1 U3410 ( .A1(n2715), .A2(REG3_REG_20__SCAN_IN), .ZN(n2716) );
  OR2_X1 U3411 ( .A1(n2717), .A2(n2716), .ZN(n3147) );
  INV_X1 U3412 ( .A(n3147), .ZN(n4178) );
  NAND2_X1 U3413 ( .A1(n2780), .A2(n4178), .ZN(n2720) );
  NAND2_X1 U3414 ( .A1(n2043), .A2(REG0_REG_20__SCAN_IN), .ZN(n2719) );
  INV_X1 U3415 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4314) );
  OR2_X1 U3416 ( .A1(n3786), .A2(n4314), .ZN(n2718) );
  NAND4_X1 U3417 ( .A1(n2721), .A2(n2720), .A3(n2719), .A4(n2718), .ZN(n4142)
         );
  NAND2_X1 U3418 ( .A1(n4142), .A2(n2048), .ZN(n2723) );
  NAND2_X1 U3419 ( .A1(n3787), .A2(DATAI_20_), .ZN(n4177) );
  OR2_X1 U3420 ( .A1(n2397), .A2(n4177), .ZN(n2722) );
  NAND2_X1 U3421 ( .A1(n2723), .A2(n2722), .ZN(n2724) );
  XNOR2_X1 U3422 ( .A(n2724), .B(n2788), .ZN(n2727) );
  NOR2_X1 U3423 ( .A1(n2853), .A2(n4177), .ZN(n2725) );
  AOI21_X1 U3424 ( .B1(n4142), .B2(n2472), .A(n2725), .ZN(n2726) );
  NOR2_X1 U3425 ( .A1(n2727), .A2(n2726), .ZN(n3143) );
  AND2_X1 U3426 ( .A1(n2727), .A2(n2726), .ZN(n3144) );
  NAND2_X1 U3427 ( .A1(n2730), .A2(REG2_REG_22__SCAN_IN), .ZN(n2737) );
  INV_X1 U3428 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3714) );
  NAND2_X1 U3429 ( .A1(n2731), .A2(n3714), .ZN(n2732) );
  AND2_X1 U3430 ( .A1(n2739), .A2(n2732), .ZN(n4132) );
  NAND2_X1 U3431 ( .A1(n2780), .A2(n4132), .ZN(n2736) );
  NAND2_X1 U3432 ( .A1(n2043), .A2(REG0_REG_22__SCAN_IN), .ZN(n2735) );
  INV_X1 U3433 ( .A(REG1_REG_22__SCAN_IN), .ZN(n2733) );
  OR2_X1 U3434 ( .A1(n3786), .A2(n2733), .ZN(n2734) );
  NAND4_X1 U3435 ( .A1(n2737), .A2(n2736), .A3(n2735), .A4(n2734), .ZN(n4143)
         );
  NAND2_X1 U3436 ( .A1(n2041), .A2(DATAI_22_), .ZN(n4129) );
  OAI22_X1 U3437 ( .A1(n3636), .A2(n2853), .B1(n2397), .B2(n4129), .ZN(n2738)
         );
  XNOR2_X1 U3438 ( .A(n2738), .B(n2042), .ZN(n2750) );
  OAI22_X1 U3439 ( .A1(n3636), .A2(n2487), .B1(n2853), .B2(n4129), .ZN(n2749)
         );
  XNOR2_X1 U3440 ( .A(n2750), .B(n2749), .ZN(n3713) );
  NAND2_X1 U3441 ( .A1(n2739), .A2(n3635), .ZN(n2740) );
  AND2_X1 U3442 ( .A1(n2754), .A2(n2740), .ZN(n4117) );
  NAND2_X1 U3443 ( .A1(n2780), .A2(n4117), .ZN(n2744) );
  NAND2_X1 U3444 ( .A1(n2730), .A2(REG2_REG_23__SCAN_IN), .ZN(n2743) );
  NAND2_X1 U3445 ( .A1(n2043), .A2(REG0_REG_23__SCAN_IN), .ZN(n2742) );
  INV_X1 U3446 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4301) );
  OR2_X1 U3447 ( .A1(n3786), .A2(n4301), .ZN(n2741) );
  NAND2_X1 U3448 ( .A1(n4126), .A2(n2047), .ZN(n2746) );
  NAND2_X1 U3449 ( .A1(n3787), .A2(DATAI_23_), .ZN(n4115) );
  OR2_X1 U3450 ( .A1(n2397), .A2(n4115), .ZN(n2745) );
  NAND2_X1 U3451 ( .A1(n2746), .A2(n2745), .ZN(n2747) );
  XNOR2_X1 U3452 ( .A(n2747), .B(n2788), .ZN(n2763) );
  NOR2_X1 U3453 ( .A1(n2853), .A2(n4115), .ZN(n2748) );
  AOI21_X1 U3454 ( .B1(n4126), .B2(n2045), .A(n2748), .ZN(n2762) );
  XNOR2_X1 U3455 ( .A(n2763), .B(n2762), .ZN(n3632) );
  NOR2_X1 U3456 ( .A1(n2750), .A2(n2749), .ZN(n3633) );
  INV_X1 U3457 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3692) );
  AND2_X1 U34580 ( .A1(n2754), .A2(n3692), .ZN(n2755) );
  OR2_X1 U34590 ( .A1(n2755), .A2(n2769), .ZN(n4094) );
  INV_X1 U3460 ( .A(n3786), .ZN(n2756) );
  AOI22_X1 U3461 ( .A1(n2756), .A2(REG1_REG_24__SCAN_IN), .B1(n2391), .B2(
        REG2_REG_24__SCAN_IN), .ZN(n2758) );
  NAND2_X1 U3462 ( .A1(n2043), .A2(REG0_REG_24__SCAN_IN), .ZN(n2757) );
  NAND2_X1 U3463 ( .A1(n4110), .A2(n2048), .ZN(n2760) );
  NAND2_X1 U3464 ( .A1(n2041), .A2(DATAI_24_), .ZN(n4092) );
  OR2_X1 U3465 ( .A1(n2397), .A2(n4092), .ZN(n2759) );
  NAND2_X1 U3466 ( .A1(n2760), .A2(n2759), .ZN(n2761) );
  XNOR2_X1 U34670 ( .A(n2761), .B(n2042), .ZN(n2767) );
  INV_X1 U3468 ( .A(n2767), .ZN(n2765) );
  NOR2_X1 U34690 ( .A1(n2763), .A2(n2762), .ZN(n2768) );
  INV_X1 U3470 ( .A(n2768), .ZN(n2764) );
  INV_X1 U34710 ( .A(n4092), .ZN(n4085) );
  AOI22_X1 U3472 ( .A1(n4110), .A2(n2045), .B1(n2048), .B2(n4085), .ZN(n3690)
         );
  OAI21_X1 U34730 ( .B1(n3631), .B2(n2768), .A(n2767), .ZN(n3688) );
  NAND2_X1 U3474 ( .A1(n2769), .A2(REG3_REG_25__SCAN_IN), .ZN(n2778) );
  OR2_X1 U34750 ( .A1(n2769), .A2(REG3_REG_25__SCAN_IN), .ZN(n2770) );
  NAND2_X1 U3476 ( .A1(n2778), .A2(n2770), .ZN(n3668) );
  AOI22_X1 U34770 ( .A1(n2756), .A2(REG1_REG_25__SCAN_IN), .B1(n2730), .B2(
        REG2_REG_25__SCAN_IN), .ZN(n2772) );
  NAND2_X1 U3478 ( .A1(n2043), .A2(REG0_REG_25__SCAN_IN), .ZN(n2771) );
  NAND2_X1 U34790 ( .A1(n3787), .A2(DATAI_25_), .ZN(n4072) );
  NOR2_X1 U3480 ( .A1(n2397), .A2(n4072), .ZN(n2773) );
  AOI21_X1 U34810 ( .B1(n4086), .B2(n2047), .A(n2773), .ZN(n2774) );
  XNOR2_X1 U3482 ( .A(n2774), .B(n2814), .ZN(n2777) );
  NOR2_X1 U34830 ( .A1(n2853), .A2(n4072), .ZN(n2775) );
  AOI21_X1 U3484 ( .B1(n4086), .B2(n2045), .A(n2775), .ZN(n2776) );
  NAND2_X1 U34850 ( .A1(n2777), .A2(n2776), .ZN(n3664) );
  NOR2_X1 U3486 ( .A1(n2777), .A2(n2776), .ZN(n3665) );
  INV_X1 U34870 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3746) );
  NAND2_X1 U3488 ( .A1(n2778), .A2(n3746), .ZN(n2779) );
  NAND2_X1 U34890 ( .A1(n4059), .A2(n2780), .ZN(n2785) );
  INV_X1 U3490 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4289) );
  NAND2_X1 U34910 ( .A1(n2043), .A2(REG0_REG_26__SCAN_IN), .ZN(n2782) );
  NAND2_X1 U3492 ( .A1(n2730), .A2(REG2_REG_26__SCAN_IN), .ZN(n2781) );
  OAI211_X1 U34930 ( .C1(n3786), .C2(n4289), .A(n2782), .B(n2781), .ZN(n2783)
         );
  INV_X1 U3494 ( .A(n2783), .ZN(n2784) );
  NAND2_X1 U34950 ( .A1(n4069), .A2(n2048), .ZN(n2787) );
  NAND2_X1 U3496 ( .A1(n2041), .A2(DATAI_26_), .ZN(n4058) );
  OR2_X1 U34970 ( .A1(n2397), .A2(n4058), .ZN(n2786) );
  NAND2_X1 U3498 ( .A1(n2787), .A2(n2786), .ZN(n2789) );
  XNOR2_X1 U34990 ( .A(n2789), .B(n2788), .ZN(n2792) );
  NOR2_X1 U3500 ( .A1(n2853), .A2(n4058), .ZN(n2790) );
  AOI21_X1 U35010 ( .B1(n4069), .B2(n2472), .A(n2790), .ZN(n2791) );
  OR2_X1 U3502 ( .A1(n2792), .A2(n2791), .ZN(n3744) );
  INV_X1 U35030 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3611) );
  AND2_X1 U3504 ( .A1(n2793), .A2(n3611), .ZN(n2794) );
  INV_X1 U35050 ( .A(REG1_REG_27__SCAN_IN), .ZN(n2797) );
  NAND2_X1 U35060 ( .A1(n2391), .A2(REG2_REG_27__SCAN_IN), .ZN(n2796) );
  NAND2_X1 U35070 ( .A1(n2043), .A2(REG0_REG_27__SCAN_IN), .ZN(n2795) );
  OAI211_X1 U35080 ( .C1(n2797), .C2(n3786), .A(n2796), .B(n2795), .ZN(n2798)
         );
  INV_X1 U35090 ( .A(n2798), .ZN(n2799) );
  NAND2_X1 U35100 ( .A1(n4052), .A2(n2047), .ZN(n2801) );
  NAND2_X1 U35110 ( .A1(n3787), .A2(DATAI_27_), .ZN(n4038) );
  OR2_X1 U35120 ( .A1(n2397), .A2(n4038), .ZN(n2800) );
  NAND2_X1 U35130 ( .A1(n2801), .A2(n2800), .ZN(n2802) );
  XNOR2_X1 U35140 ( .A(n2802), .B(n2814), .ZN(n2841) );
  NOR2_X1 U35150 ( .A1(n2853), .A2(n4038), .ZN(n2803) );
  AOI21_X1 U35160 ( .B1(n4052), .B2(n2472), .A(n2803), .ZN(n2842) );
  XNOR2_X1 U35170 ( .A(n2841), .B(n2842), .ZN(n3608) );
  NOR2_X1 U35180 ( .A1(n2804), .A2(REG3_REG_28__SCAN_IN), .ZN(n2805) );
  INV_X1 U35190 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2808) );
  NAND2_X1 U35200 ( .A1(n2391), .A2(REG2_REG_28__SCAN_IN), .ZN(n2807) );
  NAND2_X1 U35210 ( .A1(n2043), .A2(REG0_REG_28__SCAN_IN), .ZN(n2806) );
  OAI211_X1 U35220 ( .C1(n2808), .C2(n3786), .A(n2807), .B(n2806), .ZN(n2809)
         );
  INV_X1 U35230 ( .A(n2809), .ZN(n2810) );
  NAND2_X1 U35240 ( .A1(n4036), .A2(n2045), .ZN(n2813) );
  NAND2_X1 U35250 ( .A1(n3787), .A2(DATAI_28_), .ZN(n3131) );
  OR2_X1 U35260 ( .A1(n2853), .A2(n3131), .ZN(n2812) );
  NAND2_X1 U35270 ( .A1(n2813), .A2(n2812), .ZN(n2815) );
  XNOR2_X1 U35280 ( .A(n2815), .B(n2042), .ZN(n2818) );
  INV_X1 U35290 ( .A(n3131), .ZN(n3584) );
  AOI22_X1 U35300 ( .A1(n4036), .A2(n2047), .B1(n2816), .B2(n3584), .ZN(n2817)
         );
  XNOR2_X1 U35310 ( .A(n2818), .B(n2817), .ZN(n2844) );
  INV_X1 U35320 ( .A(n2844), .ZN(n2847) );
  NAND2_X1 U35330 ( .A1(n3198), .A2(B_REG_SCAN_IN), .ZN(n2820) );
  INV_X1 U35340 ( .A(n2819), .ZN(n4393) );
  MUX2_X1 U35350 ( .A(n2820), .B(B_REG_SCAN_IN), .S(n4393), .Z(n2821) );
  INV_X1 U35360 ( .A(n4392), .ZN(n2832) );
  NAND2_X1 U35370 ( .A1(n2832), .A2(n2819), .ZN(n3205) );
  NOR4_X1 U35380 ( .A1(D_REG_17__SCAN_IN), .A2(D_REG_18__SCAN_IN), .A3(
        D_REG_19__SCAN_IN), .A4(D_REG_20__SCAN_IN), .ZN(n2825) );
  NOR4_X1 U35390 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_13__SCAN_IN), .A3(
        D_REG_14__SCAN_IN), .A4(D_REG_16__SCAN_IN), .ZN(n2824) );
  NOR4_X1 U35400 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2823) );
  NOR4_X1 U35410 ( .A1(D_REG_21__SCAN_IN), .A2(D_REG_22__SCAN_IN), .A3(
        D_REG_23__SCAN_IN), .A4(D_REG_25__SCAN_IN), .ZN(n2822) );
  AND4_X1 U35420 ( .A1(n2825), .A2(n2824), .A3(n2823), .A4(n2822), .ZN(n2831)
         );
  NOR2_X1 U35430 ( .A1(D_REG_24__SCAN_IN), .A2(D_REG_12__SCAN_IN), .ZN(n2829)
         );
  NOR4_X1 U35440 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_10__SCAN_IN), .A4(D_REG_2__SCAN_IN), .ZN(n2828) );
  NOR4_X1 U35450 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_8__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_11__SCAN_IN), .ZN(n2827) );
  NOR4_X1 U35460 ( .A1(D_REG_3__SCAN_IN), .A2(D_REG_4__SCAN_IN), .A3(
        D_REG_5__SCAN_IN), .A4(D_REG_6__SCAN_IN), .ZN(n2826) );
  AND4_X1 U35470 ( .A1(n2829), .A2(n2828), .A3(n2827), .A4(n2826), .ZN(n2830)
         );
  NAND2_X1 U35480 ( .A1(n2831), .A2(n2830), .ZN(n3121) );
  INV_X1 U35490 ( .A(D_REG_1__SCAN_IN), .ZN(n3203) );
  NOR2_X1 U35500 ( .A1(n3121), .A2(n3203), .ZN(n2833) );
  NAND2_X1 U35510 ( .A1(n2832), .A2(n3198), .ZN(n3201) );
  OAI21_X1 U35520 ( .B1(n3199), .B2(n2833), .A(n3201), .ZN(n2834) );
  INV_X1 U35530 ( .A(n2834), .ZN(n3311) );
  NAND2_X1 U35540 ( .A1(n3135), .A2(n3311), .ZN(n2860) );
  INV_X1 U35550 ( .A(n2860), .ZN(n2839) );
  INV_X1 U35560 ( .A(n2360), .ZN(n4396) );
  INV_X1 U35570 ( .A(n2836), .ZN(n4621) );
  NAND2_X1 U35580 ( .A1(n4394), .A2(n4395), .ZN(n3094) );
  OAI21_X1 U35590 ( .B1(n4621), .B2(n2707), .A(n3094), .ZN(n2837) );
  NOR2_X1 U35600 ( .A1(n3207), .A2(n2848), .ZN(n2838) );
  NAND3_X1 U35610 ( .A1(n2840), .A2(n2847), .A3(n4424), .ZN(n2875) );
  INV_X1 U35620 ( .A(n2841), .ZN(n2843) );
  OR2_X1 U35630 ( .A1(n2843), .A2(n2842), .ZN(n2845) );
  INV_X1 U35640 ( .A(n2845), .ZN(n2846) );
  NAND3_X1 U35650 ( .A1(n2847), .A2(n4424), .A3(n2846), .ZN(n2872) );
  INV_X1 U35660 ( .A(n3601), .ZN(n2870) );
  NAND2_X1 U35670 ( .A1(n2848), .A2(n4267), .ZN(n2849) );
  NAND2_X1 U35680 ( .A1(n2860), .A2(n2849), .ZN(n3284) );
  AOI21_X1 U35690 ( .B1(n2360), .B2(n2707), .A(n3094), .ZN(n3120) );
  INV_X1 U35700 ( .A(n3120), .ZN(n2850) );
  NAND4_X1 U35710 ( .A1(n3284), .A2(n3163), .A3(n3208), .A4(n2850), .ZN(n2851)
         );
  NAND2_X1 U35720 ( .A1(n2851), .A2(STATE_REG_SCAN_IN), .ZN(n2854) );
  INV_X1 U35730 ( .A(n2859), .ZN(n3932) );
  NAND2_X1 U35740 ( .A1(n2860), .A2(n3932), .ZN(n3285) );
  OR2_X1 U35750 ( .A1(n3207), .A2(n4267), .ZN(n2855) );
  OR2_X1 U35760 ( .A1(n2860), .A2(n2855), .ZN(n2857) );
  INV_X1 U35770 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2858) );
  OAI22_X1 U35780 ( .A1(n3762), .A2(n3131), .B1(STATE_REG_SCAN_IN), .B2(n2858), 
        .ZN(n2869) );
  INV_X1 U35790 ( .A(n4052), .ZN(n3748) );
  NOR2_X1 U35800 ( .A1(n2860), .A2(n2859), .ZN(n2867) );
  NAND2_X1 U35810 ( .A1(n2346), .A2(n2861), .ZN(n2862) );
  NAND2_X1 U3582 ( .A1(n2862), .A2(IR_REG_31__SCAN_IN), .ZN(n2863) );
  NAND2_X2 U3583 ( .A1(n2867), .A2(n4391), .ZN(n4414) );
  INV_X1 U3584 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2899) );
  NAND2_X1 U3585 ( .A1(n2730), .A2(REG2_REG_29__SCAN_IN), .ZN(n2865) );
  NAND2_X1 U3586 ( .A1(n2043), .A2(REG0_REG_29__SCAN_IN), .ZN(n2864) );
  OAI211_X1 U3587 ( .C1(n3786), .C2(n2899), .A(n2865), .B(n2864), .ZN(n2866)
         );
  AOI21_X1 U3588 ( .B1(n3594), .B2(n2389), .A(n2866), .ZN(n3792) );
  NAND2_X2 U3589 ( .A1(n2867), .A2(n3225), .ZN(n4413) );
  OAI22_X1 U3590 ( .A1(n3748), .A2(n4414), .B1(n3792), .B2(n4413), .ZN(n2868)
         );
  AOI211_X1 U3591 ( .C1(n2870), .C2(n3751), .A(n2869), .B(n2868), .ZN(n2871)
         );
  AOI21_X1 U3592 ( .B1(n2873), .B2(n2286), .A(n2285), .ZN(n2874) );
  NAND2_X1 U3593 ( .A1(n2875), .A2(n2874), .ZN(n3047) );
  INV_X1 U3594 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4348) );
  AOI22_X1 U3595 ( .A1(n4348), .A2(keyinput123), .B1(n2877), .B2(keyinput83), 
        .ZN(n2876) );
  OAI221_X1 U3596 ( .B1(n4348), .B2(keyinput123), .C1(n2877), .C2(keyinput83), 
        .A(n2876), .ZN(n2885) );
  INV_X1 U3597 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3016) );
  AOI22_X1 U3598 ( .A1(n4134), .A2(keyinput68), .B1(keyinput81), .B2(n3016), 
        .ZN(n2878) );
  OAI221_X1 U3599 ( .B1(n4134), .B2(keyinput68), .C1(n3016), .C2(keyinput81), 
        .A(n2878), .ZN(n2884) );
  INV_X1 U3600 ( .A(ADDR_REG_11__SCAN_IN), .ZN(n2880) );
  INV_X1 U3601 ( .A(ADDR_REG_16__SCAN_IN), .ZN(n2985) );
  AOI22_X1 U3602 ( .A1(n2880), .A2(keyinput64), .B1(keyinput124), .B2(n2985), 
        .ZN(n2879) );
  OAI221_X1 U3603 ( .B1(n2880), .B2(keyinput64), .C1(n2985), .C2(keyinput124), 
        .A(n2879), .ZN(n2883) );
  INV_X1 U3604 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n3222) );
  AOI22_X1 U3605 ( .A1(n2461), .A2(keyinput88), .B1(keyinput84), .B2(n3222), 
        .ZN(n2881) );
  OAI221_X1 U3606 ( .B1(n2461), .B2(keyinput88), .C1(n3222), .C2(keyinput84), 
        .A(n2881), .ZN(n2882) );
  NOR4_X1 U3607 ( .A1(n2885), .A2(n2884), .A3(n2883), .A4(n2882), .ZN(n3044)
         );
  INV_X1 U3608 ( .A(DATAI_0_), .ZN(n4662) );
  AOI22_X1 U3609 ( .A1(n3635), .A2(keyinput127), .B1(keyinput122), .B2(n4662), 
        .ZN(n2886) );
  OAI221_X1 U3610 ( .B1(n3635), .B2(keyinput127), .C1(n4662), .C2(keyinput122), 
        .A(n2886), .ZN(n2894) );
  INV_X1 U3611 ( .A(DATAI_9_), .ZN(n2888) );
  AOI22_X1 U3612 ( .A1(n2888), .A2(keyinput74), .B1(n4642), .B2(keyinput105), 
        .ZN(n2887) );
  OAI221_X1 U3613 ( .B1(n2888), .B2(keyinput74), .C1(n4642), .C2(keyinput105), 
        .A(n2887), .ZN(n2893) );
  INV_X1 U3614 ( .A(D_REG_12__SCAN_IN), .ZN(n4636) );
  INV_X1 U3615 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4377) );
  AOI22_X1 U3616 ( .A1(n4636), .A2(keyinput120), .B1(keyinput77), .B2(n4377), 
        .ZN(n2889) );
  OAI221_X1 U3617 ( .B1(n4636), .B2(keyinput120), .C1(n4377), .C2(keyinput77), 
        .A(n2889), .ZN(n2892) );
  INV_X1 U3618 ( .A(DATAI_6_), .ZN(n4658) );
  INV_X1 U3619 ( .A(D_REG_24__SCAN_IN), .ZN(n4635) );
  AOI22_X1 U3620 ( .A1(n4658), .A2(keyinput70), .B1(n4635), .B2(keyinput100), 
        .ZN(n2890) );
  OAI221_X1 U3621 ( .B1(n4658), .B2(keyinput70), .C1(n4635), .C2(keyinput100), 
        .A(n2890), .ZN(n2891) );
  NOR4_X1 U3622 ( .A1(n2894), .A2(n2893), .A3(n2892), .A4(n2891), .ZN(n2957)
         );
  OAI22_X1 U3623 ( .A1(REG0_REG_13__SCAN_IN), .A2(keyinput114), .B1(
        keyinput110), .B2(REG0_REG_18__SCAN_IN), .ZN(n2895) );
  AOI221_X1 U3624 ( .B1(REG0_REG_13__SCAN_IN), .B2(keyinput114), .C1(
        REG0_REG_18__SCAN_IN), .C2(keyinput110), .A(n2895), .ZN(n2903) );
  OAI22_X1 U3625 ( .A1(D_REG_21__SCAN_IN), .A2(keyinput71), .B1(keyinput89), 
        .B2(REG0_REG_0__SCAN_IN), .ZN(n2896) );
  AOI221_X1 U3626 ( .B1(D_REG_21__SCAN_IN), .B2(keyinput71), .C1(
        REG0_REG_0__SCAN_IN), .C2(keyinput89), .A(n2896), .ZN(n2902) );
  INV_X1 U3627 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3381) );
  INV_X1 U3628 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4278) );
  OAI22_X1 U3629 ( .A1(n3381), .A2(keyinput66), .B1(n4278), .B2(keyinput111), 
        .ZN(n2897) );
  AOI221_X1 U3630 ( .B1(n3381), .B2(keyinput66), .C1(keyinput111), .C2(n4278), 
        .A(n2897), .ZN(n2901) );
  OAI22_X1 U3631 ( .A1(n2899), .A2(keyinput107), .B1(keyinput76), .B2(
        IR_REG_9__SCAN_IN), .ZN(n2898) );
  AOI221_X1 U3632 ( .B1(n2899), .B2(keyinput107), .C1(IR_REG_9__SCAN_IN), .C2(
        keyinput76), .A(n2898), .ZN(n2900) );
  NAND4_X1 U3633 ( .A1(n2903), .A2(n2902), .A3(n2901), .A4(n2900), .ZN(n2922)
         );
  INV_X1 U3634 ( .A(REG2_REG_31__SCAN_IN), .ZN(n4433) );
  INV_X1 U3635 ( .A(ADDR_REG_17__SCAN_IN), .ZN(n3015) );
  AOI22_X1 U3636 ( .A1(n4433), .A2(keyinput78), .B1(keyinput73), .B2(n3015), 
        .ZN(n2904) );
  OAI221_X1 U3637 ( .B1(n4433), .B2(keyinput78), .C1(n3015), .C2(keyinput73), 
        .A(n2904), .ZN(n2905) );
  INV_X1 U3638 ( .A(n2905), .ZN(n2920) );
  XNOR2_X1 U3639 ( .A(IR_REG_0__SCAN_IN), .B(keyinput103), .ZN(n2909) );
  XNOR2_X1 U3640 ( .A(IR_REG_10__SCAN_IN), .B(keyinput112), .ZN(n2908) );
  XNOR2_X1 U3641 ( .A(IR_REG_1__SCAN_IN), .B(keyinput72), .ZN(n2907) );
  XNOR2_X1 U3642 ( .A(IR_REG_18__SCAN_IN), .B(keyinput75), .ZN(n2906) );
  NAND4_X1 U3643 ( .A1(n2909), .A2(n2908), .A3(n2907), .A4(n2906), .ZN(n2915)
         );
  XNOR2_X1 U3644 ( .A(IR_REG_11__SCAN_IN), .B(keyinput121), .ZN(n2913) );
  XNOR2_X1 U3645 ( .A(IR_REG_31__SCAN_IN), .B(keyinput101), .ZN(n2912) );
  XNOR2_X1 U3646 ( .A(IR_REG_27__SCAN_IN), .B(keyinput95), .ZN(n2911) );
  XNOR2_X1 U3647 ( .A(keyinput65), .B(REG0_REG_6__SCAN_IN), .ZN(n2910) );
  NAND4_X1 U3648 ( .A1(n2913), .A2(n2912), .A3(n2911), .A4(n2910), .ZN(n2914)
         );
  NOR2_X1 U3649 ( .A1(n2915), .A2(n2914), .ZN(n2919) );
  INV_X1 U3650 ( .A(DATAO_REG_9__SCAN_IN), .ZN(n3270) );
  AOI22_X1 U3651 ( .A1(n3270), .A2(keyinput92), .B1(n2858), .B2(keyinput117), 
        .ZN(n2916) );
  OAI221_X1 U3652 ( .B1(n3270), .B2(keyinput92), .C1(n2858), .C2(keyinput117), 
        .A(n2916), .ZN(n2917) );
  INV_X1 U3653 ( .A(n2917), .ZN(n2918) );
  NAND3_X1 U3654 ( .A1(n2920), .A2(n2919), .A3(n2918), .ZN(n2921) );
  NOR2_X1 U3655 ( .A1(n2922), .A2(n2921), .ZN(n2956) );
  OAI22_X1 U3656 ( .A1(REG3_REG_15__SCAN_IN), .A2(keyinput69), .B1(keyinput109), .B2(DATAO_REG_18__SCAN_IN), .ZN(n2923) );
  AOI221_X1 U3657 ( .B1(REG3_REG_15__SCAN_IN), .B2(keyinput69), .C1(
        DATAO_REG_18__SCAN_IN), .C2(keyinput109), .A(n2923), .ZN(n2930) );
  OAI22_X1 U3658 ( .A1(DATAO_REG_22__SCAN_IN), .A2(keyinput67), .B1(
        DATAO_REG_17__SCAN_IN), .B2(keyinput115), .ZN(n2924) );
  AOI221_X1 U3659 ( .B1(DATAO_REG_22__SCAN_IN), .B2(keyinput67), .C1(
        keyinput115), .C2(DATAO_REG_17__SCAN_IN), .A(n2924), .ZN(n2929) );
  OAI22_X1 U3660 ( .A1(ADDR_REG_5__SCAN_IN), .A2(keyinput97), .B1(
        DATAO_REG_6__SCAN_IN), .B2(keyinput102), .ZN(n2925) );
  AOI221_X1 U3661 ( .B1(ADDR_REG_5__SCAN_IN), .B2(keyinput97), .C1(keyinput102), .C2(DATAO_REG_6__SCAN_IN), .A(n2925), .ZN(n2928) );
  OAI22_X1 U3662 ( .A1(B_REG_SCAN_IN), .A2(keyinput126), .B1(
        DATAO_REG_29__SCAN_IN), .B2(keyinput86), .ZN(n2926) );
  AOI221_X1 U3663 ( .B1(B_REG_SCAN_IN), .B2(keyinput126), .C1(keyinput86), 
        .C2(DATAO_REG_29__SCAN_IN), .A(n2926), .ZN(n2927) );
  NAND4_X1 U3664 ( .A1(n2930), .A2(n2929), .A3(n2928), .A4(n2927), .ZN(n2935)
         );
  INV_X1 U3665 ( .A(D_REG_10__SCAN_IN), .ZN(n4637) );
  AOI22_X1 U3666 ( .A1(n4637), .A2(keyinput91), .B1(keyinput99), .B2(n3203), 
        .ZN(n2931) );
  OAI221_X1 U3667 ( .B1(n4637), .B2(keyinput91), .C1(n3203), .C2(keyinput99), 
        .A(n2931), .ZN(n2934) );
  INV_X1 U3668 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n3213) );
  INV_X1 U3669 ( .A(DATAO_REG_16__SCAN_IN), .ZN(n3217) );
  AOI22_X1 U3670 ( .A1(n3213), .A2(keyinput82), .B1(keyinput93), .B2(n3217), 
        .ZN(n2932) );
  OAI221_X1 U3671 ( .B1(n3213), .B2(keyinput82), .C1(n3217), .C2(keyinput93), 
        .A(n2932), .ZN(n2933) );
  NOR3_X1 U3672 ( .A1(n2935), .A2(n2934), .A3(n2933), .ZN(n2955) );
  OAI22_X1 U3673 ( .A1(REG0_REG_27__SCAN_IN), .A2(keyinput118), .B1(
        keyinput125), .B2(REG2_REG_8__SCAN_IN), .ZN(n2936) );
  AOI221_X1 U3674 ( .B1(REG0_REG_27__SCAN_IN), .B2(keyinput118), .C1(
        REG2_REG_8__SCAN_IN), .C2(keyinput125), .A(n2936), .ZN(n2943) );
  OAI22_X1 U3675 ( .A1(REG2_REG_3__SCAN_IN), .A2(keyinput113), .B1(
        REG2_REG_15__SCAN_IN), .B2(keyinput106), .ZN(n2937) );
  AOI221_X1 U3676 ( .B1(REG2_REG_3__SCAN_IN), .B2(keyinput113), .C1(
        keyinput106), .C2(REG2_REG_15__SCAN_IN), .A(n2937), .ZN(n2942) );
  OAI22_X1 U3677 ( .A1(REG1_REG_22__SCAN_IN), .A2(keyinput108), .B1(
        REG1_REG_10__SCAN_IN), .B2(keyinput80), .ZN(n2938) );
  AOI221_X1 U3678 ( .B1(REG1_REG_22__SCAN_IN), .B2(keyinput108), .C1(
        keyinput80), .C2(REG1_REG_10__SCAN_IN), .A(n2938), .ZN(n2941) );
  OAI22_X1 U3679 ( .A1(REG0_REG_23__SCAN_IN), .A2(keyinput104), .B1(keyinput94), .B2(REG0_REG_21__SCAN_IN), .ZN(n2939) );
  AOI221_X1 U3680 ( .B1(REG0_REG_23__SCAN_IN), .B2(keyinput104), .C1(
        REG0_REG_21__SCAN_IN), .C2(keyinput94), .A(n2939), .ZN(n2940) );
  NAND4_X1 U3681 ( .A1(n2943), .A2(n2942), .A3(n2941), .A4(n2940), .ZN(n2953)
         );
  OAI22_X1 U3682 ( .A1(IR_REG_8__SCAN_IN), .A2(keyinput116), .B1(keyinput85), 
        .B2(REG3_REG_8__SCAN_IN), .ZN(n2944) );
  AOI221_X1 U3683 ( .B1(IR_REG_8__SCAN_IN), .B2(keyinput116), .C1(
        REG3_REG_8__SCAN_IN), .C2(keyinput85), .A(n2944), .ZN(n2951) );
  OAI22_X1 U3684 ( .A1(REG3_REG_5__SCAN_IN), .A2(keyinput96), .B1(keyinput79), 
        .B2(REG3_REG_16__SCAN_IN), .ZN(n2945) );
  AOI221_X1 U3685 ( .B1(REG3_REG_5__SCAN_IN), .B2(keyinput96), .C1(
        REG3_REG_16__SCAN_IN), .C2(keyinput79), .A(n2945), .ZN(n2950) );
  OAI22_X1 U3686 ( .A1(DATAI_3_), .A2(keyinput98), .B1(keyinput119), .B2(
        DATAI_31_), .ZN(n2946) );
  AOI221_X1 U3687 ( .B1(DATAI_3_), .B2(keyinput98), .C1(DATAI_31_), .C2(
        keyinput119), .A(n2946), .ZN(n2949) );
  OAI22_X1 U3688 ( .A1(IR_REG_3__SCAN_IN), .A2(keyinput87), .B1(DATAI_8_), 
        .B2(keyinput90), .ZN(n2947) );
  AOI221_X1 U3689 ( .B1(IR_REG_3__SCAN_IN), .B2(keyinput87), .C1(keyinput90), 
        .C2(DATAI_8_), .A(n2947), .ZN(n2948) );
  NAND4_X1 U3690 ( .A1(n2951), .A2(n2950), .A3(n2949), .A4(n2948), .ZN(n2952)
         );
  NOR2_X1 U3691 ( .A1(n2953), .A2(n2952), .ZN(n2954) );
  AND4_X1 U3692 ( .A1(n2957), .A2(n2956), .A3(n2955), .A4(n2954), .ZN(n3043)
         );
  AOI22_X1 U3693 ( .A1(DATAO_REG_18__SCAN_IN), .A2(keyinput45), .B1(
        IR_REG_31__SCAN_IN), .B2(keyinput37), .ZN(n2958) );
  OAI221_X1 U3694 ( .B1(DATAO_REG_18__SCAN_IN), .B2(keyinput45), .C1(
        IR_REG_31__SCAN_IN), .C2(keyinput37), .A(n2958), .ZN(n2965) );
  AOI22_X1 U3695 ( .A1(REG2_REG_3__SCAN_IN), .A2(keyinput49), .B1(
        REG3_REG_8__SCAN_IN), .B2(keyinput21), .ZN(n2959) );
  OAI221_X1 U3696 ( .B1(REG2_REG_3__SCAN_IN), .B2(keyinput49), .C1(
        REG3_REG_8__SCAN_IN), .C2(keyinput21), .A(n2959), .ZN(n2964) );
  AOI22_X1 U3697 ( .A1(REG0_REG_6__SCAN_IN), .A2(keyinput1), .B1(
        REG0_REG_19__SCAN_IN), .B2(keyinput13), .ZN(n2960) );
  OAI221_X1 U3698 ( .B1(REG0_REG_6__SCAN_IN), .B2(keyinput1), .C1(
        REG0_REG_19__SCAN_IN), .C2(keyinput13), .A(n2960), .ZN(n2963) );
  AOI22_X1 U3699 ( .A1(DATAI_17_), .A2(keyinput41), .B1(REG3_REG_28__SCAN_IN), 
        .B2(keyinput53), .ZN(n2961) );
  OAI221_X1 U3700 ( .B1(DATAI_17_), .B2(keyinput41), .C1(REG3_REG_28__SCAN_IN), 
        .C2(keyinput53), .A(n2961), .ZN(n2962) );
  NOR4_X1 U3701 ( .A1(n2965), .A2(n2964), .A3(n2963), .A4(n2962), .ZN(n3009)
         );
  AOI22_X1 U3702 ( .A1(REG0_REG_18__SCAN_IN), .A2(keyinput46), .B1(
        B_REG_SCAN_IN), .B2(keyinput62), .ZN(n2966) );
  OAI221_X1 U3703 ( .B1(REG0_REG_18__SCAN_IN), .B2(keyinput46), .C1(
        B_REG_SCAN_IN), .C2(keyinput62), .A(n2966), .ZN(n2973) );
  AOI22_X1 U3704 ( .A1(DATAO_REG_6__SCAN_IN), .A2(keyinput38), .B1(
        REG0_REG_13__SCAN_IN), .B2(keyinput50), .ZN(n2967) );
  OAI221_X1 U3705 ( .B1(DATAO_REG_6__SCAN_IN), .B2(keyinput38), .C1(
        REG0_REG_13__SCAN_IN), .C2(keyinput50), .A(n2967), .ZN(n2972) );
  AOI22_X1 U3706 ( .A1(DATAI_9_), .A2(keyinput10), .B1(REG0_REG_21__SCAN_IN), 
        .B2(keyinput30), .ZN(n2968) );
  OAI221_X1 U3707 ( .B1(DATAI_9_), .B2(keyinput10), .C1(REG0_REG_21__SCAN_IN), 
        .C2(keyinput30), .A(n2968), .ZN(n2971) );
  AOI22_X1 U3708 ( .A1(ADDR_REG_11__SCAN_IN), .A2(keyinput0), .B1(
        REG2_REG_7__SCAN_IN), .B2(keyinput2), .ZN(n2969) );
  OAI221_X1 U3709 ( .B1(ADDR_REG_11__SCAN_IN), .B2(keyinput0), .C1(
        REG2_REG_7__SCAN_IN), .C2(keyinput2), .A(n2969), .ZN(n2970) );
  NOR4_X1 U3710 ( .A1(n2973), .A2(n2972), .A3(n2971), .A4(n2970), .ZN(n3008)
         );
  AOI22_X1 U3711 ( .A1(REG2_REG_8__SCAN_IN), .A2(keyinput61), .B1(
        REG1_REG_22__SCAN_IN), .B2(keyinput44), .ZN(n2974) );
  OAI221_X1 U3712 ( .B1(REG2_REG_8__SCAN_IN), .B2(keyinput61), .C1(
        REG1_REG_22__SCAN_IN), .C2(keyinput44), .A(n2974), .ZN(n2981) );
  AOI22_X1 U3713 ( .A1(REG1_REG_10__SCAN_IN), .A2(keyinput16), .B1(
        REG3_REG_15__SCAN_IN), .B2(keyinput5), .ZN(n2975) );
  OAI221_X1 U3714 ( .B1(REG1_REG_10__SCAN_IN), .B2(keyinput16), .C1(
        REG3_REG_15__SCAN_IN), .C2(keyinput5), .A(n2975), .ZN(n2980) );
  AOI22_X1 U3715 ( .A1(REG3_REG_5__SCAN_IN), .A2(keyinput32), .B1(
        IR_REG_8__SCAN_IN), .B2(keyinput52), .ZN(n2976) );
  OAI221_X1 U3716 ( .B1(REG3_REG_5__SCAN_IN), .B2(keyinput32), .C1(
        IR_REG_8__SCAN_IN), .C2(keyinput52), .A(n2976), .ZN(n2979) );
  AOI22_X1 U3717 ( .A1(IR_REG_11__SCAN_IN), .A2(keyinput57), .B1(
        IR_REG_1__SCAN_IN), .B2(keyinput8), .ZN(n2977) );
  OAI221_X1 U3718 ( .B1(IR_REG_11__SCAN_IN), .B2(keyinput57), .C1(
        IR_REG_1__SCAN_IN), .C2(keyinput8), .A(n2977), .ZN(n2978) );
  NOR4_X1 U3719 ( .A1(n2981), .A2(n2980), .A3(n2979), .A4(n2978), .ZN(n3007)
         );
  INV_X1 U3720 ( .A(DATAI_3_), .ZN(n2983) );
  AOI22_X1 U3721 ( .A1(n2983), .A2(keyinput34), .B1(n3203), .B2(keyinput35), 
        .ZN(n2982) );
  OAI221_X1 U3722 ( .B1(n2983), .B2(keyinput34), .C1(n3203), .C2(keyinput35), 
        .A(n2982), .ZN(n2987) );
  AOI22_X1 U3723 ( .A1(n4635), .A2(keyinput36), .B1(keyinput60), .B2(n2985), 
        .ZN(n2984) );
  OAI221_X1 U3724 ( .B1(n4635), .B2(keyinput36), .C1(n2985), .C2(keyinput60), 
        .A(n2984), .ZN(n2986) );
  NOR2_X1 U3725 ( .A1(n2987), .A2(n2986), .ZN(n3005) );
  INV_X1 U3726 ( .A(DATAI_8_), .ZN(n4655) );
  INV_X1 U3727 ( .A(DATAO_REG_29__SCAN_IN), .ZN(n3220) );
  AOI22_X1 U3728 ( .A1(n4655), .A2(keyinput26), .B1(keyinput22), .B2(n3220), 
        .ZN(n2988) );
  OAI221_X1 U3729 ( .B1(n4655), .B2(keyinput26), .C1(n3220), .C2(keyinput22), 
        .A(n2988), .ZN(n2991) );
  INV_X1 U3730 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4411) );
  AOI22_X1 U3731 ( .A1(n4433), .A2(keyinput14), .B1(n4411), .B2(keyinput15), 
        .ZN(n2989) );
  OAI221_X1 U3732 ( .B1(n4433), .B2(keyinput14), .C1(n4411), .C2(keyinput15), 
        .A(n2989), .ZN(n2990) );
  NOR2_X1 U3733 ( .A1(n2991), .A2(n2990), .ZN(n3004) );
  AOI22_X1 U3734 ( .A1(n3222), .A2(keyinput20), .B1(n2461), .B2(keyinput24), 
        .ZN(n2992) );
  OAI221_X1 U3735 ( .B1(n3222), .B2(keyinput20), .C1(n2461), .C2(keyinput24), 
        .A(n2992), .ZN(n2994) );
  XNOR2_X1 U3736 ( .A(n3213), .B(keyinput18), .ZN(n2993) );
  NOR2_X1 U3737 ( .A1(n2994), .A2(n2993), .ZN(n3003) );
  INV_X1 U3738 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4366) );
  AOI22_X1 U3739 ( .A1(n3270), .A2(keyinput28), .B1(n4366), .B2(keyinput40), 
        .ZN(n2995) );
  OAI221_X1 U3740 ( .B1(n3270), .B2(keyinput28), .C1(n4366), .C2(keyinput40), 
        .A(n2995), .ZN(n3001) );
  XNOR2_X1 U3741 ( .A(n2996), .B(keyinput11), .ZN(n2999) );
  XNOR2_X1 U3742 ( .A(IR_REG_9__SCAN_IN), .B(keyinput12), .ZN(n2998) );
  XNOR2_X1 U3743 ( .A(IR_REG_3__SCAN_IN), .B(keyinput23), .ZN(n2997) );
  NAND3_X1 U3744 ( .A1(n2999), .A2(n2998), .A3(n2997), .ZN(n3000) );
  NOR2_X1 U3745 ( .A1(n3001), .A2(n3000), .ZN(n3002) );
  AND4_X1 U3746 ( .A1(n3005), .A2(n3004), .A3(n3003), .A4(n3002), .ZN(n3006)
         );
  NAND4_X1 U3747 ( .A1(n3009), .A2(n3008), .A3(n3007), .A4(n3006), .ZN(n3042)
         );
  INV_X1 U3748 ( .A(ADDR_REG_5__SCAN_IN), .ZN(n3011) );
  AOI22_X1 U3749 ( .A1(n4134), .A2(keyinput4), .B1(keyinput33), .B2(n3011), 
        .ZN(n3010) );
  OAI221_X1 U3750 ( .B1(n4134), .B2(keyinput4), .C1(n3011), .C2(keyinput33), 
        .A(n3010), .ZN(n3020) );
  INV_X1 U3751 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n3215) );
  AOI22_X1 U3752 ( .A1(n4658), .A2(keyinput6), .B1(keyinput3), .B2(n3215), 
        .ZN(n3012) );
  OAI221_X1 U3753 ( .B1(n4658), .B2(keyinput6), .C1(n3215), .C2(keyinput3), 
        .A(n3012), .ZN(n3019) );
  INV_X1 U3754 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4666) );
  AOI22_X1 U3755 ( .A1(n4666), .A2(keyinput25), .B1(keyinput29), .B2(n3217), 
        .ZN(n3013) );
  OAI221_X1 U3756 ( .B1(n4666), .B2(keyinput25), .C1(n3217), .C2(keyinput29), 
        .A(n3013), .ZN(n3018) );
  AOI22_X1 U3757 ( .A1(n3016), .A2(keyinput17), .B1(keyinput9), .B2(n3015), 
        .ZN(n3014) );
  OAI221_X1 U3758 ( .B1(n3016), .B2(keyinput17), .C1(n3015), .C2(keyinput9), 
        .A(n3014), .ZN(n3017) );
  NOR4_X1 U3759 ( .A1(n3020), .A2(n3019), .A3(n3018), .A4(n3017), .ZN(n3040)
         );
  AOI22_X1 U3760 ( .A1(n3635), .A2(keyinput63), .B1(keyinput58), .B2(n4662), 
        .ZN(n3021) );
  OAI221_X1 U3761 ( .B1(n3635), .B2(keyinput63), .C1(n4662), .C2(keyinput58), 
        .A(n3021), .ZN(n3029) );
  AOI22_X1 U3762 ( .A1(n4636), .A2(keyinput56), .B1(n2296), .B2(keyinput48), 
        .ZN(n3022) );
  OAI221_X1 U3763 ( .B1(n4636), .B2(keyinput56), .C1(n2296), .C2(keyinput48), 
        .A(n3022), .ZN(n3028) );
  AOI22_X1 U3764 ( .A1(n4257), .A2(keyinput42), .B1(n2377), .B2(keyinput39), 
        .ZN(n3023) );
  OAI221_X1 U3765 ( .B1(n4257), .B2(keyinput42), .C1(n2377), .C2(keyinput39), 
        .A(n3023), .ZN(n3027) );
  INV_X1 U3766 ( .A(DATAI_31_), .ZN(n3196) );
  INV_X1 U3767 ( .A(REG0_REG_27__SCAN_IN), .ZN(n3025) );
  AOI22_X1 U3768 ( .A1(n3196), .A2(keyinput55), .B1(n3025), .B2(keyinput54), 
        .ZN(n3024) );
  OAI221_X1 U3769 ( .B1(n3196), .B2(keyinput55), .C1(n3025), .C2(keyinput54), 
        .A(n3024), .ZN(n3026) );
  NOR4_X1 U3770 ( .A1(n3029), .A2(n3028), .A3(n3027), .A4(n3026), .ZN(n3039)
         );
  AOI22_X1 U3771 ( .A1(IR_REG_27__SCAN_IN), .A2(keyinput31), .B1(
        D_REG_21__SCAN_IN), .B2(keyinput7), .ZN(n3030) );
  OAI221_X1 U3772 ( .B1(IR_REG_27__SCAN_IN), .B2(keyinput31), .C1(
        D_REG_21__SCAN_IN), .C2(keyinput7), .A(n3030), .ZN(n3037) );
  AOI22_X1 U3773 ( .A1(DATAO_REG_17__SCAN_IN), .A2(keyinput51), .B1(
        REG1_REG_30__SCAN_IN), .B2(keyinput47), .ZN(n3031) );
  OAI221_X1 U3774 ( .B1(DATAO_REG_17__SCAN_IN), .B2(keyinput51), .C1(
        REG1_REG_30__SCAN_IN), .C2(keyinput47), .A(n3031), .ZN(n3036) );
  AOI22_X1 U3775 ( .A1(REG0_REG_30__SCAN_IN), .A2(keyinput59), .B1(
        REG1_REG_29__SCAN_IN), .B2(keyinput43), .ZN(n3032) );
  OAI221_X1 U3776 ( .B1(REG0_REG_30__SCAN_IN), .B2(keyinput59), .C1(
        REG1_REG_29__SCAN_IN), .C2(keyinput43), .A(n3032), .ZN(n3035) );
  AOI22_X1 U3777 ( .A1(REG1_REG_21__SCAN_IN), .A2(keyinput19), .B1(
        D_REG_10__SCAN_IN), .B2(keyinput27), .ZN(n3033) );
  OAI221_X1 U3778 ( .B1(REG1_REG_21__SCAN_IN), .B2(keyinput19), .C1(
        D_REG_10__SCAN_IN), .C2(keyinput27), .A(n3033), .ZN(n3034) );
  NOR4_X1 U3779 ( .A1(n3037), .A2(n3036), .A3(n3035), .A4(n3034), .ZN(n3038)
         );
  NAND3_X1 U3780 ( .A1(n3040), .A2(n3039), .A3(n3038), .ZN(n3041) );
  AOI211_X1 U3781 ( .C1(n3044), .C2(n3043), .A(n3042), .B(n3041), .ZN(n3045)
         );
  INV_X1 U3782 ( .A(n3045), .ZN(n3046) );
  XNOR2_X1 U3783 ( .A(n3047), .B(n3046), .ZN(U3217) );
  INV_X1 U3784 ( .A(n3939), .ZN(n4412) );
  NAND2_X1 U3785 ( .A1(n3049), .A2(n3128), .ZN(n3852) );
  NAND2_X1 U3786 ( .A1(n3095), .A2(n4606), .ZN(n4605) );
  INV_X1 U3787 ( .A(n3128), .ZN(n4613) );
  NAND2_X1 U3788 ( .A1(n3049), .A2(n4613), .ZN(n3051) );
  NAND2_X1 U3789 ( .A1(n3054), .A2(n3455), .ZN(n3857) );
  NAND2_X1 U3790 ( .A1(n3447), .A2(n3450), .ZN(n3446) );
  OR2_X1 U3791 ( .A1(n3054), .A2(n3052), .ZN(n3055) );
  NOR2_X1 U3792 ( .A1(n3948), .A2(n3860), .ZN(n3056) );
  INV_X1 U3793 ( .A(n3860), .ZN(n3407) );
  OR2_X1 U3794 ( .A1(n3947), .A2(n3322), .ZN(n3862) );
  NAND2_X1 U3795 ( .A1(n3947), .A2(n3322), .ZN(n3865) );
  NAND2_X1 U3796 ( .A1(n3862), .A2(n3865), .ZN(n3812) );
  NAND2_X1 U3797 ( .A1(n3301), .A2(n3812), .ZN(n3058) );
  INV_X1 U3798 ( .A(n3322), .ZN(n3303) );
  NAND2_X1 U3799 ( .A1(n3947), .A2(n3303), .ZN(n3057) );
  NAND2_X1 U3800 ( .A1(n3058), .A2(n3057), .ZN(n3493) );
  AND2_X1 U3801 ( .A1(n3946), .A2(n3488), .ZN(n3059) );
  NOR2_X1 U3802 ( .A1(n3945), .A2(n3364), .ZN(n3061) );
  NAND2_X1 U3803 ( .A1(n3945), .A2(n3364), .ZN(n3060) );
  OR2_X1 U3804 ( .A1(n3944), .A2(n3869), .ZN(n3098) );
  NAND2_X1 U3805 ( .A1(n3944), .A2(n3869), .ZN(n3880) );
  NAND2_X1 U3806 ( .A1(n3098), .A2(n3880), .ZN(n3813) );
  INV_X1 U3807 ( .A(n3869), .ZN(n3062) );
  AND2_X1 U3808 ( .A1(n3943), .A2(n3100), .ZN(n3063) );
  OAI22_X1 U3809 ( .A1(n3421), .A2(n3063), .B1(n3100), .B2(n3943), .ZN(n3508)
         );
  NOR2_X1 U3810 ( .A1(n3473), .A2(n3509), .ZN(n3064) );
  NAND2_X1 U3811 ( .A1(n3473), .A2(n3509), .ZN(n3065) );
  NAND2_X1 U3812 ( .A1(n3066), .A2(n3065), .ZN(n3470) );
  AND2_X1 U3813 ( .A1(n4580), .A2(n3481), .ZN(n3068) );
  OR2_X1 U3814 ( .A1(n4580), .A2(n3481), .ZN(n3067) );
  OAI21_X1 U3815 ( .B1(n3470), .B2(n3068), .A(n3067), .ZN(n4577) );
  OR2_X1 U3816 ( .A1(n3942), .A2(n3129), .ZN(n3851) );
  NAND2_X1 U3817 ( .A1(n3942), .A2(n3129), .ZN(n3892) );
  NAND2_X1 U3818 ( .A1(n3851), .A2(n3892), .ZN(n4578) );
  NAND2_X1 U3819 ( .A1(n4577), .A2(n4578), .ZN(n3070) );
  INV_X1 U3820 ( .A(n3129), .ZN(n4590) );
  OR2_X1 U3821 ( .A1(n3942), .A2(n4590), .ZN(n3069) );
  NAND2_X1 U3822 ( .A1(n3070), .A2(n3069), .ZN(n3521) );
  NOR2_X1 U3823 ( .A1(n4582), .A2(n3103), .ZN(n3071) );
  NOR2_X1 U3824 ( .A1(n3521), .A2(n3071), .ZN(n3072) );
  NOR2_X1 U3825 ( .A1(n3941), .A2(n3544), .ZN(n3534) );
  OR2_X1 U3826 ( .A1(n4252), .A2(n3625), .ZN(n3767) );
  NAND2_X1 U3827 ( .A1(n4252), .A2(n3625), .ZN(n3768) );
  AND2_X1 U3828 ( .A1(n3940), .A2(n4254), .ZN(n3073) );
  INV_X1 U3829 ( .A(n3073), .ZN(n3075) );
  OR2_X1 U3830 ( .A1(n4252), .A2(n3556), .ZN(n4241) );
  OAI22_X1 U3831 ( .A1(n3073), .A2(n4241), .B1(n4254), .B2(n3940), .ZN(n3074)
         );
  OR2_X1 U3832 ( .A1(n4224), .A2(n3576), .ZN(n3901) );
  NAND2_X1 U3833 ( .A1(n4224), .A2(n3576), .ZN(n3900) );
  NAND2_X1 U3834 ( .A1(n3901), .A2(n3900), .ZN(n3572) );
  OR2_X1 U3835 ( .A1(n4191), .A2(n4213), .ZN(n3106) );
  NAND2_X1 U3836 ( .A1(n4191), .A2(n4213), .ZN(n4184) );
  NAND2_X1 U3837 ( .A1(n3106), .A2(n4184), .ZN(n4211) );
  INV_X1 U3838 ( .A(n4213), .ZN(n4204) );
  NAND2_X1 U3839 ( .A1(n4205), .A2(n4195), .ZN(n3078) );
  INV_X1 U3840 ( .A(n4142), .ZN(n4189) );
  NAND2_X1 U3841 ( .A1(n4189), .A2(n4177), .ZN(n3080) );
  INV_X1 U3842 ( .A(n4177), .ZN(n3079) );
  INV_X1 U3843 ( .A(n4151), .ZN(n3081) );
  XNOR2_X1 U3844 ( .A(n4143), .B(n4129), .ZN(n4124) );
  NAND2_X1 U3845 ( .A1(n4100), .A2(n2066), .ZN(n3083) );
  NAND2_X1 U3846 ( .A1(n4126), .A2(n3806), .ZN(n3082) );
  NAND2_X1 U3847 ( .A1(n3083), .A2(n3082), .ZN(n4080) );
  NOR2_X1 U3848 ( .A1(n4067), .A2(n4092), .ZN(n3085) );
  NAND2_X1 U3849 ( .A1(n4067), .A2(n4092), .ZN(n3084) );
  INV_X1 U3850 ( .A(n4072), .ZN(n3086) );
  INV_X1 U3851 ( .A(n4058), .ZN(n4051) );
  NAND2_X1 U3852 ( .A1(n4029), .A2(n4058), .ZN(n3087) );
  NAND2_X1 U3853 ( .A1(n3088), .A2(n3087), .ZN(n4028) );
  INV_X1 U3854 ( .A(n4038), .ZN(n3089) );
  NOR2_X1 U3855 ( .A1(n4052), .A2(n3089), .ZN(n3091) );
  NAND2_X1 U3856 ( .A1(n4052), .A2(n3089), .ZN(n3090) );
  OR2_X1 U3857 ( .A1(n4036), .A2(n3131), .ZN(n3782) );
  NAND2_X1 U3858 ( .A1(n4036), .A2(n3131), .ZN(n3794) );
  NAND2_X1 U3859 ( .A1(n3782), .A2(n3794), .ZN(n3807) );
  XNOR2_X1 U3860 ( .A(n3585), .B(n3807), .ZN(n3607) );
  XNOR2_X1 U3861 ( .A(n3092), .B(n4394), .ZN(n3093) );
  NAND2_X1 U3862 ( .A1(n3225), .A2(n3209), .ZN(n4627) );
  OAI22_X1 U3863 ( .A1(n3792), .A2(n4627), .B1(n3131), .B2(n4267), .ZN(n3119)
         );
  INV_X1 U3864 ( .A(n4607), .ZN(n4601) );
  INV_X1 U3865 ( .A(n3450), .ZN(n3818) );
  XNOR2_X1 U3866 ( .A(n3948), .B(n3860), .ZN(n3843) );
  NAND2_X1 U3867 ( .A1(n3096), .A2(n3843), .ZN(n3410) );
  OR2_X1 U3868 ( .A1(n3948), .A2(n3407), .ZN(n3861) );
  INV_X1 U3869 ( .A(n3862), .ZN(n3097) );
  INV_X1 U3870 ( .A(n3488), .ZN(n3496) );
  AND2_X1 U3871 ( .A1(n3946), .A2(n3496), .ZN(n3486) );
  OR2_X1 U3872 ( .A1(n3946), .A2(n3496), .ZN(n3881) );
  INV_X1 U3873 ( .A(n3364), .ZN(n3358) );
  NAND2_X1 U3874 ( .A1(n3945), .A2(n3358), .ZN(n3883) );
  OR2_X1 U3875 ( .A1(n3945), .A2(n3358), .ZN(n3867) );
  INV_X1 U3876 ( .A(n3098), .ZN(n3099) );
  OR2_X1 U3877 ( .A1(n3943), .A2(n3428), .ZN(n3874) );
  NAND2_X1 U3878 ( .A1(n3943), .A2(n3428), .ZN(n3884) );
  AND2_X1 U3879 ( .A1(n3473), .A2(n2117), .ZN(n3878) );
  OR2_X1 U3880 ( .A1(n3473), .A2(n2117), .ZN(n3875) );
  INV_X1 U3881 ( .A(n3481), .ZN(n3476) );
  NAND2_X1 U3882 ( .A1(n4580), .A2(n3476), .ZN(n3893) );
  NAND2_X1 U3883 ( .A1(n3472), .A2(n3893), .ZN(n3101) );
  OR2_X1 U3884 ( .A1(n4580), .A2(n3476), .ZN(n3887) );
  NAND2_X1 U3885 ( .A1(n3101), .A2(n3887), .ZN(n4579) );
  NAND2_X1 U3886 ( .A1(n4579), .A2(n3892), .ZN(n3102) );
  NAND2_X1 U3887 ( .A1(n3102), .A2(n3851), .ZN(n3537) );
  NAND2_X1 U3888 ( .A1(n4582), .A2(n3658), .ZN(n3535) );
  INV_X1 U3889 ( .A(n3544), .ZN(n3705) );
  NAND2_X1 U3890 ( .A1(n3941), .A2(n3705), .ZN(n3104) );
  NOR2_X1 U3891 ( .A1(n4582), .A2(n3658), .ZN(n3536) );
  NOR2_X1 U3892 ( .A1(n3941), .A2(n3705), .ZN(n3105) );
  AOI21_X1 U3893 ( .B1(n3847), .B2(n3536), .A(n3105), .ZN(n3850) );
  INV_X1 U3894 ( .A(n4254), .ZN(n4244) );
  OR2_X1 U3895 ( .A1(n3940), .A2(n4244), .ZN(n3770) );
  NAND2_X1 U3896 ( .A1(n3940), .A2(n4244), .ZN(n3769) );
  NAND2_X1 U3897 ( .A1(n3770), .A2(n3769), .ZN(n4248) );
  INV_X1 U3898 ( .A(n3572), .ZN(n3819) );
  NAND2_X1 U3899 ( .A1(n4205), .A2(n4188), .ZN(n3828) );
  NAND2_X1 U3900 ( .A1(n3939), .A2(n4222), .ZN(n3903) );
  NAND3_X1 U3901 ( .A1(n4164), .A2(n3900), .A3(n3903), .ZN(n3772) );
  NOR2_X1 U3902 ( .A1(n3939), .A2(n4222), .ZN(n4161) );
  INV_X1 U3903 ( .A(n3106), .ZN(n4185) );
  NAND2_X1 U3904 ( .A1(n4164), .A2(n4185), .ZN(n3107) );
  OR2_X1 U3905 ( .A1(n4205), .A2(n4188), .ZN(n3829) );
  NAND2_X1 U3906 ( .A1(n3107), .A2(n3829), .ZN(n4165) );
  NOR2_X1 U3907 ( .A1(n4142), .A2(n4177), .ZN(n3108) );
  OR2_X1 U3908 ( .A1(n4165), .A2(n3108), .ZN(n3109) );
  AOI21_X1 U3909 ( .B1(n4164), .B2(n4161), .A(n3109), .ZN(n3906) );
  NAND2_X1 U3910 ( .A1(n4142), .A2(n4177), .ZN(n4102) );
  OR2_X1 U3911 ( .A1(n4171), .A2(n4151), .ZN(n4104) );
  OR2_X1 U3912 ( .A1(n4143), .A2(n4129), .ZN(n4106) );
  NAND2_X1 U3913 ( .A1(n4104), .A2(n4106), .ZN(n3908) );
  AND2_X1 U3914 ( .A1(n4171), .A2(n4151), .ZN(n3905) );
  NAND2_X1 U3915 ( .A1(n4126), .A2(n4115), .ZN(n3111) );
  NAND2_X1 U3916 ( .A1(n4143), .A2(n4129), .ZN(n3110) );
  NAND2_X1 U3917 ( .A1(n3111), .A2(n3110), .ZN(n3911) );
  AOI21_X1 U3918 ( .B1(n3905), .B2(n4106), .A(n3911), .ZN(n3776) );
  INV_X1 U3919 ( .A(n3776), .ZN(n3112) );
  NOR2_X1 U3920 ( .A1(n3113), .A2(n3112), .ZN(n4082) );
  NOR2_X1 U3921 ( .A1(n4110), .A2(n4092), .ZN(n3826) );
  NOR2_X1 U3922 ( .A1(n4126), .A2(n4115), .ZN(n4081) );
  NOR2_X1 U3923 ( .A1(n3826), .A2(n4081), .ZN(n3910) );
  INV_X1 U3924 ( .A(n3910), .ZN(n3114) );
  NAND2_X1 U3925 ( .A1(n4110), .A2(n4092), .ZN(n3778) );
  OAI21_X1 U3926 ( .B1(n4082), .B2(n3114), .A(n3778), .ZN(n4066) );
  AND2_X1 U3927 ( .A1(n4086), .A2(n4072), .ZN(n3834) );
  NOR2_X1 U3928 ( .A1(n4066), .A2(n3834), .ZN(n4048) );
  OR2_X1 U3929 ( .A1(n4086), .A2(n4072), .ZN(n4046) );
  OAI21_X1 U3930 ( .B1(n4069), .B2(n4058), .A(n4046), .ZN(n3916) );
  AND2_X1 U3931 ( .A1(n4069), .A2(n4058), .ZN(n3919) );
  INV_X1 U3932 ( .A(n3919), .ZN(n3115) );
  OR2_X1 U3933 ( .A1(n4052), .A2(n4038), .ZN(n3781) );
  NAND2_X1 U3934 ( .A1(n4052), .A2(n4038), .ZN(n3913) );
  NAND2_X1 U3935 ( .A1(n3781), .A2(n3913), .ZN(n4031) );
  NAND2_X1 U3936 ( .A1(n4396), .A2(n4395), .ZN(n3804) );
  NAND2_X1 U3937 ( .A1(n4397), .A2(n4394), .ZN(n3116) );
  NOR2_X1 U3938 ( .A1(n3117), .A2(n4585), .ZN(n3118) );
  OAI21_X1 U3939 ( .B1(n3199), .B2(D_REG_1__SCAN_IN), .A(n3201), .ZN(n3126) );
  INV_X1 U3940 ( .A(n3199), .ZN(n3122) );
  NAND2_X1 U3941 ( .A1(n3122), .A2(n3121), .ZN(n3125) );
  NAND2_X1 U3942 ( .A1(n4716), .A2(n3123), .ZN(n3124) );
  NAND4_X1 U3943 ( .A1(n3310), .A2(n3126), .A3(n3125), .A4(n3124), .ZN(n3136)
         );
  MUX2_X1 U3944 ( .A(REG1_REG_28__SCAN_IN), .B(n3137), .S(n4735), .Z(n3127) );
  INV_X1 U3945 ( .A(n3127), .ZN(n3134) );
  NOR2_X1 U3946 ( .A1(n4674), .A2(n3860), .ZN(n3415) );
  NAND2_X1 U3947 ( .A1(n3415), .A2(n3322), .ZN(n3494) );
  NAND2_X1 U3948 ( .A1(n4213), .A2(n4188), .ZN(n3130) );
  INV_X1 U3949 ( .A(n4129), .ZN(n4136) );
  INV_X1 U3950 ( .A(n4037), .ZN(n3132) );
  OAI21_X1 U3951 ( .B1(n3132), .B2(n3131), .A(n3588), .ZN(n3599) );
  NAND2_X1 U3952 ( .A1(n3134), .A2(n3133), .ZN(U3546) );
  NAND2_X1 U3953 ( .A1(n4375), .A2(n4715), .ZN(n4384) );
  NAND2_X1 U3954 ( .A1(n3139), .A2(n3138), .ZN(U3514) );
  INV_X1 U3955 ( .A(n3144), .ZN(n3140) );
  NAND2_X1 U3956 ( .A1(n3141), .A2(n3140), .ZN(n3146) );
  OAI21_X1 U3957 ( .B1(n3144), .B2(n3143), .A(n3142), .ZN(n3145) );
  AOI21_X1 U3958 ( .B1(n3146), .B2(n3145), .A(n3753), .ZN(n3152) );
  NOR2_X1 U3959 ( .A1(n4429), .A2(n3147), .ZN(n3151) );
  INV_X1 U3960 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3148) );
  OAI22_X1 U3961 ( .A1(n3762), .A2(n4177), .B1(STATE_REG_SCAN_IN), .B2(n3148), 
        .ZN(n3150) );
  INV_X1 U3962 ( .A(n4171), .ZN(n3715) );
  OAI22_X1 U3963 ( .A1(n3738), .A2(n4414), .B1(n4413), .B2(n3715), .ZN(n3149)
         );
  XNOR2_X1 U3964 ( .A(n3153), .B(n2158), .ZN(n3154) );
  XNOR2_X1 U3965 ( .A(n3155), .B(n3154), .ZN(n3156) );
  NOR2_X1 U3966 ( .A1(n3156), .A2(n3753), .ZN(n3162) );
  INV_X1 U3967 ( .A(n3157), .ZN(n4152) );
  NOR2_X1 U3968 ( .A1(n4429), .A2(n4152), .ZN(n3161) );
  INV_X1 U3969 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3158) );
  OAI22_X1 U3970 ( .A1(n3762), .A2(n4151), .B1(STATE_REG_SCAN_IN), .B2(n3158), 
        .ZN(n3160) );
  OAI22_X1 U3971 ( .A1(n4189), .A2(n4414), .B1(n4413), .B2(n3636), .ZN(n3159)
         );
  INV_X1 U3972 ( .A(n3164), .ZN(n3169) );
  AOI21_X1 U3973 ( .B1(n3168), .B2(n3166), .A(n3165), .ZN(n3167) );
  AOI21_X1 U3974 ( .B1(n3169), .B2(n3168), .A(n3167), .ZN(n3170) );
  NOR2_X1 U3975 ( .A1(n3170), .A2(n3753), .ZN(n3175) );
  NOR2_X1 U3976 ( .A1(n4429), .A2(n3423), .ZN(n3174) );
  INV_X1 U3977 ( .A(REG3_REG_8__SCAN_IN), .ZN(n3171) );
  OAI22_X1 U3978 ( .A1(n3762), .A2(n3428), .B1(STATE_REG_SCAN_IN), .B2(n3171), 
        .ZN(n3173) );
  INV_X1 U3979 ( .A(n3473), .ZN(n3429) );
  INV_X1 U3980 ( .A(n3944), .ZN(n3873) );
  OAI22_X1 U3981 ( .A1(n3429), .A2(n4413), .B1(n4414), .B2(n3873), .ZN(n3172)
         );
  OR4_X1 U3982 ( .A1(n3175), .A2(n3174), .A3(n3173), .A4(n3172), .ZN(U3218) );
  AOI211_X1 U3983 ( .C1(n3177), .C2(n3176), .A(n3753), .B(n2080), .ZN(n3183)
         );
  INV_X1 U3984 ( .A(n3178), .ZN(n3380) );
  NOR2_X1 U3985 ( .A1(n4429), .A2(n3380), .ZN(n3182) );
  AND2_X1 U3986 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n4482) );
  INV_X1 U3987 ( .A(n4482), .ZN(n3179) );
  OAI21_X1 U3988 ( .B1(n3762), .B2(n3869), .A(n3179), .ZN(n3181) );
  INV_X1 U3989 ( .A(n3945), .ZN(n3350) );
  INV_X1 U3990 ( .A(n3943), .ZN(n3505) );
  OAI22_X1 U3991 ( .A1(n3350), .A2(n4414), .B1(n4413), .B2(n3505), .ZN(n3180)
         );
  OR4_X1 U3992 ( .A1(n3183), .A2(n3182), .A3(n3181), .A4(n3180), .ZN(U3210) );
  INV_X1 U3993 ( .A(n3184), .ZN(n3185) );
  AOI211_X1 U3994 ( .C1(n3187), .C2(n3186), .A(n3753), .B(n3185), .ZN(n3192)
         );
  INV_X1 U3995 ( .A(n3188), .ZN(n3482) );
  NOR2_X1 U3996 ( .A1(n4429), .A2(n3482), .ZN(n3191) );
  NAND2_X1 U3997 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4499) );
  OAI21_X1 U3998 ( .B1(n3762), .B2(n3476), .A(n4499), .ZN(n3190) );
  INV_X1 U3999 ( .A(n3942), .ZN(n3656) );
  OAI22_X1 U4000 ( .A1(n3429), .A2(n4414), .B1(n4413), .B2(n3656), .ZN(n3189)
         );
  OR4_X1 U4001 ( .A1(n3192), .A2(n3191), .A3(n3190), .A4(n3189), .ZN(U3214) );
  OR4_X1 U4002 ( .A1(n3194), .A2(IR_REG_30__SCAN_IN), .A3(n3193), .A4(U3149), 
        .ZN(n3195) );
  OAI21_X1 U4003 ( .B1(STATE_REG_SCAN_IN), .B2(n3196), .A(n3195), .ZN(U3321)
         );
  NAND2_X1 U4004 ( .A1(U3149), .A2(DATAI_25_), .ZN(n3197) );
  OAI21_X1 U4005 ( .B1(n3198), .B2(U3149), .A(n3197), .ZN(U3327) );
  INV_X1 U4006 ( .A(n3207), .ZN(n3200) );
  INV_X1 U4007 ( .A(n3201), .ZN(n3202) );
  AOI22_X1 U4008 ( .A1(n4639), .A2(n3203), .B1(n3202), .B2(n4640), .ZN(U3459)
         );
  INV_X1 U4009 ( .A(n4639), .ZN(n4638) );
  OAI22_X1 U4010 ( .A1(n4638), .A2(D_REG_0__SCAN_IN), .B1(n3205), .B2(n3204), 
        .ZN(n3206) );
  INV_X1 U4011 ( .A(n3206), .ZN(U3458) );
  OR2_X1 U4012 ( .A1(n3208), .A2(U3149), .ZN(n3935) );
  NAND2_X1 U4013 ( .A1(n3207), .A2(n3935), .ZN(n3224) );
  NAND2_X1 U4014 ( .A1(n3209), .A2(n3208), .ZN(n3210) );
  AND2_X1 U4015 ( .A1(n2041), .A2(n3210), .ZN(n3223) );
  INV_X1 U4016 ( .A(n3223), .ZN(n3211) );
  NOR2_X1 U4017 ( .A1(n4563), .A2(U4043), .ZN(U3148) );
  NAND2_X1 U4018 ( .A1(n4252), .A2(U4043), .ZN(n3212) );
  OAI21_X1 U4019 ( .B1(n3213), .B2(U4043), .A(n3212), .ZN(U3564) );
  NAND2_X1 U4020 ( .A1(n4143), .A2(U4043), .ZN(n3214) );
  OAI21_X1 U4021 ( .B1(U4043), .B2(n3215), .A(n3214), .ZN(U3572) );
  NAND2_X1 U4022 ( .A1(n4224), .A2(U4043), .ZN(n3216) );
  OAI21_X1 U4023 ( .B1(U4043), .B2(n3217), .A(n3216), .ZN(U3566) );
  INV_X1 U4024 ( .A(n3792), .ZN(n3218) );
  NAND2_X1 U4025 ( .A1(n3218), .A2(U4043), .ZN(n3219) );
  OAI21_X1 U4026 ( .B1(U4043), .B2(n3220), .A(n3219), .ZN(U3579) );
  NAND2_X1 U4027 ( .A1(n4171), .A2(U4043), .ZN(n3221) );
  OAI21_X1 U4028 ( .B1(U4043), .B2(n3222), .A(n3221), .ZN(U3571) );
  INV_X1 U4029 ( .A(n4536), .ZN(n4576) );
  INV_X1 U4030 ( .A(n4399), .ZN(n3268) );
  AOI22_X1 U4031 ( .A1(REG2_REG_7__SCAN_IN), .A2(n4478), .B1(n4657), .B2(n3381), .ZN(n4486) );
  INV_X1 U4032 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3499) );
  AOI22_X1 U4033 ( .A1(n4660), .A2(REG2_REG_5__SCAN_IN), .B1(n3499), .B2(n4464), .ZN(n4461) );
  INV_X1 U4034 ( .A(REG2_REG_2__SCAN_IN), .ZN(n3972) );
  MUX2_X1 U4035 ( .A(n3972), .B(REG2_REG_2__SCAN_IN), .S(n3971), .Z(n3228) );
  INV_X1 U4036 ( .A(REG2_REG_1__SCAN_IN), .ZN(n3226) );
  MUX2_X1 U4037 ( .A(n3226), .B(REG2_REG_1__SCAN_IN), .S(n3952), .Z(n3949) );
  AND2_X1 U4038 ( .A1(REG2_REG_0__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n3961)
         );
  NAND2_X1 U4039 ( .A1(n3949), .A2(n3961), .ZN(n3974) );
  OR2_X1 U4040 ( .A1(n3952), .A2(n3226), .ZN(n3973) );
  NAND2_X1 U4041 ( .A1(n3974), .A2(n3973), .ZN(n3227) );
  INV_X1 U4042 ( .A(n3971), .ZN(n4400) );
  NAND2_X1 U40430 ( .A1(n4400), .A2(REG2_REG_2__SCAN_IN), .ZN(n3229) );
  NAND2_X1 U4044 ( .A1(n3230), .A2(n4406), .ZN(n3231) );
  NAND2_X1 U4045 ( .A1(n3231), .A2(n4404), .ZN(n3232) );
  INV_X1 U4046 ( .A(n3253), .ZN(n4444) );
  XNOR2_X1 U4047 ( .A(n3232), .B(n4444), .ZN(n4445) );
  INV_X1 U4048 ( .A(REG2_REG_4__SCAN_IN), .ZN(n3234) );
  INV_X1 U4049 ( .A(n3232), .ZN(n3233) );
  NAND2_X1 U4050 ( .A1(n4473), .A2(n3235), .ZN(n3236) );
  NAND2_X1 U4051 ( .A1(REG2_REG_6__SCAN_IN), .A2(n4472), .ZN(n4471) );
  NAND2_X1 U4052 ( .A1(n3259), .A2(n3237), .ZN(n3238) );
  NAND2_X1 U4053 ( .A1(REG2_REG_8__SCAN_IN), .A2(n4494), .ZN(n4493) );
  NAND2_X1 U4054 ( .A1(n3238), .A2(n4493), .ZN(n3243) );
  INV_X1 U4055 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3239) );
  MUX2_X1 U4056 ( .A(n3239), .B(REG2_REG_9__SCAN_IN), .S(n4399), .Z(n3240) );
  INV_X1 U4057 ( .A(n3240), .ZN(n3242) );
  XNOR2_X1 U4058 ( .A(n3241), .B(IR_REG_27__SCAN_IN), .ZN(n4438) );
  AND2_X1 U4059 ( .A1(n4391), .A2(n4438), .ZN(n3931) );
  NAND2_X1 U4060 ( .A1(n3242), .A2(n3243), .ZN(n3386) );
  OAI211_X1 U4061 ( .C1(n3243), .C2(n3242), .A(n4571), .B(n3386), .ZN(n3267)
         );
  INV_X1 U4062 ( .A(REG3_REG_9__SCAN_IN), .ZN(n3244) );
  NOR2_X1 U4063 ( .A1(STATE_REG_SCAN_IN), .A2(n3244), .ZN(n3439) );
  INV_X1 U4064 ( .A(n4473), .ZN(n4659) );
  AOI22_X1 U4065 ( .A1(n4660), .A2(REG1_REG_5__SCAN_IN), .B1(n2461), .B2(n4464), .ZN(n4458) );
  MUX2_X1 U4066 ( .A(n3245), .B(REG1_REG_2__SCAN_IN), .S(n3971), .Z(n3248) );
  AND2_X1 U4067 ( .A1(REG1_REG_0__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n3951)
         );
  OR2_X1 U4068 ( .A1(n3952), .A2(n3246), .ZN(n3964) );
  NAND2_X1 U4069 ( .A1(n3965), .A2(n3964), .ZN(n3247) );
  NAND2_X1 U4070 ( .A1(n3248), .A2(n3247), .ZN(n3968) );
  NAND2_X1 U4071 ( .A1(n4400), .A2(REG1_REG_2__SCAN_IN), .ZN(n3249) );
  NAND2_X1 U4072 ( .A1(n3968), .A2(n3249), .ZN(n3250) );
  NAND2_X1 U4073 ( .A1(n3250), .A2(n4406), .ZN(n3251) );
  INV_X1 U4074 ( .A(n3252), .ZN(n3254) );
  NAND2_X1 U4075 ( .A1(n4458), .A2(n4457), .ZN(n4456) );
  NAND2_X1 U4076 ( .A1(n4473), .A2(n3256), .ZN(n3257) );
  NOR2_X1 U4077 ( .A1(n2179), .A2(n3258), .ZN(n3260) );
  NAND2_X1 U4078 ( .A1(n4399), .A2(REG1_REG_9__SCAN_IN), .ZN(n3394) );
  OR2_X1 U4079 ( .A1(n4399), .A2(REG1_REG_9__SCAN_IN), .ZN(n3261) );
  NAND2_X1 U4080 ( .A1(n3394), .A2(n3261), .ZN(n3263) );
  INV_X1 U4081 ( .A(n3395), .ZN(n3262) );
  INV_X1 U4082 ( .A(n4438), .ZN(n3960) );
  AOI211_X1 U4083 ( .C1(n3264), .C2(n3263), .A(n3262), .B(n4540), .ZN(n3265)
         );
  AOI211_X1 U4084 ( .C1(n4563), .C2(ADDR_REG_9__SCAN_IN), .A(n3439), .B(n3265), 
        .ZN(n3266) );
  OAI211_X1 U4085 ( .C1(n4576), .C2(n3268), .A(n3267), .B(n3266), .ZN(U3249)
         );
  NAND2_X1 U4086 ( .A1(n3473), .A2(U4043), .ZN(n3269) );
  OAI21_X1 U4087 ( .B1(U4043), .B2(n3270), .A(n3269), .ZN(U3559) );
  OAI21_X1 U4088 ( .B1(n3273), .B2(n3272), .A(n3271), .ZN(n3274) );
  NAND2_X1 U4089 ( .A1(n3274), .A2(n4424), .ZN(n3279) );
  INV_X1 U4090 ( .A(n3947), .ZN(n3490) );
  OAI22_X1 U4091 ( .A1(n3053), .A2(n4414), .B1(n4413), .B2(n3490), .ZN(n3277)
         );
  NOR2_X1 U4092 ( .A1(STATE_REG_SCAN_IN), .A2(n2426), .ZN(n4401) );
  INV_X1 U4093 ( .A(n4401), .ZN(n3275) );
  OAI21_X1 U4094 ( .B1(n3762), .B2(n3407), .A(n3275), .ZN(n3276) );
  NOR2_X1 U4095 ( .A1(n3277), .A2(n3276), .ZN(n3278) );
  OAI211_X1 U4096 ( .C1(REG3_REG_3__SCAN_IN), .C2(n4429), .A(n3279), .B(n3278), 
        .ZN(U3215) );
  INV_X1 U4097 ( .A(n3280), .ZN(n3281) );
  AOI21_X1 U4098 ( .B1(n3283), .B2(n3282), .A(n3281), .ZN(n3288) );
  INV_X1 U4099 ( .A(n4413), .ZN(n3296) );
  INV_X1 U4100 ( .A(n3762), .ZN(n4417) );
  AOI22_X1 U4101 ( .A1(n3296), .A2(n3948), .B1(n4417), .B2(n3052), .ZN(n3287)
         );
  INV_X1 U4102 ( .A(n4414), .ZN(n3290) );
  NAND3_X1 U4103 ( .A1(n3285), .A2(n3284), .A3(n3310), .ZN(n3297) );
  AOI22_X1 U4104 ( .A1(n3290), .A2(n3049), .B1(REG3_REG_2__SCAN_IN), .B2(n3297), .ZN(n3286) );
  OAI211_X1 U4105 ( .C1(n3288), .C2(n3753), .A(n3287), .B(n3286), .ZN(U3234)
         );
  AOI22_X1 U4106 ( .A1(n3296), .A2(n3054), .B1(n4417), .B2(n4613), .ZN(n3292)
         );
  AOI22_X1 U4107 ( .A1(n3290), .A2(n3050), .B1(REG3_REG_1__SCAN_IN), .B2(n3297), .ZN(n3291) );
  OAI211_X1 U4108 ( .C1(n3293), .C2(n3753), .A(n3292), .B(n3291), .ZN(U3219)
         );
  XOR2_X1 U4109 ( .A(n3295), .B(n3294), .Z(n3958) );
  INV_X1 U4110 ( .A(n3958), .ZN(n3300) );
  AOI22_X1 U4111 ( .A1(n3296), .A2(n3049), .B1(n4417), .B2(n4612), .ZN(n3299)
         );
  NAND2_X1 U4112 ( .A1(n3297), .A2(REG3_REG_0__SCAN_IN), .ZN(n3298) );
  OAI211_X1 U4113 ( .C1(n3300), .C2(n3753), .A(n3299), .B(n3298), .ZN(U3229)
         );
  OAI211_X1 U4114 ( .C1(n3415), .C2(n3322), .A(n3494), .B(n4715), .ZN(n4685)
         );
  NOR2_X1 U4115 ( .A1(n4685), .A2(n4397), .ZN(n3308) );
  XNOR2_X1 U4116 ( .A(n3301), .B(n3812), .ZN(n3313) );
  XOR2_X1 U4117 ( .A(n3812), .B(n3302), .Z(n3306) );
  INV_X1 U4118 ( .A(n4603), .ZN(n4207) );
  AOI22_X1 U4119 ( .A1(n3946), .A2(n4581), .B1(n3303), .B2(n4602), .ZN(n3304)
         );
  OAI21_X1 U4120 ( .B1(n3859), .B2(n4207), .A(n3304), .ZN(n3305) );
  AOI21_X1 U4121 ( .B1(n3306), .B2(n4624), .A(n3305), .ZN(n3307) );
  OAI21_X1 U4122 ( .B1(n3313), .B2(n4608), .A(n3307), .ZN(n4686) );
  AOI211_X1 U4123 ( .C1(n4629), .C2(n3317), .A(n3308), .B(n4686), .ZN(n3316)
         );
  NAND3_X1 U4124 ( .A1(n3311), .A2(n3310), .A3(n3309), .ZN(n3312) );
  INV_X1 U4125 ( .A(n3313), .ZN(n4688) );
  OR2_X1 U4126 ( .A1(n3092), .A2(n2707), .ZN(n3375) );
  INV_X1 U4127 ( .A(n3375), .ZN(n3314) );
  AOI22_X1 U4128 ( .A1(n4688), .A2(n4630), .B1(REG2_REG_4__SCAN_IN), .B2(n4634), .ZN(n3315) );
  OAI21_X1 U4129 ( .B1(n3316), .B2(n4634), .A(n3315), .ZN(U3286) );
  INV_X1 U4130 ( .A(n3317), .ZN(n3327) );
  AND2_X1 U4131 ( .A1(n3271), .A2(n3318), .ZN(n3320) );
  OAI211_X1 U4132 ( .C1(n3320), .C2(n3319), .A(n4424), .B(n3347), .ZN(n3326)
         );
  INV_X1 U4133 ( .A(n3946), .ZN(n3336) );
  OAI22_X1 U4134 ( .A1(n3336), .A2(n4413), .B1(n4414), .B2(n3859), .ZN(n3324)
         );
  AND2_X1 U4135 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n4449) );
  INV_X1 U4136 ( .A(n4449), .ZN(n3321) );
  OAI21_X1 U4137 ( .B1(n3762), .B2(n3322), .A(n3321), .ZN(n3323) );
  NOR2_X1 U4138 ( .A1(n3324), .A2(n3323), .ZN(n3325) );
  OAI211_X1 U4139 ( .C1(n4429), .C2(n3327), .A(n3326), .B(n3325), .ZN(U3227)
         );
  INV_X1 U4140 ( .A(n4593), .ZN(n3343) );
  NAND2_X1 U4141 ( .A1(n3347), .A2(n3328), .ZN(n3330) );
  AND2_X1 U4142 ( .A1(n3330), .A2(n3329), .ZN(n3334) );
  NAND2_X1 U4143 ( .A1(n3332), .A2(n3331), .ZN(n3333) );
  XNOR2_X1 U4144 ( .A(n3334), .B(n3333), .ZN(n3335) );
  NAND2_X1 U4145 ( .A1(n3335), .A2(n4424), .ZN(n3342) );
  OAI22_X1 U4146 ( .A1(n3336), .A2(n4414), .B1(n4413), .B2(n3873), .ZN(n3340)
         );
  NOR2_X1 U4147 ( .A1(STATE_REG_SCAN_IN), .A2(n3337), .ZN(n4468) );
  INV_X1 U4148 ( .A(n4468), .ZN(n3338) );
  OAI21_X1 U4149 ( .B1(n3762), .B2(n3358), .A(n3338), .ZN(n3339) );
  NOR2_X1 U4150 ( .A1(n3340), .A2(n3339), .ZN(n3341) );
  OAI211_X1 U4151 ( .C1(n4429), .C2(n3343), .A(n3342), .B(n3341), .ZN(U3236)
         );
  INV_X1 U4152 ( .A(n3344), .ZN(n3498) );
  NAND2_X1 U4153 ( .A1(n3347), .A2(n3346), .ZN(n3348) );
  XOR2_X1 U4154 ( .A(n3345), .B(n3348), .Z(n3349) );
  NAND2_X1 U4155 ( .A1(n3349), .A2(n4424), .ZN(n3355) );
  OAI22_X1 U4156 ( .A1(n3490), .A2(n4414), .B1(n4413), .B2(n3350), .ZN(n3353)
         );
  AND2_X1 U4157 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n4466) );
  INV_X1 U4158 ( .A(n4466), .ZN(n3351) );
  OAI21_X1 U4159 ( .B1(n3762), .B2(n3496), .A(n3351), .ZN(n3352) );
  NOR2_X1 U4160 ( .A1(n3353), .A2(n3352), .ZN(n3354) );
  OAI211_X1 U4161 ( .C1(n4429), .C2(n3498), .A(n3355), .B(n3354), .ZN(U3224)
         );
  NAND2_X1 U4162 ( .A1(n3867), .A2(n3883), .ZN(n3814) );
  XNOR2_X1 U4163 ( .A(n3356), .B(n3814), .ZN(n4595) );
  INV_X1 U4164 ( .A(n4595), .ZN(n3363) );
  INV_X1 U4165 ( .A(n4608), .ZN(n4625) );
  XNOR2_X1 U4166 ( .A(n3357), .B(n3814), .ZN(n3361) );
  OAI22_X1 U4167 ( .A1(n3873), .A2(n4627), .B1(n4267), .B2(n3358), .ZN(n3359)
         );
  AOI21_X1 U4168 ( .B1(n4603), .B2(n3946), .A(n3359), .ZN(n3360) );
  OAI21_X1 U4169 ( .B1(n3361), .B2(n4585), .A(n3360), .ZN(n3362) );
  AOI21_X1 U4170 ( .B1(n4625), .B2(n4595), .A(n3362), .ZN(n4598) );
  OAI21_X1 U4171 ( .B1(n3363), .B2(n4679), .A(n4598), .ZN(n3367) );
  INV_X1 U4172 ( .A(n3367), .ZN(n3366) );
  AOI21_X1 U4173 ( .B1(n3364), .B2(n3495), .A(n3377), .ZN(n4594) );
  INV_X1 U4174 ( .A(n4384), .ZN(n4344) );
  AOI22_X1 U4175 ( .A1(n4594), .A2(n4344), .B1(REG0_REG_6__SCAN_IN), .B2(n4720), .ZN(n3365) );
  OAI21_X1 U4176 ( .B1(n3366), .B2(n4720), .A(n3365), .ZN(U3479) );
  NAND2_X1 U4177 ( .A1(n3367), .A2(n4735), .ZN(n3369) );
  INV_X1 U4178 ( .A(n4328), .ZN(n4264) );
  NAND2_X1 U4179 ( .A1(n4594), .A2(n4264), .ZN(n3368) );
  OAI211_X1 U4180 ( .C1(n4735), .C2(n2477), .A(n3369), .B(n3368), .ZN(U3524)
         );
  XNOR2_X1 U4181 ( .A(n3370), .B(n3813), .ZN(n3373) );
  OAI22_X1 U4182 ( .A1(n3505), .A2(n4627), .B1(n4267), .B2(n3869), .ZN(n3371)
         );
  AOI21_X1 U4183 ( .B1(n4603), .B2(n3945), .A(n3371), .ZN(n3372) );
  OAI21_X1 U4184 ( .B1(n3373), .B2(n4585), .A(n3372), .ZN(n4695) );
  INV_X1 U4185 ( .A(n4695), .ZN(n3385) );
  XOR2_X1 U4186 ( .A(n3374), .B(n3813), .Z(n4697) );
  NAND2_X1 U4187 ( .A1(n4608), .A2(n3375), .ZN(n3376) );
  NAND2_X1 U4188 ( .A1(n4697), .A2(n4237), .ZN(n3384) );
  OAI21_X1 U4189 ( .B1(n3377), .B2(n3869), .A(n4715), .ZN(n3378) );
  NOR2_X1 U4190 ( .A1(n3378), .A2(n3422), .ZN(n4696) );
  OAI22_X1 U4191 ( .A1(n3379), .A2(n3381), .B1(n3380), .B2(n4255), .ZN(n3382)
         );
  AOI21_X1 U4192 ( .B1(n4696), .B2(n4215), .A(n3382), .ZN(n3383) );
  OAI211_X1 U4193 ( .C1(n3385), .C2(n4634), .A(n3384), .B(n3383), .ZN(U3283)
         );
  NAND2_X1 U4194 ( .A1(n4399), .A2(REG2_REG_9__SCAN_IN), .ZN(n3387) );
  NAND2_X1 U4195 ( .A1(n3387), .A2(n3386), .ZN(n3388) );
  NAND2_X1 U4196 ( .A1(n3396), .A2(n3388), .ZN(n3389) );
  INV_X1 U4197 ( .A(n3396), .ZN(n4654) );
  XNOR2_X1 U4198 ( .A(n3388), .B(n4654), .ZN(n4503) );
  NAND2_X1 U4199 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4503), .ZN(n4502) );
  NAND2_X1 U4200 ( .A1(n3389), .A2(n4502), .ZN(n3392) );
  INV_X1 U4201 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3390) );
  MUX2_X1 U4202 ( .A(n3390), .B(REG2_REG_11__SCAN_IN), .S(n3992), .Z(n3391) );
  NAND2_X1 U4203 ( .A1(n3392), .A2(n3391), .ZN(n3982) );
  OAI211_X1 U4204 ( .C1(n3392), .C2(n3391), .A(n3982), .B(n4571), .ZN(n3405)
         );
  NOR2_X1 U4205 ( .A1(STATE_REG_SCAN_IN), .A2(n3393), .ZN(n3728) );
  NOR2_X1 U4206 ( .A1(n3397), .A2(n4654), .ZN(n3398) );
  MUX2_X1 U4207 ( .A(REG1_REG_11__SCAN_IN), .B(n3399), .S(n3992), .Z(n3401) );
  INV_X1 U4208 ( .A(n3994), .ZN(n3400) );
  AOI211_X1 U4209 ( .C1(n3402), .C2(n3401), .A(n3400), .B(n4540), .ZN(n3403)
         );
  AOI211_X1 U4210 ( .C1(n4563), .C2(ADDR_REG_11__SCAN_IN), .A(n3728), .B(n3403), .ZN(n3404) );
  OAI211_X1 U4211 ( .C1(n4576), .C2(n3992), .A(n3405), .B(n3404), .ZN(U3251)
         );
  XNOR2_X1 U4212 ( .A(n3406), .B(n3843), .ZN(n4680) );
  INV_X1 U4213 ( .A(n4630), .ZN(n3420) );
  OAI22_X1 U4214 ( .A1(n3490), .A2(n4627), .B1(n4267), .B2(n3407), .ZN(n3412)
         );
  INV_X1 U4215 ( .A(n3843), .ZN(n3408) );
  NAND3_X1 U4216 ( .A1(n3452), .A2(n3855), .A3(n3408), .ZN(n3409) );
  AOI21_X1 U4217 ( .B1(n3410), .B2(n3409), .A(n4585), .ZN(n3411) );
  AOI211_X1 U4218 ( .C1(n4603), .C2(n3054), .A(n3412), .B(n3411), .ZN(n3413)
         );
  OAI21_X1 U4219 ( .B1(n4680), .B2(n4608), .A(n3413), .ZN(n4681) );
  NAND2_X1 U4220 ( .A1(n4681), .A2(n3379), .ZN(n3419) );
  AND2_X1 U4221 ( .A1(n4674), .A2(n3860), .ZN(n3414) );
  NOR2_X1 U4222 ( .A1(n3415), .A2(n3414), .ZN(n4683) );
  INV_X1 U4223 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3416) );
  OAI22_X1 U4224 ( .A1(n3379), .A2(n3416), .B1(n4255), .B2(REG3_REG_3__SCAN_IN), .ZN(n3417) );
  AOI21_X1 U4225 ( .B1(n4683), .B2(n4617), .A(n3417), .ZN(n3418) );
  OAI211_X1 U4226 ( .C1(n4680), .C2(n3420), .A(n3419), .B(n3418), .ZN(U3287)
         );
  NAND2_X1 U4227 ( .A1(n3874), .A2(n3884), .ZN(n3815) );
  XOR2_X1 U4228 ( .A(n3815), .B(n3421), .Z(n3464) );
  INV_X1 U4229 ( .A(n3464), .ZN(n3435) );
  OAI21_X1 U4230 ( .B1(n3422), .B2(n3428), .A(n3510), .ZN(n3469) );
  INV_X1 U4231 ( .A(n3469), .ZN(n3426) );
  INV_X1 U4232 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3424) );
  OAI22_X1 U4233 ( .A1(n3379), .A2(n3424), .B1(n3423), .B2(n4255), .ZN(n3425)
         );
  AOI21_X1 U4234 ( .B1(n3426), .B2(n4617), .A(n3425), .ZN(n3434) );
  XOR2_X1 U4235 ( .A(n3815), .B(n3427), .Z(n3432) );
  OAI22_X1 U4236 ( .A1(n3429), .A2(n4627), .B1(n3428), .B2(n4267), .ZN(n3430)
         );
  AOI21_X1 U4237 ( .B1(n4603), .B2(n3944), .A(n3430), .ZN(n3431) );
  OAI21_X1 U4238 ( .B1(n3432), .B2(n4585), .A(n3431), .ZN(n3463) );
  NAND2_X1 U4239 ( .A1(n3463), .A2(n3379), .ZN(n3433) );
  OAI211_X1 U4240 ( .C1(n3435), .C2(n4262), .A(n3434), .B(n3433), .ZN(U3282)
         );
  INV_X1 U4241 ( .A(n3513), .ZN(n3445) );
  XNOR2_X1 U4242 ( .A(n3437), .B(n3436), .ZN(n3438) );
  NAND2_X1 U4243 ( .A1(n3438), .A2(n4424), .ZN(n3444) );
  INV_X1 U4244 ( .A(n4580), .ZN(n3726) );
  OAI22_X1 U4245 ( .A1(n3505), .A2(n4414), .B1(n4413), .B2(n3726), .ZN(n3442)
         );
  INV_X1 U4246 ( .A(n3439), .ZN(n3440) );
  OAI21_X1 U4247 ( .B1(n3762), .B2(n2117), .A(n3440), .ZN(n3441) );
  NOR2_X1 U4248 ( .A1(n3442), .A2(n3441), .ZN(n3443) );
  OAI211_X1 U4249 ( .C1(n4429), .C2(n3445), .A(n3444), .B(n3443), .ZN(U3228)
         );
  OAI21_X1 U4250 ( .B1(n3447), .B2(n3450), .A(n3446), .ZN(n4677) );
  INV_X1 U4251 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3449) );
  NAND2_X1 U4252 ( .A1(n4614), .A2(n3052), .ZN(n4673) );
  NAND3_X1 U4253 ( .A1(n4617), .A2(n4674), .A3(n4673), .ZN(n3448) );
  OAI21_X1 U4254 ( .B1(n4255), .B2(n3449), .A(n3448), .ZN(n3461) );
  NAND3_X1 U4255 ( .A1(n4599), .A2(n3450), .A3(n3854), .ZN(n3451) );
  NAND2_X1 U4256 ( .A1(n3452), .A2(n3451), .ZN(n3457) );
  NAND2_X1 U4257 ( .A1(n3049), .A2(n4603), .ZN(n3454) );
  NAND2_X1 U4258 ( .A1(n3948), .A2(n4581), .ZN(n3453) );
  OAI211_X1 U4259 ( .C1(n4267), .C2(n3455), .A(n3454), .B(n3453), .ZN(n3456)
         );
  AOI21_X1 U4260 ( .B1(n3457), .B2(n4624), .A(n3456), .ZN(n3459) );
  NAND2_X1 U4261 ( .A1(n4677), .A2(n4625), .ZN(n3458) );
  NAND2_X1 U4262 ( .A1(n3459), .A2(n3458), .ZN(n4675) );
  MUX2_X1 U4263 ( .A(REG2_REG_2__SCAN_IN), .B(n4675), .S(n3379), .Z(n3460) );
  AOI211_X1 U4264 ( .C1(n4630), .C2(n4677), .A(n3461), .B(n3460), .ZN(n3462)
         );
  INV_X1 U4265 ( .A(n3462), .ZN(U3288) );
  INV_X1 U4266 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3465) );
  AOI21_X1 U4267 ( .B1(n3464), .B2(n4704), .A(n3463), .ZN(n3467) );
  MUX2_X1 U4268 ( .A(n3465), .B(n3467), .S(n4722), .Z(n3466) );
  OAI21_X1 U4269 ( .B1(n3469), .B2(n4384), .A(n3466), .ZN(U3483) );
  MUX2_X1 U4270 ( .A(n2524), .B(n3467), .S(n4735), .Z(n3468) );
  OAI21_X1 U4271 ( .B1(n3469), .B2(n4328), .A(n3468), .ZN(U3526) );
  NAND2_X1 U4272 ( .A1(n3887), .A2(n3893), .ZN(n3809) );
  INV_X1 U4273 ( .A(n3809), .ZN(n3471) );
  XNOR2_X1 U4274 ( .A(n3470), .B(n3471), .ZN(n4710) );
  NAND2_X1 U4275 ( .A1(n4710), .A2(n4625), .ZN(n3480) );
  XNOR2_X1 U4276 ( .A(n3472), .B(n3471), .ZN(n3478) );
  NAND2_X1 U4277 ( .A1(n3473), .A2(n4603), .ZN(n3475) );
  NAND2_X1 U4278 ( .A1(n3942), .A2(n4581), .ZN(n3474) );
  OAI211_X1 U4279 ( .C1(n4267), .C2(n3476), .A(n3475), .B(n3474), .ZN(n3477)
         );
  AOI21_X1 U4280 ( .B1(n3478), .B2(n4624), .A(n3477), .ZN(n3479) );
  NAND2_X1 U4281 ( .A1(n3512), .A2(n3481), .ZN(n4706) );
  AND3_X1 U4282 ( .A1(n2118), .A2(n4617), .A3(n4706), .ZN(n3484) );
  OAI22_X1 U4283 ( .A1(n3379), .A2(n3016), .B1(n3482), .B2(n4255), .ZN(n3483)
         );
  AOI211_X1 U4284 ( .C1(n4710), .C2(n4630), .A(n3484), .B(n3483), .ZN(n3485)
         );
  OAI21_X1 U4285 ( .B1(n4712), .B2(n4634), .A(n3485), .ZN(U3280) );
  INV_X1 U4286 ( .A(n3486), .ZN(n3864) );
  NAND2_X1 U4287 ( .A1(n3864), .A2(n3881), .ZN(n3810) );
  XNOR2_X1 U4288 ( .A(n3487), .B(n3810), .ZN(n3492) );
  AOI22_X1 U4289 ( .A1(n3945), .A2(n4581), .B1(n4602), .B2(n3488), .ZN(n3489)
         );
  OAI21_X1 U4290 ( .B1(n3490), .B2(n4207), .A(n3489), .ZN(n3491) );
  AOI21_X1 U4291 ( .B1(n3492), .B2(n4624), .A(n3491), .ZN(n4690) );
  XOR2_X1 U4292 ( .A(n3810), .B(n3493), .Z(n4693) );
  INV_X1 U4293 ( .A(n3494), .ZN(n3497) );
  OAI21_X1 U4294 ( .B1(n3497), .B2(n3496), .A(n3495), .ZN(n4691) );
  NOR2_X1 U4295 ( .A1(n4691), .A2(n4235), .ZN(n3501) );
  OAI22_X1 U4296 ( .A1(n3379), .A2(n3499), .B1(n3498), .B2(n4255), .ZN(n3500)
         );
  AOI211_X1 U4297 ( .C1(n4693), .C2(n4237), .A(n3501), .B(n3500), .ZN(n3502)
         );
  OAI21_X1 U4298 ( .B1(n4634), .B2(n4690), .A(n3502), .ZN(U3285) );
  INV_X1 U4299 ( .A(n3878), .ZN(n3885) );
  NAND2_X1 U4300 ( .A1(n3885), .A2(n3875), .ZN(n3816) );
  XNOR2_X1 U4301 ( .A(n3503), .B(n3816), .ZN(n3507) );
  AOI22_X1 U4302 ( .A1(n4580), .A2(n4581), .B1(n4602), .B2(n3509), .ZN(n3504)
         );
  OAI21_X1 U4303 ( .B1(n3505), .B2(n4207), .A(n3504), .ZN(n3506) );
  AOI21_X1 U4304 ( .B1(n3507), .B2(n4624), .A(n3506), .ZN(n4699) );
  XNOR2_X1 U4305 ( .A(n3508), .B(n3816), .ZN(n4703) );
  NAND2_X1 U4306 ( .A1(n3510), .A2(n3509), .ZN(n3511) );
  NAND2_X1 U4307 ( .A1(n3512), .A2(n3511), .ZN(n4700) );
  AOI22_X1 U4308 ( .A1(n4634), .A2(REG2_REG_9__SCAN_IN), .B1(n3513), .B2(n4629), .ZN(n3514) );
  OAI21_X1 U4309 ( .B1(n4700), .B2(n4235), .A(n3514), .ZN(n3515) );
  AOI21_X1 U4310 ( .B1(n4703), .B2(n4237), .A(n3515), .ZN(n3516) );
  OAI21_X1 U4311 ( .B1(n4634), .B2(n4699), .A(n3516), .ZN(U3281) );
  INV_X1 U4312 ( .A(n3535), .ZN(n3517) );
  OR2_X1 U4313 ( .A1(n3536), .A2(n3517), .ZN(n3830) );
  XNOR2_X1 U4314 ( .A(n3537), .B(n3830), .ZN(n3520) );
  INV_X1 U4315 ( .A(n3941), .ZN(n3657) );
  OAI22_X1 U4316 ( .A1(n3657), .A2(n4627), .B1(n3658), .B2(n4267), .ZN(n3518)
         );
  AOI21_X1 U4317 ( .B1(n4603), .B2(n3942), .A(n3518), .ZN(n3519) );
  OAI21_X1 U4318 ( .B1(n3520), .B2(n4585), .A(n3519), .ZN(n3527) );
  INV_X1 U4319 ( .A(n3527), .ZN(n3526) );
  XNOR2_X1 U4320 ( .A(n3521), .B(n3830), .ZN(n3528) );
  OR2_X1 U4321 ( .A1(n4589), .A2(n3658), .ZN(n3522) );
  NAND2_X1 U4322 ( .A1(n3545), .A2(n3522), .ZN(n3533) );
  AOI22_X1 U4323 ( .A1(n4634), .A2(REG2_REG_12__SCAN_IN), .B1(n3649), .B2(
        n4629), .ZN(n3523) );
  OAI21_X1 U4324 ( .B1(n3533), .B2(n4235), .A(n3523), .ZN(n3524) );
  AOI21_X1 U4325 ( .B1(n3528), .B2(n4237), .A(n3524), .ZN(n3525) );
  OAI21_X1 U4326 ( .B1(n3526), .B2(n4634), .A(n3525), .ZN(U3278) );
  AOI21_X1 U4327 ( .B1(n4704), .B2(n3528), .A(n3527), .ZN(n3530) );
  MUX2_X1 U4328 ( .A(n2597), .B(n3530), .S(n4735), .Z(n3529) );
  OAI21_X1 U4329 ( .B1(n3533), .B2(n4328), .A(n3529), .ZN(U3530) );
  INV_X1 U4330 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3531) );
  MUX2_X1 U4331 ( .A(n3531), .B(n3530), .S(n4722), .Z(n3532) );
  OAI21_X1 U4332 ( .B1(n3533), .B2(n4384), .A(n3532), .ZN(U3491) );
  OR2_X1 U4333 ( .A1(n3534), .A2(n2079), .ZN(n3827) );
  XNOR2_X1 U4334 ( .A(n2063), .B(n3827), .ZN(n3543) );
  INV_X1 U4335 ( .A(n4252), .ZN(n3759) );
  OAI22_X1 U4336 ( .A1(n3759), .A2(n4627), .B1(n4267), .B2(n3705), .ZN(n3541)
         );
  OAI21_X1 U4337 ( .B1(n3537), .B2(n3536), .A(n3535), .ZN(n3538) );
  XNOR2_X1 U4338 ( .A(n3538), .B(n3827), .ZN(n3539) );
  NOR2_X1 U4339 ( .A1(n3539), .A2(n4585), .ZN(n3540) );
  AOI211_X1 U4340 ( .C1(n4603), .C2(n4582), .A(n3541), .B(n3540), .ZN(n3542)
         );
  OAI21_X1 U4341 ( .B1(n3543), .B2(n4608), .A(n3542), .ZN(n3564) );
  INV_X1 U4342 ( .A(n3564), .ZN(n3550) );
  INV_X1 U4343 ( .A(n3543), .ZN(n3565) );
  NAND2_X1 U4344 ( .A1(n3545), .A2(n3544), .ZN(n3546) );
  NAND2_X1 U4345 ( .A1(n3557), .A2(n3546), .ZN(n3570) );
  AOI22_X1 U4346 ( .A1(n4634), .A2(REG2_REG_13__SCAN_IN), .B1(n3697), .B2(
        n4629), .ZN(n3547) );
  OAI21_X1 U4347 ( .B1(n3570), .B2(n4235), .A(n3547), .ZN(n3548) );
  AOI21_X1 U4348 ( .B1(n3565), .B2(n4630), .A(n3548), .ZN(n3549) );
  OAI21_X1 U4349 ( .B1(n3550), .B2(n4634), .A(n3549), .ZN(U3277) );
  XNOR2_X1 U4350 ( .A(n3771), .B(n3808), .ZN(n3555) );
  AOI22_X1 U4351 ( .A1(n3940), .A2(n4581), .B1(n4602), .B2(n3556), .ZN(n3551)
         );
  OAI21_X1 U4352 ( .B1(n3657), .B2(n4207), .A(n3551), .ZN(n3554) );
  AOI21_X1 U4353 ( .B1(n3808), .B2(n3552), .A(n4240), .ZN(n4343) );
  NOR2_X1 U4354 ( .A1(n4343), .A2(n4608), .ZN(n3553) );
  AOI211_X1 U4355 ( .C1(n3555), .C2(n4624), .A(n3554), .B(n3553), .ZN(n4342)
         );
  INV_X1 U4356 ( .A(n4343), .ZN(n3562) );
  NAND2_X1 U4357 ( .A1(n3557), .A2(n3556), .ZN(n4339) );
  AND3_X1 U4358 ( .A1(n4340), .A2(n4617), .A3(n4339), .ZN(n3561) );
  INV_X1 U4359 ( .A(REG2_REG_14__SCAN_IN), .ZN(n3559) );
  INV_X1 U4360 ( .A(n3558), .ZN(n3630) );
  OAI22_X1 U4361 ( .A1(n3379), .A2(n3559), .B1(n3630), .B2(n4255), .ZN(n3560)
         );
  AOI211_X1 U4362 ( .C1(n3562), .C2(n4630), .A(n3561), .B(n3560), .ZN(n3563)
         );
  OAI21_X1 U4363 ( .B1(n4342), .B2(n4634), .A(n3563), .ZN(U3276) );
  INV_X1 U4364 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3566) );
  AOI21_X1 U4365 ( .B1(n4716), .B2(n3565), .A(n3564), .ZN(n3568) );
  MUX2_X1 U4366 ( .A(n3566), .B(n3568), .S(n4722), .Z(n3567) );
  OAI21_X1 U4367 ( .B1(n3570), .B2(n4384), .A(n3567), .ZN(U3493) );
  MUX2_X1 U4368 ( .A(n3998), .B(n3568), .S(n4735), .Z(n3569) );
  OAI21_X1 U4369 ( .B1(n4328), .B2(n3570), .A(n3569), .ZN(U3531) );
  OAI22_X1 U4370 ( .A1(n4412), .A2(n4627), .B1(n4267), .B2(n3576), .ZN(n3575)
         );
  INV_X1 U4371 ( .A(n3571), .ZN(n3573) );
  AOI211_X1 U4372 ( .C1(n3573), .C2(n3572), .A(n4585), .B(n4160), .ZN(n3574)
         );
  AOI211_X1 U4373 ( .C1(n4603), .C2(n3940), .A(n3575), .B(n3574), .ZN(n4331)
         );
  OR2_X1 U4374 ( .A1(n4253), .A2(n3576), .ZN(n3577) );
  NAND2_X1 U4375 ( .A1(n4230), .A2(n3577), .ZN(n4332) );
  INV_X1 U4376 ( .A(n4332), .ZN(n3580) );
  INV_X1 U4377 ( .A(REG2_REG_16__SCAN_IN), .ZN(n3578) );
  OAI22_X1 U4378 ( .A1(n3379), .A2(n3578), .B1(n4428), .B2(n4255), .ZN(n3579)
         );
  AOI21_X1 U4379 ( .B1(n3580), .B2(n4617), .A(n3579), .ZN(n3583) );
  XNOR2_X1 U4380 ( .A(n3581), .B(n3819), .ZN(n4329) );
  NAND2_X1 U4381 ( .A1(n4329), .A2(n4237), .ZN(n3582) );
  OAI211_X1 U4382 ( .C1(n4331), .C2(n4634), .A(n3583), .B(n3582), .ZN(U3274)
         );
  AOI22_X1 U4383 ( .A1(n3585), .A2(n3807), .B1(n3584), .B2(n4036), .ZN(n3586)
         );
  NAND2_X1 U4384 ( .A1(n2041), .A2(DATAI_29_), .ZN(n3587) );
  XNOR2_X1 U4385 ( .A(n3792), .B(n3587), .ZN(n3839) );
  AOI21_X1 U4386 ( .B1(n3791), .B2(n3588), .A(n4271), .ZN(n4282) );
  AOI22_X1 U4387 ( .A1(n4282), .A2(n4617), .B1(REG2_REG_29__SCAN_IN), .B2(
        n4634), .ZN(n3598) );
  XOR2_X1 U4388 ( .A(n3839), .B(n3589), .Z(n3593) );
  NAND2_X1 U4389 ( .A1(n2391), .A2(REG2_REG_30__SCAN_IN), .ZN(n3591) );
  NAND2_X1 U4390 ( .A1(n2043), .A2(REG0_REG_30__SCAN_IN), .ZN(n3590) );
  OAI211_X1 U4391 ( .C1(n3786), .C2(n4278), .A(n3591), .B(n3590), .ZN(n3937)
         );
  AOI21_X1 U4392 ( .B1(B_REG_SCAN_IN), .B2(n4438), .A(n4627), .ZN(n4265) );
  AOI22_X1 U4393 ( .A1(n3937), .A2(n4265), .B1(n4602), .B2(n3791), .ZN(n3592)
         );
  INV_X1 U4394 ( .A(n3594), .ZN(n3595) );
  NOR2_X1 U4395 ( .A1(n3595), .A2(n4255), .ZN(n3596) );
  OAI21_X1 U4396 ( .B1(n4281), .B2(n3596), .A(n3379), .ZN(n3597) );
  OAI211_X1 U4397 ( .C1(n4280), .C2(n4262), .A(n3598), .B(n3597), .ZN(U3354)
         );
  INV_X1 U4398 ( .A(n3599), .ZN(n3605) );
  INV_X1 U4399 ( .A(REG2_REG_28__SCAN_IN), .ZN(n3600) );
  OAI22_X1 U4400 ( .A1(n3601), .A2(n4255), .B1(n3600), .B2(n3379), .ZN(n3604)
         );
  NOR2_X1 U4401 ( .A1(n3602), .A2(n4634), .ZN(n3603) );
  AOI211_X1 U4402 ( .C1(n4617), .C2(n3605), .A(n3604), .B(n3603), .ZN(n3606)
         );
  OAI21_X1 U4403 ( .B1(n3607), .B2(n4262), .A(n3606), .ZN(U3262) );
  XNOR2_X1 U4404 ( .A(n3609), .B(n3608), .ZN(n3616) );
  INV_X1 U4405 ( .A(n3610), .ZN(n4039) );
  OAI22_X1 U4406 ( .A1(n3762), .A2(n4038), .B1(STATE_REG_SCAN_IN), .B2(n3611), 
        .ZN(n3614) );
  INV_X1 U4407 ( .A(n4036), .ZN(n3612) );
  OAI22_X1 U4408 ( .A1(n3612), .A2(n4413), .B1(n4029), .B2(n4414), .ZN(n3613)
         );
  AOI211_X1 U4409 ( .C1(n4039), .C2(n3751), .A(n3614), .B(n3613), .ZN(n3615)
         );
  OAI21_X1 U4410 ( .B1(n3616), .B2(n3753), .A(n3615), .ZN(U3211) );
  INV_X1 U4411 ( .A(n3701), .ZN(n3618) );
  OAI21_X1 U4412 ( .B1(n3618), .B2(n3617), .A(n3698), .ZN(n3619) );
  OAI21_X1 U4413 ( .B1(n3699), .B2(n3701), .A(n3619), .ZN(n3623) );
  NAND2_X1 U4414 ( .A1(n3621), .A2(n3620), .ZN(n3622) );
  XNOR2_X1 U4415 ( .A(n3623), .B(n3622), .ZN(n3624) );
  NAND2_X1 U4416 ( .A1(n3624), .A2(n4424), .ZN(n3629) );
  INV_X1 U4417 ( .A(n3940), .ZN(n4415) );
  OAI22_X1 U4418 ( .A1(n3657), .A2(n4414), .B1(n4413), .B2(n4415), .ZN(n3627)
         );
  NAND2_X1 U4419 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4537) );
  OAI21_X1 U4420 ( .B1(n3762), .B2(n3625), .A(n4537), .ZN(n3626) );
  NOR2_X1 U4421 ( .A1(n3627), .A2(n3626), .ZN(n3628) );
  OAI211_X1 U4422 ( .C1(n4429), .C2(n3630), .A(n3629), .B(n3628), .ZN(U3212)
         );
  OAI21_X1 U4423 ( .B1(n3711), .B2(n3633), .A(n3632), .ZN(n3634) );
  NAND3_X1 U4424 ( .A1(n2155), .A2(n4424), .A3(n3634), .ZN(n3640) );
  OAI22_X1 U4425 ( .A1(n3762), .A2(n4115), .B1(STATE_REG_SCAN_IN), .B2(n3635), 
        .ZN(n3638) );
  OAI22_X1 U4426 ( .A1(n4067), .A2(n4413), .B1(n4414), .B2(n3636), .ZN(n3637)
         );
  AOI211_X1 U4427 ( .C1(n4117), .C2(n3751), .A(n3638), .B(n3637), .ZN(n3639)
         );
  NAND2_X1 U4428 ( .A1(n3640), .A2(n3639), .ZN(U3213) );
  INV_X1 U4429 ( .A(n3641), .ZN(n4198) );
  XNOR2_X1 U4430 ( .A(n3643), .B(n3642), .ZN(n3644) );
  NAND2_X1 U4431 ( .A1(n3644), .A2(n4424), .ZN(n3648) );
  OAI22_X1 U4432 ( .A1(n3076), .A2(n4414), .B1(n4413), .B2(n4189), .ZN(n3646)
         );
  NAND2_X1 U4433 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4023) );
  OAI21_X1 U4434 ( .B1(n3762), .B2(n4188), .A(n4023), .ZN(n3645) );
  NOR2_X1 U4435 ( .A1(n3646), .A2(n3645), .ZN(n3647) );
  OAI211_X1 U4436 ( .C1(n4429), .C2(n4198), .A(n3648), .B(n3647), .ZN(U3216)
         );
  INV_X1 U4437 ( .A(n3649), .ZN(n3663) );
  INV_X1 U4438 ( .A(n3650), .ZN(n3652) );
  NAND2_X1 U4439 ( .A1(n3652), .A2(n3651), .ZN(n3653) );
  XNOR2_X1 U4440 ( .A(n3654), .B(n3653), .ZN(n3655) );
  NAND2_X1 U4441 ( .A1(n3655), .A2(n4424), .ZN(n3662) );
  OAI22_X1 U4442 ( .A1(n3657), .A2(n4413), .B1(n4414), .B2(n3656), .ZN(n3660)
         );
  NAND2_X1 U4443 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4508) );
  OAI21_X1 U4444 ( .B1(n3762), .B2(n3658), .A(n4508), .ZN(n3659) );
  NOR2_X1 U4445 ( .A1(n3660), .A2(n3659), .ZN(n3661) );
  OAI211_X1 U4446 ( .C1(n4429), .C2(n3663), .A(n3662), .B(n3661), .ZN(U3221)
         );
  NOR2_X1 U4447 ( .A1(n3665), .A2(n2141), .ZN(n3666) );
  XNOR2_X1 U4448 ( .A(n3667), .B(n3666), .ZN(n3673) );
  INV_X1 U4449 ( .A(n3668), .ZN(n4075) );
  INV_X1 U4450 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3669) );
  OAI22_X1 U4451 ( .A1(n3762), .A2(n4072), .B1(STATE_REG_SCAN_IN), .B2(n3669), 
        .ZN(n3671) );
  OAI22_X1 U4452 ( .A1(n4029), .A2(n4413), .B1(n4067), .B2(n4414), .ZN(n3670)
         );
  AOI211_X1 U4453 ( .C1(n4075), .C2(n3751), .A(n3671), .B(n3670), .ZN(n3672)
         );
  OAI21_X1 U4454 ( .B1(n3673), .B2(n3753), .A(n3672), .ZN(U3222) );
  INV_X1 U4455 ( .A(n4233), .ZN(n3685) );
  XNOR2_X1 U4456 ( .A(n3676), .B(n3675), .ZN(n3677) );
  XNOR2_X1 U4457 ( .A(n3674), .B(n3677), .ZN(n3678) );
  NAND2_X1 U4458 ( .A1(n3678), .A2(n4424), .ZN(n3684) );
  INV_X1 U4459 ( .A(n4224), .ZN(n4245) );
  OAI22_X1 U4460 ( .A1(n4245), .A2(n4414), .B1(n4413), .B2(n3076), .ZN(n3682)
         );
  INV_X1 U4461 ( .A(REG3_REG_17__SCAN_IN), .ZN(n3679) );
  NOR2_X1 U4462 ( .A1(STATE_REG_SCAN_IN), .A2(n3679), .ZN(n4562) );
  INV_X1 U4463 ( .A(n4562), .ZN(n3680) );
  OAI21_X1 U4464 ( .B1(n3762), .B2(n4222), .A(n3680), .ZN(n3681) );
  NOR2_X1 U4465 ( .A1(n3682), .A2(n3681), .ZN(n3683) );
  OAI211_X1 U4466 ( .C1(n4429), .C2(n3685), .A(n3684), .B(n3683), .ZN(U3225)
         );
  INV_X1 U4467 ( .A(n3686), .ZN(n3687) );
  NAND2_X1 U4468 ( .A1(n3688), .A2(n3687), .ZN(n3689) );
  XOR2_X1 U4469 ( .A(n3690), .B(n3689), .Z(n3691) );
  NAND2_X1 U4470 ( .A1(n3691), .A2(n4424), .ZN(n3696) );
  INV_X1 U4471 ( .A(n4086), .ZN(n3747) );
  INV_X1 U4472 ( .A(n4126), .ZN(n3716) );
  OAI22_X1 U4473 ( .A1(n3747), .A2(n4413), .B1(n4414), .B2(n3716), .ZN(n3694)
         );
  OAI22_X1 U4474 ( .A1(n3762), .A2(n4092), .B1(STATE_REG_SCAN_IN), .B2(n3692), 
        .ZN(n3693) );
  NOR2_X1 U4475 ( .A1(n3694), .A2(n3693), .ZN(n3695) );
  OAI211_X1 U4476 ( .C1(n4429), .C2(n4094), .A(n3696), .B(n3695), .ZN(U3226)
         );
  INV_X1 U4477 ( .A(n3697), .ZN(n3710) );
  XNOR2_X1 U4478 ( .A(n3699), .B(n3698), .ZN(n3700) );
  XNOR2_X1 U4479 ( .A(n3701), .B(n3700), .ZN(n3702) );
  NAND2_X1 U4480 ( .A1(n3702), .A2(n4424), .ZN(n3709) );
  INV_X1 U4481 ( .A(n4582), .ZN(n3725) );
  OAI22_X1 U4482 ( .A1(n3759), .A2(n4413), .B1(n4414), .B2(n3725), .ZN(n3707)
         );
  INV_X1 U4483 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3703) );
  NOR2_X1 U4484 ( .A1(STATE_REG_SCAN_IN), .A2(n3703), .ZN(n4519) );
  INV_X1 U4485 ( .A(n4519), .ZN(n3704) );
  OAI21_X1 U4486 ( .B1(n3762), .B2(n3705), .A(n3704), .ZN(n3706) );
  NOR2_X1 U4487 ( .A1(n3707), .A2(n3706), .ZN(n3708) );
  OAI211_X1 U4488 ( .C1(n4429), .C2(n3710), .A(n3709), .B(n3708), .ZN(U3231)
         );
  AOI21_X1 U4489 ( .B1(n3713), .B2(n3712), .A(n3711), .ZN(n3720) );
  OAI22_X1 U4490 ( .A1(n3762), .A2(n4129), .B1(STATE_REG_SCAN_IN), .B2(n3714), 
        .ZN(n3718) );
  OAI22_X1 U4491 ( .A1(n3716), .A2(n4413), .B1(n4414), .B2(n3715), .ZN(n3717)
         );
  AOI211_X1 U4492 ( .C1(n4132), .C2(n3751), .A(n3718), .B(n3717), .ZN(n3719)
         );
  OAI21_X1 U4493 ( .B1(n3720), .B2(n3753), .A(n3719), .ZN(U3232) );
  XOR2_X1 U4494 ( .A(n3722), .B(n3721), .Z(n3723) );
  XNOR2_X1 U4495 ( .A(n3724), .B(n3723), .ZN(n3731) );
  OAI22_X1 U4496 ( .A1(n3726), .A2(n4414), .B1(n4413), .B2(n3725), .ZN(n3727)
         );
  AOI211_X1 U4497 ( .C1(n4590), .C2(n4417), .A(n3728), .B(n3727), .ZN(n3730)
         );
  NAND2_X1 U4498 ( .A1(n3751), .A2(n4588), .ZN(n3729) );
  OAI211_X1 U4499 ( .C1(n3731), .C2(n3753), .A(n3730), .B(n3729), .ZN(U3233)
         );
  INV_X1 U4500 ( .A(n4216), .ZN(n3743) );
  INV_X1 U4501 ( .A(n3732), .ZN(n3734) );
  NAND2_X1 U4502 ( .A1(n3734), .A2(n3733), .ZN(n3735) );
  XNOR2_X1 U4503 ( .A(n3736), .B(n3735), .ZN(n3737) );
  NAND2_X1 U4504 ( .A1(n3737), .A2(n4424), .ZN(n3742) );
  OAI22_X1 U4505 ( .A1(n3738), .A2(n4413), .B1(n4414), .B2(n4412), .ZN(n3740)
         );
  OAI21_X1 U4506 ( .B1(n3762), .B2(n4213), .A(n2287), .ZN(n3739) );
  NOR2_X1 U4507 ( .A1(n3740), .A2(n3739), .ZN(n3741) );
  OAI211_X1 U4508 ( .C1(n4429), .C2(n3743), .A(n3742), .B(n3741), .ZN(U3235)
         );
  NAND2_X1 U4509 ( .A1(n3744), .A2(n2067), .ZN(n3745) );
  XNOR2_X1 U4510 ( .A(n2057), .B(n3745), .ZN(n3754) );
  OAI22_X1 U4511 ( .A1(n3762), .A2(n4058), .B1(STATE_REG_SCAN_IN), .B2(n3746), 
        .ZN(n3750) );
  OAI22_X1 U4512 ( .A1(n3748), .A2(n4413), .B1(n3747), .B2(n4414), .ZN(n3749)
         );
  AOI211_X1 U4513 ( .C1(n4059), .C2(n3751), .A(n3750), .B(n3749), .ZN(n3752)
         );
  OAI21_X1 U4514 ( .B1(n3754), .B2(n3753), .A(n3752), .ZN(U3237) );
  INV_X1 U4515 ( .A(n3755), .ZN(n4256) );
  INV_X1 U4516 ( .A(n4420), .ZN(n3756) );
  NOR2_X1 U4517 ( .A1(n4419), .A2(n3756), .ZN(n3757) );
  XNOR2_X1 U4518 ( .A(n3757), .B(n4421), .ZN(n3758) );
  NAND2_X1 U4519 ( .A1(n3758), .A2(n4424), .ZN(n3766) );
  OAI22_X1 U4520 ( .A1(n4245), .A2(n4413), .B1(n4414), .B2(n3759), .ZN(n3764)
         );
  NOR2_X1 U4521 ( .A1(STATE_REG_SCAN_IN), .A2(n3760), .ZN(n4544) );
  INV_X1 U4522 ( .A(n4544), .ZN(n3761) );
  OAI21_X1 U4523 ( .B1(n3762), .B2(n4244), .A(n3761), .ZN(n3763) );
  NOR2_X1 U4524 ( .A1(n3764), .A2(n3763), .ZN(n3765) );
  OAI211_X1 U4525 ( .C1(n4429), .C2(n4256), .A(n3766), .B(n3765), .ZN(U3238)
         );
  NAND2_X1 U4526 ( .A1(n3767), .A2(n3770), .ZN(n3848) );
  NAND2_X1 U4527 ( .A1(n3769), .A2(n3768), .ZN(n3879) );
  NAND2_X1 U4528 ( .A1(n3879), .A2(n3770), .ZN(n3899) );
  OAI21_X1 U4529 ( .B1(n3771), .B2(n3848), .A(n3899), .ZN(n3773) );
  AOI21_X1 U4530 ( .B1(n3773), .B2(n3901), .A(n3772), .ZN(n3774) );
  INV_X1 U4531 ( .A(n3774), .ZN(n3775) );
  AOI21_X1 U4532 ( .B1(n3775), .B2(n3906), .A(n2222), .ZN(n3777) );
  OAI21_X1 U4533 ( .B1(n3777), .B2(n3908), .A(n3776), .ZN(n3780) );
  INV_X1 U4534 ( .A(n3778), .ZN(n3825) );
  NOR2_X1 U4535 ( .A1(n3834), .A2(n3825), .ZN(n3915) );
  INV_X1 U4536 ( .A(n3915), .ZN(n3779) );
  AOI21_X1 U4537 ( .B1(n3910), .B2(n3780), .A(n3779), .ZN(n3790) );
  NAND2_X1 U4538 ( .A1(n3782), .A2(n3781), .ZN(n3797) );
  NAND2_X1 U4539 ( .A1(n3792), .A2(n3791), .ZN(n3789) );
  INV_X1 U4540 ( .A(REG1_REG_31__SCAN_IN), .ZN(n3785) );
  NAND2_X1 U4541 ( .A1(n2730), .A2(REG2_REG_31__SCAN_IN), .ZN(n3784) );
  NAND2_X1 U4542 ( .A1(n2043), .A2(REG0_REG_31__SCAN_IN), .ZN(n3783) );
  OAI211_X1 U4543 ( .C1(n3786), .C2(n3785), .A(n3784), .B(n3783), .ZN(n4266)
         );
  NAND2_X1 U4544 ( .A1(n3787), .A2(DATAI_31_), .ZN(n4268) );
  NAND2_X1 U4545 ( .A1(n4266), .A2(n4268), .ZN(n3922) );
  NAND2_X1 U4546 ( .A1(n3787), .A2(DATAI_30_), .ZN(n4263) );
  OR2_X1 U4547 ( .A1(n3937), .A2(n4263), .ZN(n3788) );
  AND2_X1 U4548 ( .A1(n3922), .A2(n3788), .ZN(n3833) );
  NAND2_X1 U4549 ( .A1(n3789), .A2(n3833), .ZN(n3795) );
  NOR4_X1 U4550 ( .A1(n3790), .A2(n3797), .A3(n3916), .A4(n3795), .ZN(n3801)
         );
  OR2_X1 U4551 ( .A1(n3792), .A2(n3791), .ZN(n3793) );
  AND2_X1 U4552 ( .A1(n3794), .A2(n3793), .ZN(n3796) );
  INV_X1 U4553 ( .A(n3796), .ZN(n3918) );
  NOR3_X1 U4554 ( .A1(n3918), .A2(n3919), .A3(n4031), .ZN(n3799) );
  AOI21_X1 U4555 ( .B1(n3797), .B2(n3796), .A(n3795), .ZN(n3923) );
  INV_X1 U4556 ( .A(n3923), .ZN(n3798) );
  NOR2_X1 U4557 ( .A1(n3799), .A2(n3798), .ZN(n3800) );
  OAI22_X1 U4558 ( .A1(n3801), .A2(n3800), .B1(n4263), .B2(n4266), .ZN(n3929)
         );
  INV_X1 U4559 ( .A(n3937), .ZN(n3802) );
  INV_X1 U4560 ( .A(n4263), .ZN(n4277) );
  NOR2_X1 U4561 ( .A1(n3802), .A2(n4277), .ZN(n3836) );
  INV_X1 U4562 ( .A(n3836), .ZN(n3803) );
  AOI21_X1 U4563 ( .B1(n3803), .B2(n4266), .A(n4268), .ZN(n3805) );
  NOR2_X1 U4564 ( .A1(n3805), .A2(n3804), .ZN(n3928) );
  XNOR2_X1 U4565 ( .A(n4126), .B(n3806), .ZN(n4101) );
  INV_X1 U4566 ( .A(n4101), .ZN(n4107) );
  NOR3_X1 U4567 ( .A1(n3807), .A2(n4031), .A3(n4107), .ZN(n3824) );
  NOR4_X1 U4568 ( .A1(n2281), .A2(n3810), .A3(n4211), .A4(n3809), .ZN(n3823)
         );
  INV_X1 U4569 ( .A(n3905), .ZN(n3811) );
  NAND2_X1 U4570 ( .A1(n3811), .A2(n4104), .ZN(n4149) );
  NOR4_X1 U4571 ( .A1(n4149), .A2(n4578), .A3(n3813), .A4(n3812), .ZN(n3822)
         );
  INV_X1 U4572 ( .A(n3903), .ZN(n4163) );
  OR2_X1 U4573 ( .A1(n4163), .A2(n4161), .ZN(n4227) );
  NOR4_X1 U4574 ( .A1(n3816), .A2(n4227), .A3(n3815), .A4(n3814), .ZN(n3820)
         );
  NOR2_X1 U4575 ( .A1(n4248), .A2(n4607), .ZN(n3817) );
  AND4_X1 U4576 ( .A1(n3820), .A2(n3819), .A3(n3818), .A4(n3817), .ZN(n3821)
         );
  NAND4_X1 U4577 ( .A1(n3824), .A2(n3823), .A3(n3822), .A4(n3821), .ZN(n3846)
         );
  NOR2_X1 U4578 ( .A1(n3826), .A2(n3825), .ZN(n4083) );
  INV_X1 U4579 ( .A(n4083), .ZN(n3832) );
  INV_X1 U4580 ( .A(n3827), .ZN(n3831) );
  NAND2_X1 U4581 ( .A1(n3829), .A2(n3828), .ZN(n4187) );
  NOR4_X1 U4582 ( .A1(n3832), .A2(n3831), .A3(n4187), .A4(n3830), .ZN(n3844)
         );
  INV_X1 U4583 ( .A(n3833), .ZN(n3841) );
  NAND2_X1 U4584 ( .A1(n3050), .A2(n4622), .ZN(n3853) );
  INV_X1 U4585 ( .A(n3834), .ZN(n3835) );
  INV_X1 U4586 ( .A(n4268), .ZN(n3838) );
  INV_X1 U4587 ( .A(n4266), .ZN(n3837) );
  AOI21_X1 U4588 ( .B1(n3838), .B2(n3837), .A(n3836), .ZN(n3920) );
  XNOR2_X1 U4589 ( .A(n4069), .B(n4051), .ZN(n4049) );
  NAND4_X1 U4590 ( .A1(n3839), .A2(n4065), .A3(n3920), .A4(n4049), .ZN(n3840)
         );
  NOR4_X1 U4591 ( .A1(n3841), .A2(n4665), .A3(n4395), .A4(n3840), .ZN(n3842)
         );
  NAND3_X1 U4592 ( .A1(n3844), .A2(n3843), .A3(n3842), .ZN(n3845) );
  XNOR2_X1 U4593 ( .A(n4142), .B(n4177), .ZN(n4168) );
  NOR4_X1 U4594 ( .A1(n3846), .A2(n3845), .A3(n4124), .A4(n4168), .ZN(n3926)
         );
  INV_X1 U4595 ( .A(n3848), .ZN(n3849) );
  OAI211_X1 U4596 ( .C1(n3851), .C2(n2090), .A(n3850), .B(n3849), .ZN(n3898)
         );
  OAI211_X1 U4597 ( .C1(n4600), .C2(n4395), .A(n3853), .B(n3852), .ZN(n3856)
         );
  NAND3_X1 U4598 ( .A1(n3856), .A2(n3855), .A3(n3854), .ZN(n3858) );
  OAI211_X1 U4599 ( .C1(n3860), .C2(n3859), .A(n3858), .B(n3857), .ZN(n3863)
         );
  NAND3_X1 U4600 ( .A1(n3863), .A2(n3862), .A3(n3861), .ZN(n3866) );
  NAND4_X1 U4601 ( .A1(n3866), .A2(n3865), .A3(n3864), .A4(n3883), .ZN(n3868)
         );
  AND2_X1 U4602 ( .A1(n3868), .A2(n3867), .ZN(n3870) );
  INV_X1 U4603 ( .A(n3870), .ZN(n3872) );
  AOI21_X1 U4604 ( .B1(n3870), .B2(n3944), .A(n3869), .ZN(n3871) );
  AOI21_X1 U4605 ( .B1(n3873), .B2(n3872), .A(n3871), .ZN(n3877) );
  INV_X1 U4606 ( .A(n3884), .ZN(n3876) );
  OAI211_X1 U4607 ( .C1(n3877), .C2(n3876), .A(n3875), .B(n3874), .ZN(n3891)
         );
  NOR2_X1 U4608 ( .A1(n3879), .A2(n3878), .ZN(n3890) );
  INV_X1 U4609 ( .A(n3880), .ZN(n3882) );
  NOR2_X1 U4610 ( .A1(n3882), .A2(n3881), .ZN(n3886) );
  NAND4_X1 U4611 ( .A1(n3886), .A2(n3885), .A3(n3884), .A4(n3883), .ZN(n3888)
         );
  NAND2_X1 U4612 ( .A1(n3888), .A2(n3887), .ZN(n3889) );
  AOI22_X1 U4613 ( .A1(n3891), .A2(n3890), .B1(n3899), .B2(n3889), .ZN(n3896)
         );
  INV_X1 U4614 ( .A(n3892), .ZN(n3895) );
  INV_X1 U4615 ( .A(n3893), .ZN(n3894) );
  NOR4_X1 U4616 ( .A1(n3896), .A2(n3895), .A3(n3894), .A4(n2090), .ZN(n3897)
         );
  AOI21_X1 U4617 ( .B1(n3899), .B2(n3898), .A(n3897), .ZN(n3902) );
  INV_X1 U4618 ( .A(n3900), .ZN(n4159) );
  OAI21_X1 U4619 ( .B1(n3902), .B2(n4159), .A(n3901), .ZN(n3904) );
  NAND3_X1 U4620 ( .A1(n3904), .A2(n4164), .A3(n3903), .ZN(n3907) );
  AOI211_X1 U4621 ( .C1(n3907), .C2(n3906), .A(n2222), .B(n3905), .ZN(n3909)
         );
  NOR2_X1 U4622 ( .A1(n3909), .A2(n3908), .ZN(n3912) );
  OAI21_X1 U4623 ( .B1(n3912), .B2(n3911), .A(n3910), .ZN(n3914) );
  OAI221_X1 U4624 ( .B1(n3916), .B2(n3915), .C1(n3916), .C2(n3914), .A(n3913), 
        .ZN(n3917) );
  OR3_X1 U4625 ( .A1(n3919), .A2(n3918), .A3(n3917), .ZN(n3924) );
  INV_X1 U4626 ( .A(n3920), .ZN(n3921) );
  AOI22_X1 U4627 ( .A1(n3924), .A2(n3923), .B1(n3922), .B2(n3921), .ZN(n3925)
         );
  MUX2_X1 U4628 ( .A(n3926), .B(n3925), .S(n2360), .Z(n3927) );
  AOI21_X1 U4629 ( .B1(n3929), .B2(n3928), .A(n3927), .ZN(n3930) );
  XNOR2_X1 U4630 ( .A(n3930), .B(n2707), .ZN(n3936) );
  NAND2_X1 U4631 ( .A1(n3932), .A2(n3931), .ZN(n3933) );
  OAI211_X1 U4632 ( .C1(n4394), .C2(n3935), .A(n3933), .B(B_REG_SCAN_IN), .ZN(
        n3934) );
  OAI21_X1 U4633 ( .B1(n3936), .B2(n3935), .A(n3934), .ZN(U3239) );
  MUX2_X1 U4634 ( .A(n4266), .B(DATAO_REG_31__SCAN_IN), .S(n3938), .Z(U3581)
         );
  MUX2_X1 U4635 ( .A(n3937), .B(DATAO_REG_30__SCAN_IN), .S(n3938), .Z(U3580)
         );
  MUX2_X1 U4636 ( .A(DATAO_REG_28__SCAN_IN), .B(n4036), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4637 ( .A(n4052), .B(DATAO_REG_27__SCAN_IN), .S(n3938), .Z(U3577)
         );
  MUX2_X1 U4638 ( .A(n4069), .B(DATAO_REG_26__SCAN_IN), .S(n3938), .Z(U3576)
         );
  MUX2_X1 U4639 ( .A(DATAO_REG_25__SCAN_IN), .B(n4086), .S(U4043), .Z(U3575)
         );
  MUX2_X1 U4640 ( .A(n4110), .B(DATAO_REG_24__SCAN_IN), .S(n3938), .Z(U3574)
         );
  MUX2_X1 U4641 ( .A(n4126), .B(DATAO_REG_23__SCAN_IN), .S(n3938), .Z(U3573)
         );
  MUX2_X1 U4642 ( .A(DATAO_REG_20__SCAN_IN), .B(n4142), .S(U4043), .Z(U3570)
         );
  MUX2_X1 U4643 ( .A(DATAO_REG_19__SCAN_IN), .B(n4205), .S(U4043), .Z(U3569)
         );
  MUX2_X1 U4644 ( .A(DATAO_REG_18__SCAN_IN), .B(n4191), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4645 ( .A(DATAO_REG_17__SCAN_IN), .B(n3939), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U4646 ( .A(DATAO_REG_15__SCAN_IN), .B(n3940), .S(U4043), .Z(U3565)
         );
  MUX2_X1 U4647 ( .A(DATAO_REG_13__SCAN_IN), .B(n3941), .S(U4043), .Z(U3563)
         );
  MUX2_X1 U4648 ( .A(DATAO_REG_12__SCAN_IN), .B(n4582), .S(U4043), .Z(U3562)
         );
  MUX2_X1 U4649 ( .A(DATAO_REG_11__SCAN_IN), .B(n3942), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4650 ( .A(DATAO_REG_10__SCAN_IN), .B(n4580), .S(U4043), .Z(U3560)
         );
  MUX2_X1 U4651 ( .A(DATAO_REG_8__SCAN_IN), .B(n3943), .S(U4043), .Z(U3558) );
  MUX2_X1 U4652 ( .A(DATAO_REG_7__SCAN_IN), .B(n3944), .S(U4043), .Z(U3557) );
  MUX2_X1 U4653 ( .A(DATAO_REG_6__SCAN_IN), .B(n3945), .S(U4043), .Z(U3556) );
  MUX2_X1 U4654 ( .A(DATAO_REG_5__SCAN_IN), .B(n3946), .S(U4043), .Z(U3555) );
  MUX2_X1 U4655 ( .A(DATAO_REG_4__SCAN_IN), .B(n3947), .S(U4043), .Z(U3554) );
  MUX2_X1 U4656 ( .A(DATAO_REG_3__SCAN_IN), .B(n3948), .S(U4043), .Z(U3553) );
  MUX2_X1 U4657 ( .A(DATAO_REG_2__SCAN_IN), .B(n3054), .S(U4043), .Z(U3552) );
  MUX2_X1 U4658 ( .A(DATAO_REG_1__SCAN_IN), .B(n3049), .S(U4043), .Z(U3551) );
  MUX2_X1 U4659 ( .A(DATAO_REG_0__SCAN_IN), .B(n3050), .S(U4043), .Z(U3550) );
  OAI211_X1 U4660 ( .C1(n3961), .C2(n3949), .A(n4571), .B(n3974), .ZN(n3956)
         );
  OAI211_X1 U4661 ( .C1(n3951), .C2(n3950), .A(n4573), .B(n3965), .ZN(n3955)
         );
  AOI22_X1 U4662 ( .A1(n4563), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3954) );
  NAND2_X1 U4663 ( .A1(n4536), .A2(n2233), .ZN(n3953) );
  NAND4_X1 U4664 ( .A1(n3956), .A2(n3955), .A3(n3954), .A4(n3953), .ZN(U3241)
         );
  INV_X1 U4665 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4632) );
  NAND2_X1 U4666 ( .A1(n4438), .A2(n4632), .ZN(n3957) );
  NAND2_X1 U4667 ( .A1(n4391), .A2(n3957), .ZN(n4439) );
  INV_X1 U4668 ( .A(n4439), .ZN(n4437) );
  NAND2_X1 U4669 ( .A1(n3958), .A2(n3960), .ZN(n3959) );
  OAI211_X1 U4670 ( .C1(n3961), .C2(n3960), .A(n3959), .B(n4391), .ZN(n3963)
         );
  OAI211_X1 U4671 ( .C1(IR_REG_0__SCAN_IN), .C2(n4437), .A(n3963), .B(U4043), 
        .ZN(n4454) );
  AOI22_X1 U4672 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4563), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3980) );
  MUX2_X1 U4673 ( .A(REG1_REG_2__SCAN_IN), .B(n3245), .S(n3971), .Z(n3966) );
  NAND3_X1 U4674 ( .A1(n3966), .A2(n3965), .A3(n3964), .ZN(n3967) );
  NAND3_X1 U4675 ( .A1(n4573), .A2(n3968), .A3(n3967), .ZN(n3970) );
  NAND2_X1 U4676 ( .A1(n4536), .A2(n4400), .ZN(n3969) );
  AND2_X1 U4677 ( .A1(n3970), .A2(n3969), .ZN(n3979) );
  MUX2_X1 U4678 ( .A(REG2_REG_2__SCAN_IN), .B(n3972), .S(n3971), .Z(n3975) );
  NAND3_X1 U4679 ( .A1(n3975), .A2(n3974), .A3(n3973), .ZN(n3977) );
  NAND3_X1 U4680 ( .A1(n4571), .A2(n3977), .A3(n3976), .ZN(n3978) );
  NAND4_X1 U4681 ( .A1(n4454), .A2(n3980), .A3(n3979), .A4(n3978), .ZN(U3242)
         );
  INV_X1 U4682 ( .A(n4014), .ZN(n4398) );
  XNOR2_X1 U4683 ( .A(n4398), .B(REG2_REG_18__SCAN_IN), .ZN(n3990) );
  NOR2_X1 U4684 ( .A1(n4005), .A2(REG2_REG_17__SCAN_IN), .ZN(n3981) );
  AOI21_X1 U4685 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4005), .A(n3981), .ZN(n4569) );
  INV_X1 U4686 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4521) );
  INV_X1 U4687 ( .A(n3999), .ZN(n4651) );
  NOR2_X1 U4688 ( .A1(n4521), .A2(n4651), .ZN(n4520) );
  NAND2_X1 U4689 ( .A1(n3996), .A2(n3983), .ZN(n3984) );
  OAI22_X1 U4690 ( .A1(n4520), .A2(n4523), .B1(REG2_REG_13__SCAN_IN), .B2(
        n3999), .ZN(n3985) );
  NOR2_X1 U4691 ( .A1(n4649), .A2(n3985), .ZN(n3986) );
  XNOR2_X1 U4692 ( .A(n4649), .B(n3985), .ZN(n4532) );
  NOR2_X1 U4693 ( .A1(n3559), .A2(n4532), .ZN(n4531) );
  NOR2_X1 U4694 ( .A1(n3986), .A2(n4531), .ZN(n4546) );
  INV_X1 U4695 ( .A(n4646), .ZN(n4551) );
  AOI22_X1 U4696 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4551), .B1(n4646), .B2(
        n4257), .ZN(n4547) );
  NOR2_X1 U4697 ( .A1(n4546), .A2(n4547), .ZN(n4545) );
  NAND2_X1 U4698 ( .A1(n3987), .A2(n4645), .ZN(n3988) );
  NAND2_X1 U4699 ( .A1(n4569), .A2(n4568), .ZN(n4567) );
  OAI21_X1 U4700 ( .B1(n4005), .B2(REG2_REG_17__SCAN_IN), .A(n4567), .ZN(n3989) );
  NOR2_X1 U4701 ( .A1(n3989), .A2(n3990), .ZN(n4018) );
  AOI21_X1 U4702 ( .B1(n3990), .B2(n3989), .A(n4018), .ZN(n3991) );
  NAND2_X1 U4703 ( .A1(n4571), .A2(n3991), .ZN(n4013) );
  AOI22_X1 U4704 ( .A1(n4005), .A2(REG1_REG_17__SCAN_IN), .B1(n4326), .B2(
        n4643), .ZN(n4566) );
  NAND2_X1 U4705 ( .A1(n2107), .A2(REG1_REG_11__SCAN_IN), .ZN(n3993) );
  NOR2_X1 U4706 ( .A1(n3995), .A2(n2105), .ZN(n3997) );
  XOR2_X1 U4707 ( .A(n3996), .B(n3995), .Z(n4507) );
  NOR2_X1 U4708 ( .A1(n2597), .A2(n4507), .ZN(n4506) );
  AOI22_X1 U4709 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4651), .B1(n3999), .B2(
        n3998), .ZN(n4516) );
  NOR2_X1 U4710 ( .A1(n4517), .A2(n4516), .ZN(n4515) );
  NOR2_X1 U4711 ( .A1(n4000), .A2(n4649), .ZN(n4001) );
  AOI22_X1 U4712 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4551), .B1(n4646), .B2(
        n4002), .ZN(n4542) );
  NAND2_X1 U4713 ( .A1(n4003), .A2(n4645), .ZN(n4004) );
  XOR2_X1 U4714 ( .A(n4645), .B(n4003), .Z(n4555) );
  NAND2_X1 U4715 ( .A1(n4555), .A2(n4554), .ZN(n4553) );
  NAND2_X1 U4716 ( .A1(n4004), .A2(n4553), .ZN(n4565) );
  NAND2_X1 U4717 ( .A1(n4566), .A2(n4565), .ZN(n4564) );
  OR2_X1 U4718 ( .A1(n4014), .A2(n4006), .ZN(n4015) );
  OAI21_X1 U4719 ( .B1(n4398), .B2(REG1_REG_18__SCAN_IN), .A(n4015), .ZN(n4007) );
  NAND2_X1 U4720 ( .A1(n4563), .A2(ADDR_REG_18__SCAN_IN), .ZN(n4009) );
  OAI211_X1 U4721 ( .C1(n4014), .C2(n4576), .A(n4013), .B(n4012), .ZN(U3258)
         );
  INV_X1 U4722 ( .A(n4015), .ZN(n4016) );
  XNOR2_X1 U4723 ( .A(n2707), .B(n4318), .ZN(n4017) );
  AOI21_X1 U4724 ( .B1(REG2_REG_18__SCAN_IN), .B2(n4398), .A(n4018), .ZN(n4021) );
  INV_X1 U4725 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4019) );
  MUX2_X1 U4726 ( .A(n4019), .B(REG2_REG_19__SCAN_IN), .S(n2707), .Z(n4020) );
  XNOR2_X1 U4727 ( .A(n4021), .B(n4020), .ZN(n4025) );
  NAND2_X1 U4728 ( .A1(n4563), .A2(ADDR_REG_19__SCAN_IN), .ZN(n4022) );
  OAI211_X1 U4729 ( .C1(n4576), .C2(n2707), .A(n4023), .B(n4022), .ZN(n4024)
         );
  AOI21_X1 U4730 ( .B1(n4025), .B2(n4571), .A(n4024), .ZN(n4026) );
  OAI21_X1 U4731 ( .B1(n4027), .B2(n4540), .A(n4026), .ZN(U3259) );
  XNOR2_X1 U4732 ( .A(n4028), .B(n4031), .ZN(n4283) );
  INV_X1 U4733 ( .A(n4283), .ZN(n4044) );
  OAI22_X1 U4734 ( .A1(n4029), .A2(n4207), .B1(n4038), .B2(n4267), .ZN(n4035)
         );
  AOI21_X1 U4735 ( .B1(n4032), .B2(n4031), .A(n4030), .ZN(n4033) );
  NOR2_X1 U4736 ( .A1(n4033), .A2(n4585), .ZN(n4034) );
  INV_X1 U4737 ( .A(n4284), .ZN(n4042) );
  OAI21_X1 U4738 ( .B1(n4056), .B2(n4038), .A(n4037), .ZN(n4286) );
  AOI22_X1 U4739 ( .A1(n4039), .A2(n4629), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4634), .ZN(n4040) );
  OAI21_X1 U4740 ( .B1(n4286), .B2(n4235), .A(n4040), .ZN(n4041) );
  AOI21_X1 U4741 ( .B1(n4042), .B2(n3379), .A(n4041), .ZN(n4043) );
  OAI21_X1 U4742 ( .B1(n4044), .B2(n4262), .A(n4043), .ZN(U3263) );
  XOR2_X1 U4743 ( .A(n4049), .B(n4045), .Z(n4288) );
  INV_X1 U4744 ( .A(n4288), .ZN(n4063) );
  INV_X1 U4745 ( .A(n4046), .ZN(n4047) );
  NOR2_X1 U4746 ( .A1(n4048), .A2(n4047), .ZN(n4050) );
  XNOR2_X1 U4747 ( .A(n4050), .B(n4049), .ZN(n4055) );
  AOI22_X1 U4748 ( .A1(n4086), .A2(n4603), .B1(n4051), .B2(n4602), .ZN(n4054)
         );
  NAND2_X1 U4749 ( .A1(n4052), .A2(n4581), .ZN(n4053) );
  OAI211_X1 U4750 ( .C1(n4055), .C2(n4585), .A(n4054), .B(n4053), .ZN(n4287)
         );
  INV_X1 U4751 ( .A(n4056), .ZN(n4057) );
  OAI21_X1 U4752 ( .B1(n4074), .B2(n4058), .A(n4057), .ZN(n4356) );
  AOI22_X1 U4753 ( .A1(n4059), .A2(n4629), .B1(n4634), .B2(
        REG2_REG_26__SCAN_IN), .ZN(n4060) );
  OAI21_X1 U4754 ( .B1(n4356), .B2(n4235), .A(n4060), .ZN(n4061) );
  AOI21_X1 U4755 ( .B1(n4287), .B2(n3379), .A(n4061), .ZN(n4062) );
  OAI21_X1 U4756 ( .B1(n4063), .B2(n4262), .A(n4062), .ZN(U3264) );
  XOR2_X1 U4757 ( .A(n4065), .B(n4064), .Z(n4292) );
  INV_X1 U4758 ( .A(n4292), .ZN(n4079) );
  XNOR2_X1 U4759 ( .A(n4066), .B(n4065), .ZN(n4071) );
  OAI22_X1 U4760 ( .A1(n4067), .A2(n4207), .B1(n4072), .B2(n4267), .ZN(n4068)
         );
  AOI21_X1 U4761 ( .B1(n4581), .B2(n4069), .A(n4068), .ZN(n4070) );
  OAI21_X1 U4762 ( .B1(n4071), .B2(n4585), .A(n4070), .ZN(n4291) );
  NOR2_X1 U4763 ( .A1(n4090), .A2(n4072), .ZN(n4073) );
  AOI22_X1 U4764 ( .A1(n4634), .A2(REG2_REG_25__SCAN_IN), .B1(n4075), .B2(
        n4629), .ZN(n4076) );
  OAI21_X1 U4765 ( .B1(n4360), .B2(n4235), .A(n4076), .ZN(n4077) );
  AOI21_X1 U4766 ( .B1(n4291), .B2(n3379), .A(n4077), .ZN(n4078) );
  OAI21_X1 U4767 ( .B1(n4079), .B2(n4262), .A(n4078), .ZN(U3265) );
  XNOR2_X1 U4768 ( .A(n4080), .B(n4083), .ZN(n4296) );
  INV_X1 U4769 ( .A(n4296), .ZN(n4099) );
  NOR2_X1 U4770 ( .A1(n4082), .A2(n4081), .ZN(n4084) );
  XNOR2_X1 U4771 ( .A(n4084), .B(n4083), .ZN(n4089) );
  AOI22_X1 U4772 ( .A1(n4126), .A2(n4603), .B1(n4085), .B2(n4602), .ZN(n4088)
         );
  NAND2_X1 U4773 ( .A1(n4086), .A2(n4581), .ZN(n4087) );
  OAI211_X1 U4774 ( .C1(n4089), .C2(n4585), .A(n4088), .B(n4087), .ZN(n4295)
         );
  INV_X1 U4775 ( .A(n4114), .ZN(n4093) );
  INV_X1 U4776 ( .A(n4090), .ZN(n4091) );
  OAI21_X1 U4777 ( .B1(n4093), .B2(n4092), .A(n4091), .ZN(n4364) );
  NOR2_X1 U4778 ( .A1(n4364), .A2(n4235), .ZN(n4097) );
  INV_X1 U4779 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4095) );
  OAI22_X1 U4780 ( .A1(n3379), .A2(n4095), .B1(n4094), .B2(n4255), .ZN(n4096)
         );
  AOI211_X1 U4781 ( .C1(n4295), .C2(n3379), .A(n4097), .B(n4096), .ZN(n4098)
         );
  OAI21_X1 U4782 ( .B1(n4099), .B2(n4262), .A(n4098), .ZN(U3266) );
  XNOR2_X1 U4783 ( .A(n4100), .B(n4101), .ZN(n4300) );
  INV_X1 U4784 ( .A(n4300), .ZN(n4121) );
  NAND2_X1 U4785 ( .A1(n4103), .A2(n4102), .ZN(n4141) );
  OR2_X1 U4786 ( .A1(n4141), .A2(n4149), .ZN(n4105) );
  OAI21_X1 U4787 ( .B1(n4125), .B2(n4124), .A(n4106), .ZN(n4108) );
  XNOR2_X1 U4788 ( .A(n4108), .B(n4107), .ZN(n4113) );
  NOR2_X1 U4789 ( .A1(n4115), .A2(n4267), .ZN(n4109) );
  AOI21_X1 U4790 ( .B1(n4110), .B2(n4581), .A(n4109), .ZN(n4112) );
  NAND2_X1 U4791 ( .A1(n4143), .A2(n4603), .ZN(n4111) );
  OAI211_X1 U4792 ( .C1(n4113), .C2(n4585), .A(n4112), .B(n4111), .ZN(n4299)
         );
  INV_X1 U4793 ( .A(n4304), .ZN(n4116) );
  OAI21_X1 U4794 ( .B1(n4116), .B2(n4115), .A(n4114), .ZN(n4368) );
  AOI22_X1 U4795 ( .A1(n4634), .A2(REG2_REG_23__SCAN_IN), .B1(n4117), .B2(
        n4629), .ZN(n4118) );
  OAI21_X1 U4796 ( .B1(n4368), .B2(n4235), .A(n4118), .ZN(n4119) );
  AOI21_X1 U4797 ( .B1(n4299), .B2(n3379), .A(n4119), .ZN(n4120) );
  OAI21_X1 U4798 ( .B1(n4121), .B2(n4262), .A(n4120), .ZN(U3267) );
  OAI21_X1 U4799 ( .B1(n4123), .B2(n4124), .A(n4122), .ZN(n4307) );
  XNOR2_X1 U4800 ( .A(n4125), .B(n4124), .ZN(n4131) );
  NAND2_X1 U4801 ( .A1(n4171), .A2(n4603), .ZN(n4128) );
  NAND2_X1 U4802 ( .A1(n4126), .A2(n4581), .ZN(n4127) );
  OAI211_X1 U4803 ( .C1(n4267), .C2(n4129), .A(n4128), .B(n4127), .ZN(n4130)
         );
  AOI21_X1 U4804 ( .B1(n4131), .B2(n4624), .A(n4130), .ZN(n4306) );
  INV_X1 U4805 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4134) );
  INV_X1 U4806 ( .A(n4132), .ZN(n4133) );
  OAI22_X1 U4807 ( .A1(n3379), .A2(n4134), .B1(n4133), .B2(n4255), .ZN(n4135)
         );
  INV_X1 U4808 ( .A(n4135), .ZN(n4138) );
  NAND2_X1 U4809 ( .A1(n4150), .A2(n4136), .ZN(n4303) );
  NAND3_X1 U4810 ( .A1(n4304), .A2(n4617), .A3(n4303), .ZN(n4137) );
  OAI211_X1 U4811 ( .C1(n4306), .C2(n4634), .A(n4138), .B(n4137), .ZN(n4139)
         );
  INV_X1 U4812 ( .A(n4139), .ZN(n4140) );
  OAI21_X1 U4813 ( .B1(n4307), .B2(n4262), .A(n4140), .ZN(U3268) );
  XNOR2_X1 U4814 ( .A(n4141), .B(n4149), .ZN(n4147) );
  NAND2_X1 U4815 ( .A1(n4142), .A2(n4603), .ZN(n4145) );
  NAND2_X1 U4816 ( .A1(n4143), .A2(n4581), .ZN(n4144) );
  OAI211_X1 U4817 ( .C1(n4267), .C2(n4151), .A(n4145), .B(n4144), .ZN(n4146)
         );
  AOI21_X1 U4818 ( .B1(n4147), .B2(n4624), .A(n4146), .ZN(n4309) );
  XNOR2_X1 U4819 ( .A(n4148), .B(n4149), .ZN(n4308) );
  NAND2_X1 U4820 ( .A1(n4308), .A2(n4237), .ZN(n4157) );
  OAI21_X1 U4821 ( .B1(n4175), .B2(n4151), .A(n4150), .ZN(n4311) );
  INV_X1 U4822 ( .A(n4311), .ZN(n4155) );
  INV_X1 U4823 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4153) );
  OAI22_X1 U4824 ( .A1(n3379), .A2(n4153), .B1(n4152), .B2(n4255), .ZN(n4154)
         );
  AOI21_X1 U4825 ( .B1(n4155), .B2(n4617), .A(n4154), .ZN(n4156) );
  OAI211_X1 U4826 ( .C1(n4634), .C2(n4309), .A(n4157), .B(n4156), .ZN(U3269)
         );
  XOR2_X1 U4827 ( .A(n4168), .B(n4158), .Z(n4313) );
  INV_X1 U4828 ( .A(n4313), .ZN(n4182) );
  INV_X1 U4829 ( .A(n4161), .ZN(n4162) );
  OAI21_X1 U4830 ( .B1(n4221), .B2(n4163), .A(n4162), .ZN(n4203) );
  NAND2_X1 U4831 ( .A1(n4203), .A2(n4164), .ZN(n4167) );
  INV_X1 U4832 ( .A(n4165), .ZN(n4166) );
  NAND2_X1 U4833 ( .A1(n4167), .A2(n4166), .ZN(n4169) );
  XNOR2_X1 U4834 ( .A(n4169), .B(n4168), .ZN(n4174) );
  NOR2_X1 U4835 ( .A1(n4177), .A2(n4267), .ZN(n4170) );
  AOI21_X1 U4836 ( .B1(n4171), .B2(n4581), .A(n4170), .ZN(n4173) );
  NAND2_X1 U4837 ( .A1(n4205), .A2(n4603), .ZN(n4172) );
  OAI211_X1 U4838 ( .C1(n4174), .C2(n4585), .A(n4173), .B(n4172), .ZN(n4312)
         );
  INV_X1 U4839 ( .A(n4175), .ZN(n4176) );
  OAI21_X1 U4840 ( .B1(n4194), .B2(n4177), .A(n4176), .ZN(n4374) );
  AOI22_X1 U4841 ( .A1(n4634), .A2(REG2_REG_20__SCAN_IN), .B1(n4178), .B2(
        n4629), .ZN(n4179) );
  OAI21_X1 U4842 ( .B1(n4374), .B2(n4235), .A(n4179), .ZN(n4180) );
  AOI21_X1 U4843 ( .B1(n4312), .B2(n3379), .A(n4180), .ZN(n4181) );
  OAI21_X1 U4844 ( .B1(n4182), .B2(n4262), .A(n4181), .ZN(U3270) );
  XNOR2_X1 U4845 ( .A(n4183), .B(n4187), .ZN(n4317) );
  INV_X1 U4846 ( .A(n4317), .ZN(n4202) );
  OAI21_X1 U4847 ( .B1(n4203), .B2(n4185), .A(n4184), .ZN(n4186) );
  XOR2_X1 U4848 ( .A(n4187), .B(n4186), .Z(n4193) );
  OAI22_X1 U4849 ( .A1(n4189), .A2(n4627), .B1(n4267), .B2(n4188), .ZN(n4190)
         );
  AOI21_X1 U4850 ( .B1(n4603), .B2(n4191), .A(n4190), .ZN(n4192) );
  OAI21_X1 U4851 ( .B1(n4193), .B2(n4585), .A(n4192), .ZN(n4316) );
  INV_X1 U4852 ( .A(n4194), .ZN(n4197) );
  OAI21_X1 U4853 ( .B1(n4232), .B2(n4204), .A(n4195), .ZN(n4196) );
  NAND2_X1 U4854 ( .A1(n4197), .A2(n4196), .ZN(n4379) );
  NOR2_X1 U4855 ( .A1(n4379), .A2(n4235), .ZN(n4200) );
  OAI22_X1 U4856 ( .A1(n3379), .A2(n4019), .B1(n4198), .B2(n4255), .ZN(n4199)
         );
  AOI211_X1 U4857 ( .C1(n4316), .C2(n3379), .A(n4200), .B(n4199), .ZN(n4201)
         );
  OAI21_X1 U4858 ( .B1(n4202), .B2(n4262), .A(n4201), .ZN(U3271) );
  XOR2_X1 U4859 ( .A(n4211), .B(n4203), .Z(n4209) );
  AOI22_X1 U4860 ( .A1(n4205), .A2(n4581), .B1(n4204), .B2(n4602), .ZN(n4206)
         );
  OAI21_X1 U4861 ( .B1(n4412), .B2(n4207), .A(n4206), .ZN(n4208) );
  AOI21_X1 U4862 ( .B1(n4209), .B2(n4624), .A(n4208), .ZN(n4322) );
  OAI21_X1 U4863 ( .B1(n4212), .B2(n4211), .A(n4210), .ZN(n4320) );
  XNOR2_X1 U4864 ( .A(n4232), .B(n4213), .ZN(n4214) );
  NAND2_X1 U4865 ( .A1(n4214), .A2(n4715), .ZN(n4321) );
  INV_X1 U4866 ( .A(n4215), .ZN(n4218) );
  AOI22_X1 U4867 ( .A1(n4634), .A2(REG2_REG_18__SCAN_IN), .B1(n4216), .B2(
        n4629), .ZN(n4217) );
  OAI21_X1 U4868 ( .B1(n4321), .B2(n4218), .A(n4217), .ZN(n4219) );
  AOI21_X1 U4869 ( .B1(n4320), .B2(n4237), .A(n4219), .ZN(n4220) );
  OAI21_X1 U4870 ( .B1(n4634), .B2(n4322), .A(n4220), .ZN(U3272) );
  XOR2_X1 U4871 ( .A(n4227), .B(n4221), .Z(n4226) );
  OAI22_X1 U4872 ( .A1(n3076), .A2(n4627), .B1(n4267), .B2(n4222), .ZN(n4223)
         );
  AOI21_X1 U4873 ( .B1(n4603), .B2(n4224), .A(n4223), .ZN(n4225) );
  OAI21_X1 U4874 ( .B1(n4226), .B2(n4585), .A(n4225), .ZN(n4324) );
  INV_X1 U4875 ( .A(n4324), .ZN(n4239) );
  XNOR2_X1 U4876 ( .A(n4228), .B(n4227), .ZN(n4325) );
  NAND2_X1 U4877 ( .A1(n4230), .A2(n4229), .ZN(n4231) );
  NAND2_X1 U4878 ( .A1(n4232), .A2(n4231), .ZN(n4385) );
  AOI22_X1 U4879 ( .A1(n4634), .A2(REG2_REG_17__SCAN_IN), .B1(n4233), .B2(
        n4629), .ZN(n4234) );
  OAI21_X1 U4880 ( .B1(n4385), .B2(n4235), .A(n4234), .ZN(n4236) );
  AOI21_X1 U4881 ( .B1(n4325), .B2(n4237), .A(n4236), .ZN(n4238) );
  OAI21_X1 U4882 ( .B1(n4634), .B2(n4239), .A(n4238), .ZN(U3273) );
  INV_X1 U4883 ( .A(n4240), .ZN(n4242) );
  NAND2_X1 U4884 ( .A1(n4242), .A2(n4241), .ZN(n4243) );
  XOR2_X1 U4885 ( .A(n4248), .B(n4243), .Z(n4338) );
  OAI22_X1 U4886 ( .A1(n4245), .A2(n4627), .B1(n4244), .B2(n4267), .ZN(n4251)
         );
  INV_X1 U4887 ( .A(n4246), .ZN(n4247) );
  AOI211_X1 U4888 ( .C1(n4249), .C2(n4248), .A(n4585), .B(n4247), .ZN(n4250)
         );
  AOI211_X1 U4889 ( .C1(n4603), .C2(n4252), .A(n4251), .B(n4250), .ZN(n4336)
         );
  INV_X1 U4890 ( .A(n4336), .ZN(n4260) );
  INV_X1 U4891 ( .A(n4253), .ZN(n4334) );
  NAND2_X1 U4892 ( .A1(n4340), .A2(n4254), .ZN(n4333) );
  AND3_X1 U4893 ( .A1(n4334), .A2(n4617), .A3(n4333), .ZN(n4259) );
  INV_X1 U4894 ( .A(REG2_REG_15__SCAN_IN), .ZN(n4257) );
  OAI22_X1 U4895 ( .A1(n3379), .A2(n4257), .B1(n4256), .B2(n4255), .ZN(n4258)
         );
  AOI211_X1 U4896 ( .C1(n4260), .C2(n3379), .A(n4259), .B(n4258), .ZN(n4261)
         );
  OAI21_X1 U4897 ( .B1(n4338), .B2(n4262), .A(n4261), .ZN(U3275) );
  XNOR2_X1 U4898 ( .A(n4272), .B(n4268), .ZN(n4431) );
  NAND2_X1 U4899 ( .A1(n4431), .A2(n4264), .ZN(n4270) );
  NAND2_X1 U4900 ( .A1(n4266), .A2(n4265), .ZN(n4275) );
  OAI21_X1 U4901 ( .B1(n4268), .B2(n4267), .A(n4275), .ZN(n4430) );
  NAND2_X1 U4902 ( .A1(n4735), .A2(n4430), .ZN(n4269) );
  OAI211_X1 U4903 ( .C1(n4735), .C2(n3785), .A(n4270), .B(n4269), .ZN(U3549)
         );
  INV_X1 U4904 ( .A(n4271), .ZN(n4274) );
  INV_X1 U4905 ( .A(n4272), .ZN(n4273) );
  AOI21_X1 U4906 ( .B1(n4277), .B2(n4274), .A(n4273), .ZN(n4434) );
  INV_X1 U4907 ( .A(n4434), .ZN(n4350) );
  INV_X1 U4908 ( .A(n4275), .ZN(n4276) );
  AOI21_X1 U4909 ( .B1(n4277), .B2(n4602), .A(n4276), .ZN(n4436) );
  MUX2_X1 U4910 ( .A(n4278), .B(n4436), .S(n4735), .Z(n4279) );
  OAI21_X1 U4911 ( .B1(n4350), .B2(n4328), .A(n4279), .ZN(U3548) );
  NAND2_X1 U4912 ( .A1(n4283), .A2(n4704), .ZN(n4285) );
  OAI211_X1 U4913 ( .C1(n4701), .C2(n4286), .A(n4285), .B(n4284), .ZN(n4352)
         );
  MUX2_X1 U4914 ( .A(REG1_REG_27__SCAN_IN), .B(n4352), .S(n4735), .Z(U3545) );
  AOI21_X1 U4915 ( .B1(n4288), .B2(n4704), .A(n4287), .ZN(n4353) );
  MUX2_X1 U4916 ( .A(n4289), .B(n4353), .S(n4735), .Z(n4290) );
  OAI21_X1 U4917 ( .B1(n4328), .B2(n4356), .A(n4290), .ZN(U3544) );
  INV_X1 U4918 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4293) );
  AOI21_X1 U4919 ( .B1(n4292), .B2(n4704), .A(n4291), .ZN(n4357) );
  MUX2_X1 U4920 ( .A(n4293), .B(n4357), .S(n4735), .Z(n4294) );
  OAI21_X1 U4921 ( .B1(n4328), .B2(n4360), .A(n4294), .ZN(U3543) );
  INV_X1 U4922 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4297) );
  AOI21_X1 U4923 ( .B1(n4296), .B2(n4704), .A(n4295), .ZN(n4361) );
  MUX2_X1 U4924 ( .A(n4297), .B(n4361), .S(n4735), .Z(n4298) );
  OAI21_X1 U4925 ( .B1(n4328), .B2(n4364), .A(n4298), .ZN(U3542) );
  AOI21_X1 U4926 ( .B1(n4300), .B2(n4704), .A(n4299), .ZN(n4365) );
  MUX2_X1 U4927 ( .A(n4301), .B(n4365), .S(n4735), .Z(n4302) );
  OAI21_X1 U4928 ( .B1(n4328), .B2(n4368), .A(n4302), .ZN(U3541) );
  NAND3_X1 U4929 ( .A1(n4304), .A2(n4715), .A3(n4303), .ZN(n4305) );
  OAI211_X1 U4930 ( .C1(n4307), .C2(n4337), .A(n4306), .B(n4305), .ZN(n4369)
         );
  MUX2_X1 U4931 ( .A(REG1_REG_22__SCAN_IN), .B(n4369), .S(n4735), .Z(U3540) );
  NAND2_X1 U4932 ( .A1(n4308), .A2(n4704), .ZN(n4310) );
  OAI211_X1 U4933 ( .C1(n4701), .C2(n4311), .A(n4310), .B(n4309), .ZN(n4370)
         );
  MUX2_X1 U4934 ( .A(REG1_REG_21__SCAN_IN), .B(n4370), .S(n4735), .Z(U3539) );
  AOI21_X1 U4935 ( .B1(n4313), .B2(n4704), .A(n4312), .ZN(n4371) );
  MUX2_X1 U4936 ( .A(n4314), .B(n4371), .S(n4735), .Z(n4315) );
  OAI21_X1 U4937 ( .B1(n4328), .B2(n4374), .A(n4315), .ZN(U3538) );
  AOI21_X1 U4938 ( .B1(n4317), .B2(n4704), .A(n4316), .ZN(n4376) );
  MUX2_X1 U4939 ( .A(n4318), .B(n4376), .S(n4735), .Z(n4319) );
  OAI21_X1 U4940 ( .B1(n4328), .B2(n4379), .A(n4319), .ZN(U3537) );
  INV_X1 U4941 ( .A(n4320), .ZN(n4323) );
  OAI211_X1 U4942 ( .C1(n4323), .C2(n4337), .A(n4322), .B(n4321), .ZN(n4380)
         );
  MUX2_X1 U4943 ( .A(REG1_REG_18__SCAN_IN), .B(n4380), .S(n4735), .Z(U3536) );
  AOI21_X1 U4944 ( .B1(n4325), .B2(n4704), .A(n4324), .ZN(n4381) );
  MUX2_X1 U4945 ( .A(n4326), .B(n4381), .S(n4735), .Z(n4327) );
  OAI21_X1 U4946 ( .B1(n4328), .B2(n4385), .A(n4327), .ZN(U3535) );
  NAND2_X1 U4947 ( .A1(n4329), .A2(n4704), .ZN(n4330) );
  OAI211_X1 U4948 ( .C1(n4701), .C2(n4332), .A(n4331), .B(n4330), .ZN(n4386)
         );
  MUX2_X1 U4949 ( .A(REG1_REG_16__SCAN_IN), .B(n4386), .S(n4735), .Z(U3534) );
  NAND3_X1 U4950 ( .A1(n4334), .A2(n4715), .A3(n4333), .ZN(n4335) );
  OAI211_X1 U4951 ( .C1(n4338), .C2(n4337), .A(n4336), .B(n4335), .ZN(n4387)
         );
  MUX2_X1 U4952 ( .A(REG1_REG_15__SCAN_IN), .B(n4387), .S(n4735), .Z(U3533) );
  NAND3_X1 U4953 ( .A1(n4340), .A2(n4715), .A3(n4339), .ZN(n4341) );
  OAI211_X1 U4954 ( .C1(n4343), .C2(n4679), .A(n4342), .B(n4341), .ZN(n4388)
         );
  MUX2_X1 U4955 ( .A(REG1_REG_14__SCAN_IN), .B(n4388), .S(n4735), .Z(U3532) );
  INV_X1 U4956 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4347) );
  NAND2_X1 U4957 ( .A1(n4431), .A2(n4344), .ZN(n4346) );
  NAND2_X1 U4958 ( .A1(n4375), .A2(n4430), .ZN(n4345) );
  OAI211_X1 U4959 ( .C1(n4375), .C2(n4347), .A(n4346), .B(n4345), .ZN(U3517)
         );
  MUX2_X1 U4960 ( .A(n4348), .B(n4436), .S(n4375), .Z(n4349) );
  OAI21_X1 U4961 ( .B1(n4350), .B2(n4384), .A(n4349), .ZN(U3516) );
  MUX2_X1 U4962 ( .A(REG0_REG_27__SCAN_IN), .B(n4352), .S(n4375), .Z(U3513) );
  INV_X1 U4963 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4354) );
  MUX2_X1 U4964 ( .A(n4354), .B(n4353), .S(n4375), .Z(n4355) );
  OAI21_X1 U4965 ( .B1(n4356), .B2(n4384), .A(n4355), .ZN(U3512) );
  INV_X1 U4966 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4358) );
  MUX2_X1 U4967 ( .A(n4358), .B(n4357), .S(n4375), .Z(n4359) );
  OAI21_X1 U4968 ( .B1(n4360), .B2(n4384), .A(n4359), .ZN(U3511) );
  INV_X1 U4969 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4362) );
  MUX2_X1 U4970 ( .A(n4362), .B(n4361), .S(n4375), .Z(n4363) );
  OAI21_X1 U4971 ( .B1(n4364), .B2(n4384), .A(n4363), .ZN(U3510) );
  MUX2_X1 U4972 ( .A(n4366), .B(n4365), .S(n4375), .Z(n4367) );
  OAI21_X1 U4973 ( .B1(n4368), .B2(n4384), .A(n4367), .ZN(U3509) );
  MUX2_X1 U4974 ( .A(REG0_REG_22__SCAN_IN), .B(n4369), .S(n4375), .Z(U3508) );
  MUX2_X1 U4975 ( .A(REG0_REG_21__SCAN_IN), .B(n4370), .S(n4375), .Z(U3507) );
  INV_X1 U4976 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4372) );
  MUX2_X1 U4977 ( .A(n4372), .B(n4371), .S(n4375), .Z(n4373) );
  OAI21_X1 U4978 ( .B1(n4374), .B2(n4384), .A(n4373), .ZN(U3506) );
  MUX2_X1 U4979 ( .A(n4377), .B(n4376), .S(n4375), .Z(n4378) );
  OAI21_X1 U4980 ( .B1(n4379), .B2(n4384), .A(n4378), .ZN(U3505) );
  MUX2_X1 U4981 ( .A(REG0_REG_18__SCAN_IN), .B(n4380), .S(n4722), .Z(U3503) );
  INV_X1 U4982 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4382) );
  MUX2_X1 U4983 ( .A(n4382), .B(n4381), .S(n4722), .Z(n4383) );
  OAI21_X1 U4984 ( .B1(n4385), .B2(n4384), .A(n4383), .ZN(U3501) );
  MUX2_X1 U4985 ( .A(REG0_REG_16__SCAN_IN), .B(n4386), .S(n4722), .Z(U3499) );
  MUX2_X1 U4986 ( .A(REG0_REG_15__SCAN_IN), .B(n4387), .S(n4722), .Z(U3497) );
  MUX2_X1 U4987 ( .A(REG0_REG_14__SCAN_IN), .B(n4388), .S(n4722), .Z(U3495) );
  MUX2_X1 U4988 ( .A(n4389), .B(DATAI_30_), .S(U3149), .Z(U3322) );
  MUX2_X1 U4989 ( .A(DATAI_29_), .B(n4390), .S(STATE_REG_SCAN_IN), .Z(U3323)
         );
  MUX2_X1 U4990 ( .A(DATAI_28_), .B(n4391), .S(STATE_REG_SCAN_IN), .Z(U3324)
         );
  MUX2_X1 U4991 ( .A(n4438), .B(DATAI_27_), .S(U3149), .Z(U3325) );
  MUX2_X1 U4992 ( .A(DATAI_26_), .B(n4392), .S(STATE_REG_SCAN_IN), .Z(U3326)
         );
  MUX2_X1 U4993 ( .A(DATAI_24_), .B(n4393), .S(STATE_REG_SCAN_IN), .Z(U3328)
         );
  MUX2_X1 U4994 ( .A(DATAI_22_), .B(n4394), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U4995 ( .A(DATAI_21_), .B(n4395), .S(STATE_REG_SCAN_IN), .Z(U3331)
         );
  MUX2_X1 U4996 ( .A(DATAI_20_), .B(n4396), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U4997 ( .A(n4397), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U4998 ( .A(n4398), .B(DATAI_18_), .S(U3149), .Z(U3334) );
  MUX2_X1 U4999 ( .A(n2107), .B(DATAI_11_), .S(U3149), .Z(U3341) );
  MUX2_X1 U5000 ( .A(DATAI_9_), .B(n4399), .S(STATE_REG_SCAN_IN), .Z(U3343) );
  MUX2_X1 U5001 ( .A(DATAI_4_), .B(n4444), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5002 ( .A(n4406), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U5003 ( .A(n4400), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5004 ( .A(n2233), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  AOI21_X1 U5005 ( .B1(n4563), .B2(ADDR_REG_3__SCAN_IN), .A(n4401), .ZN(n4410)
         );
  OAI211_X1 U5006 ( .C1(REG1_REG_3__SCAN_IN), .C2(n4403), .A(n4573), .B(n4402), 
        .ZN(n4409) );
  OAI211_X1 U5007 ( .C1(REG2_REG_3__SCAN_IN), .C2(n4405), .A(n4571), .B(n4404), 
        .ZN(n4408) );
  NAND2_X1 U5008 ( .A1(n4536), .A2(n4406), .ZN(n4407) );
  NAND4_X1 U5009 ( .A1(n4410), .A2(n4409), .A3(n4408), .A4(n4407), .ZN(U3243)
         );
  NOR2_X1 U5010 ( .A1(STATE_REG_SCAN_IN), .A2(n4411), .ZN(n4552) );
  OAI22_X1 U5011 ( .A1(n4415), .A2(n4414), .B1(n4413), .B2(n4412), .ZN(n4416)
         );
  AOI211_X1 U5012 ( .C1(n4418), .C2(n4417), .A(n4552), .B(n4416), .ZN(n4427)
         );
  AOI21_X1 U5013 ( .B1(n4421), .B2(n4420), .A(n4419), .ZN(n4422) );
  XOR2_X1 U5014 ( .A(n4423), .B(n4422), .Z(n4425) );
  NAND2_X1 U5015 ( .A1(n4425), .A2(n4424), .ZN(n4426) );
  OAI211_X1 U5016 ( .C1(n4429), .C2(n4428), .A(n4427), .B(n4426), .ZN(U3223)
         );
  AOI22_X1 U5017 ( .A1(n4431), .A2(n4617), .B1(n3379), .B2(n4430), .ZN(n4432)
         );
  OAI21_X1 U5018 ( .B1(n3379), .B2(n4433), .A(n4432), .ZN(U3260) );
  AOI22_X1 U5019 ( .A1(n4434), .A2(n4617), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4634), .ZN(n4435) );
  OAI21_X1 U5020 ( .B1(n4634), .B2(n4436), .A(n4435), .ZN(U3261) );
  OAI211_X1 U5021 ( .C1(REG1_REG_0__SCAN_IN), .C2(n4438), .A(n4440), .B(n4437), 
        .ZN(n4443) );
  AOI22_X1 U5022 ( .A1(n4440), .A2(n4439), .B1(n4573), .B2(n4723), .ZN(n4442)
         );
  AOI22_X1 U5023 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4563), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4441) );
  OAI221_X1 U5024 ( .B1(IR_REG_0__SCAN_IN), .B2(n4443), .C1(n2377), .C2(n4442), 
        .A(n4441), .ZN(U3240) );
  NAND2_X1 U5025 ( .A1(n4536), .A2(n4444), .ZN(n4453) );
  XNOR2_X1 U5026 ( .A(n4445), .B(REG2_REG_4__SCAN_IN), .ZN(n4446) );
  NAND2_X1 U5027 ( .A1(n4571), .A2(n4446), .ZN(n4452) );
  XNOR2_X1 U5028 ( .A(n4447), .B(REG1_REG_4__SCAN_IN), .ZN(n4448) );
  NAND2_X1 U5029 ( .A1(n4573), .A2(n4448), .ZN(n4451) );
  AOI21_X1 U5030 ( .B1(n4563), .B2(ADDR_REG_4__SCAN_IN), .A(n4449), .ZN(n4450)
         );
  AND4_X1 U5031 ( .A1(n4453), .A2(n4452), .A3(n4451), .A4(n4450), .ZN(n4455)
         );
  NAND2_X1 U5032 ( .A1(n4455), .A2(n4454), .ZN(U3244) );
  OAI211_X1 U5033 ( .C1(n4458), .C2(n4457), .A(n4573), .B(n4456), .ZN(n4463)
         );
  OAI211_X1 U5034 ( .C1(n4461), .C2(n4460), .A(n4571), .B(n4459), .ZN(n4462)
         );
  OAI211_X1 U5035 ( .C1(n4576), .C2(n4464), .A(n4463), .B(n4462), .ZN(n4465)
         );
  AOI211_X1 U5036 ( .C1(n4563), .C2(ADDR_REG_5__SCAN_IN), .A(n4466), .B(n4465), 
        .ZN(n4467) );
  INV_X1 U5037 ( .A(n4467), .ZN(U3245) );
  AOI21_X1 U5038 ( .B1(n4563), .B2(ADDR_REG_6__SCAN_IN), .A(n4468), .ZN(n4477)
         );
  OAI211_X1 U5039 ( .C1(REG1_REG_6__SCAN_IN), .C2(n4470), .A(n4573), .B(n4469), 
        .ZN(n4476) );
  OAI211_X1 U5040 ( .C1(REG2_REG_6__SCAN_IN), .C2(n4472), .A(n4571), .B(n4471), 
        .ZN(n4475) );
  NAND2_X1 U5041 ( .A1(n4473), .A2(n4536), .ZN(n4474) );
  NAND4_X1 U5042 ( .A1(n4477), .A2(n4476), .A3(n4475), .A4(n4474), .ZN(U3246)
         );
  AOI22_X1 U5043 ( .A1(REG1_REG_7__SCAN_IN), .A2(n4478), .B1(n4657), .B2(n2502), .ZN(n4481) );
  OAI21_X1 U5044 ( .B1(n4481), .B2(n4480), .A(n4573), .ZN(n4479) );
  AOI21_X1 U5045 ( .B1(n4481), .B2(n4480), .A(n4479), .ZN(n4483) );
  AOI211_X1 U5046 ( .C1(n4563), .C2(ADDR_REG_7__SCAN_IN), .A(n4483), .B(n4482), 
        .ZN(n4488) );
  OAI211_X1 U5047 ( .C1(n4486), .C2(n4485), .A(n4571), .B(n4484), .ZN(n4487)
         );
  OAI211_X1 U5048 ( .C1(n4576), .C2(n4657), .A(n4488), .B(n4487), .ZN(U3247)
         );
  AOI211_X1 U5049 ( .C1(n2524), .C2(n4490), .A(n4489), .B(n4540), .ZN(n4492)
         );
  AND2_X1 U5050 ( .A1(U3149), .A2(REG3_REG_8__SCAN_IN), .ZN(n4491) );
  AOI211_X1 U5051 ( .C1(n4563), .C2(ADDR_REG_8__SCAN_IN), .A(n4492), .B(n4491), 
        .ZN(n4496) );
  OAI211_X1 U5052 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4494), .A(n4571), .B(n4493), 
        .ZN(n4495) );
  OAI211_X1 U5053 ( .C1(n4576), .C2(n2179), .A(n4496), .B(n4495), .ZN(U3248)
         );
  AOI211_X1 U5054 ( .C1(n2562), .C2(n4498), .A(n4497), .B(n4540), .ZN(n4501)
         );
  INV_X1 U5055 ( .A(n4499), .ZN(n4500) );
  AOI211_X1 U5056 ( .C1(n4563), .C2(ADDR_REG_10__SCAN_IN), .A(n4501), .B(n4500), .ZN(n4505) );
  OAI211_X1 U5057 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4503), .A(n4571), .B(n4502), .ZN(n4504) );
  OAI211_X1 U5058 ( .C1(n4576), .C2(n4654), .A(n4505), .B(n4504), .ZN(U3250)
         );
  AOI211_X1 U5059 ( .C1(n2597), .C2(n4507), .A(n4506), .B(n4540), .ZN(n4510)
         );
  INV_X1 U5060 ( .A(n4508), .ZN(n4509) );
  AOI211_X1 U5061 ( .C1(n4563), .C2(ADDR_REG_12__SCAN_IN), .A(n4510), .B(n4509), .ZN(n4514) );
  OAI211_X1 U5062 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4512), .A(n4571), .B(n4511), .ZN(n4513) );
  OAI211_X1 U5063 ( .C1(n4576), .C2(n2105), .A(n4514), .B(n4513), .ZN(U3252)
         );
  AOI211_X1 U5064 ( .C1(n4517), .C2(n4516), .A(n4515), .B(n4540), .ZN(n4518)
         );
  AOI211_X1 U5065 ( .C1(n4563), .C2(ADDR_REG_13__SCAN_IN), .A(n4519), .B(n4518), .ZN(n4526) );
  AOI21_X1 U5066 ( .B1(n4521), .B2(n4651), .A(n4520), .ZN(n4524) );
  INV_X1 U5067 ( .A(n4571), .ZN(n4530) );
  AOI21_X1 U5068 ( .B1(n4524), .B2(n4523), .A(n4530), .ZN(n4522) );
  OAI21_X1 U5069 ( .B1(n4524), .B2(n4523), .A(n4522), .ZN(n4525) );
  OAI211_X1 U5070 ( .C1(n4576), .C2(n4651), .A(n4526), .B(n4525), .ZN(U3253)
         );
  NAND2_X1 U5071 ( .A1(ADDR_REG_14__SCAN_IN), .A2(n4563), .ZN(n4539) );
  AOI211_X1 U5072 ( .C1(n4529), .C2(n4528), .A(n4527), .B(n4540), .ZN(n4534)
         );
  AOI211_X1 U5073 ( .C1(n3559), .C2(n4532), .A(n4531), .B(n4530), .ZN(n4533)
         );
  AOI211_X1 U5074 ( .C1(n4536), .C2(n4535), .A(n4534), .B(n4533), .ZN(n4538)
         );
  NAND3_X1 U5075 ( .A1(n4539), .A2(n4538), .A3(n4537), .ZN(U3254) );
  AOI211_X1 U5076 ( .C1(n2054), .C2(n4542), .A(n4541), .B(n4540), .ZN(n4543)
         );
  AOI211_X1 U5077 ( .C1(n4563), .C2(ADDR_REG_15__SCAN_IN), .A(n4544), .B(n4543), .ZN(n4550) );
  AOI21_X1 U5078 ( .B1(n4547), .B2(n4546), .A(n4545), .ZN(n4548) );
  NAND2_X1 U5079 ( .A1(n4571), .A2(n4548), .ZN(n4549) );
  OAI211_X1 U5080 ( .C1(n4576), .C2(n4551), .A(n4550), .B(n4549), .ZN(U3255)
         );
  AOI21_X1 U5081 ( .B1(ADDR_REG_16__SCAN_IN), .B2(n4563), .A(n4552), .ZN(n4561) );
  OAI21_X1 U5082 ( .B1(n4555), .B2(n4554), .A(n4553), .ZN(n4559) );
  OAI21_X1 U5083 ( .B1(n4557), .B2(n3578), .A(n4556), .ZN(n4558) );
  AOI22_X1 U5084 ( .A1(n4573), .A2(n4559), .B1(n4571), .B2(n4558), .ZN(n4560)
         );
  OAI211_X1 U5085 ( .C1(n4645), .C2(n4576), .A(n4561), .B(n4560), .ZN(U3256)
         );
  AOI21_X1 U5086 ( .B1(ADDR_REG_17__SCAN_IN), .B2(n4563), .A(n4562), .ZN(n4575) );
  OAI21_X1 U5087 ( .B1(n4566), .B2(n4565), .A(n4564), .ZN(n4572) );
  OAI21_X1 U5088 ( .B1(n4569), .B2(n4568), .A(n4567), .ZN(n4570) );
  AOI22_X1 U5089 ( .A1(n4573), .A2(n4572), .B1(n4571), .B2(n4570), .ZN(n4574)
         );
  OAI211_X1 U5090 ( .C1(n4643), .C2(n4576), .A(n4575), .B(n4574), .ZN(U3257)
         );
  XNOR2_X1 U5091 ( .A(n4577), .B(n4578), .ZN(n4717) );
  XNOR2_X1 U5092 ( .A(n4579), .B(n4578), .ZN(n4586) );
  AOI22_X1 U5093 ( .A1(n4580), .A2(n4603), .B1(n4590), .B2(n4602), .ZN(n4584)
         );
  NAND2_X1 U5094 ( .A1(n4582), .A2(n4581), .ZN(n4583) );
  OAI211_X1 U5095 ( .C1(n4586), .C2(n4585), .A(n4584), .B(n4583), .ZN(n4587)
         );
  AOI21_X1 U5096 ( .B1(n4625), .B2(n4717), .A(n4587), .ZN(n4719) );
  AOI22_X1 U5097 ( .A1(n4588), .A2(n4629), .B1(REG2_REG_11__SCAN_IN), .B2(
        n4634), .ZN(n4592) );
  AOI21_X1 U5098 ( .B1(n4590), .B2(n2118), .A(n4589), .ZN(n4714) );
  AOI22_X1 U5099 ( .A1(n4717), .A2(n4630), .B1(n4617), .B2(n4714), .ZN(n4591)
         );
  OAI211_X1 U5100 ( .C1(n4634), .C2(n4719), .A(n4592), .B(n4591), .ZN(U3279)
         );
  AOI22_X1 U5101 ( .A1(n4593), .A2(n4629), .B1(REG2_REG_6__SCAN_IN), .B2(n4634), .ZN(n4597) );
  AOI22_X1 U5102 ( .A1(n4595), .A2(n4630), .B1(n4617), .B2(n4594), .ZN(n4596)
         );
  OAI211_X1 U5103 ( .C1(n4634), .C2(n4598), .A(n4597), .B(n4596), .ZN(U3284)
         );
  OAI21_X1 U5104 ( .B1(n4601), .B2(n4600), .A(n4599), .ZN(n4611) );
  AOI22_X1 U5105 ( .A1(n3050), .A2(n4603), .B1(n4602), .B2(n4613), .ZN(n4604)
         );
  OAI21_X1 U5106 ( .B1(n3053), .B2(n4627), .A(n4604), .ZN(n4610) );
  OAI21_X1 U5107 ( .B1(n4607), .B2(n4606), .A(n4605), .ZN(n4669) );
  NOR2_X1 U5108 ( .A1(n4669), .A2(n4608), .ZN(n4609) );
  AOI211_X1 U5109 ( .C1(n4624), .C2(n4611), .A(n4610), .B(n4609), .ZN(n4667)
         );
  AOI22_X1 U5110 ( .A1(REG2_REG_1__SCAN_IN), .A2(n4634), .B1(
        REG3_REG_1__SCAN_IN), .B2(n4629), .ZN(n4620) );
  INV_X1 U5111 ( .A(n4669), .ZN(n4618) );
  NAND2_X1 U5112 ( .A1(n4613), .A2(n4612), .ZN(n4615) );
  NAND2_X1 U5113 ( .A1(n4615), .A2(n4614), .ZN(n4668) );
  INV_X1 U5114 ( .A(n4668), .ZN(n4616) );
  AOI22_X1 U5115 ( .A1(n4618), .A2(n4630), .B1(n4617), .B2(n4616), .ZN(n4619)
         );
  OAI211_X1 U5116 ( .C1(n4634), .C2(n4667), .A(n4620), .B(n4619), .ZN(U3289)
         );
  NOR2_X1 U5117 ( .A1(n4622), .A2(n4621), .ZN(n4664) );
  INV_X1 U5118 ( .A(n4623), .ZN(n4628) );
  OAI21_X1 U5119 ( .B1(n4625), .B2(n4624), .A(n4665), .ZN(n4626) );
  OAI21_X1 U5120 ( .B1(n3048), .B2(n4627), .A(n4626), .ZN(n4663) );
  AOI21_X1 U5121 ( .B1(n4664), .B2(n4628), .A(n4663), .ZN(n4633) );
  AOI22_X1 U5122 ( .A1(n4665), .A2(n4630), .B1(REG3_REG_0__SCAN_IN), .B2(n4629), .ZN(n4631) );
  OAI221_X1 U5123 ( .B1(n4634), .B2(n4633), .C1(n3379), .C2(n4632), .A(n4631), 
        .ZN(U3290) );
  AND2_X1 U5124 ( .A1(D_REG_31__SCAN_IN), .A2(n4639), .ZN(U3291) );
  AND2_X1 U5125 ( .A1(D_REG_30__SCAN_IN), .A2(n4639), .ZN(U3292) );
  AND2_X1 U5126 ( .A1(D_REG_29__SCAN_IN), .A2(n4639), .ZN(U3293) );
  AND2_X1 U5127 ( .A1(D_REG_28__SCAN_IN), .A2(n4639), .ZN(U3294) );
  AND2_X1 U5128 ( .A1(D_REG_27__SCAN_IN), .A2(n4639), .ZN(U3295) );
  AND2_X1 U5129 ( .A1(D_REG_26__SCAN_IN), .A2(n4639), .ZN(U3296) );
  AND2_X1 U5130 ( .A1(D_REG_25__SCAN_IN), .A2(n4639), .ZN(U3297) );
  NOR2_X1 U5131 ( .A1(n4638), .A2(n4635), .ZN(U3298) );
  AND2_X1 U5132 ( .A1(D_REG_23__SCAN_IN), .A2(n4639), .ZN(U3299) );
  AND2_X1 U5133 ( .A1(D_REG_22__SCAN_IN), .A2(n4639), .ZN(U3300) );
  AND2_X1 U5134 ( .A1(n4639), .A2(D_REG_21__SCAN_IN), .ZN(U3301) );
  AND2_X1 U5135 ( .A1(D_REG_20__SCAN_IN), .A2(n4639), .ZN(U3302) );
  AND2_X1 U5136 ( .A1(D_REG_19__SCAN_IN), .A2(n4639), .ZN(U3303) );
  AND2_X1 U5137 ( .A1(D_REG_18__SCAN_IN), .A2(n4639), .ZN(U3304) );
  AND2_X1 U5138 ( .A1(D_REG_17__SCAN_IN), .A2(n4639), .ZN(U3305) );
  AND2_X1 U5139 ( .A1(D_REG_16__SCAN_IN), .A2(n4639), .ZN(U3306) );
  AND2_X1 U5140 ( .A1(D_REG_15__SCAN_IN), .A2(n4639), .ZN(U3307) );
  AND2_X1 U5141 ( .A1(D_REG_14__SCAN_IN), .A2(n4639), .ZN(U3308) );
  AND2_X1 U5142 ( .A1(D_REG_13__SCAN_IN), .A2(n4639), .ZN(U3309) );
  NOR2_X1 U5143 ( .A1(n4638), .A2(n4636), .ZN(U3310) );
  AND2_X1 U5144 ( .A1(D_REG_11__SCAN_IN), .A2(n4639), .ZN(U3311) );
  NOR2_X1 U5145 ( .A1(n4638), .A2(n4637), .ZN(U3312) );
  AND2_X1 U5146 ( .A1(D_REG_9__SCAN_IN), .A2(n4639), .ZN(U3313) );
  AND2_X1 U5147 ( .A1(D_REG_8__SCAN_IN), .A2(n4639), .ZN(U3314) );
  AND2_X1 U5148 ( .A1(D_REG_7__SCAN_IN), .A2(n4639), .ZN(U3315) );
  AND2_X1 U5149 ( .A1(D_REG_6__SCAN_IN), .A2(n4639), .ZN(U3316) );
  AND2_X1 U5150 ( .A1(D_REG_5__SCAN_IN), .A2(n4639), .ZN(U3317) );
  AND2_X1 U5151 ( .A1(D_REG_4__SCAN_IN), .A2(n4639), .ZN(U3318) );
  AND2_X1 U5152 ( .A1(D_REG_3__SCAN_IN), .A2(n4639), .ZN(U3319) );
  AND2_X1 U5153 ( .A1(D_REG_2__SCAN_IN), .A2(n4639), .ZN(U3320) );
  INV_X1 U5154 ( .A(DATAI_23_), .ZN(n4641) );
  AOI21_X1 U5155 ( .B1(U3149), .B2(n4641), .A(n4640), .ZN(U3329) );
  AOI22_X1 U5156 ( .A1(STATE_REG_SCAN_IN), .A2(n4643), .B1(n4642), .B2(U3149), 
        .ZN(U3335) );
  AOI22_X1 U5157 ( .A1(STATE_REG_SCAN_IN), .A2(n4645), .B1(n4644), .B2(U3149), 
        .ZN(U3336) );
  OAI22_X1 U5158 ( .A1(U3149), .A2(n4646), .B1(DATAI_15_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4647) );
  INV_X1 U5159 ( .A(n4647), .ZN(U3337) );
  AOI22_X1 U5160 ( .A1(STATE_REG_SCAN_IN), .A2(n4649), .B1(n4648), .B2(U3149), 
        .ZN(U3338) );
  INV_X1 U5161 ( .A(DATAI_13_), .ZN(n4650) );
  AOI22_X1 U5162 ( .A1(STATE_REG_SCAN_IN), .A2(n4651), .B1(n4650), .B2(U3149), 
        .ZN(U3339) );
  INV_X1 U5163 ( .A(DATAI_12_), .ZN(n4652) );
  AOI22_X1 U5164 ( .A1(STATE_REG_SCAN_IN), .A2(n2105), .B1(n4652), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U5165 ( .A(DATAI_10_), .ZN(n4653) );
  AOI22_X1 U5166 ( .A1(STATE_REG_SCAN_IN), .A2(n4654), .B1(n4653), .B2(U3149), 
        .ZN(U3342) );
  AOI22_X1 U5167 ( .A1(STATE_REG_SCAN_IN), .A2(n2179), .B1(n4655), .B2(U3149), 
        .ZN(U3344) );
  AOI22_X1 U5168 ( .A1(STATE_REG_SCAN_IN), .A2(n4657), .B1(n4656), .B2(U3149), 
        .ZN(U3345) );
  AOI22_X1 U5169 ( .A1(STATE_REG_SCAN_IN), .A2(n4659), .B1(n4658), .B2(U3149), 
        .ZN(U3346) );
  OAI22_X1 U5170 ( .A1(U3149), .A2(n4660), .B1(DATAI_5_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4661) );
  INV_X1 U5171 ( .A(n4661), .ZN(U3347) );
  AOI22_X1 U5172 ( .A1(STATE_REG_SCAN_IN), .A2(n2377), .B1(n4662), .B2(U3149), 
        .ZN(U3352) );
  AOI211_X1 U5173 ( .C1(n4716), .C2(n4665), .A(n4664), .B(n4663), .ZN(n4724)
         );
  AOI22_X1 U5174 ( .A1(n4722), .A2(n4724), .B1(n4666), .B2(n4720), .ZN(U3467)
         );
  INV_X1 U5175 ( .A(n4667), .ZN(n4671) );
  OAI22_X1 U5176 ( .A1(n4669), .A2(n4679), .B1(n4701), .B2(n4668), .ZN(n4670)
         );
  NOR2_X1 U5177 ( .A1(n4671), .A2(n4670), .ZN(n4725) );
  INV_X1 U5178 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4672) );
  AOI22_X1 U5179 ( .A1(n4722), .A2(n4725), .B1(n4672), .B2(n4720), .ZN(U3469)
         );
  AND3_X1 U5180 ( .A1(n4674), .A2(n4715), .A3(n4673), .ZN(n4676) );
  AOI211_X1 U5181 ( .C1(n4716), .C2(n4677), .A(n4676), .B(n4675), .ZN(n4726)
         );
  INV_X1 U5182 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4678) );
  AOI22_X1 U5183 ( .A1(n4722), .A2(n4726), .B1(n4678), .B2(n4720), .ZN(U3471)
         );
  NOR2_X1 U5184 ( .A1(n4680), .A2(n4679), .ZN(n4682) );
  AOI211_X1 U5185 ( .C1(n4715), .C2(n4683), .A(n4682), .B(n4681), .ZN(n4727)
         );
  INV_X1 U5186 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4684) );
  AOI22_X1 U5187 ( .A1(n4722), .A2(n4727), .B1(n4684), .B2(n4720), .ZN(U3473)
         );
  INV_X1 U5188 ( .A(n4685), .ZN(n4687) );
  AOI211_X1 U5189 ( .C1(n4688), .C2(n4716), .A(n4687), .B(n4686), .ZN(n4728)
         );
  INV_X1 U5190 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4689) );
  AOI22_X1 U5191 ( .A1(n4722), .A2(n4728), .B1(n4689), .B2(n4720), .ZN(U3475)
         );
  OAI21_X1 U5192 ( .B1(n4701), .B2(n4691), .A(n4690), .ZN(n4692) );
  AOI21_X1 U5193 ( .B1(n4693), .B2(n4704), .A(n4692), .ZN(n4729) );
  INV_X1 U5194 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4694) );
  AOI22_X1 U5195 ( .A1(n4722), .A2(n4729), .B1(n4694), .B2(n4720), .ZN(U3477)
         );
  AOI211_X1 U5196 ( .C1(n4697), .C2(n4704), .A(n4696), .B(n4695), .ZN(n4730)
         );
  INV_X1 U5197 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4698) );
  AOI22_X1 U5198 ( .A1(n4722), .A2(n4730), .B1(n4698), .B2(n4720), .ZN(U3481)
         );
  OAI21_X1 U5199 ( .B1(n4701), .B2(n4700), .A(n4699), .ZN(n4702) );
  AOI21_X1 U5200 ( .B1(n4704), .B2(n4703), .A(n4702), .ZN(n4731) );
  INV_X1 U5201 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4705) );
  AOI22_X1 U5202 ( .A1(n4722), .A2(n4731), .B1(n4705), .B2(n4720), .ZN(U3485)
         );
  NAND2_X1 U5203 ( .A1(n4706), .A2(n4715), .ZN(n4707) );
  NOR2_X1 U5204 ( .A1(n4708), .A2(n4707), .ZN(n4709) );
  AOI21_X1 U5205 ( .B1(n4710), .B2(n4716), .A(n4709), .ZN(n4711) );
  INV_X1 U5206 ( .A(REG0_REG_10__SCAN_IN), .ZN(n4713) );
  AOI22_X1 U5207 ( .A1(n4722), .A2(n4732), .B1(n4713), .B2(n4720), .ZN(U3487)
         );
  AOI22_X1 U5208 ( .A1(n4717), .A2(n4716), .B1(n4715), .B2(n4714), .ZN(n4718)
         );
  AND2_X1 U5209 ( .A1(n4719), .A2(n4718), .ZN(n4734) );
  INV_X1 U5210 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4721) );
  AOI22_X1 U5211 ( .A1(n4722), .A2(n4734), .B1(n4721), .B2(n4720), .ZN(U3489)
         );
  AOI22_X1 U5212 ( .A1(n4735), .A2(n4724), .B1(n4723), .B2(n4733), .ZN(U3518)
         );
  AOI22_X1 U5213 ( .A1(n4735), .A2(n4725), .B1(n3246), .B2(n4733), .ZN(U3519)
         );
  AOI22_X1 U5214 ( .A1(n4735), .A2(n4726), .B1(n3245), .B2(n4733), .ZN(U3520)
         );
  AOI22_X1 U5215 ( .A1(n4735), .A2(n4727), .B1(n2427), .B2(n4733), .ZN(U3521)
         );
  AOI22_X1 U5216 ( .A1(n4735), .A2(n4728), .B1(n3255), .B2(n4733), .ZN(U3522)
         );
  AOI22_X1 U5217 ( .A1(n4735), .A2(n4729), .B1(n2461), .B2(n4733), .ZN(U3523)
         );
  AOI22_X1 U5218 ( .A1(n4735), .A2(n4730), .B1(n2502), .B2(n4733), .ZN(U3525)
         );
  AOI22_X1 U5219 ( .A1(n4735), .A2(n4731), .B1(n2542), .B2(n4733), .ZN(U3527)
         );
  AOI22_X1 U5220 ( .A1(n4735), .A2(n4732), .B1(n2562), .B2(n4733), .ZN(U3528)
         );
  AOI22_X1 U5221 ( .A1(n4735), .A2(n4734), .B1(n3399), .B2(n4733), .ZN(U3529)
         );
  INV_X4 U2284 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
endmodule

