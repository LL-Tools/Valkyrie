

module b22_C_SARLock_k_64_5 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, 
        SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, 
        SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, 
        SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, 
        SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, P1_U3462, 
        P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, 
        P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, 
        P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, P2_U3292, 
        P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, 
        P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, 
        P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, 
        P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, P2_U3433, 
        P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, 
        P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, 
        P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, 
        P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, 
        P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, 
        P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3328, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, P3_U3293, 
        P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, P3_U3286, 
        P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, P3_U3279, 
        P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, P3_U3272, 
        P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, P3_U3265, 
        P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, P3_U3260, 
        P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, P3_U3253, 
        P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, P3_U3246, 
        P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, P3_U3239, 
        P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, P3_U3393, 
        P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, P3_U3414, 
        P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, P3_U3435, 
        P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, P3_U3449, 
        P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, 
        P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, 
        P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, 
        P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, 
        P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, 
        P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3233, 
        P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, P3_U3226, 
        P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, P3_U3219, 
        P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, P3_U3212, 
        P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, P3_U3205, 
        P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, P3_U3198, 
        P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, P3_U3191, 
        P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, P3_U3184, 
        P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, 
        P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, 
        P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, 
        P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, 
        P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3296, 
        P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, P3_U3175, 
        P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, P3_U3168, 
        P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, P3_U3161, 
        P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, P3_U3154, 
        P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6443, n6445, n6446, n6447, n6448, n6449, n6451, n6453, n6454, n6455,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15184, n15186;

  NAND2_X1 U7192 ( .A1(n13331), .A2(n13159), .ZN(n13332) );
  NOR2_X1 U7193 ( .A1(n10856), .A2(n14793), .ZN(n14813) );
  XNOR2_X1 U7194 ( .A(n6904), .B(n14802), .ZN(n14794) );
  INV_X2 U7195 ( .A(n8948), .ZN(n9528) );
  INV_X2 U7196 ( .A(n12247), .ZN(n12264) );
  INV_X2 U7197 ( .A(n12263), .ZN(n12255) );
  NAND2_X2 U7198 ( .A1(n9418), .A2(n9416), .ZN(n12263) );
  AND4_X1 U7199 ( .A1(n7487), .A2(n7486), .A3(n7485), .A4(n7484), .ZN(n10485)
         );
  INV_X1 U7200 ( .A(n12533), .ZN(n12543) );
  INV_X2 U7201 ( .A(n10789), .ZN(n12379) );
  CLKBUF_X2 U7202 ( .A(n8751), .Z(n6459) );
  NAND4_X1 U7203 ( .A1(n9632), .A2(n9631), .A3(n9630), .A4(n9629), .ZN(n13060)
         );
  CLKBUF_X2 U7204 ( .A(n8116), .Z(n8612) );
  INV_X1 U7205 ( .A(n14512), .ZN(n14486) );
  BUF_X4 U7206 ( .A(n8997), .Z(n6461) );
  BUF_X1 U7207 ( .A(n8120), .Z(n6457) );
  AND2_X2 U7208 ( .A1(n8039), .A2(n8730), .ZN(n13878) );
  INV_X2 U7209 ( .A(n7386), .ZN(n9335) );
  NOR2_X1 U7210 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n8964) );
  INV_X1 U7211 ( .A(n15184), .ZN(n6443) );
  INV_X2 U7212 ( .A(n6443), .ZN(P1_U3086) );
  INV_X1 U7213 ( .A(P1_STATE_REG_SCAN_IN), .ZN(n15184) );
  INV_X1 U7214 ( .A(n9279), .ZN(n6635) );
  NAND2_X1 U7215 ( .A1(n10535), .A2(n10140), .ZN(n8948) );
  NAND2_X1 U7216 ( .A1(n10065), .A2(n6461), .ZN(n9394) );
  INV_X1 U7217 ( .A(n10065), .ZN(n11898) );
  OR2_X1 U7218 ( .A1(n13402), .A2(n13404), .ZN(n7335) );
  INV_X2 U7219 ( .A(n8056), .ZN(n6454) );
  NAND2_X1 U7220 ( .A1(n6460), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7409) );
  INV_X2 U7221 ( .A(n13300), .ZN(n9633) );
  INV_X1 U7222 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9884) );
  AND3_X1 U7223 ( .A1(n8965), .A2(n8964), .A3(n9026), .ZN(n9064) );
  BUF_X1 U7224 ( .A(n8613), .Z(n8647) );
  NAND2_X1 U7225 ( .A1(n9824), .A2(n9266), .ZN(n13961) );
  NAND2_X1 U7226 ( .A1(n8001), .A2(n8037), .ZN(n8730) );
  INV_X2 U7227 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n15117) );
  NOR2_X1 U7228 ( .A1(n14794), .A2(n14795), .ZN(n14793) );
  INV_X1 U7229 ( .A(n7739), .ZN(n8761) );
  NAND2_X1 U7230 ( .A1(n11754), .A2(n11753), .ZN(n13410) );
  AND4_X1 U7231 ( .A1(n9354), .A2(n9353), .A3(n9352), .A4(n9351), .ZN(n11799)
         );
  NAND2_X1 U7232 ( .A1(n13515), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7148) );
  NAND2_X1 U7233 ( .A1(n8573), .A2(n8572), .ZN(n14028) );
  AND4_X1 U7234 ( .A1(n8087), .A2(n8088), .A3(n8086), .A4(n8089), .ZN(n8691)
         );
  INV_X1 U7235 ( .A(n10804), .ZN(n12378) );
  NAND4_X2 U7236 ( .A1(n8022), .A2(n8021), .A3(n8020), .A4(n8019), .ZN(n9279)
         );
  INV_X1 U7237 ( .A(n8007), .ZN(n8006) );
  OR2_X1 U7238 ( .A1(n14240), .A2(n14239), .ZN(n6445) );
  INV_X1 U7239 ( .A(n7386), .ZN(n8997) );
  NOR2_X1 U7240 ( .A1(n14866), .A2(n14867), .ZN(n14865) );
  BUF_X8 U7241 ( .A(n7897), .Z(n6446) );
  NAND2_X2 U7242 ( .A1(n7381), .A2(n7380), .ZN(n7897) );
  NAND2_X2 U7243 ( .A1(n7911), .A2(n9891), .ZN(n9893) );
  OAI21_X2 U7244 ( .B1(n12093), .B2(n13659), .A(n13824), .ZN(n13806) );
  INV_X1 U7245 ( .A(n8704), .ZN(n6447) );
  INV_X1 U7246 ( .A(n8704), .ZN(n6448) );
  INV_X1 U7247 ( .A(n8704), .ZN(n6449) );
  INV_X1 U7249 ( .A(n8704), .ZN(n6451) );
  INV_X4 U7251 ( .A(n6466), .ZN(n6453) );
  AND2_X2 U7252 ( .A1(n8053), .A2(n8644), .ZN(n8056) );
  INV_X1 U7254 ( .A(n8681), .ZN(n6455) );
  CLKBUF_X3 U7255 ( .A(n8113), .Z(n8681) );
  XNOR2_X2 U7256 ( .A(n11072), .B(n10864), .ZN(n10865) );
  AND2_X2 U7257 ( .A1(n8005), .A2(n6969), .ZN(n8007) );
  XNOR2_X2 U7258 ( .A(n12914), .B(n12912), .ZN(n13003) );
  NAND2_X2 U7259 ( .A1(n12305), .A2(n12306), .ZN(n11675) );
  NAND2_X2 U7260 ( .A1(n11672), .A2(n11671), .ZN(n12305) );
  AOI21_X2 U7261 ( .B1(n13003), .B2(n13002), .A(n12915), .ZN(n12916) );
  XOR2_X2 U7262 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), .Z(
        n14166) );
  XNOR2_X2 U7263 ( .A(n8519), .B(n8518), .ZN(n11961) );
  OAI221_X1 U7264 ( .B1(n15118), .B2(keyinput55), .C1(n15117), .C2(keyinput18), 
        .A(n15116), .ZN(n15123) );
  NAND2_X2 U7265 ( .A1(n10070), .A2(n10069), .ZN(n11848) );
  AND4_X2 U7266 ( .A1(n7373), .A2(n7372), .A3(n7371), .A4(n7370), .ZN(n14918)
         );
  NOR2_X2 U7267 ( .A1(n10926), .A2(n10925), .ZN(n11090) );
  AND4_X4 U7268 ( .A1(n7411), .A2(n7410), .A3(n7409), .A4(n7408), .ZN(n14920)
         );
  INV_X1 U7269 ( .A(n9624), .ZN(n9664) );
  AND2_X4 U7270 ( .A1(n9349), .A2(n11629), .ZN(n9624) );
  OAI22_X2 U7271 ( .A1(n11894), .A2(n7178), .B1(n11895), .B2(n7177), .ZN(
        n11904) );
  AND2_X2 U7272 ( .A1(n8084), .A2(n8083), .ZN(n14512) );
  OAI21_X2 U7273 ( .B1(n11675), .B2(n7013), .A(n7011), .ZN(n11697) );
  XNOR2_X2 U7274 ( .A(n8565), .B(SI_24_), .ZN(n8568) );
  NAND2_X2 U7275 ( .A1(n8544), .A2(n8543), .ZN(n8565) );
  NOR3_X2 U7276 ( .A1(n10953), .A2(n6831), .A3(n11621), .ZN(n11181) );
  NAND4_X2 U7277 ( .A1(n9672), .A2(n9671), .A3(n9670), .A4(n9669), .ZN(n13059)
         );
  AOI21_X2 U7278 ( .B1(n10514), .B2(n7916), .A(n7317), .ZN(n10422) );
  AND2_X2 U7279 ( .A1(n8797), .A2(n8796), .ZN(n8793) );
  AND2_X4 U7280 ( .A1(n10173), .A2(n12062), .ZN(n13300) );
  NAND2_X2 U7281 ( .A1(n9849), .A2(n9848), .ZN(n14702) );
  AND2_X4 U7282 ( .A1(n9349), .A2(n9350), .ZN(n7325) );
  NAND2_X2 U7283 ( .A1(n7377), .A2(n7376), .ZN(n12880) );
  MUX2_X2 U7284 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7375), .S(
        P3_IR_REG_28__SCAN_IN), .Z(n7377) );
  NOR2_X2 U7285 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n8282) );
  XNOR2_X2 U7286 ( .A(n9139), .B(n9138), .ZN(n9330) );
  NAND2_X2 U7287 ( .A1(n9137), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9139) );
  CLKBUF_X1 U7288 ( .A(n8751), .Z(n6458) );
  BUF_X4 U7289 ( .A(n8751), .Z(n6460) );
  AND2_X2 U7290 ( .A1(n7368), .A2(n7367), .ZN(n8751) );
  NAND2_X2 U7291 ( .A1(n12673), .A2(n7765), .ZN(n12657) );
  NAND2_X2 U7292 ( .A1(n7282), .A2(n6584), .ZN(n12673) );
  XNOR2_X2 U7293 ( .A(n7148), .B(n9344), .ZN(n9348) );
  NOR2_X2 U7294 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n7428) );
  OAI21_X2 U7295 ( .B1(n10288), .B2(n10287), .A(n10286), .ZN(n10455) );
  AND2_X2 U7296 ( .A1(n10277), .A2(n10278), .ZN(n10288) );
  XNOR2_X2 U7297 ( .A(n8002), .B(P1_IR_REG_30__SCAN_IN), .ZN(n12131) );
  NAND2_X1 U7298 ( .A1(n10290), .A2(n10289), .ZN(n14475) );
  NAND2_X2 U7299 ( .A1(n12611), .A2(n7828), .ZN(n12598) );
  AOI211_X2 U7300 ( .C1(n14517), .C2(n14035), .A(n14034), .B(n14033), .ZN(
        n14101) );
  AOI21_X4 U7301 ( .B1(n12657), .B2(n7780), .A(n7779), .ZN(n12645) );
  XNOR2_X2 U7302 ( .A(n11661), .B(n11659), .ZN(n12337) );
  NAND2_X2 U7303 ( .A1(n12296), .A2(n11658), .ZN(n11661) );
  NOR2_X2 U7304 ( .A1(n14209), .A2(n14420), .ZN(n14424) );
  NOR2_X2 U7305 ( .A1(n14206), .A2(n14205), .ZN(n14420) );
  OAI21_X2 U7306 ( .B1(n8568), .B2(n8567), .A(n8566), .ZN(n8586) );
  NAND2_X2 U7307 ( .A1(n7364), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7365) );
  XNOR2_X2 U7308 ( .A(n11665), .B(n11666), .ZN(n12282) );
  NAND2_X2 U7309 ( .A1(n11663), .A2(n11662), .ZN(n11665) );
  XNOR2_X2 U7310 ( .A(n7720), .B(P3_IR_REG_19__SCAN_IN), .ZN(n12533) );
  INV_X2 U7312 ( .A(n7760), .ZN(n7541) );
  NAND2_X1 U7313 ( .A1(n12110), .A2(n12091), .ZN(n13868) );
  CLKBUF_X1 U7314 ( .A(n12945), .Z(n6623) );
  NAND2_X1 U7315 ( .A1(n11744), .A2(n12055), .ZN(n11792) );
  NAND2_X1 U7316 ( .A1(n8609), .A2(n8608), .ZN(n14014) );
  XNOR2_X1 U7317 ( .A(n12182), .B(n12181), .ZN(n13645) );
  NAND2_X1 U7318 ( .A1(n11963), .A2(n11962), .ZN(n13438) );
  NAND2_X1 U7319 ( .A1(n12164), .A2(n6531), .ZN(n14345) );
  OAI21_X2 U7320 ( .B1(n8586), .B2(n6605), .A(n7213), .ZN(n8619) );
  AOI21_X1 U7321 ( .B1(n6888), .B2(n6468), .A(n6887), .ZN(n11198) );
  NAND2_X1 U7322 ( .A1(n6644), .A2(n11209), .ZN(n11277) );
  NAND2_X1 U7323 ( .A1(n10079), .A2(n7249), .ZN(n10120) );
  INV_X1 U7324 ( .A(n14467), .ZN(n6954) );
  INV_X1 U7325 ( .A(n14521), .ZN(n10615) );
  NAND2_X1 U7326 ( .A1(n8792), .A2(n8789), .ZN(n8763) );
  INV_X4 U7327 ( .A(n12174), .ZN(n12247) );
  CLKBUF_X2 U7328 ( .A(n9633), .Z(n14633) );
  INV_X2 U7329 ( .A(n11720), .ZN(n12013) );
  NAND4_X2 U7330 ( .A1(n9363), .A2(n9362), .A3(n9361), .A4(n9360), .ZN(n13064)
         );
  NAND2_X1 U7332 ( .A1(n7325), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n9362) );
  NAND2_X1 U7334 ( .A1(n7895), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7891) );
  INV_X4 U7335 ( .A(n11980), .ZN(n12001) );
  INV_X1 U7336 ( .A(n9840), .ZN(n10439) );
  NAND2_X1 U7337 ( .A1(n7892), .A2(n7889), .ZN(n7895) );
  AND2_X1 U7338 ( .A1(n7888), .A2(n7887), .ZN(n7892) );
  CLKBUF_X2 U7339 ( .A(n9332), .Z(n13154) );
  XNOR2_X1 U7340 ( .A(n6627), .B(n8016), .ZN(n8740) );
  AND2_X1 U7341 ( .A1(n7374), .A2(n7360), .ZN(n7363) );
  INV_X1 U7342 ( .A(n8111), .ZN(n7386) );
  NAND4_X1 U7343 ( .A1(n8090), .A2(n7306), .A3(n7307), .A4(n7989), .ZN(n8068)
         );
  AOI211_X1 U7344 ( .C1(n8720), .C2(n8719), .A(n8718), .B(n8717), .ZN(n8724)
         );
  OR2_X1 U7345 ( .A1(n13418), .A2(n13417), .ZN(n13499) );
  NAND2_X1 U7346 ( .A1(n13311), .A2(n13312), .ZN(n6775) );
  NOR2_X1 U7347 ( .A1(n13408), .A2(n7141), .ZN(n7140) );
  AOI21_X1 U7348 ( .B1(n14006), .B2(n14529), .A(n14005), .ZN(n14007) );
  NAND2_X1 U7349 ( .A1(n7092), .A2(n13186), .ZN(n13311) );
  NAND2_X1 U7350 ( .A1(n13325), .A2(n13185), .ZN(n7092) );
  OAI21_X1 U7351 ( .B1(n14251), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n6445), .ZN(
        n6639) );
  AND2_X1 U7352 ( .A1(n6899), .A2(n6488), .ZN(n13633) );
  NAND2_X1 U7353 ( .A1(n13806), .A2(n13820), .ZN(n13807) );
  OR2_X1 U7354 ( .A1(n13409), .A2(n7142), .ZN(n7141) );
  OR2_X1 U7355 ( .A1(n11667), .A2(n11666), .ZN(n11668) );
  AOI21_X1 U7356 ( .B1(n6868), .B2(n6870), .A(n6867), .ZN(n13826) );
  NAND2_X1 U7357 ( .A1(n13179), .A2(n13178), .ZN(n13363) );
  XNOR2_X1 U7358 ( .A(n7083), .B(n7082), .ZN(n14251) );
  OAI21_X1 U7359 ( .B1(n14280), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n6480), .ZN(
        n7083) );
  XNOR2_X1 U7360 ( .A(n8677), .B(n6609), .ZN(n11716) );
  NAND2_X1 U7361 ( .A1(n7208), .A2(n8638), .ZN(n8677) );
  NAND2_X1 U7362 ( .A1(n11462), .A2(n11461), .ZN(n11464) );
  AOI21_X1 U7363 ( .B1(n6870), .B2(n12091), .A(n6872), .ZN(n6869) );
  NAND2_X1 U7364 ( .A1(n8623), .A2(n8622), .ZN(n14009) );
  AND2_X1 U7365 ( .A1(n7079), .A2(n7078), .ZN(n14436) );
  NAND2_X1 U7366 ( .A1(n11765), .A2(n11764), .ZN(n13265) );
  NAND2_X1 U7367 ( .A1(n11776), .A2(n11775), .ZN(n13420) );
  INV_X1 U7368 ( .A(n12716), .ZN(n12717) );
  NAND2_X1 U7369 ( .A1(n14345), .A2(n12173), .ZN(n12182) );
  AOI21_X1 U7370 ( .B1(n14431), .B2(n6705), .A(n6704), .ZN(n14221) );
  XNOR2_X1 U7371 ( .A(n8619), .B(n8607), .ZN(n13522) );
  AND2_X1 U7372 ( .A1(n6707), .A2(n6706), .ZN(n14431) );
  NAND2_X1 U7373 ( .A1(n11982), .A2(n11981), .ZN(n13432) );
  NAND2_X1 U7374 ( .A1(n11623), .A2(n11622), .ZN(n12164) );
  INV_X1 U7375 ( .A(n13347), .ZN(n6463) );
  NAND2_X1 U7376 ( .A1(n11617), .A2(n11616), .ZN(n11623) );
  OR2_X1 U7377 ( .A1(n14426), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n6707) );
  NAND2_X1 U7378 ( .A1(n8486), .A2(n8485), .ZN(n14051) );
  NAND2_X1 U7379 ( .A1(n6679), .A2(n6678), .ZN(n14385) );
  AND2_X1 U7380 ( .A1(n8469), .A2(n8468), .ZN(n14114) );
  NOR2_X1 U7381 ( .A1(n14208), .A2(n14207), .ZN(n14419) );
  OAI21_X1 U7382 ( .B1(n10355), .B2(n10354), .A(n6645), .ZN(n10653) );
  AND2_X1 U7383 ( .A1(n6504), .A2(n12103), .ZN(n13950) );
  OR2_X1 U7384 ( .A1(n14300), .A2(n8836), .ZN(n7924) );
  OAI21_X1 U7385 ( .B1(n8484), .B2(n8497), .A(n6483), .ZN(n6621) );
  NAND2_X1 U7386 ( .A1(n8431), .A2(n8430), .ZN(n13967) );
  OAI21_X1 U7387 ( .B1(n8438), .B2(n8437), .A(n8440), .ZN(n8467) );
  AND2_X1 U7388 ( .A1(n8405), .A2(n8404), .ZN(n14124) );
  NAND2_X1 U7389 ( .A1(n8416), .A2(n8415), .ZN(n14372) );
  XNOR2_X1 U7390 ( .A(n10239), .B(n10240), .ZN(n10243) );
  XNOR2_X1 U7391 ( .A(n8439), .B(SI_18_), .ZN(n8438) );
  NAND2_X1 U7392 ( .A1(n13546), .A2(n6492), .ZN(n10239) );
  XNOR2_X1 U7393 ( .A(n14200), .B(n14199), .ZN(n14258) );
  INV_X1 U7394 ( .A(n7073), .ZN(n14200) );
  XNOR2_X1 U7395 ( .A(n6905), .B(n14875), .ZN(n14866) );
  NAND2_X2 U7396 ( .A1(n9857), .A2(n9856), .ZN(n14619) );
  NAND2_X1 U7397 ( .A1(n9899), .A2(n9898), .ZN(n9925) );
  NOR2_X2 U7398 ( .A1(n12148), .A2(n13878), .ZN(n14494) );
  AND2_X1 U7399 ( .A1(n8101), .A2(n10281), .ZN(n10291) );
  XNOR2_X1 U7400 ( .A(n7068), .B(P2_ADDR_REG_6__SCAN_IN), .ZN(n14256) );
  OAI21_X1 U7401 ( .B1(n15169), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6530), .ZN(
        n7068) );
  NAND2_X2 U7402 ( .A1(n12255), .A2(n13961), .ZN(n9810) );
  NAND2_X1 U7403 ( .A1(n6550), .A2(n7225), .ZN(n11806) );
  OAI211_X1 U7404 ( .C1(n9643), .C2(n9394), .A(n9642), .B(n9641), .ZN(n14634)
         );
  OR2_X1 U7405 ( .A1(n14775), .A2(n7316), .ZN(n6904) );
  AND3_X1 U7406 ( .A1(n7434), .A2(n7433), .A3(n7432), .ZN(n9890) );
  AND3_X1 U7407 ( .A1(n7400), .A2(n7399), .A3(n7398), .ZN(n10148) );
  AND4_X1 U7408 ( .A1(n8011), .A2(n8010), .A3(n8009), .A4(n8008), .ZN(n9695)
         );
  AND4_X1 U7409 ( .A1(n8065), .A2(n8064), .A3(n8063), .A4(n8062), .ZN(n9817)
         );
  XNOR2_X1 U7410 ( .A(n13878), .B(n9824), .ZN(n8052) );
  INV_X1 U7411 ( .A(n7200), .ZN(n7199) );
  AND2_X1 U7412 ( .A1(n7955), .A2(n7975), .ZN(n9089) );
  INV_X2 U7413 ( .A(n9530), .ZN(n7427) );
  NAND2_X1 U7414 ( .A1(n9273), .A2(n10586), .ZN(n9416) );
  AND2_X1 U7415 ( .A1(n8051), .A2(n8050), .ZN(n9273) );
  MUX2_X1 U7416 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8044), .S(
        P1_IR_REG_22__SCAN_IN), .Z(n8045) );
  CLKBUF_X1 U7417 ( .A(n9378), .Z(n12056) );
  AND2_X1 U7418 ( .A1(n7366), .A2(n12873), .ZN(n7367) );
  XOR2_X1 U7419 ( .A(n14165), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n15168) );
  NAND2_X1 U7420 ( .A1(n7366), .A2(n12873), .ZN(n12157) );
  NAND2_X1 U7421 ( .A1(n8733), .A2(n8734), .ZN(n11515) );
  NAND2_X1 U7422 ( .A1(n8739), .A2(n8738), .ZN(n11373) );
  MUX2_X1 U7423 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7361), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n7366) );
  OAI21_X1 U7424 ( .B1(n8726), .B2(P1_IR_REG_23__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8727) );
  INV_X2 U7425 ( .A(n9394), .ZN(n9951) );
  NAND2_X1 U7426 ( .A1(n8048), .A2(n8047), .ZN(n10586) );
  NAND2_X1 U7427 ( .A1(n7948), .A2(n7949), .ZN(n11225) );
  INV_X2 U7428 ( .A(n12875), .ZN(n12886) );
  MUX2_X1 U7429 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8004), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n8005) );
  INV_X1 U7430 ( .A(n9332), .ZN(n10176) );
  OR2_X1 U7431 ( .A1(n9133), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n9136) );
  NAND3_X1 U7432 ( .A1(n6505), .A2(n7135), .A3(n7136), .ZN(n9332) );
  NAND2_X2 U7433 ( .A1(n9335), .A2(P2_U3088), .ZN(n13526) );
  NAND2_X1 U7434 ( .A1(n6969), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8002) );
  OR2_X1 U7435 ( .A1(n8015), .A2(n14125), .ZN(n6627) );
  AND2_X1 U7436 ( .A1(n7947), .A2(n7287), .ZN(n7374) );
  XNOR2_X1 U7437 ( .A(n14142), .B(n14141), .ZN(n14178) );
  NAND2_X1 U7438 ( .A1(n8078), .A2(SI_3_), .ZN(n8109) );
  OR2_X1 U7439 ( .A1(n9197), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n9200) );
  OR2_X1 U7440 ( .A1(n9547), .A2(n7407), .ZN(n9773) );
  AND3_X1 U7441 ( .A1(n8001), .A2(n8017), .A3(n7341), .ZN(n8015) );
  XNOR2_X1 U7442 ( .A(n7431), .B(n7430), .ZN(n10851) );
  AND2_X1 U7443 ( .A1(n7332), .A2(n7358), .ZN(n6630) );
  NOR2_X1 U7444 ( .A1(n7357), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n7275) );
  INV_X1 U7445 ( .A(n7472), .ZN(n7349) );
  AOI21_X1 U7446 ( .B1(n7072), .B2(n14168), .A(n7071), .ZN(n14173) );
  AND3_X1 U7447 ( .A1(n6714), .A2(n6713), .A3(n6712), .ZN(n9325) );
  AND4_X1 U7448 ( .A1(n7352), .A2(n7645), .A3(n7351), .A4(n7350), .ZN(n7332)
         );
  AND3_X1 U7449 ( .A1(n7997), .A2(n7996), .A3(n7995), .ZN(n8728) );
  AND4_X1 U7450 ( .A1(n7347), .A2(n7346), .A3(n7345), .A4(n7344), .ZN(n7348)
         );
  INV_X1 U7451 ( .A(n8068), .ZN(n6464) );
  INV_X1 U7452 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n14245) );
  INV_X1 U7453 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7383) );
  NOR3_X1 U7454 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .A3(
        P2_IR_REG_4__SCAN_IN), .ZN(n8967) );
  NOR2_X1 U7455 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n8965) );
  NOR2_X1 U7456 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n7999) );
  NOR2_X1 U7457 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n7998) );
  INV_X1 U7458 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n8208) );
  INV_X1 U7459 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n8309) );
  NOR3_X1 U7460 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .A3(
        P2_IR_REG_12__SCAN_IN), .ZN(n8968) );
  NOR2_X1 U7461 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n6714) );
  NOR2_X1 U7462 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n6713) );
  INV_X1 U7463 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9344) );
  NOR2_X1 U7464 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n6712) );
  NOR2_X1 U7465 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n7990) );
  NOR2_X1 U7466 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n7344) );
  NOR2_X1 U7467 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n7345) );
  NOR2_X1 U7468 ( .A1(P3_IR_REG_13__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), .ZN(
        n7352) );
  INV_X4 U7469 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X4 U7470 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NOR2_X1 U7471 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n7346) );
  NOR2_X1 U7472 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n6984) );
  AND2_X1 U7473 ( .A1(n12131), .A2(n8006), .ZN(n8116) );
  NOR2_X1 U7474 ( .A1(n12131), .A2(n8007), .ZN(n8120) );
  OR2_X4 U7475 ( .A1(n11719), .A2(n12072), .ZN(n11720) );
  OAI21_X2 U7476 ( .B1(n12106), .B2(n6978), .A(n6976), .ZN(n13886) );
  NOR2_X2 U7477 ( .A1(n14898), .A2(n10863), .ZN(n11072) );
  CLKBUF_X1 U7478 ( .A(n9559), .Z(n6465) );
  XNOR2_X1 U7479 ( .A(n7403), .B(n7402), .ZN(n9559) );
  AND2_X1 U7480 ( .A1(n8053), .A2(n8644), .ZN(n6466) );
  NOR2_X2 U7481 ( .A1(n11806), .A2(n11802), .ZN(n10324) );
  NOR2_X4 U7482 ( .A1(n13856), .A2(n14028), .ZN(n13838) );
  OR2_X1 U7483 ( .A1(n7985), .A2(n12568), .ZN(n8925) );
  NAND2_X1 U7484 ( .A1(n6513), .A2(n9988), .ZN(n7108) );
  AND3_X2 U7485 ( .A1(n6837), .A2(n15186), .A3(n6464), .ZN(n8001) );
  NOR2_X1 U7486 ( .A1(n6886), .A2(n6957), .ZN(n6837) );
  NAND2_X1 U7487 ( .A1(n7994), .A2(n6959), .ZN(n6957) );
  NAND2_X1 U7488 ( .A1(n13298), .A2(n13191), .ZN(n13286) );
  NAND2_X1 U7489 ( .A1(n11543), .A2(n11542), .ZN(n11545) );
  OR2_X1 U7490 ( .A1(n7096), .A2(n11366), .ZN(n7093) );
  AND2_X1 U7491 ( .A1(n6750), .A2(n12046), .ZN(n7096) );
  NAND2_X1 U7492 ( .A1(n7098), .A2(n11305), .ZN(n6750) );
  INV_X1 U7493 ( .A(n9084), .ZN(n8444) );
  NAND2_X1 U7494 ( .A1(n8271), .A2(n8273), .ZN(n7301) );
  NOR2_X1 U7495 ( .A1(n11173), .A2(n8334), .ZN(n8351) );
  NOR2_X1 U7496 ( .A1(n8406), .A2(n8407), .ZN(n7311) );
  AOI21_X1 U7497 ( .B1(n8406), .B2(n8407), .A(n6548), .ZN(n7312) );
  NAND2_X1 U7498 ( .A1(n11880), .A2(n11883), .ZN(n6746) );
  NAND2_X1 U7499 ( .A1(n6759), .A2(n6760), .ZN(n11954) );
  AND2_X1 U7500 ( .A1(n7205), .A2(n6510), .ZN(n7204) );
  NAND2_X1 U7501 ( .A1(n6732), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n7186) );
  INV_X1 U7502 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7382) );
  OR2_X1 U7503 ( .A1(n12766), .A2(n12659), .ZN(n8891) );
  NOR2_X1 U7504 ( .A1(n7704), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n6618) );
  OR2_X1 U7505 ( .A1(n7634), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n7652) );
  AND2_X1 U7506 ( .A1(n11251), .A2(n7625), .ZN(n7278) );
  NAND2_X1 U7507 ( .A1(n10231), .A2(n7912), .ZN(n7283) );
  NAND2_X1 U7508 ( .A1(n12947), .A2(n12946), .ZN(n12945) );
  NAND2_X1 U7509 ( .A1(n6498), .A2(n7128), .ZN(n7127) );
  AOI21_X1 U7510 ( .B1(n7131), .B2(n7128), .A(n7126), .ZN(n7125) );
  NOR2_X1 U7511 ( .A1(n13416), .A2(n13222), .ZN(n7126) );
  INV_X1 U7512 ( .A(n13206), .ZN(n6790) );
  NAND2_X1 U7513 ( .A1(n9417), .A2(n9418), .ZN(n12174) );
  OR2_X1 U7514 ( .A1(n14397), .A2(n14340), .ZN(n11452) );
  XNOR2_X1 U7515 ( .A(n6954), .B(n13674), .ZN(n6955) );
  NAND2_X1 U7516 ( .A1(n10621), .A2(n10293), .ZN(n6956) );
  NAND2_X1 U7517 ( .A1(n8638), .A2(n6609), .ZN(n7211) );
  INV_X1 U7518 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8040) );
  INV_X1 U7519 ( .A(n8730), .ZN(n8041) );
  XNOR2_X1 U7520 ( .A(n8483), .B(SI_20_), .ZN(n8482) );
  INV_X1 U7521 ( .A(n8408), .ZN(n7207) );
  XNOR2_X1 U7522 ( .A(n8396), .B(SI_14_), .ZN(n8358) );
  NAND2_X1 U7523 ( .A1(n7199), .A2(n6727), .ZN(n6726) );
  INV_X1 U7524 ( .A(n8296), .ZN(n6727) );
  OAI21_X1 U7525 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n14156), .A(n14155), .ZN(
        n14213) );
  AOI21_X1 U7526 ( .B1(n7001), .B2(n11276), .A(n6475), .ZN(n6999) );
  INV_X1 U7527 ( .A(n12585), .ZN(n12555) );
  OAI21_X1 U7528 ( .B1(n12572), .B2(n8909), .A(n8910), .ZN(n8931) );
  NAND2_X1 U7529 ( .A1(n6470), .A2(n7274), .ZN(n7272) );
  INV_X1 U7530 ( .A(n12680), .ZN(n7764) );
  OR2_X1 U7531 ( .A1(n7742), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n7755) );
  OR2_X1 U7532 ( .A1(n12566), .A2(n7873), .ZN(n7886) );
  NAND2_X1 U7533 ( .A1(n7057), .A2(n7769), .ZN(n7056) );
  INV_X1 U7534 ( .A(n7782), .ZN(n7057) );
  AND2_X1 U7535 ( .A1(n13189), .A2(n13188), .ZN(n6774) );
  OR2_X1 U7536 ( .A1(n13447), .A2(n13209), .ZN(n6791) );
  OAI21_X1 U7537 ( .B1(n13389), .B2(n6536), .A(n13204), .ZN(n13368) );
  NAND2_X1 U7538 ( .A1(n13174), .A2(n13173), .ZN(n13383) );
  OAI21_X1 U7539 ( .B1(n6793), .B2(n6795), .A(n6792), .ZN(n11433) );
  AOI21_X1 U7540 ( .B1(n6794), .B2(n6796), .A(n6523), .ZN(n6792) );
  NAND2_X1 U7541 ( .A1(n11426), .A2(n11425), .ZN(n11543) );
  NAND2_X1 U7542 ( .A1(n7100), .A2(n11305), .ZN(n7094) );
  OR2_X1 U7543 ( .A1(n11306), .A2(n7099), .ZN(n7098) );
  INV_X1 U7544 ( .A(n11150), .ZN(n7099) );
  XNOR2_X1 U7545 ( .A(n13481), .B(n11343), .ZN(n12046) );
  OAI21_X1 U7546 ( .B1(n10544), .B2(n7147), .A(n7145), .ZN(n10817) );
  AOI21_X1 U7547 ( .B1(n7146), .B2(n10759), .A(n6537), .ZN(n7145) );
  NOR2_X1 U7548 ( .A1(n6806), .A2(n12034), .ZN(n6805) );
  INV_X1 U7549 ( .A(n6808), .ZN(n6806) );
  NAND2_X1 U7550 ( .A1(n7104), .A2(n7103), .ZN(n7102) );
  INV_X1 U7551 ( .A(n7108), .ZN(n7103) );
  NAND2_X1 U7552 ( .A1(n6461), .A2(n7229), .ZN(n7228) );
  INV_X1 U7553 ( .A(n9374), .ZN(n7229) );
  NAND2_X1 U7554 ( .A1(n13248), .A2(n13247), .ZN(n13246) );
  NOR2_X1 U7555 ( .A1(n7331), .A2(n6560), .ZN(n6672) );
  INV_X1 U7556 ( .A(n11022), .ZN(n6891) );
  AND2_X1 U7557 ( .A1(n11173), .A2(n11172), .ZN(n6982) );
  NAND2_X1 U7558 ( .A1(n9084), .A2(n9376), .ZN(n8094) );
  NAND2_X1 U7559 ( .A1(n9084), .A2(n9335), .ZN(n8113) );
  NAND2_X1 U7560 ( .A1(n9418), .A2(n8993), .ZN(n10305) );
  OAI21_X1 U7561 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n14225), .A(n14224), .ZN(
        n14229) );
  NAND2_X1 U7562 ( .A1(n7014), .A2(n6533), .ZN(n12317) );
  NAND2_X1 U7563 ( .A1(n13621), .A2(n6664), .ZN(n10606) );
  NAND2_X1 U7564 ( .A1(n10601), .A2(n6665), .ZN(n6664) );
  NAND2_X1 U7565 ( .A1(n8446), .A2(n8445), .ZN(n14063) );
  NAND2_X1 U7566 ( .A1(n8057), .A2(n6449), .ZN(n8058) );
  NAND2_X1 U7567 ( .A1(n8054), .A2(n6454), .ZN(n8059) );
  OAI22_X1 U7568 ( .A1(n11827), .A2(n7168), .B1(n11828), .B2(n7167), .ZN(n6766) );
  NOR2_X1 U7569 ( .A1(n11829), .A2(n11826), .ZN(n7168) );
  INV_X1 U7570 ( .A(n11826), .ZN(n7167) );
  NAND2_X1 U7571 ( .A1(n6628), .A2(n6538), .ZN(n8811) );
  OAI211_X1 U7572 ( .C1(n8804), .C2(n8805), .A(n10230), .B(n8803), .ZN(n6628)
         );
  NAND2_X1 U7573 ( .A1(n11849), .A2(n11852), .ZN(n6739) );
  NOR2_X1 U7574 ( .A1(n11856), .A2(n11853), .ZN(n7163) );
  NAND2_X1 U7575 ( .A1(n11856), .A2(n11853), .ZN(n7162) );
  INV_X1 U7576 ( .A(n11844), .ZN(n7179) );
  NOR2_X1 U7577 ( .A1(n11844), .A2(n11847), .ZN(n7180) );
  NOR2_X1 U7578 ( .A1(n7163), .A2(n6737), .ZN(n6736) );
  INV_X1 U7579 ( .A(n6739), .ZN(n6737) );
  INV_X1 U7580 ( .A(n7162), .ZN(n6734) );
  INV_X1 U7581 ( .A(n11849), .ZN(n6740) );
  NOR2_X1 U7582 ( .A1(n7311), .A2(n6539), .ZN(n7309) );
  INV_X1 U7583 ( .A(n7311), .ZN(n7308) );
  INV_X1 U7584 ( .A(n12103), .ZN(n7305) );
  INV_X1 U7585 ( .A(n11863), .ZN(n7173) );
  NOR2_X1 U7586 ( .A1(n11866), .A2(n11863), .ZN(n7174) );
  NOR2_X1 U7587 ( .A1(n11887), .A2(n11884), .ZN(n7158) );
  NAND2_X1 U7588 ( .A1(n6745), .A2(n6746), .ZN(n11885) );
  AOI21_X1 U7589 ( .B1(n6509), .B2(n6747), .A(n6742), .ZN(n6741) );
  AOI21_X1 U7590 ( .B1(n7153), .B2(n7152), .A(n7151), .ZN(n7150) );
  AOI21_X1 U7591 ( .B1(n6757), .B2(n6761), .A(n6755), .ZN(n6754) );
  NAND2_X1 U7592 ( .A1(n6625), .A2(n10742), .ZN(n7564) );
  NOR2_X1 U7593 ( .A1(n14014), .A2(n13640), .ZN(n6829) );
  NOR2_X1 U7594 ( .A1(n13934), .A2(n6865), .ZN(n6860) );
  AOI21_X1 U7595 ( .B1(n6726), .B2(n8295), .A(n6724), .ZN(n6723) );
  INV_X1 U7596 ( .A(n8342), .ZN(n6724) );
  INV_X1 U7597 ( .A(n6699), .ZN(n14144) );
  OAI21_X1 U7598 ( .B1(n14178), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n6564), .ZN(
        n6699) );
  INV_X1 U7599 ( .A(n14766), .ZN(n10882) );
  NAND2_X1 U7600 ( .A1(n14786), .A2(n6525), .ZN(n10870) );
  NAND2_X1 U7601 ( .A1(n14822), .A2(n6655), .ZN(n10872) );
  OR2_X1 U7602 ( .A1(n10897), .A2(n14999), .ZN(n6655) );
  NAND2_X1 U7603 ( .A1(n14858), .A2(n6656), .ZN(n10874) );
  OR2_X1 U7604 ( .A1(n10908), .A2(n15002), .ZN(n6656) );
  NAND2_X1 U7605 ( .A1(n14886), .A2(n10876), .ZN(n11077) );
  NAND2_X1 U7606 ( .A1(n12389), .A2(n6603), .ZN(n12410) );
  AOI21_X1 U7607 ( .B1(n12460), .B2(n12459), .A(n12501), .ZN(n6927) );
  OR2_X1 U7608 ( .A1(n12752), .A2(n12309), .ZN(n8902) );
  NAND2_X1 U7609 ( .A1(n12640), .A2(n6487), .ZN(n12623) );
  NAND2_X1 U7610 ( .A1(n7933), .A2(n6945), .ZN(n6944) );
  INV_X1 U7611 ( .A(n6946), .ZN(n6945) );
  NOR2_X1 U7612 ( .A1(n8877), .A2(n8866), .ZN(n6949) );
  OR2_X1 U7613 ( .A1(n7786), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n7806) );
  NAND2_X1 U7614 ( .A1(n12701), .A2(n7730), .ZN(n12688) );
  AND2_X1 U7615 ( .A1(n8876), .A2(n7928), .ZN(n8869) );
  NAND2_X1 U7616 ( .A1(n7618), .A2(n7617), .ZN(n7634) );
  INV_X1 U7617 ( .A(n7619), .ZN(n7618) );
  INV_X1 U7618 ( .A(n10790), .ZN(n8821) );
  NAND2_X1 U7619 ( .A1(n8827), .A2(n8826), .ZN(n7562) );
  AND2_X1 U7620 ( .A1(n10423), .A2(n8813), .ZN(n10522) );
  NAND3_X1 U7621 ( .A1(n14914), .A2(n7436), .A3(n7435), .ZN(n10142) );
  NAND2_X1 U7622 ( .A1(n7927), .A2(n6949), .ZN(n6948) );
  NOR2_X1 U7623 ( .A1(n10999), .A2(n8771), .ZN(n6942) );
  AND2_X1 U7624 ( .A1(n7289), .A2(n7288), .ZN(n7287) );
  INV_X1 U7625 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7288) );
  INV_X1 U7626 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n7351) );
  INV_X1 U7627 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n7350) );
  INV_X1 U7628 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n7354) );
  INV_X1 U7629 ( .A(n7032), .ZN(n7031) );
  OAI21_X1 U7630 ( .B1(n7663), .B2(n7033), .A(n7697), .ZN(n7032) );
  INV_X1 U7631 ( .A(n7677), .ZN(n7033) );
  INV_X1 U7632 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n8304) );
  INV_X1 U7633 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n8300) );
  NAND2_X1 U7634 ( .A1(n7608), .A2(n7607), .ZN(n7626) );
  NOR2_X1 U7635 ( .A1(n7039), .A2(n7588), .ZN(n7038) );
  INV_X1 U7636 ( .A(n7040), .ZN(n7039) );
  NOR2_X1 U7637 ( .A1(n7044), .A2(n7588), .ZN(n7036) );
  INV_X1 U7638 ( .A(n12970), .ZN(n7239) );
  INV_X1 U7639 ( .A(n12996), .ZN(n7238) );
  BUF_X1 U7640 ( .A(n9858), .Z(n12960) );
  INV_X1 U7641 ( .A(n9330), .ZN(n9378) );
  AND2_X1 U7642 ( .A1(n12055), .A2(n12054), .ZN(n12057) );
  OR2_X1 U7643 ( .A1(n11557), .A2(n11556), .ZN(n11910) );
  OR2_X1 U7644 ( .A1(n9969), .A2(n9968), .ZN(n10085) );
  INV_X1 U7645 ( .A(n11629), .ZN(n9350) );
  INV_X1 U7646 ( .A(n9348), .ZN(n9349) );
  OR2_X1 U7647 ( .A1(n11290), .A2(n11289), .ZN(n11353) );
  AND2_X2 U7648 ( .A1(n9378), .A2(n12062), .ZN(n11803) );
  NOR2_X1 U7649 ( .A1(n12035), .A2(n7114), .ZN(n7113) );
  INV_X1 U7650 ( .A(n10257), .ZN(n7114) );
  NAND2_X1 U7651 ( .A1(n6622), .A2(n13154), .ZN(n9560) );
  XNOR2_X1 U7652 ( .A(n11803), .B(n12063), .ZN(n6622) );
  NAND2_X1 U7653 ( .A1(n6773), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6772) );
  INV_X1 U7655 ( .A(n9140), .ZN(n8978) );
  AND2_X1 U7656 ( .A1(n8984), .A2(n8972), .ZN(n8980) );
  INV_X1 U7657 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8972) );
  INV_X1 U7658 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n9138) );
  NOR2_X1 U7659 ( .A1(n9200), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n9618) );
  NOR2_X1 U7660 ( .A1(n13786), .A2(n6824), .ZN(n6823) );
  INV_X1 U7661 ( .A(n6883), .ZN(n6882) );
  OAI21_X1 U7662 ( .B1(n6884), .B2(n12095), .A(n6575), .ZN(n6883) );
  NOR2_X1 U7663 ( .A1(n12108), .A2(n6980), .ZN(n6979) );
  INV_X1 U7664 ( .A(n12107), .ZN(n6980) );
  INV_X1 U7665 ( .A(n6981), .ZN(n6977) );
  OR2_X1 U7666 ( .A1(n8688), .A2(n13938), .ZN(n12085) );
  AND2_X1 U7667 ( .A1(n13917), .A2(n12105), .ZN(n6981) );
  INV_X1 U7668 ( .A(n6965), .ZN(n6964) );
  OAI21_X1 U7669 ( .B1(n11463), .B2(n6966), .A(n6539), .ZN(n6965) );
  INV_X1 U7670 ( .A(n12100), .ZN(n6966) );
  OR2_X1 U7671 ( .A1(n11226), .A2(n6843), .ZN(n6842) );
  INV_X1 U7672 ( .A(n11380), .ZN(n6840) );
  INV_X1 U7673 ( .A(n11189), .ZN(n6843) );
  OR2_X1 U7674 ( .A1(n11174), .A2(n12166), .ZN(n11380) );
  OR2_X1 U7675 ( .A1(n6832), .A2(n14390), .ZN(n6831) );
  NAND2_X1 U7676 ( .A1(n6833), .A2(n11538), .ZN(n6832) );
  NAND2_X1 U7677 ( .A1(n10630), .A2(n10629), .ZN(n6855) );
  AOI21_X1 U7678 ( .B1(n10628), .B2(n10627), .A(n10626), .ZN(n10950) );
  NAND2_X1 U7679 ( .A1(n6846), .A2(n10285), .ZN(n6845) );
  INV_X1 U7680 ( .A(n6850), .ZN(n6846) );
  NOR2_X1 U7681 ( .A1(n13547), .A2(n14521), .ZN(n6852) );
  NAND2_X1 U7682 ( .A1(n13838), .A2(n14099), .ZN(n13811) );
  OR2_X1 U7683 ( .A1(n13918), .A2(n13917), .ZN(n13920) );
  AND2_X1 U7684 ( .A1(n6955), .A2(n10294), .ZN(n6953) );
  INV_X1 U7685 ( .A(n10586), .ZN(n9272) );
  INV_X1 U7686 ( .A(n7210), .ZN(n7209) );
  AND2_X1 U7687 ( .A1(n7216), .A2(n7214), .ZN(n7213) );
  NAND2_X1 U7688 ( .A1(n7221), .A2(n7217), .ZN(n7216) );
  AND3_X1 U7689 ( .A1(n8728), .A2(n8037), .A3(n8000), .ZN(n7341) );
  INV_X1 U7690 ( .A(n7206), .ZN(n7205) );
  OAI21_X1 U7691 ( .B1(n8401), .B2(n7207), .A(n8411), .ZN(n7206) );
  NAND3_X1 U7692 ( .A1(n8396), .A2(n8399), .A3(n8395), .ZN(n8402) );
  NAND2_X1 U7693 ( .A1(n8358), .A2(n8359), .ZN(n6730) );
  OR2_X1 U7694 ( .A1(n8305), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n8306) );
  OAI21_X1 U7695 ( .B1(n9335), .B2(n6819), .A(n6818), .ZN(n6817) );
  NAND2_X1 U7696 ( .A1(n9335), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n6818) );
  OAI211_X1 U7697 ( .C1(n9377), .C2(n7186), .A(n7184), .B(n7183), .ZN(n8028)
         );
  NAND2_X1 U7698 ( .A1(n7185), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7184) );
  AND2_X1 U7699 ( .A1(n14139), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n7071) );
  XNOR2_X1 U7700 ( .A(n14144), .B(n14143), .ZN(n14164) );
  AND2_X1 U7701 ( .A1(n6702), .A2(n6573), .ZN(n14163) );
  NAND2_X1 U7702 ( .A1(n6703), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n6702) );
  INV_X1 U7703 ( .A(n14190), .ZN(n6703) );
  OAI21_X1 U7704 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n14151), .A(n14150), .ZN(
        n14153) );
  AOI21_X1 U7705 ( .B1(n12356), .B2(n7012), .A(n6519), .ZN(n7011) );
  INV_X1 U7706 ( .A(n11674), .ZN(n7012) );
  OR2_X1 U7707 ( .A1(n7545), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n7529) );
  NAND2_X1 U7708 ( .A1(n11639), .A2(n11638), .ZN(n7014) );
  NAND2_X1 U7709 ( .A1(n7021), .A2(n7017), .ZN(n7016) );
  INV_X1 U7710 ( .A(n11277), .ZN(n7003) );
  NAND2_X1 U7711 ( .A1(n11208), .A2(n11064), .ZN(n6989) );
  INV_X1 U7712 ( .A(n9890), .ZN(n14927) );
  AOI211_X1 U7713 ( .C1(n9759), .C2(n9897), .A(n9896), .B(n9895), .ZN(n9898)
         );
  INV_X1 U7714 ( .A(n7687), .ZN(n7686) );
  AOI21_X1 U7715 ( .B1(n6999), .B2(n7000), .A(n6997), .ZN(n6996) );
  INV_X1 U7716 ( .A(n11572), .ZN(n6997) );
  INV_X1 U7717 ( .A(n6999), .ZN(n6998) );
  AND4_X1 U7718 ( .A1(n7518), .A2(n7517), .A3(n7516), .A4(n7515), .ZN(n10791)
         );
  NAND2_X1 U7719 ( .A1(n10853), .A2(n10852), .ZN(n6915) );
  NAND2_X1 U7720 ( .A1(n14769), .A2(n10869), .ZN(n14788) );
  NAND2_X1 U7721 ( .A1(n14788), .A2(n14787), .ZN(n14786) );
  NAND2_X1 U7722 ( .A1(n6915), .A2(n14766), .ZN(n6914) );
  XNOR2_X1 U7723 ( .A(n10870), .B(n10893), .ZN(n14806) );
  NAND2_X1 U7724 ( .A1(n14824), .A2(n14823), .ZN(n14822) );
  XNOR2_X1 U7725 ( .A(n10872), .B(n10903), .ZN(n14842) );
  OR2_X1 U7726 ( .A1(n14811), .A2(n6913), .ZN(n6912) );
  NOR2_X1 U7727 ( .A1(n10897), .A2(n10857), .ZN(n6913) );
  NAND2_X1 U7728 ( .A1(n14860), .A2(n14859), .ZN(n14858) );
  OR2_X1 U7729 ( .A1(n14847), .A2(n6906), .ZN(n6905) );
  NOR2_X1 U7730 ( .A1(n10908), .A2(n10907), .ZN(n6906) );
  XNOR2_X1 U7731 ( .A(n10874), .B(n10914), .ZN(n14881) );
  NAND2_X1 U7732 ( .A1(n14887), .A2(n14888), .ZN(n14886) );
  XNOR2_X1 U7733 ( .A(n11077), .B(n10864), .ZN(n10877) );
  NAND2_X1 U7734 ( .A1(n11080), .A2(n11081), .ZN(n12389) );
  AOI21_X1 U7735 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n12387), .A(n12386), .ZN(
        n12406) );
  XNOR2_X1 U7736 ( .A(n12410), .B(n12407), .ZN(n12390) );
  INV_X1 U7737 ( .A(n6647), .ZN(n6646) );
  OAI22_X1 U7738 ( .A1(n6654), .A2(n12538), .B1(n12537), .B2(n12789), .ZN(
        n6647) );
  NAND2_X1 U7739 ( .A1(n7934), .A2(n8899), .ZN(n12595) );
  OAI21_X1 U7740 ( .B1(n12640), .B2(n6921), .A(n6919), .ZN(n7934) );
  OAI21_X1 U7741 ( .B1(n6487), .B2(n6921), .A(n8895), .ZN(n6920) );
  OR2_X1 U7742 ( .A1(n12681), .A2(n12690), .ZN(n12663) );
  AND2_X1 U7743 ( .A1(n12663), .A2(n12662), .ZN(n12680) );
  NAND2_X1 U7744 ( .A1(n7741), .A2(n7740), .ZN(n11652) );
  NAND2_X1 U7745 ( .A1(n11474), .A2(n11478), .ZN(n12730) );
  AND4_X1 U7746 ( .A1(n7657), .A2(n7656), .A3(n7655), .A4(n7654), .ZN(n11601)
         );
  OAI21_X1 U7747 ( .B1(n11249), .B2(n8853), .A(n8850), .ZN(n11397) );
  NAND2_X1 U7748 ( .A1(n7606), .A2(n7280), .ZN(n7279) );
  NOR2_X1 U7749 ( .A1(n6552), .A2(n7281), .ZN(n7280) );
  INV_X1 U7750 ( .A(n7605), .ZN(n7281) );
  CLKBUF_X1 U7751 ( .A(n11250), .Z(n11392) );
  AND4_X1 U7752 ( .A1(n7583), .A2(n7582), .A3(n7581), .A4(n7580), .ZN(n10998)
         );
  NAND2_X1 U7753 ( .A1(n10741), .A2(n7570), .ZN(n14302) );
  AND2_X1 U7754 ( .A1(n8801), .A2(n8802), .ZN(n10145) );
  OR2_X1 U7755 ( .A1(n9757), .A2(n8948), .ZN(n14919) );
  INV_X1 U7756 ( .A(n8793), .ZN(n14915) );
  INV_X1 U7757 ( .A(n14919), .ZN(n14286) );
  INV_X1 U7758 ( .A(n14303), .ZN(n14922) );
  NAND2_X1 U7759 ( .A1(n7880), .A2(n7879), .ZN(n7985) );
  NAND2_X1 U7760 ( .A1(n7703), .A2(n7702), .ZN(n12345) );
  NAND2_X1 U7761 ( .A1(n7684), .A2(n7683), .ZN(n12314) );
  INV_X1 U7762 ( .A(n11608), .ZN(n12795) );
  INV_X1 U7763 ( .A(n8759), .ZN(n7721) );
  NOR2_X1 U7764 ( .A1(n8955), .A2(n7982), .ZN(n9301) );
  AND2_X1 U7765 ( .A1(n12867), .A2(n9292), .ZN(n9526) );
  NAND2_X1 U7766 ( .A1(n7943), .A2(n7977), .ZN(n14979) );
  NAND2_X1 U7767 ( .A1(n9757), .A2(n9528), .ZN(n14917) );
  NAND2_X1 U7768 ( .A1(n7064), .A2(n7065), .ZN(n7874) );
  AOI21_X1 U7769 ( .B1(n7066), .B2(n7844), .A(n6611), .ZN(n7065) );
  NAND2_X1 U7770 ( .A1(n7289), .A2(n7358), .ZN(n6917) );
  XNOR2_X1 U7771 ( .A(n7954), .B(P3_IR_REG_26__SCAN_IN), .ZN(n7975) );
  AND2_X1 U7772 ( .A1(n7275), .A2(n7332), .ZN(n6918) );
  OR2_X1 U7773 ( .A1(n7800), .A2(n11979), .ZN(n7813) );
  INV_X1 U7774 ( .A(n7055), .ZN(n7054) );
  OAI21_X1 U7775 ( .B1(n7767), .B2(n7056), .A(n7781), .ZN(n7055) );
  OR2_X1 U7776 ( .A1(n7735), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7059) );
  INV_X1 U7777 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n7887) );
  NAND2_X1 U7778 ( .A1(n7664), .A2(n7663), .ZN(n7678) );
  NAND2_X1 U7779 ( .A1(n7048), .A2(n7047), .ZN(n7661) );
  NOR2_X1 U7780 ( .A1(n7321), .A2(n6602), .ZN(n7047) );
  XNOR2_X1 U7781 ( .A(n7626), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n7609) );
  AOI21_X1 U7782 ( .B1(n7044), .B2(n7042), .A(n7041), .ZN(n7040) );
  INV_X1 U7783 ( .A(n7333), .ZN(n7042) );
  INV_X1 U7784 ( .A(n7571), .ZN(n7041) );
  NAND2_X1 U7785 ( .A1(n7505), .A2(n7333), .ZN(n7045) );
  AOI21_X1 U7786 ( .B1(n7063), .B2(n7061), .A(n6561), .ZN(n7060) );
  INV_X1 U7787 ( .A(n7063), .ZN(n7062) );
  OR2_X1 U7788 ( .A1(n7551), .A2(n7550), .ZN(n7553) );
  NAND2_X1 U7789 ( .A1(n7023), .A2(n7024), .ZN(n7490) );
  INV_X1 U7790 ( .A(n7025), .ZN(n7024) );
  OAI21_X1 U7791 ( .B1(n7447), .B2(n7026), .A(n7470), .ZN(n7025) );
  NAND2_X1 U7792 ( .A1(n7027), .A2(n7447), .ZN(n7467) );
  INV_X1 U7793 ( .A(n7449), .ZN(n7027) );
  NAND2_X1 U7794 ( .A1(n7392), .A2(n7391), .ZN(n7058) );
  NAND2_X1 U7795 ( .A1(n11128), .A2(n11129), .ZN(n11331) );
  XNOR2_X1 U7796 ( .A(n12911), .B(n14634), .ZN(n9645) );
  AOI21_X1 U7797 ( .B1(n12896), .B2(n12895), .A(n7328), .ZN(n12947) );
  NAND2_X1 U7798 ( .A1(n6500), .A2(n12963), .ZN(n7270) );
  NOR2_X1 U7799 ( .A1(n7269), .A2(n7268), .ZN(n7267) );
  NOR2_X1 U7800 ( .A1(n12963), .A2(n6500), .ZN(n7268) );
  NOR2_X1 U7801 ( .A1(n7271), .A2(n7270), .ZN(n7269) );
  AOI21_X1 U7802 ( .B1(n12996), .B2(n7244), .A(n7243), .ZN(n7242) );
  INV_X1 U7803 ( .A(n12902), .ZN(n7244) );
  INV_X1 U7804 ( .A(n12908), .ZN(n7243) );
  NAND2_X1 U7805 ( .A1(n10653), .A2(n10652), .ZN(n7248) );
  AND2_X1 U7806 ( .A1(n11500), .A2(n11503), .ZN(n7245) );
  INV_X1 U7807 ( .A(n9639), .ZN(n7224) );
  AND2_X1 U7808 ( .A1(n10080), .A2(n10078), .ZN(n7249) );
  NAND2_X1 U7809 ( .A1(n10077), .A2(n10076), .ZN(n10079) );
  NAND2_X1 U7810 ( .A1(n7232), .A2(n7235), .ZN(n7231) );
  INV_X1 U7811 ( .A(n13222), .ZN(n13195) );
  INV_X1 U7812 ( .A(n11803), .ZN(n12021) );
  AND2_X1 U7813 ( .A1(n9348), .A2(n9350), .ZN(n9387) );
  NAND2_X1 U7814 ( .A1(n11709), .A2(n11708), .ZN(n13166) );
  AND2_X1 U7815 ( .A1(n6814), .A2(n7125), .ZN(n13243) );
  AND2_X1 U7816 ( .A1(n7125), .A2(n13242), .ZN(n6812) );
  NAND2_X1 U7817 ( .A1(n13286), .A2(n13192), .ZN(n7124) );
  INV_X1 U7818 ( .A(n13219), .ZN(n13285) );
  NAND2_X1 U7819 ( .A1(n13217), .A2(n13216), .ZN(n13290) );
  NOR2_X2 U7820 ( .A1(n13332), .A2(n13432), .ZN(n13318) );
  NAND2_X1 U7821 ( .A1(n13350), .A2(n13184), .ZN(n13325) );
  OAI21_X1 U7822 ( .B1(n13363), .B2(n13181), .A(n13182), .ZN(n13348) );
  NAND2_X1 U7823 ( .A1(n13383), .A2(n13175), .ZN(n6768) );
  NAND2_X1 U7824 ( .A1(n11545), .A2(n6529), .ZN(n13174) );
  NAND2_X1 U7825 ( .A1(n6716), .A2(n6477), .ZN(n11426) );
  NAND2_X1 U7826 ( .A1(n10721), .A2(n10720), .ZN(n11867) );
  NAND2_X1 U7827 ( .A1(n10821), .A2(n11055), .ZN(n11163) );
  INV_X1 U7828 ( .A(n12041), .ZN(n11154) );
  OAI21_X1 U7829 ( .B1(n6804), .B2(n10263), .A(n6802), .ZN(n10544) );
  INV_X1 U7830 ( .A(n6805), .ZN(n6804) );
  AOI21_X1 U7831 ( .B1(n6805), .B2(n6803), .A(n6546), .ZN(n6802) );
  NAND2_X1 U7832 ( .A1(n10544), .A2(n12036), .ZN(n10752) );
  AOI21_X1 U7833 ( .B1(n6809), .B2(n10262), .A(n6507), .ZN(n6808) );
  NAND2_X1 U7834 ( .A1(n10263), .A2(n6809), .ZN(n6807) );
  NAND2_X1 U7835 ( .A1(n10686), .A2(n9990), .ZN(n9992) );
  NAND2_X1 U7836 ( .A1(n9992), .A2(n9991), .ZN(n10258) );
  OAI21_X1 U7837 ( .B1(n7108), .B2(n12027), .A(n9989), .ZN(n7107) );
  NAND2_X1 U7838 ( .A1(n7102), .A2(n7101), .ZN(n10686) );
  NOR2_X1 U7839 ( .A1(n7107), .A2(n12029), .ZN(n7101) );
  NAND2_X1 U7840 ( .A1(n9987), .A2(n9986), .ZN(n10196) );
  AND2_X1 U7841 ( .A1(n9565), .A2(n9562), .ZN(n12026) );
  AND2_X1 U7842 ( .A1(n12063), .A2(n9330), .ZN(n10173) );
  NAND2_X1 U7843 ( .A1(n11920), .A2(n11919), .ZN(n13452) );
  NAND2_X1 U7844 ( .A1(n11900), .A2(n11899), .ZN(n13459) );
  NAND2_X1 U7845 ( .A1(n11429), .A2(n11428), .ZN(n13472) );
  NAND2_X1 U7846 ( .A1(n11116), .A2(n11115), .ZN(n13487) );
  AND2_X1 U7847 ( .A1(n9309), .A2(n9307), .ZN(n14654) );
  NAND3_X1 U7848 ( .A1(n8969), .A2(n7323), .A3(n7170), .ZN(n9345) );
  NOR2_X1 U7849 ( .A1(n9140), .A2(n7171), .ZN(n7170) );
  NAND2_X1 U7850 ( .A1(n6773), .A2(n7172), .ZN(n7171) );
  NAND2_X1 U7851 ( .A1(n8980), .A2(n8974), .ZN(n8982) );
  NOR2_X1 U7852 ( .A1(n9136), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n8984) );
  AOI22_X1 U7853 ( .A1(n6474), .A2(n6467), .B1(n9326), .B2(n9884), .ZN(n7136)
         );
  NAND2_X1 U7854 ( .A1(n6897), .A2(n6549), .ZN(n6896) );
  NAND2_X1 U7855 ( .A1(n13528), .A2(n6898), .ZN(n6897) );
  NOR2_X1 U7856 ( .A1(n6896), .A2(n6895), .ZN(n6894) );
  INV_X1 U7857 ( .A(n12246), .ZN(n6895) );
  NAND2_X1 U7858 ( .A1(n13552), .A2(n12212), .ZN(n6673) );
  AOI21_X1 U7859 ( .B1(n6672), .B2(n6670), .A(n6518), .ZN(n6669) );
  INV_X1 U7860 ( .A(n12212), .ZN(n6670) );
  INV_X1 U7861 ( .A(n6672), .ZN(n6671) );
  AND2_X1 U7862 ( .A1(n11319), .A2(n6596), .ZN(n6680) );
  OR2_X1 U7863 ( .A1(n9802), .A2(n9801), .ZN(n9807) );
  AND2_X1 U7864 ( .A1(n9280), .A2(n9692), .ZN(n9816) );
  AND4_X1 U7865 ( .A1(n8651), .A2(n8650), .A3(n8649), .A4(n8648), .ZN(n12273)
         );
  NOR2_X1 U7866 ( .A1(n11515), .A2(n11373), .ZN(n6682) );
  AND2_X1 U7867 ( .A1(n6688), .A2(n6687), .ZN(n13735) );
  NAND2_X1 U7868 ( .A1(n13733), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6687) );
  OR2_X1 U7869 ( .A1(n13735), .A2(n13734), .ZN(n6686) );
  NAND2_X1 U7870 ( .A1(n6876), .A2(n6878), .ZN(n6874) );
  AOI21_X1 U7871 ( .B1(n6882), .B2(n12095), .A(n6881), .ZN(n6880) );
  INV_X1 U7872 ( .A(n12138), .ZN(n6881) );
  AND2_X1 U7873 ( .A1(n6882), .A2(n6877), .ZN(n6876) );
  NAND2_X1 U7874 ( .A1(n13809), .A2(n13788), .ZN(n6877) );
  INV_X1 U7875 ( .A(n6973), .ZN(n6972) );
  NOR2_X1 U7876 ( .A1(n6575), .A2(n6974), .ZN(n6973) );
  INV_X1 U7877 ( .A(n12119), .ZN(n6974) );
  NAND2_X1 U7878 ( .A1(n6879), .A2(n6882), .ZN(n12139) );
  OR2_X1 U7879 ( .A1(n6885), .A2(n12095), .ZN(n6879) );
  INV_X1 U7880 ( .A(n13657), .ZN(n13794) );
  AND2_X1 U7881 ( .A1(n6885), .A2(n6884), .ZN(n13790) );
  AND2_X1 U7882 ( .A1(n13849), .A2(n12111), .ZN(n6983) );
  NOR2_X1 U7883 ( .A1(n13889), .A2(n13869), .ZN(n6836) );
  NAND2_X1 U7884 ( .A1(n6836), .A2(n14104), .ZN(n13856) );
  NAND2_X1 U7885 ( .A1(n13887), .A2(n8687), .ZN(n13889) );
  NAND2_X1 U7886 ( .A1(n12106), .A2(n6981), .ZN(n13915) );
  AND2_X1 U7887 ( .A1(n6863), .A2(n7318), .ZN(n6862) );
  NAND2_X1 U7888 ( .A1(n6858), .A2(n6857), .ZN(n6863) );
  NAND2_X1 U7889 ( .A1(n12079), .A2(n12078), .ZN(n13981) );
  NAND2_X1 U7890 ( .A1(n11464), .A2(n11463), .ZN(n12101) );
  NAND2_X1 U7891 ( .A1(n10950), .A2(n10949), .ZN(n10948) );
  XNOR2_X1 U7892 ( .A(n8691), .B(n10463), .ZN(n10456) );
  INV_X1 U7893 ( .A(n13983), .ZN(n13955) );
  NAND2_X1 U7894 ( .A1(n8683), .A2(n8682), .ZN(n13773) );
  NAND2_X1 U7895 ( .A1(n8640), .A2(n8639), .ZN(n13781) );
  NAND2_X1 U7896 ( .A1(n8366), .A2(n8365), .ZN(n14397) );
  NAND2_X1 U7897 ( .A1(n8331), .A2(n8330), .ZN(n11621) );
  INV_X1 U7898 ( .A(n10463), .ZN(n14504) );
  AND2_X1 U7899 ( .A1(n9270), .A2(n9269), .ZN(n10302) );
  NOR2_X1 U7900 ( .A1(n10308), .A2(n9267), .ZN(n10156) );
  INV_X1 U7901 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8016) );
  NAND2_X1 U7902 ( .A1(n8001), .A2(n7341), .ZN(n8734) );
  NOR2_X1 U7903 ( .A1(n8730), .A2(n8729), .ZN(n8735) );
  NAND2_X1 U7904 ( .A1(n8043), .A2(n6541), .ZN(n8726) );
  INV_X1 U7905 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6903) );
  INV_X1 U7906 ( .A(n6721), .ZN(n8343) );
  AOI21_X1 U7907 ( .B1(n7198), .B2(n6722), .A(n6725), .ZN(n6721) );
  INV_X1 U7908 ( .A(n6726), .ZN(n6722) );
  NAND2_X1 U7909 ( .A1(n7198), .A2(n7199), .ZN(n8297) );
  OAI21_X1 U7910 ( .B1(n6753), .B2(n8230), .A(n6751), .ZN(n8236) );
  INV_X1 U7911 ( .A(n6752), .ZN(n6751) );
  NAND2_X1 U7912 ( .A1(n8236), .A2(n8235), .ZN(n8259) );
  NAND2_X1 U7913 ( .A1(n6817), .A2(SI_6_), .ZN(n8185) );
  NAND2_X1 U7914 ( .A1(n8110), .A2(n8109), .ZN(n8141) );
  NAND2_X1 U7915 ( .A1(n8092), .A2(n8093), .ZN(n8091) );
  NAND2_X1 U7916 ( .A1(n14170), .A2(n14171), .ZN(n14174) );
  XNOR2_X1 U7917 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(n14164), .ZN(n14165) );
  INV_X1 U7918 ( .A(n6708), .ZN(n14186) );
  OAI21_X1 U7919 ( .B1(n14181), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n6567), .ZN(
        n6708) );
  NAND2_X1 U7920 ( .A1(n6638), .A2(n14193), .ZN(n14194) );
  INV_X1 U7921 ( .A(n6709), .ZN(n14210) );
  OAI21_X1 U7922 ( .B1(n14160), .B2(n14159), .A(n6710), .ZN(n6709) );
  NAND2_X1 U7923 ( .A1(n14154), .A2(P1_ADDR_REG_11__SCAN_IN), .ZN(n6710) );
  OR2_X1 U7924 ( .A1(n14423), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n7089) );
  NAND2_X1 U7925 ( .A1(n14423), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n7087) );
  AOI21_X1 U7926 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(n14158), .A(n14157), .ZN(
        n14217) );
  NAND2_X1 U7927 ( .A1(n14221), .A2(n14220), .ZN(n7080) );
  NOR2_X1 U7928 ( .A1(n14436), .A2(n7081), .ZN(n14232) );
  NAND2_X1 U7929 ( .A1(n14227), .A2(n7077), .ZN(n7076) );
  OR2_X1 U7930 ( .A1(n14438), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n7074) );
  NAND2_X1 U7931 ( .A1(n7785), .A2(n7784), .ZN(n12766) );
  AND3_X1 U7932 ( .A1(n7746), .A2(n7745), .A3(n7744), .ZN(n12677) );
  INV_X1 U7933 ( .A(n7009), .ZN(n7008) );
  INV_X1 U7934 ( .A(n12614), .ZN(n12309) );
  NAND2_X1 U7935 ( .A1(n7803), .A2(n7802), .ZN(n12634) );
  AND4_X1 U7936 ( .A1(n7639), .A2(n7638), .A3(n7637), .A4(n7636), .ZN(n11574)
         );
  AND4_X1 U7937 ( .A1(n7692), .A2(n7691), .A3(n7690), .A4(n7689), .ZN(n12721)
         );
  INV_X1 U7938 ( .A(n12865), .ZN(n11580) );
  NAND2_X1 U7939 ( .A1(n6569), .A2(n6616), .ZN(n6632) );
  NAND2_X1 U7940 ( .A1(n8939), .A2(n8938), .ZN(n6616) );
  INV_X1 U7941 ( .A(n12677), .ZN(n12704) );
  INV_X1 U7942 ( .A(n11601), .ZN(n12373) );
  INV_X1 U7943 ( .A(n10998), .ZN(n12375) );
  OAI21_X1 U7944 ( .B1(n14766), .B2(n6915), .A(n6914), .ZN(n14760) );
  NOR2_X1 U7945 ( .A1(n14760), .A2(n10881), .ZN(n14759) );
  NOR2_X1 U7946 ( .A1(n14813), .A2(n14812), .ZN(n14811) );
  XNOR2_X1 U7947 ( .A(n6912), .B(n14838), .ZN(n14830) );
  NOR2_X1 U7948 ( .A1(n14830), .A2(n14831), .ZN(n14829) );
  INV_X1 U7949 ( .A(n7985), .ZN(n12557) );
  AND2_X1 U7950 ( .A1(n12551), .A2(n14323), .ZN(n7944) );
  NOR2_X1 U7951 ( .A1(n7908), .A2(n7907), .ZN(n7909) );
  AOI21_X1 U7952 ( .B1(n12746), .B2(n14323), .A(n6951), .ZN(n12822) );
  OR2_X1 U7953 ( .A1(n14991), .A2(n14979), .ZN(n12864) );
  AND2_X1 U7954 ( .A1(n9527), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12867) );
  XNOR2_X1 U7955 ( .A(n7890), .B(P3_IR_REG_22__SCAN_IN), .ZN(n10535) );
  NAND2_X1 U7956 ( .A1(n10123), .A2(n10122), .ZN(n14720) );
  XNOR2_X1 U7957 ( .A(n9645), .B(n9644), .ZN(n9719) );
  NOR2_X1 U7958 ( .A1(n7262), .A2(n13018), .ZN(n7260) );
  NOR2_X1 U7959 ( .A1(n7263), .A2(n7265), .ZN(n7262) );
  NOR2_X1 U7960 ( .A1(n12963), .A2(n7266), .ZN(n7265) );
  INV_X1 U7961 ( .A(n7267), .ZN(n7263) );
  NAND2_X1 U7962 ( .A1(n7267), .A2(n7270), .ZN(n7264) );
  NAND2_X1 U7963 ( .A1(n13033), .A2(n13032), .ZN(n13031) );
  NAND2_X1 U7964 ( .A1(n11936), .A2(n11935), .ZN(n13447) );
  NAND2_X1 U7965 ( .A1(n12003), .A2(n12002), .ZN(n13304) );
  NAND2_X1 U7966 ( .A1(n11350), .A2(n11349), .ZN(n13476) );
  NAND2_X1 U7967 ( .A1(n9681), .A2(n9661), .ZN(n9662) );
  NAND2_X1 U7968 ( .A1(n11541), .A2(n11540), .ZN(n13466) );
  NAND2_X1 U7969 ( .A1(n6749), .A2(n11288), .ZN(n13481) );
  NAND2_X1 U7970 ( .A1(n11286), .A2(n9951), .ZN(n6749) );
  AND2_X1 U7971 ( .A1(n9675), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13025) );
  AND2_X1 U7972 ( .A1(n9165), .A2(n13525), .ZN(n14586) );
  NAND2_X1 U7973 ( .A1(n13233), .A2(n13232), .ZN(n13405) );
  AOI21_X1 U7974 ( .B1(n13224), .B2(n13004), .A(n13231), .ZN(n13232) );
  NAND2_X1 U7975 ( .A1(n6775), .A2(n13188), .ZN(n13296) );
  NAND2_X1 U7976 ( .A1(n7226), .A2(n10065), .ZN(n7225) );
  NAND2_X1 U7977 ( .A1(n7228), .A2(n7227), .ZN(n7226) );
  NAND2_X1 U7978 ( .A1(n13197), .A2(n7121), .ZN(n7120) );
  NOR2_X1 U7979 ( .A1(n13197), .A2(n7121), .ZN(n7119) );
  AND2_X1 U7980 ( .A1(n13410), .A2(n14711), .ZN(n7142) );
  NAND2_X1 U7981 ( .A1(n9343), .A2(n9342), .ZN(n13515) );
  INV_X1 U7982 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n9342) );
  INV_X1 U7983 ( .A(n9345), .ZN(n9343) );
  NAND2_X1 U7984 ( .A1(n6677), .A2(n12254), .ZN(n6676) );
  NAND2_X1 U7985 ( .A1(n6899), .A2(n6499), .ZN(n6677) );
  INV_X1 U7986 ( .A(n13528), .ZN(n6675) );
  NAND2_X1 U7987 ( .A1(n13596), .A2(n12215), .ZN(n13564) );
  NAND2_X1 U7988 ( .A1(n14385), .A2(n6532), .ZN(n11617) );
  NAND2_X1 U7989 ( .A1(n14385), .A2(n11526), .ZN(n11528) );
  AND2_X1 U7990 ( .A1(n8393), .A2(n8392), .ZN(n14366) );
  INV_X1 U7991 ( .A(n6889), .ZN(n6887) );
  INV_X1 U7992 ( .A(n10606), .ZN(n6888) );
  AOI21_X1 U7993 ( .B1(n6890), .B2(n6468), .A(n6521), .ZN(n6889) );
  NAND2_X1 U7994 ( .A1(n14136), .A2(n9084), .ZN(n8687) );
  NAND2_X1 U7995 ( .A1(n10111), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14394) );
  NAND2_X1 U7996 ( .A1(n9828), .A2(n14483), .ZN(n14389) );
  INV_X1 U7997 ( .A(n12273), .ZN(n13656) );
  OR2_X1 U7998 ( .A1(n10979), .A2(n10978), .ZN(n6688) );
  OR2_X1 U7999 ( .A1(n9211), .A2(n9424), .ZN(n13764) );
  OAI21_X1 U8000 ( .B1(n13765), .B2(n13764), .A(n6691), .ZN(n6690) );
  OR2_X1 U8001 ( .A1(n13767), .A2(n14451), .ZN(n6691) );
  OAI21_X1 U8002 ( .B1(n8428), .B2(P1_IR_REG_18__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8036) );
  OR2_X1 U8003 ( .A1(n9827), .A2(n10305), .ZN(n14483) );
  INV_X1 U8004 ( .A(n11538), .ZN(n11266) );
  NAND2_X1 U8005 ( .A1(n8270), .A2(n8269), .ZN(n11327) );
  XNOR2_X1 U8006 ( .A(n14174), .B(n6641), .ZN(n14254) );
  INV_X1 U8007 ( .A(n14175), .ZN(n6641) );
  NOR2_X1 U8008 ( .A1(n14221), .A2(n14220), .ZN(n14433) );
  AND3_X1 U8009 ( .A1(n8106), .A2(n8105), .A3(n8104), .ZN(n7319) );
  NAND2_X1 U8010 ( .A1(n7291), .A2(n8149), .ZN(n7290) );
  NAND2_X1 U8011 ( .A1(n8196), .A2(n7315), .ZN(n7314) );
  NAND2_X1 U8012 ( .A1(n6633), .A2(n8793), .ZN(n8798) );
  OR2_X1 U8013 ( .A1(n8794), .A2(n8948), .ZN(n6633) );
  INV_X1 U8014 ( .A(n11832), .ZN(n7181) );
  NOR2_X1 U8015 ( .A1(n11832), .A2(n11835), .ZN(n7182) );
  AND2_X1 U8016 ( .A1(n8351), .A2(n8347), .ZN(n8348) );
  NAND2_X1 U8017 ( .A1(n6738), .A2(n6739), .ZN(n11854) );
  MUX2_X1 U8018 ( .A(n8816), .B(n8815), .S(n9528), .Z(n8820) );
  AOI21_X1 U8019 ( .B1(n6736), .B2(n6472), .A(n6734), .ZN(n6733) );
  OAI211_X1 U8020 ( .C1(n12102), .C2(n8421), .A(n8424), .B(n6559), .ZN(n7302)
         );
  AND2_X1 U8021 ( .A1(n13931), .A2(n7304), .ZN(n7303) );
  NAND2_X1 U8022 ( .A1(n8453), .A2(n6504), .ZN(n7304) );
  OAI21_X1 U8023 ( .B1(n8844), .B2(n8843), .A(n8842), .ZN(n8849) );
  NAND2_X1 U8024 ( .A1(n11887), .A2(n11884), .ZN(n7157) );
  INV_X1 U8025 ( .A(n11876), .ZN(n7175) );
  NOR2_X1 U8026 ( .A1(n11879), .A2(n11876), .ZN(n7176) );
  AND2_X1 U8027 ( .A1(n11882), .A2(n6748), .ZN(n6747) );
  INV_X1 U8028 ( .A(n11880), .ZN(n6748) );
  INV_X1 U8029 ( .A(n7158), .ZN(n6744) );
  INV_X1 U8030 ( .A(n7157), .ZN(n6742) );
  NAND2_X1 U8031 ( .A1(n8487), .A2(n8489), .ZN(n7300) );
  INV_X1 U8032 ( .A(n11893), .ZN(n7177) );
  NOR2_X1 U8033 ( .A1(n11893), .A2(n11896), .ZN(n7178) );
  NAND2_X1 U8034 ( .A1(n11937), .A2(n11940), .ZN(n6760) );
  NOR2_X1 U8035 ( .A1(n11956), .A2(n11953), .ZN(n7153) );
  NAND2_X1 U8036 ( .A1(n11956), .A2(n11953), .ZN(n7152) );
  INV_X1 U8037 ( .A(n11921), .ZN(n7165) );
  NOR2_X1 U8038 ( .A1(n11924), .A2(n11921), .ZN(n7166) );
  NOR2_X1 U8039 ( .A1(n7153), .A2(n6758), .ZN(n6757) );
  INV_X1 U8040 ( .A(n6760), .ZN(n6758) );
  INV_X1 U8041 ( .A(n7152), .ZN(n6755) );
  AND2_X1 U8042 ( .A1(n11939), .A2(n6762), .ZN(n6761) );
  INV_X1 U8043 ( .A(n11937), .ZN(n6762) );
  NAND2_X1 U8044 ( .A1(n11742), .A2(n11741), .ZN(n11780) );
  NAND2_X1 U8045 ( .A1(n13235), .A2(n12004), .ZN(n11742) );
  INV_X1 U8046 ( .A(n10456), .ZN(n10275) );
  NAND2_X1 U8047 ( .A1(n8574), .A2(n7295), .ZN(n7294) );
  AND2_X1 U8048 ( .A1(n8584), .A2(SI_26_), .ZN(n7220) );
  AOI21_X1 U8049 ( .B1(n7054), .B2(n7056), .A(n7052), .ZN(n7051) );
  INV_X1 U8050 ( .A(n7795), .ZN(n7052) );
  NAND2_X1 U8051 ( .A1(n11983), .A2(n11986), .ZN(n7133) );
  NOR2_X1 U8052 ( .A1(n11983), .A2(n11986), .ZN(n7134) );
  AND2_X1 U8053 ( .A1(n6595), .A2(n11755), .ZN(n7194) );
  NAND2_X1 U8054 ( .A1(n13820), .A2(n6522), .ZN(n6824) );
  AOI21_X1 U8055 ( .B1(n8585), .B2(n7220), .A(n7219), .ZN(n7218) );
  INV_X1 U8056 ( .A(n8605), .ZN(n7219) );
  AOI21_X1 U8057 ( .B1(n8585), .B2(n8584), .A(SI_26_), .ZN(n7221) );
  INV_X1 U8058 ( .A(n8584), .ZN(n7217) );
  NAND2_X1 U8059 ( .A1(n7218), .A2(n7215), .ZN(n7214) );
  INV_X1 U8060 ( .A(n7220), .ZN(n7215) );
  NAND2_X1 U8061 ( .A1(n8441), .A2(n9982), .ZN(n8465) );
  NAND2_X1 U8062 ( .A1(n7202), .A2(n7203), .ZN(n8439) );
  AOI21_X1 U8063 ( .B1(n7205), .B2(n6479), .A(n6599), .ZN(n7203) );
  INV_X1 U8064 ( .A(n8109), .ZN(n7193) );
  OAI21_X1 U8065 ( .B1(n14164), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n6502), .ZN(
        n7069) );
  INV_X1 U8066 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n14149) );
  AND2_X1 U8067 ( .A1(n7018), .A2(n10162), .ZN(n7017) );
  NAND2_X1 U8068 ( .A1(n7019), .A2(n10160), .ZN(n7018) );
  AND3_X1 U8069 ( .A1(n10785), .A2(n10783), .A3(n6636), .ZN(n7021) );
  AND2_X1 U8070 ( .A1(n10486), .A2(n10487), .ZN(n6636) );
  INV_X1 U8071 ( .A(n8928), .ZN(n8929) );
  OAI21_X1 U8072 ( .B1(n8926), .B2(n12368), .A(n8927), .ZN(n8928) );
  INV_X1 U8073 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n11082) );
  INV_X1 U8074 ( .A(n8892), .ZN(n6921) );
  OR2_X1 U8075 ( .A1(n7772), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n7786) );
  NAND2_X1 U8076 ( .A1(n7929), .A2(n12646), .ZN(n8885) );
  NOR2_X1 U8077 ( .A1(n7578), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n6617) );
  INV_X1 U8078 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n7493) );
  AND2_X1 U8079 ( .A1(n8793), .A2(n10145), .ZN(n6908) );
  INV_X1 U8080 ( .A(n8801), .ZN(n6910) );
  NOR2_X1 U8081 ( .A1(n12694), .A2(n6947), .ZN(n6946) );
  INV_X1 U8082 ( .A(n7846), .ZN(n7067) );
  NOR2_X1 U8083 ( .A1(P3_IR_REG_25__SCAN_IN), .A2(P3_IR_REG_26__SCAN_IN), .ZN(
        n7289) );
  NAND2_X1 U8084 ( .A1(n7022), .A2(n6535), .ZN(n7718) );
  AOI21_X1 U8085 ( .B1(n7550), .B2(n7504), .A(n6565), .ZN(n7063) );
  INV_X1 U8086 ( .A(n7504), .ZN(n7061) );
  OR2_X1 U8087 ( .A1(n7554), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n7536) );
  NOR2_X1 U8088 ( .A1(n12958), .A2(n12927), .ZN(n7271) );
  NOR2_X1 U8089 ( .A1(n7255), .A2(n7253), .ZN(n7252) );
  INV_X1 U8090 ( .A(n9663), .ZN(n7253) );
  INV_X1 U8091 ( .A(n7343), .ZN(n7232) );
  AND2_X1 U8092 ( .A1(n12976), .A2(n12986), .ZN(n7235) );
  NAND2_X1 U8093 ( .A1(n12976), .A2(n7234), .ZN(n7233) );
  INV_X1 U8094 ( .A(n12921), .ZN(n7234) );
  INV_X1 U8095 ( .A(n7132), .ZN(n7131) );
  AOI21_X1 U8096 ( .B1(n13285), .B2(n6496), .A(n13221), .ZN(n7132) );
  INV_X1 U8097 ( .A(n11353), .ZN(n11351) );
  INV_X1 U8098 ( .A(n10127), .ZN(n10125) );
  OR2_X1 U8099 ( .A1(n10085), .A2(n14585), .ZN(n10127) );
  INV_X1 U8100 ( .A(n6809), .ZN(n6803) );
  INV_X1 U8101 ( .A(n13252), .ZN(n13266) );
  OAI21_X1 U8102 ( .B1(n13327), .B2(n13214), .A(n13213), .ZN(n13314) );
  INV_X1 U8103 ( .A(n9044), .ZN(n9065) );
  INV_X1 U8104 ( .A(n12254), .ZN(n6898) );
  INV_X1 U8105 ( .A(n9810), .ZN(n12259) );
  NAND2_X1 U8106 ( .A1(n8610), .A2(n7298), .ZN(n7297) );
  INV_X1 U8107 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n7992) );
  NAND2_X1 U8108 ( .A1(n13741), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6685) );
  NOR2_X1 U8109 ( .A1(n14009), .A2(n6828), .ZN(n6827) );
  INV_X1 U8110 ( .A(n6829), .ZN(n6828) );
  NAND2_X1 U8111 ( .A1(n13807), .A2(n13788), .ZN(n6885) );
  NOR2_X1 U8112 ( .A1(n13859), .A2(n13581), .ZN(n6872) );
  INV_X1 U8113 ( .A(n12092), .ZN(n6871) );
  INV_X1 U8114 ( .A(n14114), .ZN(n8688) );
  INV_X1 U8115 ( .A(n12083), .ZN(n6858) );
  AND2_X1 U8116 ( .A1(n11463), .A2(n12078), .ZN(n6857) );
  INV_X1 U8117 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n8251) );
  NOR2_X1 U8118 ( .A1(n10284), .A2(n6852), .ZN(n6850) );
  NAND2_X1 U8119 ( .A1(n13838), .A2(n6827), .ZN(n12142) );
  NAND2_X1 U8120 ( .A1(n13873), .A2(n13872), .ZN(n13871) );
  NAND2_X1 U8121 ( .A1(n6861), .A2(n6859), .ZN(n13918) );
  AOI21_X1 U8122 ( .B1(n6860), .B2(n6862), .A(n6526), .ZN(n6859) );
  NAND2_X1 U8123 ( .A1(n10571), .A2(n10934), .ZN(n10952) );
  INV_X1 U8124 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n7995) );
  INV_X1 U8125 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8042) );
  NOR2_X1 U8126 ( .A1(n8497), .A2(n8480), .ZN(n7189) );
  XNOR2_X1 U8127 ( .A(n8722), .B(n8721), .ZN(n9821) );
  INV_X1 U8128 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8721) );
  NOR2_X1 U8129 ( .A1(n8038), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n8413) );
  INV_X1 U8130 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n8307) );
  AOI21_X1 U8131 ( .B1(n6723), .B2(n6725), .A(n6562), .ZN(n6718) );
  INV_X1 U8132 ( .A(n6723), .ZN(n6719) );
  INV_X1 U8133 ( .A(n8295), .ZN(n6725) );
  OAI21_X1 U8134 ( .B1(n8258), .B2(n7201), .A(n8280), .ZN(n7200) );
  NOR2_X1 U8135 ( .A1(n8211), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n8238) );
  OR2_X1 U8136 ( .A1(n8207), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n8211) );
  AOI21_X1 U8137 ( .B1(n8189), .B2(n7197), .A(n7196), .ZN(n7195) );
  INV_X1 U8138 ( .A(n8204), .ZN(n7196) );
  INV_X1 U8139 ( .A(n8185), .ZN(n7197) );
  NOR2_X1 U8140 ( .A1(n8156), .A2(n8188), .ZN(n6816) );
  OR2_X1 U8141 ( .A1(n8192), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n8207) );
  NAND2_X2 U8142 ( .A1(n7186), .A2(n7187), .ZN(n8111) );
  INV_X1 U8143 ( .A(n7070), .ZN(n14142) );
  INV_X1 U8144 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n14141) );
  INV_X1 U8145 ( .A(n7069), .ZN(n14146) );
  XNOR2_X1 U8146 ( .A(n7069), .B(P3_ADDR_REG_5__SCAN_IN), .ZN(n14181) );
  OAI22_X1 U8147 ( .A1(n14186), .A2(n14147), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n14185), .ZN(n14148) );
  AND2_X1 U8148 ( .A1(n14185), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n14147) );
  INV_X1 U8149 ( .A(n6700), .ZN(n14196) );
  OAI21_X1 U8150 ( .B1(n14163), .B2(n14162), .A(n6701), .ZN(n6700) );
  NAND2_X1 U8151 ( .A1(n14149), .A2(P1_ADDR_REG_8__SCAN_IN), .ZN(n6701) );
  AND2_X1 U8152 ( .A1(n6711), .A2(n6574), .ZN(n14160) );
  OR2_X1 U8153 ( .A1(n14161), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n6711) );
  AOI21_X1 U8154 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n14219), .A(n14218), .ZN(
        n14223) );
  NOR2_X1 U8155 ( .A1(n14217), .A2(n14216), .ZN(n14218) );
  INV_X1 U8156 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7077) );
  AOI21_X1 U8157 ( .B1(n7010), .B2(n11696), .A(n11695), .ZN(n7009) );
  INV_X1 U8158 ( .A(n7011), .ZN(n7010) );
  NAND2_X1 U8159 ( .A1(n6613), .A2(n15133), .ZN(n7545) );
  INV_X1 U8160 ( .A(n7543), .ZN(n6613) );
  AND3_X1 U8161 ( .A1(n7540), .A2(n7539), .A3(n7538), .ZN(n10790) );
  OR2_X1 U8162 ( .A1(n7739), .A2(n9015), .ZN(n7540) );
  NAND2_X1 U8163 ( .A1(n6617), .A2(n11082), .ZN(n7619) );
  OR2_X1 U8164 ( .A1(n10161), .A2(n10160), .ZN(n7020) );
  INV_X1 U8165 ( .A(n11064), .ZN(n6988) );
  INV_X1 U8166 ( .A(n6618), .ZN(n7725) );
  INV_X1 U8167 ( .A(n12361), .ZN(n12338) );
  NOR2_X1 U8168 ( .A1(n8932), .A2(n8762), .ZN(n8920) );
  NAND2_X1 U8169 ( .A1(n14805), .A2(n10871), .ZN(n14824) );
  NAND2_X1 U8170 ( .A1(n14841), .A2(n10873), .ZN(n14860) );
  NOR2_X1 U8171 ( .A1(n10861), .A2(n14865), .ZN(n14900) );
  INV_X1 U8172 ( .A(n6905), .ZN(n10860) );
  NAND2_X1 U8173 ( .A1(n14880), .A2(n10875), .ZN(n14887) );
  NAND2_X1 U8174 ( .A1(n11078), .A2(n11079), .ZN(n11080) );
  OR2_X1 U8175 ( .A1(n12388), .A2(n14299), .ZN(n6933) );
  NAND2_X1 U8176 ( .A1(n12409), .A2(n6929), .ZN(n6928) );
  INV_X1 U8177 ( .A(n12422), .ZN(n6929) );
  OR2_X1 U8178 ( .A1(n12388), .A2(n6931), .ZN(n6930) );
  OR2_X1 U8179 ( .A1(n12422), .A2(n14299), .ZN(n6931) );
  NAND2_X1 U8180 ( .A1(n12411), .A2(n12412), .ZN(n12416) );
  NAND2_X1 U8181 ( .A1(n12416), .A2(n12420), .ZN(n12438) );
  NAND2_X1 U8182 ( .A1(n12438), .A2(n12441), .ZN(n12462) );
  AND3_X1 U8183 ( .A1(n6930), .A2(n6928), .A3(n12440), .ZN(n12456) );
  INV_X1 U8184 ( .A(n6927), .ZN(n6926) );
  AOI22_X1 U8185 ( .A1(n6927), .A2(n12488), .B1(n12460), .B2(n6610), .ZN(n6925) );
  NAND2_X1 U8186 ( .A1(n6924), .A2(n6927), .ZN(n12520) );
  NAND2_X1 U8187 ( .A1(n12461), .A2(n12459), .ZN(n6924) );
  NOR2_X1 U8188 ( .A1(n12563), .A2(n12575), .ZN(n12566) );
  AND2_X1 U8189 ( .A1(n8910), .A2(n7937), .ZN(n12575) );
  NAND2_X1 U8190 ( .A1(n7819), .A2(n7818), .ZN(n7836) );
  NAND2_X1 U8191 ( .A1(n12623), .A2(n8892), .ZN(n12610) );
  INV_X1 U8192 ( .A(n7794), .ZN(n7274) );
  NAND2_X1 U8193 ( .A1(n12643), .A2(n7794), .ZN(n12630) );
  NAND2_X1 U8194 ( .A1(n12640), .A2(n8891), .ZN(n12625) );
  NAND2_X1 U8195 ( .A1(n6570), .A2(n6944), .ZN(n6943) );
  NAND2_X1 U8196 ( .A1(n12645), .A2(n12644), .ZN(n12643) );
  AND2_X1 U8197 ( .A1(n8885), .A2(n8886), .ZN(n12666) );
  NAND2_X1 U8198 ( .A1(n6618), .A2(n7724), .ZN(n7742) );
  AND2_X1 U8199 ( .A1(n7763), .A2(n7762), .ZN(n12690) );
  AND2_X1 U8200 ( .A1(n12716), .A2(n7711), .ZN(n12702) );
  INV_X1 U8201 ( .A(n7652), .ZN(n7651) );
  OR2_X1 U8202 ( .A1(n7670), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n7687) );
  AND2_X1 U8203 ( .A1(n8862), .A2(n8861), .ZN(n11483) );
  INV_X1 U8204 ( .A(n6939), .ZN(n6938) );
  OAI21_X1 U8205 ( .B1(n6942), .B2(n6940), .A(n8845), .ZN(n6939) );
  NAND2_X1 U8206 ( .A1(n6941), .A2(n8840), .ZN(n6940) );
  NAND2_X1 U8207 ( .A1(n7586), .A2(n7585), .ZN(n10996) );
  OR2_X1 U8208 ( .A1(n7514), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7578) );
  INV_X1 U8209 ( .A(n6617), .ZN(n7598) );
  NAND2_X1 U8210 ( .A1(n6471), .A2(n7565), .ZN(n10739) );
  OR2_X1 U8211 ( .A1(n7567), .A2(n7566), .ZN(n7568) );
  OAI21_X1 U8212 ( .B1(n10523), .B2(n10522), .A(n7563), .ZN(n7569) );
  INV_X1 U8213 ( .A(n7562), .ZN(n10802) );
  AND4_X1 U8214 ( .A1(n7533), .A2(n7532), .A3(n7531), .A4(n7530), .ZN(n10804)
         );
  INV_X1 U8215 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n7458) );
  NAND2_X1 U8216 ( .A1(n6615), .A2(n6614), .ZN(n7543) );
  INV_X1 U8217 ( .A(n7482), .ZN(n6615) );
  AND2_X1 U8218 ( .A1(n8810), .A2(n8808), .ZN(n10214) );
  NAND2_X1 U8219 ( .A1(n7283), .A2(n7457), .ZN(n10212) );
  NAND2_X1 U8220 ( .A1(n6907), .A2(n6909), .ZN(n10514) );
  AOI21_X1 U8221 ( .B1(n10145), .B2(n6911), .A(n6910), .ZN(n6909) );
  NAND2_X1 U8222 ( .A1(n8788), .A2(n6908), .ZN(n6907) );
  INV_X1 U8223 ( .A(n8796), .ZN(n6911) );
  INV_X1 U8224 ( .A(n7912), .ZN(n10230) );
  NAND2_X1 U8225 ( .A1(n10142), .A2(n7437), .ZN(n10231) );
  NAND2_X1 U8226 ( .A1(n8793), .A2(n8788), .ZN(n14911) );
  INV_X1 U8227 ( .A(n12804), .ZN(n14925) );
  OR2_X1 U8228 ( .A1(n8759), .A2(n9050), .ZN(n7406) );
  NOR2_X1 U8229 ( .A1(n11630), .A2(n12554), .ZN(n12814) );
  NOR2_X1 U8230 ( .A1(n14919), .A2(n12555), .ZN(n7908) );
  NAND2_X1 U8231 ( .A1(n7849), .A2(n7848), .ZN(n11677) );
  NAND2_X1 U8232 ( .A1(n6948), .A2(n6946), .ZN(n12660) );
  NAND2_X1 U8233 ( .A1(n6948), .A2(n8876), .ZN(n12695) );
  NAND2_X1 U8234 ( .A1(n7924), .A2(n6942), .ZN(n6937) );
  NAND2_X1 U8235 ( .A1(n9089), .A2(n7956), .ZN(n6992) );
  NAND2_X1 U8236 ( .A1(n7878), .A2(n7877), .ZN(n8747) );
  XNOR2_X1 U8237 ( .A(n7973), .B(n7972), .ZN(n9527) );
  INV_X1 U8238 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n7972) );
  INV_X1 U8239 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n7889) );
  AND2_X1 U8240 ( .A1(n7733), .A2(n7717), .ZN(n7731) );
  NAND2_X1 U8241 ( .A1(n7030), .A2(n7028), .ZN(n7714) );
  AOI21_X1 U8242 ( .B1(n7031), .B2(n7033), .A(n7029), .ZN(n7028) );
  INV_X1 U8243 ( .A(n7699), .ZN(n7029) );
  OR2_X1 U8244 ( .A1(n7666), .A2(P3_IR_REG_15__SCAN_IN), .ZN(n7680) );
  AND2_X1 U8245 ( .A1(n7677), .A2(n7662), .ZN(n7663) );
  INV_X1 U8246 ( .A(n7641), .ZN(n7642) );
  INV_X1 U8247 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n7645) );
  NAND2_X1 U8248 ( .A1(n7037), .A2(n7034), .ZN(n7592) );
  AOI21_X1 U8249 ( .B1(n7036), .B2(n7040), .A(n7035), .ZN(n7034) );
  NOR2_X1 U8250 ( .A1(n15130), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n7035) );
  OR2_X1 U8251 ( .A1(n7592), .A2(n7591), .ZN(n7608) );
  OAI22_X1 U8252 ( .A1(n7502), .A2(n7501), .B1(P1_DATAO_REG_6__SCAN_IN), .B2(
        n6819), .ZN(n7551) );
  OR2_X1 U8253 ( .A1(n7508), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n7554) );
  XNOR2_X1 U8254 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n7500) );
  NAND2_X1 U8255 ( .A1(n7445), .A2(n7444), .ZN(n7449) );
  NAND2_X1 U8256 ( .A1(n7428), .A2(n6984), .ZN(n7472) );
  NAND2_X1 U8257 ( .A1(n7390), .A2(n7389), .ZN(n7426) );
  XNOR2_X1 U8258 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n7404) );
  NAND2_X1 U8259 ( .A1(n7387), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7417) );
  INV_X1 U8260 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n7387) );
  OR2_X1 U8261 ( .A1(n13021), .A2(n7258), .ZN(n7257) );
  INV_X1 U8262 ( .A(n9845), .ZN(n7258) );
  INV_X1 U8263 ( .A(n6624), .ZN(n11128) );
  OAI21_X1 U8264 ( .B1(n11122), .B2(n11123), .A(n6558), .ZN(n6624) );
  INV_X1 U8265 ( .A(n7271), .ZN(n7266) );
  NAND2_X1 U8266 ( .A1(n11499), .A2(n11498), .ZN(n11500) );
  NAND2_X1 U8267 ( .A1(n11496), .A2(n11495), .ZN(n11501) );
  NAND2_X1 U8268 ( .A1(n11589), .A2(n11588), .ZN(n11590) );
  NOR2_X1 U8269 ( .A1(n10660), .A2(n7247), .ZN(n7246) );
  INV_X1 U8270 ( .A(n10657), .ZN(n7247) );
  AOI21_X1 U8271 ( .B1(n6469), .B2(n7238), .A(n6557), .ZN(n7237) );
  XNOR2_X1 U8272 ( .A(n9858), .B(n11806), .ZN(n9405) );
  NAND2_X1 U8273 ( .A1(n11590), .A2(n11591), .ZN(n12890) );
  NAND2_X1 U8274 ( .A1(n11131), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n11290) );
  AND2_X1 U8275 ( .A1(n12072), .A2(n12056), .ZN(n9373) );
  AND2_X1 U8276 ( .A1(n9576), .A2(n10171), .ZN(n9359) );
  AND2_X1 U8277 ( .A1(n13125), .A2(n13124), .ZN(n13126) );
  XNOR2_X1 U8278 ( .A(n6813), .B(n13197), .ZN(n13226) );
  NAND2_X1 U8279 ( .A1(n6811), .A2(n6810), .ZN(n6813) );
  AOI21_X1 U8280 ( .B1(n6812), .B2(n7127), .A(n6568), .ZN(n6810) );
  INV_X1 U8281 ( .A(n13403), .ZN(n13235) );
  NAND2_X1 U8282 ( .A1(n13413), .A2(n6540), .ZN(n13248) );
  AND2_X1 U8283 ( .A1(n11757), .A2(n11756), .ZN(n13268) );
  AOI21_X1 U8284 ( .B1(n13290), .B2(n6498), .A(n7131), .ZN(n13260) );
  NAND2_X1 U8285 ( .A1(n6783), .A2(n6785), .ZN(n13327) );
  AOI21_X1 U8286 ( .B1(n13347), .B2(n6786), .A(n6545), .ZN(n6785) );
  NAND2_X1 U8287 ( .A1(n13207), .A2(n6784), .ZN(n6783) );
  INV_X1 U8288 ( .A(n6791), .ZN(n6786) );
  NAND2_X1 U8289 ( .A1(n6717), .A2(n6463), .ZN(n13350) );
  NAND2_X1 U8290 ( .A1(n6768), .A2(n6767), .ZN(n13179) );
  AND2_X1 U8291 ( .A1(n7339), .A2(n13176), .ZN(n6767) );
  OAI21_X1 U8292 ( .B1(n13201), .B2(n13200), .A(n7169), .ZN(n13389) );
  OR2_X1 U8293 ( .A1(n13466), .A2(n13199), .ZN(n7169) );
  NOR2_X2 U8294 ( .A1(n11442), .A2(n13472), .ZN(n11564) );
  OR2_X1 U8295 ( .A1(n11345), .A2(n6797), .ZN(n6796) );
  INV_X1 U8296 ( .A(n11284), .ZN(n6797) );
  NOR2_X2 U8297 ( .A1(n10706), .A2(n14710), .ZN(n10705) );
  INV_X1 U8298 ( .A(n12025), .ZN(n6815) );
  NAND2_X1 U8299 ( .A1(n9376), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7227) );
  NAND2_X1 U8300 ( .A1(n12026), .A2(n10329), .ZN(n10328) );
  INV_X1 U8301 ( .A(n13196), .ZN(n7121) );
  INV_X1 U8302 ( .A(n13265), .ZN(n13416) );
  NAND2_X1 U8303 ( .A1(n10258), .A2(n10257), .ZN(n10704) );
  CLKBUF_X1 U8304 ( .A(n9560), .Z(n14693) );
  INV_X1 U8305 ( .A(n9399), .ZN(n11814) );
  INV_X1 U8306 ( .A(n11806), .ZN(n14667) );
  INV_X1 U8307 ( .A(n6770), .ZN(n6769) );
  OAI21_X1 U8308 ( .B1(P2_IR_REG_31__SCAN_IN), .B2(n6773), .A(n6772), .ZN(
        n6770) );
  NAND2_X1 U8309 ( .A1(n6800), .A2(n8978), .ZN(n7222) );
  INV_X1 U8310 ( .A(n9328), .ZN(n6800) );
  XNOR2_X1 U8311 ( .A(n8991), .B(n8990), .ZN(n11219) );
  INV_X1 U8312 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8990) );
  OR2_X1 U8313 ( .A1(n9062), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n9068) );
  OR2_X1 U8314 ( .A1(n9068), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n9070) );
  OR2_X1 U8315 ( .A1(n9024), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n9044) );
  INV_X1 U8316 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8966) );
  CLKBUF_X1 U8317 ( .A(n9018), .Z(n9019) );
  AND2_X1 U8318 ( .A1(n8386), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8417) );
  INV_X1 U8319 ( .A(n10605), .ZN(n6890) );
  OR2_X1 U8320 ( .A1(n11198), .A2(n11197), .ZN(n6681) );
  OR2_X1 U8321 ( .A1(n9695), .A2(n9810), .ZN(n9420) );
  NAND2_X1 U8322 ( .A1(n6668), .A2(n6666), .ZN(n13604) );
  AOI21_X1 U8323 ( .B1(n6669), .B2(n6671), .A(n6667), .ZN(n6666) );
  INV_X1 U8324 ( .A(n13606), .ZN(n6667) );
  NOR2_X1 U8325 ( .A1(n8252), .A2(n8251), .ZN(n8274) );
  NAND2_X1 U8326 ( .A1(n13574), .A2(n12246), .ZN(n6899) );
  NOR2_X1 U8327 ( .A1(n9820), .A2(n10305), .ZN(n9826) );
  INV_X1 U8328 ( .A(n9816), .ZN(n10307) );
  OR2_X1 U8329 ( .A1(n8322), .A2(n8314), .ZN(n8368) );
  INV_X1 U8330 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n8367) );
  NOR2_X1 U8331 ( .A1(n8368), .A2(n8367), .ZN(n8386) );
  INV_X1 U8332 ( .A(n9814), .ZN(n9280) );
  XNOR2_X1 U8333 ( .A(n6820), .B(n13878), .ZN(n8712) );
  NOR2_X1 U8334 ( .A1(n12140), .A2(n6822), .ZN(n6821) );
  NOR2_X1 U8335 ( .A1(n9501), .A2(n6693), .ZN(n9494) );
  AND2_X1 U8336 ( .A1(n9506), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6693) );
  NAND2_X1 U8337 ( .A1(n9494), .A2(n9493), .ZN(n9492) );
  NAND2_X1 U8338 ( .A1(n9740), .A2(n6683), .ZN(n9742) );
  NAND2_X1 U8339 ( .A1(n9736), .A2(n9581), .ZN(n6683) );
  NAND2_X1 U8340 ( .A1(n9742), .A2(n9743), .ZN(n9935) );
  INV_X1 U8341 ( .A(n8001), .ZN(n8038) );
  XNOR2_X1 U8342 ( .A(n10974), .B(n14447), .ZN(n14444) );
  NAND2_X1 U8343 ( .A1(n10972), .A2(n6697), .ZN(n10974) );
  OR2_X1 U8344 ( .A1(n10973), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6697) );
  AND2_X1 U8345 ( .A1(n13871), .A2(n6870), .ZN(n13847) );
  NAND2_X1 U8346 ( .A1(n13871), .A2(n12092), .ZN(n13848) );
  AOI21_X1 U8347 ( .B1(n6979), .B2(n6977), .A(n6543), .ZN(n6976) );
  INV_X1 U8348 ( .A(n6979), .ZN(n6978) );
  AOI21_X1 U8349 ( .B1(n13899), .B2(n12108), .A(n12087), .ZN(n13883) );
  NOR2_X1 U8350 ( .A1(n13925), .A2(n14051), .ZN(n13887) );
  AND2_X1 U8351 ( .A1(n8417), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8432) );
  NAND2_X1 U8352 ( .A1(n8432), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n8448) );
  AOI21_X1 U8353 ( .B1(n6964), .B2(n6966), .A(n6963), .ZN(n6962) );
  INV_X1 U8354 ( .A(n12102), .ZN(n6963) );
  NAND2_X1 U8355 ( .A1(n13960), .A2(n12125), .ZN(n13962) );
  NAND2_X1 U8356 ( .A1(n11455), .A2(n11454), .ZN(n12079) );
  NAND2_X1 U8357 ( .A1(n11465), .A2(n14124), .ZN(n13975) );
  NOR2_X1 U8358 ( .A1(n11383), .A2(n14397), .ZN(n11465) );
  AOI21_X1 U8359 ( .B1(n6508), .B2(n6843), .A(n6840), .ZN(n6839) );
  AND2_X1 U8360 ( .A1(n9276), .A2(n9416), .ZN(n12177) );
  OR2_X1 U8361 ( .A1(n8337), .A2(n8320), .ZN(n8322) );
  AND4_X1 U8362 ( .A1(n8319), .A2(n8318), .A3(n8317), .A4(n8316), .ZN(n12166)
         );
  NOR2_X1 U8363 ( .A1(n10953), .A2(n11327), .ZN(n10989) );
  OAI21_X1 U8364 ( .B1(n10950), .B2(n6855), .A(n6853), .ZN(n11101) );
  AOI21_X1 U8365 ( .B1(n10630), .B2(n6478), .A(n6544), .ZN(n6853) );
  INV_X1 U8366 ( .A(n10386), .ZN(n10573) );
  OR2_X1 U8367 ( .A1(n10479), .A2(n10596), .ZN(n10572) );
  NOR2_X1 U8368 ( .A1(n10572), .A2(n14459), .ZN(n10571) );
  INV_X1 U8369 ( .A(n6852), .ZN(n6851) );
  NAND2_X1 U8370 ( .A1(n6826), .A2(n6954), .ZN(n10479) );
  OAI21_X1 U8371 ( .B1(n10457), .B2(n10456), .A(n10280), .ZN(n14477) );
  NOR2_X1 U8372 ( .A1(n14488), .A2(n14486), .ZN(n14489) );
  NAND2_X1 U8373 ( .A1(n9280), .A2(n8741), .ZN(n13983) );
  NAND2_X1 U8374 ( .A1(n9695), .A2(n9840), .ZN(n10276) );
  OR2_X1 U8375 ( .A1(n13961), .A2(n10062), .ZN(n9827) );
  AND2_X1 U8376 ( .A1(n13777), .A2(n13776), .ZN(n13994) );
  INV_X1 U8377 ( .A(n13998), .ZN(n14004) );
  AND2_X1 U8378 ( .A1(n13798), .A2(n6515), .ZN(n14016) );
  AND2_X1 U8379 ( .A1(n13855), .A2(n10480), .ZN(n14405) );
  NAND2_X1 U8380 ( .A1(n6956), .A2(n10294), .ZN(n10473) );
  AND2_X1 U8381 ( .A1(n8071), .A2(n7334), .ZN(n8084) );
  OR2_X1 U8382 ( .A1(n9643), .A2(n8266), .ZN(n8083) );
  INV_X1 U8383 ( .A(n14405), .ZN(n14518) );
  AND2_X1 U8384 ( .A1(n9821), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8993) );
  XNOR2_X1 U8385 ( .A(n7212), .B(n8679), .ZN(n13514) );
  XNOR2_X1 U8386 ( .A(n8653), .B(n8652), .ZN(n11739) );
  OAI21_X1 U8387 ( .B1(n8586), .B2(n8585), .A(n8584), .ZN(n8606) );
  INV_X1 U8388 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n8731) );
  NAND2_X1 U8389 ( .A1(n8482), .A2(n8481), .ZN(n7190) );
  OAI21_X1 U8390 ( .B1(n8402), .B2(n7207), .A(n7205), .ZN(n8427) );
  NAND2_X1 U8391 ( .A1(n8402), .A2(n8401), .ZN(n8409) );
  NAND2_X1 U8392 ( .A1(n6730), .A2(n6728), .ZN(n8361) );
  NAND2_X1 U8393 ( .A1(n8396), .A2(n6729), .ZN(n6728) );
  CLKBUF_X1 U8394 ( .A(n8068), .Z(n8069) );
  NAND2_X1 U8395 ( .A1(n8091), .A2(n8077), .ZN(n8081) );
  NAND2_X1 U8396 ( .A1(n8081), .A2(n8080), .ZN(n8110) );
  INV_X1 U8397 ( .A(n8028), .ZN(n8027) );
  AND2_X1 U8398 ( .A1(n7306), .A2(n7307), .ZN(n8024) );
  NAND2_X1 U8399 ( .A1(n6640), .A2(n14180), .ZN(n14183) );
  INV_X1 U8400 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n14185) );
  INV_X1 U8401 ( .A(n7068), .ZN(n14184) );
  OAI21_X1 U8402 ( .B1(n14257), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n6501), .ZN(
        n7073) );
  NOR2_X1 U8403 ( .A1(n14238), .A2(n14237), .ZN(n14241) );
  AND3_X1 U8404 ( .A1(n7559), .A2(n7558), .A3(n7557), .ZN(n10447) );
  NAND2_X1 U8405 ( .A1(n6995), .A2(n6999), .ZN(n11573) );
  NAND2_X1 U8406 ( .A1(n11277), .A2(n7001), .ZN(n6995) );
  NOR2_X1 U8407 ( .A1(n10838), .A2(n10837), .ZN(n11062) );
  NAND2_X1 U8408 ( .A1(n12330), .A2(n11655), .ZN(n12298) );
  NAND2_X1 U8409 ( .A1(n7752), .A2(n7751), .ZN(n12681) );
  NAND2_X1 U8410 ( .A1(n7817), .A2(n7816), .ZN(n12311) );
  INV_X1 U8411 ( .A(n7020), .ZN(n10163) );
  AND3_X1 U8412 ( .A1(n7479), .A2(n7478), .A3(n7477), .ZN(n10166) );
  NAND2_X1 U8413 ( .A1(n7014), .A2(n11642), .ZN(n12316) );
  NAND2_X1 U8414 ( .A1(n12332), .A2(n12331), .ZN(n12330) );
  NAND2_X1 U8415 ( .A1(n7002), .A2(n7004), .ZN(n11415) );
  NAND2_X1 U8416 ( .A1(n7003), .A2(n7006), .ZN(n7002) );
  AND2_X1 U8417 ( .A1(n7793), .A2(n7792), .ZN(n12659) );
  NAND2_X1 U8418 ( .A1(n7835), .A2(n7834), .ZN(n12752) );
  AND4_X1 U8419 ( .A1(n7675), .A2(n7674), .A3(n7673), .A4(n7672), .ZN(n12732)
         );
  OR2_X1 U8420 ( .A1(n9758), .A2(n9289), .ZN(n12341) );
  NAND2_X1 U8421 ( .A1(n9287), .A2(n9526), .ZN(n12366) );
  AND2_X1 U8422 ( .A1(n9290), .A2(n10030), .ZN(n12364) );
  AOI21_X1 U8423 ( .B1(n6996), .B2(n6998), .A(n6547), .ZN(n6993) );
  AND2_X1 U8424 ( .A1(n8756), .A2(n7885), .ZN(n12568) );
  NAND2_X1 U8425 ( .A1(n7872), .A2(n7871), .ZN(n12585) );
  NAND2_X1 U8426 ( .A1(n7858), .A2(n7857), .ZN(n12600) );
  NAND2_X1 U8427 ( .A1(n7842), .A2(n7841), .ZN(n12614) );
  INV_X1 U8428 ( .A(n12362), .ZN(n12627) );
  INV_X1 U8429 ( .A(n12285), .ZN(n12647) );
  INV_X1 U8430 ( .A(n11574), .ZN(n14285) );
  INV_X1 U8431 ( .A(n10791), .ZN(n12377) );
  INV_X1 U8432 ( .A(n10485), .ZN(n12380) );
  INV_X1 U8433 ( .A(n14918), .ZN(n12383) );
  CLKBUF_X1 U8434 ( .A(n7910), .Z(n12805) );
  INV_X1 U8435 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n14758) );
  INV_X1 U8436 ( .A(n14871), .ZN(n14895) );
  INV_X1 U8437 ( .A(n6914), .ZN(n10854) );
  NOR2_X1 U8438 ( .A1(n10859), .A2(n14829), .ZN(n14849) );
  INV_X1 U8439 ( .A(n6912), .ZN(n10858) );
  NOR2_X1 U8440 ( .A1(n14849), .A2(n14848), .ZN(n14847) );
  OAI21_X1 U8441 ( .B1(n10865), .B2(n6935), .A(n6934), .ZN(n12386) );
  NAND2_X1 U8442 ( .A1(n6936), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n6935) );
  NAND2_X1 U8443 ( .A1(n6930), .A2(n6928), .ZN(n12435) );
  XNOR2_X1 U8444 ( .A(n12462), .B(n12469), .ZN(n12439) );
  NOR2_X1 U8445 ( .A1(n12461), .A2(n12460), .ZN(n12489) );
  AOI21_X1 U8446 ( .B1(n12506), .B2(P3_REG1_REG_17__SCAN_IN), .A(n6649), .ZN(
        n12539) );
  INV_X1 U8447 ( .A(n6654), .ZN(n6649) );
  MUX2_X1 U8448 ( .A(n9532), .B(n12385), .S(n9531), .Z(n14876) );
  AND2_X1 U8449 ( .A1(n6651), .A2(n6650), .ZN(n12545) );
  INV_X1 U8450 ( .A(n12540), .ZN(n6652) );
  NAND2_X1 U8451 ( .A1(n7282), .A2(n7747), .ZN(n12675) );
  NAND2_X1 U8452 ( .A1(n7927), .A2(n8865), .ZN(n12707) );
  NAND2_X1 U8453 ( .A1(n7695), .A2(n7694), .ZN(n12718) );
  AND2_X1 U8454 ( .A1(n7669), .A2(n7668), .ZN(n11608) );
  AND2_X1 U8455 ( .A1(n7279), .A2(n7625), .ZN(n11252) );
  INV_X1 U8456 ( .A(n14322), .ZN(n14295) );
  NAND2_X1 U8457 ( .A1(n7924), .A2(n8835), .ZN(n11000) );
  AND3_X1 U8458 ( .A1(n7526), .A2(n7525), .A3(n7524), .ZN(n10811) );
  AND3_X1 U8459 ( .A1(n7455), .A2(n7454), .A3(n7453), .ZN(n14958) );
  NAND2_X1 U8460 ( .A1(n14914), .A2(n7435), .ZN(n10144) );
  INV_X1 U8461 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n10149) );
  INV_X1 U8462 ( .A(n11002), .ZN(n14310) );
  INV_X1 U8463 ( .A(n14936), .ZN(n14929) );
  NAND2_X1 U8464 ( .A1(n14292), .A2(n10037), .ZN(n14942) );
  AND2_X1 U8465 ( .A1(n14942), .A2(n14926), .ZN(n14939) );
  INV_X1 U8466 ( .A(n14938), .ZN(n14292) );
  NAND2_X1 U8467 ( .A1(n14310), .A2(n14957), .ZN(n14294) );
  NAND2_X1 U8468 ( .A1(n8750), .A2(n7320), .ZN(n12813) );
  INV_X1 U8469 ( .A(n11677), .ZN(n12828) );
  NAND2_X1 U8470 ( .A1(n7723), .A2(n7722), .ZN(n12853) );
  INV_X1 U8471 ( .A(n12345), .ZN(n12856) );
  INV_X1 U8472 ( .A(n12314), .ZN(n12860) );
  AND2_X1 U8473 ( .A1(n7649), .A2(n7648), .ZN(n12865) );
  AND2_X1 U8474 ( .A1(n6992), .A2(n7957), .ZN(n12868) );
  INV_X1 U8475 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n12869) );
  CLKBUF_X1 U8476 ( .A(n7364), .Z(n12873) );
  XNOR2_X1 U8477 ( .A(n7874), .B(n7863), .ZN(n12878) );
  INV_X1 U8478 ( .A(SI_27_), .ZN(n12884) );
  MUX2_X1 U8479 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7379), .S(
        P3_IR_REG_27__SCAN_IN), .Z(n7381) );
  NAND2_X1 U8480 ( .A1(n6642), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7946) );
  NAND2_X1 U8481 ( .A1(n6918), .A2(n7022), .ZN(n6642) );
  NAND2_X1 U8482 ( .A1(n7813), .A2(n7801), .ZN(n7812) );
  INV_X1 U8483 ( .A(SI_23_), .ZN(n10945) );
  OAI21_X1 U8484 ( .B1(n7768), .B2(n7056), .A(n7054), .ZN(n7796) );
  NAND2_X1 U8485 ( .A1(n7053), .A2(n7769), .ZN(n7783) );
  NAND2_X1 U8486 ( .A1(n7059), .A2(n7748), .ZN(n7737) );
  INV_X1 U8487 ( .A(SI_19_), .ZN(n9982) );
  INV_X1 U8488 ( .A(SI_16_), .ZN(n9797) );
  NAND2_X1 U8489 ( .A1(n7628), .A2(n7627), .ZN(n7640) );
  INV_X1 U8490 ( .A(SI_13_), .ZN(n9196) );
  INV_X1 U8491 ( .A(SI_12_), .ZN(n9083) );
  INV_X1 U8492 ( .A(SI_11_), .ZN(n9076) );
  OAI21_X1 U8493 ( .B1(n7505), .B2(n7043), .A(n7040), .ZN(n7589) );
  XNOR2_X1 U8494 ( .A(n7510), .B(n7509), .ZN(n10920) );
  NAND2_X1 U8495 ( .A1(n7045), .A2(n7044), .ZN(n7572) );
  NAND2_X1 U8496 ( .A1(n7058), .A2(n7393), .ZN(n7443) );
  OR3_X1 U8497 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n7395) );
  NAND2_X1 U8498 ( .A1(n7429), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7431) );
  NAND2_X1 U8499 ( .A1(n7254), .A2(n9854), .ZN(n9961) );
  NAND2_X1 U8500 ( .A1(n9846), .A2(n7256), .ZN(n7254) );
  INV_X1 U8501 ( .A(n7257), .ZN(n7256) );
  NAND2_X1 U8502 ( .A1(n13031), .A2(n12928), .ZN(n12959) );
  NAND2_X1 U8503 ( .A1(n9380), .A2(n6494), .ZN(n9381) );
  INV_X1 U8504 ( .A(n9379), .ZN(n9380) );
  NAND2_X1 U8505 ( .A1(n7240), .A2(n7242), .ZN(n12971) );
  NAND2_X1 U8506 ( .A1(n7241), .A2(n12996), .ZN(n7240) );
  NAND2_X1 U8507 ( .A1(n7248), .A2(n10657), .ZN(n10659) );
  NAND2_X1 U8508 ( .A1(n10646), .A2(n10645), .ZN(n11862) );
  NAND2_X1 U8509 ( .A1(n12985), .A2(n12921), .ZN(n12977) );
  NAND2_X1 U8510 ( .A1(n11501), .A2(n11500), .ZN(n11502) );
  NAND2_X1 U8511 ( .A1(n12984), .A2(n12986), .ZN(n12985) );
  AOI21_X1 U8512 ( .B1(n7223), .B2(n9640), .A(n6563), .ZN(n9683) );
  NAND2_X1 U8513 ( .A1(n10079), .A2(n10078), .ZN(n10082) );
  NAND2_X1 U8514 ( .A1(n12995), .A2(n12996), .ZN(n12994) );
  NAND2_X1 U8515 ( .A1(n6623), .A2(n12902), .ZN(n12995) );
  NAND2_X1 U8516 ( .A1(n10717), .A2(n10716), .ZN(n11122) );
  OR2_X1 U8517 ( .A1(n10353), .A2(n10352), .ZN(n6645) );
  NAND2_X1 U8518 ( .A1(n10358), .A2(n10357), .ZN(n13491) );
  CLKBUF_X1 U8519 ( .A(n9399), .Z(n11813) );
  NAND2_X1 U8520 ( .A1(n9359), .A2(n12019), .ZN(n13015) );
  NAND2_X1 U8521 ( .A1(n9846), .A2(n9845), .ZN(n13020) );
  INV_X1 U8522 ( .A(n12066), .ZN(n12067) );
  OAI21_X1 U8523 ( .B1(n12065), .B2(n12064), .A(n10176), .ZN(n12066) );
  INV_X1 U8524 ( .A(n12063), .ZN(n12072) );
  NAND2_X1 U8525 ( .A1(n9628), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n9361) );
  NAND2_X1 U8526 ( .A1(n13161), .A2(n13300), .ZN(n13398) );
  INV_X1 U8527 ( .A(n12022), .ZN(n13401) );
  NAND2_X1 U8528 ( .A1(n7143), .A2(n13244), .ZN(n13408) );
  NAND2_X1 U8529 ( .A1(n7144), .A2(n6493), .ZN(n7143) );
  NAND2_X1 U8530 ( .A1(n7124), .A2(n13194), .ZN(n13272) );
  NAND2_X1 U8531 ( .A1(n7124), .A2(n7123), .ZN(n13413) );
  AND2_X1 U8532 ( .A1(n13259), .A2(n13194), .ZN(n7123) );
  INV_X1 U8533 ( .A(n7130), .ZN(n13276) );
  AOI21_X1 U8534 ( .B1(n13290), .B2(n13295), .A(n6496), .ZN(n7130) );
  NAND2_X1 U8535 ( .A1(n6787), .A2(n6791), .ZN(n13339) );
  NAND2_X1 U8536 ( .A1(n13207), .A2(n6788), .ZN(n6787) );
  NAND2_X1 U8537 ( .A1(n13207), .A2(n13206), .ZN(n13354) );
  NAND2_X1 U8538 ( .A1(n6768), .A2(n13176), .ZN(n13379) );
  NAND2_X1 U8539 ( .A1(n11545), .A2(n11544), .ZN(n11548) );
  OAI21_X1 U8540 ( .B1(n11151), .B2(n7094), .A(n7093), .ZN(n11368) );
  NAND2_X1 U8541 ( .A1(n7095), .A2(n11305), .ZN(n11367) );
  NAND2_X1 U8542 ( .A1(n11151), .A2(n7097), .ZN(n7095) );
  INV_X1 U8543 ( .A(n7098), .ZN(n7097) );
  NAND2_X1 U8544 ( .A1(n11285), .A2(n11284), .ZN(n11346) );
  NAND2_X1 U8545 ( .A1(n7164), .A2(n11157), .ZN(n11160) );
  NAND2_X1 U8546 ( .A1(n11151), .A2(n11150), .ZN(n11307) );
  NAND2_X1 U8547 ( .A1(n10752), .A2(n7146), .ZN(n10777) );
  NAND2_X1 U8548 ( .A1(n6807), .A2(n6805), .ZN(n10542) );
  NAND2_X1 U8549 ( .A1(n6807), .A2(n6808), .ZN(n10265) );
  OAI21_X1 U8550 ( .B1(n10263), .B2(n10262), .A(n10261), .ZN(n10711) );
  NAND2_X1 U8551 ( .A1(n7102), .A2(n7106), .ZN(n10688) );
  INV_X1 U8552 ( .A(n7107), .ZN(n7106) );
  NAND2_X1 U8553 ( .A1(n7105), .A2(n9988), .ZN(n10184) );
  NAND2_X1 U8554 ( .A1(n10196), .A2(n12027), .ZN(n7105) );
  NAND2_X1 U8555 ( .A1(n14661), .A2(n9340), .ZN(n14646) );
  OR2_X1 U8556 ( .A1(n13429), .A2(n13428), .ZN(n13501) );
  INV_X1 U8557 ( .A(n14655), .ZN(n14656) );
  AND2_X1 U8558 ( .A1(n9337), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14661) );
  MUX2_X1 U8559 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9346), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n9347) );
  NAND2_X1 U8560 ( .A1(n7172), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6801) );
  NAND2_X1 U8561 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(n9884), .ZN(n6799) );
  INV_X1 U8562 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n11377) );
  NAND2_X1 U8563 ( .A1(n8983), .A2(n8982), .ZN(n11375) );
  NAND2_X1 U8564 ( .A1(n8988), .A2(n8987), .ZN(n11269) );
  INV_X1 U8565 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11637) );
  INV_X1 U8566 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n9794) );
  INV_X1 U8567 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n9888) );
  INV_X1 U8568 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n9253) );
  INV_X1 U8569 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9202) );
  INV_X1 U8570 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9079) );
  INV_X1 U8571 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10067) );
  INV_X1 U8572 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9073) );
  INV_X1 U8573 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9029) );
  INV_X1 U8574 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9049) );
  INV_X1 U8575 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9011) );
  INV_X1 U8576 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9039) );
  INV_X1 U8577 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9396) );
  NAND2_X1 U8578 ( .A1(n10606), .A2(n10605), .ZN(n11020) );
  NAND2_X1 U8579 ( .A1(n12164), .A2(n12163), .ZN(n14343) );
  AND4_X1 U8580 ( .A1(n8373), .A2(n8372), .A3(n8371), .A4(n8370), .ZN(n14340)
         );
  NAND2_X1 U8581 ( .A1(n6681), .A2(n6680), .ZN(n14382) );
  NAND2_X1 U8582 ( .A1(n6902), .A2(n10105), .ZN(n13546) );
  OR2_X1 U8583 ( .A1(n6571), .A2(n6896), .ZN(n6893) );
  NAND2_X1 U8584 ( .A1(n11020), .A2(n11019), .ZN(n11021) );
  OAI21_X1 U8585 ( .B1(n9804), .B2(n9803), .A(n9807), .ZN(n9836) );
  NOR2_X1 U8586 ( .A1(n9836), .A2(n9835), .ZN(n9834) );
  AND2_X1 U8587 ( .A1(n6673), .A2(n6674), .ZN(n13596) );
  AOI21_X1 U8588 ( .B1(n6680), .B2(n11197), .A(n6566), .ZN(n6678) );
  AND4_X1 U8589 ( .A1(n8341), .A2(n8340), .A3(n8339), .A4(n8338), .ZN(n14376)
         );
  OR2_X1 U8590 ( .A1(n13647), .A2(n13982), .ZN(n14378) );
  OR2_X1 U8591 ( .A1(n13647), .A2(n13983), .ZN(n14377) );
  OAI211_X1 U8592 ( .C1(n9084), .C2(n13696), .A(n8096), .B(n8095), .ZN(n10463)
         );
  OR2_X1 U8593 ( .A1(n8113), .A2(n9001), .ZN(n8096) );
  NAND2_X1 U8594 ( .A1(n6657), .A2(n6660), .ZN(n13621) );
  AND2_X1 U8595 ( .A1(n6661), .A2(n13622), .ZN(n6660) );
  NAND2_X1 U8596 ( .A1(n6662), .A2(n10600), .ZN(n6661) );
  OAI211_X1 U8597 ( .C1(n6663), .C2(n6662), .A(n6658), .B(n10600), .ZN(n13623)
         );
  NAND2_X1 U8598 ( .A1(n6659), .A2(n6484), .ZN(n6658) );
  INV_X1 U8599 ( .A(n6506), .ZN(n6659) );
  INV_X1 U8600 ( .A(n14384), .ZN(n14356) );
  AND2_X1 U8601 ( .A1(n9280), .A2(n9427), .ZN(n13954) );
  NAND4_X1 U8602 ( .A1(n8124), .A2(n8123), .A3(n8122), .A4(n8121), .ZN(n13676)
         );
  INV_X1 U8603 ( .A(n8691), .ZN(n13678) );
  NAND2_X1 U8604 ( .A1(n6695), .A2(n6694), .ZN(n13703) );
  OR2_X1 U8605 ( .A1(n13696), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6695) );
  NAND2_X1 U8606 ( .A1(n13696), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6694) );
  NOR2_X1 U8607 ( .A1(n9466), .A2(n6597), .ZN(n9503) );
  NOR2_X1 U8608 ( .A1(n9503), .A2(n9502), .ZN(n9501) );
  NOR2_X1 U8609 ( .A1(n9579), .A2(n6684), .ZN(n9583) );
  AND2_X1 U8610 ( .A1(n9580), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6684) );
  NAND2_X1 U8611 ( .A1(n9583), .A2(n9582), .ZN(n9740) );
  NOR2_X1 U8612 ( .A1(n10047), .A2(n6698), .ZN(n10050) );
  AND2_X1 U8613 ( .A1(n10055), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6698) );
  NAND2_X1 U8614 ( .A1(n10050), .A2(n10049), .ZN(n10972) );
  INV_X1 U8615 ( .A(n6686), .ZN(n13740) );
  NOR2_X1 U8616 ( .A1(n13775), .A2(n13961), .ZN(n13992) );
  XNOR2_X1 U8617 ( .A(n12141), .B(n12136), .ZN(n14006) );
  NAND2_X1 U8618 ( .A1(n6875), .A2(n6873), .ZN(n12141) );
  AND2_X1 U8619 ( .A1(n6874), .A2(n6880), .ZN(n6873) );
  NAND2_X1 U8620 ( .A1(n6972), .A2(n6491), .ZN(n6971) );
  NAND2_X1 U8621 ( .A1(n12098), .A2(n12097), .ZN(n12099) );
  NAND2_X1 U8622 ( .A1(n13868), .A2(n12111), .ZN(n13845) );
  INV_X1 U8623 ( .A(n6836), .ZN(n13858) );
  AND2_X1 U8624 ( .A1(n13868), .A2(n13867), .ZN(n14042) );
  NAND2_X1 U8625 ( .A1(n13915), .A2(n12107), .ZN(n13908) );
  NAND2_X1 U8626 ( .A1(n12106), .A2(n12105), .ZN(n13913) );
  OAI21_X1 U8627 ( .B1(n11455), .B2(n6864), .A(n6862), .ZN(n13932) );
  AND2_X1 U8628 ( .A1(n14494), .A2(n14490), .ZN(n13989) );
  NAND2_X1 U8629 ( .A1(n12101), .A2(n12100), .ZN(n13973) );
  AND2_X1 U8630 ( .A1(n11231), .A2(n11172), .ZN(n7340) );
  NAND2_X1 U8631 ( .A1(n6841), .A2(n11189), .ZN(n11379) );
  NAND2_X1 U8632 ( .A1(n11227), .A2(n11226), .ZN(n6841) );
  AND2_X1 U8633 ( .A1(n10948), .A2(n10629), .ZN(n7327) );
  NAND2_X1 U8634 ( .A1(n9648), .A2(n6835), .ZN(n8115) );
  AND2_X1 U8635 ( .A1(n10276), .A2(n8690), .ZN(n10444) );
  INV_X1 U8636 ( .A(n13991), .ZN(n14268) );
  NAND2_X1 U8637 ( .A1(n8243), .A2(n8242), .ZN(n11204) );
  AND2_X2 U8638 ( .A1(n10156), .A2(n9271), .ZN(n14540) );
  INV_X1 U8639 ( .A(n13773), .ZN(n14088) );
  OAI211_X1 U8640 ( .C1(n14018), .C2(n14405), .A(n14017), .B(n6626), .ZN(
        n14095) );
  NOR2_X1 U8641 ( .A1(n14016), .A2(n14015), .ZN(n14017) );
  INV_X1 U8642 ( .A(n14019), .ZN(n6626) );
  AND2_X1 U8643 ( .A1(n14014), .A2(n14522), .ZN(n14015) );
  INV_X1 U8644 ( .A(n13967), .ZN(n12125) );
  AND2_X1 U8645 ( .A1(n8346), .A2(n8345), .ZN(n11538) );
  AND2_X1 U8646 ( .A1(n8016), .A2(n6968), .ZN(n6967) );
  INV_X1 U8647 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n6968) );
  CLKBUF_X1 U8648 ( .A(n8740), .Z(n8741) );
  NAND2_X1 U8649 ( .A1(n8734), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8018) );
  INV_X1 U8650 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n11374) );
  INV_X1 U8651 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11273) );
  XNOR2_X1 U8652 ( .A(n8727), .B(P1_IR_REG_24__SCAN_IN), .ZN(n11270) );
  XNOR2_X1 U8653 ( .A(n6825), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14136) );
  MUX2_X1 U8654 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8046), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n8048) );
  INV_X1 U8655 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10063) );
  INV_X1 U8656 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n9833) );
  INV_X1 U8657 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n9725) );
  INV_X1 U8658 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n9907) );
  INV_X1 U8659 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9727) );
  INV_X1 U8660 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n15130) );
  INV_X1 U8661 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9081) );
  NAND2_X1 U8662 ( .A1(n8264), .A2(n8263), .ZN(n8281) );
  NAND2_X1 U8663 ( .A1(n8259), .A2(n8258), .ZN(n8264) );
  INV_X1 U8664 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9074) );
  INV_X1 U8665 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9043) );
  NAND2_X1 U8666 ( .A1(n8190), .A2(n8189), .ZN(n8205) );
  NAND2_X1 U8667 ( .A1(n8186), .A2(n8185), .ZN(n8190) );
  INV_X1 U8668 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9017) );
  INV_X1 U8669 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9005) );
  INV_X1 U8670 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n8995) );
  INV_X1 U8671 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9001) );
  XNOR2_X1 U8672 ( .A(n6696), .B(P1_IR_REG_2__SCAN_IN), .ZN(n13696) );
  NOR2_X1 U8673 ( .A1(n8024), .A2(n14125), .ZN(n6696) );
  NAND2_X1 U8674 ( .A1(n14176), .A2(n14177), .ZN(n15176) );
  NOR2_X1 U8675 ( .A1(n14261), .A2(n14260), .ZN(n14259) );
  NAND2_X1 U8676 ( .A1(n7088), .A2(n7087), .ZN(n14215) );
  NAND2_X1 U8677 ( .A1(n14424), .A2(n7089), .ZN(n7088) );
  INV_X1 U8678 ( .A(n7084), .ZN(n14426) );
  OAI21_X1 U8679 ( .B1(n14424), .B2(n7086), .A(n7085), .ZN(n7084) );
  INV_X1 U8680 ( .A(n7087), .ZN(n7086) );
  AND2_X1 U8681 ( .A1(n14214), .A2(n7089), .ZN(n7085) );
  INV_X1 U8682 ( .A(n7080), .ZN(n14434) );
  INV_X1 U8683 ( .A(n14438), .ZN(n7078) );
  INV_X1 U8684 ( .A(n14239), .ZN(n7082) );
  AND2_X1 U8685 ( .A1(n12867), .A2(n8994), .ZN(P3_U3897) );
  OAI21_X1 U8686 ( .B1(n6632), .B2(n8940), .A(n9525), .ZN(n6631) );
  OAI22_X1 U8687 ( .A1(n12557), .A2(n12803), .B1(n15164), .B2(n8960), .ZN(
        n8961) );
  OAI21_X1 U8688 ( .B1(n12822), .B2(n15162), .A(n7284), .ZN(P3_U3487) );
  AOI21_X1 U8689 ( .B1(n11704), .B2(n7286), .A(n7285), .ZN(n7284) );
  NOR2_X1 U8690 ( .A1(n15164), .A2(n12747), .ZN(n7285) );
  OAI22_X1 U8691 ( .A1(n12557), .A2(n12864), .B1(n14993), .B2(n7986), .ZN(
        n7987) );
  NAND2_X1 U8692 ( .A1(n6950), .A2(n6486), .ZN(n12823) );
  NAND2_X1 U8693 ( .A1(n9640), .A2(n9639), .ZN(n9720) );
  NAND2_X1 U8694 ( .A1(n7264), .A2(n13034), .ZN(n7261) );
  NAND2_X1 U8695 ( .A1(n14744), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6782) );
  NAND2_X1 U8696 ( .A1(n6781), .A2(n14746), .ZN(n6780) );
  NAND2_X1 U8697 ( .A1(n14744), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n7138) );
  NAND2_X1 U8698 ( .A1(n13498), .A2(n14746), .ZN(n7139) );
  OR2_X1 U8699 ( .A1(n14731), .A2(n11733), .ZN(n7122) );
  NAND2_X1 U8700 ( .A1(n14731), .A2(n14680), .ZN(n7118) );
  NAND2_X1 U8701 ( .A1(n7117), .A2(n14731), .ZN(n7116) );
  XNOR2_X1 U8702 ( .A(n6676), .B(n6675), .ZN(n13534) );
  INV_X1 U8703 ( .A(n6688), .ZN(n13732) );
  NAND2_X1 U8704 ( .A1(n6692), .A2(n6689), .ZN(P1_U3262) );
  NAND2_X1 U8705 ( .A1(n13770), .A2(n13878), .ZN(n6692) );
  AOI21_X1 U8706 ( .B1(n6690), .B2(n10062), .A(n13772), .ZN(n6689) );
  NOR2_X1 U8707 ( .A1(n14424), .A2(n14423), .ZN(n14422) );
  NOR2_X1 U8708 ( .A1(n14431), .A2(n14430), .ZN(n14429) );
  AND2_X1 U8709 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n6467) );
  CLKBUF_X3 U8710 ( .A(n7542), .Z(n7822) );
  AND2_X1 U8711 ( .A1(n11019), .A2(n6891), .ZN(n6468) );
  AND2_X1 U8712 ( .A1(n6516), .A2(n10261), .ZN(n6809) );
  INV_X1 U8713 ( .A(n13786), .ZN(n6884) );
  INV_X2 U8714 ( .A(n7616), .ZN(n7600) );
  INV_X1 U8715 ( .A(n13259), .ZN(n7128) );
  AND2_X1 U8716 ( .A1(n7242), .A2(n7239), .ZN(n6469) );
  INV_X1 U8717 ( .A(n9335), .ZN(n9376) );
  AND2_X1 U8718 ( .A1(n12629), .A2(n6517), .ZN(n6470) );
  NAND2_X1 U8719 ( .A1(n7562), .A2(n10800), .ZN(n6471) );
  AND2_X1 U8720 ( .A1(n11851), .A2(n6740), .ZN(n6472) );
  AND2_X1 U8721 ( .A1(n12117), .A2(n13786), .ZN(n6473) );
  OR2_X1 U8722 ( .A1(n7137), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n6474) );
  AND2_X1 U8723 ( .A1(n11413), .A2(n12374), .ZN(n6475) );
  NOR4_X1 U8724 ( .A1(n12091), .A2(n13907), .A3(n13885), .A4(n8700), .ZN(n6476) );
  AND2_X1 U8725 ( .A1(n6715), .A2(n12042), .ZN(n6477) );
  AND2_X1 U8726 ( .A1(n6854), .A2(n10629), .ZN(n6478) );
  AND2_X1 U8727 ( .A1(n6510), .A2(n7207), .ZN(n6479) );
  INV_X1 U8728 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n14125) );
  INV_X1 U8729 ( .A(n11859), .ZN(n7161) );
  INV_X1 U8730 ( .A(n11966), .ZN(n7151) );
  OR2_X1 U8731 ( .A1(n14232), .A2(n14233), .ZN(n6480) );
  INV_X1 U8732 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7359) );
  NAND2_X1 U8733 ( .A1(n7045), .A2(n7046), .ZN(n6481) );
  NAND2_X1 U8734 ( .A1(n7048), .A2(n7049), .ZN(n6482) );
  AND2_X1 U8735 ( .A1(n7865), .A2(n7864), .ZN(n12824) );
  INV_X1 U8736 ( .A(n12824), .ZN(n11704) );
  NAND2_X1 U8737 ( .A1(n8499), .A2(SI_21_), .ZN(n6483) );
  NAND2_X1 U8738 ( .A1(n10248), .A2(n10247), .ZN(n6484) );
  OR3_X1 U8739 ( .A1(n10953), .A2(n14390), .A3(n11327), .ZN(n6485) );
  OR2_X1 U8740 ( .A1(n14993), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n6486) );
  AND2_X1 U8741 ( .A1(n6922), .A2(n8891), .ZN(n6487) );
  INV_X1 U8742 ( .A(n10949), .ZN(n6854) );
  INV_X1 U8743 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7172) );
  NOR2_X1 U8744 ( .A1(n7326), .A2(n7336), .ZN(n6488) );
  NAND2_X1 U8745 ( .A1(n13645), .A2(n13644), .ZN(n13643) );
  OR3_X1 U8746 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .A3(
        n9546), .ZN(n6489) );
  INV_X1 U8747 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8090) );
  AND3_X1 U8748 ( .A1(n11795), .A2(n11794), .A3(n11793), .ZN(n6490) );
  NAND2_X1 U8749 ( .A1(n14009), .A2(n13657), .ZN(n6491) );
  INV_X1 U8750 ( .A(n8263), .ZN(n7201) );
  INV_X1 U8751 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n9326) );
  NAND2_X1 U8752 ( .A1(n10107), .A2(n10106), .ZN(n6492) );
  NAND2_X1 U8753 ( .A1(n6814), .A2(n6812), .ZN(n6493) );
  NAND2_X1 U8754 ( .A1(n11798), .A2(n9858), .ZN(n6494) );
  NOR2_X1 U8755 ( .A1(n13825), .A2(n12116), .ZN(n6495) );
  AND2_X1 U8756 ( .A1(n13304), .A2(n13218), .ZN(n6496) );
  AND2_X1 U8757 ( .A1(n11158), .A2(n11157), .ZN(n6497) );
  AND2_X1 U8758 ( .A1(n13285), .A2(n13295), .ZN(n6498) );
  AND2_X1 U8759 ( .A1(n6488), .A2(n13634), .ZN(n6499) );
  OR2_X1 U8760 ( .A1(n12957), .A2(n12956), .ZN(n6500) );
  OR2_X1 U8761 ( .A1(n14195), .A2(n14194), .ZN(n6501) );
  OR2_X1 U8762 ( .A1(n14144), .A2(n14143), .ZN(n6502) );
  AND2_X1 U8763 ( .A1(n8245), .A2(n8244), .ZN(n6503) );
  NOR2_X1 U8764 ( .A1(n8068), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n8145) );
  NAND2_X1 U8765 ( .A1(n8313), .A2(n8312), .ZN(n11174) );
  INV_X1 U8766 ( .A(n8266), .ZN(n6835) );
  OR2_X1 U8767 ( .A1(n13967), .A2(n13662), .ZN(n6504) );
  OR3_X1 U8768 ( .A1(n9200), .A2(n6474), .A3(P2_IR_REG_19__SCAN_IN), .ZN(n6505) );
  OR2_X1 U8769 ( .A1(n10241), .A2(n10240), .ZN(n6506) );
  NAND2_X1 U8770 ( .A1(n6682), .A2(n11270), .ZN(n9418) );
  NAND2_X1 U8771 ( .A1(n8286), .A2(n8285), .ZN(n14390) );
  INV_X1 U8772 ( .A(n13788), .ZN(n6878) );
  AND2_X1 U8773 ( .A1(n14710), .A2(n10264), .ZN(n6507) );
  AND2_X1 U8774 ( .A1(n11378), .A2(n6842), .ZN(n6508) );
  AND2_X1 U8775 ( .A1(n6746), .A2(n6744), .ZN(n6509) );
  OR2_X1 U8776 ( .A1(n8426), .A2(SI_17_), .ZN(n6510) );
  INV_X1 U8777 ( .A(n8118), .ZN(n8085) );
  INV_X1 U8778 ( .A(n13063), .ZN(n7112) );
  NAND2_X1 U8779 ( .A1(n11718), .A2(n11717), .ZN(n12022) );
  AND2_X1 U8780 ( .A1(n6686), .A2(n6685), .ZN(n6511) );
  AOI21_X1 U8781 ( .B1(n12279), .B2(n8761), .A(n8760), .ZN(n8926) );
  INV_X1 U8782 ( .A(n12356), .ZN(n7013) );
  NOR2_X1 U8783 ( .A1(n12938), .A2(n7343), .ZN(n12984) );
  INV_X1 U8784 ( .A(n8876), .ZN(n6947) );
  NOR4_X1 U8785 ( .A1(n12046), .A2(n12045), .A3(n12044), .A4(n12043), .ZN(
        n6512) );
  OR2_X1 U8786 ( .A1(n14690), .A2(n13060), .ZN(n6513) );
  INV_X1 U8787 ( .A(n12091), .ZN(n13872) );
  AND2_X1 U8788 ( .A1(n6975), .A2(n6973), .ZN(n6514) );
  INV_X1 U8789 ( .A(n8575), .ZN(n7295) );
  INV_X1 U8790 ( .A(n8197), .ZN(n7315) );
  INV_X1 U8791 ( .A(n8611), .ZN(n7298) );
  NAND2_X1 U8792 ( .A1(n13838), .A2(n6829), .ZN(n6515) );
  OR2_X1 U8793 ( .A1(n14710), .A2(n10264), .ZN(n6516) );
  NAND2_X1 U8794 ( .A1(n7188), .A2(n6620), .ZN(n8537) );
  OR2_X1 U8795 ( .A1(n12644), .A2(n7274), .ZN(n6517) );
  NOR2_X1 U8796 ( .A1(n13849), .A2(n6871), .ZN(n6870) );
  INV_X1 U8797 ( .A(n7044), .ZN(n7043) );
  NOR2_X1 U8798 ( .A1(n7322), .A2(n6598), .ZN(n7044) );
  AND2_X1 U8799 ( .A1(n12219), .A2(n12218), .ZN(n6518) );
  NAND2_X1 U8800 ( .A1(n8024), .A2(n8090), .ZN(n8066) );
  AND2_X1 U8801 ( .A1(n11676), .A2(n12309), .ZN(n6519) );
  INV_X1 U8802 ( .A(n13859), .ZN(n14104) );
  NAND2_X1 U8803 ( .A1(n8546), .A2(n8545), .ZN(n13859) );
  AND2_X1 U8804 ( .A1(n9924), .A2(n9926), .ZN(n6520) );
  AND2_X1 U8805 ( .A1(n11192), .A2(n11193), .ZN(n6521) );
  NOR2_X1 U8806 ( .A1(n13831), .A2(n13849), .ZN(n6522) );
  AND2_X1 U8807 ( .A1(n13476), .A2(n11431), .ZN(n6523) );
  INV_X1 U8808 ( .A(n13640), .ZN(n14099) );
  NAND2_X1 U8809 ( .A1(n8589), .A2(n8588), .ZN(n13640) );
  AND2_X1 U8810 ( .A1(n12571), .A2(n12570), .ZN(n6524) );
  OR2_X1 U8811 ( .A1(n10887), .A2(n14996), .ZN(n6525) );
  AND2_X1 U8812 ( .A1(n14063), .A2(n12084), .ZN(n6526) );
  NAND2_X1 U8813 ( .A1(n14459), .A2(n11023), .ZN(n6527) );
  AND2_X1 U8814 ( .A1(n6673), .A2(n6672), .ZN(n6528) );
  AND2_X1 U8815 ( .A1(n11546), .A2(n11544), .ZN(n6529) );
  OR2_X1 U8816 ( .A1(n14183), .A2(n14182), .ZN(n6530) );
  OAI21_X1 U8817 ( .B1(n6817), .B2(SI_6_), .A(n8185), .ZN(n8156) );
  AND2_X1 U8818 ( .A1(n12168), .A2(n12163), .ZN(n6531) );
  AND2_X1 U8819 ( .A1(n11530), .A2(n11526), .ZN(n6532) );
  AND2_X1 U8820 ( .A1(n11643), .A2(n11642), .ZN(n6533) );
  AND2_X1 U8821 ( .A1(n7480), .A2(n7457), .ZN(n6534) );
  AND2_X1 U8822 ( .A1(n7332), .A2(n7277), .ZN(n6535) );
  NOR2_X1 U8823 ( .A1(n13459), .A2(n13203), .ZN(n6536) );
  AND2_X1 U8824 ( .A1(n13491), .A2(n10754), .ZN(n6537) );
  AND2_X1 U8825 ( .A1(n8807), .A2(n10214), .ZN(n6538) );
  NAND2_X1 U8826 ( .A1(n14372), .A2(n13953), .ZN(n6539) );
  OR2_X1 U8827 ( .A1(n13416), .A2(n13195), .ZN(n6540) );
  AND2_X1 U8828 ( .A1(n8042), .A2(n6903), .ZN(n6541) );
  NAND2_X1 U8829 ( .A1(n12924), .A2(n12923), .ZN(n6542) );
  NOR2_X1 U8830 ( .A1(n14051), .A2(n13661), .ZN(n6543) );
  NOR2_X1 U8831 ( .A1(n11327), .A2(n14379), .ZN(n6544) );
  NOR2_X1 U8832 ( .A1(n13442), .A2(n13211), .ZN(n6545) );
  NOR2_X1 U8833 ( .A1(n11848), .A2(n10541), .ZN(n6546) );
  NOR2_X1 U8834 ( .A1(n11575), .A2(n11574), .ZN(n6547) );
  NOR2_X1 U8835 ( .A1(n8697), .A2(n6454), .ZN(n6548) );
  INV_X1 U8836 ( .A(n7005), .ZN(n7004) );
  NOR2_X1 U8837 ( .A1(n11275), .A2(n14287), .ZN(n7005) );
  NAND2_X1 U8838 ( .A1(n12262), .A2(n12261), .ZN(n6549) );
  INV_X1 U8839 ( .A(n6865), .ZN(n6864) );
  NOR2_X1 U8840 ( .A1(n12083), .A2(n6866), .ZN(n6865) );
  OR2_X1 U8841 ( .A1(n10065), .A2(n9375), .ZN(n6550) );
  AND2_X1 U8842 ( .A1(n7999), .A2(n7998), .ZN(n8037) );
  AND2_X1 U8843 ( .A1(n7467), .A2(n7466), .ZN(n6551) );
  AND2_X1 U8844 ( .A1(n14322), .A2(n12374), .ZN(n6552) );
  AND3_X1 U8845 ( .A1(n8138), .A2(n8136), .A3(n8135), .ZN(n6553) );
  INV_X1 U8846 ( .A(n6795), .ZN(n6794) );
  OAI21_X1 U8847 ( .B1(n6497), .B2(n6796), .A(n11344), .ZN(n6795) );
  AND2_X1 U8848 ( .A1(n6735), .A2(n6733), .ZN(n6554) );
  AND2_X1 U8849 ( .A1(n6743), .A2(n6741), .ZN(n6555) );
  AND2_X1 U8850 ( .A1(n6756), .A2(n6754), .ZN(n6556) );
  NOR2_X1 U8851 ( .A1(n12910), .A2(n12909), .ZN(n6557) );
  NAND2_X1 U8852 ( .A1(n11127), .A2(n11126), .ZN(n6558) );
  NAND2_X1 U8853 ( .A1(n7349), .A2(n7348), .ZN(n7276) );
  INV_X1 U8854 ( .A(n7276), .ZN(n7022) );
  OR2_X1 U8855 ( .A1(n8453), .A2(n7305), .ZN(n6559) );
  NAND2_X1 U8856 ( .A1(n12217), .A2(n12215), .ZN(n6560) );
  INV_X1 U8857 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n7277) );
  INV_X1 U8858 ( .A(n7147), .ZN(n7146) );
  NAND2_X1 U8859 ( .A1(n10753), .A2(n10751), .ZN(n7147) );
  AND2_X1 U8860 ( .A1(n9067), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n6561) );
  AND2_X1 U8861 ( .A1(n8299), .A2(n9083), .ZN(n6562) );
  AND2_X1 U8862 ( .A1(n9647), .A2(n9646), .ZN(n6563) );
  OR2_X1 U8863 ( .A1(n14142), .A2(n14141), .ZN(n6564) );
  AND2_X1 U8864 ( .A1(n9073), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n6565) );
  NAND2_X1 U8865 ( .A1(n14380), .A2(n14381), .ZN(n6566) );
  OR2_X1 U8866 ( .A1(n14146), .A2(n14145), .ZN(n6567) );
  NOR2_X1 U8867 ( .A1(n13410), .A2(n13227), .ZN(n6568) );
  NAND2_X1 U8868 ( .A1(n8941), .A2(n9754), .ZN(n6569) );
  INV_X1 U8869 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9377) );
  AND2_X1 U8870 ( .A1(n7932), .A2(n8886), .ZN(n6570) );
  INV_X1 U8871 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6773) );
  NAND2_X1 U8872 ( .A1(n7716), .A2(n7715), .ZN(n7732) );
  NAND2_X1 U8873 ( .A1(n7678), .A2(n7677), .ZN(n7698) );
  INV_X1 U8874 ( .A(n12594), .ZN(n7935) );
  AND2_X1 U8875 ( .A1(n6499), .A2(n13528), .ZN(n6571) );
  AND2_X1 U8876 ( .A1(n12356), .A2(n11696), .ZN(n6572) );
  INV_X1 U8877 ( .A(n10162), .ZN(n7019) );
  OR2_X1 U8878 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n14148), .ZN(n6573) );
  OR2_X1 U8879 ( .A1(n14152), .A2(n14153), .ZN(n6574) );
  AND2_X1 U8880 ( .A1(n12138), .A2(n8685), .ZN(n6575) );
  INV_X1 U8881 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6819) );
  AND2_X1 U8882 ( .A1(n12752), .A2(n12614), .ZN(n6576) );
  AND2_X1 U8883 ( .A1(n6827), .A2(n14001), .ZN(n6577) );
  INV_X1 U8884 ( .A(n11366), .ZN(n7100) );
  INV_X1 U8885 ( .A(n7466), .ZN(n7026) );
  AND2_X1 U8886 ( .A1(n8235), .A2(n8263), .ZN(n6578) );
  INV_X1 U8887 ( .A(n13242), .ZN(n13247) );
  AND2_X1 U8888 ( .A1(n7627), .A2(n7642), .ZN(n6579) );
  AND2_X1 U8889 ( .A1(n7933), .A2(n6949), .ZN(n6580) );
  NAND2_X1 U8890 ( .A1(n8015), .A2(n6967), .ZN(n6969) );
  INV_X1 U8891 ( .A(n12078), .ZN(n6866) );
  AND2_X1 U8892 ( .A1(n6862), .A2(n13931), .ZN(n6581) );
  AND2_X1 U8893 ( .A1(n7337), .A2(n7393), .ZN(n6582) );
  AND2_X1 U8894 ( .A1(n11656), .A2(n11655), .ZN(n6583) );
  AND2_X1 U8895 ( .A1(n7764), .A2(n7747), .ZN(n6584) );
  AND2_X1 U8896 ( .A1(n7710), .A2(n7694), .ZN(n6585) );
  OR2_X1 U8897 ( .A1(n8273), .A2(n8271), .ZN(n6586) );
  OR2_X1 U8898 ( .A1(n7295), .A2(n8574), .ZN(n6587) );
  OR2_X1 U8899 ( .A1(n7298), .A2(n8610), .ZN(n6588) );
  OR2_X1 U8900 ( .A1(n8489), .A2(n8487), .ZN(n6589) );
  OR2_X1 U8901 ( .A1(n11062), .A2(n6988), .ZN(n6590) );
  OR2_X1 U8902 ( .A1(n7315), .A2(n8196), .ZN(n6591) );
  AND2_X1 U8903 ( .A1(n7233), .A2(n6542), .ZN(n6592) );
  NAND2_X1 U8904 ( .A1(n14140), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n6593) );
  AND2_X1 U8905 ( .A1(n6473), .A2(n6491), .ZN(n6594) );
  INV_X1 U8906 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n7307) );
  NAND2_X1 U8907 ( .A1(n11778), .A2(n11777), .ZN(n6595) );
  INV_X1 U8908 ( .A(n6789), .ZN(n6788) );
  OR2_X1 U8909 ( .A1(n13210), .A2(n6790), .ZN(n6789) );
  INV_X1 U8910 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n8017) );
  NAND2_X2 U8911 ( .A1(n7369), .A2(n12157), .ZN(n7760) );
  INV_X1 U8912 ( .A(n6457), .ZN(n8630) );
  OR2_X1 U8913 ( .A1(n11313), .A2(n11312), .ZN(n6596) );
  INV_X1 U8914 ( .A(n10908), .ZN(n14855) );
  INV_X1 U8915 ( .A(n10897), .ZN(n14819) );
  NAND2_X1 U8916 ( .A1(n7606), .A2(n7605), .ZN(n14282) );
  NAND2_X1 U8917 ( .A1(n6937), .A2(n8840), .ZN(n14281) );
  INV_X1 U8918 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6959) );
  AND3_X1 U8919 ( .A1(n7349), .A2(n7348), .A3(n7277), .ZN(n7612) );
  AND2_X1 U8920 ( .A1(n9467), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6597) );
  INV_X1 U8921 ( .A(n11890), .ZN(n7156) );
  NAND2_X1 U8922 ( .A1(n7348), .A2(n7349), .ZN(n7594) );
  NAND2_X1 U8923 ( .A1(n7571), .A2(n7506), .ZN(n6598) );
  NOR2_X1 U8924 ( .A1(n13975), .A2(n14372), .ZN(n13960) );
  INV_X1 U8925 ( .A(n8359), .ZN(n8397) );
  NAND2_X1 U8926 ( .A1(n7164), .A2(n6497), .ZN(n11285) );
  AND2_X1 U8927 ( .A1(n8426), .A2(SI_17_), .ZN(n6599) );
  INV_X1 U8928 ( .A(n8847), .ZN(n6941) );
  AND2_X1 U8929 ( .A1(n6933), .A2(n6932), .ZN(n6600) );
  INV_X1 U8930 ( .A(n7322), .ZN(n7046) );
  INV_X1 U8931 ( .A(n7331), .ZN(n6674) );
  INV_X1 U8932 ( .A(n13395), .ZN(n13307) );
  AND2_X1 U8933 ( .A1(n13330), .A2(n13154), .ZN(n13395) );
  NAND2_X1 U8934 ( .A1(n7771), .A2(n7770), .ZN(n12667) );
  INV_X1 U8935 ( .A(n12667), .ZN(n7929) );
  INV_X1 U8936 ( .A(n12803), .ZN(n7286) );
  NAND2_X1 U8937 ( .A1(n14911), .A2(n8796), .ZN(n10139) );
  INV_X1 U8938 ( .A(n14748), .ZN(n6650) );
  INV_X1 U8939 ( .A(n6855), .ZN(n6856) );
  AND2_X1 U8940 ( .A1(n7020), .A2(n7019), .ZN(n6601) );
  NAND2_X1 U8941 ( .A1(n7660), .A2(n7643), .ZN(n6602) );
  INV_X1 U8942 ( .A(n7001), .ZN(n7000) );
  NOR2_X1 U8943 ( .A1(n11414), .A2(n7005), .ZN(n7001) );
  OR2_X1 U8944 ( .A1(n12394), .A2(n14317), .ZN(n6603) );
  INV_X1 U8945 ( .A(n6830), .ZN(n11232) );
  NOR2_X1 U8946 ( .A1(n10953), .A2(n6831), .ZN(n6830) );
  AND2_X1 U8947 ( .A1(n11020), .A2(n6468), .ZN(n6604) );
  NOR2_X1 U8948 ( .A1(n7221), .A2(n7218), .ZN(n6605) );
  AND2_X1 U8949 ( .A1(n6663), .A2(n6506), .ZN(n6606) );
  AND2_X1 U8950 ( .A1(n10752), .A2(n10751), .ZN(n6607) );
  AND2_X1 U8951 ( .A1(n6681), .A2(n6596), .ZN(n6608) );
  INV_X1 U8952 ( .A(n7321), .ZN(n7049) );
  INV_X1 U8953 ( .A(n6991), .ZN(n9754) );
  NAND2_X1 U8954 ( .A1(n7976), .A2(n7977), .ZN(n6991) );
  INV_X1 U8955 ( .A(n13018), .ZN(n13034) );
  XOR2_X1 U8956 ( .A(n8675), .B(SI_30_), .Z(n6609) );
  INV_X1 U8957 ( .A(n11693), .ZN(n6634) );
  AND2_X2 U8958 ( .A1(n8958), .A2(n10035), .ZN(n15164) );
  AND3_X2 U8959 ( .A1(n10015), .A2(n14661), .A3(n10170), .ZN(n14731) );
  AND2_X2 U8960 ( .A1(n9577), .A2(n9576), .ZN(n14746) );
  INV_X1 U8961 ( .A(n11327), .ZN(n6833) );
  NAND2_X1 U8962 ( .A1(n7111), .A2(n9985), .ZN(n14632) );
  NAND2_X1 U8963 ( .A1(n9359), .A2(n9358), .ZN(n13018) );
  INV_X1 U8964 ( .A(n10614), .ZN(n6826) );
  NOR2_X1 U8965 ( .A1(n12488), .A2(n12510), .ZN(n6610) );
  INV_X1 U8966 ( .A(n6484), .ZN(n6662) );
  AND2_X1 U8967 ( .A1(n14134), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6611) );
  NOR2_X1 U8968 ( .A1(n12538), .A2(n12793), .ZN(n6612) );
  NOR2_X1 U8969 ( .A1(n7861), .A2(n7067), .ZN(n7066) );
  INV_X1 U8970 ( .A(SI_26_), .ZN(n11404) );
  INV_X1 U8971 ( .A(n13878), .ZN(n10062) );
  NAND2_X1 U8972 ( .A1(n12543), .A2(n10225), .ZN(n9755) );
  INV_X1 U8973 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n6614) );
  INV_X1 U8974 ( .A(SI_14_), .ZN(n6729) );
  INV_X1 U8975 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n14140) );
  INV_X1 U8976 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7385) );
  INV_X1 U8977 ( .A(n7198), .ZN(n6720) );
  INV_X1 U8978 ( .A(n6621), .ZN(n6620) );
  INV_X1 U8979 ( .A(n13245), .ZN(n7144) );
  NAND2_X1 U8980 ( .A1(n8075), .A2(SI_2_), .ZN(n8077) );
  NOR2_X1 U8981 ( .A1(n6463), .A2(n6789), .ZN(n6784) );
  OAI21_X1 U8982 ( .B1(n8467), .B2(n8466), .A(n8465), .ZN(n8483) );
  OAI21_X1 U8983 ( .B1(n13411), .B2(n13495), .A(n7140), .ZN(n13498) );
  NAND2_X1 U8984 ( .A1(n12688), .A2(n12694), .ZN(n7282) );
  INV_X1 U8985 ( .A(n10141), .ZN(n12806) );
  NAND2_X1 U8986 ( .A1(n10210), .A2(n7481), .ZN(n10523) );
  AOI21_X1 U8987 ( .B1(n12598), .B2(n7843), .A(n6576), .ZN(n12583) );
  OR2_X1 U8988 ( .A1(n8959), .A2(n15162), .ZN(n8963) );
  NAND2_X1 U8989 ( .A1(n7805), .A2(n7804), .ZN(n7820) );
  NAND2_X1 U8990 ( .A1(n7754), .A2(n7753), .ZN(n7772) );
  NAND2_X1 U8991 ( .A1(n7494), .A2(n7493), .ZN(n7514) );
  INV_X1 U8992 ( .A(n6920), .ZN(n6919) );
  INV_X1 U8993 ( .A(n12629), .ZN(n6922) );
  NAND2_X1 U8994 ( .A1(n6631), .A2(n8945), .ZN(P3_U3296) );
  NAND3_X1 U8995 ( .A1(n13412), .A2(n13413), .A3(n14680), .ZN(n13415) );
  NAND2_X1 U8996 ( .A1(n9561), .A2(n11806), .ZN(n9565) );
  NAND2_X1 U8997 ( .A1(n10540), .A2(n10539), .ZN(n10760) );
  NAND2_X1 U8998 ( .A1(n7091), .A2(n10763), .ZN(n10816) );
  NAND2_X1 U8999 ( .A1(n7090), .A2(n10814), .ZN(n11149) );
  INV_X1 U9000 ( .A(n13348), .ZN(n6717) );
  NAND2_X1 U9001 ( .A1(n9984), .A2(n6815), .ZN(n7111) );
  NAND2_X1 U9002 ( .A1(n8043), .A2(n8042), .ZN(n8050) );
  OAI21_X1 U9003 ( .B1(n7342), .B2(n8107), .A(n7319), .ZN(n8127) );
  OAI21_X1 U9004 ( .B1(n6503), .B2(n6619), .A(n7301), .ZN(n8289) );
  OAI21_X1 U9005 ( .B1(n8672), .B2(n8671), .A(n8670), .ZN(n8717) );
  NAND2_X1 U9006 ( .A1(n8250), .A2(n6586), .ZN(n6619) );
  OAI21_X1 U9007 ( .B1(n6720), .B2(n6719), .A(n6718), .ZN(n8327) );
  NAND2_X1 U9008 ( .A1(n8303), .A2(n8302), .ZN(n8396) );
  OAI211_X1 U9009 ( .C1(n14405), .C2(n14013), .A(n14012), .B(n14011), .ZN(
        n14094) );
  OAI211_X1 U9010 ( .C1(n7291), .C2(n8149), .A(n8132), .B(n8131), .ZN(n7292)
         );
  INV_X1 U9011 ( .A(n10739), .ZN(n6625) );
  NOR2_X1 U9012 ( .A1(n7945), .A2(n7944), .ZN(n8959) );
  NAND2_X2 U9013 ( .A1(n8969), .A2(n7323), .ZN(n9327) );
  NOR2_X1 U9014 ( .A1(n9719), .A2(n7224), .ZN(n7223) );
  NAND3_X1 U9015 ( .A1(n7251), .A2(n9960), .A3(n7250), .ZN(n9966) );
  INV_X1 U9016 ( .A(n7230), .ZN(n13033) );
  NAND2_X1 U9017 ( .A1(n10120), .A2(n10119), .ZN(n10355) );
  NAND2_X1 U9018 ( .A1(n7236), .A2(n7237), .ZN(n12914) );
  NAND2_X1 U9019 ( .A1(n7553), .A2(n7504), .ZN(n7535) );
  NAND2_X2 U9020 ( .A1(n13832), .A2(n6495), .ZN(n12118) );
  NAND2_X1 U9021 ( .A1(n8117), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n8021) );
  NAND2_X1 U9022 ( .A1(n8015), .A2(n8016), .ZN(n8003) );
  NAND2_X1 U9023 ( .A1(n12104), .A2(n6504), .ZN(n13933) );
  NAND2_X1 U9024 ( .A1(n11231), .A2(n6982), .ZN(n11382) );
  NAND2_X1 U9025 ( .A1(n10633), .A2(n10632), .ZN(n10947) );
  NAND2_X1 U9026 ( .A1(n6952), .A2(n10385), .ZN(n10570) );
  NAND2_X1 U9027 ( .A1(n6975), .A2(n12119), .ZN(n12120) );
  INV_X1 U9028 ( .A(n6629), .ZN(n7947) );
  NAND4_X1 U9029 ( .A1(n6630), .A2(n7275), .A3(n7348), .A4(n7349), .ZN(n6629)
         );
  NAND2_X2 U9030 ( .A1(n13933), .A2(n13934), .ZN(n12106) );
  NAND2_X2 U9031 ( .A1(n6634), .A2(n6635), .ZN(n10277) );
  AND3_X2 U9032 ( .A1(n8032), .A2(n8031), .A3(n8033), .ZN(n11693) );
  AOI21_X1 U9033 ( .B1(n14475), .B2(n14476), .A(n10292), .ZN(n10621) );
  NAND2_X2 U9034 ( .A1(n9560), .A2(n12021), .ZN(n9858) );
  INV_X2 U9035 ( .A(n9086), .ZN(n8969) );
  NAND3_X1 U9036 ( .A1(n9064), .A2(n9006), .A3(n8967), .ZN(n9086) );
  INV_X1 U9037 ( .A(n8971), .ZN(n9137) );
  NOR2_X2 U9038 ( .A1(n9327), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n8971) );
  AOI21_X2 U9039 ( .B1(n11605), .B2(n11604), .A(n11603), .ZN(n11639) );
  NAND2_X2 U9040 ( .A1(n8817), .A2(n8818), .ZN(n10673) );
  NAND2_X1 U9041 ( .A1(n14258), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n14201) );
  INV_X1 U9042 ( .A(n14166), .ZN(n7072) );
  OAI21_X1 U9043 ( .B1(n14173), .B2(n14172), .A(n6593), .ZN(n7070) );
  NAND2_X1 U9044 ( .A1(n6637), .A2(n14601), .ZN(n14203) );
  NAND2_X1 U9045 ( .A1(n14260), .A2(n14261), .ZN(n6637) );
  NAND2_X1 U9046 ( .A1(n14256), .A2(n14255), .ZN(n14188) );
  INV_X1 U9047 ( .A(n7083), .ZN(n14240) );
  NAND2_X1 U9048 ( .A1(n15173), .A2(n15172), .ZN(n6638) );
  INV_X1 U9049 ( .A(n6639), .ZN(n14250) );
  NOR2_X1 U9050 ( .A1(n15176), .A2(n15175), .ZN(n14179) );
  NAND2_X1 U9051 ( .A1(n15167), .A2(n15168), .ZN(n6640) );
  INV_X1 U9052 ( .A(n14427), .ZN(n6706) );
  NOR2_X4 U9053 ( .A1(n13357), .A2(n13442), .ZN(n13331) );
  NOR2_X2 U9054 ( .A1(n10773), .A2(n11862), .ZN(n10821) );
  OR2_X2 U9055 ( .A1(n14635), .A2(n14634), .ZN(n14636) );
  XNOR2_X1 U9056 ( .A(n9923), .B(n12806), .ZN(n9899) );
  NAND2_X1 U9057 ( .A1(n12822), .A2(n14993), .ZN(n6950) );
  AND2_X2 U9058 ( .A1(n10203), .A2(n10192), .ZN(n10689) );
  NAND2_X1 U9059 ( .A1(n11207), .A2(n12375), .ZN(n6644) );
  NAND2_X1 U9060 ( .A1(n12571), .A2(n12570), .ZN(n6951) );
  NAND2_X1 U9061 ( .A1(n6780), .A2(n6782), .ZN(P2_U3528) );
  OAI21_X1 U9062 ( .B1(n13407), .B2(n13495), .A(n13406), .ZN(n6781) );
  INV_X1 U9063 ( .A(n6987), .ZN(n6986) );
  NAND2_X2 U9064 ( .A1(n10065), .A2(n9376), .ZN(n11980) );
  NAND3_X1 U9065 ( .A1(n6771), .A2(n8969), .A3(n7323), .ZN(n9141) );
  AOI21_X2 U9066 ( .B1(n6643), .B2(n14529), .A(n12099), .ZN(n14012) );
  NAND2_X1 U9067 ( .A1(n12096), .A2(n12139), .ZN(n6643) );
  NAND2_X1 U9068 ( .A1(n8158), .A2(n8157), .ZN(n8186) );
  INV_X1 U9069 ( .A(n6869), .ZN(n6867) );
  OAI21_X1 U9070 ( .B1(n8080), .B2(n7193), .A(n8140), .ZN(n7191) );
  OAI21_X1 U9071 ( .B1(n8081), .B2(n7193), .A(n7192), .ZN(n8143) );
  NAND2_X1 U9072 ( .A1(n6994), .A2(n6993), .ZN(n11605) );
  NOR2_X1 U9073 ( .A1(n11062), .A2(n6989), .ZN(n6987) );
  XNOR2_X2 U9074 ( .A(n10673), .B(n11664), .ZN(n10783) );
  NAND2_X1 U9075 ( .A1(n12506), .A2(n6612), .ZN(n6648) );
  NAND2_X1 U9076 ( .A1(n6648), .A2(n6646), .ZN(n6653) );
  XNOR2_X1 U9077 ( .A(n6653), .B(n6652), .ZN(n6651) );
  NAND2_X1 U9078 ( .A1(n12505), .A2(n12510), .ZN(n6654) );
  NAND2_X1 U9079 ( .A1(n10243), .A2(n10242), .ZN(n6663) );
  NAND3_X1 U9080 ( .A1(n6663), .A2(n10600), .A3(n6506), .ZN(n6657) );
  INV_X1 U9081 ( .A(n10602), .ZN(n6665) );
  OAI21_X1 U9082 ( .B1(n13552), .B2(n6671), .A(n6669), .ZN(n13605) );
  NAND2_X1 U9083 ( .A1(n13552), .A2(n6669), .ZN(n6668) );
  NAND2_X1 U9084 ( .A1(n11198), .A2(n6680), .ZN(n6679) );
  INV_X1 U9085 ( .A(n6681), .ZN(n11314) );
  AND2_X1 U9086 ( .A1(n14430), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n6704) );
  OR2_X1 U9087 ( .A1(n14430), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n6705) );
  NAND2_X1 U9088 ( .A1(n7093), .A2(n7094), .ZN(n6715) );
  NAND2_X1 U9089 ( .A1(n7093), .A2(n11151), .ZN(n6716) );
  NAND2_X2 U9090 ( .A1(n6731), .A2(n7385), .ZN(n7187) );
  NAND3_X1 U9091 ( .A1(n7384), .A2(n7383), .A3(P3_ADDR_REG_19__SCAN_IN), .ZN(
        n6731) );
  NAND3_X1 U9092 ( .A1(n14245), .A2(n7382), .A3(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n6732) );
  OR2_X1 U9093 ( .A1(n11850), .A2(n6472), .ZN(n6738) );
  NAND2_X1 U9094 ( .A1(n11850), .A2(n6736), .ZN(n6735) );
  OR2_X1 U9095 ( .A1(n11881), .A2(n6747), .ZN(n6745) );
  NAND2_X1 U9096 ( .A1(n11881), .A2(n6509), .ZN(n6743) );
  NAND2_X1 U9097 ( .A1(n6816), .A2(n8158), .ZN(n6753) );
  NAND2_X1 U9098 ( .A1(n6753), .A2(n7195), .ZN(n8231) );
  OAI21_X1 U9099 ( .B1(n7195), .B2(n8230), .A(n8232), .ZN(n6752) );
  OR2_X1 U9100 ( .A1(n11938), .A2(n6761), .ZN(n6759) );
  NAND2_X1 U9101 ( .A1(n11938), .A2(n6757), .ZN(n6756) );
  NAND2_X1 U9102 ( .A1(n6764), .A2(n6763), .ZN(n11833) );
  OR2_X1 U9103 ( .A1(n6766), .A2(n11831), .ZN(n6763) );
  NAND2_X1 U9104 ( .A1(n6765), .A2(n11830), .ZN(n6764) );
  NAND2_X1 U9105 ( .A1(n6766), .A2(n11831), .ZN(n6765) );
  NOR2_X1 U9106 ( .A1(n9140), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n6771) );
  OAI21_X2 U9107 ( .B1(n9141), .B2(n6773), .A(n6769), .ZN(n7110) );
  NAND2_X1 U9108 ( .A1(n6775), .A2(n6774), .ZN(n13298) );
  AOI21_X2 U9109 ( .B1(n6776), .B2(n6490), .A(n12018), .ZN(n12061) );
  NAND4_X1 U9110 ( .A1(n6778), .A2(n12011), .A3(n12012), .A4(n6777), .ZN(n6776) );
  OR2_X1 U9111 ( .A1(n12007), .A2(n12006), .ZN(n6777) );
  NAND2_X1 U9112 ( .A1(n6779), .A2(n12005), .ZN(n6778) );
  NAND2_X1 U9113 ( .A1(n12007), .A2(n12006), .ZN(n6779) );
  NOR2_X2 U9114 ( .A1(n13405), .A2(n7335), .ZN(n13406) );
  INV_X1 U9115 ( .A(n7164), .ZN(n6793) );
  OAI21_X1 U9116 ( .B1(n7164), .B2(n6796), .A(n6794), .ZN(n11430) );
  OAI211_X2 U9117 ( .C1(n9327), .C2(n6798), .A(n6799), .B(n6801), .ZN(n7109)
         );
  NAND2_X1 U9118 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(n8978), .ZN(n6798) );
  OR2_X1 U9119 ( .A1(n7129), .A2(n7127), .ZN(n6814) );
  NAND2_X1 U9120 ( .A1(n7129), .A2(n6812), .ZN(n6811) );
  NAND3_X1 U9121 ( .A1(n10328), .A2(n6815), .A3(n9565), .ZN(n9566) );
  XNOR2_X1 U9122 ( .A(n11813), .B(n13063), .ZN(n12025) );
  NAND2_X1 U9123 ( .A1(n8155), .A2(n8154), .ZN(n8158) );
  NAND3_X1 U9124 ( .A1(n8702), .A2(n6821), .A3(n8701), .ZN(n6820) );
  NAND3_X1 U9125 ( .A1(n6476), .A2(n6823), .A3(n6575), .ZN(n6822) );
  INV_X1 U9126 ( .A(n8687), .ZN(n13888) );
  OR2_X1 U9127 ( .A1(n11145), .A2(n9335), .ZN(n6825) );
  AND2_X2 U9128 ( .A1(n13838), .A2(n6577), .ZN(n13782) );
  CLKBUF_X1 U9129 ( .A(n6835), .Z(n6834) );
  NAND2_X1 U9130 ( .A1(n9621), .A2(n6835), .ZN(n8148) );
  NAND2_X1 U9131 ( .A1(n9952), .A2(n6834), .ZN(n8214) );
  NAND2_X1 U9132 ( .A1(n10356), .A2(n6834), .ZN(n8286) );
  NAND2_X1 U9133 ( .A1(n10643), .A2(n6834), .ZN(n8346) );
  NAND2_X1 U9134 ( .A1(n10718), .A2(n6834), .ZN(n8331) );
  NAND2_X1 U9135 ( .A1(n11113), .A2(n6834), .ZN(n8313) );
  NAND2_X1 U9136 ( .A1(n11347), .A2(n6834), .ZN(n8405) );
  NAND2_X1 U9137 ( .A1(n11427), .A2(n6834), .ZN(n8416) );
  NAND2_X1 U9138 ( .A1(n11286), .A2(n6834), .ZN(n8366) );
  NAND2_X1 U9139 ( .A1(n11539), .A2(n6834), .ZN(n8431) );
  NAND2_X1 U9140 ( .A1(n11897), .A2(n6834), .ZN(n8446) );
  NAND2_X1 U9141 ( .A1(n11918), .A2(n6834), .ZN(n8469) );
  NAND2_X1 U9142 ( .A1(n11934), .A2(n6834), .ZN(n8486) );
  NAND2_X1 U9143 ( .A1(n11978), .A2(n6834), .ZN(n8546) );
  NAND2_X1 U9144 ( .A1(n11961), .A2(n6834), .ZN(n8521) );
  NAND2_X1 U9145 ( .A1(n12000), .A2(n6834), .ZN(n8573) );
  NAND2_X1 U9146 ( .A1(n11774), .A2(n6834), .ZN(n8589) );
  NAND2_X1 U9147 ( .A1(n13522), .A2(n6834), .ZN(n8609) );
  NAND2_X1 U9148 ( .A1(n11752), .A2(n6834), .ZN(n8623) );
  AOI21_X1 U9149 ( .B1(n11739), .B2(n6834), .A(n8654), .ZN(n14001) );
  NAND2_X1 U9150 ( .A1(n13514), .A2(n6834), .ZN(n8683) );
  NAND2_X1 U9151 ( .A1(n11716), .A2(n6834), .ZN(n8640) );
  NAND2_X2 U9152 ( .A1(n8740), .A2(n14132), .ZN(n9084) );
  XNOR2_X2 U9153 ( .A(n8018), .B(n8017), .ZN(n14132) );
  NAND2_X1 U9155 ( .A1(n11227), .A2(n6508), .ZN(n6838) );
  NAND2_X1 U9156 ( .A1(n6838), .A2(n6839), .ZN(n11451) );
  NAND2_X1 U9157 ( .A1(n6844), .A2(n10285), .ZN(n10391) );
  OAI21_X1 U9158 ( .B1(n10283), .B2(n10613), .A(n6850), .ZN(n6844) );
  NAND3_X1 U9159 ( .A1(n10390), .A2(n6847), .A3(n6845), .ZN(n10394) );
  NAND3_X1 U9160 ( .A1(n6849), .A2(n10285), .A3(n6848), .ZN(n6847) );
  INV_X1 U9161 ( .A(n10613), .ZN(n6848) );
  INV_X1 U9162 ( .A(n10283), .ZN(n6849) );
  OAI21_X1 U9163 ( .B1(n10283), .B2(n10613), .A(n6851), .ZN(n10475) );
  NAND2_X1 U9164 ( .A1(n10948), .A2(n6856), .ZN(n10982) );
  NAND2_X1 U9165 ( .A1(n11455), .A2(n6581), .ZN(n6861) );
  INV_X1 U9166 ( .A(n13873), .ZN(n6868) );
  NAND2_X1 U9167 ( .A1(n13806), .A2(n6876), .ZN(n6875) );
  NOR2_X1 U9168 ( .A1(n6886), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n6958) );
  NAND4_X1 U9169 ( .A1(n8208), .A2(n7992), .A3(n8309), .A4(n7991), .ZN(n6886)
         );
  NAND2_X1 U9170 ( .A1(n13574), .A2(n6894), .ZN(n6892) );
  NAND2_X1 U9171 ( .A1(n6892), .A2(n6893), .ZN(n12270) );
  NAND2_X1 U9172 ( .A1(n6901), .A2(n6900), .ZN(n6902) );
  INV_X1 U9173 ( .A(n9812), .ZN(n6900) );
  INV_X1 U9174 ( .A(n9811), .ZN(n6901) );
  INV_X1 U9175 ( .A(n6902), .ZN(n10098) );
  NAND2_X1 U9176 ( .A1(n8050), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8044) );
  INV_X1 U9177 ( .A(n6904), .ZN(n10855) );
  NOR2_X1 U9178 ( .A1(n14777), .A2(n14776), .ZN(n14775) );
  NAND2_X1 U9179 ( .A1(n6918), .A2(n6916), .ZN(n7378) );
  NOR2_X1 U9180 ( .A1(n7276), .A2(n6917), .ZN(n6916) );
  NAND2_X1 U9181 ( .A1(n12461), .A2(n6610), .ZN(n6923) );
  OAI211_X1 U9182 ( .C1(n12461), .C2(n6926), .A(n6923), .B(n6925), .ZN(n12490)
         );
  INV_X1 U9183 ( .A(n6933), .ZN(n12408) );
  INV_X1 U9184 ( .A(n12409), .ZN(n6932) );
  NAND2_X1 U9185 ( .A1(n11074), .A2(n6936), .ZN(n6934) );
  NOR2_X1 U9186 ( .A1(n11073), .A2(n11074), .ZN(n11076) );
  NOR2_X1 U9187 ( .A1(n10865), .A2(n14312), .ZN(n11073) );
  INV_X1 U9188 ( .A(n11075), .ZN(n6936) );
  OAI21_X2 U9189 ( .B1(n7924), .B2(n6940), .A(n6938), .ZN(n11249) );
  AOI21_X1 U9190 ( .B1(n7927), .B2(n6580), .A(n6943), .ZN(n12642) );
  NAND2_X1 U9191 ( .A1(n10298), .A2(n6952), .ZN(n10321) );
  NAND2_X1 U9192 ( .A1(n10297), .A2(n10389), .ZN(n6952) );
  NAND2_X1 U9193 ( .A1(n6956), .A2(n6953), .ZN(n10471) );
  INV_X1 U9194 ( .A(n6955), .ZN(n10474) );
  NAND2_X2 U9195 ( .A1(n6553), .A2(n8137), .ZN(n13674) );
  NAND3_X1 U9196 ( .A1(n15186), .A2(n6958), .A3(n6464), .ZN(n8362) );
  NAND2_X1 U9197 ( .A1(n6961), .A2(n6962), .ZN(n13948) );
  NAND2_X1 U9198 ( .A1(n11464), .A2(n6964), .ZN(n6961) );
  NAND2_X1 U9199 ( .A1(n12118), .A2(n6594), .ZN(n6970) );
  NAND2_X1 U9200 ( .A1(n6970), .A2(n6971), .ZN(n12137) );
  NAND2_X1 U9201 ( .A1(n12118), .A2(n6473), .ZN(n6975) );
  NAND2_X1 U9202 ( .A1(n12118), .A2(n12117), .ZN(n13787) );
  NAND2_X1 U9203 ( .A1(n11382), .A2(n11381), .ZN(n11458) );
  INV_X1 U9204 ( .A(n11458), .ZN(n11460) );
  NAND2_X1 U9205 ( .A1(n13868), .A2(n6983), .ZN(n13843) );
  NAND2_X1 U9206 ( .A1(n13252), .A2(n13223), .ZN(n13253) );
  NOR2_X2 U9207 ( .A1(n14636), .A2(n14683), .ZN(n10203) );
  NAND2_X1 U9208 ( .A1(n9925), .A2(n6520), .ZN(n10020) );
  XNOR2_X1 U9209 ( .A(n11698), .B(n9890), .ZN(n9923) );
  NAND2_X1 U9210 ( .A1(n6986), .A2(n6985), .ZN(n11207) );
  OAI21_X1 U9211 ( .B1(n11062), .B2(n6988), .A(n11065), .ZN(n6985) );
  AND3_X4 U9212 ( .A1(n6990), .A2(n9756), .A3(n9755), .ZN(n11664) );
  NAND4_X1 U9213 ( .A1(n7977), .A2(n6992), .A3(n7976), .A4(n7957), .ZN(n6990)
         );
  NAND2_X1 U9214 ( .A1(n11277), .A2(n6996), .ZN(n6994) );
  INV_X1 U9215 ( .A(n11276), .ZN(n7006) );
  INV_X1 U9216 ( .A(n11675), .ZN(n7007) );
  AOI21_X1 U9217 ( .B1(n7007), .B2(n6572), .A(n7008), .ZN(n11700) );
  NAND2_X1 U9218 ( .A1(n11675), .A2(n11674), .ZN(n12355) );
  NAND2_X1 U9219 ( .A1(n12330), .A2(n6583), .ZN(n12296) );
  NOR2_X2 U9220 ( .A1(n10496), .A2(n10497), .ZN(n10838) );
  OAI211_X2 U9221 ( .C1(n7015), .C2(n10161), .A(n7016), .B(n10495), .ZN(n10496) );
  NAND2_X1 U9222 ( .A1(n7021), .A2(n7018), .ZN(n7015) );
  NOR2_X2 U9223 ( .A1(n7718), .A2(P3_IR_REG_18__SCAN_IN), .ZN(n7888) );
  NAND2_X1 U9224 ( .A1(n7449), .A2(n7466), .ZN(n7023) );
  NAND2_X1 U9225 ( .A1(n7664), .A2(n7031), .ZN(n7030) );
  NAND2_X1 U9226 ( .A1(n7505), .A2(n7038), .ZN(n7037) );
  NAND2_X1 U9227 ( .A1(n7628), .A2(n6579), .ZN(n7048) );
  NAND2_X1 U9228 ( .A1(n7050), .A2(n7051), .ZN(n7799) );
  NAND2_X1 U9229 ( .A1(n7768), .A2(n7054), .ZN(n7050) );
  NAND2_X1 U9230 ( .A1(n7768), .A2(n7767), .ZN(n7053) );
  NAND2_X1 U9231 ( .A1(n7058), .A2(n6582), .ZN(n7445) );
  NAND3_X1 U9232 ( .A1(n7059), .A2(n7736), .A3(n7748), .ZN(n7749) );
  NAND2_X1 U9233 ( .A1(n7735), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7748) );
  OAI21_X1 U9234 ( .B1(n7551), .B2(n7062), .A(n7060), .ZN(n7520) );
  NAND3_X1 U9235 ( .A1(n7813), .A2(n7801), .A3(n11273), .ZN(n7814) );
  NAND2_X1 U9236 ( .A1(n7845), .A2(n7066), .ZN(n7064) );
  OAI21_X1 U9237 ( .B1(n7845), .B2(n7844), .A(n7846), .ZN(n7862) );
  XNOR2_X1 U9238 ( .A(n14194), .B(n14195), .ZN(n14257) );
  NAND2_X1 U9239 ( .A1(n14434), .A2(n14227), .ZN(n7075) );
  INV_X1 U9240 ( .A(n7079), .ZN(n14437) );
  OAI21_X1 U9241 ( .B1(n14433), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7080), .ZN(
        n7079) );
  OAI211_X1 U9242 ( .C1(n14433), .C2(n7076), .A(n7075), .B(n7074), .ZN(n7081)
         );
  NAND2_X1 U9243 ( .A1(n10816), .A2(n10815), .ZN(n7090) );
  NAND2_X1 U9244 ( .A1(n10772), .A2(n12040), .ZN(n7091) );
  INV_X1 U9245 ( .A(n10196), .ZN(n7104) );
  NAND2_X4 U9246 ( .A1(n9144), .A2(n13525), .ZN(n10065) );
  NAND2_X2 U9247 ( .A1(n7109), .A2(n9141), .ZN(n13525) );
  NAND2_X2 U9248 ( .A1(n7110), .A2(n9345), .ZN(n9144) );
  NAND2_X1 U9249 ( .A1(n10258), .A2(n7113), .ZN(n10702) );
  INV_X1 U9250 ( .A(n13406), .ZN(n7117) );
  NAND2_X1 U9251 ( .A1(n13246), .A2(n7119), .ZN(n7115) );
  OAI211_X1 U9252 ( .C1(n13246), .C2(n13225), .A(n7120), .B(n7115), .ZN(n13407) );
  OAI211_X1 U9253 ( .C1(n13407), .C2(n7118), .A(n7122), .B(n7116), .ZN(
        P2_U3496) );
  INV_X1 U9254 ( .A(n13290), .ZN(n7129) );
  OAI21_X2 U9255 ( .B1(n11984), .B2(n7134), .A(n7133), .ZN(n12007) );
  NAND2_X1 U9256 ( .A1(n9200), .A2(n6467), .ZN(n7135) );
  INV_X1 U9257 ( .A(n9325), .ZN(n7137) );
  NAND2_X1 U9258 ( .A1(n7139), .A2(n7138), .ZN(P2_U3527) );
  AND2_X4 U9259 ( .A1(n9348), .A2(n11629), .ZN(n9628) );
  NAND2_X1 U9260 ( .A1(n9347), .A2(n13515), .ZN(n11629) );
  NAND2_X1 U9261 ( .A1(n7149), .A2(n7150), .ZN(n11965) );
  NAND2_X1 U9262 ( .A1(n11954), .A2(n7152), .ZN(n7149) );
  NAND2_X1 U9263 ( .A1(n7154), .A2(n7155), .ZN(n11889) );
  NAND2_X1 U9264 ( .A1(n11885), .A2(n7157), .ZN(n7154) );
  AOI21_X1 U9265 ( .B1(n7158), .B2(n7157), .A(n7156), .ZN(n7155) );
  NAND2_X1 U9266 ( .A1(n7159), .A2(n7160), .ZN(n11858) );
  NAND2_X1 U9267 ( .A1(n11854), .A2(n7162), .ZN(n7159) );
  AOI21_X1 U9268 ( .B1(n7163), .B2(n7162), .A(n7161), .ZN(n7160) );
  NAND2_X1 U9269 ( .A1(n11155), .A2(n11154), .ZN(n7164) );
  OAI22_X1 U9270 ( .A1(n11922), .A2(n7166), .B1(n11923), .B2(n7165), .ZN(
        n11938) );
  OAI22_X2 U9271 ( .A1(n11864), .A2(n7174), .B1(n11865), .B2(n7173), .ZN(
        n11870) );
  NAND2_X1 U9272 ( .A1(n11870), .A2(n11871), .ZN(n11869) );
  OAI22_X1 U9273 ( .A1(n11877), .A2(n7176), .B1(n11878), .B2(n7175), .ZN(
        n11881) );
  NAND2_X1 U9274 ( .A1(n11904), .A2(n11905), .ZN(n11903) );
  OAI22_X2 U9275 ( .A1(n11845), .A2(n7180), .B1(n11846), .B2(n7179), .ZN(
        n11850) );
  OAI22_X2 U9276 ( .A1(n11833), .A2(n7182), .B1(n11834), .B2(n7181), .ZN(
        n11838) );
  NAND2_X1 U9277 ( .A1(n11838), .A2(n11839), .ZN(n11837) );
  INV_X1 U9278 ( .A(n7187), .ZN(n7185) );
  NAND3_X1 U9279 ( .A1(n7186), .A2(P2_DATAO_REG_1__SCAN_IN), .A3(n7187), .ZN(
        n7183) );
  NAND2_X1 U9280 ( .A1(n8482), .A2(n7189), .ZN(n7188) );
  NAND2_X1 U9281 ( .A1(n7190), .A2(n8484), .ZN(n8498) );
  INV_X1 U9282 ( .A(n7191), .ZN(n7192) );
  NAND2_X1 U9283 ( .A1(n11792), .A2(n11755), .ZN(n11779) );
  NAND2_X1 U9284 ( .A1(n11792), .A2(n7194), .ZN(n12008) );
  NAND2_X1 U9285 ( .A1(n8236), .A2(n6578), .ZN(n7198) );
  NAND2_X1 U9286 ( .A1(n8402), .A2(n7204), .ZN(n7202) );
  NAND2_X1 U9287 ( .A1(n8653), .A2(n8652), .ZN(n7208) );
  OAI21_X1 U9288 ( .B1(n8653), .B2(n7211), .A(n7209), .ZN(n7212) );
  OAI21_X1 U9289 ( .B1(n8652), .B2(n7211), .A(n8676), .ZN(n7210) );
  NAND2_X1 U9290 ( .A1(n8619), .A2(n12884), .ZN(n8620) );
  AND2_X1 U9291 ( .A1(n8979), .A2(n7222), .ZN(n9309) );
  NAND2_X1 U9292 ( .A1(n9411), .A2(n9410), .ZN(n9640) );
  OAI21_X1 U9293 ( .B1(n7231), .B2(n12938), .A(n6592), .ZN(n7230) );
  INV_X1 U9294 ( .A(n6623), .ZN(n7241) );
  NAND2_X1 U9295 ( .A1(n6469), .A2(n12945), .ZN(n7236) );
  NAND2_X1 U9296 ( .A1(n11501), .A2(n7245), .ZN(n11589) );
  NAND2_X1 U9297 ( .A1(n7248), .A2(n7246), .ZN(n10717) );
  INV_X1 U9298 ( .A(n9854), .ZN(n7255) );
  NAND2_X1 U9299 ( .A1(n9662), .A2(n9663), .ZN(n9846) );
  NAND2_X1 U9300 ( .A1(n7257), .A2(n9854), .ZN(n7250) );
  NAND2_X1 U9301 ( .A1(n9662), .A2(n7252), .ZN(n7251) );
  NAND2_X1 U9302 ( .A1(n13031), .A2(n7260), .ZN(n7259) );
  OAI211_X1 U9303 ( .C1(n13031), .C2(n7261), .A(n7259), .B(n12969), .ZN(
        P2_U3192) );
  NAND2_X1 U9304 ( .A1(n12645), .A2(n6470), .ZN(n7273) );
  OAI21_X1 U9305 ( .B1(n12645), .B2(n7274), .A(n6470), .ZN(n12628) );
  NAND3_X1 U9306 ( .A1(n7273), .A2(n7811), .A3(n7272), .ZN(n12613) );
  NAND2_X1 U9307 ( .A1(n7279), .A2(n7278), .ZN(n11250) );
  NAND2_X1 U9308 ( .A1(n7283), .A2(n6534), .ZN(n10210) );
  NAND2_X1 U9309 ( .A1(n14915), .A2(n14916), .ZN(n14914) );
  NAND2_X1 U9310 ( .A1(n7947), .A2(n7359), .ZN(n7951) );
  NAND2_X1 U9311 ( .A1(n7695), .A2(n6585), .ZN(n12716) );
  NAND2_X1 U9312 ( .A1(n7292), .A2(n7290), .ZN(n8170) );
  INV_X1 U9313 ( .A(n8150), .ZN(n7291) );
  NAND2_X1 U9314 ( .A1(n7293), .A2(n7294), .ZN(n8592) );
  NAND3_X1 U9315 ( .A1(n8556), .A2(n6587), .A3(n8555), .ZN(n7293) );
  NAND2_X1 U9316 ( .A1(n7296), .A2(n7297), .ZN(n8658) );
  NAND3_X1 U9317 ( .A1(n8597), .A2(n6588), .A3(n8596), .ZN(n7296) );
  NAND2_X1 U9318 ( .A1(n7299), .A2(n7300), .ZN(n8502) );
  NAND3_X1 U9319 ( .A1(n8474), .A2(n6589), .A3(n8473), .ZN(n7299) );
  NAND2_X1 U9320 ( .A1(n7302), .A2(n7303), .ZN(n8457) );
  INV_X1 U9321 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7306) );
  NAND2_X1 U9322 ( .A1(n8385), .A2(n7312), .ZN(n7310) );
  AND2_X1 U9323 ( .A1(n7310), .A2(n7308), .ZN(n8421) );
  NAND2_X1 U9324 ( .A1(n7310), .A2(n7309), .ZN(n8423) );
  NAND2_X1 U9325 ( .A1(n7313), .A2(n7314), .ZN(n8217) );
  NAND3_X1 U9326 ( .A1(n8175), .A2(n6591), .A3(n8174), .ZN(n7313) );
  NAND2_X1 U9327 ( .A1(n13920), .A2(n12085), .ZN(n13899) );
  NAND2_X1 U9328 ( .A1(n7936), .A2(n7935), .ZN(n12597) );
  INV_X1 U9329 ( .A(n12595), .ZN(n7936) );
  NAND2_X1 U9330 ( .A1(n8924), .A2(n14929), .ZN(n8923) );
  OAI22_X1 U9331 ( .A1(n6635), .A2(n9810), .B1(n11693), .B2(n12174), .ZN(n9801) );
  OR2_X1 U9332 ( .A1(n9394), .A2(n9395), .ZN(n9398) );
  NAND2_X1 U9333 ( .A1(n8537), .A2(n8536), .ZN(n8544) );
  OAI21_X1 U9334 ( .B1(n8074), .B2(n8073), .A(n8072), .ZN(n8093) );
  NAND2_X1 U9335 ( .A1(n8763), .A2(n9751), .ZN(n9753) );
  OR2_X1 U9336 ( .A1(n8483), .A2(n15098), .ZN(n8484) );
  OR2_X1 U9337 ( .A1(n13818), .A2(n13825), .ZN(n13830) );
  NAND2_X1 U9338 ( .A1(n9753), .A2(n7420), .ZN(n14916) );
  NOR2_X2 U9339 ( .A1(n10024), .A2(n10023), .ZN(n10161) );
  NAND2_X1 U9340 ( .A1(n8059), .A2(n8058), .ZN(n8060) );
  XNOR2_X1 U9341 ( .A(n8568), .B(n8564), .ZN(n11978) );
  OAI21_X1 U9342 ( .B1(n13791), .B2(n13790), .A(n14529), .ZN(n13797) );
  INV_X1 U9343 ( .A(n9759), .ZN(n7419) );
  INV_X1 U9344 ( .A(n8170), .ZN(n8173) );
  NAND2_X1 U9345 ( .A1(n8055), .A2(n8690), .ZN(n8057) );
  NAND2_X1 U9346 ( .A1(n13677), .A2(n14512), .ZN(n8101) );
  NAND2_X1 U9347 ( .A1(n9817), .A2(n14486), .ZN(n10281) );
  AND2_X2 U9348 ( .A1(n10156), .A2(n10155), .ZN(n14532) );
  AND2_X1 U9349 ( .A1(n12148), .A2(n14483), .ZN(n14498) );
  INV_X1 U9350 ( .A(n14498), .ZN(n13966) );
  INV_X2 U9351 ( .A(n14991), .ZN(n14993) );
  INV_X1 U9352 ( .A(n13491), .ZN(n10764) );
  AND2_X1 U9353 ( .A1(n14783), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7316) );
  NOR2_X1 U9354 ( .A1(n7915), .A2(n10515), .ZN(n7317) );
  AND2_X1 U9355 ( .A1(n12082), .A2(n12081), .ZN(n7318) );
  NAND2_X2 U9356 ( .A1(n10172), .A2(n14646), .ZN(n13330) );
  INV_X1 U9357 ( .A(n8624), .ZN(n8180) );
  OR2_X1 U9358 ( .A1(n8759), .A2(n12871), .ZN(n7320) );
  AND2_X1 U9359 ( .A1(n8304), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n7321) );
  AND2_X1 U9360 ( .A1(n10067), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n7322) );
  AND2_X1 U9361 ( .A1(n9325), .A2(n8968), .ZN(n7323) );
  AND2_X1 U9362 ( .A1(n14779), .A2(n10885), .ZN(n7324) );
  NOR2_X1 U9363 ( .A1(n12241), .A2(n13587), .ZN(n7326) );
  AND2_X1 U9364 ( .A1(n12894), .A2(n12893), .ZN(n7328) );
  NOR2_X1 U9365 ( .A1(n8103), .A2(n6448), .ZN(n7329) );
  NOR3_X1 U9366 ( .A1(n8354), .A2(n8353), .A3(n8352), .ZN(n7330) );
  NOR2_X1 U9367 ( .A1(n12211), .A2(n13594), .ZN(n7331) );
  INV_X2 U9368 ( .A(n14942), .ZN(n14944) );
  INV_X1 U9369 ( .A(n13331), .ZN(n13342) );
  INV_X1 U9370 ( .A(n13004), .ZN(n13228) );
  INV_X1 U9371 ( .A(n13225), .ZN(n13197) );
  INV_X1 U9372 ( .A(n12646), .ZN(n12678) );
  NAND2_X1 U9373 ( .A1(n7778), .A2(n7777), .ZN(n12646) );
  INV_X1 U9374 ( .A(n9387), .ZN(n11436) );
  INV_X1 U9375 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n9968) );
  NAND2_X1 U9376 ( .A1(n9074), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n7333) );
  OR2_X1 U9377 ( .A1(n9084), .A2(n13712), .ZN(n7334) );
  INV_X1 U9378 ( .A(n12140), .ZN(n12136) );
  NOR2_X1 U9379 ( .A1(n12245), .A2(n13578), .ZN(n7336) );
  NAND2_X1 U9380 ( .A1(n8995), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7337) );
  AND2_X1 U9381 ( .A1(n12865), .A2(n11601), .ZN(n7338) );
  INV_X1 U9382 ( .A(n13887), .ZN(n13903) );
  INV_X1 U9383 ( .A(n7527), .ZN(n7616) );
  OR2_X1 U9384 ( .A1(n13452), .A2(n13177), .ZN(n7339) );
  AND2_X1 U9385 ( .A1(n8060), .A2(n10277), .ZN(n7342) );
  AND2_X1 U9386 ( .A1(n12916), .A2(n12917), .ZN(n7343) );
  INV_X1 U9387 ( .A(n13438), .ZN(n13159) );
  NAND2_X1 U9388 ( .A1(n7329), .A2(n10291), .ZN(n8104) );
  INV_X1 U9389 ( .A(n8171), .ZN(n8172) );
  MUX2_X1 U9390 ( .A(n13672), .B(n14459), .S(n6454), .Z(n8197) );
  MUX2_X1 U9391 ( .A(n13671), .B(n11027), .S(n6454), .Z(n8215) );
  MUX2_X1 U9392 ( .A(n13670), .B(n11204), .S(n6453), .Z(n8247) );
  MUX2_X1 U9393 ( .A(n13669), .B(n11327), .S(n6454), .Z(n8271) );
  MUX2_X1 U9394 ( .A(n13668), .B(n14390), .S(n6453), .Z(n8290) );
  NAND2_X1 U9395 ( .A1(n8377), .A2(n8376), .ZN(n8378) );
  MUX2_X1 U9396 ( .A(n13953), .B(n14372), .S(n6454), .Z(n8422) );
  INV_X1 U9397 ( .A(n8452), .ZN(n8453) );
  NAND2_X1 U9398 ( .A1(n6555), .A2(n7156), .ZN(n11891) );
  MUX2_X1 U9399 ( .A(n13661), .B(n14051), .S(n6453), .Z(n8488) );
  MUX2_X1 U9400 ( .A(n13901), .B(n13888), .S(n6453), .Z(n8500) );
  MUX2_X1 U9401 ( .A(n13659), .B(n14028), .S(n6454), .Z(n8575) );
  NAND2_X1 U9402 ( .A1(n13046), .A2(n12014), .ZN(n11741) );
  INV_X1 U9403 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n7991) );
  INV_X1 U9404 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n7353) );
  INV_X1 U9405 ( .A(n12719), .ZN(n7710) );
  NAND2_X1 U9406 ( .A1(n10395), .A2(n6527), .ZN(n10397) );
  INV_X1 U9407 ( .A(n8779), .ZN(n7859) );
  INV_X1 U9408 ( .A(n7755), .ZN(n7754) );
  INV_X1 U9409 ( .A(n10145), .ZN(n7436) );
  NAND2_X1 U9410 ( .A1(n7931), .A2(n7930), .ZN(n7932) );
  INV_X1 U9411 ( .A(n10214), .ZN(n7480) );
  INV_X1 U9412 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n7358) );
  INV_X1 U9413 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8970) );
  NAND2_X1 U9414 ( .A1(n13869), .A2(n13851), .ZN(n12092) );
  INV_X1 U9415 ( .A(n8425), .ZN(n8426) );
  INV_X1 U9416 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n7650) );
  OAI21_X1 U9417 ( .B1(n8931), .B2(n8930), .A(n8929), .ZN(n8935) );
  INV_X1 U9418 ( .A(n7806), .ZN(n7805) );
  NAND2_X1 U9419 ( .A1(n6462), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10852) );
  INV_X1 U9420 ( .A(n8869), .ZN(n7729) );
  AND2_X1 U9421 ( .A1(n11704), .A2(n12585), .ZN(n7873) );
  INV_X1 U9422 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7362) );
  INV_X1 U9423 ( .A(n11910), .ZN(n11725) );
  INV_X1 U9424 ( .A(n12043), .ZN(n11158) );
  INV_X1 U9425 ( .A(n12040), .ZN(n10753) );
  INV_X1 U9426 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n8223) );
  INV_X1 U9427 ( .A(n11181), .ZN(n11234) );
  INV_X1 U9428 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n7989) );
  INV_X1 U9429 ( .A(n10834), .ZN(n10835) );
  NAND2_X1 U9430 ( .A1(n7651), .A2(n7650), .ZN(n7670) );
  OR2_X1 U9431 ( .A1(n7836), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n7852) );
  AND2_X1 U9432 ( .A1(n10920), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n10863) );
  INV_X1 U9433 ( .A(n12440), .ZN(n12434) );
  NAND2_X1 U9434 ( .A1(n12735), .A2(n12734), .ZN(n12713) );
  NOR2_X1 U9435 ( .A1(n12553), .A2(n12554), .ZN(n7907) );
  OR2_X1 U9436 ( .A1(n8949), .A2(n7943), .ZN(n8946) );
  OR2_X1 U9437 ( .A1(n10523), .A2(n10522), .ZN(n10525) );
  INV_X1 U9438 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n7360) );
  OR2_X1 U9439 ( .A1(n7895), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n7971) );
  INV_X1 U9440 ( .A(n11132), .ZN(n11131) );
  OR2_X1 U9441 ( .A1(n11767), .A2(n12932), .ZN(n11757) );
  NAND2_X1 U9442 ( .A1(n11725), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n11926) );
  NAND2_X1 U9443 ( .A1(n11351), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n11557) );
  INV_X1 U9444 ( .A(n13189), .ZN(n13295) );
  INV_X1 U9445 ( .A(n12047), .ZN(n11546) );
  NAND2_X1 U9446 ( .A1(n10765), .A2(n10764), .ZN(n10773) );
  AND2_X1 U9447 ( .A1(n9373), .A2(n9144), .ZN(n12987) );
  NAND2_X1 U9448 ( .A1(n13226), .A2(n13391), .ZN(n13233) );
  OAI22_X1 U9449 ( .A1(n10817), .A2(n10756), .B1(n10755), .B2(n11862), .ZN(
        n11155) );
  NAND2_X1 U9450 ( .A1(n13064), .A2(n14667), .ZN(n9562) );
  OR2_X1 U9451 ( .A1(n9886), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n10042) );
  INV_X1 U9452 ( .A(n14342), .ZN(n12168) );
  INV_X1 U9453 ( .A(n10239), .ZN(n10241) );
  OR2_X1 U9454 ( .A1(n8224), .A2(n8223), .ZN(n8252) );
  INV_X1 U9455 ( .A(n11463), .ZN(n11454) );
  INV_X1 U9456 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n14139) );
  NOR2_X1 U9457 ( .A1(n14213), .A2(n14212), .ZN(n14157) );
  INV_X1 U9458 ( .A(n12600), .ZN(n12567) );
  NAND2_X1 U9459 ( .A1(n7686), .A2(n7685), .ZN(n7704) );
  OR2_X1 U9460 ( .A1(n9758), .A2(n9757), .ZN(n12361) );
  OR2_X1 U9461 ( .A1(n7760), .A2(n9546), .ZN(n7414) );
  INV_X1 U9462 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n10025) );
  INV_X1 U9463 ( .A(n11086), .ZN(n10864) );
  OR2_X1 U9464 ( .A1(n7866), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n11631) );
  AND2_X1 U9465 ( .A1(n8852), .A2(n8860), .ZN(n11396) );
  AND2_X1 U9466 ( .A1(n9526), .A2(n14957), .ZN(n10030) );
  OR2_X1 U9467 ( .A1(n8948), .A2(n8947), .ZN(n10034) );
  INV_X1 U9468 ( .A(n14917), .ZN(n14284) );
  NAND2_X1 U9469 ( .A1(n7942), .A2(n8946), .ZN(n12804) );
  AND2_X1 U9470 ( .A1(n7978), .A2(n8937), .ZN(n14303) );
  OAI22_X1 U9471 ( .A1(n8747), .A2(n8746), .B1(P2_DATAO_REG_29__SCAN_IN), .B2(
        n11737), .ZN(n8758) );
  OAI21_X1 U9472 ( .B1(n7971), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7973) );
  INV_X1 U9473 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7736) );
  INV_X1 U9474 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n7630) );
  INV_X1 U9475 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n7474) );
  OR2_X1 U9476 ( .A1(n10724), .A2(n10723), .ZN(n11132) );
  OR2_X1 U9477 ( .A1(n11942), .A2(n11941), .ZN(n11969) );
  NAND2_X1 U9478 ( .A1(n12918), .A2(n12920), .ZN(n12921) );
  OR2_X1 U9479 ( .A1(n11969), .A2(n11727), .ZN(n11988) );
  NAND2_X1 U9480 ( .A1(n10359), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n10724) );
  AND2_X1 U9481 ( .A1(n9404), .A2(n9639), .ZN(n9411) );
  INV_X1 U9482 ( .A(n13025), .ZN(n13038) );
  INV_X1 U9483 ( .A(n9359), .ZN(n9341) );
  INV_X1 U9484 ( .A(n7325), .ZN(n11991) );
  CLKBUF_X3 U9485 ( .A(n9387), .Z(n11971) );
  INV_X1 U9486 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n14585) );
  OR2_X1 U9487 ( .A1(n9450), .A2(n9451), .ZN(n9713) );
  AND2_X1 U9488 ( .A1(n9918), .A2(n9919), .ZN(n10339) );
  INV_X1 U9489 ( .A(n13166), .ZN(n13160) );
  NAND2_X1 U9490 ( .A1(n13372), .A2(n13377), .ZN(n13373) );
  NAND2_X1 U9491 ( .A1(n11300), .A2(n11304), .ZN(n11363) );
  INV_X1 U9492 ( .A(n14723), .ZN(n14711) );
  AND2_X1 U9493 ( .A1(n11721), .A2(n9567), .ZN(n14640) );
  INV_X1 U9494 ( .A(n14634), .ZN(n14677) );
  AND2_X1 U9495 ( .A1(n12063), .A2(n10176), .ZN(n11797) );
  INV_X1 U9496 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8974) );
  INV_X1 U9497 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8314) );
  NOR2_X1 U9498 ( .A1(n13543), .A2(n13544), .ZN(n10105) );
  NAND2_X1 U9499 ( .A1(n11018), .A2(n11017), .ZN(n11019) );
  INV_X1 U9500 ( .A(n13668), .ZN(n11532) );
  INV_X1 U9501 ( .A(n13828), .ZN(n13792) );
  AND2_X1 U9502 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n8133) );
  NOR2_X1 U9503 ( .A1(n8458), .A2(n13600), .ZN(n8475) );
  INV_X1 U9504 ( .A(n13669), .ZN(n14379) );
  AOI21_X1 U9505 ( .B1(n8712), .B2(n9825), .A(n8711), .ZN(n8713) );
  OR2_X1 U9506 ( .A1(n8448), .A2(n8447), .ZN(n8458) );
  NAND2_X1 U9507 ( .A1(n14137), .A2(n9273), .ZN(n9814) );
  INV_X1 U9508 ( .A(n13931), .ZN(n13934) );
  NAND2_X1 U9509 ( .A1(n11181), .A2(n12167), .ZN(n11383) );
  INV_X1 U9510 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n8320) );
  NOR2_X1 U9511 ( .A1(n10305), .A2(n9816), .ZN(n10153) );
  NAND2_X1 U9512 ( .A1(n14004), .A2(n14003), .ZN(n14005) );
  INV_X1 U9513 ( .A(n13961), .ZN(n14490) );
  NAND2_X1 U9514 ( .A1(n9693), .A2(n9692), .ZN(n14511) );
  INV_X1 U9515 ( .A(n10291), .ZN(n14476) );
  AND2_X1 U9516 ( .A1(n9256), .A2(n9255), .ZN(n10308) );
  AND2_X1 U9517 ( .A1(n8280), .A2(n8262), .ZN(n8263) );
  INV_X1 U9518 ( .A(n14206), .ZN(n14207) );
  OR2_X1 U9519 ( .A1(n9526), .A2(n9525), .ZN(n9551) );
  INV_X1 U9520 ( .A(n12366), .ZN(n12346) );
  AND2_X1 U9521 ( .A1(n7827), .A2(n7826), .ZN(n12362) );
  INV_X1 U9522 ( .A(n6460), .ZN(n7901) );
  INV_X1 U9523 ( .A(n14876), .ZN(n14906) );
  AND2_X1 U9524 ( .A1(n9545), .A2(n9544), .ZN(n14752) );
  INV_X1 U9525 ( .A(n12727), .ZN(n12739) );
  AND2_X2 U9526 ( .A1(n10030), .A2(n14929), .ZN(n14938) );
  INV_X1 U9527 ( .A(n14979), .ZN(n14957) );
  AND4_X1 U9528 ( .A1(n9526), .A2(n8957), .A3(n8956), .A4(n8955), .ZN(n10035)
         );
  OR2_X1 U9529 ( .A1(n12804), .A2(n14989), .ZN(n14323) );
  AND2_X1 U9530 ( .A1(n7943), .A2(n14929), .ZN(n14989) );
  NAND2_X1 U9531 ( .A1(n7960), .A2(n7959), .ZN(n10031) );
  INV_X1 U9532 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n7522) );
  INV_X1 U9533 ( .A(n13015), .ZN(n13040) );
  AND2_X1 U9534 ( .A1(n14723), .A2(n9357), .ZN(n9358) );
  OR2_X1 U9535 ( .A1(n13250), .A2(n11991), .ZN(n11751) );
  INV_X1 U9536 ( .A(n9628), .ZN(n11995) );
  INV_X1 U9537 ( .A(n14618), .ZN(n14594) );
  AND2_X1 U9538 ( .A1(n9713), .A2(n9712), .ZN(n9716) );
  INV_X1 U9539 ( .A(n14614), .ZN(n14579) );
  XNOR2_X1 U9540 ( .A(n13169), .B(n13160), .ZN(n13161) );
  INV_X1 U9541 ( .A(n14640), .ZN(n13391) );
  AND2_X1 U9542 ( .A1(n9338), .A2(n14661), .ZN(n9576) );
  NAND2_X1 U9543 ( .A1(n10173), .A2(n12071), .ZN(n14723) );
  AND2_X1 U9544 ( .A1(n14718), .A2(n14693), .ZN(n13495) );
  INV_X1 U9545 ( .A(n14693), .ZN(n14728) );
  AND2_X1 U9546 ( .A1(n11797), .A2(n12062), .ZN(n14671) );
  AND2_X1 U9547 ( .A1(n9331), .A2(n11219), .ZN(n9337) );
  INV_X1 U9548 ( .A(n8980), .ZN(n8987) );
  AND2_X1 U9549 ( .A1(n8274), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n8335) );
  AND4_X1 U9550 ( .A1(n8534), .A2(n8533), .A3(n8532), .A4(n8531), .ZN(n13581)
         );
  AND2_X1 U9551 ( .A1(n8464), .A2(n8463), .ZN(n13938) );
  INV_X1 U9552 ( .A(n13764), .ZN(n14445) );
  INV_X1 U9553 ( .A(n14451), .ZN(n13766) );
  INV_X1 U9554 ( .A(n13978), .ZN(n14487) );
  NOR2_X1 U9555 ( .A1(n13941), .A2(n14478), .ZN(n12154) );
  AND2_X1 U9556 ( .A1(n10302), .A2(n10153), .ZN(n9271) );
  INV_X1 U9557 ( .A(n14529), .ZN(n14478) );
  INV_X1 U9558 ( .A(n14511), .ZN(n14522) );
  NAND2_X1 U9559 ( .A1(n9275), .A2(n9274), .ZN(n14529) );
  NAND2_X1 U9560 ( .A1(n9118), .A2(n9121), .ZN(n9268) );
  AND2_X1 U9561 ( .A1(n8267), .A2(n8241), .ZN(n9602) );
  AND2_X1 U9562 ( .A1(n9376), .A2(P1_U3086), .ZN(n11242) );
  INV_X1 U9563 ( .A(n14198), .ZN(n14199) );
  AND2_X1 U9564 ( .A1(n9552), .A2(n9551), .ZN(n14879) );
  INV_X1 U9565 ( .A(n11652), .ZN(n12780) );
  INV_X1 U9566 ( .A(n12364), .ZN(n12354) );
  AND2_X1 U9567 ( .A1(n8756), .A2(n7904), .ZN(n12553) );
  INV_X1 U9568 ( .A(n12659), .ZN(n12626) );
  INV_X1 U9569 ( .A(n12732), .ZN(n12372) );
  INV_X1 U9570 ( .A(P3_U3897), .ZN(n12385) );
  INV_X1 U9571 ( .A(n14879), .ZN(n14910) );
  INV_X1 U9572 ( .A(n14752), .ZN(n14901) );
  INV_X1 U9573 ( .A(n12813), .ZN(n11633) );
  INV_X1 U9574 ( .A(n14939), .ZN(n12607) );
  INV_X1 U9575 ( .A(n8961), .ZN(n8962) );
  NAND2_X1 U9576 ( .A1(n15164), .A2(n14957), .ZN(n12803) );
  INV_X1 U9577 ( .A(n15164), .ZN(n15162) );
  INV_X1 U9578 ( .A(n7987), .ZN(n7988) );
  OR2_X1 U9579 ( .A1(n12782), .A2(n12781), .ZN(n12849) );
  AND2_X1 U9580 ( .A1(n7984), .A2(n7983), .ZN(n14991) );
  INV_X1 U9581 ( .A(SI_25_), .ZN(n11341) );
  INV_X1 U9582 ( .A(SI_20_), .ZN(n15098) );
  INV_X1 U9583 ( .A(n12407), .ZN(n12423) );
  INV_X1 U9584 ( .A(SI_10_), .ZN(n9061) );
  CLKBUF_X1 U9585 ( .A(n12870), .Z(n12883) );
  INV_X1 U9586 ( .A(n13026), .ZN(n13043) );
  NAND2_X1 U9587 ( .A1(n11751), .A2(n11750), .ZN(n13224) );
  INV_X1 U9588 ( .A(n14586), .ZN(n14604) );
  OR2_X1 U9589 ( .A1(n9164), .A2(n13525), .ZN(n14614) );
  OR2_X1 U9590 ( .A1(n9148), .A2(P2_U3088), .ZN(n14602) );
  NAND2_X1 U9591 ( .A1(n13330), .A2(n14650), .ZN(n13397) );
  INV_X1 U9592 ( .A(n14746), .ZN(n14744) );
  AND4_X1 U9593 ( .A1(n14698), .A2(n14697), .A3(n14696), .A4(n14695), .ZN(
        n14739) );
  INV_X1 U9594 ( .A(n14731), .ZN(n14729) );
  NOR2_X1 U9595 ( .A1(n14659), .A2(n14654), .ZN(n14655) );
  INV_X1 U9596 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n9733) );
  NAND2_X1 U9597 ( .A1(n9826), .A2(n9815), .ZN(n14384) );
  OR2_X1 U9598 ( .A1(n9122), .A2(n9418), .ZN(n13675) );
  INV_X1 U9599 ( .A(n14448), .ZN(n13722) );
  NAND2_X1 U9600 ( .A1(n13966), .A2(n10436), .ZN(n13991) );
  INV_X1 U9601 ( .A(n12154), .ZN(n14274) );
  NAND2_X1 U9602 ( .A1(n13966), .A2(n14263), .ZN(n13978) );
  NAND2_X1 U9603 ( .A1(n14540), .A2(n14522), .ZN(n14084) );
  INV_X1 U9604 ( .A(n14540), .ZN(n14537) );
  INV_X1 U9605 ( .A(n13781), .ZN(n14092) );
  INV_X1 U9606 ( .A(n14532), .ZN(n14530) );
  NAND2_X1 U9607 ( .A1(n9268), .A2(n9119), .ZN(n14500) );
  INV_X1 U9608 ( .A(n9824), .ZN(n14137) );
  INV_X1 U9609 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10046) );
  INV_X1 U9610 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9237) );
  INV_X1 U9611 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9067) );
  OAI21_X1 U9612 ( .B1(n8959), .B2(n14991), .A(n7988), .ZN(P3_U3456) );
  AND2_X1 U9613 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9143), .ZN(P2_U3947) );
  INV_X1 U9614 ( .A(n13675), .ZN(P1_U4016) );
  NOR2_X1 U9615 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n7347) );
  NOR2_X1 U9616 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), .ZN(
        n7356) );
  NOR2_X1 U9617 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), .ZN(
        n7355) );
  NAND4_X1 U9618 ( .A1(n7356), .A2(n7355), .A3(n7354), .A4(n7353), .ZN(n7357)
         );
  INV_X1 U9619 ( .A(n7363), .ZN(n7376) );
  NAND2_X1 U9620 ( .A1(n7376), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7361) );
  NAND2_X1 U9621 ( .A1(n7363), .A2(n7362), .ZN(n7364) );
  XNOR2_X2 U9622 ( .A(n7365), .B(n12869), .ZN(n7368) );
  AND2_X2 U9623 ( .A1(n12157), .A2(n7368), .ZN(n7527) );
  NAND2_X1 U9624 ( .A1(n7527), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n7373) );
  NAND2_X1 U9625 ( .A1(n6460), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n7372) );
  INV_X1 U9626 ( .A(n7368), .ZN(n7369) );
  NAND2_X1 U9627 ( .A1(n7898), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7371) );
  AND2_X2 U9628 ( .A1(n7369), .A2(n7367), .ZN(n7542) );
  NAND2_X1 U9629 ( .A1(n7542), .A2(n10149), .ZN(n7370) );
  INV_X1 U9630 ( .A(n7374), .ZN(n7380) );
  NAND2_X1 U9631 ( .A1(n7380), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7375) );
  NAND2_X1 U9632 ( .A1(n7378), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7379) );
  NAND2_X4 U9633 ( .A1(n12880), .A2(n6446), .ZN(n9530) );
  INV_X2 U9634 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7384) );
  NAND2_X4 U9635 ( .A1(n9530), .A2(n6461), .ZN(n8759) );
  OR2_X1 U9636 ( .A1(n8759), .A2(SI_3_), .ZN(n7400) );
  NAND2_X2 U9637 ( .A1(n9530), .A2(n9376), .ZN(n7739) );
  INV_X1 U9638 ( .A(n7417), .ZN(n7388) );
  NAND2_X1 U9639 ( .A1(n7404), .A2(n7388), .ZN(n7390) );
  NAND2_X1 U9640 ( .A1(n9377), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7389) );
  INV_X1 U9641 ( .A(n7426), .ZN(n7392) );
  NAND2_X1 U9642 ( .A1(n9396), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7391) );
  NAND2_X1 U9643 ( .A1(n9001), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7393) );
  XNOR2_X1 U9644 ( .A(n9039), .B(P2_DATAO_REG_3__SCAN_IN), .ZN(n7394) );
  XNOR2_X1 U9645 ( .A(n7443), .B(n7394), .ZN(n9054) );
  OR2_X1 U9646 ( .A1(n7739), .A2(n9054), .ZN(n7399) );
  INV_X1 U9647 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n7397) );
  NAND2_X1 U9648 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n7395), .ZN(n7396) );
  XNOR2_X1 U9649 ( .A(n7397), .B(n7396), .ZN(n14766) );
  NAND2_X1 U9650 ( .A1(n7427), .A2(n14766), .ZN(n7398) );
  NAND2_X1 U9651 ( .A1(n14918), .A2(n10148), .ZN(n8801) );
  INV_X1 U9652 ( .A(n10148), .ZN(n7401) );
  NAND2_X1 U9653 ( .A1(n12383), .A2(n7401), .ZN(n8802) );
  NAND2_X1 U9654 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n7403) );
  INV_X1 U9655 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7402) );
  INV_X1 U9656 ( .A(SI_1_), .ZN(n9050) );
  XNOR2_X1 U9657 ( .A(n7404), .B(n7417), .ZN(n9051) );
  OR2_X1 U9658 ( .A1(n7739), .A2(n9051), .ZN(n7405) );
  OAI211_X2 U9659 ( .C1(n9530), .C2(n6465), .A(n7406), .B(n7405), .ZN(n9759)
         );
  NAND2_X1 U9660 ( .A1(n7527), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n7411) );
  NAND2_X1 U9661 ( .A1(n7542), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n7410) );
  INV_X1 U9662 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n7407) );
  OR2_X1 U9663 ( .A1(n7760), .A2(n7407), .ZN(n7408) );
  INV_X1 U9664 ( .A(n14920), .ZN(n12384) );
  NAND2_X1 U9665 ( .A1(n7419), .A2(n12384), .ZN(n8792) );
  NAND2_X1 U9666 ( .A1(n14920), .A2(n9759), .ZN(n8789) );
  NAND2_X1 U9667 ( .A1(n6458), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n7415) );
  NAND2_X1 U9668 ( .A1(n7542), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n7413) );
  NAND2_X1 U9669 ( .A1(n7527), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n7412) );
  NAND4_X1 U9670 ( .A1(n7415), .A2(n7414), .A3(n7413), .A4(n7412), .ZN(n7910)
         );
  INV_X1 U9671 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8013) );
  NAND2_X1 U9672 ( .A1(n8013), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7416) );
  NAND2_X1 U9673 ( .A1(n7417), .A2(n7416), .ZN(n7418) );
  MUX2_X1 U9674 ( .A(n7418), .B(SI_0_), .S(n6461), .Z(n12888) );
  MUX2_X1 U9675 ( .A(P3_IR_REG_0__SCAN_IN), .B(n12888), .S(n9530), .Z(n9891)
         );
  NAND2_X1 U9676 ( .A1(n12805), .A2(n9891), .ZN(n9751) );
  NAND2_X1 U9677 ( .A1(n14920), .A2(n7419), .ZN(n7420) );
  NAND2_X1 U9678 ( .A1(n7527), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n7424) );
  NAND2_X1 U9679 ( .A1(n6460), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7423) );
  NAND2_X1 U9680 ( .A1(n7898), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7422) );
  NAND2_X1 U9681 ( .A1(n7542), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n7421) );
  AND4_X2 U9682 ( .A1(n7424), .A2(n7423), .A3(n7422), .A4(n7421), .ZN(n10141)
         );
  OR2_X1 U9683 ( .A1(n8759), .A2(SI_2_), .ZN(n7434) );
  XNOR2_X1 U9684 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n7425) );
  XNOR2_X1 U9685 ( .A(n7426), .B(n7425), .ZN(n9002) );
  OR2_X1 U9686 ( .A1(n7739), .A2(n9002), .ZN(n7433) );
  INV_X1 U9687 ( .A(n7428), .ZN(n7429) );
  INV_X1 U9688 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7430) );
  NAND2_X1 U9689 ( .A1(n7427), .A2(n6462), .ZN(n7432) );
  NAND2_X1 U9690 ( .A1(n10141), .A2(n9890), .ZN(n8796) );
  NAND2_X1 U9691 ( .A1(n12806), .A2(n14927), .ZN(n8797) );
  NAND2_X1 U9692 ( .A1(n10141), .A2(n14927), .ZN(n7435) );
  NAND2_X1 U9693 ( .A1(n12383), .A2(n10148), .ZN(n7437) );
  NAND2_X1 U9694 ( .A1(n7527), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n7442) );
  NAND2_X1 U9695 ( .A1(n7541), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7441) );
  NAND2_X1 U9696 ( .A1(n10149), .A2(n10025), .ZN(n7460) );
  NAND2_X1 U9697 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n7438) );
  NAND2_X1 U9698 ( .A1(n7460), .A2(n7438), .ZN(n10235) );
  NAND2_X1 U9699 ( .A1(n7822), .A2(n10235), .ZN(n7440) );
  NAND2_X1 U9700 ( .A1(n6460), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n7439) );
  AND4_X2 U9701 ( .A1(n7442), .A2(n7441), .A3(n7440), .A4(n7439), .ZN(n10164)
         );
  OR2_X1 U9702 ( .A1(n8759), .A2(SI_4_), .ZN(n7455) );
  NAND2_X1 U9703 ( .A1(n9039), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7444) );
  NAND2_X1 U9704 ( .A1(n9005), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n7466) );
  NAND2_X1 U9705 ( .A1(n9011), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n7446) );
  NAND2_X1 U9706 ( .A1(n7466), .A2(n7446), .ZN(n7448) );
  INV_X1 U9707 ( .A(n7448), .ZN(n7447) );
  NAND2_X1 U9708 ( .A1(n7449), .A2(n7448), .ZN(n7450) );
  AND2_X1 U9709 ( .A1(n7467), .A2(n7450), .ZN(n9057) );
  OR2_X1 U9710 ( .A1(n7739), .A2(n9057), .ZN(n7454) );
  NAND2_X1 U9711 ( .A1(n7472), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7452) );
  INV_X1 U9712 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n7451) );
  XNOR2_X1 U9713 ( .A(n7452), .B(n7451), .ZN(n14783) );
  NAND2_X1 U9714 ( .A1(n7427), .A2(n14783), .ZN(n7453) );
  NAND2_X1 U9715 ( .A1(n10164), .A2(n14958), .ZN(n10213) );
  INV_X1 U9716 ( .A(n10164), .ZN(n12382) );
  INV_X1 U9717 ( .A(n14958), .ZN(n7456) );
  NAND2_X1 U9718 ( .A1(n12382), .A2(n7456), .ZN(n8806) );
  NAND2_X1 U9719 ( .A1(n10213), .A2(n8806), .ZN(n7912) );
  NAND2_X1 U9720 ( .A1(n12382), .A2(n14958), .ZN(n7457) );
  NAND2_X1 U9721 ( .A1(n7527), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n7465) );
  NAND2_X1 U9722 ( .A1(n7898), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7464) );
  INV_X1 U9723 ( .A(n7460), .ZN(n7459) );
  NAND2_X1 U9724 ( .A1(n7459), .A2(n7458), .ZN(n7482) );
  NAND2_X1 U9725 ( .A1(n7460), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n7461) );
  NAND2_X1 U9726 ( .A1(n7482), .A2(n7461), .ZN(n10220) );
  NAND2_X1 U9727 ( .A1(n7822), .A2(n10220), .ZN(n7463) );
  NAND2_X1 U9728 ( .A1(n6459), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n7462) );
  AND4_X2 U9729 ( .A1(n7465), .A2(n7464), .A3(n7463), .A4(n7462), .ZN(n10520)
         );
  OR2_X1 U9730 ( .A1(n8759), .A2(SI_5_), .ZN(n7479) );
  NAND2_X1 U9731 ( .A1(n9017), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n7489) );
  NAND2_X1 U9732 ( .A1(n9049), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n7468) );
  NAND2_X1 U9733 ( .A1(n7489), .A2(n7468), .ZN(n7469) );
  NAND2_X1 U9734 ( .A1(n6551), .A2(n7469), .ZN(n7471) );
  INV_X1 U9735 ( .A(n7469), .ZN(n7470) );
  AND2_X1 U9736 ( .A1(n7471), .A2(n7490), .ZN(n8998) );
  OR2_X1 U9737 ( .A1(n7739), .A2(n8998), .ZN(n7478) );
  NOR2_X1 U9738 ( .A1(n7472), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n7475) );
  OR2_X1 U9739 ( .A1(n7475), .A2(n7630), .ZN(n7473) );
  MUX2_X1 U9740 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7473), .S(
        P3_IR_REG_5__SCAN_IN), .Z(n7476) );
  NAND2_X1 U9741 ( .A1(n7475), .A2(n7474), .ZN(n7508) );
  NAND2_X1 U9742 ( .A1(n7476), .A2(n7508), .ZN(n14802) );
  NAND2_X1 U9743 ( .A1(n7427), .A2(n14802), .ZN(n7477) );
  NAND2_X1 U9744 ( .A1(n10520), .A2(n10166), .ZN(n8810) );
  INV_X1 U9745 ( .A(n10520), .ZN(n12381) );
  INV_X1 U9746 ( .A(n10166), .ZN(n10219) );
  NAND2_X1 U9747 ( .A1(n12381), .A2(n10219), .ZN(n8808) );
  NAND2_X1 U9748 ( .A1(n10520), .A2(n10219), .ZN(n7481) );
  NAND2_X1 U9749 ( .A1(n7527), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n7487) );
  NAND2_X1 U9750 ( .A1(n6459), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n7486) );
  NAND2_X1 U9751 ( .A1(n7482), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7483) );
  NAND2_X1 U9752 ( .A1(n7543), .A2(n7483), .ZN(n10530) );
  NAND2_X1 U9753 ( .A1(n7822), .A2(n10530), .ZN(n7485) );
  NAND2_X1 U9754 ( .A1(n7898), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7484) );
  NAND2_X1 U9755 ( .A1(n7508), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7488) );
  XNOR2_X1 U9756 ( .A(n7488), .B(P3_IR_REG_6__SCAN_IN), .ZN(n10897) );
  INV_X1 U9757 ( .A(SI_6_), .ZN(n9052) );
  OR2_X1 U9758 ( .A1(n8759), .A2(n9052), .ZN(n7492) );
  NAND2_X1 U9759 ( .A1(n7490), .A2(n7489), .ZN(n7502) );
  XNOR2_X1 U9760 ( .A(n7502), .B(n7500), .ZN(n9053) );
  OR2_X1 U9761 ( .A1(n7739), .A2(n9053), .ZN(n7491) );
  OAI211_X1 U9762 ( .C1(n9530), .C2(n14819), .A(n7492), .B(n7491), .ZN(n10531)
         );
  NAND2_X1 U9763 ( .A1(n10485), .A2(n10531), .ZN(n10423) );
  INV_X1 U9764 ( .A(n10531), .ZN(n14967) );
  NAND2_X1 U9765 ( .A1(n12380), .A2(n14967), .ZN(n8813) );
  NAND2_X1 U9766 ( .A1(n12380), .A2(n10531), .ZN(n10421) );
  INV_X2 U9767 ( .A(n7760), .ZN(n7898) );
  NAND2_X1 U9768 ( .A1(n7541), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7499) );
  NAND2_X1 U9769 ( .A1(n7600), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n7498) );
  INV_X1 U9770 ( .A(n7529), .ZN(n7494) );
  NAND2_X1 U9771 ( .A1(n7514), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7495) );
  NAND2_X1 U9772 ( .A1(n7578), .A2(n7495), .ZN(n10841) );
  NAND2_X1 U9773 ( .A1(n7822), .A2(n10841), .ZN(n7497) );
  NAND2_X1 U9774 ( .A1(n6459), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7496) );
  NAND4_X1 U9775 ( .A1(n7499), .A2(n7498), .A3(n7497), .A4(n7496), .ZN(n12376)
         );
  INV_X1 U9776 ( .A(n7500), .ZN(n7501) );
  NAND2_X1 U9777 ( .A1(n9043), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n7504) );
  NAND2_X1 U9778 ( .A1(n9029), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n7503) );
  NAND2_X1 U9779 ( .A1(n7504), .A2(n7503), .ZN(n7550) );
  INV_X1 U9780 ( .A(n7520), .ZN(n7505) );
  NAND2_X1 U9781 ( .A1(n9081), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n7571) );
  NAND2_X1 U9782 ( .A1(n9079), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n7506) );
  NAND2_X1 U9783 ( .A1(n6481), .A2(n6598), .ZN(n7507) );
  NAND2_X1 U9784 ( .A1(n7572), .A2(n7507), .ZN(n9060) );
  NAND2_X1 U9785 ( .A1(n9060), .A2(n8761), .ZN(n7512) );
  NOR2_X1 U9786 ( .A1(n7536), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n7521) );
  NAND2_X1 U9787 ( .A1(n7521), .A2(n7522), .ZN(n7573) );
  NAND2_X1 U9788 ( .A1(n7573), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7510) );
  INV_X1 U9789 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n7509) );
  AOI22_X1 U9790 ( .A1(n7721), .A2(n9061), .B1(n7427), .B2(n10920), .ZN(n7511)
         );
  NAND2_X1 U9791 ( .A1(n7512), .A2(n7511), .ZN(n10831) );
  XNOR2_X1 U9792 ( .A(n12376), .B(n10831), .ZN(n10742) );
  INV_X1 U9793 ( .A(n10742), .ZN(n8829) );
  NAND2_X1 U9794 ( .A1(n7541), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7518) );
  NAND2_X1 U9795 ( .A1(n7527), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n7517) );
  NAND2_X1 U9796 ( .A1(n7529), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n7513) );
  NAND2_X1 U9797 ( .A1(n7514), .A2(n7513), .ZN(n10808) );
  NAND2_X1 U9798 ( .A1(n7542), .A2(n10808), .ZN(n7516) );
  NAND2_X1 U9799 ( .A1(n6460), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n7515) );
  XNOR2_X1 U9800 ( .A(n10067), .B(P2_DATAO_REG_9__SCAN_IN), .ZN(n7519) );
  XNOR2_X1 U9801 ( .A(n7520), .B(n7519), .ZN(n9040) );
  OR2_X1 U9802 ( .A1(n9040), .A2(n7739), .ZN(n7526) );
  OR2_X1 U9803 ( .A1(n8759), .A2(SI_9_), .ZN(n7525) );
  OR2_X1 U9804 ( .A1(n7521), .A2(n7630), .ZN(n7523) );
  XNOR2_X1 U9805 ( .A(n7523), .B(n7522), .ZN(n14875) );
  NAND2_X1 U9806 ( .A1(n7427), .A2(n14875), .ZN(n7524) );
  INV_X1 U9807 ( .A(n10811), .ZN(n14980) );
  NAND2_X1 U9808 ( .A1(n10791), .A2(n14980), .ZN(n7565) );
  NAND2_X1 U9809 ( .A1(n10791), .A2(n10811), .ZN(n8826) );
  NAND2_X1 U9810 ( .A1(n12377), .A2(n14980), .ZN(n8827) );
  NAND2_X1 U9811 ( .A1(n7527), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n7533) );
  NAND2_X1 U9812 ( .A1(n7541), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7532) );
  NAND2_X1 U9813 ( .A1(n7545), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n7528) );
  NAND2_X1 U9814 ( .A1(n7529), .A2(n7528), .ZN(n10794) );
  NAND2_X1 U9815 ( .A1(n7542), .A2(n10794), .ZN(n7531) );
  NAND2_X1 U9816 ( .A1(n6459), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n7530) );
  XNOR2_X1 U9817 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n7534) );
  XNOR2_X1 U9818 ( .A(n7535), .B(n7534), .ZN(n9015) );
  INV_X1 U9819 ( .A(SI_8_), .ZN(n9016) );
  OR2_X1 U9820 ( .A1(n8759), .A2(n9016), .ZN(n7539) );
  NAND2_X1 U9821 ( .A1(n7536), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7537) );
  XNOR2_X1 U9822 ( .A(n7537), .B(P3_IR_REG_8__SCAN_IN), .ZN(n10908) );
  NAND2_X1 U9823 ( .A1(n7427), .A2(n10908), .ZN(n7538) );
  NAND2_X1 U9824 ( .A1(n10804), .A2(n10790), .ZN(n8769) );
  INV_X1 U9825 ( .A(n8769), .ZN(n7561) );
  NAND2_X1 U9826 ( .A1(n12378), .A2(n8821), .ZN(n8768) );
  NAND2_X1 U9827 ( .A1(n7527), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n7549) );
  NAND2_X1 U9828 ( .A1(n7541), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7548) );
  NAND2_X1 U9829 ( .A1(n7543), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7544) );
  NAND2_X1 U9830 ( .A1(n7545), .A2(n7544), .ZN(n10448) );
  NAND2_X1 U9831 ( .A1(n7542), .A2(n10448), .ZN(n7547) );
  NAND2_X1 U9832 ( .A1(n6459), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n7546) );
  AND4_X2 U9833 ( .A1(n7549), .A2(n7548), .A3(n7547), .A4(n7546), .ZN(n10789)
         );
  OR2_X1 U9834 ( .A1(n8759), .A2(SI_7_), .ZN(n7559) );
  NAND2_X1 U9835 ( .A1(n7551), .A2(n7550), .ZN(n7552) );
  AND2_X1 U9836 ( .A1(n7553), .A2(n7552), .ZN(n9012) );
  OR2_X1 U9837 ( .A1(n7739), .A2(n9012), .ZN(n7558) );
  NAND2_X1 U9838 ( .A1(n7554), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7556) );
  INV_X1 U9839 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n7555) );
  XNOR2_X1 U9840 ( .A(n7556), .B(n7555), .ZN(n14838) );
  NAND2_X1 U9841 ( .A1(n7427), .A2(n14838), .ZN(n7557) );
  NAND2_X1 U9842 ( .A1(n12379), .A2(n10447), .ZN(n10674) );
  AND2_X1 U9843 ( .A1(n8768), .A2(n10674), .ZN(n7560) );
  OR2_X1 U9844 ( .A1(n7561), .A2(n7560), .ZN(n10800) );
  AND2_X1 U9845 ( .A1(n10421), .A2(n7564), .ZN(n7563) );
  INV_X1 U9846 ( .A(n7564), .ZN(n7567) );
  NAND2_X1 U9847 ( .A1(n10789), .A2(n10447), .ZN(n8817) );
  INV_X1 U9848 ( .A(n10447), .ZN(n10429) );
  NAND2_X1 U9849 ( .A1(n12379), .A2(n10429), .ZN(n8818) );
  AND2_X1 U9850 ( .A1(n10673), .A2(n8769), .ZN(n10798) );
  AND2_X1 U9851 ( .A1(n10798), .A2(n7565), .ZN(n10738) );
  AND2_X1 U9852 ( .A1(n10738), .A2(n10742), .ZN(n7566) );
  NAND2_X1 U9853 ( .A1(n7569), .A2(n7568), .ZN(n10741) );
  INV_X1 U9854 ( .A(n10831), .ZN(n10842) );
  NAND2_X1 U9855 ( .A1(n10842), .A2(n12376), .ZN(n7570) );
  XNOR2_X1 U9856 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n7587) );
  XNOR2_X1 U9857 ( .A(n7589), .B(n7587), .ZN(n9075) );
  NAND2_X1 U9858 ( .A1(n9075), .A2(n8761), .ZN(n7577) );
  OAI21_X1 U9859 ( .B1(n7573), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7575) );
  INV_X1 U9860 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n7574) );
  XNOR2_X1 U9861 ( .A(n7575), .B(n7574), .ZN(n11086) );
  AOI22_X1 U9862 ( .A1(n7721), .A2(n9076), .B1(n7427), .B2(n11086), .ZN(n7576)
         );
  NAND2_X1 U9863 ( .A1(n7577), .A2(n7576), .ZN(n14308) );
  NAND2_X1 U9864 ( .A1(n7600), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n7583) );
  NAND2_X1 U9865 ( .A1(n6460), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n7582) );
  NAND2_X1 U9866 ( .A1(n7578), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7579) );
  NAND2_X1 U9867 ( .A1(n7598), .A2(n7579), .ZN(n14309) );
  NAND2_X1 U9868 ( .A1(n7822), .A2(n14309), .ZN(n7581) );
  NAND2_X1 U9869 ( .A1(n7541), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n7580) );
  NAND2_X1 U9870 ( .A1(n14308), .A2(n10998), .ZN(n7584) );
  NAND2_X1 U9871 ( .A1(n14302), .A2(n7584), .ZN(n7586) );
  OR2_X1 U9872 ( .A1(n14308), .A2(n10998), .ZN(n7585) );
  INV_X1 U9873 ( .A(n7587), .ZN(n7588) );
  NAND2_X1 U9874 ( .A1(n9237), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n7607) );
  NAND2_X1 U9875 ( .A1(n9202), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n7590) );
  NAND2_X1 U9876 ( .A1(n7607), .A2(n7590), .ZN(n7591) );
  NAND2_X1 U9877 ( .A1(n7592), .A2(n7591), .ZN(n7593) );
  NAND2_X1 U9878 ( .A1(n7608), .A2(n7593), .ZN(n9082) );
  NAND2_X1 U9879 ( .A1(n9082), .A2(n8761), .ZN(n7597) );
  NAND2_X1 U9880 ( .A1(n7594), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7595) );
  XNOR2_X1 U9881 ( .A(n7595), .B(n7277), .ZN(n12387) );
  AOI22_X1 U9882 ( .A1(n7721), .A2(n9083), .B1(n7427), .B2(n12387), .ZN(n7596)
         );
  NAND2_X1 U9883 ( .A1(n7597), .A2(n7596), .ZN(n11213) );
  NAND2_X1 U9884 ( .A1(n7598), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7599) );
  NAND2_X1 U9885 ( .A1(n7619), .A2(n7599), .ZN(n11216) );
  NAND2_X1 U9886 ( .A1(n7822), .A2(n11216), .ZN(n7604) );
  NAND2_X1 U9887 ( .A1(n7600), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n7603) );
  NAND2_X1 U9888 ( .A1(n6460), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n7602) );
  NAND2_X1 U9889 ( .A1(n7898), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n7601) );
  NAND4_X1 U9890 ( .A1(n7604), .A2(n7603), .A3(n7602), .A4(n7601), .ZN(n14287)
         );
  OR2_X1 U9891 ( .A1(n11213), .A2(n14287), .ZN(n8840) );
  NAND2_X1 U9892 ( .A1(n11213), .A2(n14287), .ZN(n8841) );
  NAND2_X1 U9893 ( .A1(n8840), .A2(n8841), .ZN(n10999) );
  NAND2_X1 U9894 ( .A1(n10996), .A2(n10999), .ZN(n7606) );
  INV_X1 U9895 ( .A(n14287), .ZN(n14306) );
  OR2_X1 U9896 ( .A1(n11213), .A2(n14306), .ZN(n7605) );
  NAND2_X1 U9897 ( .A1(n7609), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7628) );
  INV_X1 U9898 ( .A(n7609), .ZN(n7610) );
  NAND2_X1 U9899 ( .A1(n7610), .A2(n9253), .ZN(n7611) );
  NAND2_X1 U9900 ( .A1(n7628), .A2(n7611), .ZN(n9195) );
  OR2_X1 U9901 ( .A1(n9195), .A2(n7739), .ZN(n7615) );
  OR2_X1 U9902 ( .A1(n7612), .A2(n7630), .ZN(n7613) );
  XNOR2_X1 U9903 ( .A(n7613), .B(P3_IR_REG_13__SCAN_IN), .ZN(n12407) );
  AOI22_X1 U9904 ( .A1(n7721), .A2(SI_13_), .B1(n7427), .B2(n12407), .ZN(n7614) );
  NAND2_X1 U9905 ( .A1(n7615), .A2(n7614), .ZN(n14322) );
  NAND2_X1 U9906 ( .A1(n7541), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n7624) );
  NAND2_X1 U9907 ( .A1(n7600), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n7623) );
  INV_X1 U9908 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n7617) );
  NAND2_X1 U9909 ( .A1(n7619), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n7620) );
  NAND2_X1 U9910 ( .A1(n7634), .A2(n7620), .ZN(n14291) );
  NAND2_X1 U9911 ( .A1(n7822), .A2(n14291), .ZN(n7622) );
  NAND2_X1 U9912 ( .A1(n6459), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n7621) );
  NAND4_X1 U9913 ( .A1(n7624), .A2(n7623), .A3(n7622), .A4(n7621), .ZN(n12374)
         );
  INV_X1 U9914 ( .A(n12374), .ZN(n11420) );
  NAND2_X1 U9915 ( .A1(n14295), .A2(n11420), .ZN(n7625) );
  NAND2_X1 U9916 ( .A1(n7626), .A2(n8300), .ZN(n7627) );
  XNOR2_X1 U9917 ( .A(n8304), .B(P2_DATAO_REG_14__SCAN_IN), .ZN(n7641) );
  XNOR2_X1 U9918 ( .A(n7640), .B(n7641), .ZN(n9442) );
  NAND2_X1 U9919 ( .A1(n9442), .A2(n8761), .ZN(n7633) );
  INV_X1 U9920 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n7629) );
  AND2_X1 U9921 ( .A1(n7612), .A2(n7629), .ZN(n7646) );
  OR2_X1 U9922 ( .A1(n7646), .A2(n7630), .ZN(n7631) );
  XNOR2_X1 U9923 ( .A(n7631), .B(n7645), .ZN(n12419) );
  INV_X1 U9924 ( .A(n12419), .ZN(n12414) );
  AOI22_X1 U9925 ( .A1(n7721), .A2(SI_14_), .B1(n7427), .B2(n12414), .ZN(n7632) );
  NAND2_X1 U9926 ( .A1(n7633), .A2(n7632), .ZN(n11422) );
  NAND2_X1 U9927 ( .A1(n7898), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n7639) );
  NAND2_X1 U9928 ( .A1(n7600), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n7638) );
  NAND2_X1 U9929 ( .A1(n7634), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n7635) );
  NAND2_X1 U9930 ( .A1(n7652), .A2(n7635), .ZN(n11417) );
  NAND2_X1 U9931 ( .A1(n7822), .A2(n11417), .ZN(n7637) );
  NAND2_X1 U9932 ( .A1(n6460), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n7636) );
  OR2_X1 U9933 ( .A1(n11422), .A2(n11574), .ZN(n7925) );
  NAND2_X1 U9934 ( .A1(n11422), .A2(n11574), .ZN(n8850) );
  NAND2_X1 U9935 ( .A1(n7925), .A2(n8850), .ZN(n11251) );
  NAND2_X1 U9936 ( .A1(n11422), .A2(n14285), .ZN(n11391) );
  NAND2_X1 U9937 ( .A1(n9907), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n7660) );
  NAND2_X1 U9938 ( .A1(n9888), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n7643) );
  NAND2_X1 U9939 ( .A1(n6482), .A2(n6602), .ZN(n7644) );
  NAND2_X1 U9940 ( .A1(n7661), .A2(n7644), .ZN(n9615) );
  OR2_X1 U9941 ( .A1(n9615), .A2(n7739), .ZN(n7649) );
  NAND2_X1 U9942 ( .A1(n7646), .A2(n7645), .ZN(n7666) );
  NAND2_X1 U9943 ( .A1(n7666), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7647) );
  XNOR2_X1 U9944 ( .A(n7647), .B(P3_IR_REG_15__SCAN_IN), .ZN(n12469) );
  AOI22_X1 U9945 ( .A1(n7721), .A2(SI_15_), .B1(n7427), .B2(n12469), .ZN(n7648) );
  NAND2_X1 U9946 ( .A1(n7898), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7657) );
  NAND2_X1 U9947 ( .A1(n7600), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n7656) );
  NAND2_X1 U9948 ( .A1(n7652), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n7653) );
  NAND2_X1 U9949 ( .A1(n7670), .A2(n7653), .ZN(n11576) );
  NAND2_X1 U9950 ( .A1(n7822), .A2(n11576), .ZN(n7655) );
  NAND2_X1 U9951 ( .A1(n6460), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n7654) );
  NAND2_X1 U9952 ( .A1(n11580), .A2(n12373), .ZN(n7658) );
  AND2_X1 U9953 ( .A1(n11391), .A2(n7658), .ZN(n7659) );
  AOI21_X2 U9954 ( .B1(n11250), .B2(n7659), .A(n7338), .ZN(n11476) );
  NAND2_X1 U9955 ( .A1(n7661), .A2(n7660), .ZN(n7664) );
  NAND2_X1 U9956 ( .A1(n9725), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n7677) );
  NAND2_X1 U9957 ( .A1(n9733), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n7662) );
  OR2_X1 U9958 ( .A1(n7664), .A2(n7663), .ZN(n7665) );
  AND2_X1 U9959 ( .A1(n7665), .A2(n7678), .ZN(n9795) );
  NAND2_X1 U9960 ( .A1(n9795), .A2(n8761), .ZN(n7669) );
  NAND2_X1 U9961 ( .A1(n7680), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7667) );
  XNOR2_X1 U9962 ( .A(n7667), .B(P3_IR_REG_16__SCAN_IN), .ZN(n12478) );
  AOI22_X1 U9963 ( .A1(n7721), .A2(SI_16_), .B1(n7427), .B2(n12478), .ZN(n7668) );
  NAND2_X1 U9964 ( .A1(n7541), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n7675) );
  NAND2_X1 U9965 ( .A1(n7600), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n7674) );
  NAND2_X1 U9966 ( .A1(n7670), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n7671) );
  NAND2_X1 U9967 ( .A1(n7687), .A2(n7671), .ZN(n11611) );
  NAND2_X1 U9968 ( .A1(n7822), .A2(n11611), .ZN(n7673) );
  NAND2_X1 U9969 ( .A1(n6459), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n7672) );
  NAND2_X1 U9970 ( .A1(n11608), .A2(n12732), .ZN(n7676) );
  NAND2_X1 U9971 ( .A1(n11476), .A2(n7676), .ZN(n11474) );
  NAND2_X1 U9972 ( .A1(n12795), .A2(n12372), .ZN(n11478) );
  NAND2_X1 U9973 ( .A1(n9833), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n7699) );
  NAND2_X1 U9974 ( .A1(n9794), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n7679) );
  NAND2_X1 U9975 ( .A1(n7699), .A2(n7679), .ZN(n7696) );
  XNOR2_X1 U9976 ( .A(n7698), .B(n7696), .ZN(n9908) );
  NAND2_X1 U9977 ( .A1(n9908), .A2(n8761), .ZN(n7684) );
  OAI21_X1 U9978 ( .B1(n7680), .B2(P3_IR_REG_16__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7681) );
  MUX2_X1 U9979 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7681), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n7682) );
  NAND2_X1 U9980 ( .A1(n7682), .A2(n7718), .ZN(n12510) );
  INV_X1 U9981 ( .A(n12510), .ZN(n12501) );
  AOI22_X1 U9982 ( .A1(n7721), .A2(SI_17_), .B1(n7427), .B2(n12501), .ZN(n7683) );
  NAND2_X1 U9983 ( .A1(n7600), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n7692) );
  NAND2_X1 U9984 ( .A1(n6459), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n7691) );
  INV_X1 U9985 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n7685) );
  NAND2_X1 U9986 ( .A1(n7687), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n7688) );
  NAND2_X1 U9987 ( .A1(n7704), .A2(n7688), .ZN(n12736) );
  NAND2_X1 U9988 ( .A1(n7822), .A2(n12736), .ZN(n7690) );
  NAND2_X1 U9989 ( .A1(n7541), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n7689) );
  NAND2_X1 U9990 ( .A1(n12314), .A2(n12721), .ZN(n12714) );
  OR2_X1 U9991 ( .A1(n12314), .A2(n12721), .ZN(n7693) );
  NAND2_X1 U9992 ( .A1(n12714), .A2(n7693), .ZN(n12729) );
  NAND2_X1 U9993 ( .A1(n12730), .A2(n12729), .ZN(n7695) );
  INV_X1 U9994 ( .A(n12721), .ZN(n12371) );
  NAND2_X1 U9995 ( .A1(n12314), .A2(n12371), .ZN(n7694) );
  INV_X1 U9996 ( .A(n7696), .ZN(n7697) );
  NAND2_X1 U9997 ( .A1(n10046), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n7715) );
  INV_X1 U9998 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10044) );
  NAND2_X1 U9999 ( .A1(n10044), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n7700) );
  NAND2_X1 U10000 ( .A1(n7715), .A2(n7700), .ZN(n7712) );
  XNOR2_X1 U10001 ( .A(n7714), .B(n7712), .ZN(n9931) );
  NAND2_X1 U10002 ( .A1(n9931), .A2(n8761), .ZN(n7703) );
  NAND2_X1 U10003 ( .A1(n7718), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7701) );
  XNOR2_X1 U10004 ( .A(n7701), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12537) );
  AOI22_X1 U10005 ( .A1(n7721), .A2(SI_18_), .B1(n7427), .B2(n12537), .ZN(
        n7702) );
  NAND2_X1 U10006 ( .A1(n7541), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n7709) );
  NAND2_X1 U10007 ( .A1(n7704), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n7705) );
  NAND2_X1 U10008 ( .A1(n7725), .A2(n7705), .ZN(n12723) );
  NAND2_X1 U10009 ( .A1(n12723), .A2(n7822), .ZN(n7708) );
  NAND2_X1 U10010 ( .A1(n7600), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n7707) );
  NAND2_X1 U10011 ( .A1(n6459), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n7706) );
  NAND4_X1 U10012 ( .A1(n7709), .A2(n7708), .A3(n7707), .A4(n7706), .ZN(n12703) );
  XNOR2_X1 U10013 ( .A(n12345), .B(n12703), .ZN(n12719) );
  OR2_X1 U10014 ( .A1(n12345), .A2(n12703), .ZN(n7711) );
  INV_X1 U10015 ( .A(n7712), .ZN(n7713) );
  NAND2_X1 U10016 ( .A1(n7714), .A2(n7713), .ZN(n7716) );
  NAND2_X1 U10017 ( .A1(n10063), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n7733) );
  NAND2_X1 U10018 ( .A1(n11637), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n7717) );
  XNOR2_X1 U10019 ( .A(n7732), .B(n7731), .ZN(n9983) );
  NAND2_X1 U10020 ( .A1(n9983), .A2(n8761), .ZN(n7723) );
  INV_X1 U10021 ( .A(n7888), .ZN(n7719) );
  NAND2_X1 U10022 ( .A1(n7719), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7720) );
  AOI22_X1 U10023 ( .A1(n7721), .A2(n9982), .B1(n7427), .B2(n12543), .ZN(n7722) );
  INV_X1 U10024 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12785) );
  INV_X1 U10025 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n7724) );
  NAND2_X1 U10026 ( .A1(n7725), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n7726) );
  NAND2_X1 U10027 ( .A1(n7742), .A2(n7726), .ZN(n12708) );
  NAND2_X1 U10028 ( .A1(n12708), .A2(n7822), .ZN(n7728) );
  AOI22_X1 U10029 ( .A1(n7541), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n7600), .B2(
        P3_REG0_REG_19__SCAN_IN), .ZN(n7727) );
  OAI211_X1 U10030 ( .C1(n7901), .C2(n12785), .A(n7728), .B(n7727), .ZN(n12370) );
  OR2_X1 U10031 ( .A1(n12853), .A2(n12370), .ZN(n8876) );
  NAND2_X1 U10032 ( .A1(n12853), .A2(n12370), .ZN(n7928) );
  NAND2_X1 U10033 ( .A1(n12702), .A2(n7729), .ZN(n12701) );
  INV_X1 U10034 ( .A(n12370), .ZN(n12722) );
  OR2_X1 U10035 ( .A1(n12853), .A2(n12722), .ZN(n7730) );
  NAND2_X1 U10036 ( .A1(n7732), .A2(n7731), .ZN(n7734) );
  NAND2_X1 U10037 ( .A1(n7734), .A2(n7733), .ZN(n7735) );
  NAND2_X1 U10038 ( .A1(n7737), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7738) );
  NAND2_X1 U10039 ( .A1(n7749), .A2(n7738), .ZN(n10226) );
  OR2_X1 U10040 ( .A1(n10226), .A2(n7739), .ZN(n7741) );
  OR2_X1 U10041 ( .A1(n8759), .A2(n15098), .ZN(n7740) );
  NAND2_X1 U10042 ( .A1(n7742), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n7743) );
  NAND2_X1 U10043 ( .A1(n7755), .A2(n7743), .ZN(n12696) );
  NAND2_X1 U10044 ( .A1(n12696), .A2(n7822), .ZN(n7746) );
  AOI22_X1 U10045 ( .A1(n7541), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n7600), .B2(
        P3_REG0_REG_20__SCAN_IN), .ZN(n7745) );
  NAND2_X1 U10046 ( .A1(n6460), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n7744) );
  XNOR2_X1 U10047 ( .A(n11652), .B(n12677), .ZN(n12694) );
  NAND2_X1 U10048 ( .A1(n11652), .A2(n12704), .ZN(n7747) );
  NAND2_X1 U10049 ( .A1(n7749), .A2(n7748), .ZN(n7768) );
  INV_X1 U10050 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n10850) );
  NAND2_X1 U10051 ( .A1(n10850), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n7769) );
  INV_X1 U10052 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11635) );
  NAND2_X1 U10053 ( .A1(n11635), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n7750) );
  NAND2_X1 U10054 ( .A1(n7769), .A2(n7750), .ZN(n7766) );
  XNOR2_X1 U10055 ( .A(n7768), .B(n7766), .ZN(n10452) );
  NAND2_X1 U10056 ( .A1(n10452), .A2(n8761), .ZN(n7752) );
  INV_X1 U10057 ( .A(SI_21_), .ZN(n10453) );
  OR2_X1 U10058 ( .A1(n8759), .A2(n10453), .ZN(n7751) );
  INV_X1 U10059 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n7753) );
  NAND2_X1 U10060 ( .A1(n7755), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n7756) );
  NAND2_X1 U10061 ( .A1(n7772), .A2(n7756), .ZN(n12682) );
  NAND2_X1 U10062 ( .A1(n12682), .A2(n7822), .ZN(n7763) );
  INV_X1 U10063 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n7759) );
  NAND2_X1 U10064 ( .A1(n6459), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n7758) );
  NAND2_X1 U10065 ( .A1(n7600), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n7757) );
  OAI211_X1 U10066 ( .C1(n7760), .C2(n7759), .A(n7758), .B(n7757), .ZN(n7761)
         );
  INV_X1 U10067 ( .A(n7761), .ZN(n7762) );
  NAND2_X1 U10068 ( .A1(n12681), .A2(n12690), .ZN(n12662) );
  INV_X1 U10069 ( .A(n12690), .ZN(n12369) );
  OR2_X1 U10070 ( .A1(n12681), .A2(n12369), .ZN(n7765) );
  INV_X1 U10071 ( .A(n7766), .ZN(n7767) );
  INV_X1 U10072 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11147) );
  XNOR2_X1 U10073 ( .A(n11147), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n7782) );
  XNOR2_X1 U10074 ( .A(n7783), .B(n7782), .ZN(n10534) );
  NAND2_X1 U10075 ( .A1(n10534), .A2(n8761), .ZN(n7771) );
  INV_X1 U10076 ( .A(SI_22_), .ZN(n8538) );
  OR2_X1 U10077 ( .A1(n8759), .A2(n8538), .ZN(n7770) );
  NAND2_X1 U10078 ( .A1(n7772), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n7773) );
  NAND2_X1 U10079 ( .A1(n7786), .A2(n7773), .ZN(n12668) );
  NAND2_X1 U10080 ( .A1(n12668), .A2(n7822), .ZN(n7778) );
  INV_X1 U10081 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12772) );
  NAND2_X1 U10082 ( .A1(n7898), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n7775) );
  NAND2_X1 U10083 ( .A1(n7600), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n7774) );
  OAI211_X1 U10084 ( .C1(n12772), .C2(n7901), .A(n7775), .B(n7774), .ZN(n7776)
         );
  INV_X1 U10085 ( .A(n7776), .ZN(n7777) );
  NAND2_X1 U10086 ( .A1(n12667), .A2(n12646), .ZN(n7780) );
  NOR2_X1 U10087 ( .A1(n12667), .A2(n12646), .ZN(n7779) );
  NAND2_X1 U10088 ( .A1(n11147), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n7781) );
  XNOR2_X1 U10089 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n7795) );
  XNOR2_X1 U10090 ( .A(n7796), .B(n7795), .ZN(n10942) );
  NAND2_X1 U10091 ( .A1(n10942), .A2(n8761), .ZN(n7785) );
  OR2_X1 U10092 ( .A1(n8759), .A2(n10945), .ZN(n7784) );
  NAND2_X1 U10093 ( .A1(n7786), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n7787) );
  NAND2_X1 U10094 ( .A1(n7806), .A2(n7787), .ZN(n12651) );
  NAND2_X1 U10095 ( .A1(n12651), .A2(n7822), .ZN(n7793) );
  INV_X1 U10096 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n7790) );
  NAND2_X1 U10097 ( .A1(n7898), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n7789) );
  NAND2_X1 U10098 ( .A1(n7600), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n7788) );
  OAI211_X1 U10099 ( .C1(n7790), .C2(n7901), .A(n7789), .B(n7788), .ZN(n7791)
         );
  INV_X1 U10100 ( .A(n7791), .ZN(n7792) );
  NAND2_X1 U10101 ( .A1(n12766), .A2(n12659), .ZN(n8787) );
  NAND2_X1 U10102 ( .A1(n8891), .A2(n8787), .ZN(n12644) );
  NAND2_X1 U10103 ( .A1(n12766), .A2(n12626), .ZN(n7794) );
  INV_X1 U10104 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7797) );
  NAND2_X1 U10105 ( .A1(n7797), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7798) );
  NAND2_X1 U10106 ( .A1(n7799), .A2(n7798), .ZN(n7800) );
  INV_X1 U10107 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11979) );
  NAND2_X1 U10108 ( .A1(n7800), .A2(n11979), .ZN(n7801) );
  XNOR2_X1 U10109 ( .A(n7812), .B(n11273), .ZN(n11222) );
  NAND2_X1 U10110 ( .A1(n11222), .A2(n8761), .ZN(n7803) );
  INV_X1 U10111 ( .A(SI_24_), .ZN(n11223) );
  OR2_X1 U10112 ( .A1(n8759), .A2(n11223), .ZN(n7802) );
  INV_X1 U10113 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n7804) );
  NAND2_X1 U10114 ( .A1(n7806), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n7807) );
  NAND2_X1 U10115 ( .A1(n7820), .A2(n7807), .ZN(n12635) );
  INV_X1 U10116 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12764) );
  NAND2_X1 U10117 ( .A1(n7600), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n7809) );
  NAND2_X1 U10118 ( .A1(n7898), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n7808) );
  OAI211_X1 U10119 ( .C1(n7901), .C2(n12764), .A(n7809), .B(n7808), .ZN(n7810)
         );
  AOI21_X1 U10120 ( .B1(n12635), .B2(n7822), .A(n7810), .ZN(n12285) );
  XNOR2_X1 U10121 ( .A(n12634), .B(n12285), .ZN(n12629) );
  NAND2_X1 U10122 ( .A1(n12634), .A2(n12647), .ZN(n7811) );
  NAND2_X1 U10123 ( .A1(n7814), .A2(n7813), .ZN(n7830) );
  XNOR2_X1 U10124 ( .A(n11377), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n7815) );
  XNOR2_X1 U10125 ( .A(n7830), .B(n7815), .ZN(n11339) );
  NAND2_X1 U10126 ( .A1(n11339), .A2(n8761), .ZN(n7817) );
  OR2_X1 U10127 ( .A1(n8759), .A2(n11341), .ZN(n7816) );
  INV_X1 U10128 ( .A(n7820), .ZN(n7819) );
  INV_X1 U10129 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n7818) );
  NAND2_X1 U10130 ( .A1(n7820), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n7821) );
  NAND2_X1 U10131 ( .A1(n7836), .A2(n7821), .ZN(n12618) );
  NAND2_X1 U10132 ( .A1(n12618), .A2(n7822), .ZN(n7827) );
  INV_X1 U10133 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n12760) );
  NAND2_X1 U10134 ( .A1(n7898), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n7824) );
  NAND2_X1 U10135 ( .A1(n7600), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n7823) );
  OAI211_X1 U10136 ( .C1(n12760), .C2(n7901), .A(n7824), .B(n7823), .ZN(n7825)
         );
  INV_X1 U10137 ( .A(n7825), .ZN(n7826) );
  XNOR2_X1 U10138 ( .A(n12311), .B(n12362), .ZN(n12612) );
  NAND2_X1 U10139 ( .A1(n12613), .A2(n12612), .ZN(n12611) );
  NAND2_X1 U10140 ( .A1(n12311), .A2(n12627), .ZN(n7828) );
  NAND2_X1 U10141 ( .A1(n11377), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n7829) );
  NAND2_X1 U10142 ( .A1(n7830), .A2(n7829), .ZN(n7832) );
  NAND2_X1 U10143 ( .A1(n11374), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n7831) );
  NAND2_X1 U10144 ( .A1(n7832), .A2(n7831), .ZN(n7845) );
  INV_X1 U10145 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n11488) );
  XNOR2_X1 U10146 ( .A(n11488), .B(P2_DATAO_REG_26__SCAN_IN), .ZN(n7833) );
  XNOR2_X1 U10147 ( .A(n7845), .B(n7833), .ZN(n11402) );
  NAND2_X1 U10148 ( .A1(n11402), .A2(n8761), .ZN(n7835) );
  OR2_X1 U10149 ( .A1(n8759), .A2(n11404), .ZN(n7834) );
  NAND2_X1 U10150 ( .A1(n7836), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n7837) );
  NAND2_X1 U10151 ( .A1(n7852), .A2(n7837), .ZN(n12603) );
  NAND2_X1 U10152 ( .A1(n12603), .A2(n7542), .ZN(n7842) );
  INV_X1 U10153 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12756) );
  NAND2_X1 U10154 ( .A1(n7541), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n7839) );
  NAND2_X1 U10155 ( .A1(n7600), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n7838) );
  OAI211_X1 U10156 ( .C1(n12756), .C2(n7901), .A(n7839), .B(n7838), .ZN(n7840)
         );
  INV_X1 U10157 ( .A(n7840), .ZN(n7841) );
  OR2_X1 U10158 ( .A1(n12752), .A2(n12614), .ZN(n7843) );
  INV_X1 U10159 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n11513) );
  AND2_X1 U10160 ( .A1(n11513), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n7844) );
  NAND2_X1 U10161 ( .A1(n11488), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n7846) );
  XNOR2_X1 U10162 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n7847) );
  XNOR2_X1 U10163 ( .A(n7862), .B(n7847), .ZN(n12882) );
  NAND2_X1 U10164 ( .A1(n12882), .A2(n8761), .ZN(n7849) );
  OR2_X1 U10165 ( .A1(n8759), .A2(n12884), .ZN(n7848) );
  INV_X1 U10166 ( .A(n7852), .ZN(n7851) );
  INV_X1 U10167 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n7850) );
  NAND2_X1 U10168 ( .A1(n7851), .A2(n7850), .ZN(n7866) );
  NAND2_X1 U10169 ( .A1(n7852), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n7853) );
  NAND2_X1 U10170 ( .A1(n7866), .A2(n7853), .ZN(n12589) );
  NAND2_X1 U10171 ( .A1(n12589), .A2(n7542), .ZN(n7858) );
  INV_X1 U10172 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n12750) );
  NAND2_X1 U10173 ( .A1(n7600), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n7855) );
  NAND2_X1 U10174 ( .A1(n7898), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n7854) );
  OAI211_X1 U10175 ( .C1(n12750), .C2(n7901), .A(n7855), .B(n7854), .ZN(n7856)
         );
  INV_X1 U10176 ( .A(n7856), .ZN(n7857) );
  XNOR2_X1 U10177 ( .A(n11677), .B(n12600), .ZN(n8779) );
  NAND2_X1 U10178 ( .A1(n12583), .A2(n7859), .ZN(n12582) );
  OR2_X1 U10179 ( .A1(n11677), .A2(n12600), .ZN(n7860) );
  NAND2_X1 U10180 ( .A1(n12582), .A2(n7860), .ZN(n12563) );
  INV_X1 U10181 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13524) );
  AND2_X1 U10182 ( .A1(n13524), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n7861) );
  INV_X1 U10183 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14134) );
  INV_X1 U10184 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n15043) );
  XNOR2_X1 U10185 ( .A(n15043), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n7863) );
  NAND2_X1 U10186 ( .A1(n12878), .A2(n8761), .ZN(n7865) );
  INV_X1 U10187 ( .A(SI_28_), .ZN(n12881) );
  OR2_X1 U10188 ( .A1(n8759), .A2(n12881), .ZN(n7864) );
  NAND2_X1 U10189 ( .A1(n7866), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n7867) );
  NAND2_X1 U10190 ( .A1(n11631), .A2(n7867), .ZN(n12577) );
  NAND2_X1 U10191 ( .A1(n12577), .A2(n7542), .ZN(n7872) );
  INV_X1 U10192 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n12747) );
  NAND2_X1 U10193 ( .A1(n7600), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n7869) );
  NAND2_X1 U10194 ( .A1(n7541), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n7868) );
  OAI211_X1 U10195 ( .C1(n7901), .C2(n12747), .A(n7869), .B(n7868), .ZN(n7870)
         );
  INV_X1 U10196 ( .A(n7870), .ZN(n7871) );
  NAND2_X1 U10197 ( .A1(n12824), .A2(n12585), .ZN(n8910) );
  NAND2_X1 U10198 ( .A1(n11704), .A2(n12555), .ZN(n7937) );
  INV_X1 U10199 ( .A(n7874), .ZN(n7876) );
  INV_X1 U10200 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n11683) );
  NAND2_X1 U10201 ( .A1(n11683), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n7875) );
  NAND2_X1 U10202 ( .A1(n7876), .A2(n7875), .ZN(n7878) );
  NAND2_X1 U10203 ( .A1(n15043), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n7877) );
  XNOR2_X1 U10204 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n8745) );
  XNOR2_X1 U10205 ( .A(n8747), .B(n8745), .ZN(n12156) );
  NAND2_X1 U10206 ( .A1(n12156), .A2(n8761), .ZN(n7880) );
  INV_X1 U10207 ( .A(SI_29_), .ZN(n12159) );
  OR2_X1 U10208 ( .A1(n8759), .A2(n12159), .ZN(n7879) );
  INV_X1 U10209 ( .A(n11631), .ZN(n7881) );
  NAND2_X1 U10210 ( .A1(n7881), .A2(n7542), .ZN(n8756) );
  INV_X1 U10211 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n8960) );
  NAND2_X1 U10212 ( .A1(n7600), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n7883) );
  NAND2_X1 U10213 ( .A1(n7898), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n7882) );
  OAI211_X1 U10214 ( .C1(n7901), .C2(n8960), .A(n7883), .B(n7882), .ZN(n7884)
         );
  INV_X1 U10215 ( .A(n7884), .ZN(n7885) );
  NAND2_X1 U10216 ( .A1(n7985), .A2(n12568), .ZN(n8927) );
  NAND2_X1 U10217 ( .A1(n8925), .A2(n8927), .ZN(n8908) );
  XNOR2_X1 U10218 ( .A(n7886), .B(n8908), .ZN(n12552) );
  NAND2_X1 U10219 ( .A1(n7971), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7890) );
  NAND2_X1 U10220 ( .A1(n10535), .A2(n12533), .ZN(n7978) );
  XNOR2_X2 U10221 ( .A(n7891), .B(P3_IR_REG_21__SCAN_IN), .ZN(n10140) );
  INV_X1 U10222 ( .A(n7892), .ZN(n7893) );
  NAND2_X1 U10223 ( .A1(n7893), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7894) );
  MUX2_X1 U10224 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7894), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n7896) );
  NAND2_X1 U10225 ( .A1(n7896), .A2(n7895), .ZN(n10225) );
  INV_X1 U10226 ( .A(n10225), .ZN(n7976) );
  NAND2_X1 U10227 ( .A1(n10140), .A2(n7976), .ZN(n8937) );
  INV_X1 U10228 ( .A(n12880), .ZN(n9531) );
  INV_X1 U10229 ( .A(n6446), .ZN(n8942) );
  NAND2_X1 U10230 ( .A1(n9531), .A2(n8942), .ZN(n9543) );
  NAND2_X1 U10231 ( .A1(n9543), .A2(n9530), .ZN(n9757) );
  INV_X1 U10232 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n7902) );
  NAND2_X1 U10233 ( .A1(n7541), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n7900) );
  NAND2_X1 U10234 ( .A1(n7600), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n7899) );
  OAI211_X1 U10235 ( .C1(n7902), .C2(n7901), .A(n7900), .B(n7899), .ZN(n7903)
         );
  INV_X1 U10236 ( .A(n7903), .ZN(n7904) );
  INV_X1 U10237 ( .A(P3_B_REG_SCAN_IN), .ZN(n7905) );
  NOR2_X1 U10238 ( .A1(n12880), .A2(n7905), .ZN(n7906) );
  OR2_X1 U10239 ( .A1(n14917), .A2(n7906), .ZN(n12554) );
  OAI21_X1 U10240 ( .B1(n12552), .B2(n14303), .A(n7909), .ZN(n7945) );
  INV_X1 U10241 ( .A(n7910), .ZN(n7911) );
  OR2_X1 U10242 ( .A1(n8763), .A2(n9893), .ZN(n9750) );
  NAND2_X1 U10243 ( .A1(n9750), .A2(n8789), .ZN(n8788) );
  AND2_X1 U10244 ( .A1(n10230), .A2(n8808), .ZN(n10513) );
  AND2_X1 U10245 ( .A1(n10513), .A2(n10522), .ZN(n7916) );
  INV_X1 U10246 ( .A(n10522), .ZN(n7915) );
  INV_X1 U10247 ( .A(n8808), .ZN(n7914) );
  AND2_X1 U10248 ( .A1(n10213), .A2(n8810), .ZN(n7913) );
  OR2_X1 U10249 ( .A1(n7914), .A2(n7913), .ZN(n10515) );
  NAND2_X1 U10250 ( .A1(n10422), .A2(n10423), .ZN(n7917) );
  INV_X1 U10251 ( .A(n10673), .ZN(n8765) );
  NAND2_X1 U10252 ( .A1(n7917), .A2(n8765), .ZN(n10425) );
  NAND2_X1 U10253 ( .A1(n10425), .A2(n8817), .ZN(n10677) );
  NAND2_X1 U10254 ( .A1(n12378), .A2(n10790), .ZN(n7918) );
  NAND2_X1 U10255 ( .A1(n10677), .A2(n7918), .ZN(n7920) );
  NAND2_X1 U10256 ( .A1(n10804), .A2(n8821), .ZN(n7919) );
  NAND2_X1 U10257 ( .A1(n7920), .A2(n7919), .ZN(n10797) );
  NAND2_X1 U10258 ( .A1(n10797), .A2(n10802), .ZN(n7921) );
  NAND2_X1 U10259 ( .A1(n7921), .A2(n8826), .ZN(n10737) );
  NAND2_X1 U10260 ( .A1(n10737), .A2(n8829), .ZN(n7923) );
  INV_X1 U10261 ( .A(n12376), .ZN(n14305) );
  NAND2_X1 U10262 ( .A1(n14305), .A2(n10842), .ZN(n7922) );
  NAND2_X1 U10263 ( .A1(n7923), .A2(n7922), .ZN(n14300) );
  NOR2_X1 U10264 ( .A1(n14308), .A2(n12375), .ZN(n8836) );
  NAND2_X1 U10265 ( .A1(n14308), .A2(n12375), .ZN(n8835) );
  AND2_X1 U10266 ( .A1(n14322), .A2(n11420), .ZN(n8847) );
  NAND2_X1 U10267 ( .A1(n14295), .A2(n12374), .ZN(n8845) );
  INV_X1 U10268 ( .A(n7925), .ZN(n8853) );
  NAND2_X1 U10269 ( .A1(n12865), .A2(n12373), .ZN(n8852) );
  NAND2_X1 U10270 ( .A1(n11580), .A2(n11601), .ZN(n8860) );
  NAND2_X1 U10271 ( .A1(n11397), .A2(n11396), .ZN(n11395) );
  NAND2_X1 U10272 ( .A1(n11395), .A2(n8860), .ZN(n11484) );
  NAND2_X1 U10273 ( .A1(n11608), .A2(n12372), .ZN(n8862) );
  NAND2_X1 U10274 ( .A1(n12795), .A2(n12732), .ZN(n8861) );
  NAND2_X1 U10275 ( .A1(n11484), .A2(n11483), .ZN(n11482) );
  NAND2_X1 U10276 ( .A1(n11482), .A2(n8861), .ZN(n12735) );
  INV_X1 U10277 ( .A(n12729), .ZN(n12734) );
  INV_X1 U10278 ( .A(n12703), .ZN(n12733) );
  NAND2_X1 U10279 ( .A1(n12345), .A2(n12733), .ZN(n7926) );
  AND2_X1 U10280 ( .A1(n7926), .A2(n12714), .ZN(n8867) );
  NAND2_X1 U10281 ( .A1(n12713), .A2(n8867), .ZN(n7927) );
  OR2_X1 U10282 ( .A1(n12345), .A2(n12733), .ZN(n8865) );
  INV_X1 U10283 ( .A(n7928), .ZN(n8877) );
  NAND2_X1 U10284 ( .A1(n12780), .A2(n12704), .ZN(n12661) );
  AND2_X1 U10285 ( .A1(n12663), .A2(n8885), .ZN(n7931) );
  AND2_X1 U10286 ( .A1(n12661), .A2(n7931), .ZN(n7933) );
  INV_X1 U10287 ( .A(n12662), .ZN(n7930) );
  NAND2_X1 U10288 ( .A1(n12667), .A2(n12678), .ZN(n8886) );
  INV_X1 U10289 ( .A(n12644), .ZN(n12641) );
  NAND2_X1 U10290 ( .A1(n12642), .A2(n12641), .ZN(n12640) );
  NAND2_X1 U10291 ( .A1(n12634), .A2(n12285), .ZN(n8892) );
  INV_X1 U10292 ( .A(n12612), .ZN(n8895) );
  NAND2_X1 U10293 ( .A1(n12311), .A2(n12362), .ZN(n8899) );
  NAND2_X1 U10294 ( .A1(n12752), .A2(n12309), .ZN(n8903) );
  NAND2_X1 U10295 ( .A1(n8902), .A2(n8903), .ZN(n12594) );
  NAND2_X1 U10296 ( .A1(n12597), .A2(n8902), .ZN(n12581) );
  NOR2_X1 U10297 ( .A1(n12581), .A2(n7859), .ZN(n12572) );
  NAND2_X1 U10298 ( .A1(n11677), .A2(n12567), .ZN(n12573) );
  NAND2_X1 U10299 ( .A1(n7937), .A2(n12573), .ZN(n8909) );
  XNOR2_X1 U10300 ( .A(n8931), .B(n8908), .ZN(n12551) );
  AND2_X1 U10301 ( .A1(n7977), .A2(n10225), .ZN(n8951) );
  INV_X1 U10302 ( .A(n8951), .ZN(n7938) );
  XNOR2_X1 U10303 ( .A(n10535), .B(n7938), .ZN(n7940) );
  NAND2_X1 U10304 ( .A1(n7977), .A2(n12543), .ZN(n7939) );
  NAND2_X1 U10305 ( .A1(n7940), .A2(n7939), .ZN(n9291) );
  INV_X1 U10306 ( .A(n10535), .ZN(n7943) );
  INV_X1 U10307 ( .A(n9755), .ZN(n8947) );
  AND2_X1 U10308 ( .A1(n14979), .A2(n8947), .ZN(n7941) );
  NAND2_X1 U10309 ( .A1(n9291), .A2(n7941), .ZN(n7942) );
  NAND2_X1 U10310 ( .A1(n7978), .A2(n9755), .ZN(n8949) );
  NAND2_X1 U10311 ( .A1(n10225), .A2(n12533), .ZN(n14936) );
  MUX2_X1 U10312 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7946), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n7948) );
  INV_X1 U10313 ( .A(n7947), .ZN(n7949) );
  XNOR2_X1 U10314 ( .A(n11225), .B(P3_B_REG_SCAN_IN), .ZN(n7953) );
  NAND2_X1 U10315 ( .A1(n7949), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7950) );
  MUX2_X1 U10316 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7950), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n7952) );
  NAND2_X1 U10317 ( .A1(n7952), .A2(n7951), .ZN(n11340) );
  NAND2_X1 U10318 ( .A1(n7953), .A2(n11340), .ZN(n7955) );
  NAND2_X1 U10319 ( .A1(n7951), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7954) );
  INV_X1 U10320 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n7956) );
  INV_X1 U10321 ( .A(n7975), .ZN(n11403) );
  NAND2_X1 U10322 ( .A1(n11403), .A2(n11225), .ZN(n7957) );
  INV_X1 U10323 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n7958) );
  NAND2_X1 U10324 ( .A1(n9089), .A2(n7958), .ZN(n7960) );
  NAND2_X1 U10325 ( .A1(n11403), .A2(n11340), .ZN(n7959) );
  INV_X1 U10326 ( .A(n10031), .ZN(n12866) );
  NAND2_X1 U10327 ( .A1(n12868), .A2(n12866), .ZN(n8957) );
  NOR2_X1 U10328 ( .A1(P3_D_REG_23__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .ZN(
        n7964) );
  NOR4_X1 U10329 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n7963) );
  NOR4_X1 U10330 ( .A1(P3_D_REG_25__SCAN_IN), .A2(P3_D_REG_20__SCAN_IN), .A3(
        P3_D_REG_19__SCAN_IN), .A4(P3_D_REG_18__SCAN_IN), .ZN(n7962) );
  NOR4_X1 U10331 ( .A1(P3_D_REG_24__SCAN_IN), .A2(P3_D_REG_15__SCAN_IN), .A3(
        P3_D_REG_22__SCAN_IN), .A4(P3_D_REG_17__SCAN_IN), .ZN(n7961) );
  NAND4_X1 U10332 ( .A1(n7964), .A2(n7963), .A3(n7962), .A4(n7961), .ZN(n7970)
         );
  NOR4_X1 U10333 ( .A1(P3_D_REG_14__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_11__SCAN_IN), .A4(P3_D_REG_9__SCAN_IN), .ZN(n7968) );
  NOR4_X1 U10334 ( .A1(P3_D_REG_10__SCAN_IN), .A2(P3_D_REG_27__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_31__SCAN_IN), .ZN(n7967) );
  NOR4_X1 U10335 ( .A1(P3_D_REG_6__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n7966) );
  NOR4_X1 U10336 ( .A1(P3_D_REG_16__SCAN_IN), .A2(P3_D_REG_30__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n7965) );
  NAND4_X1 U10337 ( .A1(n7968), .A2(n7967), .A3(n7966), .A4(n7965), .ZN(n7969)
         );
  OAI21_X1 U10338 ( .B1(n7970), .B2(n7969), .A(n9089), .ZN(n8956) );
  INV_X1 U10339 ( .A(n8956), .ZN(n7982) );
  NOR2_X1 U10340 ( .A1(n8957), .A2(n7982), .ZN(n9298) );
  NOR2_X1 U10341 ( .A1(n11340), .A2(n11225), .ZN(n7974) );
  NAND2_X1 U10342 ( .A1(n7975), .A2(n7974), .ZN(n9292) );
  NOR2_X1 U10343 ( .A1(n8948), .A2(n9755), .ZN(n9517) );
  NAND2_X1 U10344 ( .A1(n9526), .A2(n9517), .ZN(n9300) );
  NOR2_X1 U10345 ( .A1(n7978), .A2(n6991), .ZN(n9293) );
  NAND2_X1 U10346 ( .A1(n9526), .A2(n9293), .ZN(n7979) );
  NAND2_X1 U10347 ( .A1(n9300), .A2(n7979), .ZN(n7980) );
  NAND2_X1 U10348 ( .A1(n9298), .A2(n7980), .ZN(n7984) );
  INV_X1 U10349 ( .A(n12868), .ZN(n7981) );
  NAND2_X1 U10350 ( .A1(n7981), .A2(n10031), .ZN(n8955) );
  NAND3_X1 U10351 ( .A1(n9301), .A2(n9526), .A3(n9291), .ZN(n7983) );
  INV_X1 U10352 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n7986) );
  INV_X1 U10354 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n7994) );
  NOR2_X1 U10355 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n7997) );
  NOR2_X1 U10356 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), 
        .ZN(n7996) );
  NOR2_X1 U10357 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), 
        .ZN(n8000) );
  NAND2_X1 U10358 ( .A1(n8003), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8004) );
  NAND2_X2 U10359 ( .A1(n12131), .A2(n8007), .ZN(n8118) );
  NAND2_X1 U10360 ( .A1(n8085), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n8011) );
  NAND2_X1 U10361 ( .A1(n8116), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n8010) );
  NOR2_X2 U10362 ( .A1(n12131), .A2(n8006), .ZN(n8117) );
  NAND2_X1 U10363 ( .A1(n8117), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n8009) );
  NAND2_X1 U10364 ( .A1(n6457), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n8008) );
  INV_X1 U10365 ( .A(SI_0_), .ZN(n8012) );
  NOR2_X1 U10366 ( .A1(n9335), .A2(n8012), .ZN(n8014) );
  XNOR2_X1 U10367 ( .A(n8014), .B(n8013), .ZN(n14138) );
  MUX2_X1 U10368 ( .A(P1_IR_REG_0__SCAN_IN), .B(n14138), .S(n9084), .Z(n9840)
         );
  INV_X1 U10369 ( .A(n10276), .ZN(n8034) );
  NAND2_X1 U10370 ( .A1(n6457), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n8022) );
  NAND2_X1 U10371 ( .A1(n8085), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n8020) );
  NAND2_X1 U10372 ( .A1(n8116), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n8019) );
  NAND2_X1 U10373 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n8023) );
  MUX2_X1 U10374 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8023), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n8026) );
  INV_X1 U10375 ( .A(n8024), .ZN(n8025) );
  NAND2_X1 U10376 ( .A1(n8026), .A2(n8025), .ZN(n9212) );
  OR2_X1 U10377 ( .A1(n9084), .A2(n9212), .ZN(n8033) );
  INV_X1 U10378 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n8996) );
  OR2_X1 U10379 ( .A1(n8113), .A2(n8996), .ZN(n8032) );
  NAND2_X1 U10380 ( .A1(n8027), .A2(n9050), .ZN(n8029) );
  NAND2_X1 U10381 ( .A1(n8028), .A2(SI_1_), .ZN(n8072) );
  NAND2_X1 U10382 ( .A1(n8029), .A2(n8072), .ZN(n8074) );
  MUX2_X1 U10383 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(P1_DATAO_REG_0__SCAN_IN), 
        .S(n8111), .Z(n8030) );
  NAND2_X1 U10384 ( .A1(n8030), .A2(SI_0_), .ZN(n8073) );
  XNOR2_X1 U10385 ( .A(n8074), .B(n8073), .ZN(n9374) );
  OR2_X1 U10386 ( .A1(n8094), .A2(n9374), .ZN(n8031) );
  NAND2_X1 U10387 ( .A1(n9279), .A2(n11693), .ZN(n10278) );
  AND2_X1 U10388 ( .A1(n8034), .A2(n10278), .ZN(n8054) );
  INV_X1 U10389 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n8035) );
  NAND2_X1 U10390 ( .A1(n8413), .A2(n8035), .ZN(n8428) );
  MUX2_X1 U10391 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8036), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n8039) );
  NAND2_X1 U10392 ( .A1(n8041), .A2(n8040), .ZN(n8047) );
  INV_X1 U10393 ( .A(n8047), .ZN(n8043) );
  NAND2_X2 U10394 ( .A1(n8045), .A2(n8726), .ZN(n9824) );
  NAND2_X1 U10395 ( .A1(n8730), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8046) );
  OR2_X1 U10396 ( .A1(n8052), .A2(n10586), .ZN(n8053) );
  NAND2_X1 U10397 ( .A1(n8047), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8049) );
  MUX2_X1 U10398 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8049), .S(
        P1_IR_REG_21__SCAN_IN), .Z(n8051) );
  INV_X1 U10399 ( .A(n9273), .ZN(n10849) );
  NAND2_X1 U10400 ( .A1(n8052), .A2(n10849), .ZN(n8644) );
  NAND2_X1 U10401 ( .A1(n10276), .A2(n9416), .ZN(n8055) );
  INV_X1 U10402 ( .A(n9695), .ZN(n13680) );
  NAND2_X1 U10403 ( .A1(n13680), .A2(n10439), .ZN(n8690) );
  NAND2_X1 U10404 ( .A1(n8116), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n8065) );
  NAND2_X1 U10405 ( .A1(n8117), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n8064) );
  NAND2_X1 U10406 ( .A1(n6457), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n8063) );
  INV_X1 U10407 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n8061) );
  NAND2_X1 U10408 ( .A1(n8613), .A2(n8061), .ZN(n8062) );
  INV_X1 U10409 ( .A(n9817), .ZN(n13677) );
  OR2_X1 U10410 ( .A1(n8113), .A2(n8995), .ZN(n8071) );
  NAND2_X1 U10411 ( .A1(n8066), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8067) );
  MUX2_X1 U10412 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8067), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n8070) );
  NAND2_X1 U10413 ( .A1(n8070), .A2(n8069), .ZN(n13712) );
  MUX2_X1 U10414 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n8111), .Z(n8075) );
  OAI21_X1 U10415 ( .B1(n8075), .B2(SI_2_), .A(n8077), .ZN(n8076) );
  INV_X1 U10416 ( .A(n8076), .ZN(n8092) );
  MUX2_X1 U10417 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n8111), .Z(n8078) );
  OAI21_X1 U10418 ( .B1(n8078), .B2(SI_3_), .A(n8109), .ZN(n8079) );
  INV_X1 U10419 ( .A(n8079), .ZN(n8080) );
  OR2_X1 U10420 ( .A1(n8081), .A2(n8080), .ZN(n8082) );
  NAND2_X1 U10421 ( .A1(n8110), .A2(n8082), .ZN(n9643) );
  MUX2_X1 U10422 ( .A(n10278), .B(n10277), .S(n6453), .Z(n8100) );
  NAND2_X1 U10423 ( .A1(n8116), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n8089) );
  NAND2_X1 U10424 ( .A1(n6457), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n8088) );
  NAND2_X1 U10425 ( .A1(n8117), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n8087) );
  NAND2_X1 U10426 ( .A1(n8085), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n8086) );
  OAI21_X1 U10427 ( .B1(n8093), .B2(n8092), .A(n8091), .ZN(n9395) );
  OR2_X1 U10428 ( .A1(n8094), .A2(n9395), .ZN(n8095) );
  NAND2_X1 U10429 ( .A1(n8691), .A2(n10463), .ZN(n10280) );
  NAND2_X1 U10430 ( .A1(n10280), .A2(n6454), .ZN(n8098) );
  NAND2_X1 U10431 ( .A1(n13678), .A2(n14504), .ZN(n8103) );
  NAND2_X1 U10432 ( .A1(n8103), .A2(n6451), .ZN(n8097) );
  NAND2_X1 U10433 ( .A1(n8098), .A2(n8097), .ZN(n8099) );
  NAND3_X1 U10434 ( .A1(n10291), .A2(n8100), .A3(n8099), .ZN(n8107) );
  MUX2_X1 U10435 ( .A(n8101), .B(n10281), .S(n6447), .Z(n8106) );
  INV_X1 U10436 ( .A(n10280), .ZN(n8102) );
  NAND3_X1 U10437 ( .A1(n8102), .A2(n6451), .A3(n8101), .ZN(n8105) );
  NAND2_X1 U10438 ( .A1(n8069), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8108) );
  XNOR2_X1 U10439 ( .A(n8108), .B(n6959), .ZN(n9219) );
  MUX2_X1 U10440 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n8111), .Z(n8112) );
  NAND2_X1 U10441 ( .A1(n8112), .A2(SI_4_), .ZN(n8142) );
  OAI21_X1 U10442 ( .B1(n8112), .B2(SI_4_), .A(n8142), .ZN(n8139) );
  XNOR2_X1 U10443 ( .A(n8141), .B(n8139), .ZN(n9648) );
  OR2_X1 U10444 ( .A1(n8681), .A2(n9005), .ZN(n8114) );
  OAI211_X1 U10445 ( .C1(n9084), .C2(n9219), .A(n8115), .B(n8114), .ZN(n14521)
         );
  NAND2_X1 U10446 ( .A1(n8612), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n8124) );
  CLKBUF_X3 U10447 ( .A(n8117), .Z(n8624) );
  NAND2_X1 U10448 ( .A1(n8624), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n8123) );
  INV_X2 U10449 ( .A(n8118), .ZN(n8613) );
  NOR2_X1 U10450 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n8119) );
  NOR2_X1 U10451 ( .A1(n8133), .A2(n8119), .ZN(n10616) );
  NAND2_X1 U10452 ( .A1(n8613), .A2(n10616), .ZN(n8122) );
  INV_X2 U10453 ( .A(n8630), .ZN(n8625) );
  NAND2_X1 U10454 ( .A1(n8625), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n8121) );
  MUX2_X1 U10455 ( .A(n14521), .B(n13676), .S(n6453), .Z(n8128) );
  NAND2_X1 U10456 ( .A1(n8127), .A2(n8128), .ZN(n8126) );
  MUX2_X1 U10457 ( .A(n13676), .B(n14521), .S(n6454), .Z(n8125) );
  NAND2_X1 U10458 ( .A1(n8126), .A2(n8125), .ZN(n8132) );
  INV_X1 U10459 ( .A(n8127), .ZN(n8130) );
  INV_X1 U10460 ( .A(n8128), .ZN(n8129) );
  NAND2_X1 U10461 ( .A1(n8130), .A2(n8129), .ZN(n8131) );
  NAND2_X1 U10462 ( .A1(n8625), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n8138) );
  NAND2_X1 U10463 ( .A1(n8612), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n8137) );
  NAND2_X1 U10464 ( .A1(n8133), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n8178) );
  OAI21_X1 U10465 ( .B1(n8133), .B2(P1_REG3_REG_5__SCAN_IN), .A(n8178), .ZN(
        n8134) );
  INV_X1 U10466 ( .A(n8134), .ZN(n14465) );
  NAND2_X1 U10467 ( .A1(n8647), .A2(n14465), .ZN(n8136) );
  NAND2_X1 U10468 ( .A1(n8624), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n8135) );
  INV_X1 U10469 ( .A(n8139), .ZN(n8140) );
  NAND2_X1 U10470 ( .A1(n8143), .A2(n8142), .ZN(n8153) );
  MUX2_X1 U10471 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n9335), .Z(n8144) );
  NAND2_X1 U10472 ( .A1(n8144), .A2(SI_5_), .ZN(n8154) );
  OAI21_X1 U10473 ( .B1(n8144), .B2(SI_5_), .A(n8154), .ZN(n8151) );
  XNOR2_X1 U10474 ( .A(n8153), .B(n8151), .ZN(n9621) );
  OR2_X1 U10475 ( .A1(n8145), .A2(n14125), .ZN(n8146) );
  XNOR2_X1 U10476 ( .A(n8146), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9222) );
  AOI22_X1 U10477 ( .A1(n6455), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n8444), .B2(
        n9222), .ZN(n8147) );
  NAND2_X1 U10478 ( .A1(n8148), .A2(n8147), .ZN(n14467) );
  MUX2_X1 U10479 ( .A(n13674), .B(n14467), .S(n6453), .Z(n8150) );
  MUX2_X1 U10480 ( .A(n13674), .B(n14467), .S(n6451), .Z(n8149) );
  INV_X1 U10481 ( .A(n8151), .ZN(n8152) );
  NAND2_X1 U10482 ( .A1(n8153), .A2(n8152), .ZN(n8155) );
  INV_X1 U10483 ( .A(n8156), .ZN(n8157) );
  OR2_X1 U10484 ( .A1(n8158), .A2(n8157), .ZN(n8159) );
  NAND2_X1 U10485 ( .A1(n8186), .A2(n8159), .ZN(n9847) );
  OR2_X1 U10486 ( .A1(n9847), .A2(n8266), .ZN(n8163) );
  INV_X1 U10487 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n8160) );
  NAND2_X1 U10488 ( .A1(n8145), .A2(n8160), .ZN(n8192) );
  NAND2_X1 U10489 ( .A1(n8192), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8161) );
  XNOR2_X1 U10490 ( .A(n8161), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9467) );
  AOI22_X1 U10491 ( .A1(n6455), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n8444), .B2(
        n9467), .ZN(n8162) );
  NAND2_X1 U10492 ( .A1(n8163), .A2(n8162), .ZN(n10596) );
  NAND2_X1 U10493 ( .A1(n8625), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n8167) );
  NAND2_X1 U10494 ( .A1(n8612), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n8166) );
  XNOR2_X1 U10495 ( .A(n8178), .B(P1_REG3_REG_6__SCAN_IN), .ZN(n13624) );
  NAND2_X1 U10496 ( .A1(n8613), .A2(n13624), .ZN(n8165) );
  NAND2_X1 U10497 ( .A1(n8624), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n8164) );
  NAND4_X1 U10498 ( .A1(n8167), .A2(n8166), .A3(n8165), .A4(n8164), .ZN(n13673) );
  MUX2_X1 U10499 ( .A(n10596), .B(n13673), .S(n6453), .Z(n8171) );
  NAND2_X1 U10500 ( .A1(n8170), .A2(n8171), .ZN(n8169) );
  MUX2_X1 U10501 ( .A(n10596), .B(n13673), .S(n6447), .Z(n8168) );
  NAND2_X1 U10502 ( .A1(n8169), .A2(n8168), .ZN(n8175) );
  NAND2_X1 U10503 ( .A1(n8173), .A2(n8172), .ZN(n8174) );
  NAND2_X1 U10504 ( .A1(n8625), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n8184) );
  NAND2_X1 U10505 ( .A1(n8612), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n8183) );
  INV_X1 U10506 ( .A(n8178), .ZN(n8176) );
  AOI21_X1 U10507 ( .B1(n8176), .B2(P1_REG3_REG_6__SCAN_IN), .A(
        P1_REG3_REG_7__SCAN_IN), .ZN(n8179) );
  NAND2_X1 U10508 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n8177) );
  NOR2_X1 U10509 ( .A1(n8178), .A2(n8177), .ZN(n8198) );
  OR2_X1 U10510 ( .A1(n8179), .A2(n8198), .ZN(n10612) );
  INV_X1 U10511 ( .A(n10612), .ZN(n14458) );
  NAND2_X1 U10512 ( .A1(n8647), .A2(n14458), .ZN(n8182) );
  NAND2_X1 U10513 ( .A1(n8624), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n8181) );
  NAND4_X1 U10514 ( .A1(n8184), .A2(n8183), .A3(n8182), .A4(n8181), .ZN(n13672) );
  MUX2_X1 U10515 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n8111), .Z(n8187) );
  NAND2_X1 U10516 ( .A1(n8187), .A2(SI_7_), .ZN(n8204) );
  OAI21_X1 U10517 ( .B1(n8187), .B2(SI_7_), .A(n8204), .ZN(n8188) );
  INV_X1 U10518 ( .A(n8188), .ZN(n8189) );
  OR2_X1 U10519 ( .A1(n8190), .A2(n8189), .ZN(n8191) );
  NAND2_X1 U10520 ( .A1(n8205), .A2(n8191), .ZN(n9855) );
  OR2_X1 U10521 ( .A1(n9855), .A2(n8266), .ZN(n8195) );
  NAND2_X1 U10522 ( .A1(n8207), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8193) );
  XNOR2_X1 U10523 ( .A(n8193), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9506) );
  AOI22_X1 U10524 ( .A1(n6455), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n8444), .B2(
        n9506), .ZN(n8194) );
  NAND2_X1 U10525 ( .A1(n8195), .A2(n8194), .ZN(n14459) );
  MUX2_X1 U10526 ( .A(n14459), .B(n13672), .S(n6453), .Z(n8196) );
  NAND2_X1 U10527 ( .A1(n8625), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n8203) );
  NAND2_X1 U10528 ( .A1(n8612), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n8202) );
  NAND2_X1 U10529 ( .A1(n8198), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n8224) );
  OR2_X1 U10530 ( .A1(n8198), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n8199) );
  AND2_X1 U10531 ( .A1(n8224), .A2(n8199), .ZN(n11026) );
  NAND2_X1 U10532 ( .A1(n8613), .A2(n11026), .ZN(n8201) );
  NAND2_X1 U10533 ( .A1(n8624), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n8200) );
  NAND4_X1 U10534 ( .A1(n8203), .A2(n8202), .A3(n8201), .A4(n8200), .ZN(n13671) );
  MUX2_X1 U10535 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n9335), .Z(n8206) );
  NAND2_X1 U10536 ( .A1(n8206), .A2(SI_8_), .ZN(n8232) );
  OAI21_X1 U10537 ( .B1(SI_8_), .B2(n8206), .A(n8232), .ZN(n8230) );
  XNOR2_X1 U10538 ( .A(n8231), .B(n8230), .ZN(n9952) );
  NAND2_X1 U10539 ( .A1(n8211), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8209) );
  MUX2_X1 U10540 ( .A(n8209), .B(P1_IR_REG_31__SCAN_IN), .S(n8208), .Z(n8210)
         );
  INV_X1 U10541 ( .A(n8210), .ZN(n8212) );
  NOR2_X1 U10542 ( .A1(n8212), .A2(n8238), .ZN(n9477) );
  AOI22_X1 U10543 ( .A1(n6455), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n8444), .B2(
        n9477), .ZN(n8213) );
  NAND2_X1 U10544 ( .A1(n8214), .A2(n8213), .ZN(n11027) );
  MUX2_X1 U10545 ( .A(n13671), .B(n11027), .S(n6448), .Z(n8218) );
  NAND2_X1 U10546 ( .A1(n8217), .A2(n8218), .ZN(n8216) );
  NAND2_X1 U10547 ( .A1(n8216), .A2(n8215), .ZN(n8222) );
  INV_X1 U10548 ( .A(n8217), .ZN(n8220) );
  INV_X1 U10549 ( .A(n8218), .ZN(n8219) );
  NAND2_X1 U10550 ( .A1(n8220), .A2(n8219), .ZN(n8221) );
  NAND2_X1 U10551 ( .A1(n8222), .A2(n8221), .ZN(n8246) );
  NAND2_X1 U10552 ( .A1(n8612), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n8229) );
  NAND2_X1 U10553 ( .A1(n8625), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n8228) );
  NAND2_X1 U10554 ( .A1(n8224), .A2(n8223), .ZN(n8225) );
  AND2_X1 U10555 ( .A1(n8252), .A2(n8225), .ZN(n11049) );
  NAND2_X1 U10556 ( .A1(n8647), .A2(n11049), .ZN(n8227) );
  NAND2_X1 U10557 ( .A1(n8624), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n8226) );
  NAND4_X1 U10558 ( .A1(n8229), .A2(n8228), .A3(n8227), .A4(n8226), .ZN(n13670) );
  MUX2_X1 U10559 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n6461), .Z(n8233) );
  NAND2_X1 U10560 ( .A1(n8233), .A2(SI_9_), .ZN(n8258) );
  OAI21_X1 U10561 ( .B1(n8233), .B2(SI_9_), .A(n8258), .ZN(n8234) );
  INV_X1 U10562 ( .A(n8234), .ZN(n8235) );
  OR2_X1 U10563 ( .A1(n8236), .A2(n8235), .ZN(n8237) );
  NAND2_X1 U10564 ( .A1(n8259), .A2(n8237), .ZN(n10064) );
  OR2_X1 U10565 ( .A1(n10064), .A2(n8266), .ZN(n8243) );
  INV_X1 U10566 ( .A(n8238), .ZN(n8239) );
  NAND2_X1 U10567 ( .A1(n8239), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8284) );
  INV_X1 U10568 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8240) );
  NAND2_X1 U10569 ( .A1(n8284), .A2(n8240), .ZN(n8267) );
  OR2_X1 U10570 ( .A1(n8284), .A2(n8240), .ZN(n8241) );
  AOI22_X1 U10571 ( .A1(n6455), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n8444), .B2(
        n9602), .ZN(n8242) );
  NAND2_X1 U10572 ( .A1(n8246), .A2(n8247), .ZN(n8245) );
  MUX2_X1 U10573 ( .A(n13670), .B(n11204), .S(n6451), .Z(n8244) );
  INV_X1 U10574 ( .A(n8246), .ZN(n8249) );
  INV_X1 U10575 ( .A(n8247), .ZN(n8248) );
  NAND2_X1 U10576 ( .A1(n8249), .A2(n8248), .ZN(n8250) );
  NAND2_X1 U10577 ( .A1(n8625), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n8257) );
  NAND2_X1 U10578 ( .A1(n8612), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n8256) );
  AND2_X1 U10579 ( .A1(n8252), .A2(n8251), .ZN(n8253) );
  NOR2_X1 U10580 ( .A1(n8274), .A2(n8253), .ZN(n11322) );
  NAND2_X1 U10581 ( .A1(n8613), .A2(n11322), .ZN(n8255) );
  NAND2_X1 U10582 ( .A1(n8624), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n8254) );
  NAND4_X1 U10583 ( .A1(n8257), .A2(n8256), .A3(n8255), .A4(n8254), .ZN(n13669) );
  MUX2_X1 U10584 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n8997), .Z(n8260) );
  NAND2_X1 U10585 ( .A1(n8260), .A2(SI_10_), .ZN(n8280) );
  INV_X1 U10586 ( .A(n8260), .ZN(n8261) );
  NAND2_X1 U10587 ( .A1(n8261), .A2(n9061), .ZN(n8262) );
  OR2_X1 U10588 ( .A1(n8264), .A2(n8263), .ZN(n8265) );
  NAND2_X1 U10589 ( .A1(n8281), .A2(n8265), .ZN(n10121) );
  OR2_X1 U10590 ( .A1(n10121), .A2(n8266), .ZN(n8270) );
  NAND2_X1 U10591 ( .A1(n8267), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8268) );
  XNOR2_X1 U10592 ( .A(n8268), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9580) );
  AOI22_X1 U10593 ( .A1(n6455), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n9580), 
        .B2(n8444), .ZN(n8269) );
  MUX2_X1 U10594 ( .A(n13669), .B(n11327), .S(n6449), .Z(n8272) );
  INV_X1 U10595 ( .A(n8272), .ZN(n8273) );
  NOR2_X1 U10596 ( .A1(n8274), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n8275) );
  OR2_X1 U10597 ( .A1(n8335), .A2(n8275), .ZN(n14393) );
  INV_X1 U10598 ( .A(n14393), .ZN(n10990) );
  NAND2_X1 U10599 ( .A1(n8647), .A2(n10990), .ZN(n8279) );
  NAND2_X1 U10600 ( .A1(n8612), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n8278) );
  NAND2_X1 U10601 ( .A1(n8624), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n8277) );
  NAND2_X1 U10602 ( .A1(n8625), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n8276) );
  NAND4_X1 U10603 ( .A1(n8279), .A2(n8278), .A3(n8277), .A4(n8276), .ZN(n13668) );
  MUX2_X1 U10604 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n6461), .Z(n8293) );
  XNOR2_X1 U10605 ( .A(n8293), .B(SI_11_), .ZN(n8296) );
  XNOR2_X1 U10606 ( .A(n8297), .B(n8296), .ZN(n10356) );
  OR2_X1 U10607 ( .A1(n8282), .A2(n14125), .ZN(n8283) );
  NAND2_X1 U10608 ( .A1(n8284), .A2(n8283), .ZN(n8305) );
  XNOR2_X1 U10609 ( .A(n8305), .B(n15117), .ZN(n9741) );
  AOI22_X1 U10610 ( .A1(n6455), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n8444), 
        .B2(n9741), .ZN(n8285) );
  NAND2_X1 U10611 ( .A1(n8289), .A2(n8290), .ZN(n8288) );
  MUX2_X1 U10612 ( .A(n13668), .B(n14390), .S(n6447), .Z(n8287) );
  NAND2_X1 U10613 ( .A1(n8288), .A2(n8287), .ZN(n8350) );
  INV_X1 U10614 ( .A(n8289), .ZN(n8292) );
  INV_X1 U10615 ( .A(n8290), .ZN(n8291) );
  NAND2_X1 U10616 ( .A1(n8292), .A2(n8291), .ZN(n8349) );
  INV_X1 U10617 ( .A(n8293), .ZN(n8294) );
  NAND2_X1 U10618 ( .A1(n8294), .A2(n9076), .ZN(n8295) );
  MUX2_X1 U10619 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(P1_DATAO_REG_12__SCAN_IN), 
        .S(n6461), .Z(n8298) );
  XNOR2_X1 U10620 ( .A(n8298), .B(n9083), .ZN(n8342) );
  INV_X1 U10621 ( .A(n8298), .ZN(n8299) );
  MUX2_X1 U10622 ( .A(n8300), .B(n9253), .S(n6461), .Z(n8301) );
  XNOR2_X1 U10623 ( .A(n8301), .B(SI_13_), .ZN(n8328) );
  NAND2_X1 U10624 ( .A1(n8327), .A2(n8328), .ZN(n8303) );
  NAND2_X1 U10625 ( .A1(n8301), .A2(n9196), .ZN(n8302) );
  MUX2_X1 U10626 ( .A(n9727), .B(n8304), .S(n6461), .Z(n8359) );
  XNOR2_X1 U10627 ( .A(n8358), .B(n8359), .ZN(n11113) );
  NAND2_X1 U10628 ( .A1(n8306), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8344) );
  NAND2_X1 U10629 ( .A1(n8344), .A2(n8307), .ZN(n8308) );
  NAND2_X1 U10630 ( .A1(n8308), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8329) );
  NAND2_X1 U10631 ( .A1(n8329), .A2(n8309), .ZN(n8310) );
  NAND2_X1 U10632 ( .A1(n8310), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8311) );
  XNOR2_X1 U10633 ( .A(n8311), .B(P1_IR_REG_14__SCAN_IN), .ZN(n10973) );
  AOI22_X1 U10634 ( .A1(n10973), .A2(n8444), .B1(n6455), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n8312) );
  NAND2_X1 U10635 ( .A1(n8335), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8337) );
  NAND2_X1 U10636 ( .A1(n8322), .A2(n8314), .ZN(n8315) );
  NAND2_X1 U10637 ( .A1(n8368), .A2(n8315), .ZN(n14350) );
  INV_X1 U10638 ( .A(n14350), .ZN(n11177) );
  NAND2_X1 U10639 ( .A1(n8647), .A2(n11177), .ZN(n8319) );
  NAND2_X1 U10640 ( .A1(n8612), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n8318) );
  NAND2_X1 U10641 ( .A1(n8624), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n8317) );
  NAND2_X1 U10642 ( .A1(n8625), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n8316) );
  NAND2_X1 U10643 ( .A1(n11174), .A2(n12166), .ZN(n8374) );
  NAND2_X1 U10644 ( .A1(n11380), .A2(n8374), .ZN(n11173) );
  NAND2_X1 U10645 ( .A1(n8337), .A2(n8320), .ZN(n8321) );
  NAND2_X1 U10646 ( .A1(n8322), .A2(n8321), .ZN(n14279) );
  INV_X1 U10647 ( .A(n14279), .ZN(n11626) );
  NAND2_X1 U10648 ( .A1(n8613), .A2(n11626), .ZN(n8326) );
  NAND2_X1 U10649 ( .A1(n8612), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n8325) );
  NAND2_X1 U10650 ( .A1(n8624), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n8324) );
  NAND2_X1 U10651 ( .A1(n8625), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n8323) );
  NAND4_X1 U10652 ( .A1(n8326), .A2(n8325), .A3(n8324), .A4(n8323), .ZN(n13666) );
  XNOR2_X1 U10653 ( .A(n8327), .B(n8328), .ZN(n10718) );
  XNOR2_X1 U10654 ( .A(n8329), .B(P1_IR_REG_13__SCAN_IN), .ZN(n10055) );
  AOI22_X1 U10655 ( .A1(n10055), .A2(n8444), .B1(n6455), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n8330) );
  MUX2_X1 U10656 ( .A(n13666), .B(n11621), .S(n6453), .Z(n8355) );
  INV_X1 U10657 ( .A(n13666), .ZN(n14341) );
  NAND2_X1 U10658 ( .A1(n14341), .A2(n6454), .ZN(n8332) );
  OAI21_X1 U10659 ( .B1(n11621), .B2(n6453), .A(n8332), .ZN(n8333) );
  NOR2_X1 U10660 ( .A1(n8355), .A2(n8333), .ZN(n8334) );
  NAND2_X1 U10661 ( .A1(n8625), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n8341) );
  NAND2_X1 U10662 ( .A1(n8612), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n8340) );
  OR2_X1 U10663 ( .A1(n8335), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8336) );
  AND2_X1 U10664 ( .A1(n8337), .A2(n8336), .ZN(n11535) );
  NAND2_X1 U10665 ( .A1(n8647), .A2(n11535), .ZN(n8339) );
  NAND2_X1 U10666 ( .A1(n8624), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n8338) );
  XNOR2_X1 U10667 ( .A(n8343), .B(n8342), .ZN(n10643) );
  XNOR2_X1 U10668 ( .A(n8344), .B(P1_IR_REG_12__SCAN_IN), .ZN(n9936) );
  AOI22_X1 U10669 ( .A1(n9936), .A2(n8444), .B1(n6455), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n8345) );
  MUX2_X1 U10670 ( .A(n14376), .B(n11538), .S(n6454), .Z(n8353) );
  INV_X1 U10671 ( .A(n14376), .ZN(n13667) );
  MUX2_X1 U10672 ( .A(n13667), .B(n11266), .S(n6451), .Z(n8352) );
  NAND2_X1 U10673 ( .A1(n8353), .A2(n8352), .ZN(n8347) );
  NAND3_X1 U10674 ( .A1(n8350), .A2(n8349), .A3(n8348), .ZN(n8380) );
  INV_X1 U10675 ( .A(n8351), .ZN(n8354) );
  INV_X1 U10676 ( .A(n8355), .ZN(n8357) );
  MUX2_X1 U10677 ( .A(n13666), .B(n11621), .S(n6449), .Z(n8356) );
  OR3_X1 U10678 ( .A1(n11173), .A2(n8357), .A3(n8356), .ZN(n8377) );
  MUX2_X1 U10679 ( .A(n9907), .B(n9888), .S(n6461), .Z(n8398) );
  XNOR2_X1 U10680 ( .A(n8398), .B(SI_15_), .ZN(n8360) );
  XNOR2_X1 U10681 ( .A(n8361), .B(n8360), .ZN(n11286) );
  NAND2_X1 U10682 ( .A1(n8362), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8363) );
  MUX2_X1 U10683 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8363), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n8364) );
  AND2_X1 U10684 ( .A1(n8364), .A2(n8038), .ZN(n14447) );
  AOI22_X1 U10685 ( .A1(n6455), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n8444), 
        .B2(n14447), .ZN(n8365) );
  NAND2_X1 U10686 ( .A1(n8625), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n8373) );
  NAND2_X1 U10687 ( .A1(n8612), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n8372) );
  AND2_X1 U10688 ( .A1(n8368), .A2(n8367), .ZN(n8369) );
  NOR2_X1 U10689 ( .A1(n8386), .A2(n8369), .ZN(n13650) );
  NAND2_X1 U10690 ( .A1(n8647), .A2(n13650), .ZN(n8371) );
  NAND2_X1 U10691 ( .A1(n8624), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n8370) );
  NAND2_X1 U10692 ( .A1(n14397), .A2(n14340), .ZN(n8697) );
  NAND2_X1 U10693 ( .A1(n8697), .A2(n8374), .ZN(n8375) );
  NAND2_X1 U10694 ( .A1(n8375), .A2(n6453), .ZN(n8376) );
  NOR2_X1 U10695 ( .A1(n7330), .A2(n8378), .ZN(n8379) );
  NAND2_X1 U10696 ( .A1(n8380), .A2(n8379), .ZN(n8381) );
  NAND2_X1 U10697 ( .A1(n8381), .A2(n11452), .ZN(n8384) );
  NAND2_X1 U10698 ( .A1(n11452), .A2(n11380), .ZN(n8382) );
  NAND2_X1 U10699 ( .A1(n8382), .A2(n6449), .ZN(n8383) );
  NAND2_X1 U10700 ( .A1(n8384), .A2(n8383), .ZN(n8385) );
  NOR2_X1 U10701 ( .A1(n8386), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8387) );
  OR2_X1 U10702 ( .A1(n8417), .A2(n8387), .ZN(n14364) );
  NAND2_X1 U10703 ( .A1(n8624), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n8388) );
  OAI21_X1 U10704 ( .B1(n14364), .B2(n8118), .A(n8388), .ZN(n8389) );
  INV_X1 U10705 ( .A(n8389), .ZN(n8393) );
  NAND2_X1 U10706 ( .A1(n8625), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n8391) );
  NAND2_X1 U10707 ( .A1(n8612), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8390) );
  AND2_X1 U10708 ( .A1(n8391), .A2(n8390), .ZN(n8392) );
  INV_X1 U10709 ( .A(n8398), .ZN(n8394) );
  NAND2_X1 U10710 ( .A1(n8394), .A2(SI_15_), .ZN(n8399) );
  NAND2_X1 U10711 ( .A1(n8397), .A2(SI_14_), .ZN(n8395) );
  NOR2_X1 U10712 ( .A1(n8397), .A2(SI_14_), .ZN(n8400) );
  INV_X1 U10713 ( .A(SI_15_), .ZN(n9616) );
  AOI22_X1 U10714 ( .A1(n8400), .A2(n8399), .B1(n9616), .B2(n8398), .ZN(n8401)
         );
  MUX2_X1 U10715 ( .A(n9725), .B(n9733), .S(n6461), .Z(n8410) );
  XNOR2_X1 U10716 ( .A(n8410), .B(SI_16_), .ZN(n8408) );
  XNOR2_X1 U10717 ( .A(n8409), .B(n8408), .ZN(n11347) );
  NAND2_X1 U10718 ( .A1(n8038), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8403) );
  XNOR2_X1 U10719 ( .A(n8403), .B(P1_IR_REG_16__SCAN_IN), .ZN(n13733) );
  AOI22_X1 U10720 ( .A1(n6455), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n8444), 
        .B2(n13733), .ZN(n8404) );
  MUX2_X1 U10721 ( .A(n14366), .B(n14124), .S(n6454), .Z(n8407) );
  INV_X1 U10722 ( .A(n14366), .ZN(n13663) );
  INV_X1 U10723 ( .A(n14124), .ZN(n14360) );
  MUX2_X1 U10724 ( .A(n13663), .B(n14360), .S(n6448), .Z(n8406) );
  NAND2_X1 U10725 ( .A1(n8410), .A2(n9797), .ZN(n8411) );
  MUX2_X1 U10726 ( .A(n9833), .B(n9794), .S(n6461), .Z(n8425) );
  XNOR2_X1 U10727 ( .A(n8425), .B(SI_17_), .ZN(n8412) );
  XNOR2_X1 U10728 ( .A(n8427), .B(n8412), .ZN(n11427) );
  OR2_X1 U10729 ( .A1(n8413), .A2(n14125), .ZN(n8414) );
  XNOR2_X1 U10730 ( .A(n8414), .B(P1_IR_REG_17__SCAN_IN), .ZN(n13741) );
  AOI22_X1 U10731 ( .A1(n6455), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n8444), 
        .B2(n13741), .ZN(n8415) );
  NOR2_X1 U10732 ( .A1(n8417), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8418) );
  OR2_X1 U10733 ( .A1(n8432), .A2(n8418), .ZN(n14375) );
  AOI22_X1 U10734 ( .A1(n8625), .A2(P1_REG0_REG_17__SCAN_IN), .B1(n8624), .B2(
        P1_REG1_REG_17__SCAN_IN), .ZN(n8420) );
  NAND2_X1 U10735 ( .A1(n8612), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8419) );
  OAI211_X1 U10736 ( .C1(n14375), .C2(n8118), .A(n8420), .B(n8419), .ZN(n13953) );
  OR2_X1 U10737 ( .A1(n14372), .A2(n13953), .ZN(n12102) );
  NAND2_X1 U10738 ( .A1(n8423), .A2(n8422), .ZN(n8424) );
  MUX2_X1 U10739 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n6461), .Z(n8436) );
  XNOR2_X1 U10740 ( .A(n8438), .B(n8436), .ZN(n11539) );
  NAND2_X1 U10741 ( .A1(n8428), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8429) );
  XNOR2_X1 U10742 ( .A(n8429), .B(P1_IR_REG_18__SCAN_IN), .ZN(n13759) );
  AOI22_X1 U10743 ( .A1(n6455), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n8444), 
        .B2(n13759), .ZN(n8430) );
  OR2_X1 U10744 ( .A1(n8432), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n8433) );
  NAND2_X1 U10745 ( .A1(n8448), .A2(n8433), .ZN(n13964) );
  AOI22_X1 U10746 ( .A1(n8625), .A2(P1_REG0_REG_18__SCAN_IN), .B1(n8612), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n8435) );
  NAND2_X1 U10747 ( .A1(n8624), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n8434) );
  OAI211_X1 U10748 ( .C1(n13964), .C2(n8118), .A(n8435), .B(n8434), .ZN(n13662) );
  NAND2_X1 U10749 ( .A1(n13967), .A2(n13662), .ZN(n12103) );
  INV_X1 U10750 ( .A(n8436), .ZN(n8437) );
  NAND2_X1 U10751 ( .A1(n8439), .A2(SI_18_), .ZN(n8440) );
  MUX2_X1 U10752 ( .A(n10063), .B(n11637), .S(n6461), .Z(n8441) );
  INV_X1 U10753 ( .A(n8441), .ZN(n8442) );
  NAND2_X1 U10754 ( .A1(n8442), .A2(SI_19_), .ZN(n8443) );
  NAND2_X1 U10755 ( .A1(n8465), .A2(n8443), .ZN(n8466) );
  XNOR2_X1 U10756 ( .A(n8467), .B(n8466), .ZN(n11897) );
  AOI22_X1 U10757 ( .A1(n6455), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n13878), 
        .B2(n8444), .ZN(n8445) );
  INV_X1 U10758 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8447) );
  NAND2_X1 U10759 ( .A1(n8448), .A2(n8447), .ZN(n8449) );
  NAND2_X1 U10760 ( .A1(n8458), .A2(n8449), .ZN(n13939) );
  AOI22_X1 U10761 ( .A1(n8625), .A2(P1_REG0_REG_19__SCAN_IN), .B1(n8612), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n8451) );
  NAND2_X1 U10762 ( .A1(n8624), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n8450) );
  OAI211_X1 U10763 ( .C1(n13939), .C2(n8118), .A(n8451), .B(n8450), .ZN(n13956) );
  XNOR2_X1 U10764 ( .A(n14063), .B(n13956), .ZN(n13931) );
  MUX2_X1 U10765 ( .A(n13662), .B(n13967), .S(n6453), .Z(n8452) );
  NAND2_X1 U10766 ( .A1(n13956), .A2(n6451), .ZN(n8455) );
  OR2_X1 U10767 ( .A1(n13956), .A2(n6451), .ZN(n8454) );
  MUX2_X1 U10768 ( .A(n8455), .B(n8454), .S(n14063), .Z(n8456) );
  NAND2_X1 U10769 ( .A1(n8457), .A2(n8456), .ZN(n8472) );
  INV_X1 U10770 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13600) );
  AOI21_X1 U10771 ( .B1(n8458), .B2(n13600), .A(n8475), .ZN(n13916) );
  NAND2_X1 U10772 ( .A1(n13916), .A2(n8613), .ZN(n8464) );
  INV_X1 U10773 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n8461) );
  NAND2_X1 U10774 ( .A1(n8624), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n8460) );
  NAND2_X1 U10775 ( .A1(n8612), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n8459) );
  OAI211_X1 U10776 ( .C1(n8630), .C2(n8461), .A(n8460), .B(n8459), .ZN(n8462)
         );
  INV_X1 U10777 ( .A(n8462), .ZN(n8463) );
  INV_X1 U10778 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n10585) );
  MUX2_X1 U10779 ( .A(n7736), .B(n10585), .S(n6461), .Z(n8480) );
  XNOR2_X1 U10780 ( .A(n8482), .B(n8480), .ZN(n11918) );
  OR2_X1 U10781 ( .A1(n8681), .A2(n7736), .ZN(n8468) );
  MUX2_X1 U10782 ( .A(n13938), .B(n14114), .S(n6447), .Z(n8471) );
  INV_X1 U10783 ( .A(n13938), .ZN(n13900) );
  MUX2_X1 U10784 ( .A(n13900), .B(n8688), .S(n6454), .Z(n8470) );
  OAI21_X1 U10785 ( .B1(n8472), .B2(n8471), .A(n8470), .ZN(n8474) );
  NAND2_X1 U10786 ( .A1(n8472), .A2(n8471), .ZN(n8473) );
  NAND2_X1 U10787 ( .A1(n8625), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n8479) );
  NAND2_X1 U10788 ( .A1(n8612), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n8478) );
  NAND2_X1 U10789 ( .A1(n8475), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8490) );
  OAI21_X1 U10790 ( .B1(P1_REG3_REG_21__SCAN_IN), .B2(n8475), .A(n8490), .ZN(
        n13567) );
  INV_X1 U10791 ( .A(n13567), .ZN(n13904) );
  NAND2_X1 U10792 ( .A1(n8647), .A2(n13904), .ZN(n8477) );
  NAND2_X1 U10793 ( .A1(n8624), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n8476) );
  NAND4_X1 U10794 ( .A1(n8479), .A2(n8478), .A3(n8477), .A4(n8476), .ZN(n13661) );
  INV_X1 U10795 ( .A(n8480), .ZN(n8481) );
  MUX2_X1 U10796 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n6461), .Z(n8499) );
  XNOR2_X1 U10797 ( .A(n8499), .B(SI_21_), .ZN(n8497) );
  XNOR2_X1 U10798 ( .A(n8498), .B(n8497), .ZN(n11934) );
  OR2_X1 U10799 ( .A1(n8681), .A2(n10850), .ZN(n8485) );
  MUX2_X1 U10800 ( .A(n13661), .B(n14051), .S(n6449), .Z(n8487) );
  INV_X1 U10801 ( .A(n8488), .ZN(n8489) );
  NAND2_X1 U10802 ( .A1(n8612), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n8496) );
  NAND2_X1 U10803 ( .A1(n8625), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n8495) );
  INV_X1 U10804 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13610) );
  NAND2_X1 U10805 ( .A1(n13610), .A2(n8490), .ZN(n8492) );
  INV_X1 U10806 ( .A(n8490), .ZN(n8491) );
  NAND2_X1 U10807 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(n8491), .ZN(n8509) );
  AND2_X1 U10808 ( .A1(n8492), .A2(n8509), .ZN(n13891) );
  NAND2_X1 U10809 ( .A1(n8613), .A2(n13891), .ZN(n8494) );
  NAND2_X1 U10810 ( .A1(n8624), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n8493) );
  NAND4_X1 U10811 ( .A1(n8496), .A2(n8495), .A3(n8494), .A4(n8493), .ZN(n13901) );
  XNOR2_X1 U10812 ( .A(n8537), .B(SI_22_), .ZN(n11145) );
  MUX2_X1 U10813 ( .A(n13901), .B(n13888), .S(n6448), .Z(n8503) );
  NAND2_X1 U10814 ( .A1(n8502), .A2(n8503), .ZN(n8501) );
  NAND2_X1 U10815 ( .A1(n8501), .A2(n8500), .ZN(n8507) );
  INV_X1 U10816 ( .A(n8502), .ZN(n8505) );
  INV_X1 U10817 ( .A(n8503), .ZN(n8504) );
  NAND2_X1 U10818 ( .A1(n8505), .A2(n8504), .ZN(n8506) );
  NAND2_X1 U10819 ( .A1(n8507), .A2(n8506), .ZN(n8524) );
  NAND2_X1 U10820 ( .A1(n8625), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n8514) );
  NAND2_X1 U10821 ( .A1(n8612), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n8513) );
  INV_X1 U10822 ( .A(n8509), .ZN(n8508) );
  NAND2_X1 U10823 ( .A1(n8508), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n8529) );
  INV_X1 U10824 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n15040) );
  NAND2_X1 U10825 ( .A1(n8509), .A2(n15040), .ZN(n8510) );
  AND2_X1 U10826 ( .A1(n8529), .A2(n8510), .ZN(n13876) );
  NAND2_X1 U10827 ( .A1(n8647), .A2(n13876), .ZN(n8512) );
  NAND2_X1 U10828 ( .A1(n8624), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n8511) );
  NAND4_X1 U10829 ( .A1(n8514), .A2(n8513), .A3(n8512), .A4(n8511), .ZN(n13660) );
  INV_X1 U10830 ( .A(n11145), .ZN(n8515) );
  MUX2_X1 U10831 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n9335), .Z(n11144) );
  NAND2_X1 U10832 ( .A1(n8515), .A2(n11144), .ZN(n8517) );
  NAND2_X1 U10833 ( .A1(n8537), .A2(SI_22_), .ZN(n8516) );
  NAND2_X1 U10834 ( .A1(n8517), .A2(n8516), .ZN(n8519) );
  MUX2_X1 U10835 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n6461), .Z(n8541) );
  XNOR2_X1 U10836 ( .A(n8541), .B(SI_23_), .ZN(n8518) );
  INV_X1 U10837 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11245) );
  OR2_X1 U10838 ( .A1(n8681), .A2(n11245), .ZN(n8520) );
  NAND2_X2 U10839 ( .A1(n8521), .A2(n8520), .ZN(n13869) );
  MUX2_X1 U10840 ( .A(n13660), .B(n13869), .S(n6454), .Z(n8525) );
  NAND2_X1 U10841 ( .A1(n8524), .A2(n8525), .ZN(n8523) );
  MUX2_X1 U10842 ( .A(n13660), .B(n13869), .S(n6449), .Z(n8522) );
  NAND2_X1 U10843 ( .A1(n8523), .A2(n8522), .ZN(n8550) );
  INV_X1 U10844 ( .A(n8524), .ZN(n8527) );
  INV_X1 U10845 ( .A(n8525), .ZN(n8526) );
  NAND2_X1 U10846 ( .A1(n8527), .A2(n8526), .ZN(n8553) );
  NAND2_X1 U10847 ( .A1(n8550), .A2(n8553), .ZN(n8547) );
  NAND2_X1 U10848 ( .A1(n8625), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n8534) );
  NAND2_X1 U10849 ( .A1(n8612), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n8533) );
  INV_X1 U10850 ( .A(n8529), .ZN(n8528) );
  NAND2_X1 U10851 ( .A1(n8528), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n8558) );
  INV_X1 U10852 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n13588) );
  NAND2_X1 U10853 ( .A1(n8529), .A2(n13588), .ZN(n8530) );
  AND2_X1 U10854 ( .A1(n8558), .A2(n8530), .ZN(n13860) );
  NAND2_X1 U10855 ( .A1(n8613), .A2(n13860), .ZN(n8532) );
  NAND2_X1 U10856 ( .A1(n8624), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n8531) );
  INV_X1 U10857 ( .A(n11144), .ZN(n8539) );
  INV_X1 U10858 ( .A(n8541), .ZN(n8535) );
  AOI22_X1 U10859 ( .A1(n8538), .A2(n8539), .B1(n8535), .B2(n10945), .ZN(n8536) );
  OAI21_X1 U10860 ( .B1(n8539), .B2(n8538), .A(n10945), .ZN(n8542) );
  AND2_X1 U10861 ( .A1(SI_23_), .A2(SI_22_), .ZN(n8540) );
  AOI22_X1 U10862 ( .A1(n8542), .A2(n8541), .B1(n11144), .B2(n8540), .ZN(n8543) );
  MUX2_X1 U10863 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n9335), .Z(n8564) );
  OR2_X1 U10864 ( .A1(n8681), .A2(n11273), .ZN(n8545) );
  MUX2_X1 U10865 ( .A(n13581), .B(n14104), .S(n6453), .Z(n8551) );
  NAND2_X1 U10866 ( .A1(n8547), .A2(n8551), .ZN(n8549) );
  MUX2_X1 U10867 ( .A(n13581), .B(n14104), .S(n6451), .Z(n8548) );
  NAND2_X1 U10868 ( .A1(n8549), .A2(n8548), .ZN(n8556) );
  INV_X1 U10869 ( .A(n8551), .ZN(n8552) );
  AND2_X1 U10870 ( .A1(n8553), .A2(n8552), .ZN(n8554) );
  NAND2_X1 U10871 ( .A1(n8550), .A2(n8554), .ZN(n8555) );
  NAND2_X1 U10872 ( .A1(n8625), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n8563) );
  NAND2_X1 U10873 ( .A1(n8612), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n8562) );
  INV_X1 U10874 ( .A(n8558), .ZN(n8557) );
  NAND2_X1 U10875 ( .A1(n8557), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n8578) );
  INV_X1 U10876 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n13580) );
  NAND2_X1 U10877 ( .A1(n8558), .A2(n13580), .ZN(n8559) );
  AND2_X1 U10878 ( .A1(n8578), .A2(n8559), .ZN(n13579) );
  NAND2_X1 U10879 ( .A1(n8613), .A2(n13579), .ZN(n8561) );
  NAND2_X1 U10880 ( .A1(n8624), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n8560) );
  NAND4_X1 U10881 ( .A1(n8563), .A2(n8562), .A3(n8561), .A4(n8560), .ZN(n13659) );
  INV_X1 U10882 ( .A(n8564), .ZN(n8567) );
  NAND2_X1 U10883 ( .A1(n8565), .A2(SI_24_), .ZN(n8566) );
  MUX2_X1 U10884 ( .A(n11374), .B(n11377), .S(n6461), .Z(n8569) );
  NAND2_X1 U10885 ( .A1(n8569), .A2(n11341), .ZN(n8584) );
  INV_X1 U10886 ( .A(n8569), .ZN(n8570) );
  NAND2_X1 U10887 ( .A1(n8570), .A2(SI_25_), .ZN(n8571) );
  NAND2_X1 U10888 ( .A1(n8584), .A2(n8571), .ZN(n8585) );
  XNOR2_X1 U10889 ( .A(n8586), .B(n8585), .ZN(n12000) );
  OR2_X1 U10890 ( .A1(n8681), .A2(n11374), .ZN(n8572) );
  MUX2_X1 U10891 ( .A(n13659), .B(n14028), .S(n6451), .Z(n8574) );
  NAND2_X1 U10892 ( .A1(n8625), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n8583) );
  NAND2_X1 U10893 ( .A1(n8612), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n8582) );
  INV_X1 U10894 ( .A(n8578), .ZN(n8576) );
  NAND2_X1 U10895 ( .A1(n8576), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8599) );
  INV_X1 U10896 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8577) );
  NAND2_X1 U10897 ( .A1(n8578), .A2(n8577), .ZN(n8579) );
  AND2_X1 U10898 ( .A1(n8599), .A2(n8579), .ZN(n13635) );
  NAND2_X1 U10899 ( .A1(n8613), .A2(n13635), .ZN(n8581) );
  NAND2_X1 U10900 ( .A1(n8624), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n8580) );
  NAND4_X1 U10901 ( .A1(n8583), .A2(n8582), .A3(n8581), .A4(n8580), .ZN(n13828) );
  MUX2_X1 U10902 ( .A(n11513), .B(n11488), .S(n6461), .Z(n8605) );
  XNOR2_X1 U10903 ( .A(n8605), .B(SI_26_), .ZN(n8587) );
  XNOR2_X1 U10904 ( .A(n8606), .B(n8587), .ZN(n11774) );
  OR2_X1 U10905 ( .A1(n8681), .A2(n11513), .ZN(n8588) );
  MUX2_X1 U10906 ( .A(n13828), .B(n13640), .S(n6447), .Z(n8593) );
  NAND2_X1 U10907 ( .A1(n8592), .A2(n8593), .ZN(n8591) );
  MUX2_X1 U10908 ( .A(n13828), .B(n13640), .S(n6454), .Z(n8590) );
  NAND2_X1 U10909 ( .A1(n8591), .A2(n8590), .ZN(n8597) );
  INV_X1 U10910 ( .A(n8592), .ZN(n8595) );
  INV_X1 U10911 ( .A(n8593), .ZN(n8594) );
  NAND2_X1 U10912 ( .A1(n8595), .A2(n8594), .ZN(n8596) );
  NAND2_X1 U10913 ( .A1(n8625), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n8604) );
  NAND2_X1 U10914 ( .A1(n8612), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n8603) );
  INV_X1 U10915 ( .A(n8599), .ZN(n8598) );
  NAND2_X1 U10916 ( .A1(n8598), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n8646) );
  INV_X1 U10917 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n13530) );
  NAND2_X1 U10918 ( .A1(n8599), .A2(n13530), .ZN(n8600) );
  AND2_X1 U10919 ( .A1(n8646), .A2(n8600), .ZN(n13529) );
  NAND2_X1 U10920 ( .A1(n8613), .A2(n13529), .ZN(n8602) );
  NAND2_X1 U10921 ( .A1(n8624), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n8601) );
  NAND4_X1 U10922 ( .A1(n8604), .A2(n8603), .A3(n8602), .A4(n8601), .ZN(n13658) );
  MUX2_X1 U10923 ( .A(n14134), .B(n13524), .S(n6461), .Z(n8618) );
  XNOR2_X1 U10924 ( .A(n8618), .B(SI_27_), .ZN(n8607) );
  OR2_X1 U10925 ( .A1(n8681), .A2(n14134), .ZN(n8608) );
  MUX2_X1 U10926 ( .A(n13658), .B(n14014), .S(n6453), .Z(n8611) );
  MUX2_X1 U10927 ( .A(n13658), .B(n14014), .S(n6448), .Z(n8610) );
  NAND2_X1 U10928 ( .A1(n8625), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n8617) );
  NAND2_X1 U10929 ( .A1(n8612), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n8616) );
  XNOR2_X1 U10930 ( .A(n8646), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n12122) );
  NAND2_X1 U10931 ( .A1(n8613), .A2(n12122), .ZN(n8615) );
  NAND2_X1 U10932 ( .A1(n8624), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n8614) );
  NAND4_X1 U10933 ( .A1(n8617), .A2(n8616), .A3(n8615), .A4(n8614), .ZN(n13657) );
  OAI21_X1 U10934 ( .B1(n8619), .B2(n12884), .A(n8618), .ZN(n8621) );
  NAND2_X1 U10935 ( .A1(n8621), .A2(n8620), .ZN(n8633) );
  MUX2_X1 U10936 ( .A(n11683), .B(n15043), .S(n9335), .Z(n8634) );
  XNOR2_X1 U10937 ( .A(n8634), .B(SI_28_), .ZN(n8632) );
  XNOR2_X1 U10938 ( .A(n8633), .B(n8632), .ZN(n11752) );
  OR2_X1 U10939 ( .A1(n8681), .A2(n11683), .ZN(n8622) );
  MUX2_X1 U10940 ( .A(n13657), .B(n14009), .S(n6451), .Z(n8657) );
  INV_X1 U10941 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n15044) );
  NAND2_X1 U10942 ( .A1(n8612), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n8627) );
  NAND2_X1 U10943 ( .A1(n8625), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8626) );
  OAI211_X1 U10944 ( .C1(n8180), .C2(n15044), .A(n8627), .B(n8626), .ZN(n13776) );
  INV_X1 U10945 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n14090) );
  NAND2_X1 U10946 ( .A1(n8612), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8629) );
  NAND2_X1 U10947 ( .A1(n8624), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8628) );
  OAI211_X1 U10948 ( .C1(n8630), .C2(n14090), .A(n8629), .B(n8628), .ZN(n13655) );
  OAI21_X1 U10949 ( .B1(n13776), .B2(n10586), .A(n13655), .ZN(n8631) );
  INV_X1 U10950 ( .A(n8631), .ZN(n8641) );
  NAND2_X1 U10951 ( .A1(n8633), .A2(n8632), .ZN(n8636) );
  NAND2_X1 U10952 ( .A1(n8634), .A2(n12881), .ZN(n8635) );
  NAND2_X1 U10953 ( .A1(n8636), .A2(n8635), .ZN(n8653) );
  INV_X1 U10954 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14131) );
  INV_X1 U10955 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n11737) );
  MUX2_X1 U10956 ( .A(n14131), .B(n11737), .S(n6461), .Z(n8637) );
  XNOR2_X1 U10957 ( .A(n8637), .B(SI_29_), .ZN(n8652) );
  NAND2_X1 U10958 ( .A1(n8637), .A2(n12159), .ZN(n8638) );
  MUX2_X1 U10959 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n6461), .Z(n8675) );
  INV_X1 U10960 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n12132) );
  OR2_X1 U10961 ( .A1(n8681), .A2(n12132), .ZN(n8639) );
  MUX2_X1 U10962 ( .A(n8641), .B(n13781), .S(n6454), .Z(n8663) );
  NAND2_X1 U10963 ( .A1(n13776), .A2(n6454), .ZN(n8643) );
  INV_X1 U10964 ( .A(n13655), .ZN(n8642) );
  AOI21_X1 U10965 ( .B1(n8644), .B2(n8643), .A(n8642), .ZN(n8645) );
  AOI21_X1 U10966 ( .B1(n13781), .B2(n6449), .A(n8645), .ZN(n8665) );
  NAND2_X1 U10967 ( .A1(n6457), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8651) );
  NAND2_X1 U10968 ( .A1(n8612), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8650) );
  INV_X1 U10969 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n12271) );
  NOR2_X1 U10970 ( .A1(n8646), .A2(n12271), .ZN(n12146) );
  NAND2_X1 U10971 ( .A1(n8647), .A2(n12146), .ZN(n8649) );
  NAND2_X1 U10972 ( .A1(n8624), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n8648) );
  NOR2_X1 U10973 ( .A1(n8681), .A2(n14131), .ZN(n8654) );
  MUX2_X1 U10974 ( .A(n12273), .B(n14001), .S(n6448), .Z(n8660) );
  INV_X1 U10975 ( .A(n14001), .ZN(n12143) );
  MUX2_X1 U10976 ( .A(n13656), .B(n12143), .S(n6453), .Z(n8659) );
  AOI22_X1 U10977 ( .A1(n8663), .A2(n8665), .B1(n8660), .B2(n8659), .ZN(n8655)
         );
  OAI21_X1 U10978 ( .B1(n8658), .B2(n8657), .A(n8655), .ZN(n8672) );
  INV_X1 U10979 ( .A(n14009), .ZN(n12265) );
  MUX2_X1 U10980 ( .A(n13794), .B(n12265), .S(n6453), .Z(n8656) );
  AOI21_X1 U10981 ( .B1(n8658), .B2(n8657), .A(n8656), .ZN(n8671) );
  INV_X1 U10982 ( .A(n8659), .ZN(n8662) );
  INV_X1 U10983 ( .A(n8660), .ZN(n8661) );
  NAND2_X1 U10984 ( .A1(n8662), .A2(n8661), .ZN(n8664) );
  NAND2_X1 U10985 ( .A1(n8665), .A2(n8664), .ZN(n8669) );
  INV_X1 U10986 ( .A(n8663), .ZN(n8668) );
  INV_X1 U10987 ( .A(n8664), .ZN(n8667) );
  INV_X1 U10988 ( .A(n8665), .ZN(n8666) );
  AOI22_X1 U10989 ( .A1(n8669), .A2(n8668), .B1(n8667), .B2(n8666), .ZN(n8670)
         );
  NAND2_X1 U10990 ( .A1(n9824), .A2(n10586), .ZN(n8673) );
  NAND2_X1 U10991 ( .A1(n9814), .A2(n8673), .ZN(n8674) );
  INV_X1 U10992 ( .A(n9416), .ZN(n9417) );
  NAND2_X1 U10993 ( .A1(n9417), .A2(n13878), .ZN(n10311) );
  NAND2_X1 U10994 ( .A1(n8674), .A2(n10311), .ZN(n8705) );
  INV_X1 U10995 ( .A(n8705), .ZN(n8684) );
  NAND2_X1 U10996 ( .A1(n8675), .A2(SI_30_), .ZN(n8676) );
  MUX2_X1 U10997 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n6461), .Z(n8678) );
  XNOR2_X1 U10998 ( .A(n8678), .B(SI_31_), .ZN(n8679) );
  INV_X1 U10999 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n8680) );
  OR2_X1 U11000 ( .A1(n8681), .A2(n8680), .ZN(n8682) );
  XNOR2_X1 U11001 ( .A(n13773), .B(n13776), .ZN(n8702) );
  NAND3_X1 U11002 ( .A1(n8717), .A2(n8684), .A3(n8702), .ZN(n8714) );
  XNOR2_X1 U11003 ( .A(n14001), .B(n13656), .ZN(n12140) );
  INV_X1 U11004 ( .A(n13658), .ZN(n12274) );
  XNOR2_X1 U11005 ( .A(n14014), .B(n12274), .ZN(n13786) );
  NAND2_X1 U11006 ( .A1(n14009), .A2(n13794), .ZN(n12138) );
  OR2_X1 U11007 ( .A1(n14009), .A2(n13794), .ZN(n8685) );
  NAND2_X1 U11008 ( .A1(n13640), .A2(n13792), .ZN(n13788) );
  OR2_X1 U11009 ( .A1(n13640), .A2(n13792), .ZN(n8686) );
  NAND2_X1 U11010 ( .A1(n13788), .A2(n8686), .ZN(n13809) );
  XNOR2_X1 U11011 ( .A(n13859), .B(n13581), .ZN(n13849) );
  INV_X1 U11012 ( .A(n13660), .ZN(n13851) );
  XNOR2_X1 U11013 ( .A(n13869), .B(n13851), .ZN(n12091) );
  INV_X1 U11014 ( .A(n13661), .ZN(n12086) );
  XNOR2_X1 U11015 ( .A(n14051), .B(n12086), .ZN(n13907) );
  XNOR2_X1 U11016 ( .A(n8687), .B(n13901), .ZN(n13885) );
  NAND2_X1 U11017 ( .A1(n8688), .A2(n13938), .ZN(n8689) );
  NAND2_X1 U11018 ( .A1(n12085), .A2(n8689), .ZN(n13917) );
  NAND2_X1 U11019 ( .A1(n12102), .A2(n6539), .ZN(n13972) );
  XNOR2_X1 U11020 ( .A(n11266), .B(n14376), .ZN(n11104) );
  XNOR2_X1 U11021 ( .A(n14390), .B(n11532), .ZN(n11099) );
  XNOR2_X1 U11022 ( .A(n11327), .B(n14379), .ZN(n10635) );
  INV_X1 U11023 ( .A(n13671), .ZN(n11201) );
  XNOR2_X1 U11024 ( .A(n11027), .B(n11201), .ZN(n10625) );
  XNOR2_X1 U11025 ( .A(n11204), .B(n13670), .ZN(n10949) );
  NAND4_X1 U11026 ( .A1(n10291), .A2(n10288), .A3(n10444), .A4(n10275), .ZN(
        n8692) );
  INV_X1 U11027 ( .A(n13673), .ZN(n10392) );
  XNOR2_X1 U11028 ( .A(n10596), .B(n10392), .ZN(n10389) );
  INV_X1 U11029 ( .A(n13676), .ZN(n13547) );
  NAND2_X1 U11030 ( .A1(n13547), .A2(n10615), .ZN(n10293) );
  NAND2_X1 U11031 ( .A1(n13676), .A2(n14521), .ZN(n10294) );
  AND2_X1 U11032 ( .A1(n10293), .A2(n10294), .ZN(n10620) );
  NOR3_X1 U11033 ( .A1(n8692), .A2(n10389), .A3(n10620), .ZN(n8693) );
  XNOR2_X1 U11034 ( .A(n14459), .B(n13672), .ZN(n10386) );
  NAND4_X1 U11035 ( .A1(n10949), .A2(n8693), .A3(n10386), .A4(n10474), .ZN(
        n8694) );
  OR4_X1 U11036 ( .A1(n11099), .A2(n10635), .A3(n10625), .A4(n8694), .ZN(n8695) );
  NOR2_X1 U11037 ( .A1(n11104), .A2(n8695), .ZN(n8696) );
  XNOR2_X1 U11038 ( .A(n11621), .B(n13666), .ZN(n11226) );
  NAND3_X1 U11039 ( .A1(n13972), .A2(n8696), .A3(n11226), .ZN(n8698) );
  XNOR2_X1 U11040 ( .A(n14360), .B(n14366), .ZN(n11463) );
  NAND2_X1 U11041 ( .A1(n11452), .A2(n8697), .ZN(n11459) );
  OR4_X1 U11042 ( .A1(n8698), .A2(n11463), .A3(n11459), .A4(n11173), .ZN(n8699) );
  OR4_X1 U11043 ( .A1(n13917), .A2(n13950), .A3(n13934), .A4(n8699), .ZN(n8700) );
  INV_X1 U11044 ( .A(n13659), .ZN(n13850) );
  XNOR2_X1 U11045 ( .A(n14028), .B(n13850), .ZN(n13831) );
  XNOR2_X1 U11046 ( .A(n13781), .B(n13655), .ZN(n8701) );
  NAND2_X1 U11047 ( .A1(n10849), .A2(n9272), .ZN(n8706) );
  INV_X1 U11048 ( .A(n8706), .ZN(n9825) );
  AND2_X1 U11049 ( .A1(n13773), .A2(n6454), .ZN(n8719) );
  INV_X1 U11050 ( .A(n8719), .ZN(n8703) );
  OR3_X1 U11051 ( .A1(n8703), .A2(n13776), .A3(n8705), .ZN(n8710) );
  INV_X1 U11052 ( .A(n13776), .ZN(n8720) );
  AND2_X1 U11053 ( .A1(n8705), .A2(n8706), .ZN(n8715) );
  NAND4_X1 U11054 ( .A1(n8703), .A2(n8720), .A3(n8715), .A4(n13773), .ZN(n8709) );
  OR2_X1 U11055 ( .A1(n13773), .A2(n6453), .ZN(n8716) );
  XNOR2_X1 U11056 ( .A(n8716), .B(n8705), .ZN(n8707) );
  NAND4_X1 U11057 ( .A1(n8707), .A2(n14088), .A3(n13776), .A4(n8706), .ZN(
        n8708) );
  NAND3_X1 U11058 ( .A1(n8710), .A2(n8709), .A3(n8708), .ZN(n8711) );
  NAND2_X1 U11059 ( .A1(n8714), .A2(n8713), .ZN(n8725) );
  OAI21_X1 U11060 ( .B1(n8716), .B2(n8720), .A(n8715), .ZN(n8718) );
  NAND2_X1 U11061 ( .A1(n8726), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8722) );
  INV_X1 U11062 ( .A(n9821), .ZN(n9085) );
  NAND2_X1 U11063 ( .A1(n9085), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11243) );
  INV_X1 U11064 ( .A(n11243), .ZN(n8723) );
  OAI21_X1 U11065 ( .B1(n8725), .B2(n8724), .A(n8723), .ZN(n8744) );
  INV_X1 U11066 ( .A(n8728), .ZN(n8729) );
  NAND2_X1 U11067 ( .A1(n8735), .A2(n8731), .ZN(n8738) );
  NAND2_X1 U11068 ( .A1(n8738), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8732) );
  MUX2_X1 U11069 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8732), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n8733) );
  INV_X1 U11070 ( .A(n8735), .ZN(n8736) );
  NAND2_X1 U11071 ( .A1(n8736), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8737) );
  MUX2_X1 U11072 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8737), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n8739) );
  NAND2_X1 U11073 ( .A1(n10062), .A2(n10586), .ZN(n9692) );
  INV_X1 U11074 ( .A(n14132), .ZN(n9424) );
  INV_X1 U11075 ( .A(n8741), .ZN(n9427) );
  NAND3_X1 U11076 ( .A1(n10153), .A2(n9424), .A3(n13954), .ZN(n8742) );
  OAI211_X1 U11077 ( .C1(n14137), .C2(n11243), .A(n8742), .B(P1_B_REG_SCAN_IN), 
        .ZN(n8743) );
  NAND2_X1 U11078 ( .A1(n8744), .A2(n8743), .ZN(P1_U3242) );
  INV_X1 U11079 ( .A(n8745), .ZN(n8746) );
  INV_X1 U11080 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12077) );
  XNOR2_X1 U11081 ( .A(n12077), .B(P2_DATAO_REG_30__SCAN_IN), .ZN(n8757) );
  OAI22_X1 U11082 ( .A1(n8758), .A2(n8757), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(n12132), .ZN(n8749) );
  XNOR2_X1 U11083 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n8748) );
  XNOR2_X1 U11084 ( .A(n8749), .B(n8748), .ZN(n12876) );
  NAND2_X1 U11085 ( .A1(n12876), .A2(n8761), .ZN(n8750) );
  INV_X1 U11086 ( .A(SI_31_), .ZN(n12871) );
  NAND2_X1 U11087 ( .A1(n6459), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n8754) );
  NAND2_X1 U11088 ( .A1(n7541), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n8753) );
  NAND2_X1 U11089 ( .A1(n7527), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n8752) );
  AND3_X1 U11090 ( .A1(n8754), .A2(n8753), .A3(n8752), .ZN(n8755) );
  NAND2_X1 U11091 ( .A1(n8756), .A2(n8755), .ZN(n12368) );
  INV_X1 U11092 ( .A(n12368), .ZN(n11630) );
  NAND2_X1 U11093 ( .A1(n12813), .A2(n11630), .ZN(n8921) );
  XNOR2_X1 U11094 ( .A(n8758), .B(n8757), .ZN(n12279) );
  INV_X1 U11095 ( .A(SI_30_), .ZN(n12281) );
  NOR2_X1 U11096 ( .A1(n8759), .A2(n12281), .ZN(n8760) );
  INV_X1 U11097 ( .A(n8926), .ZN(n12818) );
  OR2_X1 U11098 ( .A1(n12818), .A2(n12553), .ZN(n8915) );
  NAND2_X1 U11099 ( .A1(n8921), .A2(n8915), .ZN(n8932) );
  NAND2_X1 U11100 ( .A1(n12818), .A2(n12553), .ZN(n8785) );
  INV_X1 U11101 ( .A(n8785), .ZN(n8762) );
  INV_X1 U11102 ( .A(n8920), .ZN(n8783) );
  NAND2_X1 U11103 ( .A1(n11633), .A2(n12368), .ZN(n8786) );
  INV_X1 U11104 ( .A(n8786), .ZN(n8782) );
  AND2_X1 U11105 ( .A1(n12719), .A2(n12734), .ZN(n8874) );
  INV_X1 U11106 ( .A(n8874), .ZN(n8776) );
  INV_X1 U11107 ( .A(n11483), .ZN(n11475) );
  INV_X1 U11108 ( .A(n11251), .ZN(n8774) );
  AND2_X1 U11109 ( .A1(n6941), .A2(n8845), .ZN(n14283) );
  INV_X1 U11110 ( .A(n8763), .ZN(n8764) );
  NAND4_X1 U11111 ( .A1(n8764), .A2(n8793), .A3(n10230), .A4(n10214), .ZN(
        n8767) );
  INV_X1 U11112 ( .A(n9891), .ZN(n10039) );
  NAND2_X1 U11113 ( .A1(n12805), .A2(n10039), .ZN(n8791) );
  AND2_X1 U11114 ( .A1(n9893), .A2(n8791), .ZN(n9519) );
  NAND4_X1 U11115 ( .A1(n8765), .A2(n10145), .A3(n10522), .A4(n9519), .ZN(
        n8766) );
  NOR2_X1 U11116 ( .A1(n8767), .A2(n8766), .ZN(n8770) );
  NAND2_X1 U11117 ( .A1(n8769), .A2(n8768), .ZN(n10678) );
  NAND4_X1 U11118 ( .A1(n8770), .A2(n10802), .A3(n8829), .A4(n10678), .ZN(
        n8772) );
  INV_X1 U11119 ( .A(n8835), .ZN(n8771) );
  OR2_X1 U11120 ( .A1(n8836), .A2(n8771), .ZN(n14301) );
  NOR3_X1 U11121 ( .A1(n8772), .A2(n10999), .A3(n14301), .ZN(n8773) );
  NAND4_X1 U11122 ( .A1(n11396), .A2(n8774), .A3(n14283), .A4(n8773), .ZN(
        n8775) );
  NOR4_X1 U11123 ( .A1(n7729), .A2(n8776), .A3(n11475), .A4(n8775), .ZN(n8777)
         );
  INV_X1 U11124 ( .A(n12694), .ZN(n12687) );
  NAND4_X1 U11125 ( .A1(n12666), .A2(n12680), .A3(n8777), .A4(n12687), .ZN(
        n8778) );
  NOR4_X1 U11126 ( .A1(n12594), .A2(n12629), .A3(n12644), .A4(n8778), .ZN(
        n8780) );
  NAND4_X1 U11127 ( .A1(n12575), .A2(n8780), .A3(n8895), .A4(n8779), .ZN(n8781) );
  NOR4_X1 U11128 ( .A1(n8783), .A2(n8782), .A3(n8908), .A4(n8781), .ZN(n8784)
         );
  XNOR2_X1 U11129 ( .A(n8784), .B(n12543), .ZN(n8941) );
  NAND2_X1 U11130 ( .A1(n8786), .A2(n8785), .ZN(n8934) );
  INV_X1 U11131 ( .A(n8934), .ZN(n8917) );
  INV_X1 U11132 ( .A(n8787), .ZN(n8890) );
  INV_X1 U11133 ( .A(n8788), .ZN(n14913) );
  NAND3_X1 U11134 ( .A1(n8792), .A2(n8791), .A3(n10140), .ZN(n8795) );
  INV_X1 U11135 ( .A(n8789), .ZN(n8790) );
  AOI21_X1 U11136 ( .B1(n8792), .B2(n8791), .A(n8790), .ZN(n8794) );
  AOI21_X1 U11137 ( .B1(n14913), .B2(n8795), .A(n8798), .ZN(n8805) );
  NAND2_X1 U11138 ( .A1(n8801), .A2(n8796), .ZN(n8800) );
  NAND3_X1 U11139 ( .A1(n8798), .A2(n8797), .A3(n8802), .ZN(n8799) );
  MUX2_X1 U11140 ( .A(n8800), .B(n8799), .S(n9528), .Z(n8804) );
  MUX2_X1 U11141 ( .A(n8802), .B(n8801), .S(n9528), .Z(n8803) );
  MUX2_X1 U11142 ( .A(n8806), .B(n10213), .S(n8948), .Z(n8807) );
  NAND3_X1 U11143 ( .A1(n8811), .A2(n8808), .A3(n8813), .ZN(n8809) );
  NAND2_X1 U11144 ( .A1(n8809), .A2(n10423), .ZN(n8816) );
  NAND2_X1 U11145 ( .A1(n8811), .A2(n8810), .ZN(n8814) );
  INV_X1 U11146 ( .A(n10423), .ZN(n8812) );
  AOI21_X1 U11147 ( .B1(n8814), .B2(n8813), .A(n8812), .ZN(n8815) );
  MUX2_X1 U11148 ( .A(n8818), .B(n8817), .S(n9528), .Z(n8819) );
  OAI211_X1 U11149 ( .C1(n8820), .C2(n10673), .A(n10678), .B(n8819), .ZN(n8825) );
  NAND2_X1 U11150 ( .A1(n10790), .A2(n9528), .ZN(n8823) );
  NAND2_X1 U11151 ( .A1(n8821), .A2(n8948), .ZN(n8822) );
  MUX2_X1 U11152 ( .A(n8823), .B(n8822), .S(n10804), .Z(n8824) );
  NAND3_X1 U11153 ( .A1(n8825), .A2(n10802), .A3(n8824), .ZN(n8830) );
  MUX2_X1 U11154 ( .A(n8827), .B(n8826), .S(n9528), .Z(n8828) );
  NAND3_X1 U11155 ( .A1(n8830), .A2(n8829), .A3(n8828), .ZN(n8834) );
  NAND2_X1 U11156 ( .A1(n12376), .A2(n9528), .ZN(n8832) );
  NAND2_X1 U11157 ( .A1(n14305), .A2(n8948), .ZN(n8831) );
  MUX2_X1 U11158 ( .A(n8832), .B(n8831), .S(n10842), .Z(n8833) );
  AOI21_X1 U11159 ( .B1(n8834), .B2(n8833), .A(n14301), .ZN(n8844) );
  NAND2_X1 U11160 ( .A1(n8841), .A2(n8835), .ZN(n8839) );
  INV_X1 U11161 ( .A(n8836), .ZN(n8837) );
  NAND2_X1 U11162 ( .A1(n8840), .A2(n8837), .ZN(n8838) );
  MUX2_X1 U11163 ( .A(n8839), .B(n8838), .S(n8948), .Z(n8843) );
  MUX2_X1 U11164 ( .A(n8841), .B(n8840), .S(n9528), .Z(n8842) );
  INV_X1 U11165 ( .A(n8845), .ZN(n8846) );
  MUX2_X1 U11166 ( .A(n8847), .B(n8846), .S(n8948), .Z(n8848) );
  AOI21_X1 U11167 ( .B1(n8849), .B2(n14283), .A(n8848), .ZN(n8851) );
  OAI22_X1 U11168 ( .A1(n8851), .A2(n11251), .B1(n8948), .B2(n8850), .ZN(n8857) );
  INV_X1 U11169 ( .A(n8852), .ZN(n8854) );
  OAI21_X1 U11170 ( .B1(n8854), .B2(n8853), .A(n8860), .ZN(n8855) );
  AOI21_X1 U11171 ( .B1(n8855), .B2(n8862), .A(n9528), .ZN(n8856) );
  AOI21_X1 U11172 ( .B1(n8857), .B2(n11396), .A(n8856), .ZN(n8859) );
  INV_X1 U11173 ( .A(n8861), .ZN(n8858) );
  NOR2_X1 U11174 ( .A1(n8859), .A2(n8858), .ZN(n8864) );
  AOI21_X1 U11175 ( .B1(n8861), .B2(n8860), .A(n8948), .ZN(n8863) );
  OAI22_X1 U11176 ( .A1(n8864), .A2(n8863), .B1(n8948), .B2(n8862), .ZN(n8875)
         );
  INV_X1 U11177 ( .A(n8865), .ZN(n8866) );
  NOR2_X1 U11178 ( .A1(n8867), .A2(n8866), .ZN(n8870) );
  INV_X1 U11179 ( .A(n8870), .ZN(n8868) );
  NAND2_X1 U11180 ( .A1(n8868), .A2(n8876), .ZN(n8872) );
  OAI21_X1 U11181 ( .B1(n8870), .B2(n8874), .A(n8869), .ZN(n8871) );
  MUX2_X1 U11182 ( .A(n8872), .B(n8871), .S(n9528), .Z(n8873) );
  AOI21_X1 U11183 ( .B1(n8875), .B2(n8874), .A(n8873), .ZN(n8879) );
  MUX2_X1 U11184 ( .A(n8877), .B(n6947), .S(n9528), .Z(n8878) );
  NOR2_X1 U11185 ( .A1(n8879), .A2(n8878), .ZN(n8882) );
  NAND2_X1 U11186 ( .A1(n11652), .A2(n12677), .ZN(n8880) );
  MUX2_X1 U11187 ( .A(n8880), .B(n12661), .S(n8948), .Z(n8881) );
  OAI211_X1 U11188 ( .C1(n8882), .C2(n12694), .A(n12680), .B(n8881), .ZN(n8884) );
  MUX2_X1 U11189 ( .A(n12662), .B(n12663), .S(n9528), .Z(n8883) );
  NAND3_X1 U11190 ( .A1(n8884), .A2(n12666), .A3(n8883), .ZN(n8888) );
  MUX2_X1 U11191 ( .A(n8886), .B(n8885), .S(n8948), .Z(n8887) );
  AOI21_X1 U11192 ( .B1(n8888), .B2(n8887), .A(n12644), .ZN(n8889) );
  AOI21_X1 U11193 ( .B1(n8890), .B2(n9528), .A(n8889), .ZN(n8897) );
  INV_X1 U11194 ( .A(n8891), .ZN(n8894) );
  XNOR2_X1 U11195 ( .A(n8892), .B(n8948), .ZN(n8893) );
  OAI21_X1 U11196 ( .B1(n12629), .B2(n8894), .A(n8893), .ZN(n8896) );
  OAI211_X1 U11197 ( .C1(n8897), .C2(n12629), .A(n8896), .B(n8895), .ZN(n8901)
         );
  INV_X1 U11198 ( .A(n12311), .ZN(n12836) );
  NAND2_X1 U11199 ( .A1(n12836), .A2(n12627), .ZN(n8898) );
  MUX2_X1 U11200 ( .A(n8899), .B(n8898), .S(n9528), .Z(n8900) );
  NAND3_X1 U11201 ( .A1(n8901), .A2(n7935), .A3(n8900), .ZN(n8905) );
  MUX2_X1 U11202 ( .A(n8903), .B(n8902), .S(n8948), .Z(n8904) );
  AOI21_X1 U11203 ( .B1(n8905), .B2(n8904), .A(n7859), .ZN(n8907) );
  NOR3_X1 U11204 ( .A1(n11677), .A2(n12567), .A3(n9528), .ZN(n8906) );
  OAI21_X1 U11205 ( .B1(n8907), .B2(n8906), .A(n12575), .ZN(n8914) );
  INV_X1 U11206 ( .A(n8908), .ZN(n8913) );
  NAND2_X1 U11207 ( .A1(n8909), .A2(n8910), .ZN(n8911) );
  MUX2_X1 U11208 ( .A(n8911), .B(n8910), .S(n8948), .Z(n8912) );
  NAND3_X1 U11209 ( .A1(n8914), .A2(n8913), .A3(n8912), .ZN(n8918) );
  NAND4_X1 U11210 ( .A1(n8918), .A2(n9528), .A3(n8915), .A4(n8925), .ZN(n8916)
         );
  NAND2_X1 U11211 ( .A1(n8917), .A2(n8916), .ZN(n8922) );
  AOI21_X1 U11212 ( .B1(n8918), .B2(n8927), .A(n9528), .ZN(n8919) );
  AOI22_X1 U11213 ( .A1(n8922), .A2(n8921), .B1(n8920), .B2(n8919), .ZN(n8924)
         );
  OAI21_X1 U11214 ( .B1(n8924), .B2(n9755), .A(n8923), .ZN(n8940) );
  INV_X1 U11215 ( .A(n8925), .ZN(n8930) );
  INV_X1 U11216 ( .A(n8932), .ZN(n8933) );
  OAI22_X1 U11217 ( .A1(n8935), .A2(n8934), .B1(n11633), .B2(n8933), .ZN(n8936) );
  XNOR2_X1 U11218 ( .A(n8936), .B(n12533), .ZN(n8939) );
  INV_X1 U11219 ( .A(n8937), .ZN(n8938) );
  OR2_X1 U11220 ( .A1(n9527), .A2(P3_U3151), .ZN(n10943) );
  NOR3_X1 U11221 ( .A1(n9300), .A2(n8942), .A3(n12880), .ZN(n8944) );
  OAI21_X1 U11222 ( .B1(n10943), .B2(n10535), .A(P3_B_REG_SCAN_IN), .ZN(n8943)
         );
  OR2_X1 U11223 ( .A1(n8944), .A2(n8943), .ZN(n8945) );
  NAND2_X1 U11224 ( .A1(n8946), .A2(n8948), .ZN(n10032) );
  NAND2_X1 U11225 ( .A1(n10032), .A2(n10034), .ZN(n8954) );
  NAND2_X1 U11226 ( .A1(n8949), .A2(n7977), .ZN(n8950) );
  OAI211_X1 U11227 ( .C1(n10535), .C2(n8951), .A(n8950), .B(n10031), .ZN(n8952) );
  INV_X1 U11228 ( .A(n8952), .ZN(n8953) );
  AOI21_X1 U11229 ( .B1(n12866), .B2(n8954), .A(n8953), .ZN(n8958) );
  NAND2_X1 U11230 ( .A1(n8963), .A2(n8962), .ZN(P3_U3488) );
  INV_X1 U11231 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n9026) );
  NOR2_X2 U11232 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n9018) );
  AND2_X2 U11233 ( .A1(n9018), .A2(n8966), .ZN(n9006) );
  NAND2_X1 U11234 ( .A1(n8971), .A2(n9138), .ZN(n9133) );
  NAND2_X1 U11235 ( .A1(n8982), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8973) );
  MUX2_X1 U11236 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8973), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8979) );
  NOR2_X1 U11237 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), 
        .ZN(n8977) );
  NOR2_X1 U11238 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), 
        .ZN(n8976) );
  NOR2_X1 U11239 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), 
        .ZN(n8975) );
  NAND4_X1 U11240 ( .A1(n8977), .A2(n8976), .A3(n8975), .A4(n8974), .ZN(n9140)
         );
  NAND2_X1 U11241 ( .A1(n8987), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8981) );
  MUX2_X1 U11242 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8981), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8983) );
  INV_X1 U11243 ( .A(n8984), .ZN(n8985) );
  NAND2_X1 U11244 ( .A1(n8985), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8986) );
  MUX2_X1 U11245 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8986), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n8988) );
  NOR2_X1 U11246 ( .A1(n11375), .A2(n11269), .ZN(n8989) );
  NAND2_X1 U11247 ( .A1(n9309), .A2(n8989), .ZN(n9331) );
  NAND2_X1 U11248 ( .A1(n9136), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8991) );
  INV_X1 U11249 ( .A(n11219), .ZN(n8992) );
  NOR2_X1 U11250 ( .A1(n9331), .A2(n8992), .ZN(n9143) );
  INV_X1 U11251 ( .A(n8993), .ZN(n9122) );
  INV_X1 U11252 ( .A(n9292), .ZN(n8994) );
  AND2_X1 U11253 ( .A1(n6461), .A2(P1_U3086), .ZN(n14127) );
  INV_X2 U11254 ( .A(n14127), .ZN(n14135) );
  INV_X2 U11255 ( .A(n11242), .ZN(n12134) );
  OAI222_X1 U11256 ( .A1(n14135), .A2(n8995), .B1(n12134), .B2(n9643), .C1(
        n13712), .C2(P1_U3086), .ZN(P1_U3352) );
  OAI222_X1 U11257 ( .A1(n14135), .A2(n8996), .B1(n12134), .B2(n9374), .C1(
        n9212), .C2(P1_U3086), .ZN(P1_U3354) );
  NAND2_X1 U11258 ( .A1(n6461), .A2(P3_U3151), .ZN(n12870) );
  INV_X1 U11259 ( .A(SI_5_), .ZN(n9000) );
  NOR2_X1 U11260 ( .A1(n9335), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12875) );
  INV_X1 U11261 ( .A(n8998), .ZN(n8999) );
  OAI222_X1 U11262 ( .A1(P3_U3151), .A2(n14802), .B1(n12870), .B2(n9000), .C1(
        n12886), .C2(n8999), .ZN(P3_U3290) );
  OAI222_X1 U11263 ( .A1(P1_U3086), .A2(n13696), .B1(n12134), .B2(n9395), .C1(
        n9001), .C2(n14135), .ZN(P1_U3353) );
  INV_X1 U11264 ( .A(n9002), .ZN(n9004) );
  INV_X1 U11265 ( .A(SI_2_), .ZN(n9003) );
  OAI222_X1 U11266 ( .A1(n6462), .A2(P3_U3151), .B1(n12886), .B2(n9004), .C1(
        n9003), .C2(n12883), .ZN(P3_U3293) );
  INV_X1 U11267 ( .A(n9648), .ZN(n9010) );
  OAI222_X1 U11268 ( .A1(n14135), .A2(n9005), .B1(n12134), .B2(n9010), .C1(
        P1_U3086), .C2(n9219), .ZN(P1_U3351) );
  NOR2_X1 U11269 ( .A1(n9335), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13519) );
  INV_X2 U11270 ( .A(n13519), .ZN(n13523) );
  INV_X1 U11271 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n9007) );
  AND2_X1 U11272 ( .A1(n9006), .A2(n9007), .ZN(n9037) );
  INV_X1 U11273 ( .A(n9037), .ZN(n9024) );
  NAND2_X1 U11274 ( .A1(n9024), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9008) );
  XNOR2_X1 U11275 ( .A(n9008), .B(P2_IR_REG_4__SCAN_IN), .ZN(n13084) );
  INV_X1 U11276 ( .A(n13084), .ZN(n9009) );
  OAI222_X1 U11277 ( .A1(n13523), .A2(n9011), .B1(n13526), .B2(n9010), .C1(
        P2_U3088), .C2(n9009), .ZN(P2_U3323) );
  INV_X1 U11278 ( .A(SI_7_), .ZN(n9014) );
  INV_X1 U11279 ( .A(n9012), .ZN(n9013) );
  OAI222_X1 U11280 ( .A1(P3_U3151), .A2(n14838), .B1(n12870), .B2(n9014), .C1(
        n12886), .C2(n9013), .ZN(P3_U3288) );
  OAI222_X1 U11281 ( .A1(P3_U3151), .A2(n14855), .B1(n12870), .B2(n9016), .C1(
        n12886), .C2(n9015), .ZN(P3_U3287) );
  INV_X1 U11282 ( .A(n9621), .ZN(n9048) );
  INV_X1 U11283 ( .A(n9222), .ZN(n9251) );
  OAI222_X1 U11284 ( .A1(n14135), .A2(n9017), .B1(n12134), .B2(n9048), .C1(
        P1_U3086), .C2(n9251), .ZN(P1_U3350) );
  INV_X1 U11285 ( .A(n9467), .ZN(n9474) );
  OAI222_X1 U11286 ( .A1(n14135), .A2(n6819), .B1(n12134), .B2(n9847), .C1(
        n9474), .C2(P1_U3086), .ZN(P1_U3349) );
  NOR2_X1 U11287 ( .A1(n9019), .A2(n9884), .ZN(n9020) );
  MUX2_X1 U11288 ( .A(n9884), .B(n9020), .S(P2_IR_REG_2__SCAN_IN), .Z(n9021)
         );
  INV_X1 U11289 ( .A(n9021), .ZN(n9023) );
  INV_X1 U11290 ( .A(n9006), .ZN(n9022) );
  NAND2_X1 U11291 ( .A1(n9023), .A2(n9022), .ZN(n14556) );
  OAI222_X1 U11292 ( .A1(n13526), .A2(n9395), .B1(n14556), .B2(P2_U3088), .C1(
        n9396), .C2(n13523), .ZN(P2_U3325) );
  INV_X1 U11293 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n9025) );
  NAND2_X1 U11294 ( .A1(n9065), .A2(n9025), .ZN(n9046) );
  INV_X1 U11295 ( .A(n9046), .ZN(n9027) );
  NAND2_X1 U11296 ( .A1(n9027), .A2(n9026), .ZN(n9062) );
  NAND2_X1 U11297 ( .A1(n9062), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9028) );
  XNOR2_X1 U11298 ( .A(n9028), .B(P2_IR_REG_7__SCAN_IN), .ZN(n14577) );
  INV_X1 U11299 ( .A(n14577), .ZN(n9030) );
  OAI222_X1 U11300 ( .A1(n13526), .A2(n9855), .B1(n9030), .B2(P2_U3088), .C1(
        n9029), .C2(n13523), .ZN(P2_U3320) );
  NAND2_X1 U11301 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n9031) );
  MUX2_X1 U11302 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9031), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n9033) );
  INV_X1 U11303 ( .A(n9019), .ZN(n9032) );
  NAND2_X1 U11304 ( .A1(n9033), .A2(n9032), .ZN(n9375) );
  OAI222_X1 U11305 ( .A1(n13526), .A2(n9374), .B1(n9375), .B2(P2_U3088), .C1(
        n9377), .C2(n13523), .ZN(P2_U3326) );
  NAND2_X1 U11306 ( .A1(n9046), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9034) );
  XNOR2_X1 U11307 ( .A(n9034), .B(P2_IR_REG_6__SCAN_IN), .ZN(n13112) );
  INV_X1 U11308 ( .A(n13112), .ZN(n9130) );
  INV_X1 U11309 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9035) );
  OAI222_X1 U11310 ( .A1(n13526), .A2(n9847), .B1(n9130), .B2(P2_U3088), .C1(
        n9035), .C2(n13523), .ZN(P2_U3321) );
  NOR2_X1 U11311 ( .A1(n9006), .A2(n9884), .ZN(n9036) );
  MUX2_X1 U11312 ( .A(n9884), .B(n9036), .S(P2_IR_REG_3__SCAN_IN), .Z(n9038)
         );
  NOR2_X1 U11313 ( .A1(n9038), .A2(n9037), .ZN(n13070) );
  INV_X1 U11314 ( .A(n13070), .ZN(n9126) );
  OAI222_X1 U11315 ( .A1(n13526), .A2(n9643), .B1(n9126), .B2(P2_U3088), .C1(
        n9039), .C2(n13523), .ZN(P2_U3324) );
  INV_X1 U11316 ( .A(SI_9_), .ZN(n9042) );
  INV_X1 U11317 ( .A(n9040), .ZN(n9041) );
  OAI222_X1 U11318 ( .A1(P3_U3151), .A2(n14875), .B1(n12870), .B2(n9042), .C1(
        n12886), .C2(n9041), .ZN(P3_U3286) );
  INV_X1 U11319 ( .A(n9506), .ZN(n9514) );
  OAI222_X1 U11320 ( .A1(n14135), .A2(n9043), .B1(n12134), .B2(n9855), .C1(
        n9514), .C2(P1_U3086), .ZN(P1_U3348) );
  NAND2_X1 U11321 ( .A1(n9044), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9045) );
  MUX2_X1 U11322 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9045), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n9047) );
  NAND2_X1 U11323 ( .A1(n9047), .A2(n9046), .ZN(n9160) );
  OAI222_X1 U11324 ( .A1(n13523), .A2(n9049), .B1(n13526), .B2(n9048), .C1(
        P2_U3088), .C2(n9160), .ZN(P2_U3322) );
  OAI222_X1 U11325 ( .A1(n12886), .A2(n9051), .B1(n12883), .B2(n9050), .C1(
        P3_U3151), .C2(n6465), .ZN(P3_U3294) );
  OAI222_X1 U11326 ( .A1(n12886), .A2(n9053), .B1(n12870), .B2(n9052), .C1(
        P3_U3151), .C2(n14819), .ZN(P3_U3289) );
  INV_X1 U11327 ( .A(SI_3_), .ZN(n9056) );
  INV_X1 U11328 ( .A(n9054), .ZN(n9055) );
  OAI222_X1 U11329 ( .A1(P3_U3151), .A2(n14766), .B1(n12870), .B2(n9056), .C1(
        n12886), .C2(n9055), .ZN(P3_U3292) );
  INV_X1 U11330 ( .A(SI_4_), .ZN(n9059) );
  INV_X1 U11331 ( .A(n9057), .ZN(n9058) );
  OAI222_X1 U11332 ( .A1(P3_U3151), .A2(n14783), .B1(n12870), .B2(n9059), .C1(
        n12886), .C2(n9058), .ZN(P3_U3291) );
  OAI222_X1 U11333 ( .A1(P3_U3151), .A2(n10920), .B1(n12883), .B2(n9061), .C1(
        n12886), .C2(n9060), .ZN(P3_U3285) );
  NAND2_X1 U11334 ( .A1(n9070), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9063) );
  MUX2_X1 U11335 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9063), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n9066) );
  NAND2_X1 U11336 ( .A1(n9065), .A2(n9064), .ZN(n9077) );
  NAND2_X1 U11337 ( .A1(n9066), .A2(n9077), .ZN(n10066) );
  OAI222_X1 U11338 ( .A1(n13526), .A2(n10064), .B1(n10066), .B2(P2_U3088), 
        .C1(n10067), .C2(n13523), .ZN(P2_U3318) );
  INV_X1 U11339 ( .A(n9952), .ZN(n9072) );
  INV_X1 U11340 ( .A(n9477), .ZN(n9496) );
  OAI222_X1 U11341 ( .A1(n14135), .A2(n9067), .B1(n12134), .B2(n9072), .C1(
        P1_U3086), .C2(n9496), .ZN(P1_U3347) );
  NAND2_X1 U11342 ( .A1(n9068), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9069) );
  MUX2_X1 U11343 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9069), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n9071) );
  NAND2_X1 U11344 ( .A1(n9071), .A2(n9070), .ZN(n9151) );
  OAI222_X1 U11345 ( .A1(n13523), .A2(n9073), .B1(n13526), .B2(n9072), .C1(
        P2_U3088), .C2(n9151), .ZN(P2_U3319) );
  INV_X1 U11346 ( .A(n9602), .ZN(n9611) );
  OAI222_X1 U11347 ( .A1(n14135), .A2(n9074), .B1(n12134), .B2(n10064), .C1(
        n9611), .C2(P1_U3086), .ZN(P1_U3346) );
  OAI222_X1 U11348 ( .A1(P3_U3151), .A2(n11086), .B1(n12883), .B2(n9076), .C1(
        n12886), .C2(n9075), .ZN(P3_U3284) );
  NAND2_X1 U11349 ( .A1(n9077), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9078) );
  XNOR2_X1 U11350 ( .A(n9078), .B(P2_IR_REG_10__SCAN_IN), .ZN(n14593) );
  INV_X1 U11351 ( .A(n14593), .ZN(n9080) );
  OAI222_X1 U11352 ( .A1(n13526), .A2(n10121), .B1(n9080), .B2(P2_U3088), .C1(
        n9079), .C2(n13523), .ZN(P2_U3317) );
  INV_X1 U11353 ( .A(n9580), .ZN(n9584) );
  OAI222_X1 U11354 ( .A1(n14135), .A2(n9081), .B1(n12134), .B2(n10121), .C1(
        n9584), .C2(P1_U3086), .ZN(P1_U3345) );
  OAI222_X1 U11355 ( .A1(P3_U3151), .A2(n12387), .B1(n12883), .B2(n9083), .C1(
        n12886), .C2(n9082), .ZN(P3_U3283) );
  NAND2_X1 U11356 ( .A1(n10305), .A2(n11243), .ZN(n9173) );
  OAI21_X1 U11357 ( .B1(n9085), .B2(n9814), .A(n9084), .ZN(n9171) );
  NAND2_X1 U11358 ( .A1(n9173), .A2(n9171), .ZN(n14456) );
  INV_X1 U11359 ( .A(n14456), .ZN(n13725) );
  NOR2_X1 U11360 ( .A1(n13725), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U11361 ( .A(n10356), .ZN(n9116) );
  NAND2_X1 U11363 ( .A1(n9197), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9087) );
  XNOR2_X1 U11364 ( .A(n9087), .B(P2_IR_REG_11__SCAN_IN), .ZN(n13132) );
  AOI22_X1 U11365 ( .A1(n13132), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n13519), .ZN(n9088) );
  OAI21_X1 U11366 ( .B1(n9116), .B2(n13526), .A(n9088), .ZN(P2_U3316) );
  INV_X1 U11367 ( .A(n12867), .ZN(n9090) );
  NOR2_X1 U11368 ( .A1(n9090), .A2(n9089), .ZN(n9092) );
  CLKBUF_X1 U11369 ( .A(n9092), .Z(n9114) );
  INV_X1 U11370 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n9091) );
  NOR2_X1 U11371 ( .A1(n9114), .A2(n9091), .ZN(P3_U3255) );
  INV_X1 U11372 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n15111) );
  NOR2_X1 U11373 ( .A1(n9114), .A2(n15111), .ZN(P3_U3261) );
  INV_X1 U11374 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n9093) );
  NOR2_X1 U11375 ( .A1(n9114), .A2(n9093), .ZN(P3_U3262) );
  INV_X1 U11376 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n9094) );
  NOR2_X1 U11377 ( .A1(n9092), .A2(n9094), .ZN(P3_U3258) );
  INV_X1 U11378 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n9095) );
  NOR2_X1 U11379 ( .A1(n9092), .A2(n9095), .ZN(P3_U3260) );
  INV_X1 U11380 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n9096) );
  NOR2_X1 U11381 ( .A1(n9114), .A2(n9096), .ZN(P3_U3256) );
  INV_X1 U11382 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n9097) );
  NOR2_X1 U11383 ( .A1(n9092), .A2(n9097), .ZN(P3_U3240) );
  INV_X1 U11384 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n9098) );
  NOR2_X1 U11385 ( .A1(n9114), .A2(n9098), .ZN(P3_U3254) );
  INV_X1 U11386 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n9099) );
  NOR2_X1 U11387 ( .A1(n9114), .A2(n9099), .ZN(P3_U3263) );
  INV_X1 U11388 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n9100) );
  NOR2_X1 U11389 ( .A1(n9114), .A2(n9100), .ZN(P3_U3259) );
  INV_X1 U11390 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n9101) );
  NOR2_X1 U11391 ( .A1(n9114), .A2(n9101), .ZN(P3_U3246) );
  INV_X1 U11392 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n9102) );
  NOR2_X1 U11393 ( .A1(n9092), .A2(n9102), .ZN(P3_U3245) );
  INV_X1 U11394 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n9103) );
  NOR2_X1 U11395 ( .A1(n9092), .A2(n9103), .ZN(P3_U3244) );
  INV_X1 U11396 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n15099) );
  NOR2_X1 U11397 ( .A1(n9092), .A2(n15099), .ZN(P3_U3243) );
  INV_X1 U11398 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n15076) );
  NOR2_X1 U11399 ( .A1(n9092), .A2(n15076), .ZN(P3_U3242) );
  INV_X1 U11400 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n15096) );
  NOR2_X1 U11401 ( .A1(n9092), .A2(n15096), .ZN(P3_U3241) );
  INV_X1 U11402 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n9104) );
  NOR2_X1 U11403 ( .A1(n9114), .A2(n9104), .ZN(P3_U3247) );
  INV_X1 U11404 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n15084) );
  NOR2_X1 U11405 ( .A1(n9092), .A2(n15084), .ZN(P3_U3239) );
  INV_X1 U11406 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n9105) );
  NOR2_X1 U11407 ( .A1(n9092), .A2(n9105), .ZN(P3_U3238) );
  INV_X1 U11408 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n9106) );
  NOR2_X1 U11409 ( .A1(n9114), .A2(n9106), .ZN(P3_U3257) );
  INV_X1 U11410 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n9107) );
  NOR2_X1 U11411 ( .A1(n9092), .A2(n9107), .ZN(P3_U3236) );
  INV_X1 U11412 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n9108) );
  NOR2_X1 U11413 ( .A1(n9114), .A2(n9108), .ZN(P3_U3235) );
  INV_X1 U11414 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n9109) );
  NOR2_X1 U11415 ( .A1(n9114), .A2(n9109), .ZN(P3_U3234) );
  INV_X1 U11416 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n15100) );
  NOR2_X1 U11417 ( .A1(n9114), .A2(n15100), .ZN(P3_U3253) );
  INV_X1 U11418 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n9110) );
  NOR2_X1 U11419 ( .A1(n9114), .A2(n9110), .ZN(P3_U3249) );
  INV_X1 U11420 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n9111) );
  NOR2_X1 U11421 ( .A1(n9114), .A2(n9111), .ZN(P3_U3248) );
  INV_X1 U11422 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n9112) );
  NOR2_X1 U11423 ( .A1(n9114), .A2(n9112), .ZN(P3_U3252) );
  INV_X1 U11424 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n9113) );
  NOR2_X1 U11425 ( .A1(n9114), .A2(n9113), .ZN(P3_U3251) );
  INV_X1 U11426 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n15095) );
  NOR2_X1 U11427 ( .A1(n9114), .A2(n15095), .ZN(P3_U3250) );
  INV_X1 U11428 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n9115) );
  NOR2_X1 U11429 ( .A1(n9114), .A2(n9115), .ZN(P3_U3237) );
  INV_X1 U11430 ( .A(n9741), .ZN(n9736) );
  OAI222_X1 U11431 ( .A1(n15130), .A2(n14135), .B1(P1_U3086), .B2(n9736), .C1(
        n12134), .C2(n9116), .ZN(P1_U3344) );
  NAND2_X1 U11432 ( .A1(n11373), .A2(P1_B_REG_SCAN_IN), .ZN(n9117) );
  MUX2_X1 U11433 ( .A(n9117), .B(P1_B_REG_SCAN_IN), .S(n11270), .Z(n9118) );
  INV_X1 U11434 ( .A(n11515), .ZN(n9121) );
  INV_X1 U11435 ( .A(n10305), .ZN(n9119) );
  INV_X1 U11436 ( .A(n14500), .ZN(n14499) );
  NAND2_X1 U11437 ( .A1(n11515), .A2(n11373), .ZN(n9255) );
  OAI22_X1 U11438 ( .A1(n14499), .A2(P1_D_REG_1__SCAN_IN), .B1(n9122), .B2(
        n9255), .ZN(n9120) );
  INV_X1 U11439 ( .A(n9120), .ZN(P1_U3446) );
  OR2_X1 U11440 ( .A1(n11270), .A2(n9121), .ZN(n9269) );
  OAI22_X1 U11441 ( .A1(n14499), .A2(P1_D_REG_0__SCAN_IN), .B1(n9122), .B2(
        n9269), .ZN(n9123) );
  INV_X1 U11442 ( .A(n9123), .ZN(P1_U3445) );
  INV_X1 U11443 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n13113) );
  INV_X1 U11444 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9124) );
  MUX2_X1 U11445 ( .A(n9124), .B(P2_REG2_REG_2__SCAN_IN), .S(n14556), .Z(
        n14566) );
  INV_X1 U11446 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10335) );
  XNOR2_X1 U11447 ( .A(n9375), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n14552) );
  NAND3_X1 U11448 ( .A1(n14552), .A2(P2_IR_REG_0__SCAN_IN), .A3(
        P2_REG2_REG_0__SCAN_IN), .ZN(n14550) );
  OAI21_X1 U11449 ( .B1(n10335), .B2(n9375), .A(n14550), .ZN(n14567) );
  NAND2_X1 U11450 ( .A1(n14566), .A2(n14567), .ZN(n14565) );
  INV_X1 U11451 ( .A(n14556), .ZN(n9125) );
  NAND2_X1 U11452 ( .A1(n9125), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n13072) );
  INV_X1 U11453 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n14652) );
  MUX2_X1 U11454 ( .A(n14652), .B(P2_REG2_REG_3__SCAN_IN), .S(n13070), .Z(
        n13073) );
  AOI21_X1 U11455 ( .B1(n14565), .B2(n13072), .A(n13073), .ZN(n13071) );
  NOR2_X1 U11456 ( .A1(n9126), .A2(n14652), .ZN(n13083) );
  INV_X1 U11457 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10202) );
  MUX2_X1 U11458 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n10202), .S(n13084), .Z(
        n9127) );
  OAI21_X1 U11459 ( .B1(n13071), .B2(n13083), .A(n9127), .ZN(n13101) );
  NAND2_X1 U11460 ( .A1(n13084), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n13100) );
  INV_X1 U11461 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n9128) );
  MUX2_X1 U11462 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n9128), .S(n9160), .Z(n13099) );
  AOI21_X1 U11463 ( .B1(n13101), .B2(n13100), .A(n13099), .ZN(n13098) );
  NOR2_X1 U11464 ( .A1(n9160), .A2(n9128), .ZN(n13111) );
  MUX2_X1 U11465 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n13113), .S(n13112), .Z(
        n9129) );
  OAI21_X1 U11466 ( .B1(n13098), .B2(n13111), .A(n9129), .ZN(n13118) );
  OAI21_X1 U11467 ( .B1(n13113), .B2(n9130), .A(n13118), .ZN(n14581) );
  INV_X1 U11468 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n9131) );
  MUX2_X1 U11469 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n9131), .S(n14577), .Z(
        n14580) );
  NAND2_X1 U11470 ( .A1(n14581), .A2(n14580), .ZN(n14578) );
  NAND2_X1 U11471 ( .A1(n14577), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9146) );
  INV_X1 U11472 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n9132) );
  MUX2_X1 U11473 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n9132), .S(n9151), .Z(n9145)
         );
  AOI21_X1 U11474 ( .B1(n14578), .B2(n9146), .A(n9145), .ZN(n9186) );
  NAND2_X1 U11475 ( .A1(n9133), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9134) );
  MUX2_X1 U11476 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9134), .S(
        P2_IR_REG_22__SCAN_IN), .Z(n9135) );
  NAND2_X2 U11477 ( .A1(n9136), .A2(n9135), .ZN(n12063) );
  AOI21_X1 U11478 ( .B1(n9373), .B2(n11219), .A(n11898), .ZN(n9142) );
  OR2_X1 U11479 ( .A1(n9143), .A2(n9142), .ZN(n9148) );
  NOR2_X1 U11480 ( .A1(n9144), .A2(P2_U3088), .ZN(n13518) );
  NAND2_X1 U11481 ( .A1(n9148), .A2(n13518), .ZN(n9164) );
  NAND3_X1 U11482 ( .A1(n14578), .A2(n9146), .A3(n9145), .ZN(n9147) );
  NAND2_X1 U11483 ( .A1(n14579), .A2(n9147), .ZN(n9170) );
  INV_X1 U11484 ( .A(n9151), .ZN(n9953) );
  NAND2_X1 U11485 ( .A1(n9148), .A2(n9144), .ZN(n14557) );
  OR2_X1 U11486 ( .A1(n14557), .A2(P2_U3088), .ZN(n14618) );
  INV_X1 U11487 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n9149) );
  NAND2_X1 U11488 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n9977) );
  OAI21_X1 U11489 ( .B1(n14602), .B2(n9149), .A(n9977), .ZN(n9150) );
  AOI21_X1 U11490 ( .B1(n9953), .B2(n14594), .A(n9150), .ZN(n9169) );
  INV_X1 U11491 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n14742) );
  MUX2_X1 U11492 ( .A(n14742), .B(P2_REG1_REG_8__SCAN_IN), .S(n9151), .Z(n9167) );
  INV_X1 U11493 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9152) );
  XNOR2_X1 U11494 ( .A(n13070), .B(n9152), .ZN(n13069) );
  XNOR2_X1 U11495 ( .A(n14556), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n14561) );
  XNOR2_X1 U11496 ( .A(n9375), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n14541) );
  NAND2_X1 U11497 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n14545) );
  INV_X1 U11498 ( .A(n14545), .ZN(n9153) );
  NAND2_X1 U11499 ( .A1(n14541), .A2(n9153), .ZN(n14542) );
  INV_X1 U11500 ( .A(n9375), .ZN(n14547) );
  NAND2_X1 U11501 ( .A1(n14547), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9154) );
  NAND2_X1 U11502 ( .A1(n14542), .A2(n9154), .ZN(n14560) );
  NAND2_X1 U11503 ( .A1(n14561), .A2(n14560), .ZN(n14559) );
  INV_X1 U11504 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9155) );
  OR2_X1 U11505 ( .A1(n14556), .A2(n9155), .ZN(n9156) );
  NAND2_X1 U11506 ( .A1(n14559), .A2(n9156), .ZN(n13068) );
  NAND2_X1 U11507 ( .A1(n13069), .A2(n13068), .ZN(n13067) );
  NAND2_X1 U11508 ( .A1(n13070), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9157) );
  NAND2_X1 U11509 ( .A1(n13067), .A2(n9157), .ZN(n13081) );
  INV_X1 U11510 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9158) );
  XNOR2_X1 U11511 ( .A(n13084), .B(n9158), .ZN(n13082) );
  NAND2_X1 U11512 ( .A1(n13081), .A2(n13082), .ZN(n13080) );
  NAND2_X1 U11513 ( .A1(n13084), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9159) );
  NAND2_X1 U11514 ( .A1(n13080), .A2(n9159), .ZN(n13095) );
  XNOR2_X1 U11515 ( .A(n9160), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n13096) );
  NAND2_X1 U11516 ( .A1(n13095), .A2(n13096), .ZN(n13094) );
  INV_X1 U11517 ( .A(n9160), .ZN(n13097) );
  NAND2_X1 U11518 ( .A1(n13097), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9161) );
  NAND2_X1 U11519 ( .A1(n13094), .A2(n9161), .ZN(n13109) );
  INV_X1 U11520 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n14740) );
  MUX2_X1 U11521 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n14740), .S(n13112), .Z(
        n13110) );
  NAND2_X1 U11522 ( .A1(n13109), .A2(n13110), .ZN(n13108) );
  NAND2_X1 U11523 ( .A1(n13112), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9162) );
  NAND2_X1 U11524 ( .A1(n13108), .A2(n9162), .ZN(n14572) );
  INV_X1 U11525 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10012) );
  MUX2_X1 U11526 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10012), .S(n14577), .Z(
        n14573) );
  NAND2_X1 U11527 ( .A1(n14572), .A2(n14573), .ZN(n14571) );
  NAND2_X1 U11528 ( .A1(n14577), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9163) );
  NAND2_X1 U11529 ( .A1(n14571), .A2(n9163), .ZN(n9166) );
  INV_X1 U11530 ( .A(n9164), .ZN(n9165) );
  NAND2_X1 U11531 ( .A1(n9166), .A2(n9167), .ZN(n9182) );
  OAI211_X1 U11532 ( .C1(n9167), .C2(n9166), .A(n14586), .B(n9182), .ZN(n9168)
         );
  OAI211_X1 U11533 ( .C1(n9186), .C2(n9170), .A(n9169), .B(n9168), .ZN(
        P2_U3222) );
  INV_X1 U11534 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9180) );
  INV_X1 U11535 ( .A(n9171), .ZN(n9172) );
  NAND2_X1 U11536 ( .A1(n9173), .A2(n9172), .ZN(n9211) );
  INV_X1 U11537 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9284) );
  NAND3_X1 U11538 ( .A1(n14445), .A2(P1_IR_REG_0__SCAN_IN), .A3(n9284), .ZN(
        n9179) );
  INV_X1 U11539 ( .A(n9211), .ZN(n9203) );
  INV_X1 U11540 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9174) );
  AOI21_X1 U11541 ( .B1(n9424), .B2(n9174), .A(n8741), .ZN(n9425) );
  INV_X1 U11542 ( .A(n9425), .ZN(n9175) );
  AOI21_X1 U11543 ( .B1(n9284), .B2(n14132), .A(n9175), .ZN(n9176) );
  MUX2_X1 U11544 ( .A(n9176), .B(n9175), .S(P1_IR_REG_0__SCAN_IN), .Z(n9177)
         );
  AOI22_X1 U11545 ( .A1(n9203), .A2(n9177), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n9178) );
  OAI211_X1 U11546 ( .C1(n14456), .C2(n9180), .A(n9179), .B(n9178), .ZN(
        P1_U3243) );
  INV_X1 U11547 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10270) );
  MUX2_X1 U11548 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n10270), .S(n10066), .Z(
        n9185) );
  NAND2_X1 U11549 ( .A1(n9953), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9181) );
  NAND2_X1 U11550 ( .A1(n9182), .A2(n9181), .ZN(n9184) );
  OR2_X1 U11551 ( .A1(n9184), .A2(n9185), .ZN(n9445) );
  INV_X1 U11552 ( .A(n9445), .ZN(n9183) );
  AOI21_X1 U11553 ( .B1(n9185), .B2(n9184), .A(n9183), .ZN(n9194) );
  AOI21_X1 U11554 ( .B1(n9953), .B2(P2_REG2_REG_8__SCAN_IN), .A(n9186), .ZN(
        n9189) );
  INV_X1 U11555 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n9187) );
  MUX2_X1 U11556 ( .A(n9187), .B(P2_REG2_REG_9__SCAN_IN), .S(n10066), .Z(n9188) );
  NAND2_X1 U11557 ( .A1(n9189), .A2(n9188), .ZN(n9452) );
  OAI21_X1 U11558 ( .B1(n9189), .B2(n9188), .A(n9452), .ZN(n9192) );
  INV_X1 U11559 ( .A(n14602), .ZN(n14610) );
  NAND2_X1 U11560 ( .A1(n14610), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n9190) );
  NAND2_X1 U11561 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n10094) );
  OAI211_X1 U11562 ( .C1(n14618), .C2(n10066), .A(n9190), .B(n10094), .ZN(
        n9191) );
  AOI21_X1 U11563 ( .B1(n9192), .B2(n14579), .A(n9191), .ZN(n9193) );
  OAI21_X1 U11564 ( .B1(n9194), .B2(n14604), .A(n9193), .ZN(P2_U3223) );
  OAI222_X1 U11565 ( .A1(n12883), .A2(n9196), .B1(n12886), .B2(n9195), .C1(
        n12423), .C2(P3_U3151), .ZN(P3_U3282) );
  INV_X1 U11566 ( .A(n10643), .ZN(n9236) );
  NAND2_X1 U11567 ( .A1(n9200), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9198) );
  MUX2_X1 U11568 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9198), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n9199) );
  INV_X1 U11569 ( .A(n9199), .ZN(n9201) );
  NOR2_X1 U11570 ( .A1(n9201), .A2(n9618), .ZN(n10644) );
  INV_X1 U11571 ( .A(n10644), .ZN(n9711) );
  OAI222_X1 U11572 ( .A1(n13526), .A2(n9236), .B1(n9711), .B2(P2_U3088), .C1(
        n9202), .C2(n13523), .ZN(P2_U3315) );
  AND2_X1 U11573 ( .A1(n9203), .A2(n8741), .ZN(n14448) );
  INV_X1 U11574 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9204) );
  MUX2_X1 U11575 ( .A(n9204), .B(P1_REG1_REG_6__SCAN_IN), .S(n9467), .Z(n9210)
         );
  INV_X1 U11576 ( .A(n9219), .ZN(n9433) );
  XNOR2_X1 U11577 ( .A(n9212), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n13686) );
  AND2_X1 U11578 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n13685) );
  NAND2_X1 U11579 ( .A1(n13686), .A2(n13685), .ZN(n13684) );
  INV_X1 U11580 ( .A(n9212), .ZN(n13683) );
  NAND2_X1 U11581 ( .A1(n13683), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9205) );
  NAND2_X1 U11582 ( .A1(n13684), .A2(n9205), .ZN(n13702) );
  INV_X1 U11583 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n14533) );
  NAND2_X1 U11584 ( .A1(n13702), .A2(n13703), .ZN(n13701) );
  INV_X1 U11585 ( .A(n13696), .ZN(n13695) );
  NAND2_X1 U11586 ( .A1(n13695), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9206) );
  NAND2_X1 U11587 ( .A1(n13701), .A2(n9206), .ZN(n13709) );
  XNOR2_X1 U11588 ( .A(n13712), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n13710) );
  NAND2_X1 U11589 ( .A1(n13709), .A2(n13710), .ZN(n13708) );
  INV_X1 U11590 ( .A(n13712), .ZN(n13711) );
  NAND2_X1 U11591 ( .A1(n13711), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9207) );
  NAND2_X1 U11592 ( .A1(n13708), .A2(n9207), .ZN(n9436) );
  XNOR2_X1 U11593 ( .A(n9219), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n9437) );
  AND2_X1 U11594 ( .A1(n9436), .A2(n9437), .ZN(n9434) );
  AOI21_X1 U11595 ( .B1(n9433), .B2(P1_REG1_REG_4__SCAN_IN), .A(n9434), .ZN(
        n9241) );
  INV_X1 U11596 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9208) );
  MUX2_X1 U11597 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n9208), .S(n9222), .Z(n9240)
         );
  NAND2_X1 U11598 ( .A1(n9241), .A2(n9240), .ZN(n9239) );
  OAI21_X1 U11599 ( .B1(n9222), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9239), .ZN(
        n9209) );
  NOR2_X1 U11600 ( .A1(n9209), .A2(n9210), .ZN(n9466) );
  AOI211_X1 U11601 ( .C1(n9210), .C2(n9209), .A(n9466), .B(n13764), .ZN(n9227)
         );
  OR3_X1 U11602 ( .A1(n9211), .A2(n14132), .A3(n8741), .ZN(n14451) );
  MUX2_X1 U11603 ( .A(n11684), .B(P1_REG2_REG_1__SCAN_IN), .S(n9212), .Z(
        n13687) );
  AND2_X1 U11604 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n13688) );
  NAND2_X1 U11605 ( .A1(n13687), .A2(n13688), .ZN(n13699) );
  NAND2_X1 U11606 ( .A1(n13683), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n13698) );
  NAND2_X1 U11607 ( .A1(n13699), .A2(n13698), .ZN(n9215) );
  INV_X1 U11608 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9213) );
  MUX2_X1 U11609 ( .A(n9213), .B(P1_REG2_REG_2__SCAN_IN), .S(n13696), .Z(n9214) );
  NAND2_X1 U11610 ( .A1(n9215), .A2(n9214), .ZN(n13715) );
  NAND2_X1 U11611 ( .A1(n13695), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n13714) );
  NAND2_X1 U11612 ( .A1(n13715), .A2(n13714), .ZN(n9217) );
  INV_X1 U11613 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n14484) );
  MUX2_X1 U11614 ( .A(n14484), .B(P1_REG2_REG_3__SCAN_IN), .S(n13712), .Z(
        n9216) );
  NAND2_X1 U11615 ( .A1(n9217), .A2(n9216), .ZN(n13717) );
  NAND2_X1 U11616 ( .A1(n13711), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n9218) );
  NAND2_X1 U11617 ( .A1(n13717), .A2(n9218), .ZN(n9430) );
  INV_X1 U11618 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n9220) );
  MUX2_X1 U11619 ( .A(n9220), .B(P1_REG2_REG_4__SCAN_IN), .S(n9219), .Z(n9429)
         );
  AOI22_X1 U11620 ( .A1(n9430), .A2(n9429), .B1(P1_REG2_REG_4__SCAN_IN), .B2(
        n9433), .ZN(n9245) );
  INV_X1 U11621 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9221) );
  MUX2_X1 U11622 ( .A(n9221), .B(P1_REG2_REG_5__SCAN_IN), .S(n9222), .Z(n9244)
         );
  OR2_X1 U11623 ( .A1(n9245), .A2(n9244), .ZN(n9242) );
  NAND2_X1 U11624 ( .A1(n9222), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9224) );
  INV_X1 U11625 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9473) );
  MUX2_X1 U11626 ( .A(n9473), .B(P1_REG2_REG_6__SCAN_IN), .S(n9467), .Z(n9223)
         );
  AOI21_X1 U11627 ( .B1(n9242), .B2(n9224), .A(n9223), .ZN(n9511) );
  AND3_X1 U11628 ( .A1(n9242), .A2(n9224), .A3(n9223), .ZN(n9225) );
  NOR3_X1 U11629 ( .A1(n14451), .A2(n9511), .A3(n9225), .ZN(n9226) );
  NOR2_X1 U11630 ( .A1(n9227), .A2(n9226), .ZN(n9230) );
  INV_X1 U11631 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n13626) );
  NOR2_X1 U11632 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n13626), .ZN(n9228) );
  AOI21_X1 U11633 ( .B1(n13725), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n9228), .ZN(
        n9229) );
  OAI211_X1 U11634 ( .C1(n9474), .C2(n13722), .A(n9230), .B(n9229), .ZN(
        P1_U3249) );
  INV_X1 U11635 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n14732) );
  INV_X1 U11636 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n14548) );
  OAI22_X1 U11637 ( .A1(n14604), .A2(n14732), .B1(n14548), .B2(n14614), .ZN(
        n9233) );
  NAND2_X1 U11638 ( .A1(n14586), .A2(n14732), .ZN(n9231) );
  OAI211_X1 U11639 ( .C1(P2_REG2_REG_0__SCAN_IN), .C2(n14614), .A(n9231), .B(
        n14618), .ZN(n9232) );
  MUX2_X1 U11640 ( .A(n9233), .B(n9232), .S(P2_IR_REG_0__SCAN_IN), .Z(n9235)
         );
  INV_X1 U11641 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15170) );
  INV_X1 U11642 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n9367) );
  OAI22_X1 U11643 ( .A1(n14602), .A2(n15170), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9367), .ZN(n9234) );
  OR2_X1 U11644 ( .A1(n9235), .A2(n9234), .ZN(P2_U3214) );
  INV_X1 U11645 ( .A(n9936), .ZN(n9941) );
  OAI222_X1 U11646 ( .A1(n14135), .A2(n9237), .B1(n12134), .B2(n9236), .C1(
        n9941), .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U11647 ( .A(n10718), .ZN(n9254) );
  AOI22_X1 U11648 ( .A1(n10055), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n14127), .ZN(n9238) );
  OAI21_X1 U11649 ( .B1(n9254), .B2(n12134), .A(n9238), .ZN(P1_U3342) );
  OAI21_X1 U11650 ( .B1(n9241), .B2(n9240), .A(n9239), .ZN(n9247) );
  INV_X1 U11651 ( .A(n9242), .ZN(n9243) );
  AOI211_X1 U11652 ( .C1(n9245), .C2(n9244), .A(n9243), .B(n14451), .ZN(n9246)
         );
  AOI21_X1 U11653 ( .B1(n14445), .B2(n9247), .A(n9246), .ZN(n9250) );
  NAND2_X1 U11654 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10252) );
  INV_X1 U11655 ( .A(n10252), .ZN(n9248) );
  AOI21_X1 U11656 ( .B1(n13725), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n9248), .ZN(
        n9249) );
  OAI211_X1 U11657 ( .C1(n9251), .C2(n13722), .A(n9250), .B(n9249), .ZN(
        P1_U3248) );
  OR2_X1 U11658 ( .A1(n9618), .A2(n9884), .ZN(n9252) );
  XNOR2_X1 U11659 ( .A(n9252), .B(P2_IR_REG_13__SCAN_IN), .ZN(n10719) );
  INV_X1 U11660 ( .A(n10719), .ZN(n9708) );
  OAI222_X1 U11661 ( .A1(n13526), .A2(n9254), .B1(n9708), .B2(P2_U3088), .C1(
        n9253), .C2(n13523), .ZN(P2_U3314) );
  OR2_X1 U11662 ( .A1(n9268), .A2(P1_D_REG_1__SCAN_IN), .ZN(n9256) );
  NOR4_X1 U11663 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n9265) );
  NOR4_X1 U11664 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n9264) );
  OR4_X1 U11665 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n9262) );
  NOR4_X1 U11666 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n9260) );
  NOR4_X1 U11667 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n9259) );
  NOR4_X1 U11668 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9258) );
  NOR4_X1 U11669 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n9257) );
  NAND4_X1 U11670 ( .A1(n9260), .A2(n9259), .A3(n9258), .A4(n9257), .ZN(n9261)
         );
  NOR4_X1 U11671 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n9262), .A4(n9261), .ZN(n9263) );
  AND3_X1 U11672 ( .A1(n9265), .A2(n9264), .A3(n9263), .ZN(n10303) );
  OR2_X1 U11673 ( .A1(n9268), .A2(n10303), .ZN(n9813) );
  NOR2_X1 U11674 ( .A1(n9273), .A2(n9272), .ZN(n9266) );
  NAND2_X1 U11675 ( .A1(n9813), .A2(n9827), .ZN(n9267) );
  OR2_X1 U11676 ( .A1(n9268), .A2(P1_D_REG_0__SCAN_IN), .ZN(n9270) );
  AND2_X1 U11677 ( .A1(n10849), .A2(n9824), .ZN(n9693) );
  INV_X1 U11678 ( .A(n9693), .ZN(n9282) );
  NAND2_X1 U11679 ( .A1(n14137), .A2(n13878), .ZN(n9275) );
  NAND2_X1 U11680 ( .A1(n9273), .A2(n9272), .ZN(n9274) );
  NAND2_X1 U11681 ( .A1(n14137), .A2(n10062), .ZN(n9276) );
  INV_X2 U11682 ( .A(n12177), .ZN(n10099) );
  OR2_X1 U11683 ( .A1(n9824), .A2(n9416), .ZN(n10434) );
  AND2_X1 U11684 ( .A1(n10434), .A2(n10062), .ZN(n9277) );
  NAND2_X1 U11685 ( .A1(n10099), .A2(n9277), .ZN(n13855) );
  NAND3_X1 U11686 ( .A1(n9824), .A2(n13878), .A3(n10586), .ZN(n10480) );
  INV_X1 U11687 ( .A(n10444), .ZN(n9278) );
  OAI21_X1 U11688 ( .B1(n14529), .B2(n14518), .A(n9278), .ZN(n9281) );
  NAND2_X1 U11689 ( .A1(n9279), .A2(n13955), .ZN(n10438) );
  OAI211_X1 U11690 ( .C1(n9282), .C2(n10439), .A(n9281), .B(n10438), .ZN(
        n10157) );
  NAND2_X1 U11691 ( .A1(n10157), .A2(n14540), .ZN(n9283) );
  OAI21_X1 U11692 ( .B1(n14540), .B2(n9284), .A(n9283), .ZN(P1_U3528) );
  NAND3_X1 U11693 ( .A1(n9298), .A2(n9291), .A3(n14979), .ZN(n9286) );
  NAND2_X1 U11694 ( .A1(n9301), .A2(n9293), .ZN(n9285) );
  NAND2_X1 U11695 ( .A1(n9286), .A2(n9285), .ZN(n9287) );
  INV_X1 U11696 ( .A(n9300), .ZN(n9288) );
  NAND2_X1 U11697 ( .A1(n9288), .A2(n9301), .ZN(n9758) );
  INV_X1 U11698 ( .A(n9757), .ZN(n9289) );
  INV_X1 U11699 ( .A(n12341), .ZN(n12357) );
  OR2_X1 U11700 ( .A1(n9298), .A2(n14929), .ZN(n9290) );
  AOI22_X1 U11701 ( .A1(n12384), .A2(n12357), .B1(n12364), .B2(n9891), .ZN(
        n9305) );
  INV_X1 U11702 ( .A(n9291), .ZN(n9297) );
  AND3_X1 U11703 ( .A1(n10034), .A2(n9292), .A3(n9527), .ZN(n9296) );
  INV_X1 U11704 ( .A(n9293), .ZN(n9294) );
  OR2_X1 U11705 ( .A1(n9301), .A2(n9294), .ZN(n9295) );
  OAI211_X1 U11706 ( .C1(n9298), .C2(n9297), .A(n9296), .B(n9295), .ZN(n9299)
         );
  NAND2_X1 U11707 ( .A1(n9299), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9303) );
  OR2_X1 U11708 ( .A1(n9301), .A2(n9300), .ZN(n9302) );
  NAND2_X2 U11709 ( .A1(n9303), .A2(n9302), .ZN(n12358) );
  OR2_X1 U11710 ( .A1(n12358), .A2(P3_U3151), .ZN(n9889) );
  NAND2_X1 U11711 ( .A1(n9889), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n9304) );
  OAI211_X1 U11712 ( .C1(n9519), .C2(n12366), .A(n9305), .B(n9304), .ZN(
        P3_U3172) );
  XNOR2_X1 U11713 ( .A(n11269), .B(P2_B_REG_SCAN_IN), .ZN(n9306) );
  NAND2_X1 U11714 ( .A1(n11375), .A2(n9306), .ZN(n9307) );
  INV_X1 U11715 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9308) );
  NAND2_X1 U11716 ( .A1(n14654), .A2(n9308), .ZN(n9311) );
  INV_X1 U11717 ( .A(n9309), .ZN(n11489) );
  NAND2_X1 U11718 ( .A1(n11489), .A2(n11375), .ZN(n9310) );
  NAND2_X1 U11719 ( .A1(n9311), .A2(n9310), .ZN(n14660) );
  INV_X1 U11720 ( .A(n14660), .ZN(n9322) );
  NOR4_X1 U11721 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n9315) );
  NOR4_X1 U11722 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n9314) );
  NOR4_X1 U11723 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n9313) );
  NOR4_X1 U11724 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n9312) );
  NAND4_X1 U11725 ( .A1(n9315), .A2(n9314), .A3(n9313), .A4(n9312), .ZN(n9321)
         );
  NOR2_X1 U11726 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .ZN(
        n9319) );
  NOR4_X1 U11727 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n9318) );
  NOR4_X1 U11728 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n9317) );
  NOR4_X1 U11729 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n9316) );
  NAND4_X1 U11730 ( .A1(n9319), .A2(n9318), .A3(n9317), .A4(n9316), .ZN(n9320)
         );
  OAI21_X1 U11731 ( .B1(n9321), .B2(n9320), .A(n14654), .ZN(n9574) );
  NAND2_X1 U11732 ( .A1(n9322), .A2(n9574), .ZN(n9339) );
  INV_X1 U11733 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14657) );
  NAND2_X1 U11734 ( .A1(n14654), .A2(n14657), .ZN(n9324) );
  NAND2_X1 U11735 ( .A1(n11489), .A2(n11269), .ZN(n9323) );
  NAND2_X1 U11736 ( .A1(n9324), .A2(n9323), .ZN(n14658) );
  NAND2_X1 U11737 ( .A1(n9327), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9329) );
  XNOR2_X2 U11738 ( .A(n9329), .B(n8970), .ZN(n12062) );
  NAND2_X1 U11739 ( .A1(n14671), .A2(n9330), .ZN(n9573) );
  OAI21_X1 U11740 ( .B1(n9339), .B2(n14658), .A(n9573), .ZN(n9334) );
  NAND2_X1 U11741 ( .A1(n13154), .A2(n12062), .ZN(n12071) );
  NAND2_X1 U11742 ( .A1(n9373), .A2(n12071), .ZN(n10014) );
  AND2_X1 U11743 ( .A1(n9337), .A2(n10014), .ZN(n9333) );
  NAND2_X1 U11744 ( .A1(n9334), .A2(n9333), .ZN(n9675) );
  NOR2_X1 U11745 ( .A1(n9675), .A2(P2_U3088), .ZN(n9415) );
  NAND2_X1 U11746 ( .A1(n9335), .A2(SI_0_), .ZN(n9336) );
  XNOR2_X1 U11747 ( .A(n9336), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n13527) );
  MUX2_X1 U11748 ( .A(P2_IR_REG_0__SCAN_IN), .B(n13527), .S(n10065), .Z(n11802) );
  INV_X1 U11749 ( .A(n14658), .ZN(n9338) );
  INV_X1 U11750 ( .A(n9339), .ZN(n10171) );
  INV_X1 U11751 ( .A(n12062), .ZN(n12024) );
  NAND2_X1 U11752 ( .A1(n10173), .A2(n12024), .ZN(n14645) );
  INV_X1 U11753 ( .A(n9573), .ZN(n9340) );
  OAI21_X2 U11754 ( .B1(n9341), .B2(n14645), .A(n14646), .ZN(n13026) );
  NOR2_X1 U11755 ( .A1(n11802), .A2(n13300), .ZN(n9356) );
  NAND2_X1 U11756 ( .A1(n9345), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9346) );
  NAND2_X1 U11757 ( .A1(n7325), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n9354) );
  NAND2_X1 U11758 ( .A1(n9628), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n9353) );
  NAND2_X1 U11759 ( .A1(n9624), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9352) );
  NAND2_X1 U11760 ( .A1(n9387), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n9351) );
  INV_X1 U11761 ( .A(n11799), .ZN(n13066) );
  NAND2_X1 U11762 ( .A1(n11799), .A2(n11802), .ZN(n9563) );
  NAND2_X1 U11763 ( .A1(n11802), .A2(n13300), .ZN(n9355) );
  NAND2_X1 U11764 ( .A1(n9563), .A2(n9355), .ZN(n9379) );
  AOI21_X1 U11765 ( .B1(n9356), .B2(n13066), .A(n9379), .ZN(n9364) );
  INV_X1 U11766 ( .A(n9373), .ZN(n9357) );
  INV_X1 U11767 ( .A(n12071), .ZN(n12019) );
  NAND2_X1 U11768 ( .A1(n9387), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9363) );
  NAND2_X1 U11769 ( .A1(n9624), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9360) );
  INV_X1 U11770 ( .A(n12987), .ZN(n13036) );
  INV_X1 U11771 ( .A(n13036), .ZN(n13164) );
  NAND2_X1 U11772 ( .A1(n13064), .A2(n13164), .ZN(n10178) );
  OAI22_X1 U11773 ( .A1(n9364), .A2(n13018), .B1(n13015), .B2(n10178), .ZN(
        n9365) );
  AOI21_X1 U11774 ( .B1(n11802), .B2(n13026), .A(n9365), .ZN(n9366) );
  OAI21_X1 U11775 ( .B1(n9415), .B2(n9367), .A(n9366), .ZN(P2_U3204) );
  INV_X1 U11776 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10334) );
  NAND2_X1 U11777 ( .A1(n9387), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9371) );
  NAND2_X1 U11778 ( .A1(n7325), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n9370) );
  NAND2_X1 U11779 ( .A1(n9628), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n9369) );
  NAND2_X1 U11780 ( .A1(n9624), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n9368) );
  NAND4_X2 U11781 ( .A1(n9371), .A2(n9370), .A3(n9369), .A4(n9368), .ZN(n13063) );
  INV_X1 U11782 ( .A(n9144), .ZN(n9372) );
  AND2_X2 U11783 ( .A1(n9373), .A2(n9372), .ZN(n13004) );
  OAI22_X1 U11784 ( .A1(n7112), .A2(n13036), .B1(n11799), .B2(n13228), .ZN(
        n10330) );
  AOI22_X1 U11785 ( .A1(n13040), .A2(n10330), .B1(n13026), .B2(n11806), .ZN(
        n9385) );
  NAND2_X1 U11786 ( .A1(n13064), .A2(n9633), .ZN(n9407) );
  XNOR2_X1 U11787 ( .A(n9407), .B(n9405), .ZN(n9382) );
  INV_X1 U11788 ( .A(n11802), .ZN(n11798) );
  NAND2_X1 U11789 ( .A1(n9382), .A2(n9381), .ZN(n9409) );
  OAI21_X1 U11790 ( .B1(n9382), .B2(n9381), .A(n9409), .ZN(n9383) );
  NAND2_X1 U11791 ( .A1(n13034), .A2(n9383), .ZN(n9384) );
  OAI211_X1 U11792 ( .C1(n9415), .C2(n10334), .A(n9385), .B(n9384), .ZN(
        P2_U3194) );
  INV_X1 U11793 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10506) );
  NAND2_X1 U11794 ( .A1(n13064), .A2(n13004), .ZN(n9393) );
  INV_X1 U11795 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9386) );
  NAND2_X1 U11796 ( .A1(n7325), .A2(n9386), .ZN(n9391) );
  NAND2_X1 U11797 ( .A1(n9624), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9390) );
  NAND2_X1 U11798 ( .A1(n9628), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n9389) );
  NAND2_X1 U11799 ( .A1(n9387), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9388) );
  NAND4_X1 U11800 ( .A1(n9391), .A2(n9390), .A3(n9389), .A4(n9388), .ZN(n13062) );
  NAND2_X1 U11801 ( .A1(n13062), .A2(n12987), .ZN(n9392) );
  NAND2_X1 U11802 ( .A1(n9393), .A2(n9392), .ZN(n9568) );
  OR2_X1 U11803 ( .A1(n11980), .A2(n9396), .ZN(n9397) );
  OAI211_X1 U11804 ( .C1(n10065), .C2(n14556), .A(n9398), .B(n9397), .ZN(n9399) );
  AOI22_X1 U11805 ( .A1(n13040), .A2(n9568), .B1(n13026), .B2(n11813), .ZN(
        n9414) );
  AND2_X1 U11806 ( .A1(n13063), .A2(n9633), .ZN(n9400) );
  XNOR2_X1 U11807 ( .A(n9399), .B(n9858), .ZN(n9401) );
  NAND2_X1 U11808 ( .A1(n9400), .A2(n9401), .ZN(n9404) );
  INV_X1 U11809 ( .A(n9400), .ZN(n9403) );
  INV_X1 U11810 ( .A(n9401), .ZN(n9402) );
  NAND2_X1 U11811 ( .A1(n9403), .A2(n9402), .ZN(n9639) );
  INV_X1 U11812 ( .A(n9405), .ZN(n9406) );
  NAND2_X1 U11813 ( .A1(n9407), .A2(n9406), .ZN(n9408) );
  NAND2_X1 U11814 ( .A1(n9409), .A2(n9408), .ZN(n9410) );
  OAI21_X1 U11815 ( .B1(n9411), .B2(n9410), .A(n9640), .ZN(n9412) );
  NAND2_X1 U11816 ( .A1(n13034), .A2(n9412), .ZN(n9413) );
  OAI211_X1 U11817 ( .C1(n9415), .C2(n10506), .A(n9414), .B(n9413), .ZN(
        P2_U3209) );
  INV_X1 U11818 ( .A(n9418), .ZN(n9421) );
  AOI22_X1 U11819 ( .A1(n12247), .A2(n9840), .B1(n9421), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n9419) );
  NAND2_X1 U11820 ( .A1(n9420), .A2(n9419), .ZN(n9806) );
  OR2_X1 U11821 ( .A1(n9695), .A2(n12174), .ZN(n9423) );
  AOI22_X1 U11822 ( .A1(n12255), .A2(n9840), .B1(n9421), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n9422) );
  NAND2_X1 U11823 ( .A1(n9423), .A2(n9422), .ZN(n9805) );
  XNOR2_X1 U11824 ( .A(n9806), .B(n9805), .ZN(n9844) );
  MUX2_X1 U11825 ( .A(n9844), .B(n13688), .S(n9424), .Z(n9428) );
  OAI21_X1 U11826 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(n9425), .A(P1_U4016), .ZN(
        n9426) );
  AOI21_X1 U11827 ( .B1(n9428), .B2(n9427), .A(n9426), .ZN(n13692) );
  XNOR2_X1 U11828 ( .A(n9430), .B(n9429), .ZN(n9440) );
  INV_X1 U11829 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9431) );
  NAND2_X1 U11830 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n10114) );
  OAI21_X1 U11831 ( .B1(n14456), .B2(n9431), .A(n10114), .ZN(n9432) );
  AOI21_X1 U11832 ( .B1(n9433), .B2(n14448), .A(n9432), .ZN(n9439) );
  INV_X1 U11833 ( .A(n9434), .ZN(n9435) );
  OAI211_X1 U11834 ( .C1(n9437), .C2(n9436), .A(n14445), .B(n9435), .ZN(n9438)
         );
  OAI211_X1 U11835 ( .C1(n14451), .C2(n9440), .A(n9439), .B(n9438), .ZN(n9441)
         );
  OR2_X1 U11836 ( .A1(n13692), .A2(n9441), .ZN(P1_U3247) );
  INV_X1 U11837 ( .A(n9442), .ZN(n9443) );
  OAI222_X1 U11838 ( .A1(P3_U3151), .A2(n12419), .B1(n12883), .B2(n6729), .C1(
        n12886), .C2(n9443), .ZN(P3_U3281) );
  INV_X1 U11839 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n14337) );
  MUX2_X1 U11840 ( .A(n14337), .B(P2_REG1_REG_12__SCAN_IN), .S(n10644), .Z(
        n9451) );
  NAND2_X1 U11841 ( .A1(n10066), .A2(n10270), .ZN(n9444) );
  AND2_X1 U11842 ( .A1(n9445), .A2(n9444), .ZN(n14589) );
  INV_X1 U11843 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n15068) );
  MUX2_X1 U11844 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n15068), .S(n14593), .Z(
        n14588) );
  NAND2_X1 U11845 ( .A1(n14589), .A2(n14588), .ZN(n14587) );
  NAND2_X1 U11846 ( .A1(n14593), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n9446) );
  NAND2_X1 U11847 ( .A1(n14587), .A2(n9446), .ZN(n13131) );
  INV_X1 U11848 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n9447) );
  XNOR2_X1 U11849 ( .A(n13132), .B(n9447), .ZN(n13130) );
  NAND2_X1 U11850 ( .A1(n13131), .A2(n13130), .ZN(n13129) );
  NAND2_X1 U11851 ( .A1(n13132), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n9448) );
  NAND2_X1 U11852 ( .A1(n13129), .A2(n9448), .ZN(n9450) );
  INV_X1 U11853 ( .A(n9713), .ZN(n9449) );
  AOI21_X1 U11854 ( .B1(n9451), .B2(n9450), .A(n9449), .ZN(n9464) );
  INV_X1 U11855 ( .A(n10066), .ZN(n9453) );
  OAI21_X1 U11856 ( .B1(n9453), .B2(P2_REG2_REG_9__SCAN_IN), .A(n9452), .ZN(
        n14596) );
  INV_X1 U11857 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n9454) );
  MUX2_X1 U11858 ( .A(n9454), .B(P2_REG2_REG_10__SCAN_IN), .S(n14593), .Z(
        n14597) );
  NOR2_X1 U11859 ( .A1(n14596), .A2(n14597), .ZN(n14595) );
  AOI21_X1 U11860 ( .B1(n14593), .B2(P2_REG2_REG_10__SCAN_IN), .A(n14595), 
        .ZN(n13125) );
  INV_X1 U11861 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n9455) );
  MUX2_X1 U11862 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n9455), .S(n13132), .Z(
        n13124) );
  NOR2_X1 U11863 ( .A1(n13132), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n9457) );
  INV_X1 U11864 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n9456) );
  MUX2_X1 U11865 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n9456), .S(n10644), .Z(
        n9458) );
  OAI21_X1 U11866 ( .B1(n13126), .B2(n9457), .A(n9458), .ZN(n9702) );
  INV_X1 U11867 ( .A(n9702), .ZN(n9460) );
  NOR3_X1 U11868 ( .A1(n13126), .A2(n9458), .A3(n9457), .ZN(n9459) );
  OAI21_X1 U11869 ( .B1(n9460), .B2(n9459), .A(n14579), .ZN(n9463) );
  INV_X1 U11870 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10360) );
  NOR2_X1 U11871 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10360), .ZN(n10667) );
  NOR2_X1 U11872 ( .A1(n14618), .A2(n9711), .ZN(n9461) );
  AOI211_X1 U11873 ( .C1(n14610), .C2(P2_ADDR_REG_12__SCAN_IN), .A(n10667), 
        .B(n9461), .ZN(n9462) );
  OAI211_X1 U11874 ( .C1(n9464), .C2(n14604), .A(n9463), .B(n9462), .ZN(
        P2_U3226) );
  INV_X1 U11875 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9465) );
  MUX2_X1 U11876 ( .A(n9465), .B(P1_REG1_REG_10__SCAN_IN), .S(n9580), .Z(n9472) );
  INV_X1 U11877 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9468) );
  MUX2_X1 U11878 ( .A(n9468), .B(P1_REG1_REG_7__SCAN_IN), .S(n9506), .Z(n9502)
         );
  INV_X1 U11879 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9469) );
  MUX2_X1 U11880 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n9469), .S(n9477), .Z(n9493)
         );
  OAI21_X1 U11881 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n9477), .A(n9492), .ZN(
        n9599) );
  INV_X1 U11882 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9470) );
  MUX2_X1 U11883 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n9470), .S(n9602), .Z(n9600)
         );
  NAND2_X1 U11884 ( .A1(n9599), .A2(n9600), .ZN(n9598) );
  OAI21_X1 U11885 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9602), .A(n9598), .ZN(
        n9471) );
  NOR2_X1 U11886 ( .A1(n9471), .A2(n9472), .ZN(n9579) );
  AOI211_X1 U11887 ( .C1(n9472), .C2(n9471), .A(n13764), .B(n9579), .ZN(n9488)
         );
  NOR2_X1 U11888 ( .A1(n9474), .A2(n9473), .ZN(n9505) );
  INV_X1 U11889 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9475) );
  MUX2_X1 U11890 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n9475), .S(n9506), .Z(n9476)
         );
  OAI21_X1 U11891 ( .B1(n9511), .B2(n9505), .A(n9476), .ZN(n9509) );
  NAND2_X1 U11892 ( .A1(n9506), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9490) );
  INV_X1 U11893 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n9478) );
  MUX2_X1 U11894 ( .A(n9478), .B(P1_REG2_REG_8__SCAN_IN), .S(n9477), .Z(n9489)
         );
  AOI21_X1 U11895 ( .B1(n9509), .B2(n9490), .A(n9489), .ZN(n9607) );
  NOR2_X1 U11896 ( .A1(n9496), .A2(n9478), .ZN(n9601) );
  INV_X1 U11897 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9479) );
  MUX2_X1 U11898 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n9479), .S(n9602), .Z(n9480)
         );
  OAI21_X1 U11899 ( .B1(n9607), .B2(n9601), .A(n9480), .ZN(n9605) );
  NAND2_X1 U11900 ( .A1(n9602), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9482) );
  INV_X1 U11901 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n15141) );
  MUX2_X1 U11902 ( .A(n15141), .B(P1_REG2_REG_10__SCAN_IN), .S(n9580), .Z(
        n9481) );
  AOI21_X1 U11903 ( .B1(n9605), .B2(n9482), .A(n9481), .ZN(n9591) );
  INV_X1 U11904 ( .A(n9591), .ZN(n9484) );
  NAND3_X1 U11905 ( .A1(n9605), .A2(n9482), .A3(n9481), .ZN(n9483) );
  NAND3_X1 U11906 ( .A1(n9484), .A2(n13766), .A3(n9483), .ZN(n9486) );
  AND2_X1 U11907 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11320) );
  AOI21_X1 U11908 ( .B1(n13725), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n11320), 
        .ZN(n9485) );
  OAI211_X1 U11909 ( .C1(n13722), .C2(n9584), .A(n9486), .B(n9485), .ZN(n9487)
         );
  OR2_X1 U11910 ( .A1(n9488), .A2(n9487), .ZN(P1_U3253) );
  NAND3_X1 U11911 ( .A1(n9509), .A2(n9490), .A3(n9489), .ZN(n9491) );
  NAND2_X1 U11912 ( .A1(n13766), .A2(n9491), .ZN(n9500) );
  OAI21_X1 U11913 ( .B1(n9494), .B2(n9493), .A(n9492), .ZN(n9495) );
  NAND2_X1 U11914 ( .A1(n9495), .A2(n14445), .ZN(n9499) );
  AND2_X1 U11915 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n11025) );
  NOR2_X1 U11916 ( .A1(n13722), .A2(n9496), .ZN(n9497) );
  AOI211_X1 U11917 ( .C1(n13725), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n11025), .B(
        n9497), .ZN(n9498) );
  OAI211_X1 U11918 ( .C1(n9607), .C2(n9500), .A(n9499), .B(n9498), .ZN(
        P1_U3251) );
  AOI211_X1 U11919 ( .C1(n9503), .C2(n9502), .A(n13764), .B(n9501), .ZN(n9516)
         );
  AND2_X1 U11920 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9504) );
  AOI21_X1 U11921 ( .B1(n13725), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n9504), .ZN(
        n9513) );
  INV_X1 U11922 ( .A(n9505), .ZN(n9508) );
  MUX2_X1 U11923 ( .A(n9475), .B(P1_REG2_REG_7__SCAN_IN), .S(n9506), .Z(n9507)
         );
  NAND2_X1 U11924 ( .A1(n9508), .A2(n9507), .ZN(n9510) );
  OAI211_X1 U11925 ( .C1(n9511), .C2(n9510), .A(n13766), .B(n9509), .ZN(n9512)
         );
  OAI211_X1 U11926 ( .C1(n13722), .C2(n9514), .A(n9513), .B(n9512), .ZN(n9515)
         );
  OR2_X1 U11927 ( .A1(n9516), .A2(n9515), .ZN(P1_U3250) );
  OR2_X1 U11928 ( .A1(n9517), .A2(n14957), .ZN(n9518) );
  OR2_X1 U11929 ( .A1(n9519), .A2(n9518), .ZN(n9521) );
  OR2_X1 U11930 ( .A1(n14920), .A2(n14917), .ZN(n9520) );
  NAND2_X1 U11931 ( .A1(n9521), .A2(n9520), .ZN(n10036) );
  INV_X1 U11932 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n9522) );
  OAI22_X1 U11933 ( .A1(n10039), .A2(n12864), .B1(n14993), .B2(n9522), .ZN(
        n9523) );
  AOI21_X1 U11934 ( .B1(n10036), .B2(n14993), .A(n9523), .ZN(n9524) );
  INV_X1 U11935 ( .A(n9524), .ZN(P3_U3390) );
  INV_X1 U11936 ( .A(n10943), .ZN(n9525) );
  NAND2_X1 U11937 ( .A1(n9528), .A2(n9527), .ZN(n9529) );
  AND2_X1 U11938 ( .A1(n9530), .A2(n9529), .ZN(n9550) );
  AND2_X1 U11939 ( .A1(n9551), .A2(n9550), .ZN(n9545) );
  INV_X1 U11940 ( .A(n9545), .ZN(n9532) );
  AND2_X1 U11941 ( .A1(P3_U3897), .A2(n12880), .ZN(n14871) );
  INV_X1 U11942 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n9540) );
  MUX2_X1 U11943 ( .A(n7407), .B(n9540), .S(n6446), .Z(n9534) );
  INV_X1 U11944 ( .A(n6465), .ZN(n9533) );
  NAND2_X1 U11945 ( .A1(n9534), .A2(n9533), .ZN(n9786) );
  INV_X1 U11946 ( .A(n9534), .ZN(n9535) );
  NAND2_X1 U11947 ( .A1(n9535), .A2(n6465), .ZN(n9536) );
  AND2_X1 U11948 ( .A1(n9786), .A2(n9536), .ZN(n9537) );
  MUX2_X1 U11949 ( .A(P3_REG2_REG_0__SCAN_IN), .B(P3_REG1_REG_0__SCAN_IN), .S(
        n6446), .Z(n14749) );
  INV_X1 U11950 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n9538) );
  NOR2_X1 U11951 ( .A1(n14749), .A2(n9538), .ZN(n14751) );
  NAND2_X1 U11952 ( .A1(n9537), .A2(n14751), .ZN(n9787) );
  OAI21_X1 U11953 ( .B1(n9537), .B2(n14751), .A(n9787), .ZN(n9557) );
  AND2_X1 U11954 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n9538), .ZN(n9539) );
  INV_X1 U11955 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n9765) );
  OR3_X1 U11956 ( .A1(n9765), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n9768) );
  OAI21_X1 U11957 ( .B1(n6465), .B2(n9539), .A(n9768), .ZN(n9541) );
  OR2_X1 U11958 ( .A1(n9541), .A2(n9540), .ZN(n9769) );
  NAND2_X1 U11959 ( .A1(n9541), .A2(n9540), .ZN(n9542) );
  AND2_X1 U11960 ( .A1(n9769), .A2(n9542), .ZN(n9555) );
  NAND2_X1 U11961 ( .A1(n9545), .A2(n6446), .ZN(n14748) );
  INV_X1 U11962 ( .A(n9543), .ZN(n9544) );
  INV_X1 U11963 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n9546) );
  NOR2_X1 U11964 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n9546), .ZN(n14747) );
  OAI21_X1 U11965 ( .B1(n9559), .B2(n14747), .A(n6489), .ZN(n9547) );
  NAND2_X1 U11966 ( .A1(n9547), .A2(n7407), .ZN(n9548) );
  NAND2_X1 U11967 ( .A1(n9773), .A2(n9548), .ZN(n9549) );
  NAND2_X1 U11968 ( .A1(n14752), .A2(n9549), .ZN(n9554) );
  INV_X1 U11969 ( .A(n9550), .ZN(n9552) );
  AOI22_X1 U11970 ( .A1(n14879), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n9553) );
  OAI211_X1 U11971 ( .C1(n9555), .C2(n14748), .A(n9554), .B(n9553), .ZN(n9556)
         );
  AOI21_X1 U11972 ( .B1(n14871), .B2(n9557), .A(n9556), .ZN(n9558) );
  OAI21_X1 U11973 ( .B1(n6465), .B2(n14876), .A(n9558), .ZN(P3_U3183) );
  INV_X1 U11974 ( .A(n13064), .ZN(n9561) );
  OR2_X1 U11975 ( .A1(n11799), .A2(n11798), .ZN(n10175) );
  INV_X1 U11976 ( .A(n10175), .ZN(n10326) );
  OAI22_X1 U11977 ( .A1(n12026), .A2(n10326), .B1(n11806), .B2(n13064), .ZN(
        n9984) );
  XNOR2_X1 U11978 ( .A(n9984), .B(n12025), .ZN(n10512) );
  INV_X1 U11979 ( .A(n10512), .ZN(n9572) );
  INV_X1 U11980 ( .A(n14671), .ZN(n14718) );
  NOR2_X1 U11981 ( .A1(n10512), .A2(n14718), .ZN(n9571) );
  INV_X1 U11982 ( .A(n9563), .ZN(n10329) );
  NAND2_X1 U11983 ( .A1(n10328), .A2(n9565), .ZN(n9564) );
  NAND2_X1 U11984 ( .A1(n9564), .A2(n12025), .ZN(n9993) );
  NAND2_X1 U11985 ( .A1(n9993), .A2(n9566), .ZN(n9569) );
  NAND2_X1 U11986 ( .A1(n12072), .A2(n10176), .ZN(n11721) );
  OR2_X1 U11987 ( .A1(n9330), .A2(n12062), .ZN(n9567) );
  AOI21_X1 U11988 ( .B1(n9569), .B2(n13391), .A(n9568), .ZN(n10505) );
  NAND2_X1 U11989 ( .A1(n10324), .A2(n11814), .ZN(n14635) );
  OAI211_X1 U11990 ( .C1(n10324), .C2(n11814), .A(n13300), .B(n14635), .ZN(
        n10507) );
  OAI211_X1 U11991 ( .C1(n11814), .C2(n14723), .A(n10505), .B(n10507), .ZN(
        n9570) );
  AOI211_X1 U11992 ( .C1(n14728), .C2(n9572), .A(n9571), .B(n9570), .ZN(n14674) );
  NAND3_X1 U11993 ( .A1(n14660), .A2(n9574), .A3(n9573), .ZN(n10013) );
  INV_X1 U11994 ( .A(n10014), .ZN(n9575) );
  NOR2_X1 U11995 ( .A1(n10013), .A2(n9575), .ZN(n9577) );
  NAND2_X1 U11996 ( .A1(n14744), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9578) );
  OAI21_X1 U11997 ( .B1(n14674), .B2(n14744), .A(n9578), .ZN(P2_U3501) );
  INV_X1 U11998 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9581) );
  MUX2_X1 U11999 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n9581), .S(n9741), .Z(n9582) );
  OAI21_X1 U12000 ( .B1(n9583), .B2(n9582), .A(n9740), .ZN(n9596) );
  NOR2_X1 U12001 ( .A1(n9584), .A2(n15141), .ZN(n9589) );
  INV_X1 U12002 ( .A(n9589), .ZN(n9586) );
  MUX2_X1 U12003 ( .A(n9587), .B(P1_REG2_REG_11__SCAN_IN), .S(n9741), .Z(n9585) );
  NAND2_X1 U12004 ( .A1(n9586), .A2(n9585), .ZN(n9590) );
  INV_X1 U12005 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9587) );
  MUX2_X1 U12006 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n9587), .S(n9741), .Z(n9588) );
  OAI21_X1 U12007 ( .B1(n9591), .B2(n9589), .A(n9588), .ZN(n9735) );
  OAI211_X1 U12008 ( .C1(n9591), .C2(n9590), .A(n9735), .B(n13766), .ZN(n9594)
         );
  NAND2_X1 U12009 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14391)
         );
  INV_X1 U12010 ( .A(n14391), .ZN(n9592) );
  AOI21_X1 U12011 ( .B1(n13725), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n9592), .ZN(
        n9593) );
  OAI211_X1 U12012 ( .C1(n9736), .C2(n13722), .A(n9594), .B(n9593), .ZN(n9595)
         );
  AOI21_X1 U12013 ( .B1(n9596), .B2(n14445), .A(n9595), .ZN(n9597) );
  INV_X1 U12014 ( .A(n9597), .ZN(P1_U3254) );
  OAI21_X1 U12015 ( .B1(n9600), .B2(n9599), .A(n9598), .ZN(n9613) );
  INV_X1 U12016 ( .A(n9601), .ZN(n9604) );
  MUX2_X1 U12017 ( .A(n9479), .B(P1_REG2_REG_9__SCAN_IN), .S(n9602), .Z(n9603)
         );
  NAND2_X1 U12018 ( .A1(n9604), .A2(n9603), .ZN(n9606) );
  OAI211_X1 U12019 ( .C1(n9607), .C2(n9606), .A(n9605), .B(n13766), .ZN(n9610)
         );
  NAND2_X1 U12020 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n11199) );
  INV_X1 U12021 ( .A(n11199), .ZN(n9608) );
  AOI21_X1 U12022 ( .B1(n13725), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n9608), .ZN(
        n9609) );
  OAI211_X1 U12023 ( .C1(n13722), .C2(n9611), .A(n9610), .B(n9609), .ZN(n9612)
         );
  AOI21_X1 U12024 ( .B1(n9613), .B2(n14445), .A(n9612), .ZN(n9614) );
  INV_X1 U12025 ( .A(n9614), .ZN(P1_U3252) );
  INV_X1 U12026 ( .A(n12469), .ZN(n12463) );
  OAI222_X1 U12027 ( .A1(P3_U3151), .A2(n12463), .B1(n12883), .B2(n9616), .C1(
        n12886), .C2(n9615), .ZN(P3_U3280) );
  INV_X1 U12028 ( .A(n11113), .ZN(n9726) );
  INV_X1 U12029 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n9617) );
  AND2_X1 U12030 ( .A1(n9618), .A2(n9617), .ZN(n9729) );
  OR2_X1 U12031 ( .A1(n9729), .A2(n9884), .ZN(n9619) );
  XNOR2_X1 U12032 ( .A(n9619), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11114) );
  AOI22_X1 U12033 ( .A1(n11114), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n13519), .ZN(n9620) );
  OAI21_X1 U12034 ( .B1(n9726), .B2(n13526), .A(n9620), .ZN(P2_U3313) );
  NAND2_X1 U12035 ( .A1(n9621), .A2(n9951), .ZN(n9623) );
  AOI22_X1 U12036 ( .A1(n12001), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n11898), 
        .B2(n13097), .ZN(n9622) );
  NAND2_X1 U12037 ( .A1(n9623), .A2(n9622), .ZN(n14690) );
  INV_X4 U12038 ( .A(n9858), .ZN(n12911) );
  XNOR2_X1 U12039 ( .A(n14690), .B(n12911), .ZN(n9634) );
  INV_X2 U12040 ( .A(n9664), .ZN(n11992) );
  NAND2_X1 U12041 ( .A1(n11992), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9632) );
  NAND2_X1 U12042 ( .A1(n9387), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9631) );
  NAND3_X1 U12043 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n9667) );
  INV_X1 U12044 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9626) );
  NAND2_X1 U12045 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n9625) );
  NAND2_X1 U12046 ( .A1(n9626), .A2(n9625), .ZN(n9627) );
  AND2_X1 U12047 ( .A1(n9667), .A2(n9627), .ZN(n10190) );
  NAND2_X1 U12048 ( .A1(n7325), .A2(n10190), .ZN(n9630) );
  NAND2_X1 U12049 ( .A1(n9628), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n9629) );
  NAND2_X1 U12050 ( .A1(n13060), .A2(n9633), .ZN(n9635) );
  NAND2_X1 U12051 ( .A1(n9634), .A2(n9635), .ZN(n9845) );
  INV_X1 U12052 ( .A(n9634), .ZN(n9637) );
  INV_X1 U12053 ( .A(n9635), .ZN(n9636) );
  NAND2_X1 U12054 ( .A1(n9637), .A2(n9636), .ZN(n9638) );
  AND2_X1 U12055 ( .A1(n9845), .A2(n9638), .ZN(n9663) );
  NAND2_X1 U12056 ( .A1(n11898), .A2(n13070), .ZN(n9642) );
  NAND2_X1 U12057 ( .A1(n12001), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n9641) );
  NAND2_X1 U12058 ( .A1(n13062), .A2(n9633), .ZN(n9644) );
  INV_X1 U12059 ( .A(n9644), .ZN(n9647) );
  INV_X1 U12060 ( .A(n9645), .ZN(n9646) );
  NAND2_X1 U12061 ( .A1(n9648), .A2(n9951), .ZN(n9650) );
  AOI22_X1 U12062 ( .A1(n12001), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n11898), 
        .B2(n13084), .ZN(n9649) );
  NAND2_X1 U12063 ( .A1(n9650), .A2(n9649), .ZN(n14683) );
  XNOR2_X1 U12064 ( .A(n14683), .B(n12911), .ZN(n9656) );
  NAND2_X1 U12065 ( .A1(n9387), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9655) );
  NAND2_X1 U12066 ( .A1(n9628), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n9654) );
  INV_X1 U12067 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n9651) );
  XNOR2_X1 U12068 ( .A(n9651), .B(P2_REG3_REG_3__SCAN_IN), .ZN(n10204) );
  NAND2_X1 U12069 ( .A1(n7325), .A2(n10204), .ZN(n9653) );
  NAND2_X1 U12070 ( .A1(n11992), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9652) );
  NAND4_X1 U12071 ( .A1(n9655), .A2(n9654), .A3(n9653), .A4(n9652), .ZN(n13061) );
  NAND2_X1 U12072 ( .A1(n13061), .A2(n9633), .ZN(n9657) );
  NAND2_X1 U12073 ( .A1(n9656), .A2(n9657), .ZN(n9661) );
  INV_X1 U12074 ( .A(n9656), .ZN(n9659) );
  INV_X1 U12075 ( .A(n9657), .ZN(n9658) );
  NAND2_X1 U12076 ( .A1(n9659), .A2(n9658), .ZN(n9660) );
  AND2_X1 U12077 ( .A1(n9661), .A2(n9660), .ZN(n9682) );
  NAND2_X1 U12078 ( .A1(n9683), .A2(n9682), .ZN(n9681) );
  OAI21_X1 U12079 ( .B1(n9663), .B2(n9662), .A(n9846), .ZN(n9679) );
  INV_X1 U12080 ( .A(n14690), .ZN(n10192) );
  NAND2_X1 U12081 ( .A1(n13061), .A2(n13004), .ZN(n9674) );
  NAND2_X1 U12082 ( .A1(n11992), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n9672) );
  NAND2_X1 U12083 ( .A1(n11971), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9671) );
  INV_X1 U12084 ( .A(n9667), .ZN(n9665) );
  NAND2_X1 U12085 ( .A1(n9665), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n9861) );
  INV_X1 U12086 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9666) );
  NAND2_X1 U12087 ( .A1(n9667), .A2(n9666), .ZN(n9668) );
  AND2_X1 U12088 ( .A1(n9861), .A2(n9668), .ZN(n13024) );
  NAND2_X1 U12089 ( .A1(n7325), .A2(n13024), .ZN(n9670) );
  NAND2_X1 U12090 ( .A1(n9628), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n9669) );
  NAND2_X1 U12091 ( .A1(n13059), .A2(n12987), .ZN(n9673) );
  NAND2_X1 U12092 ( .A1(n9674), .A2(n9673), .ZN(n10186) );
  AND2_X1 U12093 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n13103) );
  AOI21_X1 U12094 ( .B1(n13040), .B2(n10186), .A(n13103), .ZN(n9677) );
  NAND2_X1 U12095 ( .A1(n13025), .A2(n10190), .ZN(n9676) );
  OAI211_X1 U12096 ( .C1(n10192), .C2(n13043), .A(n9677), .B(n9676), .ZN(n9678) );
  AOI21_X1 U12097 ( .B1(n9679), .B2(n13034), .A(n9678), .ZN(n9680) );
  INV_X1 U12098 ( .A(n9680), .ZN(P2_U3199) );
  OAI21_X1 U12099 ( .B1(n9683), .B2(n9682), .A(n9681), .ZN(n9689) );
  INV_X1 U12100 ( .A(n14683), .ZN(n10206) );
  NAND2_X1 U12101 ( .A1(n13062), .A2(n13004), .ZN(n9685) );
  NAND2_X1 U12102 ( .A1(n13060), .A2(n12987), .ZN(n9684) );
  NAND2_X1 U12103 ( .A1(n9685), .A2(n9684), .ZN(n10200) );
  AND2_X1 U12104 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n13089) );
  AOI21_X1 U12105 ( .B1(n13040), .B2(n10200), .A(n13089), .ZN(n9687) );
  NAND2_X1 U12106 ( .A1(n13025), .A2(n10204), .ZN(n9686) );
  OAI211_X1 U12107 ( .C1(n10206), .C2(n13043), .A(n9687), .B(n9686), .ZN(n9688) );
  AOI21_X1 U12108 ( .B1(n9689), .B2(n13034), .A(n9688), .ZN(n9690) );
  INV_X1 U12109 ( .A(n9690), .ZN(P2_U3202) );
  NOR2_X1 U12110 ( .A1(n9695), .A2(n10439), .ZN(n10287) );
  XNOR2_X1 U12111 ( .A(n10288), .B(n10287), .ZN(n11688) );
  NAND2_X1 U12112 ( .A1(n10439), .A2(n11693), .ZN(n10464) );
  OR2_X1 U12113 ( .A1(n10439), .A2(n11693), .ZN(n9691) );
  NAND2_X1 U12114 ( .A1(n10464), .A2(n9691), .ZN(n11685) );
  NOR2_X1 U12115 ( .A1(n8691), .A2(n13983), .ZN(n11689) );
  AOI21_X1 U12116 ( .B1(n14522), .B2(n6634), .A(n11689), .ZN(n9694) );
  OAI21_X1 U12117 ( .B1(n13961), .B2(n11685), .A(n9694), .ZN(n9700) );
  INV_X1 U12118 ( .A(n10288), .ZN(n9696) );
  OAI21_X1 U12119 ( .B1(n9696), .B2(n9695), .A(n14529), .ZN(n9699) );
  INV_X1 U12120 ( .A(n13954), .ZN(n13982) );
  XNOR2_X1 U12121 ( .A(n11685), .B(n9279), .ZN(n9697) );
  AOI21_X1 U12122 ( .B1(n9697), .B2(n14529), .A(n13680), .ZN(n9698) );
  AOI21_X1 U12123 ( .B1(n9699), .B2(n13982), .A(n9698), .ZN(n11690) );
  AOI211_X1 U12124 ( .C1(n14518), .C2(n11688), .A(n9700), .B(n11690), .ZN(
        n14502) );
  NAND2_X1 U12125 ( .A1(n14537), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9701) );
  OAI21_X1 U12126 ( .B1(n14502), .B2(n14537), .A(n9701), .ZN(P1_U3529) );
  OAI21_X1 U12127 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n10644), .A(n9702), .ZN(
        n9705) );
  INV_X1 U12128 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n9703) );
  MUX2_X1 U12129 ( .A(n9703), .B(P2_REG2_REG_13__SCAN_IN), .S(n10719), .Z(
        n9704) );
  NOR2_X1 U12130 ( .A1(n9705), .A2(n9704), .ZN(n9911) );
  AOI211_X1 U12131 ( .C1(n9705), .C2(n9704), .A(n14614), .B(n9911), .ZN(n9710)
         );
  INV_X1 U12132 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n10732) );
  NOR2_X1 U12133 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10732), .ZN(n9706) );
  AOI21_X1 U12134 ( .B1(n14610), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n9706), .ZN(
        n9707) );
  OAI21_X1 U12135 ( .B1(n9708), .B2(n14618), .A(n9707), .ZN(n9709) );
  NOR2_X1 U12136 ( .A1(n9710), .A2(n9709), .ZN(n9718) );
  NAND2_X1 U12137 ( .A1(n9711), .A2(n14337), .ZN(n9712) );
  INV_X1 U12138 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9714) );
  XNOR2_X1 U12139 ( .A(n10719), .B(n9714), .ZN(n9715) );
  NAND2_X1 U12140 ( .A1(n9716), .A2(n9715), .ZN(n9916) );
  OAI211_X1 U12141 ( .C1(n9716), .C2(n9715), .A(n9916), .B(n14586), .ZN(n9717)
         );
  NAND2_X1 U12142 ( .A1(n9718), .A2(n9717), .ZN(P2_U3227) );
  XNOR2_X1 U12143 ( .A(n9720), .B(n9719), .ZN(n9724) );
  INV_X1 U12144 ( .A(n13061), .ZN(n9997) );
  OAI22_X1 U12145 ( .A1(n7112), .A2(n13228), .B1(n9997), .B2(n13036), .ZN(
        n14643) );
  AOI22_X1 U12146 ( .A1(n13040), .A2(n14643), .B1(P2_U3088), .B2(
        P2_REG3_REG_3__SCAN_IN), .ZN(n9721) );
  OAI21_X1 U12147 ( .B1(n14677), .B2(n13043), .A(n9721), .ZN(n9722) );
  AOI21_X1 U12148 ( .B1(n13025), .B2(n9386), .A(n9722), .ZN(n9723) );
  OAI21_X1 U12149 ( .B1(n9724), .B2(n13018), .A(n9723), .ZN(P2_U3190) );
  INV_X1 U12150 ( .A(n11347), .ZN(n9732) );
  INV_X1 U12151 ( .A(n13733), .ZN(n13729) );
  OAI222_X1 U12152 ( .A1(n14135), .A2(n9725), .B1(n12134), .B2(n9732), .C1(
        n13729), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U12153 ( .A(n10973), .ZN(n10964) );
  OAI222_X1 U12154 ( .A1(n14135), .A2(n9727), .B1(n12134), .B2(n9726), .C1(
        n10964), .C2(P1_U3086), .ZN(P1_U3341) );
  INV_X1 U12155 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n9728) );
  AND2_X1 U12156 ( .A1(n9729), .A2(n9728), .ZN(n9882) );
  INV_X1 U12157 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n9730) );
  NAND2_X1 U12158 ( .A1(n9882), .A2(n9730), .ZN(n9886) );
  NAND2_X1 U12159 ( .A1(n9886), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9731) );
  XNOR2_X1 U12160 ( .A(n9731), .B(P2_IR_REG_16__SCAN_IN), .ZN(n11348) );
  INV_X1 U12161 ( .A(n11348), .ZN(n11039) );
  OAI222_X1 U12162 ( .A1(n13523), .A2(n9733), .B1(n11039), .B2(P2_U3088), .C1(
        n13526), .C2(n9732), .ZN(P2_U3311) );
  INV_X1 U12163 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n9734) );
  MUX2_X1 U12164 ( .A(n9734), .B(P1_REG2_REG_12__SCAN_IN), .S(n9936), .Z(n9738) );
  OAI21_X1 U12165 ( .B1(n9736), .B2(n9587), .A(n9735), .ZN(n9737) );
  NOR2_X1 U12166 ( .A1(n9737), .A2(n9738), .ZN(n9940) );
  AOI21_X1 U12167 ( .B1(n9738), .B2(n9737), .A(n9940), .ZN(n9748) );
  INV_X1 U12168 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9739) );
  MUX2_X1 U12169 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9739), .S(n9936), .Z(n9743) );
  OAI21_X1 U12170 ( .B1(n9743), .B2(n9742), .A(n9935), .ZN(n9744) );
  NAND2_X1 U12171 ( .A1(n9744), .A2(n14445), .ZN(n9747) );
  AND2_X1 U12172 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n11534) );
  NOR2_X1 U12173 ( .A1(n13722), .A2(n9941), .ZN(n9745) );
  AOI211_X1 U12174 ( .C1(n13725), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n11534), 
        .B(n9745), .ZN(n9746) );
  OAI211_X1 U12175 ( .C1(n9748), .C2(n14451), .A(n9747), .B(n9746), .ZN(
        P1_U3255) );
  NAND2_X1 U12176 ( .A1(n8763), .A2(n9893), .ZN(n9749) );
  NAND2_X1 U12177 ( .A1(n9750), .A2(n9749), .ZN(n14940) );
  OR2_X1 U12178 ( .A1(n8763), .A2(n9751), .ZN(n9752) );
  NAND2_X1 U12179 ( .A1(n9753), .A2(n9752), .ZN(n12807) );
  NAND2_X1 U12180 ( .A1(n10140), .A2(n10225), .ZN(n9756) );
  MUX2_X1 U12181 ( .A(n14940), .B(n12807), .S(n11664), .Z(n9763) );
  NAND2_X1 U12182 ( .A1(n9889), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n9761) );
  AOI22_X1 U12183 ( .A1(n12338), .A2(n12805), .B1(n12364), .B2(n9759), .ZN(
        n9760) );
  OAI211_X1 U12184 ( .C1(n10141), .C2(n12341), .A(n9761), .B(n9760), .ZN(n9762) );
  AOI21_X1 U12185 ( .B1(n9763), .B2(n12346), .A(n9762), .ZN(n9764) );
  INV_X1 U12186 ( .A(n9764), .ZN(P3_U3162) );
  OAI22_X1 U12187 ( .A1(n12803), .A2(n10039), .B1(n15164), .B2(n9765), .ZN(
        n9766) );
  AOI21_X1 U12188 ( .B1(n10036), .B2(n15164), .A(n9766), .ZN(n9767) );
  INV_X1 U12189 ( .A(n9767), .ZN(P3_U3459) );
  INV_X1 U12190 ( .A(n6462), .ZN(n10867) );
  INV_X1 U12191 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n9781) );
  MUX2_X1 U12192 ( .A(P3_REG1_REG_2__SCAN_IN), .B(n9781), .S(n6462), .Z(n9771)
         );
  NAND2_X1 U12193 ( .A1(n9769), .A2(n9768), .ZN(n9770) );
  NAND2_X1 U12194 ( .A1(n9771), .A2(n9770), .ZN(n10866) );
  OAI21_X1 U12195 ( .B1(n9771), .B2(n9770), .A(n10866), .ZN(n9772) );
  INV_X1 U12196 ( .A(n9772), .ZN(n9780) );
  INV_X1 U12197 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n14933) );
  XNOR2_X1 U12198 ( .A(n10851), .B(n14933), .ZN(n9775) );
  NAND2_X1 U12199 ( .A1(n9773), .A2(n6489), .ZN(n9774) );
  NAND2_X1 U12200 ( .A1(n9775), .A2(n9774), .ZN(n10853) );
  OAI21_X1 U12201 ( .B1(n9775), .B2(n9774), .A(n10853), .ZN(n9776) );
  NAND2_X1 U12202 ( .A1(n14752), .A2(n9776), .ZN(n9779) );
  INV_X1 U12203 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n9904) );
  NOR2_X1 U12204 ( .A1(n9904), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9777) );
  AOI21_X1 U12205 ( .B1(n14879), .B2(P3_ADDR_REG_2__SCAN_IN), .A(n9777), .ZN(
        n9778) );
  OAI211_X1 U12206 ( .C1(n9780), .C2(n14748), .A(n9779), .B(n9778), .ZN(n9791)
         );
  MUX2_X1 U12207 ( .A(n14933), .B(n9781), .S(n6446), .Z(n9782) );
  NAND2_X1 U12208 ( .A1(n9782), .A2(n10867), .ZN(n10879) );
  INV_X1 U12209 ( .A(n9782), .ZN(n9783) );
  NAND2_X1 U12210 ( .A1(n9783), .A2(n6462), .ZN(n9784) );
  NAND2_X1 U12211 ( .A1(n10879), .A2(n9784), .ZN(n9785) );
  AOI21_X1 U12212 ( .B1(n9787), .B2(n9786), .A(n9785), .ZN(n14762) );
  INV_X1 U12213 ( .A(n14762), .ZN(n9789) );
  NAND3_X1 U12214 ( .A1(n9787), .A2(n9786), .A3(n9785), .ZN(n9788) );
  AOI21_X1 U12215 ( .B1(n9789), .B2(n9788), .A(n14895), .ZN(n9790) );
  AOI211_X1 U12216 ( .C1(n14906), .C2(n10867), .A(n9791), .B(n9790), .ZN(n9792) );
  INV_X1 U12217 ( .A(n9792), .ZN(P3_U3184) );
  INV_X1 U12218 ( .A(n11427), .ZN(n9832) );
  NAND2_X1 U12219 ( .A1(n10042), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9793) );
  XNOR2_X1 U12220 ( .A(n9793), .B(P2_IR_REG_17__SCAN_IN), .ZN(n13138) );
  INV_X1 U12221 ( .A(n13138), .ZN(n13145) );
  OAI222_X1 U12222 ( .A1(n13526), .A2(n9832), .B1(n13145), .B2(P2_U3088), .C1(
        n9794), .C2(n13523), .ZN(P2_U3310) );
  INV_X1 U12223 ( .A(n9795), .ZN(n9796) );
  INV_X1 U12224 ( .A(n12478), .ZN(n12485) );
  OAI222_X1 U12225 ( .A1(n12883), .A2(n9797), .B1(n12886), .B2(n9796), .C1(
        n12485), .C2(P3_U3151), .ZN(P3_U3279) );
  NAND2_X1 U12226 ( .A1(n9279), .A2(n12247), .ZN(n9799) );
  OR2_X1 U12227 ( .A1(n12263), .A2(n11693), .ZN(n9798) );
  NAND2_X1 U12228 ( .A1(n9799), .A2(n9798), .ZN(n9800) );
  XNOR2_X1 U12229 ( .A(n9800), .B(n10099), .ZN(n9802) );
  INV_X1 U12230 ( .A(n9802), .ZN(n9804) );
  INV_X1 U12231 ( .A(n9801), .ZN(n9803) );
  MUX2_X1 U12232 ( .A(n12177), .B(n9806), .S(n9805), .Z(n9835) );
  INV_X1 U12233 ( .A(n9807), .ZN(n9808) );
  NOR2_X1 U12234 ( .A1(n9834), .A2(n9808), .ZN(n9811) );
  OAI22_X1 U12235 ( .A1(n8691), .A2(n12264), .B1(n14504), .B2(n12263), .ZN(
        n9809) );
  XNOR2_X1 U12236 ( .A(n9809), .B(n10099), .ZN(n10104) );
  OAI22_X1 U12237 ( .A1(n8691), .A2(n9810), .B1(n14504), .B2(n12264), .ZN(
        n10103) );
  XNOR2_X1 U12238 ( .A(n10104), .B(n10103), .ZN(n9812) );
  AOI21_X1 U12239 ( .B1(n9811), .B2(n9812), .A(n10098), .ZN(n9831) );
  NAND3_X1 U12240 ( .A1(n10302), .A2(n10308), .A3(n9813), .ZN(n9820) );
  AND2_X1 U12241 ( .A1(n14511), .A2(n9814), .ZN(n9815) );
  NAND2_X1 U12242 ( .A1(n9826), .A2(n10307), .ZN(n13647) );
  INV_X1 U12243 ( .A(n13647), .ZN(n14358) );
  OR2_X1 U12244 ( .A1(n9817), .A2(n13983), .ZN(n9819) );
  NAND2_X1 U12245 ( .A1(n9279), .A2(n13954), .ZN(n9818) );
  NAND2_X1 U12246 ( .A1(n9819), .A2(n9818), .ZN(n10459) );
  NAND2_X1 U12247 ( .A1(n9820), .A2(n9827), .ZN(n9823) );
  AND3_X1 U12248 ( .A1(n9418), .A2(n10307), .A3(n9821), .ZN(n9822) );
  NAND2_X1 U12249 ( .A1(n9823), .A2(n9822), .ZN(n10111) );
  OR2_X1 U12250 ( .A1(n10111), .A2(P1_U3086), .ZN(n9841) );
  AOI22_X1 U12251 ( .A1(n14358), .A2(n10459), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n9841), .ZN(n9830) );
  AND2_X1 U12252 ( .A1(n9825), .A2(n9824), .ZN(n14263) );
  NAND2_X1 U12253 ( .A1(n9826), .A2(n14263), .ZN(n9828) );
  NAND2_X1 U12254 ( .A1(n14389), .A2(n10463), .ZN(n9829) );
  OAI211_X1 U12255 ( .C1(n9831), .C2(n14384), .A(n9830), .B(n9829), .ZN(
        P1_U3237) );
  INV_X1 U12256 ( .A(n13741), .ZN(n13748) );
  OAI222_X1 U12257 ( .A1(n14135), .A2(n9833), .B1(n12134), .B2(n9832), .C1(
        n13748), .C2(P1_U3086), .ZN(P1_U3338) );
  AOI21_X1 U12258 ( .B1(n9836), .B2(n9835), .A(n9834), .ZN(n9839) );
  INV_X1 U12259 ( .A(n14378), .ZN(n13629) );
  INV_X1 U12260 ( .A(n14377), .ZN(n13625) );
  AOI22_X1 U12261 ( .A1(n13629), .A2(n13680), .B1(n13625), .B2(n13678), .ZN(
        n9838) );
  AOI22_X1 U12262 ( .A1(n14389), .A2(n6634), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n9841), .ZN(n9837) );
  OAI211_X1 U12263 ( .C1(n9839), .C2(n14384), .A(n9838), .B(n9837), .ZN(
        P1_U3222) );
  AOI22_X1 U12264 ( .A1(n13625), .A2(n9279), .B1(n9840), .B2(n14389), .ZN(
        n9843) );
  NAND2_X1 U12265 ( .A1(n9841), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n9842) );
  OAI211_X1 U12266 ( .C1(n9844), .C2(n14384), .A(n9843), .B(n9842), .ZN(
        P1_U3232) );
  OR2_X1 U12267 ( .A1(n9847), .A2(n9394), .ZN(n9849) );
  AOI22_X1 U12268 ( .A1(n12001), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n11898), 
        .B2(n13112), .ZN(n9848) );
  XNOR2_X1 U12269 ( .A(n14702), .B(n12911), .ZN(n9850) );
  NAND2_X1 U12270 ( .A1(n13059), .A2(n9633), .ZN(n9851) );
  XNOR2_X1 U12271 ( .A(n9850), .B(n9851), .ZN(n13021) );
  INV_X1 U12272 ( .A(n9850), .ZN(n9853) );
  INV_X1 U12273 ( .A(n9851), .ZN(n9852) );
  NAND2_X1 U12274 ( .A1(n9853), .A2(n9852), .ZN(n9854) );
  OR2_X1 U12275 ( .A1(n9855), .A2(n9394), .ZN(n9857) );
  AOI22_X1 U12276 ( .A1(n12001), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n11898), 
        .B2(n14577), .ZN(n9856) );
  XNOR2_X1 U12277 ( .A(n14619), .B(n12960), .ZN(n9964) );
  NAND2_X1 U12278 ( .A1(n11992), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9866) );
  NAND2_X1 U12279 ( .A1(n11971), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9865) );
  INV_X1 U12280 ( .A(n9861), .ZN(n9859) );
  NAND2_X1 U12281 ( .A1(n9859), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n9869) );
  INV_X1 U12282 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9860) );
  NAND2_X1 U12283 ( .A1(n9861), .A2(n9860), .ZN(n9862) );
  AND2_X1 U12284 ( .A1(n9869), .A2(n9862), .ZN(n14622) );
  NAND2_X1 U12285 ( .A1(n7325), .A2(n14622), .ZN(n9864) );
  NAND2_X1 U12286 ( .A1(n9628), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n9863) );
  NAND4_X1 U12287 ( .A1(n9866), .A2(n9865), .A3(n9864), .A4(n9863), .ZN(n13058) );
  NAND2_X1 U12288 ( .A1(n13058), .A2(n9633), .ZN(n9962) );
  XNOR2_X1 U12289 ( .A(n9964), .B(n9962), .ZN(n9960) );
  XNOR2_X1 U12290 ( .A(n9960), .B(n9961), .ZN(n9881) );
  NAND2_X1 U12291 ( .A1(n13059), .A2(n13004), .ZN(n9876) );
  NAND2_X1 U12292 ( .A1(n11971), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9874) );
  NAND2_X1 U12293 ( .A1(n11992), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9873) );
  INV_X1 U12294 ( .A(n9869), .ZN(n9867) );
  NAND2_X1 U12295 ( .A1(n9867), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n9969) );
  INV_X1 U12296 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9868) );
  NAND2_X1 U12297 ( .A1(n9869), .A2(n9868), .ZN(n9870) );
  AND2_X1 U12298 ( .A1(n9969), .A2(n9870), .ZN(n10707) );
  NAND2_X1 U12299 ( .A1(n7325), .A2(n10707), .ZN(n9872) );
  NAND2_X1 U12300 ( .A1(n9628), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n9871) );
  NAND4_X1 U12301 ( .A1(n9874), .A2(n9873), .A3(n9872), .A4(n9871), .ZN(n13057) );
  NAND2_X1 U12302 ( .A1(n13057), .A2(n12987), .ZN(n9875) );
  NAND2_X1 U12303 ( .A1(n9876), .A2(n9875), .ZN(n10006) );
  INV_X1 U12304 ( .A(n10006), .ZN(n9877) );
  OAI22_X1 U12305 ( .A1(n13015), .A2(n9877), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9860), .ZN(n9878) );
  AOI21_X1 U12306 ( .B1(n14622), .B2(n13025), .A(n9878), .ZN(n9880) );
  NAND2_X1 U12307 ( .A1(n13026), .A2(n14619), .ZN(n9879) );
  OAI211_X1 U12308 ( .C1(n9881), .C2(n13018), .A(n9880), .B(n9879), .ZN(
        P2_U3185) );
  INV_X1 U12309 ( .A(n11286), .ZN(n9906) );
  NOR2_X1 U12310 ( .A1(n9882), .A2(n9884), .ZN(n9883) );
  MUX2_X1 U12311 ( .A(n9884), .B(n9883), .S(P2_IR_REG_15__SCAN_IN), .Z(n9885)
         );
  INV_X1 U12312 ( .A(n9885), .ZN(n9887) );
  AND2_X1 U12313 ( .A1(n9887), .A2(n9886), .ZN(n11287) );
  INV_X1 U12314 ( .A(n11287), .ZN(n10404) );
  OAI222_X1 U12315 ( .A1(n13526), .A2(n9906), .B1(n10404), .B2(P2_U3088), .C1(
        n9888), .C2(n13523), .ZN(P2_U3312) );
  INV_X1 U12316 ( .A(n9889), .ZN(n9905) );
  INV_X4 U12317 ( .A(n11664), .ZN(n11698) );
  NAND3_X1 U12318 ( .A1(n12805), .A2(n11664), .A3(n9891), .ZN(n9892) );
  OAI21_X1 U12319 ( .B1(n14920), .B2(n11698), .A(n9892), .ZN(n9897) );
  INV_X1 U12320 ( .A(n9893), .ZN(n9894) );
  AOI211_X1 U12321 ( .C1(n11664), .C2(n10039), .A(n14920), .B(n9894), .ZN(
        n9896) );
  AOI211_X1 U12322 ( .C1(n9894), .C2(n14920), .A(n11664), .B(n9759), .ZN(n9895) );
  OAI21_X1 U12323 ( .B1(n9899), .B2(n9898), .A(n9925), .ZN(n9900) );
  NAND2_X1 U12324 ( .A1(n9900), .A2(n12346), .ZN(n9903) );
  OAI22_X1 U12325 ( .A1(n14920), .A2(n12361), .B1(n12354), .B2(n14927), .ZN(
        n9901) );
  AOI21_X1 U12326 ( .B1(n12357), .B2(n12383), .A(n9901), .ZN(n9902) );
  OAI211_X1 U12327 ( .C1(n9905), .C2(n9904), .A(n9903), .B(n9902), .ZN(
        P3_U3177) );
  INV_X1 U12328 ( .A(n14447), .ZN(n10975) );
  OAI222_X1 U12329 ( .A1(n14135), .A2(n9907), .B1(n12134), .B2(n9906), .C1(
        n10975), .C2(P1_U3086), .ZN(P1_U3340) );
  INV_X1 U12330 ( .A(n9908), .ZN(n9910) );
  INV_X1 U12331 ( .A(SI_17_), .ZN(n9909) );
  OAI222_X1 U12332 ( .A1(n12510), .A2(P3_U3151), .B1(n12886), .B2(n9910), .C1(
        n9909), .C2(n12883), .ZN(P3_U3278) );
  AOI21_X1 U12333 ( .B1(n10719), .B2(P2_REG2_REG_13__SCAN_IN), .A(n9911), .ZN(
        n10345) );
  XNOR2_X1 U12334 ( .A(n10345), .B(n11114), .ZN(n10346) );
  XNOR2_X1 U12335 ( .A(n10346), .B(P2_REG2_REG_14__SCAN_IN), .ZN(n9922) );
  NAND2_X1 U12336 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n11140)
         );
  INV_X1 U12337 ( .A(n11140), .ZN(n9913) );
  INV_X1 U12338 ( .A(n11114), .ZN(n10344) );
  NOR2_X1 U12339 ( .A1(n14618), .A2(n10344), .ZN(n9912) );
  AOI211_X1 U12340 ( .C1(n14610), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n9913), .B(
        n9912), .ZN(n9921) );
  INV_X1 U12341 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9914) );
  XNOR2_X1 U12342 ( .A(n11114), .B(n9914), .ZN(n9919) );
  NAND2_X1 U12343 ( .A1(n10719), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n9915) );
  NAND2_X1 U12344 ( .A1(n9916), .A2(n9915), .ZN(n9918) );
  INV_X1 U12345 ( .A(n10339), .ZN(n9917) );
  OAI211_X1 U12346 ( .C1(n9919), .C2(n9918), .A(n9917), .B(n14586), .ZN(n9920)
         );
  OAI211_X1 U12347 ( .C1(n9922), .C2(n14614), .A(n9921), .B(n9920), .ZN(
        P2_U3228) );
  INV_X1 U12348 ( .A(n12358), .ZN(n10381) );
  NAND2_X1 U12349 ( .A1(n10141), .A2(n9923), .ZN(n9924) );
  AND2_X1 U12350 ( .A1(n9925), .A2(n9924), .ZN(n9927) );
  XNOR2_X1 U12351 ( .A(n10148), .B(n11664), .ZN(n10019) );
  XNOR2_X1 U12352 ( .A(n14918), .B(n10019), .ZN(n9926) );
  OAI211_X1 U12353 ( .C1(n9927), .C2(n9926), .A(n12346), .B(n10020), .ZN(n9930) );
  NOR2_X1 U12354 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10149), .ZN(n14768) );
  OAI22_X1 U12355 ( .A1(n10141), .A2(n12361), .B1(n10164), .B2(n12341), .ZN(
        n9928) );
  AOI211_X1 U12356 ( .C1(n12364), .C2(n10148), .A(n14768), .B(n9928), .ZN(
        n9929) );
  OAI211_X1 U12357 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n10381), .A(n9930), .B(
        n9929), .ZN(P3_U3158) );
  INV_X1 U12358 ( .A(n12537), .ZN(n9934) );
  INV_X1 U12359 ( .A(n9931), .ZN(n9933) );
  INV_X1 U12360 ( .A(SI_18_), .ZN(n9932) );
  OAI222_X1 U12361 ( .A1(n9934), .A2(P3_U3151), .B1(n12886), .B2(n9933), .C1(
        n9932), .C2(n12883), .ZN(P3_U3277) );
  OAI21_X1 U12362 ( .B1(n9936), .B2(P1_REG1_REG_12__SCAN_IN), .A(n9935), .ZN(
        n9939) );
  INV_X1 U12363 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9937) );
  MUX2_X1 U12364 ( .A(n9937), .B(P1_REG1_REG_13__SCAN_IN), .S(n10055), .Z(
        n9938) );
  NOR2_X1 U12365 ( .A1(n9939), .A2(n9938), .ZN(n10047) );
  AOI211_X1 U12366 ( .C1(n9939), .C2(n9938), .A(n10047), .B(n13764), .ZN(n9950) );
  INV_X1 U12367 ( .A(n10055), .ZN(n9948) );
  AOI21_X1 U12368 ( .B1(n9734), .B2(n9941), .A(n9940), .ZN(n9944) );
  INV_X1 U12369 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9942) );
  MUX2_X1 U12370 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n9942), .S(n10055), .Z(
        n9943) );
  NAND2_X1 U12371 ( .A1(n9943), .A2(n9944), .ZN(n10053) );
  OAI211_X1 U12372 ( .C1(n9944), .C2(n9943), .A(n13766), .B(n10053), .ZN(n9947) );
  NAND2_X1 U12373 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n11624)
         );
  INV_X1 U12374 ( .A(n11624), .ZN(n9945) );
  AOI21_X1 U12375 ( .B1(n13725), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n9945), .ZN(
        n9946) );
  OAI211_X1 U12376 ( .C1(n13722), .C2(n9948), .A(n9947), .B(n9946), .ZN(n9949)
         );
  OR2_X1 U12377 ( .A1(n9950), .A2(n9949), .ZN(P1_U3256) );
  NAND2_X1 U12378 ( .A1(n9952), .A2(n9951), .ZN(n9955) );
  AOI22_X1 U12379 ( .A1(n12001), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n11898), 
        .B2(n9953), .ZN(n9954) );
  NAND2_X1 U12380 ( .A1(n9955), .A2(n9954), .ZN(n14710) );
  XNOR2_X1 U12381 ( .A(n14710), .B(n12911), .ZN(n9956) );
  NAND2_X1 U12382 ( .A1(n13057), .A2(n9633), .ZN(n9957) );
  NAND2_X1 U12383 ( .A1(n9956), .A2(n9957), .ZN(n10076) );
  INV_X1 U12384 ( .A(n9956), .ZN(n9959) );
  INV_X1 U12385 ( .A(n9957), .ZN(n9958) );
  NAND2_X1 U12386 ( .A1(n9959), .A2(n9958), .ZN(n10078) );
  NAND2_X1 U12387 ( .A1(n10076), .A2(n10078), .ZN(n9967) );
  INV_X1 U12388 ( .A(n9962), .ZN(n9963) );
  NAND2_X1 U12389 ( .A1(n9964), .A2(n9963), .ZN(n9965) );
  NAND2_X1 U12390 ( .A1(n9966), .A2(n9965), .ZN(n10077) );
  XOR2_X1 U12391 ( .A(n9967), .B(n10077), .Z(n9981) );
  NAND2_X1 U12392 ( .A1(n13058), .A2(n13004), .ZN(n9976) );
  NAND2_X1 U12393 ( .A1(n11971), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n9974) );
  NAND2_X1 U12394 ( .A1(n9628), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n9973) );
  NAND2_X1 U12395 ( .A1(n9969), .A2(n9968), .ZN(n9970) );
  AND2_X1 U12396 ( .A1(n10085), .A2(n9970), .ZN(n10084) );
  NAND2_X1 U12397 ( .A1(n7325), .A2(n10084), .ZN(n9972) );
  NAND2_X1 U12398 ( .A1(n9624), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n9971) );
  NAND4_X1 U12399 ( .A1(n9974), .A2(n9973), .A3(n9972), .A4(n9971), .ZN(n13056) );
  NAND2_X1 U12400 ( .A1(n13056), .A2(n12987), .ZN(n9975) );
  AND2_X1 U12401 ( .A1(n9976), .A2(n9975), .ZN(n10712) );
  NAND2_X1 U12402 ( .A1(n13025), .A2(n10707), .ZN(n9978) );
  OAI211_X1 U12403 ( .C1(n10712), .C2(n13015), .A(n9978), .B(n9977), .ZN(n9979) );
  AOI21_X1 U12404 ( .B1(n14710), .B2(n13026), .A(n9979), .ZN(n9980) );
  OAI21_X1 U12405 ( .B1(n9981), .B2(n13018), .A(n9980), .ZN(P2_U3193) );
  OAI222_X1 U12406 ( .A1(P3_U3151), .A2(n12543), .B1(n12886), .B2(n9983), .C1(
        n9982), .C2(n12883), .ZN(P3_U3276) );
  NAND2_X1 U12407 ( .A1(n7112), .A2(n11814), .ZN(n9985) );
  XNOR2_X1 U12408 ( .A(n13062), .B(n14634), .ZN(n11818) );
  INV_X1 U12409 ( .A(n11818), .ZN(n14639) );
  NAND2_X1 U12410 ( .A1(n14632), .A2(n14639), .ZN(n9987) );
  INV_X1 U12411 ( .A(n13062), .ZN(n9995) );
  NAND2_X1 U12412 ( .A1(n9995), .A2(n14677), .ZN(n9986) );
  XNOR2_X1 U12413 ( .A(n9997), .B(n14683), .ZN(n12027) );
  NAND2_X1 U12414 ( .A1(n10206), .A2(n9997), .ZN(n9988) );
  NAND2_X1 U12415 ( .A1(n14690), .A2(n13060), .ZN(n9989) );
  XNOR2_X1 U12416 ( .A(n14702), .B(n13059), .ZN(n12029) );
  OR2_X1 U12417 ( .A1(n14702), .A2(n13059), .ZN(n9990) );
  XNOR2_X1 U12418 ( .A(n14619), .B(n13058), .ZN(n12032) );
  INV_X1 U12419 ( .A(n12032), .ZN(n9991) );
  OAI21_X1 U12420 ( .B1(n9992), .B2(n9991), .A(n10258), .ZN(n14629) );
  INV_X1 U12421 ( .A(n14629), .ZN(n10010) );
  NAND2_X1 U12422 ( .A1(n7112), .A2(n11813), .ZN(n14638) );
  NAND2_X1 U12423 ( .A1(n9993), .A2(n14638), .ZN(n9994) );
  NAND2_X1 U12424 ( .A1(n9994), .A2(n11818), .ZN(n14642) );
  NAND2_X1 U12425 ( .A1(n9995), .A2(n14634), .ZN(n9996) );
  NAND2_X1 U12426 ( .A1(n14642), .A2(n9996), .ZN(n10199) );
  INV_X1 U12427 ( .A(n12027), .ZN(n10198) );
  NAND2_X1 U12428 ( .A1(n10199), .A2(n10198), .ZN(n10197) );
  NAND2_X1 U12429 ( .A1(n9997), .A2(n14683), .ZN(n9998) );
  NAND2_X1 U12430 ( .A1(n10197), .A2(n9998), .ZN(n10185) );
  INV_X1 U12431 ( .A(n13060), .ZN(n10000) );
  OR2_X1 U12432 ( .A1(n10000), .A2(n14690), .ZN(n9999) );
  NAND2_X1 U12433 ( .A1(n10185), .A2(n9999), .ZN(n10002) );
  NAND2_X1 U12434 ( .A1(n14690), .A2(n10000), .ZN(n10001) );
  NAND2_X1 U12435 ( .A1(n10002), .A2(n10001), .ZN(n10696) );
  NAND2_X1 U12436 ( .A1(n10696), .A2(n12029), .ZN(n10005) );
  INV_X1 U12437 ( .A(n13059), .ZN(n10003) );
  NAND2_X1 U12438 ( .A1(n14702), .A2(n10003), .ZN(n10004) );
  NAND2_X1 U12439 ( .A1(n10005), .A2(n10004), .ZN(n10263) );
  XNOR2_X1 U12440 ( .A(n10263), .B(n12032), .ZN(n10007) );
  AOI21_X1 U12441 ( .B1(n10007), .B2(n13391), .A(n10006), .ZN(n14631) );
  INV_X1 U12442 ( .A(n14702), .ZN(n10694) );
  NAND2_X1 U12443 ( .A1(n10689), .A2(n10694), .ZN(n10690) );
  OR2_X1 U12444 ( .A1(n10690), .A2(n14619), .ZN(n10706) );
  INV_X1 U12445 ( .A(n10706), .ZN(n10008) );
  AOI211_X1 U12446 ( .C1(n14619), .C2(n10690), .A(n14633), .B(n10008), .ZN(
        n14620) );
  AOI21_X1 U12447 ( .B1(n14711), .B2(n14619), .A(n14620), .ZN(n10009) );
  OAI211_X1 U12448 ( .C1(n10010), .C2(n13495), .A(n14631), .B(n10009), .ZN(
        n10016) );
  NAND2_X1 U12449 ( .A1(n10016), .A2(n14746), .ZN(n10011) );
  OAI21_X1 U12450 ( .B1(n14746), .B2(n10012), .A(n10011), .ZN(P2_U3506) );
  INV_X1 U12451 ( .A(n10013), .ZN(n10015) );
  AND2_X1 U12452 ( .A1(n14658), .A2(n10014), .ZN(n10170) );
  INV_X1 U12453 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10018) );
  NAND2_X1 U12454 ( .A1(n10016), .A2(n14731), .ZN(n10017) );
  OAI21_X1 U12455 ( .B1(n14731), .B2(n10018), .A(n10017), .ZN(P2_U3451) );
  INV_X1 U12456 ( .A(n10019), .ZN(n10021) );
  OAI21_X1 U12457 ( .B1(n14918), .B2(n10021), .A(n10020), .ZN(n10024) );
  XNOR2_X1 U12458 ( .A(n14958), .B(n11698), .ZN(n10022) );
  NAND2_X1 U12459 ( .A1(n10164), .A2(n10022), .ZN(n10159) );
  OAI21_X1 U12460 ( .B1(n10164), .B2(n10022), .A(n10159), .ZN(n10023) );
  AOI21_X1 U12461 ( .B1(n10024), .B2(n10023), .A(n10161), .ZN(n10029) );
  NOR2_X1 U12462 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10025), .ZN(n14785) );
  OAI22_X1 U12463 ( .A1(n10520), .A2(n12341), .B1(n14918), .B2(n12361), .ZN(
        n10026) );
  AOI211_X1 U12464 ( .C1(n12364), .C2(n14958), .A(n14785), .B(n10026), .ZN(
        n10028) );
  NAND2_X1 U12465 ( .A1(n12358), .A2(n10235), .ZN(n10027) );
  OAI211_X1 U12466 ( .C1(n10029), .C2(n12366), .A(n10028), .B(n10027), .ZN(
        P3_U3170) );
  XNOR2_X1 U12467 ( .A(n10032), .B(n10031), .ZN(n10033) );
  NAND3_X1 U12468 ( .A1(n10035), .A2(n10034), .A3(n10033), .ZN(n10037) );
  MUX2_X1 U12469 ( .A(n10036), .B(P3_REG2_REG_0__SCAN_IN), .S(n14944), .Z(
        n10041) );
  OR2_X1 U12470 ( .A1(n10037), .A2(n14929), .ZN(n11002) );
  INV_X1 U12471 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10038) );
  OAI22_X1 U12472 ( .A1(n14294), .A2(n10039), .B1(n14292), .B2(n10038), .ZN(
        n10040) );
  OR2_X1 U12473 ( .A1(n10041), .A2(n10040), .ZN(P3_U3233) );
  INV_X1 U12474 ( .A(n11539), .ZN(n10045) );
  OAI21_X1 U12475 ( .B1(n10042), .B2(P2_IR_REG_17__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n10043) );
  XNOR2_X1 U12476 ( .A(n10043), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13147) );
  INV_X1 U12477 ( .A(n13147), .ZN(n14617) );
  OAI222_X1 U12478 ( .A1(n13523), .A2(n10044), .B1(n13526), .B2(n10045), .C1(
        P2_U3088), .C2(n14617), .ZN(P2_U3309) );
  INV_X1 U12479 ( .A(n13759), .ZN(n13754) );
  OAI222_X1 U12480 ( .A1(n14135), .A2(n10046), .B1(n12134), .B2(n10045), .C1(
        P1_U3086), .C2(n13754), .ZN(P1_U3337) );
  INV_X1 U12481 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n10048) );
  MUX2_X1 U12482 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10048), .S(n10973), .Z(
        n10049) );
  OAI21_X1 U12483 ( .B1(n10050), .B2(n10049), .A(n10972), .ZN(n10060) );
  NAND2_X1 U12484 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14348)
         );
  INV_X1 U12485 ( .A(n14348), .ZN(n10051) );
  AOI21_X1 U12486 ( .B1(n13725), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n10051), 
        .ZN(n10052) );
  OAI21_X1 U12487 ( .B1(n13722), .B2(n10964), .A(n10052), .ZN(n10059) );
  INV_X1 U12488 ( .A(n10053), .ZN(n10054) );
  AOI21_X1 U12489 ( .B1(n10055), .B2(P1_REG2_REG_13__SCAN_IN), .A(n10054), 
        .ZN(n10057) );
  INV_X1 U12490 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11180) );
  MUX2_X1 U12491 ( .A(n11180), .B(P1_REG2_REG_14__SCAN_IN), .S(n10973), .Z(
        n10056) );
  NOR2_X1 U12492 ( .A1(n10056), .A2(n10057), .ZN(n10962) );
  AOI211_X1 U12493 ( .C1(n10057), .C2(n10056), .A(n14451), .B(n10962), .ZN(
        n10058) );
  AOI211_X1 U12494 ( .C1(n14445), .C2(n10060), .A(n10059), .B(n10058), .ZN(
        n10061) );
  INV_X1 U12495 ( .A(n10061), .ZN(P1_U3257) );
  INV_X1 U12496 ( .A(n11897), .ZN(n11636) );
  OAI222_X1 U12497 ( .A1(n14135), .A2(n10063), .B1(n12134), .B2(n11636), .C1(
        P1_U3086), .C2(n10062), .ZN(P1_U3336) );
  OR2_X1 U12498 ( .A1(n10064), .A2(n9394), .ZN(n10070) );
  OAI22_X1 U12499 ( .A1(n11980), .A2(n10067), .B1(n10066), .B2(n10065), .ZN(
        n10068) );
  INV_X1 U12500 ( .A(n10068), .ZN(n10069) );
  XNOR2_X1 U12501 ( .A(n11848), .B(n12911), .ZN(n10071) );
  NAND2_X1 U12502 ( .A1(n13056), .A2(n9633), .ZN(n10072) );
  NAND2_X1 U12503 ( .A1(n10071), .A2(n10072), .ZN(n10119) );
  INV_X1 U12504 ( .A(n10071), .ZN(n10074) );
  INV_X1 U12505 ( .A(n10072), .ZN(n10073) );
  NAND2_X1 U12506 ( .A1(n10074), .A2(n10073), .ZN(n10075) );
  NAND2_X1 U12507 ( .A1(n10119), .A2(n10075), .ZN(n10083) );
  INV_X1 U12508 ( .A(n10083), .ZN(n10080) );
  INV_X1 U12509 ( .A(n10120), .ZN(n10081) );
  AOI21_X1 U12510 ( .B1(n10083), .B2(n10082), .A(n10081), .ZN(n10097) );
  INV_X1 U12511 ( .A(n10084), .ZN(n10561) );
  NAND2_X1 U12512 ( .A1(n13057), .A2(n13004), .ZN(n10092) );
  NAND2_X1 U12513 ( .A1(n9624), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n10090) );
  NAND2_X1 U12514 ( .A1(n11971), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10089) );
  NAND2_X1 U12515 ( .A1(n10085), .A2(n14585), .ZN(n10086) );
  AND2_X1 U12516 ( .A1(n10127), .A2(n10086), .ZN(n10124) );
  NAND2_X1 U12517 ( .A1(n7325), .A2(n10124), .ZN(n10088) );
  NAND2_X1 U12518 ( .A1(n9628), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n10087) );
  NAND4_X1 U12519 ( .A1(n10090), .A2(n10089), .A3(n10088), .A4(n10087), .ZN(
        n13055) );
  NAND2_X1 U12520 ( .A1(n13055), .A2(n13164), .ZN(n10091) );
  NAND2_X1 U12521 ( .A1(n10092), .A2(n10091), .ZN(n10266) );
  NAND2_X1 U12522 ( .A1(n13040), .A2(n10266), .ZN(n10093) );
  OAI211_X1 U12523 ( .C1(n13038), .C2(n10561), .A(n10094), .B(n10093), .ZN(
        n10095) );
  AOI21_X1 U12524 ( .B1(n11848), .B2(n13026), .A(n10095), .ZN(n10096) );
  OAI21_X1 U12525 ( .B1(n10097), .B2(n13018), .A(n10096), .ZN(P2_U3203) );
  OAI22_X1 U12526 ( .A1(n9817), .A2(n12264), .B1(n14512), .B2(n12263), .ZN(
        n10100) );
  XNOR2_X1 U12527 ( .A(n10100), .B(n10099), .ZN(n10106) );
  OR2_X1 U12528 ( .A1(n9817), .A2(n9810), .ZN(n10102) );
  NAND2_X1 U12529 ( .A1(n12247), .A2(n14486), .ZN(n10101) );
  NAND2_X1 U12530 ( .A1(n10102), .A2(n10101), .ZN(n10107) );
  XNOR2_X1 U12531 ( .A(n10106), .B(n10107), .ZN(n13543) );
  NOR2_X1 U12532 ( .A1(n10104), .A2(n10103), .ZN(n13544) );
  AOI22_X1 U12533 ( .A1(n12259), .A2(n13676), .B1(n12247), .B2(n14521), .ZN(
        n10240) );
  NAND2_X1 U12534 ( .A1(n13676), .A2(n12247), .ZN(n10109) );
  NAND2_X1 U12535 ( .A1(n12255), .A2(n14521), .ZN(n10108) );
  NAND2_X1 U12536 ( .A1(n10109), .A2(n10108), .ZN(n10110) );
  XNOR2_X1 U12537 ( .A(n10110), .B(n10099), .ZN(n10242) );
  XNOR2_X1 U12538 ( .A(n10243), .B(n10242), .ZN(n10118) );
  INV_X1 U12539 ( .A(n14394), .ZN(n13649) );
  INV_X1 U12540 ( .A(n14389), .ZN(n13653) );
  OR2_X1 U12541 ( .A1(n9817), .A2(n13982), .ZN(n10113) );
  NAND2_X1 U12542 ( .A1(n13674), .A2(n13955), .ZN(n10112) );
  NAND2_X1 U12543 ( .A1(n10113), .A2(n10112), .ZN(n14520) );
  NAND2_X1 U12544 ( .A1(n14358), .A2(n14520), .ZN(n10115) );
  OAI211_X1 U12545 ( .C1(n13653), .C2(n10615), .A(n10115), .B(n10114), .ZN(
        n10116) );
  AOI21_X1 U12546 ( .B1(n10616), .B2(n13649), .A(n10116), .ZN(n10117) );
  OAI21_X1 U12547 ( .B1(n10118), .B2(n14384), .A(n10117), .ZN(P1_U3230) );
  OR2_X1 U12548 ( .A1(n10121), .A2(n9394), .ZN(n10123) );
  AOI22_X1 U12549 ( .A1(n12001), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n11898), 
        .B2(n14593), .ZN(n10122) );
  XNOR2_X1 U12550 ( .A(n14720), .B(n12911), .ZN(n10353) );
  NAND2_X1 U12551 ( .A1(n13055), .A2(n9633), .ZN(n10352) );
  XNOR2_X1 U12552 ( .A(n10353), .B(n10352), .ZN(n10354) );
  XNOR2_X1 U12553 ( .A(n10355), .B(n10354), .ZN(n10138) );
  INV_X1 U12554 ( .A(n10124), .ZN(n10549) );
  NAND2_X1 U12555 ( .A1(n13056), .A2(n13004), .ZN(n10134) );
  NAND2_X1 U12556 ( .A1(n11971), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n10132) );
  NAND2_X1 U12557 ( .A1(n10125), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n10361) );
  INV_X1 U12558 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10126) );
  NAND2_X1 U12559 ( .A1(n10127), .A2(n10126), .ZN(n10128) );
  AND2_X1 U12560 ( .A1(n10361), .A2(n10128), .ZN(n10775) );
  NAND2_X1 U12561 ( .A1(n7325), .A2(n10775), .ZN(n10131) );
  NAND2_X1 U12562 ( .A1(n9628), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n10130) );
  NAND2_X1 U12563 ( .A1(n9624), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n10129) );
  NAND4_X1 U12564 ( .A1(n10132), .A2(n10131), .A3(n10130), .A4(n10129), .ZN(
        n13054) );
  NAND2_X1 U12565 ( .A1(n13054), .A2(n13164), .ZN(n10133) );
  NAND2_X1 U12566 ( .A1(n10134), .A2(n10133), .ZN(n10545) );
  AOI22_X1 U12567 ( .A1(n13040), .A2(n10545), .B1(P2_REG3_REG_10__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10135) );
  OAI21_X1 U12568 ( .B1(n13038), .B2(n10549), .A(n10135), .ZN(n10136) );
  AOI21_X1 U12569 ( .B1(n14720), .B2(n13026), .A(n10136), .ZN(n10137) );
  OAI21_X1 U12570 ( .B1(n10138), .B2(n13018), .A(n10137), .ZN(P2_U3189) );
  XNOR2_X1 U12571 ( .A(n10145), .B(n10139), .ZN(n14955) );
  INV_X1 U12572 ( .A(n14955), .ZN(n10152) );
  AND2_X1 U12573 ( .A1(n14929), .A2(n10140), .ZN(n14926) );
  INV_X1 U12574 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10881) );
  OAI22_X1 U12575 ( .A1(n10141), .A2(n14919), .B1(n10164), .B2(n14917), .ZN(
        n10147) );
  INV_X1 U12576 ( .A(n10142), .ZN(n10143) );
  AOI211_X1 U12577 ( .C1(n10145), .C2(n10144), .A(n14303), .B(n10143), .ZN(
        n10146) );
  AOI211_X1 U12578 ( .C1(n14955), .C2(n12804), .A(n10147), .B(n10146), .ZN(
        n14952) );
  MUX2_X1 U12579 ( .A(n10881), .B(n14952), .S(n14942), .Z(n10151) );
  AND2_X1 U12580 ( .A1(n10148), .A2(n14957), .ZN(n14954) );
  AOI22_X1 U12581 ( .A1(n14310), .A2(n14954), .B1(n14938), .B2(n10149), .ZN(
        n10150) );
  OAI211_X1 U12582 ( .C1(n10152), .C2(n12607), .A(n10151), .B(n10150), .ZN(
        P3_U3230) );
  INV_X1 U12583 ( .A(n10153), .ZN(n10154) );
  NOR2_X1 U12584 ( .A1(n10302), .A2(n10154), .ZN(n10155) );
  INV_X1 U12585 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n15038) );
  NAND2_X1 U12586 ( .A1(n10157), .A2(n14532), .ZN(n10158) );
  OAI21_X1 U12587 ( .B1(n14532), .B2(n15038), .A(n10158), .ZN(P1_U3459) );
  INV_X1 U12588 ( .A(n10159), .ZN(n10160) );
  XNOR2_X1 U12589 ( .A(n10166), .B(n11698), .ZN(n10374) );
  XNOR2_X1 U12590 ( .A(n10520), .B(n10374), .ZN(n10162) );
  AOI21_X1 U12591 ( .B1(n10163), .B2(n10162), .A(n6601), .ZN(n10169) );
  AND2_X1 U12592 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n14804) );
  OAI22_X1 U12593 ( .A1(n10485), .A2(n12341), .B1(n10164), .B2(n12361), .ZN(
        n10165) );
  AOI211_X1 U12594 ( .C1(n12364), .C2(n10166), .A(n14804), .B(n10165), .ZN(
        n10168) );
  NAND2_X1 U12595 ( .A1(n12358), .A2(n10220), .ZN(n10167) );
  OAI211_X1 U12596 ( .C1(n10169), .C2(n12366), .A(n10168), .B(n10167), .ZN(
        P3_U3167) );
  NAND3_X1 U12597 ( .A1(n10171), .A2(n14661), .A3(n10170), .ZN(n10172) );
  AOI21_X1 U12598 ( .B1(n12024), .B2(n13330), .A(n13395), .ZN(n10183) );
  NAND2_X1 U12599 ( .A1(n11802), .A2(n10173), .ZN(n14662) );
  NAND2_X1 U12600 ( .A1(n11799), .A2(n11798), .ZN(n10174) );
  NAND2_X1 U12601 ( .A1(n10175), .A2(n10174), .ZN(n12023) );
  INV_X1 U12602 ( .A(n12023), .ZN(n14665) );
  NAND2_X1 U12603 ( .A1(n10176), .A2(n11803), .ZN(n11719) );
  INV_X1 U12604 ( .A(n11719), .ZN(n10177) );
  NAND2_X1 U12605 ( .A1(n13330), .A2(n10177), .ZN(n10830) );
  INV_X1 U12606 ( .A(n10830), .ZN(n10327) );
  NOR2_X1 U12607 ( .A1(n13391), .A2(n14728), .ZN(n10179) );
  OAI21_X1 U12608 ( .B1(n12023), .B2(n10179), .A(n10178), .ZN(n14663) );
  INV_X1 U12609 ( .A(n14646), .ZN(n14621) );
  AOI22_X1 U12610 ( .A1(n13330), .A2(n14663), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n14621), .ZN(n10180) );
  OAI21_X1 U12611 ( .B1(n14548), .B2(n13330), .A(n10180), .ZN(n10181) );
  AOI21_X1 U12612 ( .B1(n14665), .B2(n10327), .A(n10181), .ZN(n10182) );
  OAI21_X1 U12613 ( .B1(n10183), .B2(n14662), .A(n10182), .ZN(P2_U3265) );
  NAND2_X1 U12614 ( .A1(n14693), .A2(n11719), .ZN(n14650) );
  XNOR2_X1 U12615 ( .A(n14690), .B(n13060), .ZN(n12030) );
  XNOR2_X1 U12616 ( .A(n10184), .B(n12030), .ZN(n14694) );
  XNOR2_X1 U12617 ( .A(n10185), .B(n12030), .ZN(n10187) );
  AOI21_X1 U12618 ( .B1(n10187), .B2(n13391), .A(n10186), .ZN(n14698) );
  MUX2_X1 U12619 ( .A(n9128), .B(n14698), .S(n13330), .Z(n10195) );
  OAI21_X1 U12620 ( .B1(n10203), .B2(n10192), .A(n13300), .ZN(n10188) );
  NOR2_X1 U12621 ( .A1(n10188), .A2(n10689), .ZN(n14692) );
  INV_X1 U12622 ( .A(n14645), .ZN(n10189) );
  NAND2_X2 U12623 ( .A1(n13330), .A2(n10189), .ZN(n14625) );
  INV_X1 U12624 ( .A(n10190), .ZN(n10191) );
  OAI22_X1 U12625 ( .A1(n14625), .A2(n10192), .B1(n14646), .B2(n10191), .ZN(
        n10193) );
  AOI21_X1 U12626 ( .B1(n13395), .B2(n14692), .A(n10193), .ZN(n10194) );
  OAI211_X1 U12627 ( .C1(n13397), .C2(n14694), .A(n10195), .B(n10194), .ZN(
        P2_U3260) );
  XNOR2_X1 U12628 ( .A(n10196), .B(n10198), .ZN(n14686) );
  OAI21_X1 U12629 ( .B1(n10199), .B2(n10198), .A(n10197), .ZN(n10201) );
  AOI21_X1 U12630 ( .B1(n10201), .B2(n13391), .A(n10200), .ZN(n14685) );
  MUX2_X1 U12631 ( .A(n10202), .B(n14685), .S(n13330), .Z(n10209) );
  AOI211_X1 U12632 ( .C1(n14683), .C2(n14636), .A(n14633), .B(n10203), .ZN(
        n14682) );
  INV_X1 U12633 ( .A(n10204), .ZN(n10205) );
  OAI22_X1 U12634 ( .A1(n14625), .A2(n10206), .B1(n10205), .B2(n14646), .ZN(
        n10207) );
  AOI21_X1 U12635 ( .B1(n13395), .B2(n14682), .A(n10207), .ZN(n10208) );
  OAI211_X1 U12636 ( .C1(n13397), .C2(n14686), .A(n10209), .B(n10208), .ZN(
        P2_U3261) );
  INV_X1 U12637 ( .A(n10210), .ZN(n10211) );
  AOI21_X1 U12638 ( .B1(n10214), .B2(n10212), .A(n10211), .ZN(n10218) );
  AOI22_X1 U12639 ( .A1(n14284), .A2(n12380), .B1(n12382), .B2(n14286), .ZN(
        n10217) );
  NAND2_X1 U12640 ( .A1(n10514), .A2(n10230), .ZN(n10228) );
  NAND2_X1 U12641 ( .A1(n10228), .A2(n10213), .ZN(n10215) );
  XNOR2_X1 U12642 ( .A(n10215), .B(n10214), .ZN(n14965) );
  NAND2_X1 U12643 ( .A1(n14965), .A2(n12804), .ZN(n10216) );
  OAI211_X1 U12644 ( .C1(n10218), .C2(n14303), .A(n10217), .B(n10216), .ZN(
        n14963) );
  INV_X1 U12645 ( .A(n14963), .ZN(n10224) );
  INV_X1 U12646 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n14795) );
  NOR2_X1 U12647 ( .A1(n10219), .A2(n14979), .ZN(n14964) );
  AOI22_X1 U12648 ( .A1(n14964), .A2(n14310), .B1(n14938), .B2(n10220), .ZN(
        n10221) );
  OAI21_X1 U12649 ( .B1(n14795), .B2(n14942), .A(n10221), .ZN(n10222) );
  AOI21_X1 U12650 ( .B1(n14965), .B2(n14939), .A(n10222), .ZN(n10223) );
  OAI21_X1 U12651 ( .B1(n10224), .B2(n14944), .A(n10223), .ZN(P3_U3228) );
  OAI222_X1 U12652 ( .A1(n12886), .A2(n10226), .B1(n12883), .B2(n15098), .C1(
        P3_U3151), .C2(n10225), .ZN(P3_U3275) );
  OR2_X1 U12653 ( .A1(n10514), .A2(n10230), .ZN(n10227) );
  NAND2_X1 U12654 ( .A1(n10228), .A2(n10227), .ZN(n14959) );
  INV_X1 U12655 ( .A(n14959), .ZN(n10238) );
  INV_X1 U12656 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10886) );
  OAI22_X1 U12657 ( .A1(n10520), .A2(n14917), .B1(n14918), .B2(n14919), .ZN(
        n10229) );
  AOI21_X1 U12658 ( .B1(n14959), .B2(n12804), .A(n10229), .ZN(n10234) );
  XNOR2_X1 U12659 ( .A(n10231), .B(n10230), .ZN(n10232) );
  NAND2_X1 U12660 ( .A1(n10232), .A2(n14922), .ZN(n10233) );
  AND2_X1 U12661 ( .A1(n10234), .A2(n10233), .ZN(n14961) );
  MUX2_X1 U12662 ( .A(n10886), .B(n14961), .S(n14942), .Z(n10237) );
  INV_X1 U12663 ( .A(n14294), .ZN(n12604) );
  AOI22_X1 U12664 ( .A1(n12604), .A2(n14958), .B1(n14938), .B2(n10235), .ZN(
        n10236) );
  OAI211_X1 U12665 ( .C1(n10238), .C2(n12607), .A(n10237), .B(n10236), .ZN(
        P3_U3229) );
  NAND2_X1 U12666 ( .A1(n14467), .A2(n12255), .ZN(n10245) );
  NAND2_X1 U12667 ( .A1(n13674), .A2(n12247), .ZN(n10244) );
  NAND2_X1 U12668 ( .A1(n10245), .A2(n10244), .ZN(n10246) );
  XNOR2_X1 U12669 ( .A(n10246), .B(n12177), .ZN(n10248) );
  AOI22_X1 U12670 ( .A1(n12259), .A2(n13674), .B1(n12247), .B2(n14467), .ZN(
        n10247) );
  OR2_X1 U12671 ( .A1(n10248), .A2(n10247), .ZN(n10600) );
  NAND2_X1 U12672 ( .A1(n6484), .A2(n10600), .ZN(n10249) );
  XNOR2_X1 U12673 ( .A(n6606), .B(n10249), .ZN(n10256) );
  NAND2_X1 U12674 ( .A1(n13676), .A2(n13954), .ZN(n10251) );
  NAND2_X1 U12675 ( .A1(n13673), .A2(n13955), .ZN(n10250) );
  NAND2_X1 U12676 ( .A1(n10251), .A2(n10250), .ZN(n10477) );
  NAND2_X1 U12677 ( .A1(n14358), .A2(n10477), .ZN(n10253) );
  OAI211_X1 U12678 ( .C1(n13653), .C2(n6954), .A(n10253), .B(n10252), .ZN(
        n10254) );
  AOI21_X1 U12679 ( .B1(n14465), .B2(n13649), .A(n10254), .ZN(n10255) );
  OAI21_X1 U12680 ( .B1(n10256), .B2(n14384), .A(n10255), .ZN(P1_U3227) );
  INV_X1 U12681 ( .A(n13495), .ZN(n14680) );
  OR2_X1 U12682 ( .A1(n14619), .A2(n13058), .ZN(n10257) );
  XNOR2_X1 U12683 ( .A(n14710), .B(n13057), .ZN(n12035) );
  NAND2_X1 U12684 ( .A1(n14710), .A2(n13057), .ZN(n10259) );
  NAND2_X1 U12685 ( .A1(n10702), .A2(n10259), .ZN(n10538) );
  INV_X1 U12686 ( .A(n13056), .ZN(n10541) );
  XNOR2_X1 U12687 ( .A(n11848), .B(n10541), .ZN(n12034) );
  XOR2_X1 U12688 ( .A(n10538), .B(n12034), .Z(n10559) );
  INV_X1 U12689 ( .A(n11848), .ZN(n10268) );
  INV_X1 U12690 ( .A(n13058), .ZN(n10260) );
  AND2_X1 U12691 ( .A1(n14619), .A2(n10260), .ZN(n10262) );
  OR2_X1 U12692 ( .A1(n14619), .A2(n10260), .ZN(n10261) );
  INV_X1 U12693 ( .A(n13057), .ZN(n10264) );
  AOI21_X1 U12694 ( .B1(n10265), .B2(n12034), .A(n14640), .ZN(n10267) );
  AOI21_X1 U12695 ( .B1(n10267), .B2(n10542), .A(n10266), .ZN(n10560) );
  NAND2_X1 U12696 ( .A1(n10705), .A2(n10268), .ZN(n10547) );
  OAI211_X1 U12697 ( .C1(n10705), .C2(n10268), .A(n13300), .B(n10547), .ZN(
        n10564) );
  OAI211_X1 U12698 ( .C1(n10268), .C2(n14723), .A(n10560), .B(n10564), .ZN(
        n10269) );
  AOI21_X1 U12699 ( .B1(n14680), .B2(n10559), .A(n10269), .ZN(n10274) );
  OR2_X1 U12700 ( .A1(n14746), .A2(n10270), .ZN(n10271) );
  OAI21_X1 U12701 ( .B1(n10274), .B2(n14744), .A(n10271), .ZN(P2_U3508) );
  INV_X1 U12702 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10272) );
  OR2_X1 U12703 ( .A1(n14731), .A2(n10272), .ZN(n10273) );
  OAI21_X1 U12704 ( .B1(n10274), .B2(n14729), .A(n10273), .ZN(P2_U3457) );
  NAND2_X1 U12705 ( .A1(n10277), .A2(n10276), .ZN(n10279) );
  NAND2_X1 U12706 ( .A1(n10279), .A2(n10278), .ZN(n10457) );
  NAND2_X1 U12707 ( .A1(n14477), .A2(n10291), .ZN(n10282) );
  NAND2_X1 U12708 ( .A1(n10282), .A2(n10281), .ZN(n10613) );
  NOR2_X1 U12709 ( .A1(n13676), .A2(n10615), .ZN(n10283) );
  AND2_X1 U12710 ( .A1(n6954), .A2(n13674), .ZN(n10284) );
  INV_X1 U12711 ( .A(n13674), .ZN(n10295) );
  NAND2_X1 U12712 ( .A1(n10295), .A2(n14467), .ZN(n10285) );
  XNOR2_X1 U12713 ( .A(n10391), .B(n10389), .ZN(n10301) );
  NAND2_X1 U12714 ( .A1(n6635), .A2(n11693), .ZN(n10286) );
  NAND2_X1 U12715 ( .A1(n10455), .A2(n10456), .ZN(n10290) );
  NAND2_X1 U12716 ( .A1(n8691), .A2(n14504), .ZN(n10289) );
  AND2_X1 U12717 ( .A1(n9817), .A2(n14512), .ZN(n10292) );
  NAND2_X1 U12718 ( .A1(n6954), .A2(n10295), .ZN(n10296) );
  NAND2_X1 U12719 ( .A1(n10471), .A2(n10296), .ZN(n10297) );
  OR2_X1 U12720 ( .A1(n10297), .A2(n10389), .ZN(n10298) );
  INV_X1 U12721 ( .A(n13855), .ZN(n14482) );
  NAND2_X1 U12722 ( .A1(n10321), .A2(n14482), .ZN(n10300) );
  AOI22_X1 U12723 ( .A1(n13954), .A2(n13674), .B1(n13672), .B2(n13955), .ZN(
        n10299) );
  OAI211_X1 U12724 ( .C1(n14478), .C2(n10301), .A(n10300), .B(n10299), .ZN(
        n10319) );
  INV_X1 U12725 ( .A(n10302), .ZN(n10309) );
  INV_X1 U12726 ( .A(n10303), .ZN(n10304) );
  OAI21_X1 U12727 ( .B1(n10305), .B2(n10304), .A(n14500), .ZN(n10306) );
  NAND4_X1 U12728 ( .A1(n10309), .A2(n10308), .A3(n10307), .A4(n10306), .ZN(
        n12148) );
  MUX2_X1 U12729 ( .A(n10319), .B(P1_REG2_REG_6__SCAN_IN), .S(n14498), .Z(
        n10310) );
  INV_X1 U12730 ( .A(n10310), .ZN(n10318) );
  INV_X1 U12731 ( .A(n10311), .ZN(n10312) );
  NAND2_X1 U12732 ( .A1(n13966), .A2(n10312), .ZN(n13865) );
  INV_X1 U12733 ( .A(n13865), .ZN(n14495) );
  INV_X1 U12734 ( .A(n10596), .ZN(n13627) );
  INV_X1 U12735 ( .A(n14483), .ZN(n14466) );
  NAND2_X1 U12736 ( .A1(n14466), .A2(n13624), .ZN(n10315) );
  OR2_X1 U12737 ( .A1(n10464), .A2(n10463), .ZN(n14488) );
  NAND2_X1 U12738 ( .A1(n14489), .A2(n10615), .ZN(n10614) );
  AOI21_X1 U12739 ( .B1(n10479), .B2(n10596), .A(n13961), .ZN(n10313) );
  AND2_X1 U12740 ( .A1(n10572), .A2(n10313), .ZN(n10320) );
  NAND2_X1 U12741 ( .A1(n10320), .A2(n14494), .ZN(n10314) );
  OAI211_X1 U12742 ( .C1(n13978), .C2(n13627), .A(n10315), .B(n10314), .ZN(
        n10316) );
  AOI21_X1 U12743 ( .B1(n10321), .B2(n14495), .A(n10316), .ZN(n10317) );
  NAND2_X1 U12744 ( .A1(n10318), .A2(n10317), .ZN(P1_U3287) );
  INV_X1 U12745 ( .A(n10480), .ZN(n14517) );
  AOI211_X1 U12746 ( .C1(n14517), .C2(n10321), .A(n10320), .B(n10319), .ZN(
        n10558) );
  OAI22_X1 U12747 ( .A1(n14084), .A2(n13627), .B1(n14540), .B2(n9204), .ZN(
        n10322) );
  INV_X1 U12748 ( .A(n10322), .ZN(n10323) );
  OAI21_X1 U12749 ( .B1(n10558), .B2(n14537), .A(n10323), .ZN(P1_U3534) );
  INV_X1 U12750 ( .A(n10324), .ZN(n10325) );
  OAI211_X1 U12751 ( .C1(n14667), .C2(n11798), .A(n10325), .B(n13300), .ZN(
        n14666) );
  XNOR2_X1 U12752 ( .A(n12026), .B(n10326), .ZN(n14670) );
  INV_X1 U12753 ( .A(n14625), .ZN(n13303) );
  AOI22_X1 U12754 ( .A1(n10327), .A2(n14670), .B1(n13303), .B2(n11806), .ZN(
        n10338) );
  INV_X1 U12755 ( .A(n14670), .ZN(n10333) );
  OAI21_X1 U12756 ( .B1(n12026), .B2(n10329), .A(n10328), .ZN(n10331) );
  AOI21_X1 U12757 ( .B1(n10331), .B2(n13391), .A(n10330), .ZN(n10332) );
  OAI21_X1 U12758 ( .B1(n10333), .B2(n14693), .A(n10332), .ZN(n14668) );
  OAI22_X1 U12759 ( .A1(n13330), .A2(n10335), .B1(n10334), .B2(n14646), .ZN(
        n10336) );
  AOI21_X1 U12760 ( .B1(n13330), .B2(n14668), .A(n10336), .ZN(n10337) );
  OAI211_X1 U12761 ( .C1(n13307), .C2(n14666), .A(n10338), .B(n10337), .ZN(
        P2_U3264) );
  INV_X1 U12762 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n11332) );
  NOR2_X1 U12763 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11332), .ZN(n10343) );
  AOI21_X1 U12764 ( .B1(n11114), .B2(P2_REG1_REG_14__SCAN_IN), .A(n10339), 
        .ZN(n10405) );
  XNOR2_X1 U12765 ( .A(n10404), .B(n10405), .ZN(n10341) );
  INV_X1 U12766 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n10340) );
  NOR2_X1 U12767 ( .A1(n10340), .A2(n10341), .ZN(n10406) );
  AOI211_X1 U12768 ( .C1(n10341), .C2(n10340), .A(n10406), .B(n14604), .ZN(
        n10342) );
  AOI211_X1 U12769 ( .C1(n14610), .C2(P2_ADDR_REG_15__SCAN_IN), .A(n10343), 
        .B(n10342), .ZN(n10351) );
  OR2_X1 U12770 ( .A1(n10345), .A2(n10344), .ZN(n10348) );
  NAND2_X1 U12771 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n10346), .ZN(n10347) );
  NAND2_X1 U12772 ( .A1(n10348), .A2(n10347), .ZN(n10410) );
  XNOR2_X1 U12773 ( .A(n10404), .B(n10410), .ZN(n10349) );
  NAND2_X1 U12774 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n10349), .ZN(n10411) );
  OAI211_X1 U12775 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n10349), .A(n14579), 
        .B(n10411), .ZN(n10350) );
  OAI211_X1 U12776 ( .C1(n14618), .C2(n10404), .A(n10351), .B(n10350), .ZN(
        P2_U3229) );
  NAND2_X1 U12777 ( .A1(n10356), .A2(n9951), .ZN(n10358) );
  AOI22_X1 U12778 ( .A1(n12001), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n11898), 
        .B2(n13132), .ZN(n10357) );
  XNOR2_X1 U12779 ( .A(n13491), .B(n12960), .ZN(n10656) );
  NAND2_X1 U12780 ( .A1(n13054), .A2(n9633), .ZN(n10654) );
  XNOR2_X1 U12781 ( .A(n10656), .B(n10654), .ZN(n10652) );
  XNOR2_X1 U12782 ( .A(n10653), .B(n10652), .ZN(n10373) );
  INV_X1 U12783 ( .A(n10775), .ZN(n10370) );
  NAND2_X1 U12784 ( .A1(n13055), .A2(n13004), .ZN(n10368) );
  NAND2_X1 U12785 ( .A1(n11971), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n10366) );
  NAND2_X1 U12786 ( .A1(n9628), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n10365) );
  INV_X1 U12787 ( .A(n10361), .ZN(n10359) );
  NAND2_X1 U12788 ( .A1(n10361), .A2(n10360), .ZN(n10362) );
  AND2_X1 U12789 ( .A1(n10724), .A2(n10362), .ZN(n10824) );
  NAND2_X1 U12790 ( .A1(n7325), .A2(n10824), .ZN(n10364) );
  NAND2_X1 U12791 ( .A1(n9624), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n10363) );
  NAND4_X1 U12792 ( .A1(n10366), .A2(n10365), .A3(n10364), .A4(n10363), .ZN(
        n13053) );
  NAND2_X1 U12793 ( .A1(n13053), .A2(n12987), .ZN(n10367) );
  NAND2_X1 U12794 ( .A1(n10368), .A2(n10367), .ZN(n10778) );
  NOR2_X1 U12795 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10126), .ZN(n13128) );
  AOI21_X1 U12796 ( .B1(n13040), .B2(n10778), .A(n13128), .ZN(n10369) );
  OAI21_X1 U12797 ( .B1(n13038), .B2(n10370), .A(n10369), .ZN(n10371) );
  AOI21_X1 U12798 ( .B1(n13491), .B2(n13026), .A(n10371), .ZN(n10372) );
  OAI21_X1 U12799 ( .B1(n10373), .B2(n13018), .A(n10372), .ZN(P2_U3208) );
  INV_X1 U12800 ( .A(n10530), .ZN(n10382) );
  NAND2_X1 U12801 ( .A1(n10520), .A2(n10374), .ZN(n10487) );
  INV_X1 U12802 ( .A(n10487), .ZN(n10375) );
  NOR2_X1 U12803 ( .A1(n6601), .A2(n10375), .ZN(n10377) );
  XNOR2_X1 U12804 ( .A(n10531), .B(n11664), .ZN(n10483) );
  XNOR2_X1 U12805 ( .A(n10485), .B(n10483), .ZN(n10376) );
  NAND2_X1 U12806 ( .A1(n10377), .A2(n10376), .ZN(n10445) );
  OAI211_X1 U12807 ( .C1(n10377), .C2(n10376), .A(n10445), .B(n12346), .ZN(
        n10380) );
  NOR2_X1 U12808 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n6614), .ZN(n14821) );
  OAI22_X1 U12809 ( .A1(n10789), .A2(n12341), .B1(n10520), .B2(n12361), .ZN(
        n10378) );
  AOI211_X1 U12810 ( .C1(n12364), .C2(n10531), .A(n14821), .B(n10378), .ZN(
        n10379) );
  OAI211_X1 U12811 ( .C1(n10382), .C2(n10381), .A(n10380), .B(n10379), .ZN(
        P3_U3179) );
  NAND2_X1 U12812 ( .A1(n12385), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n10383) );
  OAI21_X1 U12813 ( .B1(n12568), .B2(n12385), .A(n10383), .ZN(P3_U3520) );
  NAND2_X1 U12814 ( .A1(n12385), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n10384) );
  OAI21_X1 U12815 ( .B1(n12553), .B2(n12385), .A(n10384), .ZN(P3_U3521) );
  NAND2_X1 U12816 ( .A1(n13627), .A2(n10392), .ZN(n10385) );
  NAND2_X1 U12817 ( .A1(n10570), .A2(n10573), .ZN(n10569) );
  OR2_X1 U12818 ( .A1(n14459), .A2(n13672), .ZN(n10387) );
  NAND2_X1 U12819 ( .A1(n10569), .A2(n10387), .ZN(n10388) );
  NAND2_X1 U12820 ( .A1(n10388), .A2(n10625), .ZN(n10633) );
  OAI21_X1 U12821 ( .B1(n10388), .B2(n10625), .A(n10633), .ZN(n10940) );
  INV_X1 U12822 ( .A(n10940), .ZN(n10401) );
  INV_X1 U12823 ( .A(n10389), .ZN(n10390) );
  NAND2_X1 U12824 ( .A1(n10596), .A2(n10392), .ZN(n10393) );
  NAND2_X1 U12825 ( .A1(n10394), .A2(n10393), .ZN(n10574) );
  INV_X1 U12826 ( .A(n10574), .ZN(n10395) );
  INV_X1 U12827 ( .A(n13672), .ZN(n11023) );
  OR2_X1 U12828 ( .A1(n14459), .A2(n11023), .ZN(n10396) );
  NAND2_X1 U12829 ( .A1(n10397), .A2(n10396), .ZN(n10628) );
  XNOR2_X1 U12830 ( .A(n10628), .B(n10625), .ZN(n10398) );
  NAND2_X1 U12831 ( .A1(n10398), .A2(n14529), .ZN(n10400) );
  AOI22_X1 U12832 ( .A1(n13954), .A2(n13672), .B1(n13670), .B2(n13955), .ZN(
        n10399) );
  AND2_X1 U12833 ( .A1(n10400), .A2(n10399), .ZN(n10935) );
  INV_X1 U12834 ( .A(n11027), .ZN(n10934) );
  OAI211_X1 U12835 ( .C1(n10571), .C2(n10934), .A(n14490), .B(n10952), .ZN(
        n10936) );
  OAI211_X1 U12836 ( .C1(n10401), .C2(n14405), .A(n10935), .B(n10936), .ZN(
        n10594) );
  OAI22_X1 U12837 ( .A1(n14084), .A2(n10934), .B1(n14540), .B2(n9469), .ZN(
        n10402) );
  AOI21_X1 U12838 ( .B1(n10594), .B2(n14540), .A(n10402), .ZN(n10403) );
  INV_X1 U12839 ( .A(n10403), .ZN(P1_U3536) );
  NOR2_X1 U12840 ( .A1(n10405), .A2(n10404), .ZN(n10407) );
  NOR2_X1 U12841 ( .A1(n10407), .A2(n10406), .ZN(n10409) );
  XNOR2_X1 U12842 ( .A(n11348), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n10408) );
  NOR2_X1 U12843 ( .A1(n10409), .A2(n10408), .ZN(n11031) );
  AOI211_X1 U12844 ( .C1(n10409), .C2(n10408), .A(n11031), .B(n14604), .ZN(
        n10420) );
  NAND2_X1 U12845 ( .A1(n11287), .A2(n10410), .ZN(n10412) );
  NAND2_X1 U12846 ( .A1(n10412), .A2(n10411), .ZN(n10415) );
  NOR2_X1 U12847 ( .A1(n11348), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n10413) );
  AOI21_X1 U12848 ( .B1(n11348), .B2(P2_REG2_REG_16__SCAN_IN), .A(n10413), 
        .ZN(n10414) );
  NAND2_X1 U12849 ( .A1(n10414), .A2(n10415), .ZN(n11037) );
  OAI211_X1 U12850 ( .C1(n10415), .C2(n10414), .A(n14579), .B(n11037), .ZN(
        n10418) );
  NAND2_X1 U12851 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n11507)
         );
  INV_X1 U12852 ( .A(n11507), .ZN(n10416) );
  AOI21_X1 U12853 ( .B1(n14610), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n10416), 
        .ZN(n10417) );
  OAI211_X1 U12854 ( .C1(n14618), .C2(n11039), .A(n10418), .B(n10417), .ZN(
        n10419) );
  OR2_X1 U12855 ( .A1(n10420), .A2(n10419), .ZN(P2_U3230) );
  NAND2_X1 U12856 ( .A1(n10525), .A2(n10421), .ZN(n10799) );
  XNOR2_X1 U12857 ( .A(n10799), .B(n10673), .ZN(n10428) );
  NAND3_X1 U12858 ( .A1(n10422), .A2(n10673), .A3(n10423), .ZN(n10424) );
  NAND2_X1 U12859 ( .A1(n10425), .A2(n10424), .ZN(n14973) );
  OAI22_X1 U12860 ( .A1(n10485), .A2(n14919), .B1(n10804), .B2(n14917), .ZN(
        n10426) );
  AOI21_X1 U12861 ( .B1(n14973), .B2(n12804), .A(n10426), .ZN(n10427) );
  OAI21_X1 U12862 ( .B1(n10428), .B2(n14303), .A(n10427), .ZN(n14971) );
  INV_X1 U12863 ( .A(n14971), .ZN(n10433) );
  INV_X1 U12864 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n14831) );
  NOR2_X1 U12865 ( .A1(n10429), .A2(n14979), .ZN(n14972) );
  AOI22_X1 U12866 ( .A1(n14972), .A2(n14310), .B1(n14938), .B2(n10448), .ZN(
        n10430) );
  OAI21_X1 U12867 ( .B1(n14831), .B2(n14942), .A(n10430), .ZN(n10431) );
  AOI21_X1 U12868 ( .B1(n14973), .B2(n14939), .A(n10431), .ZN(n10432) );
  OAI21_X1 U12869 ( .B1(n10433), .B2(n14944), .A(n10432), .ZN(P3_U3226) );
  INV_X1 U12870 ( .A(n10434), .ZN(n10435) );
  NOR2_X1 U12871 ( .A1(n12177), .A2(n10435), .ZN(n10436) );
  NOR2_X1 U12872 ( .A1(n14268), .A2(n12154), .ZN(n10443) );
  INV_X2 U12873 ( .A(n13966), .ZN(n13941) );
  INV_X1 U12874 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10437) );
  OAI22_X1 U12875 ( .A1(n13941), .A2(n10438), .B1(n10437), .B2(n14483), .ZN(
        n10441) );
  INV_X1 U12876 ( .A(n13989), .ZN(n14270) );
  AOI21_X1 U12877 ( .B1(n14270), .B2(n13978), .A(n10439), .ZN(n10440) );
  AOI211_X1 U12878 ( .C1(n14498), .C2(P1_REG2_REG_0__SCAN_IN), .A(n10441), .B(
        n10440), .ZN(n10442) );
  OAI21_X1 U12879 ( .B1(n10444), .B2(n10443), .A(n10442), .ZN(P1_U3293) );
  NAND2_X1 U12880 ( .A1(n12380), .A2(n10483), .ZN(n10488) );
  NAND2_X1 U12881 ( .A1(n10445), .A2(n10488), .ZN(n10784) );
  XNOR2_X1 U12882 ( .A(n10784), .B(n10783), .ZN(n10451) );
  INV_X1 U12883 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n15133) );
  NOR2_X1 U12884 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15133), .ZN(n14840) );
  OAI22_X1 U12885 ( .A1(n10485), .A2(n12361), .B1(n10804), .B2(n12341), .ZN(
        n10446) );
  AOI211_X1 U12886 ( .C1(n12364), .C2(n10447), .A(n14840), .B(n10446), .ZN(
        n10450) );
  NAND2_X1 U12887 ( .A1(n12358), .A2(n10448), .ZN(n10449) );
  OAI211_X1 U12888 ( .C1(n10451), .C2(n12366), .A(n10450), .B(n10449), .ZN(
        P3_U3153) );
  INV_X1 U12889 ( .A(n10452), .ZN(n10454) );
  OAI222_X1 U12890 ( .A1(n7977), .A2(P3_U3151), .B1(n12886), .B2(n10454), .C1(
        n10453), .C2(n12883), .ZN(P3_U3274) );
  XNOR2_X1 U12891 ( .A(n10455), .B(n10456), .ZN(n14506) );
  XNOR2_X1 U12892 ( .A(n10457), .B(n10456), .ZN(n10458) );
  NAND2_X1 U12893 ( .A1(n10458), .A2(n14529), .ZN(n10461) );
  INV_X1 U12894 ( .A(n10459), .ZN(n10460) );
  NAND2_X1 U12895 ( .A1(n10461), .A2(n10460), .ZN(n10462) );
  AOI21_X1 U12896 ( .B1(n14506), .B2(n14482), .A(n10462), .ZN(n14508) );
  NAND2_X1 U12897 ( .A1(n14487), .A2(n10463), .ZN(n10468) );
  AOI21_X1 U12898 ( .B1(n10464), .B2(n10463), .A(n13961), .ZN(n10465) );
  NAND2_X1 U12899 ( .A1(n10465), .A2(n14488), .ZN(n14503) );
  INV_X1 U12900 ( .A(n14503), .ZN(n10466) );
  AOI22_X1 U12901 ( .A1(n14494), .A2(n10466), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n14466), .ZN(n10467) );
  OAI211_X1 U12902 ( .C1(n9213), .C2(n13966), .A(n10468), .B(n10467), .ZN(
        n10469) );
  AOI21_X1 U12903 ( .B1(n14495), .B2(n14506), .A(n10469), .ZN(n10470) );
  OAI21_X1 U12904 ( .B1(n14498), .B2(n14508), .A(n10470), .ZN(P1_U3291) );
  INV_X1 U12905 ( .A(n10471), .ZN(n10472) );
  AOI21_X1 U12906 ( .B1(n10474), .B2(n10473), .A(n10472), .ZN(n14468) );
  XOR2_X1 U12907 ( .A(n10475), .B(n10474), .Z(n10478) );
  NOR2_X1 U12908 ( .A1(n14468), .A2(n13855), .ZN(n10476) );
  AOI211_X1 U12909 ( .C1(n10478), .C2(n14529), .A(n10477), .B(n10476), .ZN(
        n14474) );
  OAI211_X1 U12910 ( .C1(n6826), .C2(n6954), .A(n14490), .B(n10479), .ZN(
        n14469) );
  OAI211_X1 U12911 ( .C1(n14468), .C2(n10480), .A(n14474), .B(n14469), .ZN(
        n10590) );
  OAI22_X1 U12912 ( .A1(n14084), .A2(n6954), .B1(n14540), .B2(n9208), .ZN(
        n10481) );
  AOI21_X1 U12913 ( .B1(n10590), .B2(n14540), .A(n10481), .ZN(n10482) );
  INV_X1 U12914 ( .A(n10482), .ZN(P1_U3533) );
  XNOR2_X1 U12915 ( .A(n10811), .B(n11698), .ZN(n10832) );
  XNOR2_X1 U12916 ( .A(n10832), .B(n10791), .ZN(n10497) );
  XNOR2_X1 U12917 ( .A(n10790), .B(n11664), .ZN(n10491) );
  XNOR2_X1 U12918 ( .A(n10804), .B(n10491), .ZN(n10490) );
  INV_X1 U12919 ( .A(n10490), .ZN(n10785) );
  INV_X1 U12920 ( .A(n10483), .ZN(n10484) );
  NAND2_X1 U12921 ( .A1(n10485), .A2(n10484), .ZN(n10486) );
  OAI21_X1 U12922 ( .B1(n10490), .B2(n10488), .A(n10783), .ZN(n10494) );
  INV_X1 U12923 ( .A(n10783), .ZN(n10489) );
  OAI21_X1 U12924 ( .B1(n10490), .B2(n10789), .A(n10489), .ZN(n10493) );
  INV_X1 U12925 ( .A(n10491), .ZN(n10492) );
  AOI22_X1 U12926 ( .A1(n10494), .A2(n10493), .B1(n10492), .B2(n12378), .ZN(
        n10495) );
  AOI21_X1 U12927 ( .B1(n10497), .B2(n10496), .A(n10838), .ZN(n10498) );
  NOR2_X1 U12928 ( .A1(n10498), .A2(n12366), .ZN(n10504) );
  AND2_X1 U12929 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n14878) );
  AOI21_X1 U12930 ( .B1(n12378), .B2(n12338), .A(n14878), .ZN(n10502) );
  NAND2_X1 U12931 ( .A1(n12364), .A2(n10811), .ZN(n10501) );
  NAND2_X1 U12932 ( .A1(n12358), .A2(n10808), .ZN(n10500) );
  NAND2_X1 U12933 ( .A1(n12357), .A2(n12376), .ZN(n10499) );
  NAND4_X1 U12934 ( .A1(n10502), .A2(n10501), .A3(n10500), .A4(n10499), .ZN(
        n10503) );
  OR2_X1 U12935 ( .A1(n10504), .A2(n10503), .ZN(P3_U3171) );
  INV_X1 U12936 ( .A(n10505), .ZN(n10510) );
  OAI22_X1 U12937 ( .A1(n13330), .A2(n9124), .B1(n10506), .B2(n14646), .ZN(
        n10509) );
  OAI22_X1 U12938 ( .A1(n13307), .A2(n10507), .B1(n11814), .B2(n14625), .ZN(
        n10508) );
  AOI211_X1 U12939 ( .C1(n13330), .C2(n10510), .A(n10509), .B(n10508), .ZN(
        n10511) );
  OAI21_X1 U12940 ( .B1(n13397), .B2(n10512), .A(n10511), .ZN(P2_U3263) );
  NAND2_X1 U12941 ( .A1(n10514), .A2(n10513), .ZN(n10516) );
  NAND2_X1 U12942 ( .A1(n10516), .A2(n10515), .ZN(n10517) );
  OR2_X1 U12943 ( .A1(n10517), .A2(n10522), .ZN(n10518) );
  NAND2_X1 U12944 ( .A1(n10422), .A2(n10518), .ZN(n10519) );
  INV_X1 U12945 ( .A(n10519), .ZN(n14968) );
  NAND2_X1 U12946 ( .A1(n10519), .A2(n12804), .ZN(n10528) );
  OAI22_X1 U12947 ( .A1(n10789), .A2(n14917), .B1(n10520), .B2(n14919), .ZN(
        n10521) );
  INV_X1 U12948 ( .A(n10521), .ZN(n10527) );
  NAND2_X1 U12949 ( .A1(n10523), .A2(n10522), .ZN(n10524) );
  NAND3_X1 U12950 ( .A1(n10525), .A2(n14922), .A3(n10524), .ZN(n10526) );
  NAND3_X1 U12951 ( .A1(n10528), .A2(n10527), .A3(n10526), .ZN(n14969) );
  MUX2_X1 U12952 ( .A(n14969), .B(P3_REG2_REG_6__SCAN_IN), .S(n14944), .Z(
        n10529) );
  INV_X1 U12953 ( .A(n10529), .ZN(n10533) );
  AOI22_X1 U12954 ( .A1(n12604), .A2(n10531), .B1(n14938), .B2(n10530), .ZN(
        n10532) );
  OAI211_X1 U12955 ( .C1(n14968), .C2(n12607), .A(n10533), .B(n10532), .ZN(
        P3_U3227) );
  INV_X1 U12956 ( .A(n10534), .ZN(n10537) );
  OAI22_X1 U12957 ( .A1(n10535), .A2(P3_U3151), .B1(SI_22_), .B2(n12870), .ZN(
        n10536) );
  AOI21_X1 U12958 ( .B1(n10537), .B2(n12875), .A(n10536), .ZN(P3_U3273) );
  NAND2_X1 U12959 ( .A1(n10538), .A2(n12034), .ZN(n10540) );
  NAND2_X1 U12960 ( .A1(n11848), .A2(n13056), .ZN(n10539) );
  XNOR2_X1 U12961 ( .A(n14720), .B(n13055), .ZN(n12036) );
  INV_X1 U12962 ( .A(n12036), .ZN(n10759) );
  XNOR2_X1 U12963 ( .A(n10760), .B(n10759), .ZN(n14719) );
  INV_X1 U12964 ( .A(n10544), .ZN(n10543) );
  AOI21_X1 U12965 ( .B1(n10543), .B2(n10759), .A(n14640), .ZN(n10546) );
  AOI21_X1 U12966 ( .B1(n10546), .B2(n10752), .A(n10545), .ZN(n14722) );
  INV_X1 U12967 ( .A(n14722), .ZN(n10553) );
  AOI21_X1 U12968 ( .B1(n10547), .B2(n14720), .A(n14633), .ZN(n10548) );
  NOR2_X2 U12969 ( .A1(n10547), .A2(n14720), .ZN(n10765) );
  INV_X1 U12970 ( .A(n10765), .ZN(n10774) );
  NAND2_X1 U12971 ( .A1(n10548), .A2(n10774), .ZN(n14721) );
  OAI22_X1 U12972 ( .A1(n13330), .A2(n9454), .B1(n10549), .B2(n14646), .ZN(
        n10550) );
  AOI21_X1 U12973 ( .B1(n14720), .B2(n13303), .A(n10550), .ZN(n10551) );
  OAI21_X1 U12974 ( .B1(n14721), .B2(n13307), .A(n10551), .ZN(n10552) );
  AOI21_X1 U12975 ( .B1(n10553), .B2(n13330), .A(n10552), .ZN(n10554) );
  OAI21_X1 U12976 ( .B1(n14719), .B2(n13397), .A(n10554), .ZN(P2_U3255) );
  NAND2_X1 U12977 ( .A1(n14532), .A2(n14522), .ZN(n14123) );
  INV_X1 U12978 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10555) );
  OAI22_X1 U12979 ( .A1(n14123), .A2(n13627), .B1(n14532), .B2(n10555), .ZN(
        n10556) );
  INV_X1 U12980 ( .A(n10556), .ZN(n10557) );
  OAI21_X1 U12981 ( .B1(n10558), .B2(n14530), .A(n10557), .ZN(P1_U3477) );
  INV_X1 U12982 ( .A(n10559), .ZN(n10568) );
  INV_X1 U12983 ( .A(n10560), .ZN(n10566) );
  OAI22_X1 U12984 ( .A1(n13330), .A2(n9187), .B1(n10561), .B2(n14646), .ZN(
        n10562) );
  AOI21_X1 U12985 ( .B1(n13303), .B2(n11848), .A(n10562), .ZN(n10563) );
  OAI21_X1 U12986 ( .B1(n10564), .B2(n13307), .A(n10563), .ZN(n10565) );
  AOI21_X1 U12987 ( .B1(n10566), .B2(n13330), .A(n10565), .ZN(n10567) );
  OAI21_X1 U12988 ( .B1(n10568), .B2(n13397), .A(n10567), .ZN(P2_U3256) );
  OAI21_X1 U12989 ( .B1(n10570), .B2(n10573), .A(n10569), .ZN(n14461) );
  AOI211_X1 U12990 ( .C1(n14459), .C2(n10572), .A(n13961), .B(n10571), .ZN(
        n14460) );
  XNOR2_X1 U12991 ( .A(n10574), .B(n10573), .ZN(n10575) );
  AOI22_X1 U12992 ( .A1(n13954), .A2(n13673), .B1(n13671), .B2(n13955), .ZN(
        n10608) );
  OAI21_X1 U12993 ( .B1(n10575), .B2(n14478), .A(n10608), .ZN(n10576) );
  AOI21_X1 U12994 ( .B1(n14461), .B2(n14482), .A(n10576), .ZN(n14464) );
  INV_X1 U12995 ( .A(n14464), .ZN(n10577) );
  AOI211_X1 U12996 ( .C1(n14517), .C2(n14461), .A(n14460), .B(n10577), .ZN(
        n10584) );
  INV_X1 U12997 ( .A(n14459), .ZN(n10581) );
  INV_X1 U12998 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10578) );
  OAI22_X1 U12999 ( .A1(n14123), .A2(n10581), .B1(n14532), .B2(n10578), .ZN(
        n10579) );
  INV_X1 U13000 ( .A(n10579), .ZN(n10580) );
  OAI21_X1 U13001 ( .B1(n10584), .B2(n14530), .A(n10580), .ZN(P1_U3480) );
  OAI22_X1 U13002 ( .A1(n14084), .A2(n10581), .B1(n14540), .B2(n9468), .ZN(
        n10582) );
  INV_X1 U13003 ( .A(n10582), .ZN(n10583) );
  OAI21_X1 U13004 ( .B1(n10584), .B2(n14537), .A(n10583), .ZN(P1_U3535) );
  INV_X1 U13005 ( .A(n11918), .ZN(n10587) );
  OAI222_X1 U13006 ( .A1(n13526), .A2(n10587), .B1(n12062), .B2(P2_U3088), 
        .C1(n10585), .C2(n13523), .ZN(P2_U3307) );
  OAI222_X1 U13007 ( .A1(n14135), .A2(n7736), .B1(n12134), .B2(n10587), .C1(
        n10586), .C2(P1_U3086), .ZN(P1_U3335) );
  INV_X1 U13008 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10588) );
  OAI22_X1 U13009 ( .A1(n14123), .A2(n6954), .B1(n14532), .B2(n10588), .ZN(
        n10589) );
  AOI21_X1 U13010 ( .B1(n10590), .B2(n14532), .A(n10589), .ZN(n10591) );
  INV_X1 U13011 ( .A(n10591), .ZN(P1_U3474) );
  INV_X1 U13012 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10592) );
  OAI22_X1 U13013 ( .A1(n14123), .A2(n10934), .B1(n14532), .B2(n10592), .ZN(
        n10593) );
  AOI21_X1 U13014 ( .B1(n10594), .B2(n14532), .A(n10593), .ZN(n10595) );
  INV_X1 U13015 ( .A(n10595), .ZN(P1_U3483) );
  AOI22_X1 U13016 ( .A1(n12247), .A2(n10596), .B1(n12259), .B2(n13673), .ZN(
        n10602) );
  NAND2_X1 U13017 ( .A1(n10596), .A2(n12255), .ZN(n10598) );
  NAND2_X1 U13018 ( .A1(n13673), .A2(n12247), .ZN(n10597) );
  NAND2_X1 U13019 ( .A1(n10598), .A2(n10597), .ZN(n10599) );
  XNOR2_X1 U13020 ( .A(n10599), .B(n10099), .ZN(n10601) );
  XNOR2_X1 U13021 ( .A(n10601), .B(n10602), .ZN(n13622) );
  NOR2_X1 U13022 ( .A1(n11023), .A2(n9810), .ZN(n10603) );
  AOI21_X1 U13023 ( .B1(n14459), .B2(n12247), .A(n10603), .ZN(n11016) );
  AOI22_X1 U13024 ( .A1(n14459), .A2(n12255), .B1(n12247), .B2(n13672), .ZN(
        n10604) );
  XNOR2_X1 U13025 ( .A(n10604), .B(n10099), .ZN(n11015) );
  XOR2_X1 U13026 ( .A(n11016), .B(n11015), .Z(n10605) );
  OAI211_X1 U13027 ( .C1(n10606), .C2(n10605), .A(n11020), .B(n14356), .ZN(
        n10611) );
  INV_X1 U13028 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n10607) );
  OAI22_X1 U13029 ( .A1(n13647), .A2(n10608), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10607), .ZN(n10609) );
  AOI21_X1 U13030 ( .B1(n14459), .B2(n14389), .A(n10609), .ZN(n10610) );
  OAI211_X1 U13031 ( .C1(n14394), .C2(n10612), .A(n10611), .B(n10610), .ZN(
        P1_U3213) );
  XOR2_X1 U13032 ( .A(n10613), .B(n10620), .Z(n14528) );
  INV_X1 U13033 ( .A(n14528), .ZN(n10624) );
  MUX2_X1 U13034 ( .A(n14520), .B(P1_REG2_REG_4__SCAN_IN), .S(n13941), .Z(
        n10619) );
  INV_X1 U13035 ( .A(n14494), .ZN(n13896) );
  OAI211_X1 U13036 ( .C1(n14489), .C2(n10615), .A(n14490), .B(n10614), .ZN(
        n14524) );
  INV_X1 U13037 ( .A(n10616), .ZN(n10617) );
  OAI22_X1 U13038 ( .A1(n13896), .A2(n14524), .B1(n10617), .B2(n14483), .ZN(
        n10618) );
  AOI211_X1 U13039 ( .C1(n14487), .C2(n14521), .A(n10619), .B(n10618), .ZN(
        n10623) );
  XOR2_X1 U13040 ( .A(n10621), .B(n10620), .Z(n14519) );
  NAND2_X1 U13041 ( .A1(n14519), .A2(n14268), .ZN(n10622) );
  OAI211_X1 U13042 ( .C1(n10624), .C2(n14274), .A(n10623), .B(n10622), .ZN(
        P1_U3289) );
  INV_X1 U13043 ( .A(n13670), .ZN(n11325) );
  INV_X1 U13044 ( .A(n10625), .ZN(n10627) );
  NOR2_X1 U13045 ( .A1(n11027), .A2(n11201), .ZN(n10626) );
  NAND2_X1 U13046 ( .A1(n11204), .A2(n11325), .ZN(n10629) );
  INV_X1 U13047 ( .A(n10635), .ZN(n10630) );
  OAI211_X1 U13048 ( .C1(n7327), .C2(n10630), .A(n14529), .B(n10982), .ZN(
        n10631) );
  OAI21_X1 U13049 ( .B1(n11325), .B2(n13982), .A(n10631), .ZN(n11007) );
  INV_X1 U13050 ( .A(n11007), .ZN(n10642) );
  OR2_X1 U13051 ( .A1(n11027), .A2(n13671), .ZN(n10632) );
  NAND2_X1 U13052 ( .A1(n10947), .A2(n6854), .ZN(n10946) );
  OR2_X1 U13053 ( .A1(n11204), .A2(n13670), .ZN(n10634) );
  NAND2_X1 U13054 ( .A1(n10946), .A2(n10634), .ZN(n10636) );
  NAND2_X1 U13055 ( .A1(n10636), .A2(n10635), .ZN(n10987) );
  OAI21_X1 U13056 ( .B1(n10636), .B2(n10635), .A(n10987), .ZN(n11009) );
  OR2_X2 U13057 ( .A1(n10952), .A2(n11204), .ZN(n10953) );
  AOI211_X1 U13058 ( .C1(n11327), .C2(n10953), .A(n13961), .B(n10989), .ZN(
        n10637) );
  AND2_X1 U13059 ( .A1(n13668), .A2(n13955), .ZN(n11321) );
  OR2_X1 U13060 ( .A1(n10637), .A2(n11321), .ZN(n11008) );
  NAND2_X1 U13061 ( .A1(n11008), .A2(n14494), .ZN(n10639) );
  AOI22_X1 U13062 ( .A1(n13941), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n11322), 
        .B2(n14466), .ZN(n10638) );
  OAI211_X1 U13063 ( .C1(n6833), .C2(n13978), .A(n10639), .B(n10638), .ZN(
        n10640) );
  AOI21_X1 U13064 ( .B1(n11009), .B2(n14268), .A(n10640), .ZN(n10641) );
  OAI21_X1 U13065 ( .B1(n10642), .B2(n14498), .A(n10641), .ZN(P1_U3283) );
  NAND2_X1 U13066 ( .A1(n10643), .A2(n9951), .ZN(n10646) );
  AOI22_X1 U13067 ( .A1(n12001), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n11898), 
        .B2(n10644), .ZN(n10645) );
  XNOR2_X1 U13068 ( .A(n11862), .B(n12911), .ZN(n10647) );
  NAND2_X1 U13069 ( .A1(n13053), .A2(n14633), .ZN(n10648) );
  NAND2_X1 U13070 ( .A1(n10647), .A2(n10648), .ZN(n10716) );
  INV_X1 U13071 ( .A(n10647), .ZN(n10650) );
  INV_X1 U13072 ( .A(n10648), .ZN(n10649) );
  NAND2_X1 U13073 ( .A1(n10650), .A2(n10649), .ZN(n10651) );
  NAND2_X1 U13074 ( .A1(n10716), .A2(n10651), .ZN(n10660) );
  INV_X1 U13075 ( .A(n10654), .ZN(n10655) );
  NAND2_X1 U13076 ( .A1(n10656), .A2(n10655), .ZN(n10657) );
  INV_X1 U13077 ( .A(n10717), .ZN(n10658) );
  AOI21_X1 U13078 ( .B1(n10660), .B2(n10659), .A(n10658), .ZN(n10672) );
  INV_X1 U13079 ( .A(n10824), .ZN(n10669) );
  NAND2_X1 U13080 ( .A1(n13054), .A2(n13004), .ZN(n10666) );
  NAND2_X1 U13081 ( .A1(n9624), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n10664) );
  NAND2_X1 U13082 ( .A1(n11971), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n10663) );
  XNOR2_X1 U13083 ( .A(n10724), .B(P2_REG3_REG_13__SCAN_IN), .ZN(n10766) );
  NAND2_X1 U13084 ( .A1(n7325), .A2(n10766), .ZN(n10662) );
  NAND2_X1 U13085 ( .A1(n9628), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n10661) );
  NAND4_X1 U13086 ( .A1(n10664), .A2(n10663), .A3(n10662), .A4(n10661), .ZN(
        n13052) );
  NAND2_X1 U13087 ( .A1(n13052), .A2(n12987), .ZN(n10665) );
  NAND2_X1 U13088 ( .A1(n10666), .A2(n10665), .ZN(n10818) );
  AOI21_X1 U13089 ( .B1(n13040), .B2(n10818), .A(n10667), .ZN(n10668) );
  OAI21_X1 U13090 ( .B1(n13038), .B2(n10669), .A(n10668), .ZN(n10670) );
  AOI21_X1 U13091 ( .B1(n11862), .B2(n13026), .A(n10670), .ZN(n10671) );
  OAI21_X1 U13092 ( .B1(n10672), .B2(n13018), .A(n10671), .ZN(P2_U3196) );
  NAND2_X1 U13093 ( .A1(n10799), .A2(n10673), .ZN(n10675) );
  NAND2_X1 U13094 ( .A1(n10675), .A2(n10674), .ZN(n10676) );
  XOR2_X1 U13095 ( .A(n10678), .B(n10676), .Z(n10681) );
  AOI22_X1 U13096 ( .A1(n14286), .A2(n12379), .B1(n12377), .B2(n14284), .ZN(
        n10680) );
  XNOR2_X1 U13097 ( .A(n10677), .B(n10678), .ZN(n14977) );
  NAND2_X1 U13098 ( .A1(n14977), .A2(n12804), .ZN(n10679) );
  OAI211_X1 U13099 ( .C1(n10681), .C2(n14303), .A(n10680), .B(n10679), .ZN(
        n14975) );
  INV_X1 U13100 ( .A(n14975), .ZN(n10685) );
  INV_X1 U13101 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n10907) );
  NOR2_X1 U13102 ( .A1(n10790), .A2(n14979), .ZN(n14976) );
  AOI22_X1 U13103 ( .A1(n14310), .A2(n14976), .B1(n14938), .B2(n10794), .ZN(
        n10682) );
  OAI21_X1 U13104 ( .B1(n10907), .B2(n14942), .A(n10682), .ZN(n10683) );
  AOI21_X1 U13105 ( .B1(n14977), .B2(n14939), .A(n10683), .ZN(n10684) );
  OAI21_X1 U13106 ( .B1(n10685), .B2(n14944), .A(n10684), .ZN(P3_U3225) );
  INV_X1 U13107 ( .A(n10686), .ZN(n10687) );
  AOI21_X1 U13108 ( .B1(n12029), .B2(n10688), .A(n10687), .ZN(n14704) );
  INV_X1 U13109 ( .A(n10689), .ZN(n10692) );
  INV_X1 U13110 ( .A(n10690), .ZN(n10691) );
  AOI211_X1 U13111 ( .C1(n14702), .C2(n10692), .A(n14633), .B(n10691), .ZN(
        n14701) );
  INV_X1 U13112 ( .A(n13024), .ZN(n10693) );
  OAI22_X1 U13113 ( .A1(n14625), .A2(n10694), .B1(n10693), .B2(n14646), .ZN(
        n10695) );
  AOI21_X1 U13114 ( .B1(n14701), .B2(n13395), .A(n10695), .ZN(n10701) );
  XNOR2_X1 U13115 ( .A(n10696), .B(n12029), .ZN(n10699) );
  NAND2_X1 U13116 ( .A1(n13060), .A2(n13004), .ZN(n10698) );
  NAND2_X1 U13117 ( .A1(n13058), .A2(n12987), .ZN(n10697) );
  NAND2_X1 U13118 ( .A1(n10698), .A2(n10697), .ZN(n13023) );
  AOI21_X1 U13119 ( .B1(n10699), .B2(n13391), .A(n13023), .ZN(n14700) );
  MUX2_X1 U13120 ( .A(n13113), .B(n14700), .S(n13330), .Z(n10700) );
  OAI211_X1 U13121 ( .C1(n14704), .C2(n13397), .A(n10701), .B(n10700), .ZN(
        P2_U3259) );
  INV_X1 U13122 ( .A(n10702), .ZN(n10703) );
  AOI21_X1 U13123 ( .B1(n12035), .B2(n10704), .A(n10703), .ZN(n14716) );
  INV_X1 U13124 ( .A(n14716), .ZN(n14713) );
  AOI211_X1 U13125 ( .C1(n14710), .C2(n10706), .A(n14633), .B(n10705), .ZN(
        n14709) );
  INV_X1 U13126 ( .A(n14710), .ZN(n10709) );
  AOI22_X1 U13127 ( .A1(n14653), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n10707), 
        .B2(n14621), .ZN(n10708) );
  OAI21_X1 U13128 ( .B1(n10709), .B2(n14625), .A(n10708), .ZN(n10710) );
  AOI21_X1 U13129 ( .B1(n14709), .B2(n13395), .A(n10710), .ZN(n10715) );
  XNOR2_X1 U13130 ( .A(n10711), .B(n12035), .ZN(n10713) );
  OAI21_X1 U13131 ( .B1(n10713), .B2(n14640), .A(n10712), .ZN(n14715) );
  NAND2_X1 U13132 ( .A1(n14715), .A2(n13330), .ZN(n10714) );
  OAI211_X1 U13133 ( .C1(n14713), .C2(n13397), .A(n10715), .B(n10714), .ZN(
        P2_U3257) );
  NAND2_X1 U13134 ( .A1(n10718), .A2(n9951), .ZN(n10721) );
  AOI22_X1 U13135 ( .A1(n12001), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n11898), 
        .B2(n10719), .ZN(n10720) );
  XNOR2_X1 U13136 ( .A(n11867), .B(n12911), .ZN(n11124) );
  NAND2_X1 U13137 ( .A1(n13052), .A2(n14633), .ZN(n11125) );
  XNOR2_X1 U13138 ( .A(n11124), .B(n11125), .ZN(n11123) );
  XNOR2_X1 U13139 ( .A(n11122), .B(n11123), .ZN(n10736) );
  NAND2_X1 U13140 ( .A1(n11971), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n10729) );
  NAND2_X1 U13141 ( .A1(n9624), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n10728) );
  INV_X1 U13142 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10722) );
  OAI21_X1 U13143 ( .B1(n10724), .B2(n10732), .A(n10722), .ZN(n10725) );
  NAND2_X1 U13144 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_REG3_REG_14__SCAN_IN), 
        .ZN(n10723) );
  AND2_X1 U13145 ( .A1(n10725), .A2(n11132), .ZN(n11164) );
  NAND2_X1 U13146 ( .A1(n7325), .A2(n11164), .ZN(n10727) );
  NAND2_X1 U13147 ( .A1(n9628), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n10726) );
  NAND4_X1 U13148 ( .A1(n10729), .A2(n10728), .A3(n10727), .A4(n10726), .ZN(
        n13051) );
  NAND2_X1 U13149 ( .A1(n13051), .A2(n12987), .ZN(n10731) );
  NAND2_X1 U13150 ( .A1(n13053), .A2(n13004), .ZN(n10730) );
  AND2_X1 U13151 ( .A1(n10731), .A2(n10730), .ZN(n10757) );
  OAI22_X1 U13152 ( .A1(n13015), .A2(n10757), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10732), .ZN(n10734) );
  INV_X1 U13153 ( .A(n11867), .ZN(n11055) );
  NOR2_X1 U13154 ( .A1(n11055), .A2(n13043), .ZN(n10733) );
  AOI211_X1 U13155 ( .C1(n13025), .C2(n10766), .A(n10734), .B(n10733), .ZN(
        n10735) );
  OAI21_X1 U13156 ( .B1(n10736), .B2(n13018), .A(n10735), .ZN(P2_U3206) );
  XNOR2_X1 U13157 ( .A(n10737), .B(n10742), .ZN(n14986) );
  AOI22_X1 U13158 ( .A1(n14286), .A2(n12377), .B1(n12375), .B2(n14284), .ZN(
        n10745) );
  NAND2_X1 U13159 ( .A1(n10799), .A2(n10738), .ZN(n10740) );
  NAND2_X1 U13160 ( .A1(n10740), .A2(n10739), .ZN(n10743) );
  OAI211_X1 U13161 ( .C1(n10743), .C2(n10742), .A(n10741), .B(n14922), .ZN(
        n10744) );
  OAI211_X1 U13162 ( .C1(n14986), .C2(n14925), .A(n10745), .B(n10744), .ZN(
        n14987) );
  NAND2_X1 U13163 ( .A1(n14987), .A2(n14942), .ZN(n10749) );
  NOR2_X1 U13164 ( .A1(n10831), .A2(n14979), .ZN(n14988) );
  INV_X1 U13165 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n10918) );
  INV_X1 U13166 ( .A(n10841), .ZN(n10746) );
  OAI22_X1 U13167 ( .A1(n14942), .A2(n10918), .B1(n10746), .B2(n14292), .ZN(
        n10747) );
  AOI21_X1 U13168 ( .B1(n14310), .B2(n14988), .A(n10747), .ZN(n10748) );
  OAI211_X1 U13169 ( .C1(n14986), .C2(n12607), .A(n10749), .B(n10748), .ZN(
        P3_U3223) );
  INV_X1 U13170 ( .A(n13055), .ZN(n10750) );
  OR2_X1 U13171 ( .A1(n14720), .A2(n10750), .ZN(n10751) );
  INV_X1 U13172 ( .A(n13054), .ZN(n10754) );
  XNOR2_X1 U13173 ( .A(n13491), .B(n10754), .ZN(n12040) );
  INV_X1 U13174 ( .A(n13053), .ZN(n10755) );
  AND2_X1 U13175 ( .A1(n11862), .A2(n10755), .ZN(n10756) );
  INV_X1 U13176 ( .A(n13052), .ZN(n11156) );
  XNOR2_X1 U13177 ( .A(n11867), .B(n11156), .ZN(n12041) );
  XNOR2_X1 U13178 ( .A(n11155), .B(n11154), .ZN(n10758) );
  OAI21_X1 U13179 ( .B1(n10758), .B2(n14640), .A(n10757), .ZN(n11056) );
  INV_X1 U13180 ( .A(n11056), .ZN(n10771) );
  INV_X2 U13181 ( .A(n13330), .ZN(n14653) );
  NAND2_X1 U13182 ( .A1(n10760), .A2(n10759), .ZN(n10762) );
  NAND2_X1 U13183 ( .A1(n14720), .A2(n13055), .ZN(n10761) );
  NAND2_X1 U13184 ( .A1(n10762), .A2(n10761), .ZN(n10772) );
  NAND2_X1 U13185 ( .A1(n13491), .A2(n13054), .ZN(n10763) );
  OR2_X1 U13186 ( .A1(n11862), .A2(n13053), .ZN(n10815) );
  NAND2_X1 U13187 ( .A1(n11862), .A2(n13053), .ZN(n10814) );
  XNOR2_X1 U13188 ( .A(n11149), .B(n11154), .ZN(n11058) );
  INV_X1 U13189 ( .A(n13397), .ZN(n14628) );
  OAI211_X1 U13190 ( .C1(n11055), .C2(n10821), .A(n13300), .B(n11163), .ZN(
        n11054) );
  AOI22_X1 U13191 ( .A1(n14653), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n10766), 
        .B2(n14621), .ZN(n10768) );
  NAND2_X1 U13192 ( .A1(n11867), .A2(n13303), .ZN(n10767) );
  OAI211_X1 U13193 ( .C1(n11054), .C2(n13307), .A(n10768), .B(n10767), .ZN(
        n10769) );
  AOI21_X1 U13194 ( .B1(n11058), .B2(n14628), .A(n10769), .ZN(n10770) );
  OAI21_X1 U13195 ( .B1(n10771), .B2(n14653), .A(n10770), .ZN(P2_U3252) );
  XNOR2_X1 U13196 ( .A(n10772), .B(n12040), .ZN(n13494) );
  INV_X1 U13197 ( .A(n10773), .ZN(n10823) );
  AOI211_X1 U13198 ( .C1(n13491), .C2(n10774), .A(n9633), .B(n10823), .ZN(
        n13490) );
  AOI22_X1 U13199 ( .A1(n14653), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n10775), 
        .B2(n14621), .ZN(n10776) );
  OAI21_X1 U13200 ( .B1(n10764), .B2(n14625), .A(n10776), .ZN(n10781) );
  OAI21_X1 U13201 ( .B1(n6607), .B2(n10753), .A(n10777), .ZN(n10779) );
  AOI21_X1 U13202 ( .B1(n10779), .B2(n13391), .A(n10778), .ZN(n13493) );
  NOR2_X1 U13203 ( .A1(n13493), .A2(n14653), .ZN(n10780) );
  AOI211_X1 U13204 ( .C1(n13490), .C2(n13395), .A(n10781), .B(n10780), .ZN(
        n10782) );
  OAI21_X1 U13205 ( .B1(n13397), .B2(n13494), .A(n10782), .ZN(P2_U3254) );
  MUX2_X1 U13206 ( .A(n12379), .B(n10784), .S(n10783), .Z(n10786) );
  XNOR2_X1 U13207 ( .A(n10786), .B(n10785), .ZN(n10796) );
  INV_X1 U13208 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n10787) );
  NOR2_X1 U13209 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10787), .ZN(n14857) );
  INV_X1 U13210 ( .A(n14857), .ZN(n10788) );
  OAI21_X1 U13211 ( .B1(n10789), .B2(n12361), .A(n10788), .ZN(n10793) );
  OAI22_X1 U13212 ( .A1(n10791), .A2(n12341), .B1(n12354), .B2(n10790), .ZN(
        n10792) );
  AOI211_X1 U13213 ( .C1(n10794), .C2(n12358), .A(n10793), .B(n10792), .ZN(
        n10795) );
  OAI21_X1 U13214 ( .B1(n10796), .B2(n12366), .A(n10795), .ZN(P3_U3161) );
  XOR2_X1 U13215 ( .A(n10797), .B(n10802), .Z(n14982) );
  NAND2_X1 U13216 ( .A1(n10799), .A2(n10798), .ZN(n10801) );
  NAND2_X1 U13217 ( .A1(n10801), .A2(n10800), .ZN(n10803) );
  XNOR2_X1 U13218 ( .A(n10803), .B(n10802), .ZN(n10806) );
  OAI22_X1 U13219 ( .A1(n14305), .A2(n14917), .B1(n10804), .B2(n14919), .ZN(
        n10805) );
  AOI21_X1 U13220 ( .B1(n10806), .B2(n14922), .A(n10805), .ZN(n10807) );
  OAI21_X1 U13221 ( .B1(n14982), .B2(n14925), .A(n10807), .ZN(n14984) );
  NAND2_X1 U13222 ( .A1(n14984), .A2(n14942), .ZN(n10813) );
  INV_X1 U13223 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n14867) );
  INV_X1 U13224 ( .A(n10808), .ZN(n10809) );
  OAI22_X1 U13225 ( .A1(n14942), .A2(n14867), .B1(n10809), .B2(n14292), .ZN(
        n10810) );
  AOI21_X1 U13226 ( .B1(n12604), .B2(n10811), .A(n10810), .ZN(n10812) );
  OAI211_X1 U13227 ( .C1(n14982), .C2(n12607), .A(n10813), .B(n10812), .ZN(
        P3_U3224) );
  NAND2_X1 U13228 ( .A1(n10815), .A2(n10814), .ZN(n12038) );
  XOR2_X1 U13229 ( .A(n10816), .B(n12038), .Z(n14331) );
  XNOR2_X1 U13230 ( .A(n10817), .B(n12038), .ZN(n10819) );
  AOI21_X1 U13231 ( .B1(n10819), .B2(n13391), .A(n10818), .ZN(n10820) );
  OAI21_X1 U13232 ( .B1(n14331), .B2(n14693), .A(n10820), .ZN(n14334) );
  NAND2_X1 U13233 ( .A1(n14334), .A2(n13330), .ZN(n10829) );
  INV_X1 U13234 ( .A(n11862), .ZN(n14333) );
  INV_X1 U13235 ( .A(n10821), .ZN(n10822) );
  OAI211_X1 U13236 ( .C1(n14333), .C2(n10823), .A(n10822), .B(n13300), .ZN(
        n14332) );
  INV_X1 U13237 ( .A(n14332), .ZN(n10827) );
  AOI22_X1 U13238 ( .A1(n14653), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n10824), 
        .B2(n14621), .ZN(n10825) );
  OAI21_X1 U13239 ( .B1(n14333), .B2(n14625), .A(n10825), .ZN(n10826) );
  AOI21_X1 U13240 ( .B1(n10827), .B2(n13395), .A(n10826), .ZN(n10828) );
  OAI211_X1 U13241 ( .C1(n14331), .C2(n10830), .A(n10829), .B(n10828), .ZN(
        P2_U3253) );
  XNOR2_X1 U13242 ( .A(n10831), .B(n11698), .ZN(n11063) );
  XNOR2_X1 U13243 ( .A(n11063), .B(n12376), .ZN(n10840) );
  INV_X1 U13244 ( .A(n10832), .ZN(n10833) );
  NOR2_X1 U13245 ( .A1(n12377), .A2(n10833), .ZN(n10834) );
  OR2_X1 U13246 ( .A1(n10838), .A2(n10834), .ZN(n10839) );
  INV_X1 U13247 ( .A(n10840), .ZN(n10836) );
  NAND2_X1 U13248 ( .A1(n10836), .A2(n10835), .ZN(n10837) );
  AOI211_X1 U13249 ( .C1(n10840), .C2(n10839), .A(n12366), .B(n11062), .ZN(
        n10848) );
  INV_X1 U13250 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n15052) );
  NOR2_X1 U13251 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15052), .ZN(n14889) );
  AOI21_X1 U13252 ( .B1(n12377), .B2(n12338), .A(n14889), .ZN(n10846) );
  NAND2_X1 U13253 ( .A1(n12358), .A2(n10841), .ZN(n10845) );
  NAND2_X1 U13254 ( .A1(n10842), .A2(n12364), .ZN(n10844) );
  OR2_X1 U13255 ( .A1(n10998), .A2(n12341), .ZN(n10843) );
  NAND4_X1 U13256 ( .A1(n10846), .A2(n10845), .A3(n10844), .A4(n10843), .ZN(
        n10847) );
  OR2_X1 U13257 ( .A1(n10848), .A2(n10847), .ZN(P3_U3157) );
  INV_X1 U13258 ( .A(n11934), .ZN(n11634) );
  OAI222_X1 U13259 ( .A1(n14135), .A2(n10850), .B1(n12134), .B2(n11634), .C1(
        P1_U3086), .C2(n10849), .ZN(P1_U3334) );
  INV_X1 U13260 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n14312) );
  INV_X1 U13261 ( .A(n14875), .ZN(n10914) );
  INV_X1 U13262 ( .A(n14838), .ZN(n10903) );
  INV_X1 U13263 ( .A(n14802), .ZN(n10893) );
  NOR2_X1 U13264 ( .A1(n14759), .A2(n10854), .ZN(n14777) );
  INV_X1 U13265 ( .A(n14783), .ZN(n10887) );
  AOI22_X1 U13266 ( .A1(n10887), .A2(P3_REG2_REG_4__SCAN_IN), .B1(n10886), 
        .B2(n14783), .ZN(n14776) );
  NOR2_X1 U13267 ( .A1(n10893), .A2(n10855), .ZN(n10856) );
  INV_X1 U13268 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n10857) );
  AOI22_X1 U13269 ( .A1(n10897), .A2(P3_REG2_REG_6__SCAN_IN), .B1(n10857), 
        .B2(n14819), .ZN(n14812) );
  NOR2_X1 U13270 ( .A1(n10903), .A2(n10858), .ZN(n10859) );
  AOI22_X1 U13271 ( .A1(n10908), .A2(P3_REG2_REG_8__SCAN_IN), .B1(n10907), 
        .B2(n14855), .ZN(n14848) );
  NOR2_X1 U13272 ( .A1(n10914), .A2(n10860), .ZN(n10861) );
  NAND2_X1 U13273 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n10920), .ZN(n10862) );
  OAI21_X1 U13274 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n10920), .A(n10862), 
        .ZN(n14899) );
  NOR2_X1 U13275 ( .A1(n14900), .A2(n14899), .ZN(n14898) );
  AOI21_X1 U13276 ( .B1(n14312), .B2(n10865), .A(n11073), .ZN(n10932) );
  NAND2_X1 U13277 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n10920), .ZN(n10876) );
  INV_X1 U13278 ( .A(n10920), .ZN(n14905) );
  INV_X1 U13279 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n15005) );
  AOI22_X1 U13280 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n10920), .B1(n14905), 
        .B2(n15005), .ZN(n14888) );
  INV_X1 U13281 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15002) );
  AOI22_X1 U13282 ( .A1(n10908), .A2(n15002), .B1(P3_REG1_REG_8__SCAN_IN), 
        .B2(n14855), .ZN(n14859) );
  INV_X1 U13283 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n14999) );
  AOI22_X1 U13284 ( .A1(n10897), .A2(n14999), .B1(P3_REG1_REG_6__SCAN_IN), 
        .B2(n14819), .ZN(n14823) );
  INV_X1 U13285 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n14996) );
  AOI22_X1 U13286 ( .A1(n10887), .A2(n14996), .B1(P3_REG1_REG_4__SCAN_IN), 
        .B2(n14783), .ZN(n14787) );
  OAI21_X1 U13287 ( .B1(n10867), .B2(n9781), .A(n10866), .ZN(n10868) );
  NAND2_X1 U13288 ( .A1(n10868), .A2(n14766), .ZN(n10869) );
  XNOR2_X1 U13289 ( .A(n10868), .B(n10882), .ZN(n14770) );
  NAND2_X1 U13290 ( .A1(P3_REG1_REG_3__SCAN_IN), .A2(n14770), .ZN(n14769) );
  NAND2_X1 U13291 ( .A1(n14802), .A2(n10870), .ZN(n10871) );
  NAND2_X1 U13292 ( .A1(P3_REG1_REG_5__SCAN_IN), .A2(n14806), .ZN(n14805) );
  NAND2_X1 U13293 ( .A1(n14838), .A2(n10872), .ZN(n10873) );
  NAND2_X1 U13294 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n14842), .ZN(n14841) );
  NAND2_X1 U13295 ( .A1(n14875), .A2(n10874), .ZN(n10875) );
  NAND2_X1 U13296 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n14881), .ZN(n14880) );
  NAND2_X1 U13297 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n10877), .ZN(n11078) );
  OAI21_X1 U13298 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n10877), .A(n11078), 
        .ZN(n10930) );
  AND2_X1 U13299 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n11066) );
  AOI21_X1 U13300 ( .B1(n14879), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n11066), 
        .ZN(n10878) );
  OAI21_X1 U13301 ( .B1(n14876), .B2(n11086), .A(n10878), .ZN(n10929) );
  INV_X1 U13302 ( .A(n10879), .ZN(n14761) );
  INV_X1 U13303 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10880) );
  MUX2_X1 U13304 ( .A(n10881), .B(n10880), .S(n6446), .Z(n10883) );
  NAND2_X1 U13305 ( .A1(n10883), .A2(n10882), .ZN(n14779) );
  INV_X1 U13306 ( .A(n10883), .ZN(n10884) );
  NAND2_X1 U13307 ( .A1(n10884), .A2(n14766), .ZN(n10885) );
  OAI21_X1 U13308 ( .B1(n14762), .B2(n14761), .A(n7324), .ZN(n14780) );
  MUX2_X1 U13309 ( .A(n10886), .B(n14996), .S(n6446), .Z(n10888) );
  NAND2_X1 U13310 ( .A1(n10888), .A2(n10887), .ZN(n10891) );
  INV_X1 U13311 ( .A(n10888), .ZN(n10889) );
  NAND2_X1 U13312 ( .A1(n10889), .A2(n14783), .ZN(n10890) );
  NAND2_X1 U13313 ( .A1(n10891), .A2(n10890), .ZN(n14778) );
  AOI21_X1 U13314 ( .B1(n14780), .B2(n14779), .A(n14778), .ZN(n14798) );
  INV_X1 U13315 ( .A(n10891), .ZN(n14797) );
  INV_X1 U13316 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n10892) );
  MUX2_X1 U13317 ( .A(n14795), .B(n10892), .S(n6446), .Z(n10894) );
  NAND2_X1 U13318 ( .A1(n10894), .A2(n10893), .ZN(n14815) );
  INV_X1 U13319 ( .A(n10894), .ZN(n10895) );
  NAND2_X1 U13320 ( .A1(n10895), .A2(n14802), .ZN(n10896) );
  AND2_X1 U13321 ( .A1(n14815), .A2(n10896), .ZN(n14796) );
  OAI21_X1 U13322 ( .B1(n14798), .B2(n14797), .A(n14796), .ZN(n14816) );
  MUX2_X1 U13323 ( .A(n10857), .B(n14999), .S(n6446), .Z(n10898) );
  NAND2_X1 U13324 ( .A1(n10898), .A2(n10897), .ZN(n10901) );
  INV_X1 U13325 ( .A(n10898), .ZN(n10899) );
  NAND2_X1 U13326 ( .A1(n10899), .A2(n14819), .ZN(n10900) );
  NAND2_X1 U13327 ( .A1(n10901), .A2(n10900), .ZN(n14814) );
  AOI21_X1 U13328 ( .B1(n14816), .B2(n14815), .A(n14814), .ZN(n14834) );
  INV_X1 U13329 ( .A(n10901), .ZN(n14833) );
  INV_X1 U13330 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n10902) );
  MUX2_X1 U13331 ( .A(n14831), .B(n10902), .S(n6446), .Z(n10904) );
  NAND2_X1 U13332 ( .A1(n10904), .A2(n10903), .ZN(n14851) );
  INV_X1 U13333 ( .A(n10904), .ZN(n10905) );
  NAND2_X1 U13334 ( .A1(n10905), .A2(n14838), .ZN(n10906) );
  AND2_X1 U13335 ( .A1(n14851), .A2(n10906), .ZN(n14832) );
  OAI21_X1 U13336 ( .B1(n14834), .B2(n14833), .A(n14832), .ZN(n14852) );
  MUX2_X1 U13337 ( .A(n10907), .B(n15002), .S(n6446), .Z(n10909) );
  NAND2_X1 U13338 ( .A1(n10909), .A2(n10908), .ZN(n10912) );
  INV_X1 U13339 ( .A(n10909), .ZN(n10910) );
  NAND2_X1 U13340 ( .A1(n10910), .A2(n14855), .ZN(n10911) );
  NAND2_X1 U13341 ( .A1(n10912), .A2(n10911), .ZN(n14850) );
  AOI21_X1 U13342 ( .B1(n14852), .B2(n14851), .A(n14850), .ZN(n14870) );
  INV_X1 U13343 ( .A(n10912), .ZN(n14869) );
  INV_X1 U13344 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n10913) );
  MUX2_X1 U13345 ( .A(n14867), .B(n10913), .S(n6446), .Z(n10915) );
  NAND2_X1 U13346 ( .A1(n10915), .A2(n10914), .ZN(n14893) );
  INV_X1 U13347 ( .A(n10915), .ZN(n10916) );
  NAND2_X1 U13348 ( .A1(n10916), .A2(n14875), .ZN(n10917) );
  AND2_X1 U13349 ( .A1(n14893), .A2(n10917), .ZN(n14868) );
  OAI21_X1 U13350 ( .B1(n14870), .B2(n14869), .A(n14868), .ZN(n14894) );
  MUX2_X1 U13351 ( .A(n10918), .B(n15005), .S(n6446), .Z(n10919) );
  NAND2_X1 U13352 ( .A1(n10919), .A2(n14905), .ZN(n10923) );
  INV_X1 U13353 ( .A(n10919), .ZN(n10921) );
  NAND2_X1 U13354 ( .A1(n10921), .A2(n10920), .ZN(n10922) );
  NAND2_X1 U13355 ( .A1(n10923), .A2(n10922), .ZN(n14892) );
  AOI21_X1 U13356 ( .B1(n14894), .B2(n14893), .A(n14892), .ZN(n14891) );
  INV_X1 U13357 ( .A(n10923), .ZN(n10924) );
  NOR2_X1 U13358 ( .A1(n14891), .A2(n10924), .ZN(n10926) );
  MUX2_X1 U13359 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n6446), .Z(n11087) );
  XNOR2_X1 U13360 ( .A(n11087), .B(n11086), .ZN(n10925) );
  AOI21_X1 U13361 ( .B1(n10926), .B2(n10925), .A(n11090), .ZN(n10927) );
  NOR2_X1 U13362 ( .A1(n10927), .A2(n14895), .ZN(n10928) );
  AOI211_X1 U13363 ( .C1(n6650), .C2(n10930), .A(n10929), .B(n10928), .ZN(
        n10931) );
  OAI21_X1 U13364 ( .B1(n10932), .B2(n14901), .A(n10931), .ZN(P3_U3193) );
  INV_X1 U13365 ( .A(n11026), .ZN(n10933) );
  OAI22_X1 U13366 ( .A1(n13978), .A2(n10934), .B1(n10933), .B2(n14483), .ZN(
        n10939) );
  OAI21_X1 U13367 ( .B1(n13878), .B2(n10936), .A(n10935), .ZN(n10937) );
  MUX2_X1 U13368 ( .A(n10937), .B(P1_REG2_REG_8__SCAN_IN), .S(n13941), .Z(
        n10938) );
  AOI211_X1 U13369 ( .C1(n14268), .C2(n10940), .A(n10939), .B(n10938), .ZN(
        n10941) );
  INV_X1 U13370 ( .A(n10941), .ZN(P1_U3285) );
  NAND2_X1 U13371 ( .A1(n10942), .A2(n12875), .ZN(n10944) );
  OAI211_X1 U13372 ( .C1(n10945), .C2(n12870), .A(n10944), .B(n10943), .ZN(
        P3_U3272) );
  OAI21_X1 U13373 ( .B1(n10947), .B2(n6854), .A(n10946), .ZN(n11045) );
  OAI21_X1 U13374 ( .B1(n10950), .B2(n10949), .A(n10948), .ZN(n10951) );
  AOI222_X1 U13375 ( .A1(n14529), .A2(n10951), .B1(n13669), .B2(n13955), .C1(
        n13671), .C2(n13954), .ZN(n11047) );
  INV_X1 U13376 ( .A(n11204), .ZN(n10957) );
  INV_X1 U13377 ( .A(n10952), .ZN(n10954) );
  OAI211_X1 U13378 ( .C1(n10957), .C2(n10954), .A(n10953), .B(n14490), .ZN(
        n10955) );
  NAND2_X1 U13379 ( .A1(n11047), .A2(n10955), .ZN(n11044) );
  AOI21_X1 U13380 ( .B1(n14518), .B2(n11045), .A(n11044), .ZN(n10961) );
  INV_X1 U13381 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10956) );
  OAI22_X1 U13382 ( .A1(n10957), .A2(n14123), .B1(n14532), .B2(n10956), .ZN(
        n10958) );
  INV_X1 U13383 ( .A(n10958), .ZN(n10959) );
  OAI21_X1 U13384 ( .B1(n10961), .B2(n14530), .A(n10959), .ZN(P1_U3486) );
  INV_X1 U13385 ( .A(n14084), .ZN(n11265) );
  AOI22_X1 U13386 ( .A1(n11265), .A2(n11204), .B1(n14537), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n10960) );
  OAI21_X1 U13387 ( .B1(n10961), .B2(n14537), .A(n10960), .ZN(P1_U3537) );
  INV_X1 U13388 ( .A(n10962), .ZN(n10963) );
  OAI21_X1 U13389 ( .B1(n11180), .B2(n10964), .A(n10963), .ZN(n10965) );
  NOR2_X1 U13390 ( .A1(n14447), .A2(n10965), .ZN(n10966) );
  XNOR2_X1 U13391 ( .A(n14447), .B(n10965), .ZN(n14441) );
  NOR2_X1 U13392 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14441), .ZN(n14440) );
  NOR2_X1 U13393 ( .A1(n10966), .A2(n14440), .ZN(n10969) );
  INV_X1 U13394 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n13728) );
  NOR2_X1 U13395 ( .A1(n13729), .A2(n13728), .ZN(n10967) );
  AOI21_X1 U13396 ( .B1(n13728), .B2(n13729), .A(n10967), .ZN(n10968) );
  NAND2_X1 U13397 ( .A1(n10968), .A2(n10969), .ZN(n13727) );
  OAI211_X1 U13398 ( .C1(n10969), .C2(n10968), .A(n13766), .B(n13727), .ZN(
        n10971) );
  INV_X1 U13399 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n15065) );
  NOR2_X1 U13400 ( .A1(n15065), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14361) );
  AOI21_X1 U13401 ( .B1(n13725), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n14361), 
        .ZN(n10970) );
  OAI211_X1 U13402 ( .C1(n13722), .C2(n13729), .A(n10971), .B(n10970), .ZN(
        n10981) );
  NAND2_X1 U13403 ( .A1(n10975), .A2(n10974), .ZN(n10976) );
  INV_X1 U13404 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14443) );
  NAND2_X1 U13405 ( .A1(n14444), .A2(n14443), .ZN(n14442) );
  NAND2_X1 U13406 ( .A1(n10976), .A2(n14442), .ZN(n10979) );
  INV_X1 U13407 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n14082) );
  NOR2_X1 U13408 ( .A1(n13733), .A2(n14082), .ZN(n10977) );
  AOI21_X1 U13409 ( .B1(n14082), .B2(n13733), .A(n10977), .ZN(n10978) );
  AOI211_X1 U13410 ( .C1(n10979), .C2(n10978), .A(n13732), .B(n13764), .ZN(
        n10980) );
  OR2_X1 U13411 ( .A1(n10981), .A2(n10980), .ZN(P1_U3259) );
  XNOR2_X1 U13412 ( .A(n11101), .B(n11099), .ZN(n10983) );
  NAND2_X1 U13413 ( .A1(n10983), .A2(n14529), .ZN(n10985) );
  AOI22_X1 U13414 ( .A1(n13667), .A2(n13955), .B1(n13954), .B2(n13669), .ZN(
        n10984) );
  NAND2_X1 U13415 ( .A1(n10985), .A2(n10984), .ZN(n14411) );
  INV_X1 U13416 ( .A(n14411), .ZN(n10995) );
  OR2_X1 U13417 ( .A1(n11327), .A2(n13669), .ZN(n10986) );
  NAND2_X1 U13418 ( .A1(n10987), .A2(n10986), .ZN(n10988) );
  NAND2_X1 U13419 ( .A1(n10988), .A2(n11099), .ZN(n11097) );
  OAI21_X1 U13420 ( .B1(n10988), .B2(n11099), .A(n11097), .ZN(n14413) );
  INV_X1 U13421 ( .A(n14390), .ZN(n14410) );
  OAI211_X1 U13422 ( .C1(n14410), .C2(n10989), .A(n6485), .B(n14490), .ZN(
        n14409) );
  AOI22_X1 U13423 ( .A1(n13941), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n10990), 
        .B2(n14466), .ZN(n10992) );
  NAND2_X1 U13424 ( .A1(n14390), .A2(n14487), .ZN(n10991) );
  OAI211_X1 U13425 ( .C1(n14409), .C2(n13896), .A(n10992), .B(n10991), .ZN(
        n10993) );
  AOI21_X1 U13426 ( .B1(n14413), .B2(n14268), .A(n10993), .ZN(n10994) );
  OAI21_X1 U13427 ( .B1(n14498), .B2(n10995), .A(n10994), .ZN(P1_U3282) );
  XNOR2_X1 U13428 ( .A(n10996), .B(n10999), .ZN(n10997) );
  OAI222_X1 U13429 ( .A1(n14917), .A2(n11420), .B1(n14919), .B2(n10998), .C1(
        n10997), .C2(n14303), .ZN(n14314) );
  INV_X1 U13430 ( .A(n14314), .ZN(n11006) );
  XNOR2_X1 U13431 ( .A(n11000), .B(n10999), .ZN(n14316) );
  OR2_X1 U13432 ( .A1(n12804), .A2(n14926), .ZN(n14307) );
  NAND2_X1 U13433 ( .A1(n14942), .A2(n14307), .ZN(n12727) );
  NOR2_X1 U13434 ( .A1(n11213), .A2(n14979), .ZN(n14315) );
  INV_X1 U13435 ( .A(n14315), .ZN(n11003) );
  AOI22_X1 U13436 ( .A1(n14944), .A2(P3_REG2_REG_12__SCAN_IN), .B1(n14938), 
        .B2(n11216), .ZN(n11001) );
  OAI21_X1 U13437 ( .B1(n11003), .B2(n11002), .A(n11001), .ZN(n11004) );
  AOI21_X1 U13438 ( .B1(n14316), .B2(n12739), .A(n11004), .ZN(n11005) );
  OAI21_X1 U13439 ( .B1(n11006), .B2(n14944), .A(n11005), .ZN(P3_U3221) );
  AOI211_X1 U13440 ( .C1(n14518), .C2(n11009), .A(n11008), .B(n11007), .ZN(
        n11013) );
  INV_X1 U13441 ( .A(n14123), .ZN(n11010) );
  AOI22_X1 U13442 ( .A1(n11327), .A2(n11010), .B1(n14530), .B2(
        P1_REG0_REG_10__SCAN_IN), .ZN(n11011) );
  OAI21_X1 U13443 ( .B1(n11013), .B2(n14530), .A(n11011), .ZN(P1_U3489) );
  AOI22_X1 U13444 ( .A1(n11327), .A2(n11265), .B1(n14537), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n11012) );
  OAI21_X1 U13445 ( .B1(n11013), .B2(n14537), .A(n11012), .ZN(P1_U3538) );
  AOI22_X1 U13446 ( .A1(n11027), .A2(n12255), .B1(n12247), .B2(n13671), .ZN(
        n11014) );
  XNOR2_X1 U13447 ( .A(n11014), .B(n10099), .ZN(n11192) );
  AOI22_X1 U13448 ( .A1(n11027), .A2(n12247), .B1(n12259), .B2(n13671), .ZN(
        n11193) );
  XNOR2_X1 U13449 ( .A(n11192), .B(n11193), .ZN(n11022) );
  INV_X1 U13450 ( .A(n11015), .ZN(n11018) );
  INV_X1 U13451 ( .A(n11016), .ZN(n11017) );
  AOI21_X1 U13452 ( .B1(n11022), .B2(n11021), .A(n6604), .ZN(n11030) );
  OAI22_X1 U13453 ( .A1(n11023), .A2(n14378), .B1(n14377), .B2(n11325), .ZN(
        n11024) );
  AOI211_X1 U13454 ( .C1(n13649), .C2(n11026), .A(n11025), .B(n11024), .ZN(
        n11029) );
  NAND2_X1 U13455 ( .A1(n14389), .A2(n11027), .ZN(n11028) );
  OAI211_X1 U13456 ( .C1(n11030), .C2(n14384), .A(n11029), .B(n11028), .ZN(
        P1_U3221) );
  NAND2_X1 U13457 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n11593)
         );
  INV_X1 U13458 ( .A(n11593), .ZN(n11035) );
  AOI21_X1 U13459 ( .B1(n11348), .B2(P2_REG1_REG_16__SCAN_IN), .A(n11031), 
        .ZN(n11033) );
  XNOR2_X1 U13460 ( .A(n13138), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n11032) );
  NOR2_X1 U13461 ( .A1(n11033), .A2(n11032), .ZN(n13137) );
  AOI211_X1 U13462 ( .C1(n11033), .C2(n11032), .A(n13137), .B(n14604), .ZN(
        n11034) );
  AOI211_X1 U13463 ( .C1(n14610), .C2(P2_ADDR_REG_17__SCAN_IN), .A(n11035), 
        .B(n11034), .ZN(n11043) );
  INV_X1 U13464 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13144) );
  NOR2_X1 U13465 ( .A1(n13145), .A2(n13144), .ZN(n11036) );
  AOI21_X1 U13466 ( .B1(n13144), .B2(n13145), .A(n11036), .ZN(n11041) );
  INV_X1 U13467 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n11038) );
  OAI21_X1 U13468 ( .B1(n11039), .B2(n11038), .A(n11037), .ZN(n11040) );
  NAND2_X1 U13469 ( .A1(n11041), .A2(n11040), .ZN(n13143) );
  OAI211_X1 U13470 ( .C1(n11041), .C2(n11040), .A(n14579), .B(n13143), .ZN(
        n11042) );
  OAI211_X1 U13471 ( .C1(n14618), .C2(n13145), .A(n11043), .B(n11042), .ZN(
        P2_U3231) );
  INV_X1 U13472 ( .A(n11045), .ZN(n11053) );
  AOI21_X1 U13473 ( .B1(n14482), .B2(n11045), .A(n11044), .ZN(n11046) );
  AOI211_X1 U13474 ( .C1(n13878), .C2(n11047), .A(n13941), .B(n11046), .ZN(
        n11048) );
  INV_X1 U13475 ( .A(n11048), .ZN(n11052) );
  INV_X1 U13476 ( .A(n11049), .ZN(n11200) );
  OAI22_X1 U13477 ( .A1(n13966), .A2(n9479), .B1(n11200), .B2(n14483), .ZN(
        n11050) );
  AOI21_X1 U13478 ( .B1(n14487), .B2(n11204), .A(n11050), .ZN(n11051) );
  OAI211_X1 U13479 ( .C1(n11053), .C2(n13865), .A(n11052), .B(n11051), .ZN(
        P1_U3284) );
  OAI21_X1 U13480 ( .B1(n11055), .B2(n14723), .A(n11054), .ZN(n11057) );
  AOI211_X1 U13481 ( .C1(n14680), .C2(n11058), .A(n11057), .B(n11056), .ZN(
        n11061) );
  NAND2_X1 U13482 ( .A1(n14729), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n11059) );
  OAI21_X1 U13483 ( .B1(n11061), .B2(n14729), .A(n11059), .ZN(P2_U3469) );
  NAND2_X1 U13484 ( .A1(n14744), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n11060) );
  OAI21_X1 U13485 ( .B1(n11061), .B2(n14744), .A(n11060), .ZN(P2_U3512) );
  NAND2_X1 U13486 ( .A1(n11063), .A2(n12376), .ZN(n11064) );
  XNOR2_X1 U13487 ( .A(n14308), .B(n11698), .ZN(n11208) );
  INV_X1 U13488 ( .A(n11208), .ZN(n11065) );
  XNOR2_X1 U13489 ( .A(n11207), .B(n12375), .ZN(n11071) );
  AOI21_X1 U13490 ( .B1(n12338), .B2(n12376), .A(n11066), .ZN(n11067) );
  OAI21_X1 U13491 ( .B1(n14306), .B2(n12341), .A(n11067), .ZN(n11069) );
  NOR2_X1 U13492 ( .A1(n14308), .A2(n12354), .ZN(n11068) );
  AOI211_X1 U13493 ( .C1(n14309), .C2(n12358), .A(n11069), .B(n11068), .ZN(
        n11070) );
  OAI21_X1 U13494 ( .B1(n11071), .B2(n12366), .A(n11070), .ZN(P3_U3176) );
  NOR2_X1 U13495 ( .A1(n10864), .A2(n11072), .ZN(n11074) );
  INV_X1 U13496 ( .A(n12387), .ZN(n12394) );
  INV_X1 U13497 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n15041) );
  AOI22_X1 U13498 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n12394), .B1(n12387), 
        .B2(n15041), .ZN(n11075) );
  AOI21_X1 U13499 ( .B1(n11076), .B2(n11075), .A(n12386), .ZN(n11095) );
  INV_X1 U13500 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14317) );
  AOI22_X1 U13501 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n12387), .B1(n12394), 
        .B2(n14317), .ZN(n11081) );
  NAND2_X1 U13502 ( .A1(n11086), .A2(n11077), .ZN(n11079) );
  OAI21_X1 U13503 ( .B1(n11081), .B2(n11080), .A(n12389), .ZN(n11085) );
  NOR2_X1 U13504 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11082), .ZN(n11211) );
  AOI21_X1 U13505 ( .B1(n14879), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n11211), 
        .ZN(n11083) );
  OAI21_X1 U13506 ( .B1(n14876), .B2(n12387), .A(n11083), .ZN(n11084) );
  AOI21_X1 U13507 ( .B1(n11085), .B2(n6650), .A(n11084), .ZN(n11094) );
  NOR2_X1 U13508 ( .A1(n11087), .A2(n11086), .ZN(n11089) );
  MUX2_X1 U13509 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n6446), .Z(n12393) );
  XNOR2_X1 U13510 ( .A(n12393), .B(n12387), .ZN(n11088) );
  NOR3_X1 U13511 ( .A1(n11090), .A2(n11089), .A3(n11088), .ZN(n12398) );
  INV_X1 U13512 ( .A(n12398), .ZN(n11092) );
  OAI21_X1 U13513 ( .B1(n11090), .B2(n11089), .A(n11088), .ZN(n11091) );
  NAND3_X1 U13514 ( .A1(n11092), .A2(n14871), .A3(n11091), .ZN(n11093) );
  OAI211_X1 U13515 ( .C1(n11095), .C2(n14901), .A(n11094), .B(n11093), .ZN(
        P3_U3194) );
  OR2_X1 U13516 ( .A1(n14390), .A2(n13668), .ZN(n11096) );
  NAND2_X1 U13517 ( .A1(n11097), .A2(n11096), .ZN(n11098) );
  NAND2_X1 U13518 ( .A1(n11098), .A2(n11104), .ZN(n11171) );
  OAI21_X1 U13519 ( .B1(n11098), .B2(n11104), .A(n11171), .ZN(n11261) );
  INV_X1 U13520 ( .A(n11261), .ZN(n11112) );
  INV_X1 U13521 ( .A(n11099), .ZN(n11100) );
  NAND2_X1 U13522 ( .A1(n11101), .A2(n11100), .ZN(n11103) );
  OR2_X1 U13523 ( .A1(n14390), .A2(n11532), .ZN(n11102) );
  NAND2_X1 U13524 ( .A1(n11103), .A2(n11102), .ZN(n11186) );
  INV_X1 U13525 ( .A(n11104), .ZN(n11185) );
  XNOR2_X1 U13526 ( .A(n11186), .B(n11185), .ZN(n11107) );
  NAND2_X1 U13527 ( .A1(n11261), .A2(n14482), .ZN(n11106) );
  AOI22_X1 U13528 ( .A1(n13954), .A2(n13668), .B1(n13666), .B2(n13955), .ZN(
        n11105) );
  OAI211_X1 U13529 ( .C1(n14478), .C2(n11107), .A(n11106), .B(n11105), .ZN(
        n11259) );
  NAND2_X1 U13530 ( .A1(n11259), .A2(n13966), .ZN(n11111) );
  AOI211_X1 U13531 ( .C1(n11266), .C2(n6485), .A(n13961), .B(n6830), .ZN(
        n11260) );
  AOI22_X1 U13532 ( .A1(n13941), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n11535), 
        .B2(n14466), .ZN(n11108) );
  OAI21_X1 U13533 ( .B1(n11538), .B2(n13978), .A(n11108), .ZN(n11109) );
  AOI21_X1 U13534 ( .B1(n11260), .B2(n14494), .A(n11109), .ZN(n11110) );
  OAI211_X1 U13535 ( .C1(n11112), .C2(n13865), .A(n11111), .B(n11110), .ZN(
        P1_U3281) );
  NAND2_X1 U13536 ( .A1(n11113), .A2(n9951), .ZN(n11116) );
  AOI22_X1 U13537 ( .A1(n12001), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n11898), 
        .B2(n11114), .ZN(n11115) );
  INV_X1 U13538 ( .A(n13487), .ZN(n11167) );
  XNOR2_X1 U13539 ( .A(n13487), .B(n12911), .ZN(n11117) );
  NAND2_X1 U13540 ( .A1(n13051), .A2(n14633), .ZN(n11118) );
  NAND2_X1 U13541 ( .A1(n11117), .A2(n11118), .ZN(n11330) );
  INV_X1 U13542 ( .A(n11117), .ZN(n11120) );
  INV_X1 U13543 ( .A(n11118), .ZN(n11119) );
  NAND2_X1 U13544 ( .A1(n11120), .A2(n11119), .ZN(n11121) );
  AND2_X1 U13545 ( .A1(n11330), .A2(n11121), .ZN(n11129) );
  INV_X1 U13546 ( .A(n11124), .ZN(n11127) );
  INV_X1 U13547 ( .A(n11125), .ZN(n11126) );
  OAI21_X1 U13548 ( .B1(n11129), .B2(n11128), .A(n11331), .ZN(n11130) );
  NAND2_X1 U13549 ( .A1(n11130), .A2(n13034), .ZN(n11143) );
  NAND2_X1 U13550 ( .A1(n11971), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n11137) );
  NAND2_X1 U13551 ( .A1(n9624), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n11136) );
  NAND2_X1 U13552 ( .A1(n11132), .A2(n11332), .ZN(n11133) );
  AND2_X1 U13553 ( .A1(n11290), .A2(n11133), .ZN(n11335) );
  NAND2_X1 U13554 ( .A1(n7325), .A2(n11335), .ZN(n11135) );
  NAND2_X1 U13555 ( .A1(n9628), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n11134) );
  NAND4_X1 U13556 ( .A1(n11137), .A2(n11136), .A3(n11135), .A4(n11134), .ZN(
        n13050) );
  NAND2_X1 U13557 ( .A1(n13050), .A2(n12987), .ZN(n11139) );
  NAND2_X1 U13558 ( .A1(n13052), .A2(n13004), .ZN(n11138) );
  AND2_X1 U13559 ( .A1(n11139), .A2(n11138), .ZN(n11161) );
  OAI21_X1 U13560 ( .B1(n13015), .B2(n11161), .A(n11140), .ZN(n11141) );
  AOI21_X1 U13561 ( .B1(n11164), .B2(n13025), .A(n11141), .ZN(n11142) );
  OAI211_X1 U13562 ( .C1(n11167), .C2(n13043), .A(n11143), .B(n11142), .ZN(
        P2_U3187) );
  XNOR2_X1 U13563 ( .A(n11145), .B(n11144), .ZN(n11950) );
  INV_X1 U13564 ( .A(n11950), .ZN(n11146) );
  OAI222_X1 U13565 ( .A1(n13523), .A2(n11147), .B1(n13526), .B2(n11146), .C1(
        P2_U3088), .C2(n12063), .ZN(P2_U3305) );
  OR2_X1 U13566 ( .A1(n11867), .A2(n13052), .ZN(n11148) );
  NAND2_X1 U13567 ( .A1(n11149), .A2(n11148), .ZN(n11151) );
  NAND2_X1 U13568 ( .A1(n11867), .A2(n13052), .ZN(n11150) );
  INV_X1 U13569 ( .A(n13051), .ZN(n11152) );
  NAND2_X1 U13570 ( .A1(n13487), .A2(n11152), .ZN(n11284) );
  OR2_X1 U13571 ( .A1(n13487), .A2(n11152), .ZN(n11153) );
  NAND2_X1 U13572 ( .A1(n11284), .A2(n11153), .ZN(n12043) );
  XNOR2_X1 U13573 ( .A(n11307), .B(n12043), .ZN(n13489) );
  OR2_X1 U13574 ( .A1(n11867), .A2(n11156), .ZN(n11157) );
  INV_X1 U13575 ( .A(n11285), .ZN(n11159) );
  AOI21_X1 U13576 ( .B1(n12043), .B2(n11160), .A(n11159), .ZN(n11162) );
  OAI21_X1 U13577 ( .B1(n11162), .B2(n14640), .A(n11161), .ZN(n13485) );
  NOR2_X2 U13578 ( .A1(n11163), .A2(n13487), .ZN(n11300) );
  INV_X1 U13579 ( .A(n11300), .ZN(n11302) );
  AOI211_X1 U13580 ( .C1(n13487), .C2(n11163), .A(n14633), .B(n11300), .ZN(
        n13486) );
  NAND2_X1 U13581 ( .A1(n13486), .A2(n13395), .ZN(n11166) );
  AOI22_X1 U13582 ( .A1(n14653), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n11164), 
        .B2(n14621), .ZN(n11165) );
  OAI211_X1 U13583 ( .C1(n11167), .C2(n14625), .A(n11166), .B(n11165), .ZN(
        n11168) );
  AOI21_X1 U13584 ( .B1(n13485), .B2(n13330), .A(n11168), .ZN(n11169) );
  OAI21_X1 U13585 ( .B1(n13397), .B2(n13489), .A(n11169), .ZN(P2_U3251) );
  NAND2_X1 U13586 ( .A1(n11538), .A2(n14376), .ZN(n11170) );
  NAND2_X1 U13587 ( .A1(n11171), .A2(n11170), .ZN(n11229) );
  INV_X1 U13588 ( .A(n11226), .ZN(n11228) );
  NAND2_X1 U13589 ( .A1(n11229), .A2(n11228), .ZN(n11231) );
  OR2_X1 U13590 ( .A1(n11621), .A2(n13666), .ZN(n11172) );
  INV_X1 U13591 ( .A(n11173), .ZN(n11378) );
  OAI21_X1 U13592 ( .B1(n7340), .B2(n11173), .A(n11382), .ZN(n14406) );
  OR2_X1 U13593 ( .A1(n14340), .A2(n13983), .ZN(n11176) );
  NAND2_X1 U13594 ( .A1(n13666), .A2(n13954), .ZN(n11175) );
  NAND2_X1 U13595 ( .A1(n11176), .A2(n11175), .ZN(n14402) );
  NAND2_X1 U13596 ( .A1(n13966), .A2(n14402), .ZN(n11179) );
  NAND2_X1 U13597 ( .A1(n14466), .A2(n11177), .ZN(n11178) );
  OAI211_X1 U13598 ( .C1(n13966), .C2(n11180), .A(n11179), .B(n11178), .ZN(
        n11184) );
  AOI21_X1 U13599 ( .B1(n11174), .B2(n11234), .A(n13961), .ZN(n11182) );
  NAND2_X1 U13600 ( .A1(n11182), .A2(n11383), .ZN(n14403) );
  NOR2_X1 U13601 ( .A1(n14403), .A2(n13896), .ZN(n11183) );
  AOI211_X1 U13602 ( .C1(n14487), .C2(n11174), .A(n11184), .B(n11183), .ZN(
        n11191) );
  NAND2_X1 U13603 ( .A1(n11186), .A2(n11185), .ZN(n11188) );
  NAND2_X1 U13604 ( .A1(n11538), .A2(n13667), .ZN(n11187) );
  NAND2_X1 U13605 ( .A1(n11188), .A2(n11187), .ZN(n11227) );
  OR2_X1 U13606 ( .A1(n11621), .A2(n14341), .ZN(n11189) );
  XNOR2_X1 U13607 ( .A(n11379), .B(n11173), .ZN(n14408) );
  NAND2_X1 U13608 ( .A1(n14408), .A2(n12154), .ZN(n11190) );
  OAI211_X1 U13609 ( .C1(n14406), .C2(n13991), .A(n11191), .B(n11190), .ZN(
        P1_U3279) );
  AOI22_X1 U13610 ( .A1(n11204), .A2(n12247), .B1(n12259), .B2(n13670), .ZN(
        n11311) );
  NAND2_X1 U13611 ( .A1(n11204), .A2(n12255), .ZN(n11195) );
  NAND2_X1 U13612 ( .A1(n13670), .A2(n12247), .ZN(n11194) );
  NAND2_X1 U13613 ( .A1(n11195), .A2(n11194), .ZN(n11196) );
  XNOR2_X1 U13614 ( .A(n11196), .B(n10099), .ZN(n11313) );
  XOR2_X1 U13615 ( .A(n11311), .B(n11313), .Z(n11197) );
  AOI21_X1 U13616 ( .B1(n11198), .B2(n11197), .A(n11314), .ZN(n11206) );
  OAI21_X1 U13617 ( .B1(n14394), .B2(n11200), .A(n11199), .ZN(n11203) );
  OAI22_X1 U13618 ( .A1(n11201), .A2(n14378), .B1(n14377), .B2(n14379), .ZN(
        n11202) );
  AOI211_X1 U13619 ( .C1(n11204), .C2(n14389), .A(n11203), .B(n11202), .ZN(
        n11205) );
  OAI21_X1 U13620 ( .B1(n11206), .B2(n14384), .A(n11205), .ZN(P1_U3231) );
  NAND2_X1 U13621 ( .A1(n6590), .A2(n11208), .ZN(n11209) );
  XNOR2_X1 U13622 ( .A(n11213), .B(n11664), .ZN(n11274) );
  XNOR2_X1 U13623 ( .A(n11274), .B(n14287), .ZN(n11210) );
  XNOR2_X1 U13624 ( .A(n11277), .B(n11210), .ZN(n11218) );
  AOI21_X1 U13625 ( .B1(n12375), .B2(n12338), .A(n11211), .ZN(n11212) );
  OAI21_X1 U13626 ( .B1(n11420), .B2(n12341), .A(n11212), .ZN(n11215) );
  NOR2_X1 U13627 ( .A1(n11213), .A2(n12354), .ZN(n11214) );
  AOI211_X1 U13628 ( .C1(n11216), .C2(n12358), .A(n11215), .B(n11214), .ZN(
        n11217) );
  OAI21_X1 U13629 ( .B1(n11218), .B2(n12366), .A(n11217), .ZN(P3_U3164) );
  INV_X1 U13630 ( .A(n11961), .ZN(n11221) );
  OR2_X1 U13631 ( .A1(n11219), .A2(P2_U3088), .ZN(n12075) );
  NAND2_X1 U13632 ( .A1(n13519), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n11220) );
  OAI211_X1 U13633 ( .C1(n11221), .C2(n13526), .A(n12075), .B(n11220), .ZN(
        P2_U3304) );
  INV_X1 U13634 ( .A(n11222), .ZN(n11224) );
  OAI222_X1 U13635 ( .A1(P3_U3151), .A2(n11225), .B1(n12886), .B2(n11224), 
        .C1(n11223), .C2(n12883), .ZN(P3_U3271) );
  XNOR2_X1 U13636 ( .A(n11227), .B(n11226), .ZN(n14275) );
  OR2_X1 U13637 ( .A1(n11229), .A2(n11228), .ZN(n11230) );
  NAND2_X1 U13638 ( .A1(n11231), .A2(n11230), .ZN(n14269) );
  NAND2_X1 U13639 ( .A1(n11232), .A2(n11621), .ZN(n11233) );
  NAND2_X1 U13640 ( .A1(n11234), .A2(n11233), .ZN(n14271) );
  OR2_X1 U13641 ( .A1(n14376), .A2(n13982), .ZN(n11236) );
  OR2_X1 U13642 ( .A1(n12166), .A2(n13983), .ZN(n11235) );
  AND2_X1 U13643 ( .A1(n11236), .A2(n11235), .ZN(n14264) );
  INV_X1 U13644 ( .A(n14264), .ZN(n11237) );
  AOI21_X1 U13645 ( .B1(n11621), .B2(n14522), .A(n11237), .ZN(n11238) );
  OAI21_X1 U13646 ( .B1(n14271), .B2(n13961), .A(n11238), .ZN(n11239) );
  AOI21_X1 U13647 ( .B1(n14269), .B2(n14518), .A(n11239), .ZN(n11240) );
  OAI21_X1 U13648 ( .B1(n14478), .B2(n14275), .A(n11240), .ZN(n11246) );
  NAND2_X1 U13649 ( .A1(n11246), .A2(n14540), .ZN(n11241) );
  OAI21_X1 U13650 ( .B1(n14540), .B2(n9937), .A(n11241), .ZN(P1_U3541) );
  NAND2_X1 U13651 ( .A1(n11961), .A2(n11242), .ZN(n11244) );
  OAI211_X1 U13652 ( .C1(n11245), .C2(n14135), .A(n11244), .B(n11243), .ZN(
        P1_U3332) );
  INV_X1 U13653 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n11248) );
  NAND2_X1 U13654 ( .A1(n11246), .A2(n14532), .ZN(n11247) );
  OAI21_X1 U13655 ( .B1(n14532), .B2(n11248), .A(n11247), .ZN(P1_U3498) );
  XNOR2_X1 U13656 ( .A(n11249), .B(n11251), .ZN(n11407) );
  INV_X1 U13657 ( .A(n11407), .ZN(n11258) );
  OAI211_X1 U13658 ( .C1(n11252), .C2(n11251), .A(n11392), .B(n14922), .ZN(
        n11254) );
  AOI22_X1 U13659 ( .A1(n12373), .A2(n14284), .B1(n14286), .B2(n12374), .ZN(
        n11253) );
  NAND2_X1 U13660 ( .A1(n11254), .A2(n11253), .ZN(n11406) );
  INV_X1 U13661 ( .A(n11422), .ZN(n11412) );
  AOI22_X1 U13662 ( .A1(n14944), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n14938), 
        .B2(n11417), .ZN(n11255) );
  OAI21_X1 U13663 ( .B1(n11412), .B2(n14294), .A(n11255), .ZN(n11256) );
  AOI21_X1 U13664 ( .B1(n11406), .B2(n14942), .A(n11256), .ZN(n11257) );
  OAI21_X1 U13665 ( .B1(n11258), .B2(n12727), .A(n11257), .ZN(P3_U3219) );
  AOI211_X1 U13666 ( .C1(n14517), .C2(n11261), .A(n11260), .B(n11259), .ZN(
        n11268) );
  INV_X1 U13667 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n11262) );
  OAI22_X1 U13668 ( .A1(n11538), .A2(n14123), .B1(n14532), .B2(n11262), .ZN(
        n11263) );
  INV_X1 U13669 ( .A(n11263), .ZN(n11264) );
  OAI21_X1 U13670 ( .B1(n11268), .B2(n14530), .A(n11264), .ZN(P1_U3495) );
  AOI22_X1 U13671 ( .A1(n11266), .A2(n11265), .B1(n14537), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n11267) );
  OAI21_X1 U13672 ( .B1(n11268), .B2(n14537), .A(n11267), .ZN(P1_U3540) );
  INV_X1 U13673 ( .A(n11978), .ZN(n11272) );
  OAI222_X1 U13674 ( .A1(n13523), .A2(n11979), .B1(n13526), .B2(n11272), .C1(
        P2_U3088), .C2(n11269), .ZN(P2_U3303) );
  INV_X1 U13675 ( .A(n11270), .ZN(n11271) );
  OAI222_X1 U13676 ( .A1(n14135), .A2(n11273), .B1(n12134), .B2(n11272), .C1(
        P1_U3086), .C2(n11271), .ZN(P1_U3331) );
  NOR2_X1 U13677 ( .A1(n11274), .A2(n14306), .ZN(n11276) );
  INV_X1 U13678 ( .A(n11274), .ZN(n11275) );
  XNOR2_X1 U13679 ( .A(n14295), .B(n11698), .ZN(n11413) );
  XNOR2_X1 U13680 ( .A(n11413), .B(n12374), .ZN(n11278) );
  XNOR2_X1 U13681 ( .A(n11415), .B(n11278), .ZN(n11283) );
  AND2_X1 U13682 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n12391) );
  AOI21_X1 U13683 ( .B1(n12338), .B2(n14287), .A(n12391), .ZN(n11280) );
  NAND2_X1 U13684 ( .A1(n12358), .A2(n14291), .ZN(n11279) );
  OAI211_X1 U13685 ( .C1(n11574), .C2(n12341), .A(n11280), .B(n11279), .ZN(
        n11281) );
  AOI21_X1 U13686 ( .B1(n14322), .B2(n12364), .A(n11281), .ZN(n11282) );
  OAI21_X1 U13687 ( .B1(n11283), .B2(n12366), .A(n11282), .ZN(P3_U3174) );
  AOI22_X1 U13688 ( .A1(n11287), .A2(n11898), .B1(n12001), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n11288) );
  INV_X1 U13689 ( .A(n13050), .ZN(n11343) );
  XOR2_X1 U13690 ( .A(n11346), .B(n12046), .Z(n11299) );
  INV_X1 U13691 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n11289) );
  NAND2_X1 U13692 ( .A1(n11290), .A2(n11289), .ZN(n11291) );
  AND2_X1 U13693 ( .A1(n11353), .A2(n11291), .ZN(n11506) );
  NAND2_X1 U13694 ( .A1(n11506), .A2(n7325), .ZN(n11295) );
  NAND2_X1 U13695 ( .A1(n9624), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n11294) );
  NAND2_X1 U13696 ( .A1(n11971), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n11293) );
  NAND2_X1 U13697 ( .A1(n9628), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n11292) );
  NAND4_X1 U13698 ( .A1(n11295), .A2(n11294), .A3(n11293), .A4(n11292), .ZN(
        n13049) );
  NAND2_X1 U13699 ( .A1(n13049), .A2(n12987), .ZN(n11297) );
  NAND2_X1 U13700 ( .A1(n13051), .A2(n13004), .ZN(n11296) );
  AND2_X1 U13701 ( .A1(n11297), .A2(n11296), .ZN(n11333) );
  INV_X1 U13702 ( .A(n11333), .ZN(n11298) );
  AOI21_X1 U13703 ( .B1(n11299), .B2(n13391), .A(n11298), .ZN(n13483) );
  INV_X1 U13704 ( .A(n11363), .ZN(n11301) );
  AOI211_X1 U13705 ( .C1(n13481), .C2(n11302), .A(n14633), .B(n11301), .ZN(
        n13480) );
  INV_X1 U13706 ( .A(n13481), .ZN(n11304) );
  AOI22_X1 U13707 ( .A1(n14653), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n11335), 
        .B2(n14621), .ZN(n11303) );
  OAI21_X1 U13708 ( .B1(n11304), .B2(n14625), .A(n11303), .ZN(n11309) );
  AND2_X1 U13709 ( .A1(n13487), .A2(n13051), .ZN(n11306) );
  OR2_X1 U13710 ( .A1(n13487), .A2(n13051), .ZN(n11305) );
  XOR2_X1 U13711 ( .A(n11367), .B(n12046), .Z(n13484) );
  NOR2_X1 U13712 ( .A1(n13484), .A2(n13397), .ZN(n11308) );
  AOI211_X1 U13713 ( .C1(n13480), .C2(n13395), .A(n11309), .B(n11308), .ZN(
        n11310) );
  OAI21_X1 U13714 ( .B1(n14653), .B2(n13483), .A(n11310), .ZN(P2_U3250) );
  INV_X1 U13715 ( .A(n11311), .ZN(n11312) );
  NAND2_X1 U13716 ( .A1(n11327), .A2(n12255), .ZN(n11316) );
  NAND2_X1 U13717 ( .A1(n13669), .A2(n12247), .ZN(n11315) );
  NAND2_X1 U13718 ( .A1(n11316), .A2(n11315), .ZN(n11317) );
  XNOR2_X1 U13719 ( .A(n11317), .B(n10099), .ZN(n11522) );
  NOR2_X1 U13720 ( .A1(n14379), .A2(n9810), .ZN(n11318) );
  AOI21_X1 U13721 ( .B1(n11327), .B2(n12247), .A(n11318), .ZN(n11520) );
  XNOR2_X1 U13722 ( .A(n11522), .B(n11520), .ZN(n11319) );
  OAI211_X1 U13723 ( .C1(n6608), .C2(n11319), .A(n14382), .B(n14356), .ZN(
        n11329) );
  AOI21_X1 U13724 ( .B1(n14358), .B2(n11321), .A(n11320), .ZN(n11324) );
  NAND2_X1 U13725 ( .A1(n13649), .A2(n11322), .ZN(n11323) );
  OAI211_X1 U13726 ( .C1(n11325), .C2(n14378), .A(n11324), .B(n11323), .ZN(
        n11326) );
  AOI21_X1 U13727 ( .B1(n11327), .B2(n14389), .A(n11326), .ZN(n11328) );
  NAND2_X1 U13728 ( .A1(n11329), .A2(n11328), .ZN(P1_U3217) );
  NAND2_X1 U13729 ( .A1(n11331), .A2(n11330), .ZN(n11497) );
  XNOR2_X1 U13730 ( .A(n13481), .B(n12960), .ZN(n11498) );
  XNOR2_X1 U13731 ( .A(n11497), .B(n11498), .ZN(n11496) );
  AND2_X1 U13732 ( .A1(n13050), .A2(n14633), .ZN(n11495) );
  XNOR2_X1 U13733 ( .A(n11496), .B(n11495), .ZN(n11338) );
  OAI22_X1 U13734 ( .A1(n13015), .A2(n11333), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11332), .ZN(n11334) );
  AOI21_X1 U13735 ( .B1(n11335), .B2(n13025), .A(n11334), .ZN(n11337) );
  NAND2_X1 U13736 ( .A1(n13481), .A2(n13026), .ZN(n11336) );
  OAI211_X1 U13737 ( .C1(n11338), .C2(n13018), .A(n11337), .B(n11336), .ZN(
        P2_U3213) );
  INV_X1 U13738 ( .A(n11339), .ZN(n11342) );
  OAI222_X1 U13739 ( .A1(n12886), .A2(n11342), .B1(n12883), .B2(n11341), .C1(
        P3_U3151), .C2(n11340), .ZN(P3_U3270) );
  AND2_X1 U13740 ( .A1(n13481), .A2(n11343), .ZN(n11345) );
  OR2_X1 U13741 ( .A1(n13481), .A2(n11343), .ZN(n11344) );
  NAND2_X1 U13742 ( .A1(n11347), .A2(n9951), .ZN(n11350) );
  AOI22_X1 U13743 ( .A1(n11898), .A2(n11348), .B1(n12001), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n11349) );
  INV_X1 U13744 ( .A(n13049), .ZN(n11431) );
  XNOR2_X1 U13745 ( .A(n13476), .B(n11431), .ZN(n12042) );
  XNOR2_X1 U13746 ( .A(n11430), .B(n12042), .ZN(n11361) );
  INV_X1 U13747 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n11359) );
  INV_X1 U13748 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n11352) );
  NAND2_X1 U13749 ( .A1(n11353), .A2(n11352), .ZN(n11354) );
  NAND2_X1 U13750 ( .A1(n11557), .A2(n11354), .ZN(n11445) );
  OR2_X1 U13751 ( .A1(n11445), .A2(n11991), .ZN(n11358) );
  NAND2_X1 U13752 ( .A1(n9624), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n11356) );
  NAND2_X1 U13753 ( .A1(n11971), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n11355) );
  AND2_X1 U13754 ( .A1(n11356), .A2(n11355), .ZN(n11357) );
  OAI211_X1 U13755 ( .C1(n11995), .C2(n11359), .A(n11358), .B(n11357), .ZN(
        n13048) );
  AOI22_X1 U13756 ( .A1(n13048), .A2(n13164), .B1(n13004), .B2(n13050), .ZN(
        n11509) );
  INV_X1 U13757 ( .A(n11509), .ZN(n11360) );
  AOI21_X1 U13758 ( .B1(n11361), .B2(n13391), .A(n11360), .ZN(n13478) );
  OR2_X2 U13759 ( .A1(n11363), .A2(n13476), .ZN(n11442) );
  INV_X1 U13760 ( .A(n11442), .ZN(n11362) );
  AOI211_X1 U13761 ( .C1(n13476), .C2(n11363), .A(n14633), .B(n11362), .ZN(
        n13475) );
  INV_X1 U13762 ( .A(n13476), .ZN(n11365) );
  AOI22_X1 U13763 ( .A1(n14653), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n11506), 
        .B2(n14621), .ZN(n11364) );
  OAI21_X1 U13764 ( .B1(n11365), .B2(n14625), .A(n11364), .ZN(n11371) );
  NOR2_X1 U13765 ( .A1(n13481), .A2(n13050), .ZN(n11366) );
  OR2_X1 U13766 ( .A1(n11368), .A2(n12042), .ZN(n11369) );
  NAND2_X1 U13767 ( .A1(n11426), .A2(n11369), .ZN(n13479) );
  NOR2_X1 U13768 ( .A1(n13479), .A2(n13397), .ZN(n11370) );
  AOI211_X1 U13769 ( .C1(n13475), .C2(n13395), .A(n11371), .B(n11370), .ZN(
        n11372) );
  OAI21_X1 U13770 ( .B1(n14653), .B2(n13478), .A(n11372), .ZN(P2_U3249) );
  INV_X1 U13771 ( .A(n12000), .ZN(n11376) );
  OAI222_X1 U13772 ( .A1(n14135), .A2(n11374), .B1(n12134), .B2(n11376), .C1(
        P1_U3086), .C2(n11373), .ZN(P1_U3330) );
  OAI222_X1 U13773 ( .A1(n13523), .A2(n11377), .B1(n13526), .B2(n11376), .C1(
        P2_U3088), .C2(n11375), .ZN(P2_U3302) );
  INV_X1 U13774 ( .A(n11459), .ZN(n11450) );
  XNOR2_X1 U13775 ( .A(n11451), .B(n11450), .ZN(n14399) );
  INV_X1 U13776 ( .A(n12166), .ZN(n13665) );
  NAND2_X1 U13777 ( .A1(n11174), .A2(n13665), .ZN(n11381) );
  XNOR2_X1 U13778 ( .A(n11458), .B(n11450), .ZN(n14401) );
  NAND2_X1 U13779 ( .A1(n14401), .A2(n14268), .ZN(n11390) );
  AOI211_X1 U13780 ( .C1(n14397), .C2(n11383), .A(n13961), .B(n11465), .ZN(
        n14395) );
  INV_X1 U13781 ( .A(n14397), .ZN(n13654) );
  OR2_X1 U13782 ( .A1(n14366), .A2(n13983), .ZN(n11385) );
  OR2_X1 U13783 ( .A1(n12166), .A2(n13982), .ZN(n11384) );
  NAND2_X1 U13784 ( .A1(n11385), .A2(n11384), .ZN(n14396) );
  AOI22_X1 U13785 ( .A1(n13966), .A2(n14396), .B1(n13650), .B2(n14466), .ZN(
        n11387) );
  NAND2_X1 U13786 ( .A1(n13941), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n11386) );
  OAI211_X1 U13787 ( .C1(n13654), .C2(n13978), .A(n11387), .B(n11386), .ZN(
        n11388) );
  AOI21_X1 U13788 ( .B1(n14395), .B2(n14494), .A(n11388), .ZN(n11389) );
  OAI211_X1 U13789 ( .C1(n14399), .C2(n14274), .A(n11390), .B(n11389), .ZN(
        P1_U3278) );
  NAND2_X1 U13790 ( .A1(n11392), .A2(n11391), .ZN(n11393) );
  XOR2_X1 U13791 ( .A(n11396), .B(n11393), .Z(n11394) );
  OAI222_X1 U13792 ( .A1(n14917), .A2(n12732), .B1(n14919), .B2(n11574), .C1(
        n11394), .C2(n14303), .ZN(n12799) );
  INV_X1 U13793 ( .A(n12799), .ZN(n11401) );
  OAI21_X1 U13794 ( .B1(n11397), .B2(n11396), .A(n11395), .ZN(n12800) );
  AOI22_X1 U13795 ( .A1(n14944), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n14938), 
        .B2(n11576), .ZN(n11398) );
  OAI21_X1 U13796 ( .B1(n12865), .B2(n14294), .A(n11398), .ZN(n11399) );
  AOI21_X1 U13797 ( .B1(n12800), .B2(n12739), .A(n11399), .ZN(n11400) );
  OAI21_X1 U13798 ( .B1(n11401), .B2(n14944), .A(n11400), .ZN(P3_U3218) );
  INV_X1 U13799 ( .A(n11402), .ZN(n11405) );
  OAI222_X1 U13800 ( .A1(n12886), .A2(n11405), .B1(n12883), .B2(n11404), .C1(
        P3_U3151), .C2(n11403), .ZN(P3_U3269) );
  INV_X1 U13801 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12413) );
  AOI21_X1 U13802 ( .B1(n14323), .B2(n11407), .A(n11406), .ZN(n11409) );
  MUX2_X1 U13803 ( .A(n12413), .B(n11409), .S(n15164), .Z(n11408) );
  OAI21_X1 U13804 ( .B1(n11412), .B2(n12803), .A(n11408), .ZN(P3_U3473) );
  INV_X1 U13805 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n11410) );
  MUX2_X1 U13806 ( .A(n11410), .B(n11409), .S(n14993), .Z(n11411) );
  OAI21_X1 U13807 ( .B1(n11412), .B2(n12864), .A(n11411), .ZN(P3_U3432) );
  NOR2_X1 U13808 ( .A1(n11413), .A2(n12374), .ZN(n11414) );
  XNOR2_X1 U13809 ( .A(n11422), .B(n11698), .ZN(n11575) );
  XNOR2_X1 U13810 ( .A(n11575), .B(n14285), .ZN(n11572) );
  XNOR2_X1 U13811 ( .A(n11573), .B(n11572), .ZN(n11424) );
  INV_X1 U13812 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n11416) );
  NOR2_X1 U13813 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11416), .ZN(n12417) );
  AOI21_X1 U13814 ( .B1(n12373), .B2(n12357), .A(n12417), .ZN(n11419) );
  NAND2_X1 U13815 ( .A1(n12358), .A2(n11417), .ZN(n11418) );
  OAI211_X1 U13816 ( .C1(n11420), .C2(n12361), .A(n11419), .B(n11418), .ZN(
        n11421) );
  AOI21_X1 U13817 ( .B1(n11422), .B2(n12364), .A(n11421), .ZN(n11423) );
  OAI21_X1 U13818 ( .B1(n11424), .B2(n12366), .A(n11423), .ZN(P3_U3155) );
  NAND2_X1 U13819 ( .A1(n13476), .A2(n13049), .ZN(n11425) );
  NAND2_X1 U13820 ( .A1(n11427), .A2(n9951), .ZN(n11429) );
  AOI22_X1 U13821 ( .A1(n13138), .A2(n11898), .B1(n12001), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n11428) );
  INV_X1 U13822 ( .A(n13048), .ZN(n11549) );
  XNOR2_X1 U13823 ( .A(n13472), .B(n11549), .ZN(n12044) );
  XNOR2_X1 U13824 ( .A(n11543), .B(n12044), .ZN(n13474) );
  OR2_X1 U13825 ( .A1(n13476), .A2(n11431), .ZN(n11432) );
  NAND2_X1 U13826 ( .A1(n11433), .A2(n11432), .ZN(n11552) );
  XOR2_X1 U13827 ( .A(n11552), .B(n12044), .Z(n11441) );
  XNOR2_X1 U13828 ( .A(n11557), .B(P2_REG3_REG_18__SCAN_IN), .ZN(n13013) );
  NAND2_X1 U13829 ( .A1(n13013), .A2(n7325), .ZN(n11439) );
  INV_X1 U13830 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n14606) );
  NAND2_X1 U13831 ( .A1(n11992), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n11435) );
  NAND2_X1 U13832 ( .A1(n9628), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n11434) );
  OAI211_X1 U13833 ( .C1(n11436), .C2(n14606), .A(n11435), .B(n11434), .ZN(
        n11437) );
  INV_X1 U13834 ( .A(n11437), .ZN(n11438) );
  NAND2_X1 U13835 ( .A1(n11439), .A2(n11438), .ZN(n13198) );
  AND2_X1 U13836 ( .A1(n13049), .A2(n13004), .ZN(n11440) );
  AOI21_X1 U13837 ( .B1(n13198), .B2(n13164), .A(n11440), .ZN(n11594) );
  OAI21_X1 U13838 ( .B1(n11441), .B2(n14640), .A(n11594), .ZN(n13470) );
  INV_X1 U13839 ( .A(n13472), .ZN(n11599) );
  NAND2_X1 U13840 ( .A1(n11442), .A2(n13472), .ZN(n11443) );
  NAND2_X1 U13841 ( .A1(n11443), .A2(n13300), .ZN(n11444) );
  NOR2_X1 U13842 ( .A1(n11564), .A2(n11444), .ZN(n13471) );
  NAND2_X1 U13843 ( .A1(n13471), .A2(n13395), .ZN(n11447) );
  INV_X1 U13844 ( .A(n11445), .ZN(n11596) );
  AOI22_X1 U13845 ( .A1(n14653), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n11596), 
        .B2(n14621), .ZN(n11446) );
  OAI211_X1 U13846 ( .C1(n11599), .C2(n14625), .A(n11447), .B(n11446), .ZN(
        n11448) );
  AOI21_X1 U13847 ( .B1(n13470), .B2(n13330), .A(n11448), .ZN(n11449) );
  OAI21_X1 U13848 ( .B1(n13474), .B2(n13397), .A(n11449), .ZN(P2_U3248) );
  NAND2_X1 U13849 ( .A1(n11451), .A2(n11450), .ZN(n11453) );
  NAND2_X1 U13850 ( .A1(n11453), .A2(n11452), .ZN(n11457) );
  INV_X1 U13851 ( .A(n11457), .ZN(n11455) );
  INV_X1 U13852 ( .A(n12079), .ZN(n11456) );
  AOI21_X1 U13853 ( .B1(n11463), .B2(n11457), .A(n11456), .ZN(n14079) );
  NAND2_X1 U13854 ( .A1(n11460), .A2(n11459), .ZN(n11462) );
  INV_X1 U13855 ( .A(n14340), .ZN(n13664) );
  OR2_X1 U13856 ( .A1(n14397), .A2(n13664), .ZN(n11461) );
  OAI21_X1 U13857 ( .B1(n11464), .B2(n11463), .A(n12101), .ZN(n14081) );
  NAND2_X1 U13858 ( .A1(n14081), .A2(n14268), .ZN(n11473) );
  OAI211_X1 U13859 ( .C1(n11465), .C2(n14124), .A(n13975), .B(n14490), .ZN(
        n14077) );
  INV_X1 U13860 ( .A(n14077), .ZN(n11471) );
  NAND2_X1 U13861 ( .A1(n13953), .A2(n13955), .ZN(n11467) );
  OR2_X1 U13862 ( .A1(n14340), .A2(n13982), .ZN(n11466) );
  NAND2_X1 U13863 ( .A1(n11467), .A2(n11466), .ZN(n14359) );
  INV_X1 U13864 ( .A(n14359), .ZN(n14078) );
  OAI22_X1 U13865 ( .A1(n13941), .A2(n14078), .B1(n14364), .B2(n14483), .ZN(
        n11468) );
  AOI21_X1 U13866 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n13941), .A(n11468), 
        .ZN(n11469) );
  OAI21_X1 U13867 ( .B1(n14124), .B2(n13978), .A(n11469), .ZN(n11470) );
  AOI21_X1 U13868 ( .B1(n11471), .B2(n14494), .A(n11470), .ZN(n11472) );
  OAI211_X1 U13869 ( .C1(n14079), .C2(n14274), .A(n11473), .B(n11472), .ZN(
        P1_U3277) );
  INV_X1 U13870 ( .A(n11474), .ZN(n11479) );
  OAI21_X1 U13871 ( .B1(n11476), .B2(n11475), .A(n14922), .ZN(n11477) );
  AOI21_X1 U13872 ( .B1(n11479), .B2(n11478), .A(n11477), .ZN(n11481) );
  OAI22_X1 U13873 ( .A1(n11601), .A2(n14919), .B1(n12721), .B2(n14917), .ZN(
        n11480) );
  NOR2_X1 U13874 ( .A1(n11481), .A2(n11480), .ZN(n12798) );
  OAI21_X1 U13875 ( .B1(n11484), .B2(n11483), .A(n11482), .ZN(n12796) );
  AOI22_X1 U13876 ( .A1(n14944), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n14938), 
        .B2(n11611), .ZN(n11485) );
  OAI21_X1 U13877 ( .B1(n11608), .B2(n14294), .A(n11485), .ZN(n11486) );
  AOI21_X1 U13878 ( .B1(n12796), .B2(n12739), .A(n11486), .ZN(n11487) );
  OAI21_X1 U13879 ( .B1(n12798), .B2(n14944), .A(n11487), .ZN(P3_U3217) );
  INV_X1 U13880 ( .A(n11774), .ZN(n11514) );
  OAI222_X1 U13881 ( .A1(n13526), .A2(n11514), .B1(n11489), .B2(P2_U3088), 
        .C1(n11488), .C2(n13523), .ZN(P2_U3301) );
  XNOR2_X1 U13882 ( .A(n13476), .B(n12911), .ZN(n11490) );
  NAND2_X1 U13883 ( .A1(n13049), .A2(n14633), .ZN(n11491) );
  NAND2_X1 U13884 ( .A1(n11490), .A2(n11491), .ZN(n11588) );
  INV_X1 U13885 ( .A(n11490), .ZN(n11493) );
  INV_X1 U13886 ( .A(n11491), .ZN(n11492) );
  NAND2_X1 U13887 ( .A1(n11493), .A2(n11492), .ZN(n11494) );
  NAND2_X1 U13888 ( .A1(n11588), .A2(n11494), .ZN(n11505) );
  INV_X1 U13889 ( .A(n11497), .ZN(n11499) );
  INV_X1 U13890 ( .A(n11505), .ZN(n11503) );
  INV_X1 U13891 ( .A(n11589), .ZN(n11504) );
  AOI21_X1 U13892 ( .B1(n11505), .B2(n11502), .A(n11504), .ZN(n11512) );
  NAND2_X1 U13893 ( .A1(n13025), .A2(n11506), .ZN(n11508) );
  OAI211_X1 U13894 ( .C1(n11509), .C2(n13015), .A(n11508), .B(n11507), .ZN(
        n11510) );
  AOI21_X1 U13895 ( .B1(n13476), .B2(n13026), .A(n11510), .ZN(n11511) );
  OAI21_X1 U13896 ( .B1(n11512), .B2(n13018), .A(n11511), .ZN(P2_U3198) );
  OAI222_X1 U13897 ( .A1(P1_U3086), .A2(n11515), .B1(n12134), .B2(n11514), 
        .C1(n11513), .C2(n14135), .ZN(P1_U3329) );
  NAND2_X1 U13898 ( .A1(n14390), .A2(n12255), .ZN(n11517) );
  NAND2_X1 U13899 ( .A1(n13668), .A2(n12247), .ZN(n11516) );
  NAND2_X1 U13900 ( .A1(n11517), .A2(n11516), .ZN(n11518) );
  XNOR2_X1 U13901 ( .A(n11518), .B(n10099), .ZN(n11523) );
  NOR2_X1 U13902 ( .A1(n11532), .A2(n9810), .ZN(n11519) );
  AOI21_X1 U13903 ( .B1(n14390), .B2(n12247), .A(n11519), .ZN(n11524) );
  XNOR2_X1 U13904 ( .A(n11523), .B(n11524), .ZN(n14380) );
  INV_X1 U13905 ( .A(n11520), .ZN(n11521) );
  NAND2_X1 U13906 ( .A1(n11522), .A2(n11521), .ZN(n14381) );
  INV_X1 U13907 ( .A(n11523), .ZN(n11525) );
  NAND2_X1 U13908 ( .A1(n11525), .A2(n11524), .ZN(n11526) );
  OAI22_X1 U13909 ( .A1(n11538), .A2(n12263), .B1(n14376), .B2(n12264), .ZN(
        n11527) );
  XNOR2_X1 U13910 ( .A(n11527), .B(n10099), .ZN(n11615) );
  OAI22_X1 U13911 ( .A1(n11538), .A2(n12264), .B1(n14376), .B2(n9810), .ZN(
        n11614) );
  XNOR2_X1 U13912 ( .A(n11615), .B(n11614), .ZN(n11529) );
  AOI21_X1 U13913 ( .B1(n11528), .B2(n11529), .A(n14384), .ZN(n11531) );
  INV_X1 U13914 ( .A(n11529), .ZN(n11530) );
  NAND2_X1 U13915 ( .A1(n11531), .A2(n11617), .ZN(n11537) );
  OAI22_X1 U13916 ( .A1(n11532), .A2(n14378), .B1(n14377), .B2(n14341), .ZN(
        n11533) );
  AOI211_X1 U13917 ( .C1(n13649), .C2(n11535), .A(n11534), .B(n11533), .ZN(
        n11536) );
  OAI211_X1 U13918 ( .C1(n11538), .C2(n13653), .A(n11537), .B(n11536), .ZN(
        P1_U3224) );
  NAND2_X1 U13919 ( .A1(n11539), .A2(n9951), .ZN(n11541) );
  AOI22_X1 U13920 ( .A1(n13147), .A2(n11898), .B1(n12001), .B2(
        P1_DATAO_REG_18__SCAN_IN), .ZN(n11540) );
  XNOR2_X1 U13921 ( .A(n13466), .B(n13198), .ZN(n12047) );
  OR2_X1 U13922 ( .A1(n13472), .A2(n13048), .ZN(n11542) );
  NAND2_X1 U13923 ( .A1(n13472), .A2(n13048), .ZN(n11544) );
  INV_X1 U13924 ( .A(n13174), .ZN(n11547) );
  AOI21_X1 U13925 ( .B1(n12047), .B2(n11548), .A(n11547), .ZN(n13469) );
  INV_X1 U13926 ( .A(n13013), .ZN(n11562) );
  NOR2_X1 U13927 ( .A1(n13472), .A2(n11549), .ZN(n11551) );
  NAND2_X1 U13928 ( .A1(n13472), .A2(n11549), .ZN(n11550) );
  OAI21_X2 U13929 ( .B1(n11552), .B2(n11551), .A(n11550), .ZN(n13201) );
  XNOR2_X1 U13930 ( .A(n13201), .B(n12047), .ZN(n11553) );
  NAND2_X1 U13931 ( .A1(n11553), .A2(n13391), .ZN(n13467) );
  INV_X1 U13932 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n11561) );
  INV_X1 U13933 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n11555) );
  INV_X1 U13934 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n11554) );
  OAI21_X1 U13935 ( .B1(n11557), .B2(n11555), .A(n11554), .ZN(n11558) );
  NAND2_X1 U13936 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_REG3_REG_19__SCAN_IN), 
        .ZN(n11556) );
  NAND2_X1 U13937 ( .A1(n11558), .A2(n11910), .ZN(n12949) );
  OR2_X1 U13938 ( .A1(n12949), .A2(n11991), .ZN(n11560) );
  AOI22_X1 U13939 ( .A1(n9628), .A2(P2_REG0_REG_19__SCAN_IN), .B1(n11971), 
        .B2(P2_REG1_REG_19__SCAN_IN), .ZN(n11559) );
  OAI211_X1 U13940 ( .C1(n9664), .C2(n11561), .A(n11560), .B(n11559), .ZN(
        n13202) );
  AOI22_X1 U13941 ( .A1(n13202), .A2(n13164), .B1(n13004), .B2(n13048), .ZN(
        n13463) );
  OAI211_X1 U13942 ( .C1(n14646), .C2(n11562), .A(n13467), .B(n13463), .ZN(
        n11563) );
  NAND2_X1 U13943 ( .A1(n11563), .A2(n13330), .ZN(n11571) );
  INV_X1 U13944 ( .A(n11564), .ZN(n11566) );
  INV_X1 U13945 ( .A(n13466), .ZN(n11568) );
  NAND2_X1 U13946 ( .A1(n11568), .A2(n11564), .ZN(n13385) );
  INV_X1 U13947 ( .A(n13385), .ZN(n11565) );
  AOI211_X1 U13948 ( .C1(n13466), .C2(n11566), .A(n14633), .B(n11565), .ZN(
        n13464) );
  INV_X1 U13949 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n11567) );
  OAI22_X1 U13950 ( .A1(n11568), .A2(n14625), .B1(n11567), .B2(n13330), .ZN(
        n11569) );
  AOI21_X1 U13951 ( .B1(n13464), .B2(n13395), .A(n11569), .ZN(n11570) );
  OAI211_X1 U13952 ( .C1(n13469), .C2(n13397), .A(n11571), .B(n11570), .ZN(
        P2_U3247) );
  XNOR2_X1 U13953 ( .A(n12865), .B(n11698), .ZN(n11600) );
  XNOR2_X1 U13954 ( .A(n11600), .B(n11601), .ZN(n11604) );
  XNOR2_X1 U13955 ( .A(n11605), .B(n11604), .ZN(n11582) );
  AND2_X1 U13956 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12449) );
  AOI21_X1 U13957 ( .B1(n14285), .B2(n12338), .A(n12449), .ZN(n11578) );
  NAND2_X1 U13958 ( .A1(n12358), .A2(n11576), .ZN(n11577) );
  OAI211_X1 U13959 ( .C1(n12732), .C2(n12341), .A(n11578), .B(n11577), .ZN(
        n11579) );
  AOI21_X1 U13960 ( .B1(n11580), .B2(n12364), .A(n11579), .ZN(n11581) );
  OAI21_X1 U13961 ( .B1(n11582), .B2(n12366), .A(n11581), .ZN(P3_U3181) );
  XNOR2_X1 U13962 ( .A(n13472), .B(n12911), .ZN(n11583) );
  NAND2_X1 U13963 ( .A1(n13048), .A2(n14633), .ZN(n11584) );
  NAND2_X1 U13964 ( .A1(n11583), .A2(n11584), .ZN(n12889) );
  INV_X1 U13965 ( .A(n11583), .ZN(n11586) );
  INV_X1 U13966 ( .A(n11584), .ZN(n11585) );
  NAND2_X1 U13967 ( .A1(n11586), .A2(n11585), .ZN(n11587) );
  AND2_X1 U13968 ( .A1(n12889), .A2(n11587), .ZN(n11591) );
  OAI21_X1 U13969 ( .B1(n11591), .B2(n11590), .A(n12890), .ZN(n11592) );
  NAND2_X1 U13970 ( .A1(n11592), .A2(n13034), .ZN(n11598) );
  OAI21_X1 U13971 ( .B1(n13015), .B2(n11594), .A(n11593), .ZN(n11595) );
  AOI21_X1 U13972 ( .B1(n11596), .B2(n13025), .A(n11595), .ZN(n11597) );
  OAI211_X1 U13973 ( .C1(n11599), .C2(n13043), .A(n11598), .B(n11597), .ZN(
        P2_U3200) );
  INV_X1 U13974 ( .A(n11600), .ZN(n11602) );
  NOR2_X1 U13975 ( .A1(n11602), .A2(n11601), .ZN(n11603) );
  XNOR2_X1 U13976 ( .A(n11608), .B(n11698), .ZN(n11640) );
  XNOR2_X1 U13977 ( .A(n11640), .B(n12372), .ZN(n11606) );
  XNOR2_X1 U13978 ( .A(n11639), .B(n11606), .ZN(n11613) );
  NAND2_X1 U13979 ( .A1(n12373), .A2(n12338), .ZN(n11607) );
  NAND2_X1 U13980 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12476)
         );
  OAI211_X1 U13981 ( .C1(n12721), .C2(n12341), .A(n11607), .B(n12476), .ZN(
        n11610) );
  NOR2_X1 U13982 ( .A1(n11608), .A2(n12354), .ZN(n11609) );
  AOI211_X1 U13983 ( .C1(n11611), .C2(n12358), .A(n11610), .B(n11609), .ZN(
        n11612) );
  OAI21_X1 U13984 ( .B1(n11613), .B2(n12366), .A(n11612), .ZN(P3_U3166) );
  INV_X1 U13985 ( .A(n11621), .ZN(n14266) );
  NAND2_X1 U13986 ( .A1(n11615), .A2(n11614), .ZN(n11616) );
  NAND2_X1 U13987 ( .A1(n11621), .A2(n12255), .ZN(n11619) );
  NAND2_X1 U13988 ( .A1(n13666), .A2(n12247), .ZN(n11618) );
  NAND2_X1 U13989 ( .A1(n11619), .A2(n11618), .ZN(n11620) );
  XNOR2_X1 U13990 ( .A(n11620), .B(n10099), .ZN(n12162) );
  AOI22_X1 U13991 ( .A1(n11621), .A2(n12247), .B1(n12259), .B2(n13666), .ZN(
        n12160) );
  XNOR2_X1 U13992 ( .A(n12162), .B(n12160), .ZN(n11622) );
  OAI211_X1 U13993 ( .C1(n11623), .C2(n11622), .A(n12164), .B(n14356), .ZN(
        n11628) );
  OAI21_X1 U13994 ( .B1(n13647), .B2(n14264), .A(n11624), .ZN(n11625) );
  AOI21_X1 U13995 ( .B1(n11626), .B2(n13649), .A(n11625), .ZN(n11627) );
  OAI211_X1 U13996 ( .C1(n14266), .C2(n13653), .A(n11628), .B(n11627), .ZN(
        P1_U3234) );
  INV_X1 U13997 ( .A(n11739), .ZN(n14130) );
  OAI222_X1 U13998 ( .A1(n13526), .A2(n14130), .B1(n11629), .B2(P2_U3088), 
        .C1(n11737), .C2(n13523), .ZN(P2_U3298) );
  NOR2_X1 U13999 ( .A1(n11631), .A2(n14292), .ZN(n12559) );
  AOI21_X1 U14000 ( .B1(n12814), .B2(n14942), .A(n12559), .ZN(n12550) );
  NAND2_X1 U14001 ( .A1(n14944), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n11632) );
  OAI211_X1 U14002 ( .C1(n11633), .C2(n14294), .A(n12550), .B(n11632), .ZN(
        P3_U3202) );
  OAI222_X1 U14003 ( .A1(n13523), .A2(n11635), .B1(n13526), .B2(n11634), .C1(
        P2_U3088), .C2(n9330), .ZN(P2_U3306) );
  OAI222_X1 U14004 ( .A1(n13523), .A2(n11637), .B1(n13526), .B2(n11636), .C1(
        P2_U3088), .C2(n13154), .ZN(P2_U3308) );
  NAND2_X1 U14005 ( .A1(n11640), .A2(n12372), .ZN(n11638) );
  INV_X1 U14006 ( .A(n11640), .ZN(n11641) );
  NAND2_X1 U14007 ( .A1(n11641), .A2(n12732), .ZN(n11642) );
  XNOR2_X1 U14008 ( .A(n12314), .B(n11698), .ZN(n11644) );
  XNOR2_X1 U14009 ( .A(n11644), .B(n12721), .ZN(n12315) );
  INV_X1 U14010 ( .A(n12315), .ZN(n11643) );
  INV_X1 U14011 ( .A(n11644), .ZN(n11645) );
  NAND2_X1 U14012 ( .A1(n11645), .A2(n12371), .ZN(n11646) );
  NAND2_X1 U14013 ( .A1(n12317), .A2(n11646), .ZN(n12349) );
  XNOR2_X1 U14014 ( .A(n12345), .B(n11698), .ZN(n11647) );
  XNOR2_X1 U14015 ( .A(n11647), .B(n12703), .ZN(n12348) );
  NAND2_X1 U14016 ( .A1(n12349), .A2(n12348), .ZN(n12347) );
  INV_X1 U14017 ( .A(n11647), .ZN(n11648) );
  NAND2_X1 U14018 ( .A1(n11648), .A2(n12703), .ZN(n11649) );
  NAND2_X1 U14019 ( .A1(n12347), .A2(n11649), .ZN(n12291) );
  XNOR2_X1 U14020 ( .A(n12853), .B(n11698), .ZN(n11650) );
  XNOR2_X1 U14021 ( .A(n11650), .B(n12722), .ZN(n12290) );
  NAND2_X1 U14022 ( .A1(n12291), .A2(n12290), .ZN(n12289) );
  NAND2_X1 U14023 ( .A1(n11650), .A2(n12370), .ZN(n11651) );
  NAND2_X1 U14024 ( .A1(n12289), .A2(n11651), .ZN(n12332) );
  XNOR2_X1 U14025 ( .A(n11652), .B(n11698), .ZN(n11653) );
  XNOR2_X1 U14026 ( .A(n11653), .B(n12704), .ZN(n12331) );
  INV_X1 U14027 ( .A(n11653), .ZN(n11654) );
  NAND2_X1 U14028 ( .A1(n11654), .A2(n12704), .ZN(n11655) );
  XNOR2_X1 U14029 ( .A(n12681), .B(n11698), .ZN(n11657) );
  XNOR2_X1 U14030 ( .A(n11657), .B(n12690), .ZN(n12299) );
  INV_X1 U14031 ( .A(n12299), .ZN(n11656) );
  NAND2_X1 U14032 ( .A1(n11657), .A2(n12690), .ZN(n11658) );
  XNOR2_X1 U14033 ( .A(n12667), .B(n11664), .ZN(n11659) );
  NAND2_X1 U14034 ( .A1(n12337), .A2(n12678), .ZN(n11663) );
  INV_X1 U14035 ( .A(n11659), .ZN(n11660) );
  NAND2_X1 U14036 ( .A1(n11661), .A2(n11660), .ZN(n11662) );
  XNOR2_X1 U14037 ( .A(n12766), .B(n11664), .ZN(n11666) );
  NAND2_X1 U14038 ( .A1(n12282), .A2(n12659), .ZN(n11669) );
  INV_X1 U14039 ( .A(n11665), .ZN(n11667) );
  NAND2_X1 U14040 ( .A1(n11669), .A2(n11668), .ZN(n12323) );
  XNOR2_X1 U14041 ( .A(n12634), .B(n11698), .ZN(n11670) );
  XNOR2_X1 U14042 ( .A(n11670), .B(n12647), .ZN(n12324) );
  NAND2_X1 U14043 ( .A1(n12323), .A2(n12324), .ZN(n11672) );
  NAND2_X1 U14044 ( .A1(n11670), .A2(n12285), .ZN(n11671) );
  XNOR2_X1 U14045 ( .A(n12311), .B(n11698), .ZN(n11673) );
  XNOR2_X1 U14046 ( .A(n11673), .B(n12627), .ZN(n12306) );
  NAND2_X1 U14047 ( .A1(n11673), .A2(n12362), .ZN(n11674) );
  XNOR2_X1 U14048 ( .A(n12752), .B(n11698), .ZN(n11676) );
  XNOR2_X1 U14049 ( .A(n11676), .B(n12614), .ZN(n12356) );
  XNOR2_X1 U14050 ( .A(n11677), .B(n11698), .ZN(n11694) );
  XNOR2_X1 U14051 ( .A(n11694), .B(n12600), .ZN(n11696) );
  XNOR2_X1 U14052 ( .A(n11697), .B(n11696), .ZN(n11678) );
  NAND2_X1 U14053 ( .A1(n11678), .A2(n12346), .ZN(n11682) );
  AOI22_X1 U14054 ( .A1(n12589), .A2(n12358), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11679) );
  OAI21_X1 U14055 ( .B1(n12309), .B2(n12361), .A(n11679), .ZN(n11680) );
  AOI21_X1 U14056 ( .B1(n12357), .B2(n12585), .A(n11680), .ZN(n11681) );
  OAI211_X1 U14057 ( .C1(n12828), .C2(n12354), .A(n11682), .B(n11681), .ZN(
        P3_U3154) );
  INV_X1 U14058 ( .A(n11752), .ZN(n13521) );
  OAI222_X1 U14059 ( .A1(n14135), .A2(n11683), .B1(n12134), .B2(n13521), .C1(
        n8741), .C2(P1_U3086), .ZN(P1_U3327) );
  INV_X1 U14060 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n11684) );
  INV_X1 U14061 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n13681) );
  OAI22_X1 U14062 ( .A1(n13966), .A2(n11684), .B1(n13681), .B2(n14483), .ZN(
        n11687) );
  NOR2_X1 U14063 ( .A1(n14270), .A2(n11685), .ZN(n11686) );
  AOI211_X1 U14064 ( .C1(n14268), .C2(n11688), .A(n11687), .B(n11686), .ZN(
        n11692) );
  OAI21_X1 U14065 ( .B1(n11690), .B2(n11689), .A(n13966), .ZN(n11691) );
  OAI211_X1 U14066 ( .C1(n11693), .C2(n13978), .A(n11692), .B(n11691), .ZN(
        P1_U3292) );
  AND2_X1 U14067 ( .A1(n11694), .A2(n12567), .ZN(n11695) );
  XNOR2_X1 U14068 ( .A(n12575), .B(n11698), .ZN(n11699) );
  XNOR2_X1 U14069 ( .A(n11700), .B(n11699), .ZN(n11706) );
  NOR2_X1 U14070 ( .A1(n12568), .A2(n12341), .ZN(n11703) );
  AOI22_X1 U14071 ( .A1(n12577), .A2(n12358), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11701) );
  OAI21_X1 U14072 ( .B1(n12567), .B2(n12361), .A(n11701), .ZN(n11702) );
  AOI211_X1 U14073 ( .C1(n11704), .C2(n12364), .A(n11703), .B(n11702), .ZN(
        n11705) );
  OAI21_X1 U14074 ( .B1(n11706), .B2(n12366), .A(n11705), .ZN(P3_U3160) );
  NAND2_X1 U14075 ( .A1(n13514), .A2(n9951), .ZN(n11709) );
  INV_X1 U14076 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n11707) );
  OR2_X1 U14077 ( .A1(n11980), .A2(n11707), .ZN(n11708) );
  NAND2_X1 U14078 ( .A1(n11971), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n11712) );
  NAND2_X1 U14079 ( .A1(n9624), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n11711) );
  NAND2_X1 U14080 ( .A1(n9628), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n11710) );
  NAND3_X1 U14081 ( .A1(n11712), .A2(n11711), .A3(n11710), .ZN(n13044) );
  XNOR2_X1 U14082 ( .A(n13166), .B(n13044), .ZN(n12055) );
  NAND2_X1 U14083 ( .A1(n11971), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n11715) );
  NAND2_X1 U14084 ( .A1(n9624), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n11714) );
  NAND2_X1 U14085 ( .A1(n9628), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n11713) );
  NAND3_X1 U14086 ( .A1(n11715), .A2(n11714), .A3(n11713), .ZN(n13045) );
  NAND2_X1 U14087 ( .A1(n11716), .A2(n9951), .ZN(n11718) );
  OR2_X1 U14088 ( .A1(n11980), .A2(n12077), .ZN(n11717) );
  MUX2_X1 U14089 ( .A(n13045), .B(n12022), .S(n11720), .Z(n11789) );
  INV_X4 U14090 ( .A(n12013), .ZN(n12014) );
  OAI211_X1 U14091 ( .C1(n11721), .C2(n12024), .A(n12056), .B(n12071), .ZN(
        n11722) );
  AOI21_X1 U14092 ( .B1(n13044), .B2(n12014), .A(n11722), .ZN(n11723) );
  INV_X1 U14093 ( .A(n13045), .ZN(n13230) );
  NOR2_X1 U14094 ( .A1(n11723), .A2(n13230), .ZN(n11724) );
  AOI21_X1 U14095 ( .B1(n12022), .B2(n12013), .A(n11724), .ZN(n11790) );
  INV_X1 U14096 ( .A(n11926), .ZN(n11726) );
  NAND2_X1 U14097 ( .A1(n11726), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n11942) );
  INV_X1 U14098 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n11941) );
  NAND2_X1 U14099 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(P2_REG3_REG_23__SCAN_IN), 
        .ZN(n11727) );
  INV_X1 U14100 ( .A(n11988), .ZN(n11728) );
  NAND2_X1 U14101 ( .A1(n11728), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n11990) );
  INV_X1 U14102 ( .A(n11990), .ZN(n11729) );
  NAND2_X1 U14103 ( .A1(n11729), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n11767) );
  INV_X1 U14104 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n12932) );
  INV_X1 U14105 ( .A(n11757), .ZN(n11730) );
  NAND2_X1 U14106 ( .A1(n11730), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n13236) );
  OR2_X1 U14107 ( .A1(n13236), .A2(n11991), .ZN(n11736) );
  INV_X1 U14108 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n11733) );
  NAND2_X1 U14109 ( .A1(n11971), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n11732) );
  NAND2_X1 U14110 ( .A1(n11992), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n11731) );
  OAI211_X1 U14111 ( .C1(n11995), .C2(n11733), .A(n11732), .B(n11731), .ZN(
        n11734) );
  INV_X1 U14112 ( .A(n11734), .ZN(n11735) );
  NAND2_X1 U14113 ( .A1(n11736), .A2(n11735), .ZN(n13046) );
  INV_X1 U14114 ( .A(n13046), .ZN(n11740) );
  NOR2_X1 U14115 ( .A1(n11980), .A2(n11737), .ZN(n11738) );
  AOI21_X2 U14116 ( .B1(n11739), .B2(n9951), .A(n11738), .ZN(n13403) );
  MUX2_X1 U14117 ( .A(n11740), .B(n13403), .S(n12014), .Z(n11781) );
  INV_X1 U14118 ( .A(n11720), .ZN(n12004) );
  NAND2_X1 U14119 ( .A1(n11781), .A2(n11780), .ZN(n11743) );
  OAI21_X1 U14120 ( .B1(n11789), .B2(n11790), .A(n11743), .ZN(n11744) );
  INV_X1 U14121 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n11745) );
  NAND2_X1 U14122 ( .A1(n11757), .A2(n11745), .ZN(n11746) );
  NAND2_X1 U14123 ( .A1(n13236), .A2(n11746), .ZN(n13250) );
  INV_X1 U14124 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13249) );
  NAND2_X1 U14125 ( .A1(n11971), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n11748) );
  NAND2_X1 U14126 ( .A1(n9628), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n11747) );
  OAI211_X1 U14127 ( .C1(n13249), .C2(n9664), .A(n11748), .B(n11747), .ZN(
        n11749) );
  INV_X1 U14128 ( .A(n11749), .ZN(n11750) );
  INV_X1 U14129 ( .A(n13224), .ZN(n13227) );
  NAND2_X1 U14130 ( .A1(n11752), .A2(n9951), .ZN(n11754) );
  OR2_X1 U14131 ( .A1(n11980), .A2(n15043), .ZN(n11753) );
  INV_X1 U14132 ( .A(n13410), .ZN(n13223) );
  MUX2_X1 U14133 ( .A(n13227), .B(n13223), .S(n11720), .Z(n11783) );
  MUX2_X1 U14134 ( .A(n13224), .B(n13410), .S(n12004), .Z(n11782) );
  NAND2_X1 U14135 ( .A1(n11783), .A2(n11782), .ZN(n11755) );
  NAND2_X1 U14136 ( .A1(n11767), .A2(n12932), .ZN(n11756) );
  NAND2_X1 U14137 ( .A1(n13268), .A2(n7325), .ZN(n11763) );
  INV_X1 U14138 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n11760) );
  NAND2_X1 U14139 ( .A1(n11992), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n11759) );
  NAND2_X1 U14140 ( .A1(n11971), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n11758) );
  OAI211_X1 U14141 ( .C1(n11760), .C2(n11995), .A(n11759), .B(n11758), .ZN(
        n11761) );
  INV_X1 U14142 ( .A(n11761), .ZN(n11762) );
  NAND2_X1 U14143 ( .A1(n11763), .A2(n11762), .ZN(n13222) );
  NAND2_X1 U14144 ( .A1(n13522), .A2(n9951), .ZN(n11765) );
  NAND2_X1 U14145 ( .A1(n12001), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n11764) );
  MUX2_X1 U14146 ( .A(n13195), .B(n13416), .S(n11720), .Z(n11778) );
  MUX2_X1 U14147 ( .A(n13222), .B(n13265), .S(n12004), .Z(n11777) );
  INV_X1 U14148 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n13037) );
  NAND2_X1 U14149 ( .A1(n11990), .A2(n13037), .ZN(n11766) );
  NAND2_X1 U14150 ( .A1(n11767), .A2(n11766), .ZN(n13281) );
  OR2_X1 U14151 ( .A1(n13281), .A2(n11991), .ZN(n11773) );
  INV_X1 U14152 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n11770) );
  NAND2_X1 U14153 ( .A1(n11971), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n11769) );
  NAND2_X1 U14154 ( .A1(n11992), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n11768) );
  OAI211_X1 U14155 ( .C1(n11995), .C2(n11770), .A(n11769), .B(n11768), .ZN(
        n11771) );
  INV_X1 U14156 ( .A(n11771), .ZN(n11772) );
  NAND2_X1 U14157 ( .A1(n11773), .A2(n11772), .ZN(n13193) );
  INV_X1 U14158 ( .A(n13193), .ZN(n13220) );
  NAND2_X1 U14159 ( .A1(n11774), .A2(n9951), .ZN(n11776) );
  NAND2_X1 U14160 ( .A1(n12001), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n11775) );
  INV_X1 U14161 ( .A(n13420), .ZN(n13284) );
  MUX2_X1 U14162 ( .A(n13220), .B(n13284), .S(n12014), .Z(n12010) );
  MUX2_X1 U14163 ( .A(n13193), .B(n13420), .S(n12013), .Z(n12009) );
  OR3_X1 U14164 ( .A1(n12008), .A2(n12010), .A3(n12009), .ZN(n11795) );
  OR3_X1 U14165 ( .A1(n11779), .A2(n11778), .A3(n11777), .ZN(n11794) );
  INV_X1 U14166 ( .A(n11780), .ZN(n11787) );
  INV_X1 U14167 ( .A(n11781), .ZN(n11786) );
  INV_X1 U14168 ( .A(n11782), .ZN(n11785) );
  INV_X1 U14169 ( .A(n11783), .ZN(n11784) );
  AOI22_X1 U14170 ( .A1(n11787), .A2(n11786), .B1(n11785), .B2(n11784), .ZN(
        n11788) );
  NAND2_X1 U14171 ( .A1(n12055), .A2(n11788), .ZN(n11791) );
  AOI22_X1 U14172 ( .A1(n11792), .A2(n11791), .B1(n11790), .B2(n11789), .ZN(
        n11793) );
  NAND2_X1 U14173 ( .A1(n11802), .A2(n11803), .ZN(n11796) );
  NAND2_X1 U14174 ( .A1(n11796), .A2(n11720), .ZN(n11801) );
  NAND2_X1 U14175 ( .A1(n11798), .A2(n11797), .ZN(n11800) );
  MUX2_X1 U14176 ( .A(n11801), .B(n11800), .S(n11799), .Z(n11805) );
  MUX2_X1 U14177 ( .A(n11803), .B(n11720), .S(n11802), .Z(n11804) );
  NAND2_X1 U14178 ( .A1(n11805), .A2(n11804), .ZN(n11809) );
  INV_X1 U14179 ( .A(n11809), .ZN(n11812) );
  MUX2_X1 U14180 ( .A(n13064), .B(n11806), .S(n11720), .Z(n11811) );
  INV_X1 U14181 ( .A(n11811), .ZN(n11808) );
  MUX2_X1 U14182 ( .A(n13064), .B(n11806), .S(n12013), .Z(n11807) );
  OAI21_X1 U14183 ( .B1(n11809), .B2(n11808), .A(n11807), .ZN(n11810) );
  OAI211_X1 U14184 ( .C1(n11812), .C2(n11811), .A(n11810), .B(n12025), .ZN(
        n11820) );
  OAI21_X1 U14185 ( .B1(n13063), .B2(n12013), .A(n11813), .ZN(n11817) );
  NAND2_X1 U14186 ( .A1(n13063), .A2(n12004), .ZN(n11815) );
  NAND2_X1 U14187 ( .A1(n11815), .A2(n11814), .ZN(n11816) );
  NAND2_X1 U14188 ( .A1(n11817), .A2(n11816), .ZN(n11819) );
  NAND3_X1 U14189 ( .A1(n11820), .A2(n11819), .A3(n11818), .ZN(n11825) );
  NAND2_X1 U14190 ( .A1(n13062), .A2(n12014), .ZN(n11821) );
  NAND2_X1 U14191 ( .A1(n11821), .A2(n14677), .ZN(n11823) );
  OAI21_X1 U14192 ( .B1(n13062), .B2(n12014), .A(n14634), .ZN(n11822) );
  NAND2_X1 U14193 ( .A1(n11823), .A2(n11822), .ZN(n11824) );
  NAND2_X1 U14194 ( .A1(n11825), .A2(n11824), .ZN(n11827) );
  MUX2_X1 U14195 ( .A(n13061), .B(n14683), .S(n12013), .Z(n11828) );
  MUX2_X1 U14196 ( .A(n13061), .B(n14683), .S(n12014), .Z(n11826) );
  INV_X1 U14197 ( .A(n11828), .ZN(n11829) );
  MUX2_X1 U14198 ( .A(n13060), .B(n14690), .S(n11720), .Z(n11831) );
  MUX2_X1 U14199 ( .A(n13060), .B(n14690), .S(n12004), .Z(n11830) );
  MUX2_X1 U14200 ( .A(n14702), .B(n13059), .S(n12014), .Z(n11834) );
  INV_X1 U14201 ( .A(n11720), .ZN(n11901) );
  MUX2_X1 U14202 ( .A(n14702), .B(n13059), .S(n11901), .Z(n11832) );
  INV_X1 U14203 ( .A(n11834), .ZN(n11835) );
  MUX2_X1 U14204 ( .A(n13058), .B(n14619), .S(n12014), .Z(n11839) );
  MUX2_X1 U14205 ( .A(n14619), .B(n13058), .S(n12014), .Z(n11836) );
  NAND2_X1 U14206 ( .A1(n11837), .A2(n11836), .ZN(n11843) );
  INV_X1 U14207 ( .A(n11838), .ZN(n11841) );
  INV_X1 U14208 ( .A(n11839), .ZN(n11840) );
  NAND2_X1 U14209 ( .A1(n11841), .A2(n11840), .ZN(n11842) );
  NAND2_X1 U14210 ( .A1(n11843), .A2(n11842), .ZN(n11845) );
  MUX2_X1 U14211 ( .A(n13057), .B(n14710), .S(n11901), .Z(n11846) );
  MUX2_X1 U14212 ( .A(n13057), .B(n14710), .S(n11720), .Z(n11844) );
  INV_X1 U14213 ( .A(n11846), .ZN(n11847) );
  MUX2_X1 U14214 ( .A(n13056), .B(n11848), .S(n12014), .Z(n11851) );
  MUX2_X1 U14215 ( .A(n13056), .B(n11848), .S(n11901), .Z(n11849) );
  INV_X1 U14216 ( .A(n11851), .ZN(n11852) );
  MUX2_X1 U14217 ( .A(n13055), .B(n14720), .S(n11901), .Z(n11855) );
  MUX2_X1 U14218 ( .A(n13055), .B(n14720), .S(n12014), .Z(n11853) );
  INV_X1 U14219 ( .A(n11855), .ZN(n11856) );
  MUX2_X1 U14220 ( .A(n13054), .B(n13491), .S(n12014), .Z(n11859) );
  MUX2_X1 U14221 ( .A(n13054), .B(n13491), .S(n11901), .Z(n11857) );
  NAND2_X1 U14222 ( .A1(n11858), .A2(n11857), .ZN(n11861) );
  NAND2_X1 U14223 ( .A1(n6554), .A2(n7161), .ZN(n11860) );
  NAND2_X1 U14224 ( .A1(n11861), .A2(n11860), .ZN(n11864) );
  MUX2_X1 U14225 ( .A(n13053), .B(n11862), .S(n11901), .Z(n11865) );
  MUX2_X1 U14226 ( .A(n13053), .B(n11862), .S(n12014), .Z(n11863) );
  INV_X1 U14227 ( .A(n11865), .ZN(n11866) );
  MUX2_X1 U14228 ( .A(n13052), .B(n11867), .S(n12014), .Z(n11871) );
  MUX2_X1 U14229 ( .A(n13052), .B(n11867), .S(n11901), .Z(n11868) );
  NAND2_X1 U14230 ( .A1(n11869), .A2(n11868), .ZN(n11875) );
  INV_X1 U14231 ( .A(n11870), .ZN(n11873) );
  INV_X1 U14232 ( .A(n11871), .ZN(n11872) );
  NAND2_X1 U14233 ( .A1(n11873), .A2(n11872), .ZN(n11874) );
  NAND2_X1 U14234 ( .A1(n11875), .A2(n11874), .ZN(n11877) );
  MUX2_X1 U14235 ( .A(n13051), .B(n13487), .S(n11901), .Z(n11878) );
  MUX2_X1 U14236 ( .A(n13051), .B(n13487), .S(n11720), .Z(n11876) );
  INV_X1 U14237 ( .A(n11878), .ZN(n11879) );
  MUX2_X1 U14238 ( .A(n13050), .B(n13481), .S(n12014), .Z(n11882) );
  MUX2_X1 U14239 ( .A(n13050), .B(n13481), .S(n11901), .Z(n11880) );
  INV_X1 U14240 ( .A(n11882), .ZN(n11883) );
  MUX2_X1 U14241 ( .A(n13049), .B(n13476), .S(n11901), .Z(n11886) );
  MUX2_X1 U14242 ( .A(n13049), .B(n13476), .S(n11720), .Z(n11884) );
  INV_X1 U14243 ( .A(n11886), .ZN(n11887) );
  MUX2_X1 U14244 ( .A(n13048), .B(n13472), .S(n11720), .Z(n11890) );
  MUX2_X1 U14245 ( .A(n13048), .B(n13472), .S(n11901), .Z(n11888) );
  NAND2_X1 U14246 ( .A1(n11889), .A2(n11888), .ZN(n11892) );
  NAND2_X1 U14247 ( .A1(n11892), .A2(n11891), .ZN(n11894) );
  MUX2_X1 U14248 ( .A(n13198), .B(n13466), .S(n11901), .Z(n11895) );
  MUX2_X1 U14249 ( .A(n13198), .B(n13466), .S(n12014), .Z(n11893) );
  INV_X1 U14250 ( .A(n11895), .ZN(n11896) );
  NAND2_X1 U14251 ( .A1(n11897), .A2(n9951), .ZN(n11900) );
  AOI22_X1 U14252 ( .A1(n12001), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n10176), 
        .B2(n11898), .ZN(n11899) );
  MUX2_X1 U14253 ( .A(n13202), .B(n13459), .S(n11720), .Z(n11905) );
  MUX2_X1 U14254 ( .A(n13202), .B(n13459), .S(n11901), .Z(n11902) );
  NAND2_X1 U14255 ( .A1(n11903), .A2(n11902), .ZN(n11909) );
  INV_X1 U14256 ( .A(n11904), .ZN(n11907) );
  INV_X1 U14257 ( .A(n11905), .ZN(n11906) );
  NAND2_X1 U14258 ( .A1(n11907), .A2(n11906), .ZN(n11908) );
  NAND2_X1 U14259 ( .A1(n11909), .A2(n11908), .ZN(n11922) );
  INV_X1 U14260 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n15055) );
  NAND2_X1 U14261 ( .A1(n11910), .A2(n15055), .ZN(n11911) );
  NAND2_X1 U14262 ( .A1(n11926), .A2(n11911), .ZN(n12998) );
  OR2_X1 U14263 ( .A1(n12998), .A2(n11991), .ZN(n11917) );
  INV_X1 U14264 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n11914) );
  NAND2_X1 U14265 ( .A1(n11971), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n11913) );
  NAND2_X1 U14266 ( .A1(n11992), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n11912) );
  OAI211_X1 U14267 ( .C1(n11914), .C2(n11995), .A(n11913), .B(n11912), .ZN(
        n11915) );
  INV_X1 U14268 ( .A(n11915), .ZN(n11916) );
  NAND2_X1 U14269 ( .A1(n11917), .A2(n11916), .ZN(n13177) );
  NAND2_X1 U14270 ( .A1(n11918), .A2(n9951), .ZN(n11920) );
  NAND2_X1 U14271 ( .A1(n12001), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n11919) );
  MUX2_X1 U14272 ( .A(n13177), .B(n13452), .S(n12004), .Z(n11923) );
  MUX2_X1 U14273 ( .A(n13177), .B(n13452), .S(n12014), .Z(n11921) );
  INV_X1 U14274 ( .A(n11923), .ZN(n11924) );
  INV_X1 U14275 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n11925) );
  NAND2_X1 U14276 ( .A1(n11926), .A2(n11925), .ZN(n11927) );
  NAND2_X1 U14277 ( .A1(n11942), .A2(n11927), .ZN(n13359) );
  OR2_X1 U14278 ( .A1(n13359), .A2(n11991), .ZN(n11933) );
  INV_X1 U14279 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n11930) );
  NAND2_X1 U14280 ( .A1(n11971), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n11929) );
  NAND2_X1 U14281 ( .A1(n11992), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n11928) );
  OAI211_X1 U14282 ( .C1(n11995), .C2(n11930), .A(n11929), .B(n11928), .ZN(
        n11931) );
  INV_X1 U14283 ( .A(n11931), .ZN(n11932) );
  NAND2_X1 U14284 ( .A1(n11933), .A2(n11932), .ZN(n13208) );
  NAND2_X1 U14285 ( .A1(n11934), .A2(n9951), .ZN(n11936) );
  NAND2_X1 U14286 ( .A1(n12001), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n11935) );
  MUX2_X1 U14287 ( .A(n13208), .B(n13447), .S(n12014), .Z(n11939) );
  MUX2_X1 U14288 ( .A(n13208), .B(n13447), .S(n12004), .Z(n11937) );
  INV_X1 U14289 ( .A(n11939), .ZN(n11940) );
  NAND2_X1 U14290 ( .A1(n11942), .A2(n11941), .ZN(n11943) );
  NAND2_X1 U14291 ( .A1(n11969), .A2(n11943), .ZN(n13343) );
  OR2_X1 U14292 ( .A1(n13343), .A2(n11991), .ZN(n11949) );
  INV_X1 U14293 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n11946) );
  NAND2_X1 U14294 ( .A1(n11992), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n11945) );
  NAND2_X1 U14295 ( .A1(n11971), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n11944) );
  OAI211_X1 U14296 ( .C1(n11946), .C2(n11995), .A(n11945), .B(n11944), .ZN(
        n11947) );
  INV_X1 U14297 ( .A(n11947), .ZN(n11948) );
  NAND2_X1 U14298 ( .A1(n11949), .A2(n11948), .ZN(n13183) );
  NAND2_X1 U14299 ( .A1(n11950), .A2(n9951), .ZN(n11952) );
  NAND2_X1 U14300 ( .A1(n12001), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n11951) );
  NAND2_X2 U14301 ( .A1(n11952), .A2(n11951), .ZN(n13442) );
  MUX2_X1 U14302 ( .A(n13183), .B(n13442), .S(n12004), .Z(n11955) );
  MUX2_X1 U14303 ( .A(n13183), .B(n13442), .S(n11720), .Z(n11953) );
  INV_X1 U14304 ( .A(n11955), .ZN(n11956) );
  XNOR2_X1 U14305 ( .A(n11969), .B(P2_REG3_REG_23__SCAN_IN), .ZN(n13334) );
  INV_X1 U14306 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n11959) );
  NAND2_X1 U14307 ( .A1(n11992), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n11958) );
  NAND2_X1 U14308 ( .A1(n11971), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n11957) );
  OAI211_X1 U14309 ( .C1(n11959), .C2(n11995), .A(n11958), .B(n11957), .ZN(
        n11960) );
  AOI21_X1 U14310 ( .B1(n13334), .B2(n7325), .A(n11960), .ZN(n13212) );
  INV_X1 U14311 ( .A(n13212), .ZN(n13047) );
  NAND2_X1 U14312 ( .A1(n11961), .A2(n9951), .ZN(n11963) );
  NAND2_X1 U14313 ( .A1(n12001), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n11962) );
  MUX2_X1 U14314 ( .A(n13047), .B(n13438), .S(n12014), .Z(n11966) );
  MUX2_X1 U14315 ( .A(n13047), .B(n13438), .S(n12004), .Z(n11964) );
  NAND2_X1 U14316 ( .A1(n11965), .A2(n11964), .ZN(n11968) );
  NAND2_X1 U14317 ( .A1(n6556), .A2(n7151), .ZN(n11967) );
  NAND2_X1 U14318 ( .A1(n11968), .A2(n11967), .ZN(n11984) );
  INV_X1 U14319 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n12940) );
  INV_X1 U14320 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n12990) );
  OAI21_X1 U14321 ( .B1(n11969), .B2(n12940), .A(n12990), .ZN(n11970) );
  AND2_X1 U14322 ( .A1(n11988), .A2(n11970), .ZN(n13319) );
  NAND2_X1 U14323 ( .A1(n13319), .A2(n7325), .ZN(n11977) );
  INV_X1 U14324 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n11974) );
  NAND2_X1 U14325 ( .A1(n9628), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n11973) );
  NAND2_X1 U14326 ( .A1(n11971), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n11972) );
  OAI211_X1 U14327 ( .C1(n9664), .C2(n11974), .A(n11973), .B(n11972), .ZN(
        n11975) );
  INV_X1 U14328 ( .A(n11975), .ZN(n11976) );
  NAND2_X1 U14329 ( .A1(n11977), .A2(n11976), .ZN(n13187) );
  NAND2_X1 U14330 ( .A1(n11978), .A2(n9951), .ZN(n11982) );
  OR2_X1 U14331 ( .A1(n11980), .A2(n11979), .ZN(n11981) );
  MUX2_X1 U14332 ( .A(n13187), .B(n13432), .S(n12004), .Z(n11985) );
  MUX2_X1 U14333 ( .A(n13187), .B(n13432), .S(n12014), .Z(n11983) );
  INV_X1 U14334 ( .A(n11985), .ZN(n11986) );
  INV_X1 U14335 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n11987) );
  NAND2_X1 U14336 ( .A1(n11988), .A2(n11987), .ZN(n11989) );
  NAND2_X1 U14337 ( .A1(n11990), .A2(n11989), .ZN(n13301) );
  OR2_X1 U14338 ( .A1(n13301), .A2(n11991), .ZN(n11999) );
  INV_X1 U14339 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n11996) );
  NAND2_X1 U14340 ( .A1(n11992), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n11994) );
  NAND2_X1 U14341 ( .A1(n11971), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n11993) );
  OAI211_X1 U14342 ( .C1(n11996), .C2(n11995), .A(n11994), .B(n11993), .ZN(
        n11997) );
  INV_X1 U14343 ( .A(n11997), .ZN(n11998) );
  NAND2_X1 U14344 ( .A1(n11999), .A2(n11998), .ZN(n13190) );
  NAND2_X1 U14345 ( .A1(n12000), .A2(n9951), .ZN(n12003) );
  NAND2_X1 U14346 ( .A1(n12001), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n12002) );
  MUX2_X1 U14347 ( .A(n13190), .B(n13304), .S(n12014), .Z(n12006) );
  MUX2_X1 U14348 ( .A(n13190), .B(n13304), .S(n12004), .Z(n12005) );
  INV_X1 U14349 ( .A(n12008), .ZN(n12012) );
  NAND2_X1 U14350 ( .A1(n12010), .A2(n12009), .ZN(n12011) );
  NAND2_X1 U14351 ( .A1(n13044), .A2(n12013), .ZN(n12016) );
  INV_X1 U14352 ( .A(n13044), .ZN(n13165) );
  NAND2_X1 U14353 ( .A1(n13165), .A2(n12014), .ZN(n12015) );
  MUX2_X1 U14354 ( .A(n12016), .B(n12015), .S(n13166), .Z(n12017) );
  INV_X1 U14355 ( .A(n12017), .ZN(n12018) );
  AOI21_X1 U14356 ( .B1(n12056), .B2(n13154), .A(n12019), .ZN(n12020) );
  OAI21_X1 U14357 ( .B1(n12072), .B2(n12021), .A(n12020), .ZN(n12060) );
  XNOR2_X1 U14358 ( .A(n12022), .B(n13045), .ZN(n12053) );
  XNOR2_X1 U14359 ( .A(n13265), .B(n13195), .ZN(n13259) );
  XNOR2_X1 U14360 ( .A(n13420), .B(n13220), .ZN(n13219) );
  INV_X1 U14361 ( .A(n13190), .ZN(n13218) );
  XNOR2_X1 U14362 ( .A(n13304), .B(n13218), .ZN(n13189) );
  INV_X1 U14363 ( .A(n13187), .ZN(n13215) );
  XNOR2_X1 U14364 ( .A(n13432), .B(n13215), .ZN(n13312) );
  OR2_X1 U14365 ( .A1(n13438), .A2(n13047), .ZN(n13185) );
  NAND2_X1 U14366 ( .A1(n13438), .A2(n13047), .ZN(n13186) );
  NAND2_X1 U14367 ( .A1(n13185), .A2(n13186), .ZN(n13326) );
  OR2_X1 U14368 ( .A1(n13447), .A2(n13208), .ZN(n13182) );
  NAND2_X1 U14369 ( .A1(n13447), .A2(n13208), .ZN(n13180) );
  NAND2_X1 U14370 ( .A1(n13182), .A2(n13180), .ZN(n13364) );
  NAND4_X1 U14371 ( .A1(n12026), .A2(n12025), .A3(n12024), .A4(n12023), .ZN(
        n12028) );
  NOR3_X1 U14372 ( .A1(n12028), .A2(n12027), .A3(n14639), .ZN(n12031) );
  NAND4_X1 U14373 ( .A1(n12032), .A2(n12031), .A3(n12030), .A4(n12029), .ZN(
        n12033) );
  NOR2_X1 U14374 ( .A1(n12034), .A2(n12033), .ZN(n12037) );
  NAND4_X1 U14375 ( .A1(n12038), .A2(n12037), .A3(n12036), .A4(n12035), .ZN(
        n12039) );
  OR4_X1 U14376 ( .A1(n12042), .A2(n12041), .A3(n12040), .A4(n12039), .ZN(
        n12045) );
  OR2_X1 U14377 ( .A1(n13459), .A2(n13202), .ZN(n13176) );
  NAND2_X1 U14378 ( .A1(n13459), .A2(n13202), .ZN(n13175) );
  NAND2_X1 U14379 ( .A1(n13176), .A2(n13175), .ZN(n13390) );
  AND4_X1 U14380 ( .A1(n13364), .A2(n6512), .A3(n12047), .A4(n13390), .ZN(
        n12048) );
  XNOR2_X1 U14381 ( .A(n13442), .B(n13183), .ZN(n13347) );
  XNOR2_X1 U14382 ( .A(n13452), .B(n13177), .ZN(n13378) );
  NAND4_X1 U14383 ( .A1(n13326), .A2(n12048), .A3(n13347), .A4(n13378), .ZN(
        n12049) );
  OR4_X1 U14384 ( .A1(n13219), .A2(n13189), .A3(n13312), .A4(n12049), .ZN(
        n12050) );
  NOR2_X1 U14385 ( .A1(n13259), .A2(n12050), .ZN(n12052) );
  XNOR2_X1 U14386 ( .A(n13235), .B(n13046), .ZN(n13225) );
  NAND2_X1 U14387 ( .A1(n13410), .A2(n13224), .ZN(n13196) );
  OR2_X1 U14388 ( .A1(n13410), .A2(n13224), .ZN(n12051) );
  NAND2_X1 U14389 ( .A1(n13196), .A2(n12051), .ZN(n13242) );
  AND4_X1 U14390 ( .A1(n12053), .A2(n12052), .A3(n13225), .A4(n13242), .ZN(
        n12054) );
  AOI21_X1 U14391 ( .B1(n12057), .B2(n10176), .A(n12056), .ZN(n12065) );
  INV_X1 U14392 ( .A(n12057), .ZN(n12058) );
  OAI21_X1 U14393 ( .B1(n13154), .B2(n12062), .A(n12058), .ZN(n12059) );
  AOI22_X1 U14394 ( .A1(n12061), .A2(n12060), .B1(n12065), .B2(n12059), .ZN(
        n12070) );
  INV_X1 U14395 ( .A(n12061), .ZN(n12068) );
  AOI21_X1 U14396 ( .B1(n12063), .B2(n12062), .A(n9330), .ZN(n12064) );
  NAND2_X1 U14397 ( .A1(n12068), .A2(n12067), .ZN(n12069) );
  AND2_X1 U14398 ( .A1(n12070), .A2(n12069), .ZN(n12076) );
  INV_X1 U14399 ( .A(n14661), .ZN(n14659) );
  NOR4_X1 U14400 ( .A1(n14659), .A2(n13228), .A3(n12071), .A4(n13525), .ZN(
        n12074) );
  OAI21_X1 U14401 ( .B1(n12075), .B2(n12072), .A(P2_B_REG_SCAN_IN), .ZN(n12073) );
  OAI22_X1 U14402 ( .A1(n12076), .A2(n12075), .B1(n12074), .B2(n12073), .ZN(
        P2_U3328) );
  INV_X1 U14403 ( .A(n11716), .ZN(n12133) );
  OAI222_X1 U14404 ( .A1(n13526), .A2(n12133), .B1(n9348), .B2(P2_U3088), .C1(
        n12077), .C2(n13523), .ZN(P2_U3297) );
  INV_X1 U14405 ( .A(n14028), .ZN(n12093) );
  INV_X1 U14406 ( .A(n13581), .ZN(n13827) );
  OR2_X1 U14407 ( .A1(n14124), .A2(n13663), .ZN(n12078) );
  INV_X1 U14408 ( .A(n13972), .ZN(n13980) );
  OR2_X1 U14409 ( .A1(n13980), .A2(n13950), .ZN(n12083) );
  INV_X1 U14410 ( .A(n13953), .ZN(n12080) );
  OR2_X1 U14411 ( .A1(n14372), .A2(n12080), .ZN(n13949) );
  OR2_X1 U14412 ( .A1(n13950), .A2(n13949), .ZN(n12082) );
  INV_X1 U14413 ( .A(n13662), .ZN(n14365) );
  OR2_X1 U14414 ( .A1(n13967), .A2(n14365), .ZN(n12081) );
  INV_X1 U14415 ( .A(n13956), .ZN(n12084) );
  INV_X1 U14416 ( .A(n13907), .ZN(n12108) );
  NOR2_X1 U14417 ( .A1(n14051), .A2(n12086), .ZN(n12087) );
  INV_X1 U14418 ( .A(n13885), .ZN(n12088) );
  NAND2_X1 U14419 ( .A1(n13883), .A2(n12088), .ZN(n12090) );
  INV_X1 U14420 ( .A(n13901), .ZN(n13568) );
  NAND2_X1 U14421 ( .A1(n13888), .A2(n13568), .ZN(n12089) );
  NAND2_X1 U14422 ( .A1(n12090), .A2(n12089), .ZN(n13873) );
  INV_X1 U14423 ( .A(n13869), .ZN(n14108) );
  INV_X1 U14424 ( .A(n13831), .ZN(n13825) );
  NAND2_X1 U14425 ( .A1(n13826), .A2(n13825), .ZN(n13824) );
  INV_X1 U14426 ( .A(n13809), .ZN(n13820) );
  INV_X1 U14427 ( .A(n14014), .ZN(n12094) );
  NOR2_X1 U14428 ( .A1(n12094), .A2(n13658), .ZN(n12095) );
  OR3_X1 U14429 ( .A1(n13790), .A2(n6575), .A3(n12095), .ZN(n12096) );
  NAND2_X1 U14430 ( .A1(n13656), .A2(n13955), .ZN(n12098) );
  NAND2_X1 U14431 ( .A1(n13658), .A2(n13954), .ZN(n12097) );
  NAND2_X1 U14432 ( .A1(n14124), .A2(n14366), .ZN(n12100) );
  NAND2_X1 U14433 ( .A1(n13948), .A2(n12103), .ZN(n12104) );
  OR2_X1 U14434 ( .A1(n14063), .A2(n13956), .ZN(n12105) );
  INV_X1 U14435 ( .A(n13917), .ZN(n13912) );
  OR2_X1 U14436 ( .A1(n14114), .A2(n13938), .ZN(n12107) );
  NAND2_X1 U14437 ( .A1(n13886), .A2(n13885), .ZN(n13884) );
  OR2_X1 U14438 ( .A1(n13888), .A2(n13901), .ZN(n12109) );
  NAND2_X1 U14439 ( .A1(n13884), .A2(n12109), .ZN(n13866) );
  INV_X1 U14440 ( .A(n13866), .ZN(n12110) );
  NAND2_X1 U14441 ( .A1(n13869), .A2(n13660), .ZN(n12111) );
  INV_X1 U14442 ( .A(n13849), .ZN(n13846) );
  NAND2_X1 U14443 ( .A1(n14104), .A2(n13581), .ZN(n12112) );
  NAND2_X1 U14444 ( .A1(n13843), .A2(n12112), .ZN(n13818) );
  INV_X1 U14445 ( .A(n13818), .ZN(n13832) );
  NAND2_X1 U14446 ( .A1(n13640), .A2(n13828), .ZN(n12114) );
  INV_X1 U14447 ( .A(n12114), .ZN(n12113) );
  NOR2_X1 U14448 ( .A1(n12113), .A2(n13809), .ZN(n12116) );
  NAND2_X1 U14449 ( .A1(n14028), .A2(n13659), .ZN(n13819) );
  AND2_X1 U14450 ( .A1(n13819), .A2(n12114), .ZN(n12115) );
  OR2_X1 U14451 ( .A1(n12116), .A2(n12115), .ZN(n12117) );
  OR2_X1 U14452 ( .A1(n14014), .A2(n13658), .ZN(n12119) );
  AND2_X1 U14453 ( .A1(n12120), .A2(n6575), .ZN(n12121) );
  OR2_X2 U14454 ( .A1(n6514), .A2(n12121), .ZN(n14013) );
  INV_X1 U14455 ( .A(n12122), .ZN(n12272) );
  NAND2_X1 U14456 ( .A1(n13941), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n12123) );
  OAI21_X1 U14457 ( .B1(n14483), .B2(n12272), .A(n12123), .ZN(n12124) );
  AOI21_X1 U14458 ( .B1(n14009), .B2(n14487), .A(n12124), .ZN(n12128) );
  NOR2_X1 U14459 ( .A1(n13962), .A2(n14063), .ZN(n13937) );
  NAND2_X1 U14460 ( .A1(n14114), .A2(n13937), .ZN(n13925) );
  NAND2_X1 U14461 ( .A1(n14009), .A2(n6515), .ZN(n12126) );
  AND2_X1 U14462 ( .A1(n12142), .A2(n12126), .ZN(n14010) );
  NAND2_X1 U14463 ( .A1(n14010), .A2(n13989), .ZN(n12127) );
  OAI211_X1 U14464 ( .C1(n14013), .C2(n13991), .A(n12128), .B(n12127), .ZN(
        n12129) );
  INV_X1 U14465 ( .A(n12129), .ZN(n12130) );
  OAI21_X1 U14466 ( .B1(n14012), .B2(n14498), .A(n12130), .ZN(P1_U3265) );
  INV_X1 U14467 ( .A(n12131), .ZN(n12135) );
  OAI222_X1 U14468 ( .A1(n12135), .A2(P1_U3086), .B1(n12134), .B2(n12133), 
        .C1(n12132), .C2(n14135), .ZN(P1_U3325) );
  XNOR2_X1 U14469 ( .A(n12137), .B(n12136), .ZN(n14008) );
  AOI211_X1 U14470 ( .C1(n12143), .C2(n12142), .A(n13961), .B(n13782), .ZN(
        n13998) );
  NAND2_X1 U14471 ( .A1(n13998), .A2(n14494), .ZN(n12152) );
  INV_X1 U14472 ( .A(P1_B_REG_SCAN_IN), .ZN(n12144) );
  NOR2_X1 U14473 ( .A1(n14132), .A2(n12144), .ZN(n12145) );
  NOR2_X1 U14474 ( .A1(n13983), .A2(n12145), .ZN(n13777) );
  NAND2_X1 U14475 ( .A1(n13777), .A2(n13655), .ZN(n14000) );
  INV_X1 U14476 ( .A(n12146), .ZN(n12147) );
  OAI22_X1 U14477 ( .A1(n12148), .A2(n14000), .B1(n12147), .B2(n14483), .ZN(
        n12150) );
  NAND2_X1 U14478 ( .A1(n13657), .A2(n13954), .ZN(n13999) );
  NOR2_X1 U14479 ( .A1(n13941), .A2(n13999), .ZN(n12149) );
  AOI211_X1 U14480 ( .C1(n14498), .C2(P1_REG2_REG_29__SCAN_IN), .A(n12150), 
        .B(n12149), .ZN(n12151) );
  OAI211_X1 U14481 ( .C1(n14001), .C2(n13978), .A(n12152), .B(n12151), .ZN(
        n12153) );
  AOI21_X1 U14482 ( .B1(n14006), .B2(n12154), .A(n12153), .ZN(n12155) );
  OAI21_X1 U14483 ( .B1(n14008), .B2(n13991), .A(n12155), .ZN(P1_U3356) );
  INV_X1 U14484 ( .A(n12156), .ZN(n12158) );
  OAI222_X1 U14485 ( .A1(n12883), .A2(n12159), .B1(n12886), .B2(n12158), .C1(
        n12157), .C2(P3_U3151), .ZN(P3_U3266) );
  INV_X1 U14486 ( .A(n12160), .ZN(n12161) );
  NAND2_X1 U14487 ( .A1(n12162), .A2(n12161), .ZN(n12163) );
  INV_X1 U14488 ( .A(n11174), .ZN(n12167) );
  OAI22_X1 U14489 ( .A1(n12167), .A2(n12263), .B1(n12166), .B2(n12264), .ZN(
        n12165) );
  XNOR2_X1 U14490 ( .A(n12165), .B(n10099), .ZN(n12169) );
  OAI22_X1 U14491 ( .A1(n12167), .A2(n12264), .B1(n12166), .B2(n9810), .ZN(
        n12170) );
  XNOR2_X1 U14492 ( .A(n12169), .B(n12170), .ZN(n14342) );
  INV_X1 U14493 ( .A(n12169), .ZN(n12172) );
  INV_X1 U14494 ( .A(n12170), .ZN(n12171) );
  NAND2_X1 U14495 ( .A1(n12172), .A2(n12171), .ZN(n12173) );
  NAND2_X1 U14496 ( .A1(n14397), .A2(n12255), .ZN(n12176) );
  OR2_X1 U14497 ( .A1(n14340), .A2(n12174), .ZN(n12175) );
  NAND2_X1 U14498 ( .A1(n12176), .A2(n12175), .ZN(n12178) );
  XNOR2_X1 U14499 ( .A(n12178), .B(n12177), .ZN(n12180) );
  NOR2_X1 U14500 ( .A1(n12182), .A2(n12180), .ZN(n14352) );
  OAI22_X1 U14501 ( .A1(n14124), .A2(n12263), .B1(n14366), .B2(n12264), .ZN(
        n12179) );
  XNOR2_X1 U14502 ( .A(n12179), .B(n10099), .ZN(n12185) );
  OAI22_X1 U14503 ( .A1(n14124), .A2(n12264), .B1(n14366), .B2(n9810), .ZN(
        n12184) );
  XNOR2_X1 U14504 ( .A(n12185), .B(n12184), .ZN(n14351) );
  NOR2_X1 U14505 ( .A1(n14352), .A2(n14351), .ZN(n12183) );
  INV_X1 U14506 ( .A(n12180), .ZN(n12181) );
  OAI22_X1 U14507 ( .A1(n13654), .A2(n12264), .B1(n14340), .B2(n9810), .ZN(
        n13644) );
  NAND2_X1 U14508 ( .A1(n12183), .A2(n13643), .ZN(n14354) );
  OR2_X1 U14509 ( .A1(n12185), .A2(n12184), .ZN(n12186) );
  NAND2_X1 U14510 ( .A1(n14354), .A2(n12186), .ZN(n14367) );
  NAND2_X1 U14511 ( .A1(n14372), .A2(n12255), .ZN(n12188) );
  NAND2_X1 U14512 ( .A1(n13953), .A2(n12247), .ZN(n12187) );
  NAND2_X1 U14513 ( .A1(n12188), .A2(n12187), .ZN(n12189) );
  XNOR2_X1 U14514 ( .A(n12189), .B(n10099), .ZN(n12190) );
  AOI22_X1 U14515 ( .A1(n14372), .A2(n12247), .B1(n12259), .B2(n13953), .ZN(
        n12191) );
  XNOR2_X1 U14516 ( .A(n12190), .B(n12191), .ZN(n14368) );
  NAND2_X1 U14517 ( .A1(n14367), .A2(n14368), .ZN(n13552) );
  INV_X1 U14518 ( .A(n12190), .ZN(n12192) );
  NAND2_X1 U14519 ( .A1(n12192), .A2(n12191), .ZN(n13614) );
  NAND2_X1 U14520 ( .A1(n13967), .A2(n12255), .ZN(n12194) );
  NAND2_X1 U14521 ( .A1(n13662), .A2(n12247), .ZN(n12193) );
  NAND2_X1 U14522 ( .A1(n12194), .A2(n12193), .ZN(n12195) );
  XNOR2_X1 U14523 ( .A(n12195), .B(n10099), .ZN(n12208) );
  INV_X1 U14524 ( .A(n12208), .ZN(n12196) );
  AOI22_X1 U14525 ( .A1(n13967), .A2(n12247), .B1(n12259), .B2(n13662), .ZN(
        n12207) );
  NAND2_X1 U14526 ( .A1(n12196), .A2(n12207), .ZN(n12206) );
  AND2_X1 U14527 ( .A1(n13614), .A2(n12206), .ZN(n13553) );
  AND2_X1 U14528 ( .A1(n13956), .A2(n12259), .ZN(n12197) );
  AOI21_X1 U14529 ( .B1(n14063), .B2(n12247), .A(n12197), .ZN(n12203) );
  NAND2_X1 U14530 ( .A1(n14063), .A2(n12255), .ZN(n12199) );
  NAND2_X1 U14531 ( .A1(n13956), .A2(n12247), .ZN(n12198) );
  NAND2_X1 U14532 ( .A1(n12199), .A2(n12198), .ZN(n12200) );
  XNOR2_X1 U14533 ( .A(n12200), .B(n10099), .ZN(n12205) );
  XOR2_X1 U14534 ( .A(n12203), .B(n12205), .Z(n13560) );
  INV_X1 U14535 ( .A(n13560), .ZN(n12201) );
  AND2_X1 U14536 ( .A1(n13553), .A2(n12201), .ZN(n13556) );
  OAI22_X1 U14537 ( .A1(n14114), .A2(n12264), .B1(n13938), .B2(n9810), .ZN(
        n12213) );
  OAI22_X1 U14538 ( .A1(n14114), .A2(n12263), .B1(n13938), .B2(n12264), .ZN(
        n12202) );
  XNOR2_X1 U14539 ( .A(n12202), .B(n10099), .ZN(n12214) );
  XOR2_X1 U14540 ( .A(n12213), .B(n12214), .Z(n13597) );
  AND2_X1 U14541 ( .A1(n13556), .A2(n13597), .ZN(n12212) );
  INV_X1 U14542 ( .A(n13597), .ZN(n12211) );
  INV_X1 U14543 ( .A(n12203), .ZN(n12204) );
  NAND2_X1 U14544 ( .A1(n12205), .A2(n12204), .ZN(n12210) );
  INV_X1 U14545 ( .A(n12206), .ZN(n12209) );
  XNOR2_X1 U14546 ( .A(n12208), .B(n12207), .ZN(n13616) );
  OR2_X1 U14547 ( .A1(n12209), .A2(n13616), .ZN(n13554) );
  OR2_X1 U14548 ( .A1(n13560), .A2(n13554), .ZN(n13557) );
  AND2_X1 U14549 ( .A1(n12210), .A2(n13557), .ZN(n13594) );
  NAND2_X1 U14550 ( .A1(n12214), .A2(n12213), .ZN(n12215) );
  AOI22_X1 U14551 ( .A1(n14051), .A2(n12255), .B1(n12247), .B2(n13661), .ZN(
        n12216) );
  XNOR2_X1 U14552 ( .A(n12216), .B(n10099), .ZN(n12219) );
  AOI22_X1 U14553 ( .A1(n14051), .A2(n12247), .B1(n12259), .B2(n13661), .ZN(
        n12218) );
  XNOR2_X1 U14554 ( .A(n12219), .B(n12218), .ZN(n13565) );
  INV_X1 U14555 ( .A(n13565), .ZN(n12217) );
  NOR2_X1 U14556 ( .A1(n13568), .A2(n9810), .ZN(n12220) );
  AOI21_X1 U14557 ( .B1(n13888), .B2(n12247), .A(n12220), .ZN(n12222) );
  AOI22_X1 U14558 ( .A1(n13888), .A2(n12255), .B1(n12247), .B2(n13901), .ZN(
        n12221) );
  XNOR2_X1 U14559 ( .A(n12221), .B(n10099), .ZN(n12223) );
  XOR2_X1 U14560 ( .A(n12222), .B(n12223), .Z(n13606) );
  NAND2_X1 U14561 ( .A1(n12223), .A2(n12222), .ZN(n12224) );
  NAND2_X1 U14562 ( .A1(n13604), .A2(n12224), .ZN(n13535) );
  NAND2_X1 U14563 ( .A1(n13869), .A2(n12255), .ZN(n12226) );
  NAND2_X1 U14564 ( .A1(n13660), .A2(n12247), .ZN(n12225) );
  NAND2_X1 U14565 ( .A1(n12226), .A2(n12225), .ZN(n12227) );
  XNOR2_X1 U14566 ( .A(n12227), .B(n10099), .ZN(n12228) );
  AOI22_X1 U14567 ( .A1(n13869), .A2(n12247), .B1(n12259), .B2(n13660), .ZN(
        n12229) );
  XNOR2_X1 U14568 ( .A(n12228), .B(n12229), .ZN(n13536) );
  NAND2_X1 U14569 ( .A1(n13535), .A2(n13536), .ZN(n13574) );
  INV_X1 U14570 ( .A(n12228), .ZN(n12230) );
  NAND2_X1 U14571 ( .A1(n12230), .A2(n12229), .ZN(n13573) );
  OAI22_X1 U14572 ( .A1(n14104), .A2(n12263), .B1(n13581), .B2(n12264), .ZN(
        n12231) );
  XNOR2_X1 U14573 ( .A(n12231), .B(n10099), .ZN(n12239) );
  INV_X1 U14574 ( .A(n12239), .ZN(n12233) );
  OAI22_X1 U14575 ( .A1(n14104), .A2(n12264), .B1(n13581), .B2(n9810), .ZN(
        n12240) );
  INV_X1 U14576 ( .A(n12240), .ZN(n12232) );
  NAND2_X1 U14577 ( .A1(n12233), .A2(n12232), .ZN(n13575) );
  NAND2_X1 U14578 ( .A1(n14028), .A2(n12255), .ZN(n12235) );
  NAND2_X1 U14579 ( .A1(n13659), .A2(n12247), .ZN(n12234) );
  NAND2_X1 U14580 ( .A1(n12235), .A2(n12234), .ZN(n12236) );
  XNOR2_X1 U14581 ( .A(n12236), .B(n10099), .ZN(n12244) );
  INV_X1 U14582 ( .A(n12244), .ZN(n12237) );
  AOI22_X1 U14583 ( .A1(n14028), .A2(n12247), .B1(n12259), .B2(n13659), .ZN(
        n12243) );
  NAND2_X1 U14584 ( .A1(n12237), .A2(n12243), .ZN(n12242) );
  AND2_X1 U14585 ( .A1(n13575), .A2(n12242), .ZN(n12238) );
  AND2_X1 U14586 ( .A1(n13573), .A2(n12238), .ZN(n12246) );
  INV_X1 U14587 ( .A(n12238), .ZN(n12241) );
  XOR2_X1 U14588 ( .A(n12240), .B(n12239), .Z(n13587) );
  INV_X1 U14589 ( .A(n12242), .ZN(n12245) );
  XNOR2_X1 U14590 ( .A(n12244), .B(n12243), .ZN(n13578) );
  NAND2_X1 U14591 ( .A1(n13640), .A2(n12255), .ZN(n12249) );
  NAND2_X1 U14592 ( .A1(n13828), .A2(n12247), .ZN(n12248) );
  NAND2_X1 U14593 ( .A1(n12249), .A2(n12248), .ZN(n12250) );
  XNOR2_X1 U14594 ( .A(n12250), .B(n10099), .ZN(n12251) );
  AOI22_X1 U14595 ( .A1(n13640), .A2(n12247), .B1(n12259), .B2(n13828), .ZN(
        n12252) );
  XNOR2_X1 U14596 ( .A(n12251), .B(n12252), .ZN(n13634) );
  INV_X1 U14597 ( .A(n12251), .ZN(n12253) );
  NAND2_X1 U14598 ( .A1(n12253), .A2(n12252), .ZN(n12254) );
  NAND2_X1 U14599 ( .A1(n14014), .A2(n12255), .ZN(n12257) );
  NAND2_X1 U14600 ( .A1(n13658), .A2(n12247), .ZN(n12256) );
  NAND2_X1 U14601 ( .A1(n12257), .A2(n12256), .ZN(n12258) );
  XNOR2_X1 U14602 ( .A(n12258), .B(n10099), .ZN(n12260) );
  AOI22_X1 U14603 ( .A1(n14014), .A2(n12247), .B1(n12259), .B2(n13658), .ZN(
        n12261) );
  XNOR2_X1 U14604 ( .A(n12260), .B(n12261), .ZN(n13528) );
  INV_X1 U14605 ( .A(n12260), .ZN(n12262) );
  OAI22_X1 U14606 ( .A1(n12265), .A2(n12263), .B1(n13794), .B2(n12264), .ZN(
        n12268) );
  OAI22_X1 U14607 ( .A1(n12265), .A2(n12264), .B1(n13794), .B2(n9810), .ZN(
        n12266) );
  XNOR2_X1 U14608 ( .A(n12266), .B(n10099), .ZN(n12267) );
  XOR2_X1 U14609 ( .A(n12268), .B(n12267), .Z(n12269) );
  XNOR2_X1 U14610 ( .A(n12270), .B(n12269), .ZN(n12278) );
  OAI22_X1 U14611 ( .A1(n14394), .A2(n12272), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12271), .ZN(n12276) );
  OAI22_X1 U14612 ( .A1(n12274), .A2(n14378), .B1(n14377), .B2(n12273), .ZN(
        n12275) );
  AOI211_X1 U14613 ( .C1(n14009), .C2(n14389), .A(n12276), .B(n12275), .ZN(
        n12277) );
  OAI21_X1 U14614 ( .B1(n12278), .B2(n14384), .A(n12277), .ZN(P1_U3220) );
  INV_X1 U14615 ( .A(n12279), .ZN(n12280) );
  OAI222_X1 U14616 ( .A1(n7368), .A2(P3_U3151), .B1(n12870), .B2(n12281), .C1(
        n12886), .C2(n12280), .ZN(P3_U3265) );
  XNOR2_X1 U14617 ( .A(n12282), .B(n12626), .ZN(n12288) );
  AOI22_X1 U14618 ( .A1(n12646), .A2(n12338), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12284) );
  NAND2_X1 U14619 ( .A1(n12651), .A2(n12358), .ZN(n12283) );
  OAI211_X1 U14620 ( .C1(n12285), .C2(n12341), .A(n12284), .B(n12283), .ZN(
        n12286) );
  AOI21_X1 U14621 ( .B1(n12766), .B2(n12364), .A(n12286), .ZN(n12287) );
  OAI21_X1 U14622 ( .B1(n12288), .B2(n12366), .A(n12287), .ZN(P3_U3156) );
  OAI211_X1 U14623 ( .C1(n12291), .C2(n12290), .A(n12289), .B(n12346), .ZN(
        n12295) );
  NAND2_X1 U14624 ( .A1(n12338), .A2(n12703), .ZN(n12292) );
  NAND2_X1 U14625 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12542)
         );
  OAI211_X1 U14626 ( .C1(n12677), .C2(n12341), .A(n12292), .B(n12542), .ZN(
        n12293) );
  AOI21_X1 U14627 ( .B1(n12708), .B2(n12358), .A(n12293), .ZN(n12294) );
  OAI211_X1 U14628 ( .C1(n12354), .C2(n12853), .A(n12295), .B(n12294), .ZN(
        P3_U3159) );
  INV_X1 U14629 ( .A(n12296), .ZN(n12297) );
  AOI21_X1 U14630 ( .B1(n12299), .B2(n12298), .A(n12297), .ZN(n12304) );
  AOI22_X1 U14631 ( .A1(n12704), .A2(n12338), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12301) );
  NAND2_X1 U14632 ( .A1(n12682), .A2(n12358), .ZN(n12300) );
  OAI211_X1 U14633 ( .C1(n12678), .C2(n12341), .A(n12301), .B(n12300), .ZN(
        n12302) );
  AOI21_X1 U14634 ( .B1(n12681), .B2(n12364), .A(n12302), .ZN(n12303) );
  OAI21_X1 U14635 ( .B1(n12304), .B2(n12366), .A(n12303), .ZN(P3_U3163) );
  XOR2_X1 U14636 ( .A(n12306), .B(n12305), .Z(n12313) );
  AOI22_X1 U14637 ( .A1(n12647), .A2(n12338), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12308) );
  NAND2_X1 U14638 ( .A1(n12618), .A2(n12358), .ZN(n12307) );
  OAI211_X1 U14639 ( .C1(n12309), .C2(n12341), .A(n12308), .B(n12307), .ZN(
        n12310) );
  AOI21_X1 U14640 ( .B1(n12311), .B2(n12364), .A(n12310), .ZN(n12312) );
  OAI21_X1 U14641 ( .B1(n12313), .B2(n12366), .A(n12312), .ZN(P3_U3165) );
  AOI21_X1 U14642 ( .B1(n12316), .B2(n12315), .A(n12366), .ZN(n12318) );
  NAND2_X1 U14643 ( .A1(n12318), .A2(n12317), .ZN(n12322) );
  NAND2_X1 U14644 ( .A1(n12357), .A2(n12703), .ZN(n12319) );
  NAND2_X1 U14645 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n12493)
         );
  OAI211_X1 U14646 ( .C1(n12732), .C2(n12361), .A(n12319), .B(n12493), .ZN(
        n12320) );
  AOI21_X1 U14647 ( .B1(n12736), .B2(n12358), .A(n12320), .ZN(n12321) );
  OAI211_X1 U14648 ( .C1(n12860), .C2(n12354), .A(n12322), .B(n12321), .ZN(
        P3_U3168) );
  XOR2_X1 U14649 ( .A(n12324), .B(n12323), .Z(n12329) );
  AOI22_X1 U14650 ( .A1(n12626), .A2(n12338), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12326) );
  NAND2_X1 U14651 ( .A1(n12635), .A2(n12358), .ZN(n12325) );
  OAI211_X1 U14652 ( .C1(n12362), .C2(n12341), .A(n12326), .B(n12325), .ZN(
        n12327) );
  AOI21_X1 U14653 ( .B1(n12634), .B2(n12364), .A(n12327), .ZN(n12328) );
  OAI21_X1 U14654 ( .B1(n12329), .B2(n12366), .A(n12328), .ZN(P3_U3169) );
  OAI211_X1 U14655 ( .C1(n12332), .C2(n12331), .A(n12330), .B(n12346), .ZN(
        n12336) );
  AOI22_X1 U14656 ( .A1(n12369), .A2(n12357), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12333) );
  OAI21_X1 U14657 ( .B1(n12722), .B2(n12361), .A(n12333), .ZN(n12334) );
  AOI21_X1 U14658 ( .B1(n12696), .B2(n12358), .A(n12334), .ZN(n12335) );
  OAI211_X1 U14659 ( .C1(n12780), .C2(n12354), .A(n12336), .B(n12335), .ZN(
        P3_U3173) );
  XNOR2_X1 U14660 ( .A(n12337), .B(n12646), .ZN(n12344) );
  AOI22_X1 U14661 ( .A1(n12369), .A2(n12338), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12340) );
  NAND2_X1 U14662 ( .A1(n12668), .A2(n12358), .ZN(n12339) );
  OAI211_X1 U14663 ( .C1(n12659), .C2(n12341), .A(n12340), .B(n12339), .ZN(
        n12342) );
  AOI21_X1 U14664 ( .B1(n12667), .B2(n12364), .A(n12342), .ZN(n12343) );
  OAI21_X1 U14665 ( .B1(n12344), .B2(n12366), .A(n12343), .ZN(P3_U3175) );
  OAI211_X1 U14666 ( .C1(n12349), .C2(n12348), .A(n12347), .B(n12346), .ZN(
        n12353) );
  NAND2_X1 U14667 ( .A1(n12370), .A2(n12357), .ZN(n12350) );
  NAND2_X1 U14668 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12507)
         );
  OAI211_X1 U14669 ( .C1(n12721), .C2(n12361), .A(n12350), .B(n12507), .ZN(
        n12351) );
  AOI21_X1 U14670 ( .B1(n12723), .B2(n12358), .A(n12351), .ZN(n12352) );
  OAI211_X1 U14671 ( .C1(n12856), .C2(n12354), .A(n12353), .B(n12352), .ZN(
        P3_U3178) );
  XOR2_X1 U14672 ( .A(n12356), .B(n12355), .Z(n12367) );
  NAND2_X1 U14673 ( .A1(n12600), .A2(n12357), .ZN(n12360) );
  AOI22_X1 U14674 ( .A1(n12603), .A2(n12358), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12359) );
  OAI211_X1 U14675 ( .C1(n12362), .C2(n12361), .A(n12360), .B(n12359), .ZN(
        n12363) );
  AOI21_X1 U14676 ( .B1(n12752), .B2(n12364), .A(n12363), .ZN(n12365) );
  OAI21_X1 U14677 ( .B1(n12367), .B2(n12366), .A(n12365), .ZN(P3_U3180) );
  MUX2_X1 U14678 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12368), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U14679 ( .A(n12585), .B(P3_DATAO_REG_28__SCAN_IN), .S(n12385), .Z(
        P3_U3519) );
  MUX2_X1 U14680 ( .A(n12600), .B(P3_DATAO_REG_27__SCAN_IN), .S(n12385), .Z(
        P3_U3518) );
  MUX2_X1 U14681 ( .A(n12614), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12385), .Z(
        P3_U3517) );
  MUX2_X1 U14682 ( .A(n12627), .B(P3_DATAO_REG_25__SCAN_IN), .S(n12385), .Z(
        P3_U3516) );
  MUX2_X1 U14683 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n12647), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U14684 ( .A(n12626), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12385), .Z(
        P3_U3514) );
  MUX2_X1 U14685 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12646), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U14686 ( .A(n12369), .B(P3_DATAO_REG_21__SCAN_IN), .S(n12385), .Z(
        P3_U3512) );
  MUX2_X1 U14687 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12704), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14688 ( .A(n12370), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12385), .Z(
        P3_U3510) );
  MUX2_X1 U14689 ( .A(n12703), .B(P3_DATAO_REG_18__SCAN_IN), .S(n12385), .Z(
        P3_U3509) );
  MUX2_X1 U14690 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n12371), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14691 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n12372), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14692 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n12373), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U14693 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n14285), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U14694 ( .A(n12374), .B(P3_DATAO_REG_13__SCAN_IN), .S(n12385), .Z(
        P3_U3504) );
  MUX2_X1 U14695 ( .A(n14287), .B(P3_DATAO_REG_12__SCAN_IN), .S(n12385), .Z(
        P3_U3503) );
  MUX2_X1 U14696 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n12375), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U14697 ( .A(n12376), .B(P3_DATAO_REG_10__SCAN_IN), .S(n12385), .Z(
        P3_U3501) );
  MUX2_X1 U14698 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n12377), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U14699 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12378), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U14700 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12379), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14701 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12380), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14702 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12381), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U14703 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12382), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U14704 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n12383), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U14705 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n12806), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U14706 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n12384), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U14707 ( .A(n12805), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12385), .Z(
        P3_U3491) );
  INV_X1 U14708 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n14299) );
  XNOR2_X1 U14709 ( .A(n12406), .B(n12407), .ZN(n12388) );
  AOI21_X1 U14710 ( .B1(n14299), .B2(n12388), .A(n12408), .ZN(n12405) );
  NAND2_X1 U14711 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n12390), .ZN(n12411) );
  OAI21_X1 U14712 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n12390), .A(n12411), 
        .ZN(n12403) );
  AOI21_X1 U14713 ( .B1(n14879), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n12391), 
        .ZN(n12392) );
  OAI21_X1 U14714 ( .B1(n14876), .B2(n12423), .A(n12392), .ZN(n12402) );
  INV_X1 U14715 ( .A(n12393), .ZN(n12395) );
  NOR2_X1 U14716 ( .A1(n12395), .A2(n12394), .ZN(n12397) );
  MUX2_X1 U14717 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n6446), .Z(n12424) );
  XNOR2_X1 U14718 ( .A(n12424), .B(n12423), .ZN(n12396) );
  NOR3_X1 U14719 ( .A1(n12398), .A2(n12397), .A3(n12396), .ZN(n12426) );
  INV_X1 U14720 ( .A(n12426), .ZN(n12400) );
  OAI21_X1 U14721 ( .B1(n12398), .B2(n12397), .A(n12396), .ZN(n12399) );
  AOI21_X1 U14722 ( .B1(n12400), .B2(n12399), .A(n14895), .ZN(n12401) );
  AOI211_X1 U14723 ( .C1(n12403), .C2(n6650), .A(n12402), .B(n12401), .ZN(
        n12404) );
  OAI21_X1 U14724 ( .B1(n12405), .B2(n14901), .A(n12404), .ZN(P3_U3195) );
  NOR2_X1 U14725 ( .A1(n12407), .A2(n12406), .ZN(n12409) );
  NAND2_X1 U14726 ( .A1(n12419), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12440) );
  OAI21_X1 U14727 ( .B1(P3_REG2_REG_14__SCAN_IN), .B2(n12419), .A(n12440), 
        .ZN(n12422) );
  AOI21_X1 U14728 ( .B1(n6600), .B2(n12422), .A(n12435), .ZN(n12433) );
  NAND2_X1 U14729 ( .A1(n12423), .A2(n12410), .ZN(n12412) );
  NAND2_X1 U14730 ( .A1(n12414), .A2(n12413), .ZN(n12415) );
  NAND2_X1 U14731 ( .A1(n12419), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12441) );
  AND2_X1 U14732 ( .A1(n12415), .A2(n12441), .ZN(n12420) );
  OAI21_X1 U14733 ( .B1(n12416), .B2(n12420), .A(n12438), .ZN(n12431) );
  AOI21_X1 U14734 ( .B1(n14879), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n12417), 
        .ZN(n12418) );
  OAI21_X1 U14735 ( .B1(n14876), .B2(n12419), .A(n12418), .ZN(n12430) );
  INV_X1 U14736 ( .A(n12420), .ZN(n12421) );
  MUX2_X1 U14737 ( .A(n12422), .B(n12421), .S(n6446), .Z(n12428) );
  NOR2_X1 U14738 ( .A1(n12424), .A2(n12423), .ZN(n12425) );
  OR2_X1 U14739 ( .A1(n12426), .A2(n12425), .ZN(n12427) );
  NOR3_X1 U14740 ( .A1(n12426), .A2(n12425), .A3(n12428), .ZN(n12444) );
  AOI211_X1 U14741 ( .C1(n12428), .C2(n12427), .A(n14895), .B(n12444), .ZN(
        n12429) );
  AOI211_X1 U14742 ( .C1(n6650), .C2(n12431), .A(n12430), .B(n12429), .ZN(
        n12432) );
  OAI21_X1 U14743 ( .B1(n12433), .B2(n14901), .A(n12432), .ZN(P3_U3196) );
  INV_X1 U14744 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12437) );
  XOR2_X1 U14745 ( .A(n12463), .B(n12456), .Z(n12436) );
  NOR2_X1 U14746 ( .A1(n12437), .A2(n12436), .ZN(n12457) );
  AOI21_X1 U14747 ( .B1(n12437), .B2(n12436), .A(n12457), .ZN(n12455) );
  NAND2_X1 U14748 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n12439), .ZN(n12464) );
  OAI21_X1 U14749 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n12439), .A(n12464), 
        .ZN(n12453) );
  INV_X1 U14750 ( .A(n12441), .ZN(n12442) );
  MUX2_X1 U14751 ( .A(n12434), .B(n12442), .S(n6446), .Z(n12443) );
  NOR2_X1 U14752 ( .A1(n12444), .A2(n12443), .ZN(n12470) );
  INV_X1 U14753 ( .A(n12470), .ZN(n12445) );
  XNOR2_X1 U14754 ( .A(n12445), .B(n12463), .ZN(n12447) );
  MUX2_X1 U14755 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n6446), .Z(n12446) );
  NOR2_X1 U14756 ( .A1(n12447), .A2(n12446), .ZN(n12468) );
  AOI21_X1 U14757 ( .B1(n12447), .B2(n12446), .A(n12468), .ZN(n12451) );
  INV_X1 U14758 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14225) );
  NOR2_X1 U14759 ( .A1(n14910), .A2(n14225), .ZN(n12448) );
  AOI211_X1 U14760 ( .C1(n14906), .C2(n12469), .A(n12449), .B(n12448), .ZN(
        n12450) );
  OAI21_X1 U14761 ( .B1(n12451), .B2(n14895), .A(n12450), .ZN(n12452) );
  AOI21_X1 U14762 ( .B1(n6650), .B2(n12453), .A(n12452), .ZN(n12454) );
  OAI21_X1 U14763 ( .B1(n12455), .B2(n14901), .A(n12454), .ZN(P3_U3197) );
  NOR2_X1 U14764 ( .A1(n12469), .A2(n12456), .ZN(n12458) );
  NOR2_X2 U14765 ( .A1(n12458), .A2(n12457), .ZN(n12461) );
  INV_X1 U14766 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12472) );
  NOR2_X1 U14767 ( .A1(n12478), .A2(n12472), .ZN(n12488) );
  INV_X1 U14768 ( .A(n12488), .ZN(n12459) );
  OAI21_X1 U14769 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(n12485), .A(n12459), 
        .ZN(n12460) );
  AOI21_X1 U14770 ( .B1(n12461), .B2(n12460), .A(n12489), .ZN(n12484) );
  INV_X1 U14771 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12471) );
  AOI22_X1 U14772 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12485), .B1(n12478), 
        .B2(n12471), .ZN(n12467) );
  NAND2_X1 U14773 ( .A1(n12463), .A2(n12462), .ZN(n12465) );
  NAND2_X1 U14774 ( .A1(n12465), .A2(n12464), .ZN(n12466) );
  NAND2_X1 U14775 ( .A1(n12467), .A2(n12466), .ZN(n12486) );
  OAI21_X1 U14776 ( .B1(n12467), .B2(n12466), .A(n12486), .ZN(n12482) );
  AOI21_X1 U14777 ( .B1(n12470), .B2(n12469), .A(n12468), .ZN(n12496) );
  MUX2_X1 U14778 ( .A(n12472), .B(n12471), .S(n6446), .Z(n12473) );
  NOR2_X1 U14779 ( .A1(n12473), .A2(n12478), .ZN(n12495) );
  NAND2_X1 U14780 ( .A1(n12473), .A2(n12478), .ZN(n12494) );
  INV_X1 U14781 ( .A(n12494), .ZN(n12474) );
  NOR2_X1 U14782 ( .A1(n12495), .A2(n12474), .ZN(n12475) );
  XNOR2_X1 U14783 ( .A(n12496), .B(n12475), .ZN(n12480) );
  INV_X1 U14784 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14228) );
  OAI21_X1 U14785 ( .B1(n14910), .B2(n14228), .A(n12476), .ZN(n12477) );
  AOI21_X1 U14786 ( .B1(n14906), .B2(n12478), .A(n12477), .ZN(n12479) );
  OAI21_X1 U14787 ( .B1(n12480), .B2(n14895), .A(n12479), .ZN(n12481) );
  AOI21_X1 U14788 ( .B1(n6650), .B2(n12482), .A(n12481), .ZN(n12483) );
  OAI21_X1 U14789 ( .B1(n12484), .B2(n14901), .A(n12483), .ZN(P3_U3198) );
  NAND2_X1 U14790 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12485), .ZN(n12487) );
  NAND2_X1 U14791 ( .A1(n12487), .A2(n12486), .ZN(n12505) );
  XNOR2_X1 U14792 ( .A(n12505), .B(n12501), .ZN(n12506) );
  XOR2_X1 U14793 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n12506), .Z(n12504) );
  INV_X1 U14794 ( .A(n12490), .ZN(n12491) );
  NAND2_X1 U14795 ( .A1(n12491), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n12521) );
  OAI21_X1 U14796 ( .B1(P3_REG2_REG_17__SCAN_IN), .B2(n12491), .A(n12521), 
        .ZN(n12492) );
  NAND2_X1 U14797 ( .A1(n12492), .A2(n14752), .ZN(n12503) );
  INV_X1 U14798 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14236) );
  OAI21_X1 U14799 ( .B1(n14910), .B2(n14236), .A(n12493), .ZN(n12500) );
  MUX2_X1 U14800 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n6446), .Z(n12511) );
  XNOR2_X1 U14801 ( .A(n12511), .B(n12510), .ZN(n12498) );
  OAI21_X1 U14802 ( .B1(n12496), .B2(n12495), .A(n12494), .ZN(n12497) );
  NOR2_X1 U14803 ( .A1(n12497), .A2(n12498), .ZN(n12509) );
  AOI211_X1 U14804 ( .C1(n12498), .C2(n12497), .A(n14895), .B(n12509), .ZN(
        n12499) );
  AOI211_X1 U14805 ( .C1(n14906), .C2(n12501), .A(n12500), .B(n12499), .ZN(
        n12502) );
  OAI211_X1 U14806 ( .C1(n14748), .C2(n12504), .A(n12503), .B(n12502), .ZN(
        P3_U3199) );
  XOR2_X1 U14807 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n12537), .Z(n12538) );
  XOR2_X1 U14808 ( .A(n12538), .B(n12539), .Z(n12525) );
  INV_X1 U14809 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n12508) );
  OAI21_X1 U14810 ( .B1(n14910), .B2(n12508), .A(n12507), .ZN(n12516) );
  MUX2_X1 U14811 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n6446), .Z(n12513) );
  AOI21_X1 U14812 ( .B1(n12511), .B2(n12510), .A(n12509), .ZN(n12531) );
  XNOR2_X1 U14813 ( .A(n12531), .B(n12537), .ZN(n12512) );
  NOR2_X1 U14814 ( .A1(n12512), .A2(n12513), .ZN(n12530) );
  AOI21_X1 U14815 ( .B1(n12513), .B2(n12512), .A(n12530), .ZN(n12514) );
  NOR2_X1 U14816 ( .A1(n12514), .A2(n14895), .ZN(n12515) );
  AOI211_X1 U14817 ( .C1(n14906), .C2(n12537), .A(n12516), .B(n12515), .ZN(
        n12524) );
  INV_X1 U14818 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12517) );
  OR2_X1 U14819 ( .A1(n12537), .A2(n12517), .ZN(n12526) );
  NAND2_X1 U14820 ( .A1(n12537), .A2(n12517), .ZN(n12518) );
  NAND2_X1 U14821 ( .A1(n12526), .A2(n12518), .ZN(n12519) );
  AOI21_X1 U14822 ( .B1(n12521), .B2(n12520), .A(n12519), .ZN(n12528) );
  AND3_X1 U14823 ( .A1(n12521), .A2(n12520), .A3(n12519), .ZN(n12522) );
  OAI21_X1 U14824 ( .B1(n12528), .B2(n12522), .A(n14752), .ZN(n12523) );
  OAI211_X1 U14825 ( .C1(n12525), .C2(n14748), .A(n12524), .B(n12523), .ZN(
        P3_U3200) );
  INV_X1 U14826 ( .A(n12526), .ZN(n12527) );
  NOR2_X1 U14827 ( .A1(n12528), .A2(n12527), .ZN(n12529) );
  XNOR2_X1 U14828 ( .A(n12533), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12532) );
  XNOR2_X1 U14829 ( .A(n12529), .B(n12532), .ZN(n12548) );
  AOI21_X1 U14830 ( .B1(n12531), .B2(n12537), .A(n12530), .ZN(n12536) );
  INV_X1 U14831 ( .A(n12532), .ZN(n12534) );
  XNOR2_X1 U14832 ( .A(n12533), .B(n12785), .ZN(n12540) );
  MUX2_X1 U14833 ( .A(n12534), .B(n12540), .S(n6446), .Z(n12535) );
  XNOR2_X1 U14834 ( .A(n12536), .B(n12535), .ZN(n12546) );
  INV_X1 U14835 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12789) );
  NAND2_X1 U14836 ( .A1(n14879), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12541) );
  OAI211_X1 U14837 ( .C1(n14876), .C2(n12543), .A(n12542), .B(n12541), .ZN(
        n12544) );
  AOI211_X1 U14838 ( .C1(n12546), .C2(n14871), .A(n12545), .B(n12544), .ZN(
        n12547) );
  OAI21_X1 U14839 ( .B1(n12548), .B2(n14901), .A(n12547), .ZN(P3_U3201) );
  NAND2_X1 U14840 ( .A1(n14944), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n12549) );
  OAI211_X1 U14841 ( .C1(n8926), .C2(n14294), .A(n12550), .B(n12549), .ZN(
        P3_U3203) );
  INV_X1 U14842 ( .A(n12551), .ZN(n12562) );
  OAI222_X1 U14843 ( .A1(n14919), .A2(n12555), .B1(n12552), .B2(n14303), .C1(
        n12554), .C2(n12553), .ZN(n12556) );
  NAND2_X1 U14844 ( .A1(n12556), .A2(n14942), .ZN(n12561) );
  NOR2_X1 U14845 ( .A1(n12557), .A2(n14294), .ZN(n12558) );
  AOI211_X1 U14846 ( .C1(n14944), .C2(P3_REG2_REG_29__SCAN_IN), .A(n12559), 
        .B(n12558), .ZN(n12560) );
  OAI211_X1 U14847 ( .C1(n12562), .C2(n12727), .A(n12561), .B(n12560), .ZN(
        P3_U3204) );
  NAND2_X1 U14848 ( .A1(n12563), .A2(n12575), .ZN(n12564) );
  NAND2_X1 U14849 ( .A1(n12564), .A2(n14922), .ZN(n12565) );
  OR2_X1 U14850 ( .A1(n12566), .A2(n12565), .ZN(n12571) );
  OAI22_X1 U14851 ( .A1(n12568), .A2(n14917), .B1(n12567), .B2(n14919), .ZN(
        n12569) );
  INV_X1 U14852 ( .A(n12569), .ZN(n12570) );
  INV_X1 U14853 ( .A(n12573), .ZN(n12574) );
  OR2_X1 U14854 ( .A1(n12572), .A2(n12574), .ZN(n12576) );
  XNOR2_X1 U14855 ( .A(n12576), .B(n12575), .ZN(n12746) );
  AOI22_X1 U14856 ( .A1(n12577), .A2(n14938), .B1(n14944), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n12578) );
  OAI21_X1 U14857 ( .B1(n12824), .B2(n14294), .A(n12578), .ZN(n12579) );
  AOI21_X1 U14858 ( .B1(n12746), .B2(n12739), .A(n12579), .ZN(n12580) );
  OAI21_X1 U14859 ( .B1(n6524), .B2(n14944), .A(n12580), .ZN(P3_U3205) );
  AOI21_X1 U14860 ( .B1(n7859), .B2(n12581), .A(n12572), .ZN(n12588) );
  OAI21_X1 U14861 ( .B1(n12583), .B2(n7859), .A(n12582), .ZN(n12584) );
  NAND2_X1 U14862 ( .A1(n12584), .A2(n14922), .ZN(n12587) );
  AOI22_X1 U14863 ( .A1(n12585), .A2(n14284), .B1(n14286), .B2(n12614), .ZN(
        n12586) );
  OAI211_X1 U14864 ( .C1(n12588), .C2(n14925), .A(n12587), .B(n12586), .ZN(
        n12748) );
  INV_X1 U14865 ( .A(n12748), .ZN(n12593) );
  INV_X1 U14866 ( .A(n12588), .ZN(n12749) );
  AOI22_X1 U14867 ( .A1(n12589), .A2(n14938), .B1(n14944), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12590) );
  OAI21_X1 U14868 ( .B1(n12828), .B2(n14294), .A(n12590), .ZN(n12591) );
  AOI21_X1 U14869 ( .B1(n12749), .B2(n14939), .A(n12591), .ZN(n12592) );
  OAI21_X1 U14870 ( .B1(n12593), .B2(n14944), .A(n12592), .ZN(P3_U3206) );
  NAND2_X1 U14871 ( .A1(n12595), .A2(n12594), .ZN(n12596) );
  NAND2_X1 U14872 ( .A1(n12597), .A2(n12596), .ZN(n12753) );
  XNOR2_X1 U14873 ( .A(n12598), .B(n7935), .ZN(n12599) );
  NAND2_X1 U14874 ( .A1(n12599), .A2(n14922), .ZN(n12602) );
  AOI22_X1 U14875 ( .A1(n12600), .A2(n14284), .B1(n14286), .B2(n12627), .ZN(
        n12601) );
  OAI211_X1 U14876 ( .C1(n14925), .C2(n12753), .A(n12602), .B(n12601), .ZN(
        n12754) );
  AOI22_X1 U14877 ( .A1(n12603), .A2(n14938), .B1(n14944), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n12606) );
  NAND2_X1 U14878 ( .A1(n12752), .A2(n12604), .ZN(n12605) );
  OAI211_X1 U14879 ( .C1(n12753), .C2(n12607), .A(n12606), .B(n12605), .ZN(
        n12608) );
  AOI21_X1 U14880 ( .B1(n12754), .B2(n14942), .A(n12608), .ZN(n12609) );
  INV_X1 U14881 ( .A(n12609), .ZN(P3_U3207) );
  XNOR2_X1 U14882 ( .A(n12610), .B(n12612), .ZN(n12617) );
  OAI211_X1 U14883 ( .C1(n12613), .C2(n12612), .A(n12611), .B(n14922), .ZN(
        n12616) );
  AOI22_X1 U14884 ( .A1(n12614), .A2(n14284), .B1(n12647), .B2(n14286), .ZN(
        n12615) );
  OAI211_X1 U14885 ( .C1(n14925), .C2(n12617), .A(n12616), .B(n12615), .ZN(
        n12758) );
  INV_X1 U14886 ( .A(n12758), .ZN(n12622) );
  INV_X1 U14887 ( .A(n12617), .ZN(n12759) );
  AOI22_X1 U14888 ( .A1(n12618), .A2(n14938), .B1(n14944), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n12619) );
  OAI21_X1 U14889 ( .B1(n12836), .B2(n14294), .A(n12619), .ZN(n12620) );
  AOI21_X1 U14890 ( .B1(n12759), .B2(n14939), .A(n12620), .ZN(n12621) );
  OAI21_X1 U14891 ( .B1(n12622), .B2(n14944), .A(n12621), .ZN(P3_U3208) );
  INV_X1 U14892 ( .A(n12623), .ZN(n12624) );
  AOI21_X1 U14893 ( .B1(n12629), .B2(n12625), .A(n12624), .ZN(n12633) );
  AOI22_X1 U14894 ( .A1(n12627), .A2(n14284), .B1(n14286), .B2(n12626), .ZN(
        n12632) );
  OAI211_X1 U14895 ( .C1(n12630), .C2(n12629), .A(n12628), .B(n14922), .ZN(
        n12631) );
  OAI211_X1 U14896 ( .C1(n12633), .C2(n14925), .A(n12632), .B(n12631), .ZN(
        n12762) );
  INV_X1 U14897 ( .A(n12762), .ZN(n12639) );
  INV_X1 U14898 ( .A(n12633), .ZN(n12763) );
  INV_X1 U14899 ( .A(n12634), .ZN(n12840) );
  AOI22_X1 U14900 ( .A1(n12635), .A2(n14938), .B1(n14944), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n12636) );
  OAI21_X1 U14901 ( .B1(n12840), .B2(n14294), .A(n12636), .ZN(n12637) );
  AOI21_X1 U14902 ( .B1(n12763), .B2(n14939), .A(n12637), .ZN(n12638) );
  OAI21_X1 U14903 ( .B1(n12639), .B2(n14944), .A(n12638), .ZN(P3_U3209) );
  OAI21_X1 U14904 ( .B1(n12642), .B2(n12641), .A(n12640), .ZN(n12769) );
  OAI211_X1 U14905 ( .C1(n12645), .C2(n12644), .A(n12643), .B(n14922), .ZN(
        n12649) );
  AOI22_X1 U14906 ( .A1(n12647), .A2(n14284), .B1(n14286), .B2(n12646), .ZN(
        n12648) );
  OAI211_X1 U14907 ( .C1(n14925), .C2(n12769), .A(n12649), .B(n12648), .ZN(
        n12650) );
  INV_X1 U14908 ( .A(n12650), .ZN(n12768) );
  INV_X1 U14909 ( .A(n12769), .ZN(n12655) );
  INV_X1 U14910 ( .A(n12766), .ZN(n12653) );
  AOI22_X1 U14911 ( .A1(n12651), .A2(n14938), .B1(n14944), .B2(
        P3_REG2_REG_23__SCAN_IN), .ZN(n12652) );
  OAI21_X1 U14912 ( .B1(n12653), .B2(n14294), .A(n12652), .ZN(n12654) );
  AOI21_X1 U14913 ( .B1(n12655), .B2(n14939), .A(n12654), .ZN(n12656) );
  OAI21_X1 U14914 ( .B1(n12768), .B2(n14944), .A(n12656), .ZN(P3_U3210) );
  XNOR2_X1 U14915 ( .A(n12657), .B(n12666), .ZN(n12658) );
  OAI222_X1 U14916 ( .A1(n14917), .A2(n12659), .B1(n14919), .B2(n12690), .C1(
        n14303), .C2(n12658), .ZN(n12770) );
  INV_X1 U14917 ( .A(n12770), .ZN(n12672) );
  NAND2_X1 U14918 ( .A1(n12660), .A2(n12661), .ZN(n12679) );
  NAND2_X1 U14919 ( .A1(n12679), .A2(n12662), .ZN(n12664) );
  NAND2_X1 U14920 ( .A1(n12664), .A2(n12663), .ZN(n12665) );
  XOR2_X1 U14921 ( .A(n12666), .B(n12665), .Z(n12771) );
  AOI22_X1 U14922 ( .A1(n12668), .A2(n14938), .B1(n14944), .B2(
        P3_REG2_REG_22__SCAN_IN), .ZN(n12669) );
  OAI21_X1 U14923 ( .B1(n7929), .B2(n14294), .A(n12669), .ZN(n12670) );
  AOI21_X1 U14924 ( .B1(n12771), .B2(n12739), .A(n12670), .ZN(n12671) );
  OAI21_X1 U14925 ( .B1(n12672), .B2(n14944), .A(n12671), .ZN(P3_U3211) );
  INV_X1 U14926 ( .A(n12673), .ZN(n12674) );
  AOI21_X1 U14927 ( .B1(n12680), .B2(n12675), .A(n12674), .ZN(n12676) );
  OAI222_X1 U14928 ( .A1(n14917), .A2(n12678), .B1(n14919), .B2(n12677), .C1(
        n14303), .C2(n12676), .ZN(n12774) );
  INV_X1 U14929 ( .A(n12774), .ZN(n12686) );
  XOR2_X1 U14930 ( .A(n12680), .B(n12679), .Z(n12775) );
  INV_X1 U14931 ( .A(n12681), .ZN(n12848) );
  AOI22_X1 U14932 ( .A1(n14938), .A2(n12682), .B1(n14944), .B2(
        P3_REG2_REG_21__SCAN_IN), .ZN(n12683) );
  OAI21_X1 U14933 ( .B1(n12848), .B2(n14294), .A(n12683), .ZN(n12684) );
  AOI21_X1 U14934 ( .B1(n12775), .B2(n12739), .A(n12684), .ZN(n12685) );
  OAI21_X1 U14935 ( .B1(n12686), .B2(n14944), .A(n12685), .ZN(P3_U3212) );
  XNOR2_X1 U14936 ( .A(n12688), .B(n12687), .ZN(n12689) );
  NAND2_X1 U14937 ( .A1(n12689), .A2(n14922), .ZN(n12693) );
  OAI22_X1 U14938 ( .A1(n12690), .A2(n14917), .B1(n12722), .B2(n14919), .ZN(
        n12691) );
  INV_X1 U14939 ( .A(n12691), .ZN(n12692) );
  NAND2_X1 U14940 ( .A1(n12693), .A2(n12692), .ZN(n12782) );
  NAND2_X1 U14941 ( .A1(n12695), .A2(n12694), .ZN(n12778) );
  NAND3_X1 U14942 ( .A1(n12660), .A2(n12778), .A3(n12739), .ZN(n12698) );
  AOI22_X1 U14943 ( .A1(n14944), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n14938), 
        .B2(n12696), .ZN(n12697) );
  OAI211_X1 U14944 ( .C1(n12780), .C2(n14294), .A(n12698), .B(n12697), .ZN(
        n12699) );
  AOI21_X1 U14945 ( .B1(n12782), .B2(n14942), .A(n12699), .ZN(n12700) );
  INV_X1 U14946 ( .A(n12700), .ZN(P3_U3213) );
  OAI211_X1 U14947 ( .C1(n12702), .C2(n7729), .A(n12701), .B(n14922), .ZN(
        n12706) );
  AOI22_X1 U14948 ( .A1(n12704), .A2(n14284), .B1(n14286), .B2(n12703), .ZN(
        n12705) );
  NAND2_X1 U14949 ( .A1(n12706), .A2(n12705), .ZN(n12783) );
  INV_X1 U14950 ( .A(n12783), .ZN(n12712) );
  XNOR2_X1 U14951 ( .A(n12707), .B(n7729), .ZN(n12784) );
  AOI22_X1 U14952 ( .A1(n14944), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n14938), 
        .B2(n12708), .ZN(n12709) );
  OAI21_X1 U14953 ( .B1(n12853), .B2(n14294), .A(n12709), .ZN(n12710) );
  AOI21_X1 U14954 ( .B1(n12784), .B2(n12739), .A(n12710), .ZN(n12711) );
  OAI21_X1 U14955 ( .B1(n12712), .B2(n14944), .A(n12711), .ZN(P3_U3214) );
  NAND2_X1 U14956 ( .A1(n12713), .A2(n12714), .ZN(n12715) );
  XNOR2_X1 U14957 ( .A(n12715), .B(n12719), .ZN(n12788) );
  INV_X1 U14958 ( .A(n12788), .ZN(n12728) );
  AOI21_X1 U14959 ( .B1(n12719), .B2(n12718), .A(n12717), .ZN(n12720) );
  OAI222_X1 U14960 ( .A1(n14917), .A2(n12722), .B1(n14919), .B2(n12721), .C1(
        n14303), .C2(n12720), .ZN(n12787) );
  AOI22_X1 U14961 ( .A1(n14944), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n14938), 
        .B2(n12723), .ZN(n12724) );
  OAI21_X1 U14962 ( .B1(n12856), .B2(n14294), .A(n12724), .ZN(n12725) );
  AOI21_X1 U14963 ( .B1(n12787), .B2(n14942), .A(n12725), .ZN(n12726) );
  OAI21_X1 U14964 ( .B1(n12728), .B2(n12727), .A(n12726), .ZN(P3_U3215) );
  XNOR2_X1 U14965 ( .A(n12730), .B(n12729), .ZN(n12731) );
  OAI222_X1 U14966 ( .A1(n14917), .A2(n12733), .B1(n14919), .B2(n12732), .C1(
        n12731), .C2(n14303), .ZN(n12791) );
  INV_X1 U14967 ( .A(n12791), .ZN(n12741) );
  OAI21_X1 U14968 ( .B1(n12735), .B2(n12734), .A(n12713), .ZN(n12792) );
  AOI22_X1 U14969 ( .A1(n14944), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n14938), 
        .B2(n12736), .ZN(n12737) );
  OAI21_X1 U14970 ( .B1(n12860), .B2(n14294), .A(n12737), .ZN(n12738) );
  AOI21_X1 U14971 ( .B1(n12792), .B2(n12739), .A(n12738), .ZN(n12740) );
  OAI21_X1 U14972 ( .B1(n12741), .B2(n14944), .A(n12740), .ZN(P3_U3216) );
  INV_X1 U14973 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n12743) );
  NAND2_X1 U14974 ( .A1(n12813), .A2(n7286), .ZN(n12742) );
  NAND2_X1 U14975 ( .A1(n12814), .A2(n15164), .ZN(n12744) );
  OAI211_X1 U14976 ( .C1(n15164), .C2(n12743), .A(n12742), .B(n12744), .ZN(
        P3_U3490) );
  NAND2_X1 U14977 ( .A1(n12818), .A2(n7286), .ZN(n12745) );
  OAI211_X1 U14978 ( .C1(n15164), .C2(n7902), .A(n12745), .B(n12744), .ZN(
        P3_U3489) );
  AOI21_X1 U14979 ( .B1(n14989), .B2(n12749), .A(n12748), .ZN(n12825) );
  MUX2_X1 U14980 ( .A(n12750), .B(n12825), .S(n15164), .Z(n12751) );
  OAI21_X1 U14981 ( .B1(n12828), .B2(n12803), .A(n12751), .ZN(P3_U3486) );
  INV_X1 U14982 ( .A(n12752), .ZN(n12832) );
  INV_X1 U14983 ( .A(n12753), .ZN(n12755) );
  AOI21_X1 U14984 ( .B1(n14989), .B2(n12755), .A(n12754), .ZN(n12829) );
  MUX2_X1 U14985 ( .A(n12756), .B(n12829), .S(n15164), .Z(n12757) );
  OAI21_X1 U14986 ( .B1(n12832), .B2(n12803), .A(n12757), .ZN(P3_U3485) );
  AOI21_X1 U14987 ( .B1(n14989), .B2(n12759), .A(n12758), .ZN(n12833) );
  MUX2_X1 U14988 ( .A(n12760), .B(n12833), .S(n15164), .Z(n12761) );
  OAI21_X1 U14989 ( .B1(n12836), .B2(n12803), .A(n12761), .ZN(P3_U3484) );
  AOI21_X1 U14990 ( .B1(n14989), .B2(n12763), .A(n12762), .ZN(n12837) );
  MUX2_X1 U14991 ( .A(n12764), .B(n12837), .S(n15164), .Z(n12765) );
  OAI21_X1 U14992 ( .B1(n12840), .B2(n12803), .A(n12765), .ZN(P3_U3483) );
  INV_X1 U14993 ( .A(n14989), .ZN(n14981) );
  NAND2_X1 U14994 ( .A1(n12766), .A2(n14957), .ZN(n12767) );
  OAI211_X1 U14995 ( .C1(n12769), .C2(n14981), .A(n12768), .B(n12767), .ZN(
        n12841) );
  MUX2_X1 U14996 ( .A(P3_REG1_REG_23__SCAN_IN), .B(n12841), .S(n15164), .Z(
        P3_U3482) );
  AOI21_X1 U14997 ( .B1(n14323), .B2(n12771), .A(n12770), .ZN(n12842) );
  MUX2_X1 U14998 ( .A(n12772), .B(n12842), .S(n15164), .Z(n12773) );
  OAI21_X1 U14999 ( .B1(n7929), .B2(n12803), .A(n12773), .ZN(P3_U3481) );
  INV_X1 U15000 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12776) );
  AOI21_X1 U15001 ( .B1(n14323), .B2(n12775), .A(n12774), .ZN(n12845) );
  MUX2_X1 U15002 ( .A(n12776), .B(n12845), .S(n15164), .Z(n12777) );
  OAI21_X1 U15003 ( .B1(n12848), .B2(n12803), .A(n12777), .ZN(P3_U3480) );
  NAND3_X1 U15004 ( .A1(n12660), .A2(n12778), .A3(n14323), .ZN(n12779) );
  OAI21_X1 U15005 ( .B1(n12780), .B2(n14979), .A(n12779), .ZN(n12781) );
  MUX2_X1 U15006 ( .A(n12849), .B(P3_REG1_REG_20__SCAN_IN), .S(n15162), .Z(
        P3_U3479) );
  AOI21_X1 U15007 ( .B1(n14323), .B2(n12784), .A(n12783), .ZN(n12850) );
  MUX2_X1 U15008 ( .A(n12785), .B(n12850), .S(n15164), .Z(n12786) );
  OAI21_X1 U15009 ( .B1(n12803), .B2(n12853), .A(n12786), .ZN(P3_U3478) );
  AOI21_X1 U15010 ( .B1(n14323), .B2(n12788), .A(n12787), .ZN(n12854) );
  MUX2_X1 U15011 ( .A(n12789), .B(n12854), .S(n15164), .Z(n12790) );
  OAI21_X1 U15012 ( .B1(n12856), .B2(n12803), .A(n12790), .ZN(P3_U3477) );
  INV_X1 U15013 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12793) );
  AOI21_X1 U15014 ( .B1(n14323), .B2(n12792), .A(n12791), .ZN(n12857) );
  MUX2_X1 U15015 ( .A(n12793), .B(n12857), .S(n15164), .Z(n12794) );
  OAI21_X1 U15016 ( .B1(n12860), .B2(n12803), .A(n12794), .ZN(P3_U3476) );
  AOI22_X1 U15017 ( .A1(n12796), .A2(n14323), .B1(n14957), .B2(n12795), .ZN(
        n12797) );
  NAND2_X1 U15018 ( .A1(n12798), .A2(n12797), .ZN(n12861) );
  MUX2_X1 U15019 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n12861), .S(n15164), .Z(
        P3_U3475) );
  INV_X1 U15020 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12801) );
  AOI21_X1 U15021 ( .B1(n14323), .B2(n12800), .A(n12799), .ZN(n12862) );
  MUX2_X1 U15022 ( .A(n12801), .B(n12862), .S(n15164), .Z(n12802) );
  OAI21_X1 U15023 ( .B1(n12865), .B2(n12803), .A(n12802), .ZN(P3_U3474) );
  NAND2_X1 U15024 ( .A1(n14940), .A2(n12804), .ZN(n12810) );
  AOI22_X1 U15025 ( .A1(n12806), .A2(n14284), .B1(n14286), .B2(n12805), .ZN(
        n12809) );
  NAND2_X1 U15026 ( .A1(n12807), .A2(n14922), .ZN(n12808) );
  AND3_X1 U15027 ( .A1(n12810), .A2(n12809), .A3(n12808), .ZN(n14934) );
  AND2_X1 U15028 ( .A1(n9759), .A2(n14957), .ZN(n14937) );
  AOI21_X1 U15029 ( .B1(n14940), .B2(n14989), .A(n14937), .ZN(n12811) );
  AND2_X1 U15030 ( .A1(n14934), .A2(n12811), .ZN(n14946) );
  INV_X1 U15031 ( .A(n14946), .ZN(n12812) );
  MUX2_X1 U15032 ( .A(P3_REG1_REG_1__SCAN_IN), .B(n12812), .S(n15164), .Z(
        P3_U3460) );
  INV_X1 U15033 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n12816) );
  INV_X1 U15034 ( .A(n12864), .ZN(n12817) );
  NAND2_X1 U15035 ( .A1(n12813), .A2(n12817), .ZN(n12815) );
  NAND2_X1 U15036 ( .A1(n12814), .A2(n14993), .ZN(n12819) );
  OAI211_X1 U15037 ( .C1(n12816), .C2(n14993), .A(n12815), .B(n12819), .ZN(
        P3_U3458) );
  INV_X1 U15038 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n12821) );
  NAND2_X1 U15039 ( .A1(n12818), .A2(n12817), .ZN(n12820) );
  OAI211_X1 U15040 ( .C1(n12821), .C2(n14993), .A(n12820), .B(n12819), .ZN(
        P3_U3457) );
  OAI21_X1 U15041 ( .B1(n12824), .B2(n12864), .A(n12823), .ZN(P3_U3455) );
  INV_X1 U15042 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n12826) );
  MUX2_X1 U15043 ( .A(n12826), .B(n12825), .S(n14993), .Z(n12827) );
  OAI21_X1 U15044 ( .B1(n12828), .B2(n12864), .A(n12827), .ZN(P3_U3454) );
  INV_X1 U15045 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n12830) );
  MUX2_X1 U15046 ( .A(n12830), .B(n12829), .S(n14993), .Z(n12831) );
  OAI21_X1 U15047 ( .B1(n12832), .B2(n12864), .A(n12831), .ZN(P3_U3453) );
  INV_X1 U15048 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n12834) );
  MUX2_X1 U15049 ( .A(n12834), .B(n12833), .S(n14993), .Z(n12835) );
  OAI21_X1 U15050 ( .B1(n12836), .B2(n12864), .A(n12835), .ZN(P3_U3452) );
  INV_X1 U15051 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n12838) );
  MUX2_X1 U15052 ( .A(n12838), .B(n12837), .S(n14993), .Z(n12839) );
  OAI21_X1 U15053 ( .B1(n12840), .B2(n12864), .A(n12839), .ZN(P3_U3451) );
  MUX2_X1 U15054 ( .A(P3_REG0_REG_23__SCAN_IN), .B(n12841), .S(n14993), .Z(
        P3_U3450) );
  INV_X1 U15055 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n12843) );
  MUX2_X1 U15056 ( .A(n12843), .B(n12842), .S(n14993), .Z(n12844) );
  OAI21_X1 U15057 ( .B1(n7929), .B2(n12864), .A(n12844), .ZN(P3_U3449) );
  INV_X1 U15058 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12846) );
  MUX2_X1 U15059 ( .A(n12846), .B(n12845), .S(n14993), .Z(n12847) );
  OAI21_X1 U15060 ( .B1(n12848), .B2(n12864), .A(n12847), .ZN(P3_U3448) );
  MUX2_X1 U15061 ( .A(n12849), .B(P3_REG0_REG_20__SCAN_IN), .S(n14991), .Z(
        P3_U3447) );
  INV_X1 U15062 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n12851) );
  MUX2_X1 U15063 ( .A(n12851), .B(n12850), .S(n14993), .Z(n12852) );
  OAI21_X1 U15064 ( .B1(n12864), .B2(n12853), .A(n12852), .ZN(P3_U3446) );
  INV_X1 U15065 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n15037) );
  MUX2_X1 U15066 ( .A(n15037), .B(n12854), .S(n14993), .Z(n12855) );
  OAI21_X1 U15067 ( .B1(n12856), .B2(n12864), .A(n12855), .ZN(P3_U3444) );
  INV_X1 U15068 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n12858) );
  MUX2_X1 U15069 ( .A(n12858), .B(n12857), .S(n14993), .Z(n12859) );
  OAI21_X1 U15070 ( .B1(n12860), .B2(n12864), .A(n12859), .ZN(P3_U3441) );
  MUX2_X1 U15071 ( .A(P3_REG0_REG_16__SCAN_IN), .B(n12861), .S(n14993), .Z(
        P3_U3438) );
  INV_X1 U15072 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n15112) );
  MUX2_X1 U15073 ( .A(n15112), .B(n12862), .S(n14993), .Z(n12863) );
  OAI21_X1 U15074 ( .B1(n12865), .B2(n12864), .A(n12863), .ZN(P3_U3435) );
  MUX2_X1 U15075 ( .A(P3_D_REG_1__SCAN_IN), .B(n12866), .S(n12867), .Z(
        P3_U3377) );
  MUX2_X1 U15076 ( .A(P3_D_REG_0__SCAN_IN), .B(n12868), .S(n12867), .Z(
        P3_U3376) );
  NAND3_X1 U15077 ( .A1(n12869), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .ZN(n12872) );
  OAI22_X1 U15078 ( .A1(n12873), .A2(n12872), .B1(n12871), .B2(n12870), .ZN(
        n12874) );
  AOI21_X1 U15079 ( .B1(n12876), .B2(n12875), .A(n12874), .ZN(n12877) );
  INV_X1 U15080 ( .A(n12877), .ZN(P3_U3264) );
  INV_X1 U15081 ( .A(n12878), .ZN(n12879) );
  OAI222_X1 U15082 ( .A1(n12883), .A2(n12881), .B1(P3_U3151), .B2(n12880), 
        .C1(n12886), .C2(n12879), .ZN(P3_U3267) );
  INV_X1 U15083 ( .A(n12882), .ZN(n12885) );
  OAI222_X1 U15084 ( .A1(P3_U3151), .A2(n6446), .B1(n12886), .B2(n12885), .C1(
        n12884), .C2(n12883), .ZN(P3_U3268) );
  MUX2_X1 U15085 ( .A(n12888), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  NAND2_X1 U15086 ( .A1(n12890), .A2(n12889), .ZN(n13012) );
  INV_X1 U15087 ( .A(n13012), .ZN(n12896) );
  XNOR2_X1 U15088 ( .A(n13466), .B(n12911), .ZN(n12891) );
  NAND2_X1 U15089 ( .A1(n13198), .A2(n14633), .ZN(n12892) );
  XNOR2_X1 U15090 ( .A(n12891), .B(n12892), .ZN(n13011) );
  INV_X1 U15091 ( .A(n13011), .ZN(n12895) );
  INV_X1 U15092 ( .A(n12891), .ZN(n12894) );
  INV_X1 U15093 ( .A(n12892), .ZN(n12893) );
  XNOR2_X1 U15094 ( .A(n13459), .B(n12911), .ZN(n12897) );
  NAND2_X1 U15095 ( .A1(n13202), .A2(n14633), .ZN(n12898) );
  NAND2_X1 U15096 ( .A1(n12897), .A2(n12898), .ZN(n12902) );
  INV_X1 U15097 ( .A(n12897), .ZN(n12900) );
  INV_X1 U15098 ( .A(n12898), .ZN(n12899) );
  NAND2_X1 U15099 ( .A1(n12900), .A2(n12899), .ZN(n12901) );
  AND2_X1 U15100 ( .A1(n12902), .A2(n12901), .ZN(n12946) );
  XNOR2_X1 U15101 ( .A(n13452), .B(n12911), .ZN(n12903) );
  NAND2_X1 U15102 ( .A1(n13177), .A2(n14633), .ZN(n12904) );
  NAND2_X1 U15103 ( .A1(n12903), .A2(n12904), .ZN(n12908) );
  INV_X1 U15104 ( .A(n12903), .ZN(n12906) );
  INV_X1 U15105 ( .A(n12904), .ZN(n12905) );
  NAND2_X1 U15106 ( .A1(n12906), .A2(n12905), .ZN(n12907) );
  AND2_X1 U15107 ( .A1(n12908), .A2(n12907), .ZN(n12996) );
  XNOR2_X1 U15108 ( .A(n13447), .B(n12911), .ZN(n12910) );
  NAND2_X1 U15109 ( .A1(n13208), .A2(n14633), .ZN(n12909) );
  XNOR2_X1 U15110 ( .A(n12910), .B(n12909), .ZN(n12970) );
  XNOR2_X1 U15111 ( .A(n13442), .B(n12911), .ZN(n12912) );
  AND2_X1 U15112 ( .A1(n13183), .A2(n14633), .ZN(n13002) );
  INV_X1 U15113 ( .A(n12912), .ZN(n12913) );
  AND2_X1 U15114 ( .A1(n12914), .A2(n12913), .ZN(n12915) );
  XOR2_X1 U15115 ( .A(n12960), .B(n13438), .Z(n12917) );
  XNOR2_X1 U15116 ( .A(n12916), .B(n12917), .ZN(n12937) );
  NOR2_X1 U15117 ( .A1(n13212), .A2(n13300), .ZN(n12939) );
  NOR2_X1 U15118 ( .A1(n12937), .A2(n12939), .ZN(n12938) );
  XNOR2_X1 U15119 ( .A(n13432), .B(n12960), .ZN(n12918) );
  NAND2_X1 U15120 ( .A1(n13187), .A2(n9633), .ZN(n12919) );
  XNOR2_X1 U15121 ( .A(n12918), .B(n12919), .ZN(n12986) );
  INV_X1 U15122 ( .A(n12919), .ZN(n12920) );
  XNOR2_X1 U15123 ( .A(n13304), .B(n12960), .ZN(n12924) );
  NAND2_X1 U15124 ( .A1(n13190), .A2(n14633), .ZN(n12922) );
  XNOR2_X1 U15125 ( .A(n12924), .B(n12922), .ZN(n12976) );
  INV_X1 U15126 ( .A(n12922), .ZN(n12923) );
  AND2_X1 U15127 ( .A1(n13193), .A2(n14633), .ZN(n12926) );
  XNOR2_X1 U15128 ( .A(n13420), .B(n12960), .ZN(n12925) );
  NOR2_X1 U15129 ( .A1(n12925), .A2(n12926), .ZN(n12927) );
  AOI21_X1 U15130 ( .B1(n12926), .B2(n12925), .A(n12927), .ZN(n13032) );
  INV_X1 U15131 ( .A(n12927), .ZN(n12928) );
  NAND2_X1 U15132 ( .A1(n13222), .A2(n14633), .ZN(n12956) );
  XNOR2_X1 U15133 ( .A(n13265), .B(n12960), .ZN(n12955) );
  XOR2_X1 U15134 ( .A(n12956), .B(n12955), .Z(n12958) );
  XNOR2_X1 U15135 ( .A(n12959), .B(n12958), .ZN(n12936) );
  NAND2_X1 U15136 ( .A1(n13224), .A2(n12987), .ZN(n12930) );
  NAND2_X1 U15137 ( .A1(n13193), .A2(n13004), .ZN(n12929) );
  NAND2_X1 U15138 ( .A1(n12930), .A2(n12929), .ZN(n13262) );
  NAND2_X1 U15139 ( .A1(n13268), .A2(n13025), .ZN(n12931) );
  OAI21_X1 U15140 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n12932), .A(n12931), .ZN(
        n12933) );
  AOI21_X1 U15141 ( .B1(n13262), .B2(n13040), .A(n12933), .ZN(n12935) );
  NAND2_X1 U15142 ( .A1(n13265), .A2(n13026), .ZN(n12934) );
  OAI211_X1 U15143 ( .C1(n12936), .C2(n13018), .A(n12935), .B(n12934), .ZN(
        P2_U3186) );
  AOI21_X1 U15144 ( .B1(n12939), .B2(n12937), .A(n12938), .ZN(n12944) );
  AOI22_X1 U15145 ( .A1(n13187), .A2(n13164), .B1(n13004), .B2(n13183), .ZN(
        n13328) );
  OAI22_X1 U15146 ( .A1(n13328), .A2(n13015), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12940), .ZN(n12941) );
  AOI21_X1 U15147 ( .B1(n13334), .B2(n13025), .A(n12941), .ZN(n12943) );
  NAND2_X1 U15148 ( .A1(n13438), .A2(n13026), .ZN(n12942) );
  OAI211_X1 U15149 ( .C1(n12944), .C2(n13018), .A(n12943), .B(n12942), .ZN(
        P2_U3188) );
  INV_X1 U15150 ( .A(n13459), .ZN(n13388) );
  OAI21_X1 U15151 ( .B1(n12947), .B2(n12946), .A(n6623), .ZN(n12948) );
  NAND2_X1 U15152 ( .A1(n12948), .A2(n13034), .ZN(n12954) );
  INV_X1 U15153 ( .A(n12949), .ZN(n13386) );
  NAND2_X1 U15154 ( .A1(n13177), .A2(n12987), .ZN(n12951) );
  NAND2_X1 U15155 ( .A1(n13198), .A2(n13004), .ZN(n12950) );
  AND2_X1 U15156 ( .A1(n12951), .A2(n12950), .ZN(n13456) );
  NAND2_X1 U15157 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13157)
         );
  OAI21_X1 U15158 ( .B1(n13015), .B2(n13456), .A(n13157), .ZN(n12952) );
  AOI21_X1 U15159 ( .B1(n13386), .B2(n13025), .A(n12952), .ZN(n12953) );
  OAI211_X1 U15160 ( .C1(n13388), .C2(n13043), .A(n12954), .B(n12953), .ZN(
        P2_U3191) );
  INV_X1 U15161 ( .A(n12955), .ZN(n12957) );
  NAND2_X1 U15162 ( .A1(n13224), .A2(n14633), .ZN(n12961) );
  XNOR2_X1 U15163 ( .A(n12961), .B(n12960), .ZN(n12962) );
  XNOR2_X1 U15164 ( .A(n13410), .B(n12962), .ZN(n12963) );
  NAND2_X1 U15165 ( .A1(n13046), .A2(n12987), .ZN(n12965) );
  NAND2_X1 U15166 ( .A1(n13222), .A2(n13004), .ZN(n12964) );
  AND2_X1 U15167 ( .A1(n12965), .A2(n12964), .ZN(n13244) );
  INV_X1 U15168 ( .A(n13250), .ZN(n12966) );
  AOI22_X1 U15169 ( .A1(n12966), .A2(n13025), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12967) );
  OAI21_X1 U15170 ( .B1(n13244), .B2(n13015), .A(n12967), .ZN(n12968) );
  AOI21_X1 U15171 ( .B1(n13410), .B2(n13026), .A(n12968), .ZN(n12969) );
  XNOR2_X1 U15172 ( .A(n12971), .B(n12970), .ZN(n12975) );
  INV_X1 U15173 ( .A(n13183), .ZN(n13211) );
  INV_X1 U15174 ( .A(n13177), .ZN(n13205) );
  OAI22_X1 U15175 ( .A1(n13211), .A2(n13036), .B1(n13205), .B2(n13228), .ZN(
        n13355) );
  AOI22_X1 U15176 ( .A1(n13355), .A2(n13040), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12972) );
  OAI21_X1 U15177 ( .B1(n13359), .B2(n13038), .A(n12972), .ZN(n12973) );
  AOI21_X1 U15178 ( .B1(n13447), .B2(n13026), .A(n12973), .ZN(n12974) );
  OAI21_X1 U15179 ( .B1(n12975), .B2(n13018), .A(n12974), .ZN(P2_U3195) );
  XNOR2_X1 U15180 ( .A(n12977), .B(n12976), .ZN(n12983) );
  NAND2_X1 U15181 ( .A1(n13193), .A2(n12987), .ZN(n12979) );
  NAND2_X1 U15182 ( .A1(n13187), .A2(n13004), .ZN(n12978) );
  NAND2_X1 U15183 ( .A1(n12979), .A2(n12978), .ZN(n13292) );
  AOI22_X1 U15184 ( .A1(n13292), .A2(n13040), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12980) );
  OAI21_X1 U15185 ( .B1(n13301), .B2(n13038), .A(n12980), .ZN(n12981) );
  AOI21_X1 U15186 ( .B1(n13304), .B2(n13026), .A(n12981), .ZN(n12982) );
  OAI21_X1 U15187 ( .B1(n12983), .B2(n13018), .A(n12982), .ZN(P2_U3197) );
  INV_X1 U15188 ( .A(n13432), .ZN(n13321) );
  OAI211_X1 U15189 ( .C1(n12984), .C2(n12986), .A(n12985), .B(n13034), .ZN(
        n12993) );
  NAND2_X1 U15190 ( .A1(n13190), .A2(n12987), .ZN(n12989) );
  OR2_X1 U15191 ( .A1(n13212), .A2(n13228), .ZN(n12988) );
  AND2_X1 U15192 ( .A1(n12989), .A2(n12988), .ZN(n13316) );
  OAI22_X1 U15193 ( .A1(n13316), .A2(n13015), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12990), .ZN(n12991) );
  AOI21_X1 U15194 ( .B1(n13319), .B2(n13025), .A(n12991), .ZN(n12992) );
  OAI211_X1 U15195 ( .C1(n13321), .C2(n13043), .A(n12993), .B(n12992), .ZN(
        P2_U3201) );
  INV_X1 U15196 ( .A(n13452), .ZN(n13377) );
  OAI21_X1 U15197 ( .B1(n12996), .B2(n12995), .A(n12994), .ZN(n12997) );
  NAND2_X1 U15198 ( .A1(n12997), .A2(n13034), .ZN(n13001) );
  INV_X1 U15199 ( .A(n12998), .ZN(n13375) );
  AOI22_X1 U15200 ( .A1(n13208), .A2(n13164), .B1(n13004), .B2(n13202), .ZN(
        n13369) );
  OAI22_X1 U15201 ( .A1(n13015), .A2(n13369), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15055), .ZN(n12999) );
  AOI21_X1 U15202 ( .B1(n13375), .B2(n13025), .A(n12999), .ZN(n13000) );
  OAI211_X1 U15203 ( .C1(n13377), .C2(n13043), .A(n13001), .B(n13000), .ZN(
        P2_U3205) );
  XNOR2_X1 U15204 ( .A(n13003), .B(n13002), .ZN(n13010) );
  OR2_X1 U15205 ( .A1(n13212), .A2(n13036), .ZN(n13006) );
  NAND2_X1 U15206 ( .A1(n13208), .A2(n13004), .ZN(n13005) );
  NAND2_X1 U15207 ( .A1(n13006), .A2(n13005), .ZN(n13340) );
  AOI22_X1 U15208 ( .A1(n13340), .A2(n13040), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13007) );
  OAI21_X1 U15209 ( .B1(n13343), .B2(n13038), .A(n13007), .ZN(n13008) );
  AOI21_X1 U15210 ( .B1(n13442), .B2(n13026), .A(n13008), .ZN(n13009) );
  OAI21_X1 U15211 ( .B1(n13010), .B2(n13018), .A(n13009), .ZN(P2_U3207) );
  XNOR2_X1 U15212 ( .A(n13012), .B(n13011), .ZN(n13019) );
  NAND2_X1 U15213 ( .A1(n13025), .A2(n13013), .ZN(n13014) );
  NAND2_X1 U15214 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n14603)
         );
  OAI211_X1 U15215 ( .C1(n13463), .C2(n13015), .A(n13014), .B(n14603), .ZN(
        n13016) );
  AOI21_X1 U15216 ( .B1(n13466), .B2(n13026), .A(n13016), .ZN(n13017) );
  OAI21_X1 U15217 ( .B1(n13019), .B2(n13018), .A(n13017), .ZN(P2_U3210) );
  XOR2_X1 U15218 ( .A(n13021), .B(n13020), .Z(n13022) );
  NAND2_X1 U15219 ( .A1(n13022), .A2(n13034), .ZN(n13030) );
  AND2_X1 U15220 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n13119) );
  AOI21_X1 U15221 ( .B1(n13040), .B2(n13023), .A(n13119), .ZN(n13029) );
  NAND2_X1 U15222 ( .A1(n13025), .A2(n13024), .ZN(n13028) );
  NAND2_X1 U15223 ( .A1(n13026), .A2(n14702), .ZN(n13027) );
  NAND4_X1 U15224 ( .A1(n13030), .A2(n13029), .A3(n13028), .A4(n13027), .ZN(
        P2_U3211) );
  OAI21_X1 U15225 ( .B1(n13033), .B2(n13032), .A(n13031), .ZN(n13035) );
  NAND2_X1 U15226 ( .A1(n13035), .A2(n13034), .ZN(n13042) );
  OAI22_X1 U15227 ( .A1(n13195), .A2(n13036), .B1(n13218), .B2(n13228), .ZN(
        n13277) );
  OAI22_X1 U15228 ( .A1(n13038), .A2(n13281), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13037), .ZN(n13039) );
  AOI21_X1 U15229 ( .B1(n13277), .B2(n13040), .A(n13039), .ZN(n13041) );
  OAI211_X1 U15230 ( .C1(n13284), .C2(n13043), .A(n13042), .B(n13041), .ZN(
        P2_U3212) );
  MUX2_X1 U15231 ( .A(n13044), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13065), .Z(
        P2_U3562) );
  MUX2_X1 U15232 ( .A(n13045), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13065), .Z(
        P2_U3561) );
  MUX2_X1 U15233 ( .A(n13046), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13065), .Z(
        P2_U3560) );
  MUX2_X1 U15234 ( .A(n13224), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13065), .Z(
        P2_U3559) );
  MUX2_X1 U15235 ( .A(n13222), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13065), .Z(
        P2_U3558) );
  MUX2_X1 U15236 ( .A(n13193), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13065), .Z(
        P2_U3557) );
  MUX2_X1 U15237 ( .A(n13190), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13065), .Z(
        P2_U3556) );
  MUX2_X1 U15238 ( .A(n13187), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13065), .Z(
        P2_U3555) );
  MUX2_X1 U15239 ( .A(n13047), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13065), .Z(
        P2_U3554) );
  MUX2_X1 U15240 ( .A(n13183), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13065), .Z(
        P2_U3553) );
  MUX2_X1 U15241 ( .A(n13208), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13065), .Z(
        P2_U3552) );
  MUX2_X1 U15242 ( .A(n13177), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13065), .Z(
        P2_U3551) );
  MUX2_X1 U15243 ( .A(n13202), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13065), .Z(
        P2_U3550) );
  MUX2_X1 U15244 ( .A(n13198), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13065), .Z(
        P2_U3549) );
  INV_X2 U15245 ( .A(P2_U3947), .ZN(n13065) );
  MUX2_X1 U15246 ( .A(n13048), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13065), .Z(
        P2_U3548) );
  MUX2_X1 U15247 ( .A(n13049), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13065), .Z(
        P2_U3547) );
  MUX2_X1 U15248 ( .A(n13050), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13065), .Z(
        P2_U3546) );
  MUX2_X1 U15249 ( .A(n13051), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13065), .Z(
        P2_U3545) );
  MUX2_X1 U15250 ( .A(n13052), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13065), .Z(
        P2_U3544) );
  MUX2_X1 U15251 ( .A(n13053), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13065), .Z(
        P2_U3543) );
  MUX2_X1 U15252 ( .A(n13054), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13065), .Z(
        P2_U3542) );
  MUX2_X1 U15253 ( .A(n13055), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13065), .Z(
        P2_U3541) );
  MUX2_X1 U15254 ( .A(n13056), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13065), .Z(
        P2_U3540) );
  MUX2_X1 U15255 ( .A(n13057), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13065), .Z(
        P2_U3539) );
  MUX2_X1 U15256 ( .A(n13058), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13065), .Z(
        P2_U3538) );
  MUX2_X1 U15257 ( .A(n13059), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13065), .Z(
        P2_U3537) );
  MUX2_X1 U15258 ( .A(n13060), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13065), .Z(
        P2_U3536) );
  MUX2_X1 U15259 ( .A(n13061), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13065), .Z(
        P2_U3535) );
  MUX2_X1 U15260 ( .A(n13062), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13065), .Z(
        P2_U3534) );
  MUX2_X1 U15261 ( .A(n13063), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13065), .Z(
        P2_U3533) );
  MUX2_X1 U15262 ( .A(n13064), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13065), .Z(
        P2_U3532) );
  MUX2_X1 U15263 ( .A(n13066), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13065), .Z(
        P2_U3531) );
  OAI211_X1 U15264 ( .C1(n13069), .C2(n13068), .A(n14586), .B(n13067), .ZN(
        n13079) );
  NAND2_X1 U15265 ( .A1(n14594), .A2(n13070), .ZN(n13078) );
  INV_X1 U15266 ( .A(n13071), .ZN(n13087) );
  NAND3_X1 U15267 ( .A1(n13073), .A2(n14565), .A3(n13072), .ZN(n13074) );
  NAND3_X1 U15268 ( .A1(n14579), .A2(n13087), .A3(n13074), .ZN(n13077) );
  NOR2_X1 U15269 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9386), .ZN(n13075) );
  AOI21_X1 U15270 ( .B1(n14610), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n13075), .ZN(
        n13076) );
  NAND4_X1 U15271 ( .A1(n13079), .A2(n13078), .A3(n13077), .A4(n13076), .ZN(
        P2_U3217) );
  OAI211_X1 U15272 ( .C1(n13082), .C2(n13081), .A(n14586), .B(n13080), .ZN(
        n13093) );
  NAND2_X1 U15273 ( .A1(n14594), .A2(n13084), .ZN(n13092) );
  INV_X1 U15274 ( .A(n13083), .ZN(n13086) );
  MUX2_X1 U15275 ( .A(n10202), .B(P2_REG2_REG_4__SCAN_IN), .S(n13084), .Z(
        n13085) );
  NAND3_X1 U15276 ( .A1(n13087), .A2(n13086), .A3(n13085), .ZN(n13088) );
  NAND3_X1 U15277 ( .A1(n14579), .A2(n13101), .A3(n13088), .ZN(n13091) );
  AOI21_X1 U15278 ( .B1(n14610), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n13089), .ZN(
        n13090) );
  NAND4_X1 U15279 ( .A1(n13093), .A2(n13092), .A3(n13091), .A4(n13090), .ZN(
        P2_U3218) );
  OAI211_X1 U15280 ( .C1(n13096), .C2(n13095), .A(n14586), .B(n13094), .ZN(
        n13107) );
  NAND2_X1 U15281 ( .A1(n14594), .A2(n13097), .ZN(n13106) );
  INV_X1 U15282 ( .A(n13098), .ZN(n13116) );
  NAND3_X1 U15283 ( .A1(n13101), .A2(n13100), .A3(n13099), .ZN(n13102) );
  NAND3_X1 U15284 ( .A1(n14579), .A2(n13116), .A3(n13102), .ZN(n13105) );
  AOI21_X1 U15285 ( .B1(n14610), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n13103), .ZN(
        n13104) );
  NAND4_X1 U15286 ( .A1(n13107), .A2(n13106), .A3(n13105), .A4(n13104), .ZN(
        P2_U3219) );
  OAI211_X1 U15287 ( .C1(n13110), .C2(n13109), .A(n14586), .B(n13108), .ZN(
        n13123) );
  NAND2_X1 U15288 ( .A1(n14594), .A2(n13112), .ZN(n13122) );
  INV_X1 U15289 ( .A(n13111), .ZN(n13115) );
  MUX2_X1 U15290 ( .A(n13113), .B(P2_REG2_REG_6__SCAN_IN), .S(n13112), .Z(
        n13114) );
  NAND3_X1 U15291 ( .A1(n13116), .A2(n13115), .A3(n13114), .ZN(n13117) );
  NAND3_X1 U15292 ( .A1(n14579), .A2(n13118), .A3(n13117), .ZN(n13121) );
  AOI21_X1 U15293 ( .B1(n14610), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n13119), .ZN(
        n13120) );
  NAND4_X1 U15294 ( .A1(n13123), .A2(n13122), .A3(n13121), .A4(n13120), .ZN(
        P2_U3220) );
  NOR2_X1 U15295 ( .A1(n13125), .A2(n13124), .ZN(n13127) );
  OAI21_X1 U15296 ( .B1(n13127), .B2(n13126), .A(n14579), .ZN(n13136) );
  AOI21_X1 U15297 ( .B1(n14610), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n13128), 
        .ZN(n13135) );
  OAI211_X1 U15298 ( .C1(n13131), .C2(n13130), .A(n13129), .B(n14586), .ZN(
        n13134) );
  NAND2_X1 U15299 ( .A1(n14594), .A2(n13132), .ZN(n13133) );
  NAND4_X1 U15300 ( .A1(n13136), .A2(n13135), .A3(n13134), .A4(n13133), .ZN(
        P2_U3225) );
  AOI21_X1 U15301 ( .B1(n13138), .B2(P2_REG1_REG_17__SCAN_IN), .A(n13137), 
        .ZN(n13139) );
  XNOR2_X1 U15302 ( .A(n14617), .B(n13139), .ZN(n14607) );
  NOR2_X1 U15303 ( .A1(n14606), .A2(n14607), .ZN(n14605) );
  NOR2_X1 U15304 ( .A1(n13139), .A2(n14617), .ZN(n13140) );
  NOR2_X1 U15305 ( .A1(n14605), .A2(n13140), .ZN(n13142) );
  INV_X1 U15306 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n13141) );
  XOR2_X1 U15307 ( .A(n13142), .B(n13141), .Z(n13153) );
  INV_X1 U15308 ( .A(n13153), .ZN(n13151) );
  OAI21_X1 U15309 ( .B1(n13145), .B2(n13144), .A(n13143), .ZN(n13146) );
  XNOR2_X1 U15310 ( .A(n13147), .B(n13146), .ZN(n14612) );
  NOR2_X1 U15311 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n14612), .ZN(n14611) );
  NOR2_X1 U15312 ( .A1(n13147), .A2(n13146), .ZN(n13148) );
  NOR2_X1 U15313 ( .A1(n14611), .A2(n13148), .ZN(n13149) );
  XOR2_X1 U15314 ( .A(n13149), .B(P2_REG2_REG_19__SCAN_IN), .Z(n13152) );
  OAI21_X1 U15315 ( .B1(n13152), .B2(n14614), .A(n14618), .ZN(n13150) );
  AOI21_X1 U15316 ( .B1(n13151), .B2(n14586), .A(n13150), .ZN(n13156) );
  AOI22_X1 U15317 ( .A1(n13153), .A2(n14586), .B1(n14579), .B2(n13152), .ZN(
        n13155) );
  MUX2_X1 U15318 ( .A(n13156), .B(n13155), .S(n13154), .Z(n13158) );
  OAI211_X1 U15319 ( .C1(n7384), .C2(n14602), .A(n13158), .B(n13157), .ZN(
        P2_U3233) );
  NOR2_X2 U15320 ( .A1(n13385), .A2(n13459), .ZN(n13372) );
  OR2_X2 U15321 ( .A1(n13447), .A2(n13373), .ZN(n13357) );
  INV_X1 U15322 ( .A(n13304), .ZN(n13427) );
  NAND2_X1 U15323 ( .A1(n13318), .A2(n13427), .ZN(n13299) );
  OR2_X2 U15324 ( .A1(n13299), .A2(n13420), .ZN(n13279) );
  NOR2_X2 U15325 ( .A1(n13279), .A2(n13265), .ZN(n13252) );
  NOR2_X2 U15326 ( .A1(n13253), .A2(n13235), .ZN(n13234) );
  NAND2_X1 U15327 ( .A1(n13234), .A2(n13401), .ZN(n13169) );
  INV_X1 U15328 ( .A(n13525), .ZN(n13162) );
  NAND2_X1 U15329 ( .A1(n13162), .A2(P2_B_REG_SCAN_IN), .ZN(n13163) );
  NAND2_X1 U15330 ( .A1(n13164), .A2(n13163), .ZN(n13229) );
  OR2_X1 U15331 ( .A1(n13165), .A2(n13229), .ZN(n13399) );
  NOR2_X1 U15332 ( .A1(n14653), .A2(n13399), .ZN(n13171) );
  NOR2_X1 U15333 ( .A1(n13160), .A2(n14625), .ZN(n13167) );
  AOI211_X1 U15334 ( .C1(n14653), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13171), 
        .B(n13167), .ZN(n13168) );
  OAI21_X1 U15335 ( .B1(n13398), .B2(n13307), .A(n13168), .ZN(P2_U3234) );
  OAI211_X1 U15336 ( .C1(n13234), .C2(n13401), .A(n13300), .B(n13169), .ZN(
        n13400) );
  NOR2_X1 U15337 ( .A1(n13401), .A2(n14625), .ZN(n13170) );
  AOI211_X1 U15338 ( .C1(n14653), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13171), 
        .B(n13170), .ZN(n13172) );
  OAI21_X1 U15339 ( .B1(n13307), .B2(n13400), .A(n13172), .ZN(P2_U3235) );
  OR2_X1 U15340 ( .A1(n13466), .A2(n13198), .ZN(n13173) );
  NAND2_X1 U15341 ( .A1(n13452), .A2(n13177), .ZN(n13178) );
  INV_X1 U15342 ( .A(n13180), .ZN(n13181) );
  NAND2_X1 U15343 ( .A1(n13442), .A2(n13183), .ZN(n13184) );
  NAND2_X1 U15344 ( .A1(n13432), .A2(n13187), .ZN(n13188) );
  OR2_X1 U15345 ( .A1(n13304), .A2(n13190), .ZN(n13191) );
  NAND2_X1 U15346 ( .A1(n13420), .A2(n13193), .ZN(n13192) );
  OR2_X1 U15347 ( .A1(n13420), .A2(n13193), .ZN(n13194) );
  INV_X1 U15348 ( .A(n13198), .ZN(n13199) );
  AND2_X1 U15349 ( .A1(n13466), .A2(n13199), .ZN(n13200) );
  INV_X1 U15350 ( .A(n13202), .ZN(n13203) );
  NAND2_X1 U15351 ( .A1(n13459), .A2(n13203), .ZN(n13204) );
  NAND2_X1 U15352 ( .A1(n13368), .A2(n13378), .ZN(n13207) );
  NAND2_X1 U15353 ( .A1(n13452), .A2(n13205), .ZN(n13206) );
  INV_X1 U15354 ( .A(n13208), .ZN(n13209) );
  AND2_X1 U15355 ( .A1(n13447), .A2(n13209), .ZN(n13210) );
  NOR2_X1 U15356 ( .A1(n13438), .A2(n13212), .ZN(n13214) );
  NAND2_X1 U15357 ( .A1(n13438), .A2(n13212), .ZN(n13213) );
  INV_X1 U15358 ( .A(n13312), .ZN(n13313) );
  NAND2_X1 U15359 ( .A1(n13314), .A2(n13313), .ZN(n13217) );
  NAND2_X1 U15360 ( .A1(n13432), .A2(n13215), .ZN(n13216) );
  AND2_X1 U15361 ( .A1(n13420), .A2(n13220), .ZN(n13221) );
  NOR2_X1 U15362 ( .A1(n13230), .A2(n13229), .ZN(n13231) );
  NAND2_X1 U15363 ( .A1(n13405), .A2(n13330), .ZN(n13241) );
  AOI211_X1 U15364 ( .C1(n13235), .C2(n13253), .A(n14633), .B(n13234), .ZN(
        n13402) );
  INV_X1 U15365 ( .A(n13236), .ZN(n13237) );
  AOI22_X1 U15366 ( .A1(n13237), .A2(n14621), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n14653), .ZN(n13238) );
  OAI21_X1 U15367 ( .B1(n13403), .B2(n14625), .A(n13238), .ZN(n13239) );
  AOI21_X1 U15368 ( .B1(n13402), .B2(n13395), .A(n13239), .ZN(n13240) );
  OAI211_X1 U15369 ( .C1(n13407), .C2(n13397), .A(n13241), .B(n13240), .ZN(
        P2_U3236) );
  OAI21_X1 U15370 ( .B1(n13243), .B2(n13242), .A(n13391), .ZN(n13245) );
  OAI21_X1 U15371 ( .B1(n13248), .B2(n13247), .A(n13246), .ZN(n13411) );
  OAI22_X1 U15372 ( .A1(n13250), .A2(n14646), .B1(n13249), .B2(n13330), .ZN(
        n13251) );
  AOI21_X1 U15373 ( .B1(n13410), .B2(n13303), .A(n13251), .ZN(n13256) );
  AOI21_X1 U15374 ( .B1(n13410), .B2(n13266), .A(n14633), .ZN(n13254) );
  AND2_X1 U15375 ( .A1(n13254), .A2(n13253), .ZN(n13409) );
  NAND2_X1 U15376 ( .A1(n13409), .A2(n13395), .ZN(n13255) );
  OAI211_X1 U15377 ( .C1(n13411), .C2(n13397), .A(n13256), .B(n13255), .ZN(
        n13257) );
  AOI21_X1 U15378 ( .B1(n13408), .B2(n13330), .A(n13257), .ZN(n13258) );
  INV_X1 U15379 ( .A(n13258), .ZN(P2_U3237) );
  XNOR2_X1 U15380 ( .A(n13260), .B(n13259), .ZN(n13261) );
  NAND2_X1 U15381 ( .A1(n13261), .A2(n13391), .ZN(n13264) );
  INV_X1 U15382 ( .A(n13262), .ZN(n13263) );
  NAND2_X1 U15383 ( .A1(n13264), .A2(n13263), .ZN(n13418) );
  INV_X1 U15384 ( .A(n13418), .ZN(n13275) );
  AOI21_X1 U15385 ( .B1(n13265), .B2(n13279), .A(n14633), .ZN(n13267) );
  NAND2_X1 U15386 ( .A1(n13267), .A2(n13266), .ZN(n13414) );
  INV_X1 U15387 ( .A(n13414), .ZN(n13271) );
  AOI22_X1 U15388 ( .A1(n13268), .A2(n14621), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n14653), .ZN(n13269) );
  OAI21_X1 U15389 ( .B1(n13416), .B2(n14625), .A(n13269), .ZN(n13270) );
  AOI21_X1 U15390 ( .B1(n13271), .B2(n13395), .A(n13270), .ZN(n13274) );
  NAND2_X1 U15391 ( .A1(n13272), .A2(n7128), .ZN(n13412) );
  NAND3_X1 U15392 ( .A1(n13413), .A2(n13412), .A3(n14628), .ZN(n13273) );
  OAI211_X1 U15393 ( .C1(n13275), .C2(n14653), .A(n13274), .B(n13273), .ZN(
        P2_U3238) );
  XNOR2_X1 U15394 ( .A(n13276), .B(n13285), .ZN(n13278) );
  AOI21_X1 U15395 ( .B1(n13278), .B2(n13391), .A(n13277), .ZN(n13422) );
  INV_X1 U15396 ( .A(n13279), .ZN(n13280) );
  AOI211_X1 U15397 ( .C1(n13420), .C2(n13299), .A(n14633), .B(n13280), .ZN(
        n13419) );
  INV_X1 U15398 ( .A(n13281), .ZN(n13282) );
  AOI22_X1 U15399 ( .A1(n13282), .A2(n14621), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n14653), .ZN(n13283) );
  OAI21_X1 U15400 ( .B1(n13284), .B2(n14625), .A(n13283), .ZN(n13288) );
  XNOR2_X1 U15401 ( .A(n13286), .B(n13285), .ZN(n13423) );
  NOR2_X1 U15402 ( .A1(n13423), .A2(n13397), .ZN(n13287) );
  AOI211_X1 U15403 ( .C1(n13419), .C2(n13395), .A(n13288), .B(n13287), .ZN(
        n13289) );
  OAI21_X1 U15404 ( .B1(n14653), .B2(n13422), .A(n13289), .ZN(P2_U3239) );
  XNOR2_X1 U15405 ( .A(n13290), .B(n13295), .ZN(n13291) );
  NAND2_X1 U15406 ( .A1(n13291), .A2(n13391), .ZN(n13294) );
  INV_X1 U15407 ( .A(n13292), .ZN(n13293) );
  NAND2_X1 U15408 ( .A1(n13294), .A2(n13293), .ZN(n13429) );
  INV_X1 U15409 ( .A(n13429), .ZN(n13310) );
  NAND2_X1 U15410 ( .A1(n13296), .A2(n13295), .ZN(n13297) );
  NAND2_X1 U15411 ( .A1(n13298), .A2(n13297), .ZN(n13424) );
  OAI211_X1 U15412 ( .C1(n13318), .C2(n13427), .A(n13300), .B(n13299), .ZN(
        n13425) );
  INV_X1 U15413 ( .A(n13301), .ZN(n13302) );
  AOI22_X1 U15414 ( .A1(P2_REG2_REG_25__SCAN_IN), .A2(n14653), .B1(n13302), 
        .B2(n14621), .ZN(n13306) );
  NAND2_X1 U15415 ( .A1(n13304), .A2(n13303), .ZN(n13305) );
  OAI211_X1 U15416 ( .C1(n13425), .C2(n13307), .A(n13306), .B(n13305), .ZN(
        n13308) );
  AOI21_X1 U15417 ( .B1(n13424), .B2(n14628), .A(n13308), .ZN(n13309) );
  OAI21_X1 U15418 ( .B1(n13310), .B2(n14653), .A(n13309), .ZN(P2_U3240) );
  XNOR2_X1 U15419 ( .A(n13311), .B(n13312), .ZN(n13435) );
  XNOR2_X1 U15420 ( .A(n13314), .B(n13313), .ZN(n13315) );
  NAND2_X1 U15421 ( .A1(n13315), .A2(n13391), .ZN(n13433) );
  INV_X1 U15422 ( .A(n13433), .ZN(n13317) );
  INV_X1 U15423 ( .A(n13316), .ZN(n13431) );
  OAI21_X1 U15424 ( .B1(n13317), .B2(n13431), .A(n13330), .ZN(n13324) );
  AOI211_X1 U15425 ( .C1(n13432), .C2(n13332), .A(n14633), .B(n13318), .ZN(
        n13430) );
  AOI22_X1 U15426 ( .A1(n14653), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n13319), 
        .B2(n14621), .ZN(n13320) );
  OAI21_X1 U15427 ( .B1(n13321), .B2(n14625), .A(n13320), .ZN(n13322) );
  AOI21_X1 U15428 ( .B1(n13430), .B2(n13395), .A(n13322), .ZN(n13323) );
  OAI211_X1 U15429 ( .C1(n13435), .C2(n13397), .A(n13324), .B(n13323), .ZN(
        P2_U3241) );
  XOR2_X1 U15430 ( .A(n13325), .B(n13326), .Z(n13440) );
  XNOR2_X1 U15431 ( .A(n13327), .B(n13326), .ZN(n13329) );
  OAI21_X1 U15432 ( .B1(n13329), .B2(n14640), .A(n13328), .ZN(n13436) );
  NAND2_X1 U15433 ( .A1(n13436), .A2(n13330), .ZN(n13338) );
  INV_X1 U15434 ( .A(n13332), .ZN(n13333) );
  AOI211_X1 U15435 ( .C1(n13438), .C2(n13342), .A(n14633), .B(n13333), .ZN(
        n13437) );
  AOI22_X1 U15436 ( .A1(n14653), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n13334), 
        .B2(n14621), .ZN(n13335) );
  OAI21_X1 U15437 ( .B1(n13159), .B2(n14625), .A(n13335), .ZN(n13336) );
  AOI21_X1 U15438 ( .B1(n13437), .B2(n13395), .A(n13336), .ZN(n13337) );
  OAI211_X1 U15439 ( .C1(n13440), .C2(n13397), .A(n13338), .B(n13337), .ZN(
        P2_U3242) );
  XOR2_X1 U15440 ( .A(n13339), .B(n13347), .Z(n13341) );
  AOI21_X1 U15441 ( .B1(n13341), .B2(n13391), .A(n13340), .ZN(n13444) );
  AOI211_X1 U15442 ( .C1(n13442), .C2(n13357), .A(n14633), .B(n13331), .ZN(
        n13441) );
  INV_X1 U15443 ( .A(n13442), .ZN(n13346) );
  INV_X1 U15444 ( .A(n13343), .ZN(n13344) );
  AOI22_X1 U15445 ( .A1(n14653), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n13344), 
        .B2(n14621), .ZN(n13345) );
  OAI21_X1 U15446 ( .B1(n13346), .B2(n14625), .A(n13345), .ZN(n13352) );
  NAND2_X1 U15447 ( .A1(n13348), .A2(n13347), .ZN(n13349) );
  NAND2_X1 U15448 ( .A1(n13350), .A2(n13349), .ZN(n13445) );
  NOR2_X1 U15449 ( .A1(n13445), .A2(n13397), .ZN(n13351) );
  AOI211_X1 U15450 ( .C1(n13441), .C2(n13395), .A(n13352), .B(n13351), .ZN(
        n13353) );
  OAI21_X1 U15451 ( .B1(n14653), .B2(n13444), .A(n13353), .ZN(P2_U3243) );
  XNOR2_X1 U15452 ( .A(n13354), .B(n13364), .ZN(n13356) );
  AOI21_X1 U15453 ( .B1(n13356), .B2(n13391), .A(n13355), .ZN(n13449) );
  INV_X1 U15454 ( .A(n13357), .ZN(n13358) );
  AOI211_X1 U15455 ( .C1(n13447), .C2(n13373), .A(n14633), .B(n13358), .ZN(
        n13446) );
  INV_X1 U15456 ( .A(n13447), .ZN(n13362) );
  INV_X1 U15457 ( .A(n13359), .ZN(n13360) );
  AOI22_X1 U15458 ( .A1(n14653), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n13360), 
        .B2(n14621), .ZN(n13361) );
  OAI21_X1 U15459 ( .B1(n13362), .B2(n14625), .A(n13361), .ZN(n13366) );
  XOR2_X1 U15460 ( .A(n13364), .B(n13363), .Z(n13450) );
  NOR2_X1 U15461 ( .A1(n13450), .A2(n13397), .ZN(n13365) );
  AOI211_X1 U15462 ( .C1(n13446), .C2(n13395), .A(n13366), .B(n13365), .ZN(
        n13367) );
  OAI21_X1 U15463 ( .B1(n14653), .B2(n13449), .A(n13367), .ZN(P2_U3244) );
  XNOR2_X1 U15464 ( .A(n13368), .B(n13378), .ZN(n13371) );
  INV_X1 U15465 ( .A(n13369), .ZN(n13370) );
  AOI21_X1 U15466 ( .B1(n13371), .B2(n13391), .A(n13370), .ZN(n13454) );
  INV_X1 U15467 ( .A(n13372), .ZN(n13384) );
  INV_X1 U15468 ( .A(n13373), .ZN(n13374) );
  AOI211_X1 U15469 ( .C1(n13452), .C2(n13384), .A(n14633), .B(n13374), .ZN(
        n13451) );
  AOI22_X1 U15470 ( .A1(n14653), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n13375), 
        .B2(n14621), .ZN(n13376) );
  OAI21_X1 U15471 ( .B1(n13377), .B2(n14625), .A(n13376), .ZN(n13381) );
  XNOR2_X1 U15472 ( .A(n13379), .B(n13378), .ZN(n13455) );
  NOR2_X1 U15473 ( .A1(n13455), .A2(n13397), .ZN(n13380) );
  AOI211_X1 U15474 ( .C1(n13451), .C2(n13395), .A(n13381), .B(n13380), .ZN(
        n13382) );
  OAI21_X1 U15475 ( .B1(n14653), .B2(n13454), .A(n13382), .ZN(P2_U3245) );
  XNOR2_X1 U15476 ( .A(n13383), .B(n13390), .ZN(n13462) );
  AOI211_X1 U15477 ( .C1(n13459), .C2(n13385), .A(n14633), .B(n13372), .ZN(
        n13457) );
  AOI22_X1 U15478 ( .A1(n14653), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13386), 
        .B2(n14621), .ZN(n13387) );
  OAI21_X1 U15479 ( .B1(n13388), .B2(n14625), .A(n13387), .ZN(n13394) );
  XOR2_X1 U15480 ( .A(n13390), .B(n13389), .Z(n13392) );
  NAND2_X1 U15481 ( .A1(n13392), .A2(n13391), .ZN(n13461) );
  AOI21_X1 U15482 ( .B1(n13461), .B2(n13456), .A(n14653), .ZN(n13393) );
  AOI211_X1 U15483 ( .C1(n13457), .C2(n13395), .A(n13394), .B(n13393), .ZN(
        n13396) );
  OAI21_X1 U15484 ( .B1(n13397), .B2(n13462), .A(n13396), .ZN(P2_U3246) );
  OAI211_X1 U15485 ( .C1(n13160), .C2(n14723), .A(n13398), .B(n13399), .ZN(
        n13496) );
  MUX2_X1 U15486 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13496), .S(n14746), .Z(
        P2_U3530) );
  OAI211_X1 U15487 ( .C1(n13401), .C2(n14723), .A(n13400), .B(n13399), .ZN(
        n13497) );
  MUX2_X1 U15488 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13497), .S(n14746), .Z(
        P2_U3529) );
  NOR2_X1 U15489 ( .A1(n13403), .A2(n14723), .ZN(n13404) );
  OAI211_X1 U15490 ( .C1(n13416), .C2(n14723), .A(n13415), .B(n13414), .ZN(
        n13417) );
  MUX2_X1 U15491 ( .A(n13499), .B(P2_REG1_REG_27__SCAN_IN), .S(n14744), .Z(
        P2_U3526) );
  AOI21_X1 U15492 ( .B1(n14711), .B2(n13420), .A(n13419), .ZN(n13421) );
  OAI211_X1 U15493 ( .C1(n13495), .C2(n13423), .A(n13422), .B(n13421), .ZN(
        n13500) );
  MUX2_X1 U15494 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13500), .S(n14746), .Z(
        P2_U3525) );
  NAND2_X1 U15495 ( .A1(n13424), .A2(n14680), .ZN(n13426) );
  OAI211_X1 U15496 ( .C1(n13427), .C2(n14723), .A(n13426), .B(n13425), .ZN(
        n13428) );
  MUX2_X1 U15497 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13501), .S(n14746), .Z(
        P2_U3524) );
  AOI211_X1 U15498 ( .C1(n14711), .C2(n13432), .A(n13431), .B(n13430), .ZN(
        n13434) );
  OAI211_X1 U15499 ( .C1(n13495), .C2(n13435), .A(n13434), .B(n13433), .ZN(
        n13502) );
  MUX2_X1 U15500 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13502), .S(n14746), .Z(
        P2_U3523) );
  AOI211_X1 U15501 ( .C1(n14711), .C2(n13438), .A(n13437), .B(n13436), .ZN(
        n13439) );
  OAI21_X1 U15502 ( .B1(n13495), .B2(n13440), .A(n13439), .ZN(n13503) );
  MUX2_X1 U15503 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13503), .S(n14746), .Z(
        P2_U3522) );
  AOI21_X1 U15504 ( .B1(n14711), .B2(n13442), .A(n13441), .ZN(n13443) );
  OAI211_X1 U15505 ( .C1(n13495), .C2(n13445), .A(n13444), .B(n13443), .ZN(
        n13504) );
  MUX2_X1 U15506 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13504), .S(n14746), .Z(
        P2_U3521) );
  AOI21_X1 U15507 ( .B1(n14711), .B2(n13447), .A(n13446), .ZN(n13448) );
  OAI211_X1 U15508 ( .C1(n13495), .C2(n13450), .A(n13449), .B(n13448), .ZN(
        n13505) );
  MUX2_X1 U15509 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13505), .S(n14746), .Z(
        P2_U3520) );
  AOI21_X1 U15510 ( .B1(n14711), .B2(n13452), .A(n13451), .ZN(n13453) );
  OAI211_X1 U15511 ( .C1(n13495), .C2(n13455), .A(n13454), .B(n13453), .ZN(
        n13506) );
  MUX2_X1 U15512 ( .A(n13506), .B(P2_REG1_REG_20__SCAN_IN), .S(n14744), .Z(
        P2_U3519) );
  INV_X1 U15513 ( .A(n13456), .ZN(n13458) );
  AOI211_X1 U15514 ( .C1(n14711), .C2(n13459), .A(n13458), .B(n13457), .ZN(
        n13460) );
  OAI211_X1 U15515 ( .C1(n13495), .C2(n13462), .A(n13461), .B(n13460), .ZN(
        n13507) );
  MUX2_X1 U15516 ( .A(n13507), .B(P2_REG1_REG_19__SCAN_IN), .S(n14744), .Z(
        P2_U3518) );
  INV_X1 U15517 ( .A(n13463), .ZN(n13465) );
  AOI211_X1 U15518 ( .C1(n14711), .C2(n13466), .A(n13465), .B(n13464), .ZN(
        n13468) );
  OAI211_X1 U15519 ( .C1(n13469), .C2(n13495), .A(n13468), .B(n13467), .ZN(
        n13508) );
  MUX2_X1 U15520 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13508), .S(n14746), .Z(
        P2_U3517) );
  AOI211_X1 U15521 ( .C1(n14711), .C2(n13472), .A(n13471), .B(n13470), .ZN(
        n13473) );
  OAI21_X1 U15522 ( .B1(n13495), .B2(n13474), .A(n13473), .ZN(n13509) );
  MUX2_X1 U15523 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13509), .S(n14746), .Z(
        P2_U3516) );
  AOI21_X1 U15524 ( .B1(n14711), .B2(n13476), .A(n13475), .ZN(n13477) );
  OAI211_X1 U15525 ( .C1(n13495), .C2(n13479), .A(n13478), .B(n13477), .ZN(
        n13510) );
  MUX2_X1 U15526 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13510), .S(n14746), .Z(
        P2_U3515) );
  AOI21_X1 U15527 ( .B1(n14711), .B2(n13481), .A(n13480), .ZN(n13482) );
  OAI211_X1 U15528 ( .C1(n13495), .C2(n13484), .A(n13483), .B(n13482), .ZN(
        n13511) );
  MUX2_X1 U15529 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n13511), .S(n14746), .Z(
        P2_U3514) );
  AOI211_X1 U15530 ( .C1(n14711), .C2(n13487), .A(n13486), .B(n13485), .ZN(
        n13488) );
  OAI21_X1 U15531 ( .B1(n13495), .B2(n13489), .A(n13488), .ZN(n13512) );
  MUX2_X1 U15532 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n13512), .S(n14746), .Z(
        P2_U3513) );
  AOI21_X1 U15533 ( .B1(n14711), .B2(n13491), .A(n13490), .ZN(n13492) );
  OAI211_X1 U15534 ( .C1(n13495), .C2(n13494), .A(n13493), .B(n13492), .ZN(
        n13513) );
  MUX2_X1 U15535 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n13513), .S(n14746), .Z(
        P2_U3510) );
  MUX2_X1 U15536 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13496), .S(n14731), .Z(
        P2_U3498) );
  MUX2_X1 U15537 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13497), .S(n14731), .Z(
        P2_U3497) );
  MUX2_X1 U15538 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13498), .S(n14731), .Z(
        P2_U3495) );
  MUX2_X1 U15539 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13499), .S(n14731), .Z(
        P2_U3494) );
  MUX2_X1 U15540 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13500), .S(n14731), .Z(
        P2_U3493) );
  MUX2_X1 U15541 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13501), .S(n14731), .Z(
        P2_U3492) );
  MUX2_X1 U15542 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13502), .S(n14731), .Z(
        P2_U3491) );
  MUX2_X1 U15543 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13503), .S(n14731), .Z(
        P2_U3490) );
  MUX2_X1 U15544 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13504), .S(n14731), .Z(
        P2_U3489) );
  MUX2_X1 U15545 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13505), .S(n14731), .Z(
        P2_U3488) );
  MUX2_X1 U15546 ( .A(n13506), .B(P2_REG0_REG_20__SCAN_IN), .S(n14729), .Z(
        P2_U3487) );
  MUX2_X1 U15547 ( .A(n13507), .B(P2_REG0_REG_19__SCAN_IN), .S(n14729), .Z(
        P2_U3486) );
  MUX2_X1 U15548 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13508), .S(n14731), .Z(
        P2_U3484) );
  MUX2_X1 U15549 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13509), .S(n14731), .Z(
        P2_U3481) );
  MUX2_X1 U15550 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13510), .S(n14731), .Z(
        P2_U3478) );
  MUX2_X1 U15551 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n13511), .S(n14731), .Z(
        P2_U3475) );
  MUX2_X1 U15552 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n13512), .S(n14731), .Z(
        P2_U3472) );
  MUX2_X1 U15553 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n13513), .S(n14731), .Z(
        P2_U3463) );
  INV_X1 U15554 ( .A(n13514), .ZN(n14129) );
  NOR4_X1 U15555 ( .A1(n13515), .A2(P2_IR_REG_30__SCAN_IN), .A3(n9884), .A4(
        P2_U3088), .ZN(n13516) );
  AOI21_X1 U15556 ( .B1(n13519), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n13516), 
        .ZN(n13517) );
  OAI21_X1 U15557 ( .B1(n14129), .B2(n13526), .A(n13517), .ZN(P2_U3296) );
  AOI21_X1 U15558 ( .B1(n13519), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n13518), 
        .ZN(n13520) );
  OAI21_X1 U15559 ( .B1(n13521), .B2(n13526), .A(n13520), .ZN(P2_U3299) );
  INV_X1 U15560 ( .A(n13522), .ZN(n14133) );
  OAI222_X1 U15561 ( .A1(n13526), .A2(n14133), .B1(n13525), .B2(P2_U3088), 
        .C1(n13524), .C2(n13523), .ZN(P2_U3300) );
  MUX2_X1 U15562 ( .A(n13527), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  INV_X1 U15563 ( .A(n13529), .ZN(n13800) );
  OAI22_X1 U15564 ( .A1(n14394), .A2(n13800), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13530), .ZN(n13532) );
  OAI22_X1 U15565 ( .A1(n13792), .A2(n14378), .B1(n14377), .B2(n13794), .ZN(
        n13531) );
  AOI211_X1 U15566 ( .C1(n14014), .C2(n14389), .A(n13532), .B(n13531), .ZN(
        n13533) );
  OAI21_X1 U15567 ( .B1(n13534), .B2(n14384), .A(n13533), .ZN(P1_U3214) );
  XOR2_X1 U15568 ( .A(n13536), .B(n13535), .Z(n13542) );
  OR2_X1 U15569 ( .A1(n13581), .A2(n13983), .ZN(n13538) );
  NAND2_X1 U15570 ( .A1(n13901), .A2(n13954), .ZN(n13537) );
  AND2_X1 U15571 ( .A1(n13538), .A2(n13537), .ZN(n14039) );
  OAI22_X1 U15572 ( .A1(n13647), .A2(n14039), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15040), .ZN(n13539) );
  AOI21_X1 U15573 ( .B1(n13876), .B2(n13649), .A(n13539), .ZN(n13541) );
  NAND2_X1 U15574 ( .A1(n13869), .A2(n14389), .ZN(n13540) );
  OAI211_X1 U15575 ( .C1(n13542), .C2(n14384), .A(n13541), .B(n13540), .ZN(
        P1_U3216) );
  OAI21_X1 U15576 ( .B1(n10098), .B2(n13544), .A(n13543), .ZN(n13545) );
  NAND3_X1 U15577 ( .A1(n13546), .A2(n14356), .A3(n13545), .ZN(n13550) );
  OAI22_X1 U15578 ( .A1(n13547), .A2(n13983), .B1(n8691), .B2(n13982), .ZN(
        n14481) );
  AOI22_X1 U15579 ( .A1(n14358), .A2(n14481), .B1(n14389), .B2(n14486), .ZN(
        n13549) );
  MUX2_X1 U15580 ( .A(n14394), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n13548) );
  NAND3_X1 U15581 ( .A1(n13550), .A2(n13549), .A3(n13548), .ZN(P1_U3218) );
  AOI22_X1 U15582 ( .A1(n13629), .A2(n13662), .B1(n13625), .B2(n13900), .ZN(
        n13551) );
  NAND2_X1 U15583 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13771)
         );
  OAI211_X1 U15584 ( .C1(n14394), .C2(n13939), .A(n13551), .B(n13771), .ZN(
        n13562) );
  NAND2_X1 U15585 ( .A1(n13552), .A2(n13553), .ZN(n13555) );
  AND2_X1 U15586 ( .A1(n13555), .A2(n13554), .ZN(n13559) );
  NAND2_X1 U15587 ( .A1(n13552), .A2(n13556), .ZN(n13595) );
  NAND2_X1 U15588 ( .A1(n13595), .A2(n13557), .ZN(n13558) );
  AOI211_X1 U15589 ( .C1(n13560), .C2(n13559), .A(n14384), .B(n13558), .ZN(
        n13561) );
  AOI211_X1 U15590 ( .C1(n14063), .C2(n14389), .A(n13562), .B(n13561), .ZN(
        n13563) );
  INV_X1 U15591 ( .A(n13563), .ZN(P1_U3219) );
  AOI21_X1 U15592 ( .B1(n13565), .B2(n13564), .A(n6528), .ZN(n13572) );
  INV_X1 U15593 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n13566) );
  OAI22_X1 U15594 ( .A1(n14394), .A2(n13567), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13566), .ZN(n13570) );
  OAI22_X1 U15595 ( .A1(n13938), .A2(n14378), .B1(n14377), .B2(n13568), .ZN(
        n13569) );
  AOI211_X1 U15596 ( .C1(n14051), .C2(n14389), .A(n13570), .B(n13569), .ZN(
        n13571) );
  OAI21_X1 U15597 ( .B1(n13572), .B2(n14384), .A(n13571), .ZN(P1_U3223) );
  NAND2_X1 U15598 ( .A1(n13574), .A2(n13573), .ZN(n13586) );
  NAND2_X1 U15599 ( .A1(n13586), .A2(n13587), .ZN(n13576) );
  NAND2_X1 U15600 ( .A1(n13576), .A2(n13575), .ZN(n13577) );
  XOR2_X1 U15601 ( .A(n13578), .B(n13577), .Z(n13585) );
  INV_X1 U15602 ( .A(n13579), .ZN(n13834) );
  OAI22_X1 U15603 ( .A1(n14394), .A2(n13834), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13580), .ZN(n13583) );
  OAI22_X1 U15604 ( .A1(n13581), .A2(n14378), .B1(n14377), .B2(n13792), .ZN(
        n13582) );
  AOI211_X1 U15605 ( .C1(n14028), .C2(n14389), .A(n13583), .B(n13582), .ZN(
        n13584) );
  OAI21_X1 U15606 ( .B1(n13585), .B2(n14384), .A(n13584), .ZN(P1_U3225) );
  XOR2_X1 U15607 ( .A(n13587), .B(n13586), .Z(n13593) );
  INV_X1 U15608 ( .A(n13860), .ZN(n13589) );
  OAI22_X1 U15609 ( .A1(n14394), .A2(n13589), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13588), .ZN(n13591) );
  OAI22_X1 U15610 ( .A1(n13851), .A2(n14378), .B1(n14377), .B2(n13850), .ZN(
        n13590) );
  AOI211_X1 U15611 ( .C1(n13859), .C2(n14389), .A(n13591), .B(n13590), .ZN(
        n13592) );
  OAI21_X1 U15612 ( .B1(n13593), .B2(n14384), .A(n13592), .ZN(P1_U3229) );
  NAND2_X1 U15613 ( .A1(n13595), .A2(n13594), .ZN(n13598) );
  OAI211_X1 U15614 ( .C1(n13598), .C2(n13597), .A(n13596), .B(n14356), .ZN(
        n13603) );
  AND2_X1 U15615 ( .A1(n13661), .A2(n13955), .ZN(n13599) );
  AOI21_X1 U15616 ( .B1(n13956), .B2(n13954), .A(n13599), .ZN(n13921) );
  OAI22_X1 U15617 ( .A1(n13647), .A2(n13921), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13600), .ZN(n13601) );
  AOI21_X1 U15618 ( .B1(n13916), .B2(n13649), .A(n13601), .ZN(n13602) );
  OAI211_X1 U15619 ( .C1(n14114), .C2(n13653), .A(n13603), .B(n13602), .ZN(
        P1_U3233) );
  OAI21_X1 U15620 ( .B1(n13606), .B2(n13605), .A(n13604), .ZN(n13607) );
  NAND2_X1 U15621 ( .A1(n13607), .A2(n14356), .ZN(n13613) );
  NAND2_X1 U15622 ( .A1(n13661), .A2(n13954), .ZN(n13609) );
  NAND2_X1 U15623 ( .A1(n13660), .A2(n13955), .ZN(n13608) );
  AND2_X1 U15624 ( .A1(n13609), .A2(n13608), .ZN(n14044) );
  OAI22_X1 U15625 ( .A1(n13647), .A2(n14044), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13610), .ZN(n13611) );
  AOI21_X1 U15626 ( .B1(n13891), .B2(n13649), .A(n13611), .ZN(n13612) );
  OAI211_X1 U15627 ( .C1(n13653), .C2(n8687), .A(n13613), .B(n13612), .ZN(
        P1_U3235) );
  NAND2_X1 U15628 ( .A1(n13552), .A2(n13614), .ZN(n13615) );
  XOR2_X1 U15629 ( .A(n13616), .B(n13615), .Z(n13620) );
  AOI22_X1 U15630 ( .A1(n13629), .A2(n13953), .B1(n13625), .B2(n13956), .ZN(
        n13617) );
  NAND2_X1 U15631 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n13744)
         );
  OAI211_X1 U15632 ( .C1(n14394), .C2(n13964), .A(n13617), .B(n13744), .ZN(
        n13618) );
  AOI21_X1 U15633 ( .B1(n13967), .B2(n14389), .A(n13618), .ZN(n13619) );
  OAI21_X1 U15634 ( .B1(n13620), .B2(n14384), .A(n13619), .ZN(P1_U3238) );
  OAI211_X1 U15635 ( .C1(n13623), .C2(n13622), .A(n13621), .B(n14356), .ZN(
        n13632) );
  AOI22_X1 U15636 ( .A1(n13625), .A2(n13672), .B1(n13649), .B2(n13624), .ZN(
        n13631) );
  OAI22_X1 U15637 ( .A1(n13653), .A2(n13627), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13626), .ZN(n13628) );
  AOI21_X1 U15638 ( .B1(n13629), .B2(n13674), .A(n13628), .ZN(n13630) );
  NAND3_X1 U15639 ( .A1(n13632), .A2(n13631), .A3(n13630), .ZN(P1_U3239) );
  XOR2_X1 U15640 ( .A(n13634), .B(n13633), .Z(n13642) );
  INV_X1 U15641 ( .A(n13635), .ZN(n13813) );
  NAND2_X1 U15642 ( .A1(n13659), .A2(n13954), .ZN(n13637) );
  NAND2_X1 U15643 ( .A1(n13658), .A2(n13955), .ZN(n13636) );
  NAND2_X1 U15644 ( .A1(n13637), .A2(n13636), .ZN(n13812) );
  AOI22_X1 U15645 ( .A1(n14358), .A2(n13812), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13638) );
  OAI21_X1 U15646 ( .B1(n13813), .B2(n14394), .A(n13638), .ZN(n13639) );
  AOI21_X1 U15647 ( .B1(n13640), .B2(n14389), .A(n13639), .ZN(n13641) );
  OAI21_X1 U15648 ( .B1(n13642), .B2(n14384), .A(n13641), .ZN(P1_U3240) );
  OAI211_X1 U15649 ( .C1(n13645), .C2(n13644), .A(n13643), .B(n14356), .ZN(
        n13652) );
  INV_X1 U15650 ( .A(n14396), .ZN(n13646) );
  NAND2_X1 U15651 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n14454)
         );
  OAI21_X1 U15652 ( .B1(n13647), .B2(n13646), .A(n14454), .ZN(n13648) );
  AOI21_X1 U15653 ( .B1(n13650), .B2(n13649), .A(n13648), .ZN(n13651) );
  OAI211_X1 U15654 ( .C1(n13654), .C2(n13653), .A(n13652), .B(n13651), .ZN(
        P1_U3241) );
  MUX2_X1 U15655 ( .A(n13776), .B(P1_DATAO_REG_31__SCAN_IN), .S(n13675), .Z(
        P1_U3591) );
  INV_X1 U15656 ( .A(P1_U4016), .ZN(n13679) );
  MUX2_X1 U15657 ( .A(n13655), .B(P1_DATAO_REG_30__SCAN_IN), .S(n13679), .Z(
        P1_U3590) );
  MUX2_X1 U15658 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13656), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U15659 ( .A(n13657), .B(P1_DATAO_REG_28__SCAN_IN), .S(n13675), .Z(
        P1_U3588) );
  MUX2_X1 U15660 ( .A(n13658), .B(P1_DATAO_REG_27__SCAN_IN), .S(n13679), .Z(
        P1_U3587) );
  MUX2_X1 U15661 ( .A(n13828), .B(P1_DATAO_REG_26__SCAN_IN), .S(n13679), .Z(
        P1_U3586) );
  MUX2_X1 U15662 ( .A(n13659), .B(P1_DATAO_REG_25__SCAN_IN), .S(n13679), .Z(
        P1_U3585) );
  MUX2_X1 U15663 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n13827), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15664 ( .A(n13660), .B(P1_DATAO_REG_23__SCAN_IN), .S(n13675), .Z(
        P1_U3583) );
  MUX2_X1 U15665 ( .A(n13901), .B(P1_DATAO_REG_22__SCAN_IN), .S(n13679), .Z(
        P1_U3582) );
  MUX2_X1 U15666 ( .A(n13661), .B(P1_DATAO_REG_21__SCAN_IN), .S(n13675), .Z(
        P1_U3581) );
  MUX2_X1 U15667 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n13900), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U15668 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n13956), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U15669 ( .A(n13662), .B(P1_DATAO_REG_18__SCAN_IN), .S(n13679), .Z(
        P1_U3578) );
  MUX2_X1 U15670 ( .A(n13953), .B(P1_DATAO_REG_17__SCAN_IN), .S(n13679), .Z(
        P1_U3577) );
  MUX2_X1 U15671 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n13663), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U15672 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n13664), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U15673 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n13665), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U15674 ( .A(n13666), .B(P1_DATAO_REG_13__SCAN_IN), .S(n13679), .Z(
        P1_U3573) );
  MUX2_X1 U15675 ( .A(n13667), .B(P1_DATAO_REG_12__SCAN_IN), .S(n13675), .Z(
        P1_U3572) );
  MUX2_X1 U15676 ( .A(n13668), .B(P1_DATAO_REG_11__SCAN_IN), .S(n13679), .Z(
        P1_U3571) );
  MUX2_X1 U15677 ( .A(n13669), .B(P1_DATAO_REG_10__SCAN_IN), .S(n13675), .Z(
        P1_U3570) );
  MUX2_X1 U15678 ( .A(n13670), .B(P1_DATAO_REG_9__SCAN_IN), .S(n13679), .Z(
        P1_U3569) );
  MUX2_X1 U15679 ( .A(n13671), .B(P1_DATAO_REG_8__SCAN_IN), .S(n13679), .Z(
        P1_U3568) );
  MUX2_X1 U15680 ( .A(n13672), .B(P1_DATAO_REG_7__SCAN_IN), .S(n13675), .Z(
        P1_U3567) );
  MUX2_X1 U15681 ( .A(n13673), .B(P1_DATAO_REG_6__SCAN_IN), .S(n13675), .Z(
        P1_U3566) );
  MUX2_X1 U15682 ( .A(n13674), .B(P1_DATAO_REG_5__SCAN_IN), .S(n13679), .Z(
        P1_U3565) );
  MUX2_X1 U15683 ( .A(n13676), .B(P1_DATAO_REG_4__SCAN_IN), .S(n13675), .Z(
        P1_U3564) );
  MUX2_X1 U15684 ( .A(n13677), .B(P1_DATAO_REG_3__SCAN_IN), .S(n13679), .Z(
        P1_U3563) );
  MUX2_X1 U15685 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n13678), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U15686 ( .A(n9279), .B(P1_DATAO_REG_1__SCAN_IN), .S(n13679), .Z(
        P1_U3561) );
  MUX2_X1 U15687 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n13680), .S(P1_U4016), .Z(
        P1_U3560) );
  OAI22_X1 U15688 ( .A1(n14456), .A2(n14139), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13681), .ZN(n13682) );
  AOI21_X1 U15689 ( .B1(n13683), .B2(n14448), .A(n13682), .ZN(n13691) );
  OAI211_X1 U15690 ( .C1(n13686), .C2(n13685), .A(n14445), .B(n13684), .ZN(
        n13690) );
  OAI211_X1 U15691 ( .C1(n13688), .C2(n13687), .A(n13766), .B(n13699), .ZN(
        n13689) );
  NAND3_X1 U15692 ( .A1(n13691), .A2(n13690), .A3(n13689), .ZN(P1_U3244) );
  INV_X1 U15693 ( .A(n13692), .ZN(n13707) );
  INV_X1 U15694 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n13693) );
  OAI22_X1 U15695 ( .A1(n14456), .A2(n14140), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13693), .ZN(n13694) );
  AOI21_X1 U15696 ( .B1(n13695), .B2(n14448), .A(n13694), .ZN(n13706) );
  MUX2_X1 U15697 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n9213), .S(n13696), .Z(
        n13697) );
  NAND3_X1 U15698 ( .A1(n13699), .A2(n13698), .A3(n13697), .ZN(n13700) );
  NAND3_X1 U15699 ( .A1(n13766), .A2(n13715), .A3(n13700), .ZN(n13705) );
  OAI211_X1 U15700 ( .C1(n13703), .C2(n13702), .A(n14445), .B(n13701), .ZN(
        n13704) );
  NAND4_X1 U15701 ( .A1(n13707), .A2(n13706), .A3(n13705), .A4(n13704), .ZN(
        P1_U3245) );
  OAI211_X1 U15702 ( .C1(n13710), .C2(n13709), .A(n14445), .B(n13708), .ZN(
        n13721) );
  AOI22_X1 U15703 ( .A1(n13725), .A2(P1_ADDR_REG_3__SCAN_IN), .B1(
        P1_REG3_REG_3__SCAN_IN), .B2(P1_U3086), .ZN(n13720) );
  NAND2_X1 U15704 ( .A1(n14448), .A2(n13711), .ZN(n13719) );
  MUX2_X1 U15705 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n14484), .S(n13712), .Z(
        n13713) );
  NAND3_X1 U15706 ( .A1(n13715), .A2(n13714), .A3(n13713), .ZN(n13716) );
  NAND3_X1 U15707 ( .A1(n13766), .A2(n13717), .A3(n13716), .ZN(n13718) );
  NAND4_X1 U15708 ( .A1(n13721), .A2(n13720), .A3(n13719), .A4(n13718), .ZN(
        P1_U3246) );
  NAND2_X1 U15709 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3086), .ZN(n14373)
         );
  INV_X1 U15710 ( .A(n14373), .ZN(n13724) );
  NOR2_X1 U15711 ( .A1(n13722), .A2(n13748), .ZN(n13723) );
  AOI211_X1 U15712 ( .C1(n13725), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n13724), 
        .B(n13723), .ZN(n13739) );
  INV_X1 U15713 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n13749) );
  NOR2_X1 U15714 ( .A1(n13748), .A2(n13749), .ZN(n13726) );
  AOI21_X1 U15715 ( .B1(n13749), .B2(n13748), .A(n13726), .ZN(n13731) );
  OAI21_X1 U15716 ( .B1(n13729), .B2(n13728), .A(n13727), .ZN(n13730) );
  NAND2_X1 U15717 ( .A1(n13731), .A2(n13730), .ZN(n13747) );
  OAI211_X1 U15718 ( .C1(n13731), .C2(n13730), .A(n13766), .B(n13747), .ZN(
        n13738) );
  XNOR2_X1 U15719 ( .A(n13741), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n13734) );
  AOI211_X1 U15720 ( .C1(n13735), .C2(n13734), .A(n13740), .B(n13764), .ZN(
        n13736) );
  INV_X1 U15721 ( .A(n13736), .ZN(n13737) );
  NAND3_X1 U15722 ( .A1(n13739), .A2(n13738), .A3(n13737), .ZN(P1_U3260) );
  XNOR2_X1 U15723 ( .A(n13754), .B(n6511), .ZN(n13742) );
  INV_X1 U15724 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n14071) );
  NOR2_X1 U15725 ( .A1(n14071), .A2(n13742), .ZN(n13756) );
  AOI211_X1 U15726 ( .C1(n13742), .C2(n14071), .A(n13756), .B(n13764), .ZN(
        n13743) );
  INV_X1 U15727 ( .A(n13743), .ZN(n13753) );
  INV_X1 U15728 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n13745) );
  OAI21_X1 U15729 ( .B1(n14456), .B2(n13745), .A(n13744), .ZN(n13746) );
  AOI21_X1 U15730 ( .B1(n13759), .B2(n14448), .A(n13746), .ZN(n13752) );
  OAI21_X1 U15731 ( .B1(n13749), .B2(n13748), .A(n13747), .ZN(n13758) );
  XNOR2_X1 U15732 ( .A(n13754), .B(n13758), .ZN(n13750) );
  NAND2_X1 U15733 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n13750), .ZN(n13761) );
  OAI211_X1 U15734 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n13750), .A(n13766), 
        .B(n13761), .ZN(n13751) );
  NAND3_X1 U15735 ( .A1(n13753), .A2(n13752), .A3(n13751), .ZN(P1_U3261) );
  NOR2_X1 U15736 ( .A1(n6511), .A2(n13754), .ZN(n13755) );
  NOR2_X1 U15737 ( .A1(n13756), .A2(n13755), .ZN(n13757) );
  XOR2_X1 U15738 ( .A(n13757), .B(P1_REG1_REG_19__SCAN_IN), .Z(n13765) );
  NAND2_X1 U15739 ( .A1(n13759), .A2(n13758), .ZN(n13760) );
  NAND2_X1 U15740 ( .A1(n13761), .A2(n13760), .ZN(n13763) );
  INV_X1 U15741 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n13762) );
  XOR2_X1 U15742 ( .A(n13763), .B(n13762), .Z(n13767) );
  NAND2_X1 U15743 ( .A1(n13765), .A2(n14445), .ZN(n13769) );
  AOI21_X1 U15744 ( .B1(n13767), .B2(n13766), .A(n14448), .ZN(n13768) );
  NAND2_X1 U15745 ( .A1(n13769), .A2(n13768), .ZN(n13770) );
  OAI21_X1 U15746 ( .B1(n14456), .B2(n7385), .A(n13771), .ZN(n13772) );
  NAND2_X1 U15747 ( .A1(n13782), .A2(n14092), .ZN(n13774) );
  XNOR2_X1 U15748 ( .A(n13774), .B(n13773), .ZN(n13775) );
  NAND2_X1 U15749 ( .A1(n13992), .A2(n14494), .ZN(n13780) );
  INV_X1 U15750 ( .A(n13994), .ZN(n13778) );
  NOR2_X1 U15751 ( .A1(n13941), .A2(n13778), .ZN(n13783) );
  AOI21_X1 U15752 ( .B1(n14498), .B2(P1_REG2_REG_31__SCAN_IN), .A(n13783), 
        .ZN(n13779) );
  OAI211_X1 U15753 ( .C1(n14088), .C2(n13978), .A(n13780), .B(n13779), .ZN(
        P1_U3263) );
  XNOR2_X1 U15754 ( .A(n13782), .B(n13781), .ZN(n13995) );
  NAND2_X1 U15755 ( .A1(n13995), .A2(n13989), .ZN(n13785) );
  AOI21_X1 U15756 ( .B1(n14498), .B2(P1_REG2_REG_30__SCAN_IN), .A(n13783), 
        .ZN(n13784) );
  OAI211_X1 U15757 ( .C1(n14092), .C2(n13978), .A(n13785), .B(n13784), .ZN(
        P1_U3264) );
  XNOR2_X1 U15758 ( .A(n13787), .B(n13786), .ZN(n14018) );
  NOR2_X1 U15759 ( .A1(n6884), .A2(n6878), .ZN(n13789) );
  AND2_X1 U15760 ( .A1(n13807), .A2(n13789), .ZN(n13791) );
  OR2_X1 U15761 ( .A1(n13792), .A2(n13982), .ZN(n13793) );
  OAI21_X1 U15762 ( .B1(n13794), .B2(n13983), .A(n13793), .ZN(n13795) );
  INV_X1 U15763 ( .A(n13795), .ZN(n13796) );
  NAND2_X1 U15764 ( .A1(n13797), .A2(n13796), .ZN(n14019) );
  AOI21_X1 U15765 ( .B1(n14014), .B2(n13811), .A(n13961), .ZN(n13798) );
  NAND2_X1 U15766 ( .A1(n14016), .A2(n14494), .ZN(n13803) );
  NAND2_X1 U15767 ( .A1(n13941), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n13799) );
  OAI21_X1 U15768 ( .B1(n14483), .B2(n13800), .A(n13799), .ZN(n13801) );
  AOI21_X1 U15769 ( .B1(n14014), .B2(n14487), .A(n13801), .ZN(n13802) );
  NAND2_X1 U15770 ( .A1(n13803), .A2(n13802), .ZN(n13804) );
  AOI21_X1 U15771 ( .B1(n14019), .B2(n13966), .A(n13804), .ZN(n13805) );
  OAI21_X1 U15772 ( .B1(n14018), .B2(n13991), .A(n13805), .ZN(P1_U3266) );
  INV_X1 U15773 ( .A(n13806), .ZN(n13810) );
  INV_X1 U15774 ( .A(n13807), .ZN(n13808) );
  AOI21_X1 U15775 ( .B1(n13810), .B2(n13809), .A(n13808), .ZN(n14022) );
  OAI211_X1 U15776 ( .C1(n13838), .C2(n14099), .A(n13811), .B(n14490), .ZN(
        n14020) );
  INV_X1 U15777 ( .A(n14020), .ZN(n13817) );
  INV_X1 U15778 ( .A(n13812), .ZN(n14021) );
  OAI22_X1 U15779 ( .A1(n13941), .A2(n14021), .B1(n13813), .B2(n14483), .ZN(
        n13814) );
  AOI21_X1 U15780 ( .B1(P1_REG2_REG_26__SCAN_IN), .B2(n13941), .A(n13814), 
        .ZN(n13815) );
  OAI21_X1 U15781 ( .B1(n14099), .B2(n13978), .A(n13815), .ZN(n13816) );
  AOI21_X1 U15782 ( .B1(n13817), .B2(n14494), .A(n13816), .ZN(n13823) );
  NAND2_X1 U15783 ( .A1(n13830), .A2(n13819), .ZN(n13821) );
  XNOR2_X1 U15784 ( .A(n13821), .B(n13820), .ZN(n14024) );
  NAND2_X1 U15785 ( .A1(n14024), .A2(n14268), .ZN(n13822) );
  OAI211_X1 U15786 ( .C1(n14022), .C2(n14274), .A(n13823), .B(n13822), .ZN(
        P1_U3267) );
  OAI21_X1 U15787 ( .B1(n13826), .B2(n13825), .A(n13824), .ZN(n13829) );
  AOI222_X1 U15788 ( .A1(n14529), .A2(n13829), .B1(n13828), .B2(n13955), .C1(
        n13827), .C2(n13954), .ZN(n14030) );
  OAI21_X1 U15789 ( .B1(n13832), .B2(n13831), .A(n13830), .ZN(n14031) );
  NAND2_X1 U15790 ( .A1(n13941), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n13833) );
  OAI21_X1 U15791 ( .B1(n14483), .B2(n13834), .A(n13833), .ZN(n13835) );
  AOI21_X1 U15792 ( .B1(n14028), .B2(n14487), .A(n13835), .ZN(n13840) );
  NAND2_X1 U15793 ( .A1(n13856), .A2(n14028), .ZN(n13836) );
  NAND2_X1 U15794 ( .A1(n13836), .A2(n14490), .ZN(n13837) );
  NOR2_X1 U15795 ( .A1(n13838), .A2(n13837), .ZN(n14027) );
  NAND2_X1 U15796 ( .A1(n14027), .A2(n14494), .ZN(n13839) );
  OAI211_X1 U15797 ( .C1(n14031), .C2(n13991), .A(n13840), .B(n13839), .ZN(
        n13841) );
  INV_X1 U15798 ( .A(n13841), .ZN(n13842) );
  OAI21_X1 U15799 ( .B1(n14030), .B2(n14498), .A(n13842), .ZN(P1_U3268) );
  INV_X1 U15800 ( .A(n13843), .ZN(n13844) );
  AOI21_X1 U15801 ( .B1(n13846), .B2(n13845), .A(n13844), .ZN(n14032) );
  AOI211_X1 U15802 ( .C1(n13849), .C2(n13848), .A(n14478), .B(n13847), .ZN(
        n13853) );
  OAI22_X1 U15803 ( .A1(n13851), .A2(n13982), .B1(n13850), .B2(n13983), .ZN(
        n13852) );
  NOR2_X1 U15804 ( .A1(n13853), .A2(n13852), .ZN(n13854) );
  OAI21_X1 U15805 ( .B1(n14032), .B2(n13855), .A(n13854), .ZN(n14033) );
  NAND2_X1 U15806 ( .A1(n14033), .A2(n13966), .ZN(n13864) );
  INV_X1 U15807 ( .A(n13856), .ZN(n13857) );
  AOI211_X1 U15808 ( .C1(n13859), .C2(n13858), .A(n13961), .B(n13857), .ZN(
        n14034) );
  AOI22_X1 U15809 ( .A1(n13941), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n13860), 
        .B2(n14466), .ZN(n13861) );
  OAI21_X1 U15810 ( .B1(n14104), .B2(n13978), .A(n13861), .ZN(n13862) );
  AOI21_X1 U15811 ( .B1(n14034), .B2(n14494), .A(n13862), .ZN(n13863) );
  OAI211_X1 U15812 ( .C1(n14032), .C2(n13865), .A(n13864), .B(n13863), .ZN(
        P1_U3269) );
  NAND2_X1 U15813 ( .A1(n13866), .A2(n13872), .ZN(n13867) );
  INV_X1 U15814 ( .A(n14042), .ZN(n13882) );
  AOI22_X1 U15815 ( .A1(n13869), .A2(n14487), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n14498), .ZN(n13881) );
  XNOR2_X1 U15816 ( .A(n13889), .B(n13869), .ZN(n13870) );
  OR2_X1 U15817 ( .A1(n13870), .A2(n13961), .ZN(n14038) );
  OAI21_X1 U15818 ( .B1(n13873), .B2(n13872), .A(n13871), .ZN(n13874) );
  NAND2_X1 U15819 ( .A1(n13874), .A2(n14529), .ZN(n14040) );
  INV_X1 U15820 ( .A(n14039), .ZN(n13875) );
  AOI21_X1 U15821 ( .B1(n13876), .B2(n14466), .A(n13875), .ZN(n13877) );
  OAI211_X1 U15822 ( .C1(n13878), .C2(n14038), .A(n14040), .B(n13877), .ZN(
        n13879) );
  NAND2_X1 U15823 ( .A1(n13879), .A2(n13966), .ZN(n13880) );
  OAI211_X1 U15824 ( .C1(n13882), .C2(n13991), .A(n13881), .B(n13880), .ZN(
        P1_U3270) );
  XNOR2_X1 U15825 ( .A(n13883), .B(n13885), .ZN(n14049) );
  OAI21_X1 U15826 ( .B1(n13886), .B2(n13885), .A(n13884), .ZN(n14047) );
  AOI21_X1 U15827 ( .B1(n13888), .B2(n13903), .A(n13961), .ZN(n13890) );
  NAND2_X1 U15828 ( .A1(n13890), .A2(n13889), .ZN(n14045) );
  INV_X1 U15829 ( .A(n13891), .ZN(n13892) );
  OAI22_X1 U15830 ( .A1(n13941), .A2(n14044), .B1(n13892), .B2(n14483), .ZN(
        n13894) );
  NOR2_X1 U15831 ( .A1(n8687), .A2(n13978), .ZN(n13893) );
  AOI211_X1 U15832 ( .C1(n14498), .C2(P1_REG2_REG_22__SCAN_IN), .A(n13894), 
        .B(n13893), .ZN(n13895) );
  OAI21_X1 U15833 ( .B1(n13896), .B2(n14045), .A(n13895), .ZN(n13897) );
  AOI21_X1 U15834 ( .B1(n14047), .B2(n14268), .A(n13897), .ZN(n13898) );
  OAI21_X1 U15835 ( .B1(n14049), .B2(n14274), .A(n13898), .ZN(P1_U3271) );
  XNOR2_X1 U15836 ( .A(n13899), .B(n13907), .ZN(n13902) );
  AOI222_X1 U15837 ( .A1(n14529), .A2(n13902), .B1(n13901), .B2(n13955), .C1(
        n13900), .C2(n13954), .ZN(n14053) );
  AOI211_X1 U15838 ( .C1(n14051), .C2(n13925), .A(n13961), .B(n13887), .ZN(
        n14050) );
  INV_X1 U15839 ( .A(n14051), .ZN(n13906) );
  AOI22_X1 U15840 ( .A1(n13941), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n13904), 
        .B2(n14466), .ZN(n13905) );
  OAI21_X1 U15841 ( .B1(n13906), .B2(n13978), .A(n13905), .ZN(n13910) );
  XNOR2_X1 U15842 ( .A(n13908), .B(n13907), .ZN(n14054) );
  NOR2_X1 U15843 ( .A1(n14054), .A2(n13991), .ZN(n13909) );
  AOI211_X1 U15844 ( .C1(n14050), .C2(n14494), .A(n13910), .B(n13909), .ZN(
        n13911) );
  OAI21_X1 U15845 ( .B1(n14498), .B2(n14053), .A(n13911), .ZN(P1_U3272) );
  NAND2_X1 U15846 ( .A1(n13913), .A2(n13912), .ZN(n13914) );
  NAND2_X1 U15847 ( .A1(n13915), .A2(n13914), .ZN(n14057) );
  INV_X1 U15848 ( .A(n13916), .ZN(n13923) );
  NAND2_X1 U15849 ( .A1(n13918), .A2(n13917), .ZN(n13919) );
  NAND3_X1 U15850 ( .A1(n13920), .A2(n14529), .A3(n13919), .ZN(n13922) );
  AND2_X1 U15851 ( .A1(n13922), .A2(n13921), .ZN(n14056) );
  OAI21_X1 U15852 ( .B1(n13923), .B2(n14483), .A(n14056), .ZN(n13924) );
  NAND2_X1 U15853 ( .A1(n13924), .A2(n13966), .ZN(n13930) );
  OAI211_X1 U15854 ( .C1(n14114), .C2(n13937), .A(n14490), .B(n13925), .ZN(
        n14055) );
  INV_X1 U15855 ( .A(n14055), .ZN(n13928) );
  INV_X1 U15856 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n13926) );
  OAI22_X1 U15857 ( .A1(n14114), .A2(n13978), .B1(n13966), .B2(n13926), .ZN(
        n13927) );
  AOI21_X1 U15858 ( .B1(n13928), .B2(n14494), .A(n13927), .ZN(n13929) );
  OAI211_X1 U15859 ( .C1(n14057), .C2(n13991), .A(n13930), .B(n13929), .ZN(
        P1_U3273) );
  XNOR2_X1 U15860 ( .A(n13932), .B(n13931), .ZN(n14066) );
  XNOR2_X1 U15861 ( .A(n13933), .B(n13934), .ZN(n14060) );
  NAND2_X1 U15862 ( .A1(n14060), .A2(n14268), .ZN(n13947) );
  NAND2_X1 U15863 ( .A1(n13962), .A2(n14063), .ZN(n13935) );
  NAND2_X1 U15864 ( .A1(n13935), .A2(n14490), .ZN(n13936) );
  NOR2_X1 U15865 ( .A1(n13937), .A2(n13936), .ZN(n14061) );
  INV_X1 U15866 ( .A(n14063), .ZN(n13944) );
  OAI22_X1 U15867 ( .A1(n13938), .A2(n13983), .B1(n14365), .B2(n13982), .ZN(
        n14062) );
  INV_X1 U15868 ( .A(n13939), .ZN(n13940) );
  AOI22_X1 U15869 ( .A1(n13966), .A2(n14062), .B1(n13940), .B2(n14466), .ZN(
        n13943) );
  NAND2_X1 U15870 ( .A1(n13941), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n13942) );
  OAI211_X1 U15871 ( .C1(n13944), .C2(n13978), .A(n13943), .B(n13942), .ZN(
        n13945) );
  AOI21_X1 U15872 ( .B1(n14061), .B2(n14494), .A(n13945), .ZN(n13946) );
  OAI211_X1 U15873 ( .C1(n14066), .C2(n14274), .A(n13947), .B(n13946), .ZN(
        P1_U3274) );
  XNOR2_X1 U15874 ( .A(n13948), .B(n13950), .ZN(n14068) );
  OR2_X1 U15875 ( .A1(n13981), .A2(n13980), .ZN(n13985) );
  NAND2_X1 U15876 ( .A1(n13985), .A2(n13949), .ZN(n13952) );
  INV_X1 U15877 ( .A(n13950), .ZN(n13951) );
  XNOR2_X1 U15878 ( .A(n13952), .B(n13951), .ZN(n13958) );
  AOI22_X1 U15879 ( .A1(n13956), .A2(n13955), .B1(n13954), .B2(n13953), .ZN(
        n13957) );
  OAI21_X1 U15880 ( .B1(n13958), .B2(n14478), .A(n13957), .ZN(n13959) );
  AOI21_X1 U15881 ( .B1(n14068), .B2(n14482), .A(n13959), .ZN(n14070) );
  INV_X1 U15882 ( .A(n13960), .ZN(n13974) );
  AOI21_X1 U15883 ( .B1(n13974), .B2(n13967), .A(n13961), .ZN(n13963) );
  AND2_X1 U15884 ( .A1(n13963), .A2(n13962), .ZN(n14067) );
  INV_X1 U15885 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n13965) );
  OAI22_X1 U15886 ( .A1(n13966), .A2(n13965), .B1(n13964), .B2(n14483), .ZN(
        n13969) );
  NOR2_X1 U15887 ( .A1(n12125), .A2(n13978), .ZN(n13968) );
  AOI211_X1 U15888 ( .C1(n14067), .C2(n14494), .A(n13969), .B(n13968), .ZN(
        n13971) );
  NAND2_X1 U15889 ( .A1(n14068), .A2(n14495), .ZN(n13970) );
  OAI211_X1 U15890 ( .C1(n14070), .C2(n13941), .A(n13971), .B(n13970), .ZN(
        P1_U3275) );
  XNOR2_X1 U15891 ( .A(n13973), .B(n13972), .ZN(n14076) );
  AOI21_X1 U15892 ( .B1(n14372), .B2(n13975), .A(n13960), .ZN(n14073) );
  INV_X1 U15893 ( .A(n14372), .ZN(n13979) );
  INV_X1 U15894 ( .A(n14375), .ZN(n13976) );
  AOI22_X1 U15895 ( .A1(n13941), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n13976), 
        .B2(n14466), .ZN(n13977) );
  OAI21_X1 U15896 ( .B1(n13979), .B2(n13978), .A(n13977), .ZN(n13988) );
  AOI21_X1 U15897 ( .B1(n13981), .B2(n13980), .A(n14478), .ZN(n13986) );
  OAI22_X1 U15898 ( .A1(n14365), .A2(n13983), .B1(n14366), .B2(n13982), .ZN(
        n13984) );
  AOI21_X1 U15899 ( .B1(n13986), .B2(n13985), .A(n13984), .ZN(n14075) );
  NOR2_X1 U15900 ( .A1(n14075), .A2(n14498), .ZN(n13987) );
  AOI211_X1 U15901 ( .C1(n14073), .C2(n13989), .A(n13988), .B(n13987), .ZN(
        n13990) );
  OAI21_X1 U15902 ( .B1(n13991), .B2(n14076), .A(n13990), .ZN(P1_U3276) );
  NOR2_X1 U15903 ( .A1(n13992), .A2(n13994), .ZN(n14085) );
  MUX2_X1 U15904 ( .A(n15044), .B(n14085), .S(n14540), .Z(n13993) );
  OAI21_X1 U15905 ( .B1(n14088), .B2(n14084), .A(n13993), .ZN(P1_U3559) );
  INV_X1 U15906 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n13996) );
  AOI21_X1 U15907 ( .B1(n13995), .B2(n14490), .A(n13994), .ZN(n14089) );
  MUX2_X1 U15908 ( .A(n13996), .B(n14089), .S(n14540), .Z(n13997) );
  OAI21_X1 U15909 ( .B1(n14092), .B2(n14084), .A(n13997), .ZN(P1_U3558) );
  OAI211_X1 U15910 ( .C1(n14001), .C2(n14511), .A(n14000), .B(n13999), .ZN(
        n14002) );
  INV_X1 U15911 ( .A(n14002), .ZN(n14003) );
  OAI21_X1 U15912 ( .B1(n14008), .B2(n14405), .A(n14007), .ZN(n14093) );
  MUX2_X1 U15913 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14093), .S(n14540), .Z(
        P1_U3557) );
  AOI22_X1 U15914 ( .A1(n14010), .A2(n14490), .B1(n14522), .B2(n14009), .ZN(
        n14011) );
  MUX2_X1 U15915 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14094), .S(n14540), .Z(
        P1_U3556) );
  MUX2_X1 U15916 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14095), .S(n14540), .Z(
        P1_U3555) );
  INV_X1 U15917 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n14025) );
  OAI211_X1 U15918 ( .C1(n14022), .C2(n14478), .A(n14021), .B(n14020), .ZN(
        n14023) );
  AOI21_X1 U15919 ( .B1(n14024), .B2(n14518), .A(n14023), .ZN(n14096) );
  MUX2_X1 U15920 ( .A(n14025), .B(n14096), .S(n14540), .Z(n14026) );
  OAI21_X1 U15921 ( .B1(n14099), .B2(n14084), .A(n14026), .ZN(P1_U3554) );
  AOI21_X1 U15922 ( .B1(n14522), .B2(n14028), .A(n14027), .ZN(n14029) );
  OAI211_X1 U15923 ( .C1(n14405), .C2(n14031), .A(n14030), .B(n14029), .ZN(
        n14100) );
  MUX2_X1 U15924 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14100), .S(n14540), .Z(
        P1_U3553) );
  INV_X1 U15925 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n14036) );
  INV_X1 U15926 ( .A(n14032), .ZN(n14035) );
  MUX2_X1 U15927 ( .A(n14036), .B(n14101), .S(n14540), .Z(n14037) );
  OAI21_X1 U15928 ( .B1(n14104), .B2(n14084), .A(n14037), .ZN(P1_U3552) );
  INV_X1 U15929 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n15118) );
  NAND3_X1 U15930 ( .A1(n14040), .A2(n14039), .A3(n14038), .ZN(n14041) );
  AOI21_X1 U15931 ( .B1(n14042), .B2(n14518), .A(n14041), .ZN(n14105) );
  MUX2_X1 U15932 ( .A(n15118), .B(n14105), .S(n14540), .Z(n14043) );
  OAI21_X1 U15933 ( .B1(n14108), .B2(n14084), .A(n14043), .ZN(P1_U3551) );
  OAI211_X1 U15934 ( .C1(n14511), .C2(n8687), .A(n14045), .B(n14044), .ZN(
        n14046) );
  AOI21_X1 U15935 ( .B1(n14047), .B2(n14518), .A(n14046), .ZN(n14048) );
  OAI21_X1 U15936 ( .B1(n14478), .B2(n14049), .A(n14048), .ZN(n14109) );
  MUX2_X1 U15937 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14109), .S(n14540), .Z(
        P1_U3550) );
  AOI21_X1 U15938 ( .B1(n14522), .B2(n14051), .A(n14050), .ZN(n14052) );
  OAI211_X1 U15939 ( .C1(n14405), .C2(n14054), .A(n14053), .B(n14052), .ZN(
        n14110) );
  MUX2_X1 U15940 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14110), .S(n14540), .Z(
        P1_U3549) );
  OAI211_X1 U15941 ( .C1(n14057), .C2(n14405), .A(n14056), .B(n14055), .ZN(
        n14111) );
  MUX2_X1 U15942 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14111), .S(n14540), .Z(
        n14058) );
  INV_X1 U15943 ( .A(n14058), .ZN(n14059) );
  OAI21_X1 U15944 ( .B1(n14114), .B2(n14084), .A(n14059), .ZN(P1_U3548) );
  NAND2_X1 U15945 ( .A1(n14060), .A2(n14518), .ZN(n14065) );
  AOI211_X1 U15946 ( .C1(n14522), .C2(n14063), .A(n14062), .B(n14061), .ZN(
        n14064) );
  OAI211_X1 U15947 ( .C1(n14478), .C2(n14066), .A(n14065), .B(n14064), .ZN(
        n14115) );
  MUX2_X1 U15948 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14115), .S(n14540), .Z(
        P1_U3547) );
  AOI21_X1 U15949 ( .B1(n14068), .B2(n14517), .A(n14067), .ZN(n14069) );
  AND2_X1 U15950 ( .A1(n14070), .A2(n14069), .ZN(n14116) );
  MUX2_X1 U15951 ( .A(n14071), .B(n14116), .S(n14540), .Z(n14072) );
  OAI21_X1 U15952 ( .B1(n12125), .B2(n14084), .A(n14072), .ZN(P1_U3546) );
  AOI22_X1 U15953 ( .A1(n14073), .A2(n14490), .B1(n14522), .B2(n14372), .ZN(
        n14074) );
  OAI211_X1 U15954 ( .C1(n14076), .C2(n14405), .A(n14075), .B(n14074), .ZN(
        n14119) );
  MUX2_X1 U15955 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14119), .S(n14540), .Z(
        P1_U3545) );
  OAI211_X1 U15956 ( .C1(n14079), .C2(n14478), .A(n14078), .B(n14077), .ZN(
        n14080) );
  AOI21_X1 U15957 ( .B1(n14518), .B2(n14081), .A(n14080), .ZN(n14120) );
  MUX2_X1 U15958 ( .A(n14082), .B(n14120), .S(n14540), .Z(n14083) );
  OAI21_X1 U15959 ( .B1(n14124), .B2(n14084), .A(n14083), .ZN(P1_U3544) );
  INV_X1 U15960 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n14086) );
  MUX2_X1 U15961 ( .A(n14086), .B(n14085), .S(n14532), .Z(n14087) );
  OAI21_X1 U15962 ( .B1(n14088), .B2(n14123), .A(n14087), .ZN(P1_U3527) );
  MUX2_X1 U15963 ( .A(n14090), .B(n14089), .S(n14532), .Z(n14091) );
  OAI21_X1 U15964 ( .B1(n14092), .B2(n14123), .A(n14091), .ZN(P1_U3526) );
  MUX2_X1 U15965 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14093), .S(n14532), .Z(
        P1_U3525) );
  MUX2_X1 U15966 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14094), .S(n14532), .Z(
        P1_U3524) );
  MUX2_X1 U15967 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14095), .S(n14532), .Z(
        P1_U3523) );
  INV_X1 U15968 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n14097) );
  MUX2_X1 U15969 ( .A(n14097), .B(n14096), .S(n14532), .Z(n14098) );
  OAI21_X1 U15970 ( .B1(n14099), .B2(n14123), .A(n14098), .ZN(P1_U3522) );
  MUX2_X1 U15971 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14100), .S(n14532), .Z(
        P1_U3521) );
  INV_X1 U15972 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n14102) );
  MUX2_X1 U15973 ( .A(n14102), .B(n14101), .S(n14532), .Z(n14103) );
  OAI21_X1 U15974 ( .B1(n14104), .B2(n14123), .A(n14103), .ZN(P1_U3520) );
  INV_X1 U15975 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n14106) );
  MUX2_X1 U15976 ( .A(n14106), .B(n14105), .S(n14532), .Z(n14107) );
  OAI21_X1 U15977 ( .B1(n14108), .B2(n14123), .A(n14107), .ZN(P1_U3519) );
  MUX2_X1 U15978 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14109), .S(n14532), .Z(
        P1_U3518) );
  MUX2_X1 U15979 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14110), .S(n14532), .Z(
        P1_U3517) );
  MUX2_X1 U15980 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14111), .S(n14532), .Z(
        n14112) );
  INV_X1 U15981 ( .A(n14112), .ZN(n14113) );
  OAI21_X1 U15982 ( .B1(n14114), .B2(n14123), .A(n14113), .ZN(P1_U3516) );
  MUX2_X1 U15983 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14115), .S(n14532), .Z(
        P1_U3515) );
  INV_X1 U15984 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n14117) );
  MUX2_X1 U15985 ( .A(n14117), .B(n14116), .S(n14532), .Z(n14118) );
  OAI21_X1 U15986 ( .B1(n12125), .B2(n14123), .A(n14118), .ZN(P1_U3513) );
  MUX2_X1 U15987 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14119), .S(n14532), .Z(
        P1_U3510) );
  INV_X1 U15988 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n14121) );
  MUX2_X1 U15989 ( .A(n14121), .B(n14120), .S(n14532), .Z(n14122) );
  OAI21_X1 U15990 ( .B1(n14124), .B2(n14123), .A(n14122), .ZN(P1_U3507) );
  NOR4_X1 U15991 ( .A1(n6969), .A2(P1_IR_REG_30__SCAN_IN), .A3(n14125), .A4(
        P1_U3086), .ZN(n14126) );
  AOI21_X1 U15992 ( .B1(n14127), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n14126), 
        .ZN(n14128) );
  OAI21_X1 U15993 ( .B1(n14129), .B2(n12134), .A(n14128), .ZN(P1_U3324) );
  OAI222_X1 U15994 ( .A1(n14135), .A2(n14131), .B1(n12134), .B2(n14130), .C1(
        n8006), .C2(P1_U3086), .ZN(P1_U3326) );
  OAI222_X1 U15995 ( .A1(n14135), .A2(n14134), .B1(n12134), .B2(n14133), .C1(
        n14132), .C2(P1_U3086), .ZN(P1_U3328) );
  MUX2_X1 U15996 ( .A(n14137), .B(n14136), .S(P1_U3086), .Z(P1_U3333) );
  MUX2_X1 U15997 ( .A(n14138), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U15998 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n14227) );
  INV_X1 U15999 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14158) );
  INV_X1 U16000 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n14156) );
  XOR2_X1 U16001 ( .A(n14156), .B(P1_ADDR_REG_12__SCAN_IN), .Z(n14211) );
  INV_X1 U16002 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14154) );
  INV_X1 U16003 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n14152) );
  INV_X1 U16004 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n14151) );
  XOR2_X1 U16005 ( .A(n14151), .B(P1_ADDR_REG_9__SCAN_IN), .Z(n14197) );
  NOR2_X1 U16006 ( .A1(n14758), .A2(P1_ADDR_REG_0__SCAN_IN), .ZN(n14168) );
  INV_X1 U16007 ( .A(n14168), .ZN(n14167) );
  XNOR2_X1 U16008 ( .A(n14140), .B(P3_ADDR_REG_2__SCAN_IN), .ZN(n14172) );
  INV_X1 U16009 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n14143) );
  INV_X1 U16010 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n14145) );
  XNOR2_X1 U16011 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n14148), .ZN(n14190) );
  INV_X1 U16012 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n14191) );
  XNOR2_X1 U16013 ( .A(n14149), .B(P1_ADDR_REG_8__SCAN_IN), .ZN(n14162) );
  NAND2_X1 U16014 ( .A1(n14197), .A2(n14196), .ZN(n14150) );
  XOR2_X1 U16015 ( .A(P1_ADDR_REG_10__SCAN_IN), .B(n14153), .Z(n14161) );
  XOR2_X1 U16016 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .Z(n14159) );
  NAND2_X1 U16017 ( .A1(n14211), .A2(n14210), .ZN(n14155) );
  XNOR2_X1 U16018 ( .A(n14158), .B(P1_ADDR_REG_13__SCAN_IN), .ZN(n14212) );
  XOR2_X1 U16019 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .Z(n14216) );
  XOR2_X1 U16020 ( .A(n14217), .B(n14216), .Z(n14430) );
  XOR2_X1 U16021 ( .A(n14160), .B(n14159), .Z(n14206) );
  XOR2_X1 U16022 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(n14161), .Z(n14261) );
  XOR2_X1 U16023 ( .A(n14163), .B(n14162), .Z(n14195) );
  NAND2_X1 U16024 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n14165), .ZN(n14180) );
  XNOR2_X1 U16025 ( .A(n14167), .B(n14166), .ZN(n14169) );
  NAND2_X1 U16026 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14169), .ZN(n14171) );
  AOI21_X1 U16027 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n14758), .A(n14168), .ZN(
        n15171) );
  NOR2_X1 U16028 ( .A1(n15171), .A2(n15170), .ZN(n15180) );
  XOR2_X1 U16029 ( .A(n14169), .B(P2_ADDR_REG_1__SCAN_IN), .Z(n15179) );
  NAND2_X1 U16030 ( .A1(n15180), .A2(n15179), .ZN(n14170) );
  XNOR2_X1 U16031 ( .A(n14173), .B(n14172), .ZN(n14175) );
  NAND2_X1 U16032 ( .A1(n14174), .A2(n14175), .ZN(n14177) );
  NAND2_X1 U16033 ( .A1(n14254), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n14176) );
  XNOR2_X1 U16034 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n14178), .ZN(n15175) );
  INV_X1 U16035 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15177) );
  NAND2_X1 U16036 ( .A1(n15176), .A2(n15175), .ZN(n15174) );
  OAI21_X1 U16037 ( .B1(n14179), .B2(n15177), .A(n15174), .ZN(n15167) );
  XNOR2_X1 U16038 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n14181), .ZN(n14182) );
  XNOR2_X1 U16039 ( .A(n14183), .B(n14182), .ZN(n15169) );
  NAND2_X1 U16040 ( .A1(n14184), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14189) );
  XOR2_X1 U16041 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n14185), .Z(n14187) );
  XOR2_X1 U16042 ( .A(n14187), .B(n14186), .Z(n14255) );
  NAND2_X1 U16043 ( .A1(n14189), .A2(n14188), .ZN(n14192) );
  NAND2_X1 U16044 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n14192), .ZN(n14193) );
  XOR2_X1 U16045 ( .A(n14191), .B(n14190), .Z(n15172) );
  INV_X1 U16046 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n14584) );
  XNOR2_X1 U16047 ( .A(n14584), .B(n14192), .ZN(n15173) );
  XNOR2_X1 U16048 ( .A(n14197), .B(n14196), .ZN(n14198) );
  NAND2_X1 U16049 ( .A1(n14200), .A2(n14198), .ZN(n14202) );
  NAND2_X1 U16050 ( .A1(n14202), .A2(n14201), .ZN(n14260) );
  INV_X1 U16051 ( .A(n14259), .ZN(n14204) );
  INV_X1 U16052 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n14601) );
  NAND2_X1 U16053 ( .A1(n14204), .A2(n14203), .ZN(n14208) );
  INV_X1 U16054 ( .A(n14208), .ZN(n14205) );
  NOR2_X1 U16055 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n14419), .ZN(n14209) );
  XNOR2_X1 U16056 ( .A(n14211), .B(n14210), .ZN(n14423) );
  XOR2_X1 U16057 ( .A(n14213), .B(n14212), .Z(n14214) );
  NOR2_X1 U16058 ( .A1(n14215), .A2(n14214), .ZN(n14427) );
  INV_X1 U16059 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n14219) );
  INV_X1 U16060 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14457) );
  XOR2_X1 U16061 ( .A(n14457), .B(P3_ADDR_REG_15__SCAN_IN), .Z(n14222) );
  XOR2_X1 U16062 ( .A(n14223), .B(n14222), .Z(n14220) );
  INV_X1 U16063 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n14231) );
  XOR2_X1 U16064 ( .A(n14231), .B(P3_ADDR_REG_16__SCAN_IN), .Z(n14226) );
  NAND2_X1 U16065 ( .A1(n14223), .A2(n14222), .ZN(n14224) );
  XNOR2_X1 U16066 ( .A(n14226), .B(n14229), .ZN(n14438) );
  NOR2_X1 U16067 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14228), .ZN(n14230) );
  OAI22_X1 U16068 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n14231), .B1(n14230), 
        .B2(n14229), .ZN(n14234) );
  XNOR2_X1 U16069 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n14234), .ZN(n14235) );
  XNOR2_X1 U16070 ( .A(n14236), .B(n14235), .ZN(n14233) );
  XNOR2_X1 U16071 ( .A(n14233), .B(n14232), .ZN(n14280) );
  NOR2_X1 U16072 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n14234), .ZN(n14238) );
  NOR2_X1 U16073 ( .A1(n14236), .A2(n14235), .ZN(n14237) );
  XNOR2_X1 U16074 ( .A(n12508), .B(n14241), .ZN(n14242) );
  XNOR2_X1 U16075 ( .A(P1_ADDR_REG_18__SCAN_IN), .B(n14242), .ZN(n14239) );
  NOR2_X1 U16076 ( .A1(n14241), .A2(n12508), .ZN(n14244) );
  NOR2_X1 U16077 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n14242), .ZN(n14243) );
  NOR2_X1 U16078 ( .A1(n14244), .A2(n14243), .ZN(n14248) );
  XNOR2_X1 U16079 ( .A(n14245), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n14246) );
  XNOR2_X1 U16080 ( .A(n14246), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n14247) );
  XNOR2_X1 U16081 ( .A(n14248), .B(n14247), .ZN(n14249) );
  XNOR2_X1 U16082 ( .A(n14250), .B(n14249), .ZN(SUB_1596_U4) );
  XNOR2_X1 U16083 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n14251), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16084 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14252) );
  OAI21_X1 U16085 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14252), 
        .ZN(U28) );
  AOI21_X1 U16086 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14253) );
  OAI21_X1 U16087 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14253), 
        .ZN(U29) );
  XOR2_X1 U16088 ( .A(n14254), .B(P2_ADDR_REG_2__SCAN_IN), .Z(SUB_1596_U61) );
  XOR2_X1 U16089 ( .A(n14256), .B(n14255), .Z(SUB_1596_U57) );
  XNOR2_X1 U16090 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n14257), .ZN(SUB_1596_U55)
         );
  XOR2_X1 U16091 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n14258), .Z(SUB_1596_U54) );
  AOI21_X1 U16092 ( .B1(n14261), .B2(n14260), .A(n14259), .ZN(n14262) );
  XOR2_X1 U16093 ( .A(n14262), .B(P2_ADDR_REG_10__SCAN_IN), .Z(SUB_1596_U70)
         );
  INV_X1 U16094 ( .A(n14263), .ZN(n14265) );
  OAI211_X1 U16095 ( .C1(n14266), .C2(n14265), .A(n14264), .B(n13966), .ZN(
        n14267) );
  OAI21_X1 U16096 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n13966), .A(n14267), 
        .ZN(n14278) );
  NAND2_X1 U16097 ( .A1(n14269), .A2(n14268), .ZN(n14273) );
  OR2_X1 U16098 ( .A1(n14271), .A2(n14270), .ZN(n14272) );
  OAI211_X1 U16099 ( .C1(n14275), .C2(n14274), .A(n14273), .B(n14272), .ZN(
        n14276) );
  INV_X1 U16100 ( .A(n14276), .ZN(n14277) );
  OAI211_X1 U16101 ( .C1(n14483), .C2(n14279), .A(n14278), .B(n14277), .ZN(
        P1_U3280) );
  XNOR2_X1 U16102 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n14280), .ZN(SUB_1596_U63)
         );
  INV_X1 U16103 ( .A(n14307), .ZN(n14290) );
  XNOR2_X1 U16104 ( .A(n14281), .B(n14283), .ZN(n14324) );
  INV_X1 U16105 ( .A(n14324), .ZN(n14289) );
  XNOR2_X1 U16106 ( .A(n14282), .B(n14283), .ZN(n14288) );
  AOI222_X1 U16107 ( .A1(n14922), .A2(n14288), .B1(n14287), .B2(n14286), .C1(
        n14285), .C2(n14284), .ZN(n14326) );
  OAI21_X1 U16108 ( .B1(n14290), .B2(n14289), .A(n14326), .ZN(n14297) );
  INV_X1 U16109 ( .A(n14291), .ZN(n14293) );
  OAI22_X1 U16110 ( .A1(n14295), .A2(n14294), .B1(n14293), .B2(n14292), .ZN(
        n14296) );
  AOI21_X1 U16111 ( .B1(n14297), .B2(n14942), .A(n14296), .ZN(n14298) );
  OAI21_X1 U16112 ( .B1(n14942), .B2(n14299), .A(n14298), .ZN(P3_U3220) );
  XOR2_X1 U16113 ( .A(n14300), .B(n14301), .Z(n14320) );
  XNOR2_X1 U16114 ( .A(n14302), .B(n14301), .ZN(n14304) );
  OAI222_X1 U16115 ( .A1(n14917), .A2(n14306), .B1(n14919), .B2(n14305), .C1(
        n14304), .C2(n14303), .ZN(n14318) );
  AOI21_X1 U16116 ( .B1(n14320), .B2(n14307), .A(n14318), .ZN(n14313) );
  NOR2_X1 U16117 ( .A1(n14308), .A2(n14979), .ZN(n14319) );
  AOI22_X1 U16118 ( .A1(n14319), .A2(n14310), .B1(n14938), .B2(n14309), .ZN(
        n14311) );
  OAI221_X1 U16119 ( .B1(n14944), .B2(n14313), .C1(n14942), .C2(n14312), .A(
        n14311), .ZN(P3_U3222) );
  AOI211_X1 U16120 ( .C1(n14323), .C2(n14316), .A(n14315), .B(n14314), .ZN(
        n14328) );
  AOI22_X1 U16121 ( .A1(n15164), .A2(n14328), .B1(n14317), .B2(n15162), .ZN(
        P3_U3471) );
  AOI211_X1 U16122 ( .C1(n14320), .C2(n14323), .A(n14319), .B(n14318), .ZN(
        n14330) );
  INV_X1 U16123 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14321) );
  AOI22_X1 U16124 ( .A1(n15164), .A2(n14330), .B1(n14321), .B2(n15162), .ZN(
        P3_U3470) );
  AOI22_X1 U16125 ( .A1(n14324), .A2(n14323), .B1(n14957), .B2(n14322), .ZN(
        n14325) );
  NAND2_X1 U16126 ( .A1(n14326), .A2(n14325), .ZN(n15163) );
  MUX2_X1 U16127 ( .A(n15163), .B(P3_REG0_REG_13__SCAN_IN), .S(n14991), .Z(
        P3_U3429) );
  INV_X1 U16128 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14327) );
  AOI22_X1 U16129 ( .A1(n14993), .A2(n14328), .B1(n14327), .B2(n14991), .ZN(
        P3_U3426) );
  INV_X1 U16130 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14329) );
  AOI22_X1 U16131 ( .A1(n14993), .A2(n14330), .B1(n14329), .B2(n14991), .ZN(
        P3_U3423) );
  INV_X1 U16132 ( .A(n14331), .ZN(n14336) );
  OAI21_X1 U16133 ( .B1(n14333), .B2(n14723), .A(n14332), .ZN(n14335) );
  AOI211_X1 U16134 ( .C1(n14671), .C2(n14336), .A(n14335), .B(n14334), .ZN(
        n14339) );
  AOI22_X1 U16135 ( .A1(n14746), .A2(n14339), .B1(n14337), .B2(n14744), .ZN(
        P2_U3511) );
  INV_X1 U16136 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14338) );
  AOI22_X1 U16137 ( .A1(n14731), .A2(n14339), .B1(n14338), .B2(n14729), .ZN(
        P2_U3466) );
  OAI22_X1 U16138 ( .A1(n14341), .A2(n14378), .B1(n14377), .B2(n14340), .ZN(
        n14347) );
  NAND2_X1 U16139 ( .A1(n14343), .A2(n14342), .ZN(n14344) );
  AOI21_X1 U16140 ( .B1(n14345), .B2(n14344), .A(n14384), .ZN(n14346) );
  AOI211_X1 U16141 ( .C1(n11174), .C2(n14389), .A(n14347), .B(n14346), .ZN(
        n14349) );
  OAI211_X1 U16142 ( .C1(n14394), .C2(n14350), .A(n14349), .B(n14348), .ZN(
        P1_U3215) );
  INV_X1 U16143 ( .A(n13643), .ZN(n14353) );
  OAI21_X1 U16144 ( .B1(n14353), .B2(n14352), .A(n14351), .ZN(n14355) );
  NAND2_X1 U16145 ( .A1(n14355), .A2(n14354), .ZN(n14357) );
  AOI222_X1 U16146 ( .A1(n14389), .A2(n14360), .B1(n14359), .B2(n14358), .C1(
        n14357), .C2(n14356), .ZN(n14363) );
  INV_X1 U16147 ( .A(n14361), .ZN(n14362) );
  OAI211_X1 U16148 ( .C1(n14394), .C2(n14364), .A(n14363), .B(n14362), .ZN(
        P1_U3226) );
  OAI22_X1 U16149 ( .A1(n14366), .A2(n14378), .B1(n14377), .B2(n14365), .ZN(
        n14371) );
  XOR2_X1 U16150 ( .A(n14368), .B(n14367), .Z(n14369) );
  NOR2_X1 U16151 ( .A1(n14369), .A2(n14384), .ZN(n14370) );
  AOI211_X1 U16152 ( .C1(n14372), .C2(n14389), .A(n14371), .B(n14370), .ZN(
        n14374) );
  OAI211_X1 U16153 ( .C1(n14394), .C2(n14375), .A(n14374), .B(n14373), .ZN(
        P1_U3228) );
  OAI22_X1 U16154 ( .A1(n14379), .A2(n14378), .B1(n14377), .B2(n14376), .ZN(
        n14388) );
  AOI21_X1 U16155 ( .B1(n14382), .B2(n14381), .A(n14380), .ZN(n14383) );
  INV_X1 U16156 ( .A(n14383), .ZN(n14386) );
  AOI21_X1 U16157 ( .B1(n14386), .B2(n14385), .A(n14384), .ZN(n14387) );
  AOI211_X1 U16158 ( .C1(n14390), .C2(n14389), .A(n14388), .B(n14387), .ZN(
        n14392) );
  OAI211_X1 U16159 ( .C1(n14394), .C2(n14393), .A(n14392), .B(n14391), .ZN(
        P1_U3236) );
  AOI211_X1 U16160 ( .C1(n14522), .C2(n14397), .A(n14396), .B(n14395), .ZN(
        n14398) );
  OAI21_X1 U16161 ( .B1(n14478), .B2(n14399), .A(n14398), .ZN(n14400) );
  AOI21_X1 U16162 ( .B1(n14401), .B2(n14518), .A(n14400), .ZN(n14415) );
  AOI22_X1 U16163 ( .A1(n14540), .A2(n14415), .B1(n14443), .B2(n14537), .ZN(
        P1_U3543) );
  AOI21_X1 U16164 ( .B1(n11174), .B2(n14522), .A(n14402), .ZN(n14404) );
  OAI211_X1 U16165 ( .C1(n14406), .C2(n14405), .A(n14404), .B(n14403), .ZN(
        n14407) );
  AOI21_X1 U16166 ( .B1(n14529), .B2(n14408), .A(n14407), .ZN(n14416) );
  AOI22_X1 U16167 ( .A1(n14540), .A2(n14416), .B1(n10048), .B2(n14537), .ZN(
        P1_U3542) );
  OAI21_X1 U16168 ( .B1(n14410), .B2(n14511), .A(n14409), .ZN(n14412) );
  AOI211_X1 U16169 ( .C1(n14518), .C2(n14413), .A(n14412), .B(n14411), .ZN(
        n14418) );
  AOI22_X1 U16170 ( .A1(n14540), .A2(n14418), .B1(n9581), .B2(n14537), .ZN(
        P1_U3539) );
  INV_X1 U16171 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n14414) );
  AOI22_X1 U16172 ( .A1(n14532), .A2(n14415), .B1(n14414), .B2(n14530), .ZN(
        P1_U3504) );
  INV_X1 U16173 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n15115) );
  AOI22_X1 U16174 ( .A1(n14532), .A2(n14416), .B1(n15115), .B2(n14530), .ZN(
        P1_U3501) );
  INV_X1 U16175 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14417) );
  AOI22_X1 U16176 ( .A1(n14532), .A2(n14418), .B1(n14417), .B2(n14530), .ZN(
        P1_U3492) );
  NOR2_X1 U16177 ( .A1(n14420), .A2(n14419), .ZN(n14421) );
  XOR2_X1 U16178 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n14421), .Z(SUB_1596_U69)
         );
  AOI21_X1 U16179 ( .B1(n14424), .B2(n14423), .A(n14422), .ZN(n14425) );
  XOR2_X1 U16180 ( .A(n14425), .B(P2_ADDR_REG_12__SCAN_IN), .Z(SUB_1596_U68)
         );
  NOR2_X1 U16181 ( .A1(n14427), .A2(n14426), .ZN(n14428) );
  XOR2_X1 U16182 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(n14428), .Z(SUB_1596_U67)
         );
  AOI21_X1 U16183 ( .B1(n14431), .B2(n14430), .A(n14429), .ZN(n14432) );
  XOR2_X1 U16184 ( .A(n14432), .B(P2_ADDR_REG_14__SCAN_IN), .Z(SUB_1596_U66)
         );
  NOR2_X1 U16185 ( .A1(n14434), .A2(n14433), .ZN(n14435) );
  XOR2_X1 U16186 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n14435), .Z(SUB_1596_U65)
         );
  AOI21_X1 U16187 ( .B1(n14438), .B2(n14437), .A(n14436), .ZN(n14439) );
  XOR2_X1 U16188 ( .A(n14439), .B(P2_ADDR_REG_16__SCAN_IN), .Z(SUB_1596_U64)
         );
  AOI21_X1 U16189 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14441), .A(n14440), 
        .ZN(n14452) );
  OAI21_X1 U16190 ( .B1(n14444), .B2(n14443), .A(n14442), .ZN(n14446) );
  NAND2_X1 U16191 ( .A1(n14446), .A2(n14445), .ZN(n14450) );
  NAND2_X1 U16192 ( .A1(n14448), .A2(n14447), .ZN(n14449) );
  OAI211_X1 U16193 ( .C1(n14452), .C2(n14451), .A(n14450), .B(n14449), .ZN(
        n14453) );
  INV_X1 U16194 ( .A(n14453), .ZN(n14455) );
  OAI211_X1 U16195 ( .C1(n14457), .C2(n14456), .A(n14455), .B(n14454), .ZN(
        P1_U3258) );
  AOI222_X1 U16196 ( .A1(n14459), .A2(n14487), .B1(n14458), .B2(n14466), .C1(
        P1_REG2_REG_7__SCAN_IN), .C2(n13941), .ZN(n14463) );
  AOI22_X1 U16197 ( .A1(n14461), .A2(n14495), .B1(n14494), .B2(n14460), .ZN(
        n14462) );
  OAI211_X1 U16198 ( .C1(n14498), .C2(n14464), .A(n14463), .B(n14462), .ZN(
        P1_U3286) );
  AOI222_X1 U16199 ( .A1(n14467), .A2(n14487), .B1(P1_REG2_REG_5__SCAN_IN), 
        .B2(n13941), .C1(n14466), .C2(n14465), .ZN(n14473) );
  INV_X1 U16200 ( .A(n14468), .ZN(n14471) );
  INV_X1 U16201 ( .A(n14469), .ZN(n14470) );
  AOI22_X1 U16202 ( .A1(n14471), .A2(n14495), .B1(n14494), .B2(n14470), .ZN(
        n14472) );
  OAI211_X1 U16203 ( .C1(n14498), .C2(n14474), .A(n14473), .B(n14472), .ZN(
        P1_U3288) );
  XNOR2_X1 U16204 ( .A(n14475), .B(n14476), .ZN(n14516) );
  XNOR2_X1 U16205 ( .A(n14477), .B(n14476), .ZN(n14479) );
  NOR2_X1 U16206 ( .A1(n14479), .A2(n14478), .ZN(n14480) );
  AOI211_X1 U16207 ( .C1(n14482), .C2(n14516), .A(n14481), .B(n14480), .ZN(
        n14513) );
  OAI22_X1 U16208 ( .A1(n13966), .A2(n14484), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n14483), .ZN(n14485) );
  AOI21_X1 U16209 ( .B1(n14487), .B2(n14486), .A(n14485), .ZN(n14497) );
  INV_X1 U16210 ( .A(n14488), .ZN(n14492) );
  INV_X1 U16211 ( .A(n14489), .ZN(n14491) );
  OAI211_X1 U16212 ( .C1(n14512), .C2(n14492), .A(n14491), .B(n14490), .ZN(
        n14510) );
  INV_X1 U16213 ( .A(n14510), .ZN(n14493) );
  AOI22_X1 U16214 ( .A1(n14495), .A2(n14516), .B1(n14494), .B2(n14493), .ZN(
        n14496) );
  OAI211_X1 U16215 ( .C1(n14498), .C2(n14513), .A(n14497), .B(n14496), .ZN(
        P1_U3290) );
  AND2_X1 U16216 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14500), .ZN(P1_U3294) );
  AND2_X1 U16217 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14500), .ZN(P1_U3295) );
  AND2_X1 U16218 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14500), .ZN(P1_U3296) );
  AND2_X1 U16219 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14500), .ZN(P1_U3297) );
  AND2_X1 U16220 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14500), .ZN(P1_U3298) );
  AND2_X1 U16221 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14500), .ZN(P1_U3299) );
  AND2_X1 U16222 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14500), .ZN(P1_U3300) );
  AND2_X1 U16223 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14500), .ZN(P1_U3301) );
  AND2_X1 U16224 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14500), .ZN(P1_U3302) );
  INV_X1 U16225 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n15135) );
  NOR2_X1 U16226 ( .A1(n14499), .A2(n15135), .ZN(P1_U3303) );
  AND2_X1 U16227 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14500), .ZN(P1_U3304) );
  AND2_X1 U16228 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14500), .ZN(P1_U3305) );
  AND2_X1 U16229 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14500), .ZN(P1_U3306) );
  AND2_X1 U16230 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14500), .ZN(P1_U3307) );
  AND2_X1 U16231 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14500), .ZN(P1_U3308) );
  AND2_X1 U16232 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14500), .ZN(P1_U3309) );
  AND2_X1 U16233 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14500), .ZN(P1_U3310) );
  AND2_X1 U16234 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14500), .ZN(P1_U3311) );
  AND2_X1 U16235 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14500), .ZN(P1_U3312) );
  AND2_X1 U16236 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14500), .ZN(P1_U3313) );
  AND2_X1 U16237 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14500), .ZN(P1_U3314) );
  AND2_X1 U16238 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14500), .ZN(P1_U3315) );
  AND2_X1 U16239 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14500), .ZN(P1_U3316) );
  AND2_X1 U16240 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14500), .ZN(P1_U3317) );
  AND2_X1 U16241 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14500), .ZN(P1_U3318) );
  INV_X1 U16242 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n15083) );
  NOR2_X1 U16243 ( .A1(n14499), .A2(n15083), .ZN(P1_U3319) );
  INV_X1 U16244 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n15105) );
  NOR2_X1 U16245 ( .A1(n14499), .A2(n15105), .ZN(P1_U3320) );
  AND2_X1 U16246 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14500), .ZN(P1_U3321) );
  AND2_X1 U16247 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14500), .ZN(P1_U3322) );
  AND2_X1 U16248 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14500), .ZN(P1_U3323) );
  INV_X1 U16249 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n14501) );
  AOI22_X1 U16250 ( .A1(n14532), .A2(n14502), .B1(n14501), .B2(n14530), .ZN(
        P1_U3462) );
  OAI21_X1 U16251 ( .B1(n14504), .B2(n14511), .A(n14503), .ZN(n14505) );
  AOI21_X1 U16252 ( .B1(n14506), .B2(n14517), .A(n14505), .ZN(n14507) );
  AND2_X1 U16253 ( .A1(n14508), .A2(n14507), .ZN(n14534) );
  INV_X1 U16254 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n14509) );
  AOI22_X1 U16255 ( .A1(n14532), .A2(n14534), .B1(n14509), .B2(n14530), .ZN(
        P1_U3465) );
  OAI21_X1 U16256 ( .B1(n14512), .B2(n14511), .A(n14510), .ZN(n14515) );
  INV_X1 U16257 ( .A(n14513), .ZN(n14514) );
  AOI211_X1 U16258 ( .C1(n14517), .C2(n14516), .A(n14515), .B(n14514), .ZN(
        n14536) );
  INV_X1 U16259 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n15132) );
  AOI22_X1 U16260 ( .A1(n14532), .A2(n14536), .B1(n15132), .B2(n14530), .ZN(
        P1_U3468) );
  NAND2_X1 U16261 ( .A1(n14519), .A2(n14518), .ZN(n14526) );
  INV_X1 U16262 ( .A(n14520), .ZN(n14525) );
  NAND2_X1 U16263 ( .A1(n14522), .A2(n14521), .ZN(n14523) );
  NAND4_X1 U16264 ( .A1(n14526), .A2(n14525), .A3(n14524), .A4(n14523), .ZN(
        n14527) );
  AOI21_X1 U16265 ( .B1(n14529), .B2(n14528), .A(n14527), .ZN(n14539) );
  INV_X1 U16266 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n14531) );
  AOI22_X1 U16267 ( .A1(n14532), .A2(n14539), .B1(n14531), .B2(n14530), .ZN(
        P1_U3471) );
  AOI22_X1 U16268 ( .A1(n14540), .A2(n14534), .B1(n14533), .B2(n14537), .ZN(
        P1_U3530) );
  INV_X1 U16269 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n14535) );
  AOI22_X1 U16270 ( .A1(n14540), .A2(n14536), .B1(n14535), .B2(n14537), .ZN(
        P1_U3531) );
  INV_X1 U16271 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n14538) );
  AOI22_X1 U16272 ( .A1(n14540), .A2(n14539), .B1(n14538), .B2(n14537), .ZN(
        P1_U3532) );
  NOR2_X1 U16273 ( .A1(n14610), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U16274 ( .A1(n14610), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n14555) );
  INV_X1 U16275 ( .A(n14541), .ZN(n14544) );
  INV_X1 U16276 ( .A(n14542), .ZN(n14543) );
  AOI211_X1 U16277 ( .C1(n14545), .C2(n14544), .A(n14543), .B(n14604), .ZN(
        n14546) );
  AOI21_X1 U16278 ( .B1(n14594), .B2(n14547), .A(n14546), .ZN(n14554) );
  INV_X1 U16279 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n14549) );
  NOR2_X1 U16280 ( .A1(n14549), .A2(n14548), .ZN(n14551) );
  OAI211_X1 U16281 ( .C1(n14552), .C2(n14551), .A(n14579), .B(n14550), .ZN(
        n14553) );
  NAND3_X1 U16282 ( .A1(n14555), .A2(n14554), .A3(n14553), .ZN(P2_U3215) );
  OAI21_X1 U16283 ( .B1(n14557), .B2(n14556), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n14558) );
  OAI21_X1 U16284 ( .B1(P2_STATE_REG_SCAN_IN), .B2(P2_REG3_REG_2__SCAN_IN), 
        .A(n14558), .ZN(n14570) );
  OAI21_X1 U16285 ( .B1(n14561), .B2(n14560), .A(n14559), .ZN(n14562) );
  INV_X1 U16286 ( .A(n14562), .ZN(n14563) );
  AND2_X1 U16287 ( .A1(n14586), .A2(n14563), .ZN(n14564) );
  AOI21_X1 U16288 ( .B1(n14610), .B2(P2_ADDR_REG_2__SCAN_IN), .A(n14564), .ZN(
        n14569) );
  OAI211_X1 U16289 ( .C1(n14567), .C2(n14566), .A(n14579), .B(n14565), .ZN(
        n14568) );
  NAND3_X1 U16290 ( .A1(n14570), .A2(n14569), .A3(n14568), .ZN(P2_U3216) );
  NOR2_X1 U16291 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9860), .ZN(n14576) );
  OAI211_X1 U16292 ( .C1(n14573), .C2(n14572), .A(n14586), .B(n14571), .ZN(
        n14574) );
  INV_X1 U16293 ( .A(n14574), .ZN(n14575) );
  AOI211_X1 U16294 ( .C1(n14594), .C2(n14577), .A(n14576), .B(n14575), .ZN(
        n14583) );
  OAI211_X1 U16295 ( .C1(n14581), .C2(n14580), .A(n14579), .B(n14578), .ZN(
        n14582) );
  OAI211_X1 U16296 ( .C1(n14602), .C2(n14584), .A(n14583), .B(n14582), .ZN(
        P2_U3221) );
  NOR2_X1 U16297 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n14585), .ZN(n14592) );
  OAI211_X1 U16298 ( .C1(n14589), .C2(n14588), .A(n14587), .B(n14586), .ZN(
        n14590) );
  INV_X1 U16299 ( .A(n14590), .ZN(n14591) );
  AOI211_X1 U16300 ( .C1(n14594), .C2(n14593), .A(n14592), .B(n14591), .ZN(
        n14600) );
  AOI211_X1 U16301 ( .C1(n14597), .C2(n14596), .A(n14614), .B(n14595), .ZN(
        n14598) );
  INV_X1 U16302 ( .A(n14598), .ZN(n14599) );
  OAI211_X1 U16303 ( .C1(n14602), .C2(n14601), .A(n14600), .B(n14599), .ZN(
        P2_U3224) );
  INV_X1 U16304 ( .A(n14603), .ZN(n14609) );
  AOI211_X1 U16305 ( .C1(n14607), .C2(n14606), .A(n14605), .B(n14604), .ZN(
        n14608) );
  AOI211_X1 U16306 ( .C1(P2_ADDR_REG_18__SCAN_IN), .C2(n14610), .A(n14609), 
        .B(n14608), .ZN(n14616) );
  AOI21_X1 U16307 ( .B1(n14612), .B2(P2_REG2_REG_18__SCAN_IN), .A(n14611), 
        .ZN(n14613) );
  OR2_X1 U16308 ( .A1(n14614), .A2(n14613), .ZN(n14615) );
  OAI211_X1 U16309 ( .C1(n14618), .C2(n14617), .A(n14616), .B(n14615), .ZN(
        P2_U3232) );
  INV_X1 U16310 ( .A(n14619), .ZN(n14626) );
  NAND2_X1 U16311 ( .A1(n14620), .A2(n13395), .ZN(n14624) );
  AOI22_X1 U16312 ( .A1(n14653), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n14622), 
        .B2(n14621), .ZN(n14623) );
  OAI211_X1 U16313 ( .C1(n14626), .C2(n14625), .A(n14624), .B(n14623), .ZN(
        n14627) );
  AOI21_X1 U16314 ( .B1(n14629), .B2(n14628), .A(n14627), .ZN(n14630) );
  OAI21_X1 U16315 ( .B1(n14653), .B2(n14631), .A(n14630), .ZN(P2_U3258) );
  XNOR2_X1 U16316 ( .A(n14632), .B(n14639), .ZN(n14679) );
  AOI21_X1 U16317 ( .B1(n14635), .B2(n14634), .A(n14633), .ZN(n14637) );
  NAND2_X1 U16318 ( .A1(n14637), .A2(n14636), .ZN(n14675) );
  NAND3_X1 U16319 ( .A1(n9993), .A2(n14639), .A3(n14638), .ZN(n14641) );
  AOI21_X1 U16320 ( .B1(n14642), .B2(n14641), .A(n14640), .ZN(n14644) );
  NOR2_X1 U16321 ( .A1(n14644), .A2(n14643), .ZN(n14676) );
  OAI22_X1 U16322 ( .A1(n14646), .A2(P2_REG3_REG_3__SCAN_IN), .B1(n14677), 
        .B2(n14645), .ZN(n14647) );
  INV_X1 U16323 ( .A(n14647), .ZN(n14648) );
  OAI211_X1 U16324 ( .C1(n10176), .C2(n14675), .A(n14676), .B(n14648), .ZN(
        n14649) );
  AOI21_X1 U16325 ( .B1(n14650), .B2(n14679), .A(n14649), .ZN(n14651) );
  AOI22_X1 U16326 ( .A1(n14653), .A2(n14652), .B1(n14651), .B2(n13330), .ZN(
        P2_U3262) );
  AND2_X1 U16327 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14656), .ZN(P2_U3266) );
  AND2_X1 U16328 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14656), .ZN(P2_U3267) );
  AND2_X1 U16329 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14656), .ZN(P2_U3268) );
  INV_X1 U16330 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n15127) );
  NOR2_X1 U16331 ( .A1(n14655), .A2(n15127), .ZN(P2_U3269) );
  AND2_X1 U16332 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14656), .ZN(P2_U3270) );
  AND2_X1 U16333 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14656), .ZN(P2_U3271) );
  AND2_X1 U16334 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14656), .ZN(P2_U3272) );
  AND2_X1 U16335 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14656), .ZN(P2_U3273) );
  AND2_X1 U16336 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14656), .ZN(P2_U3274) );
  AND2_X1 U16337 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14656), .ZN(P2_U3275) );
  AND2_X1 U16338 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14656), .ZN(P2_U3276) );
  AND2_X1 U16339 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14656), .ZN(P2_U3277) );
  AND2_X1 U16340 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14656), .ZN(P2_U3278) );
  AND2_X1 U16341 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14656), .ZN(P2_U3279) );
  AND2_X1 U16342 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14656), .ZN(P2_U3280) );
  AND2_X1 U16343 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14656), .ZN(P2_U3281) );
  AND2_X1 U16344 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14656), .ZN(P2_U3282) );
  AND2_X1 U16345 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n14656), .ZN(P2_U3283) );
  AND2_X1 U16346 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14656), .ZN(P2_U3284) );
  AND2_X1 U16347 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14656), .ZN(P2_U3285) );
  AND2_X1 U16348 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14656), .ZN(P2_U3286) );
  AND2_X1 U16349 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14656), .ZN(P2_U3287) );
  AND2_X1 U16350 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14656), .ZN(P2_U3288) );
  AND2_X1 U16351 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n14656), .ZN(P2_U3289) );
  AND2_X1 U16352 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14656), .ZN(P2_U3290) );
  AND2_X1 U16353 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14656), .ZN(P2_U3291) );
  AND2_X1 U16354 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14656), .ZN(P2_U3292) );
  AND2_X1 U16355 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14656), .ZN(P2_U3293) );
  INV_X1 U16356 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n15067) );
  NOR2_X1 U16357 ( .A1(n14655), .A2(n15067), .ZN(P2_U3294) );
  AND2_X1 U16358 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14656), .ZN(P2_U3295) );
  AOI22_X1 U16359 ( .A1(n14661), .A2(n14658), .B1(n14657), .B2(n14659), .ZN(
        P2_U3416) );
  AOI22_X1 U16360 ( .A1(n14661), .A2(n14660), .B1(n9308), .B2(n14659), .ZN(
        P2_U3417) );
  INV_X1 U16361 ( .A(n14662), .ZN(n14664) );
  AOI211_X1 U16362 ( .C1(n14671), .C2(n14665), .A(n14664), .B(n14663), .ZN(
        n14733) );
  INV_X1 U16363 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n15119) );
  AOI22_X1 U16364 ( .A1(n14731), .A2(n14733), .B1(n15119), .B2(n14729), .ZN(
        P2_U3430) );
  OAI21_X1 U16365 ( .B1(n14667), .B2(n14723), .A(n14666), .ZN(n14669) );
  AOI211_X1 U16366 ( .C1(n14671), .C2(n14670), .A(n14669), .B(n14668), .ZN(
        n14735) );
  INV_X1 U16367 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n14672) );
  AOI22_X1 U16368 ( .A1(n14731), .A2(n14735), .B1(n14672), .B2(n14729), .ZN(
        P2_U3433) );
  INV_X1 U16369 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n14673) );
  AOI22_X1 U16370 ( .A1(n14731), .A2(n14674), .B1(n14673), .B2(n14729), .ZN(
        P2_U3436) );
  OAI211_X1 U16371 ( .C1(n14677), .C2(n14723), .A(n14676), .B(n14675), .ZN(
        n14678) );
  AOI21_X1 U16372 ( .B1(n14680), .B2(n14679), .A(n14678), .ZN(n14736) );
  INV_X1 U16373 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n14681) );
  AOI22_X1 U16374 ( .A1(n14731), .A2(n14736), .B1(n14681), .B2(n14729), .ZN(
        P2_U3439) );
  INV_X1 U16375 ( .A(n14686), .ZN(n14688) );
  AOI21_X1 U16376 ( .B1(n14711), .B2(n14683), .A(n14682), .ZN(n14684) );
  OAI211_X1 U16377 ( .C1(n14718), .C2(n14686), .A(n14685), .B(n14684), .ZN(
        n14687) );
  AOI21_X1 U16378 ( .B1(n14728), .B2(n14688), .A(n14687), .ZN(n14737) );
  INV_X1 U16379 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n14689) );
  AOI22_X1 U16380 ( .A1(n14731), .A2(n14737), .B1(n14689), .B2(n14729), .ZN(
        P2_U3442) );
  AND2_X1 U16381 ( .A1(n14690), .A2(n14711), .ZN(n14691) );
  NOR2_X1 U16382 ( .A1(n14692), .A2(n14691), .ZN(n14697) );
  OR2_X1 U16383 ( .A1(n14694), .A2(n14718), .ZN(n14696) );
  OR2_X1 U16384 ( .A1(n14694), .A2(n14693), .ZN(n14695) );
  INV_X1 U16385 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n14699) );
  AOI22_X1 U16386 ( .A1(n14731), .A2(n14739), .B1(n14699), .B2(n14729), .ZN(
        P2_U3445) );
  INV_X1 U16387 ( .A(n14704), .ZN(n14707) );
  INV_X1 U16388 ( .A(n14700), .ZN(n14706) );
  AOI21_X1 U16389 ( .B1(n14711), .B2(n14702), .A(n14701), .ZN(n14703) );
  OAI21_X1 U16390 ( .B1(n14704), .B2(n14718), .A(n14703), .ZN(n14705) );
  AOI211_X1 U16391 ( .C1(n14728), .C2(n14707), .A(n14706), .B(n14705), .ZN(
        n14741) );
  INV_X1 U16392 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n14708) );
  AOI22_X1 U16393 ( .A1(n14731), .A2(n14741), .B1(n14708), .B2(n14729), .ZN(
        P2_U3448) );
  AOI21_X1 U16394 ( .B1(n14711), .B2(n14710), .A(n14709), .ZN(n14712) );
  OAI21_X1 U16395 ( .B1(n14713), .B2(n14718), .A(n14712), .ZN(n14714) );
  AOI211_X1 U16396 ( .C1(n14728), .C2(n14716), .A(n14715), .B(n14714), .ZN(
        n14743) );
  INV_X1 U16397 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n14717) );
  AOI22_X1 U16398 ( .A1(n14731), .A2(n14743), .B1(n14717), .B2(n14729), .ZN(
        P2_U3454) );
  INV_X1 U16399 ( .A(n14719), .ZN(n14727) );
  NOR2_X1 U16400 ( .A1(n14719), .A2(n14718), .ZN(n14726) );
  INV_X1 U16401 ( .A(n14720), .ZN(n14724) );
  OAI211_X1 U16402 ( .C1(n14724), .C2(n14723), .A(n14722), .B(n14721), .ZN(
        n14725) );
  AOI211_X1 U16403 ( .C1(n14728), .C2(n14727), .A(n14726), .B(n14725), .ZN(
        n14745) );
  INV_X1 U16404 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n14730) );
  AOI22_X1 U16405 ( .A1(n14731), .A2(n14745), .B1(n14730), .B2(n14729), .ZN(
        P2_U3460) );
  AOI22_X1 U16406 ( .A1(n14746), .A2(n14733), .B1(n14732), .B2(n14744), .ZN(
        P2_U3499) );
  INV_X1 U16407 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n14734) );
  AOI22_X1 U16408 ( .A1(n14746), .A2(n14735), .B1(n14734), .B2(n14744), .ZN(
        P2_U3500) );
  AOI22_X1 U16409 ( .A1(n14746), .A2(n14736), .B1(n9152), .B2(n14744), .ZN(
        P2_U3502) );
  AOI22_X1 U16410 ( .A1(n14746), .A2(n14737), .B1(n9158), .B2(n14744), .ZN(
        P2_U3503) );
  INV_X1 U16411 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n14738) );
  AOI22_X1 U16412 ( .A1(n14746), .A2(n14739), .B1(n14738), .B2(n14744), .ZN(
        P2_U3504) );
  AOI22_X1 U16413 ( .A1(n14746), .A2(n14741), .B1(n14740), .B2(n14744), .ZN(
        P2_U3505) );
  AOI22_X1 U16414 ( .A1(n14746), .A2(n14743), .B1(n14742), .B2(n14744), .ZN(
        P2_U3507) );
  AOI22_X1 U16415 ( .A1(n14746), .A2(n14745), .B1(n15068), .B2(n14744), .ZN(
        P2_U3509) );
  NOR2_X1 U16416 ( .A1(P3_U3897), .A2(n14879), .ZN(P3_U3150) );
  AOI22_X1 U16417 ( .A1(n14747), .A2(n14752), .B1(P3_REG3_REG_0__SCAN_IN), 
        .B2(P3_U3151), .ZN(n14757) );
  NAND2_X1 U16418 ( .A1(n14748), .A2(n14895), .ZN(n14753) );
  NAND2_X1 U16419 ( .A1(n14753), .A2(n14749), .ZN(n14750) );
  MUX2_X1 U16420 ( .A(n14750), .B(n14876), .S(P3_IR_REG_0__SCAN_IN), .Z(n14755) );
  OAI21_X1 U16421 ( .B1(n14753), .B2(n14752), .A(n14751), .ZN(n14754) );
  AND2_X1 U16422 ( .A1(n14755), .A2(n14754), .ZN(n14756) );
  OAI211_X1 U16423 ( .C1(n14910), .C2(n14758), .A(n14757), .B(n14756), .ZN(
        P3_U3182) );
  AOI21_X1 U16424 ( .B1(n10881), .B2(n14760), .A(n14759), .ZN(n14774) );
  INV_X1 U16425 ( .A(n14780), .ZN(n14764) );
  NOR3_X1 U16426 ( .A1(n14762), .A2(n14761), .A3(n7324), .ZN(n14763) );
  OAI21_X1 U16427 ( .B1(n14764), .B2(n14763), .A(n14871), .ZN(n14765) );
  OAI21_X1 U16428 ( .B1(n14876), .B2(n14766), .A(n14765), .ZN(n14767) );
  AOI211_X1 U16429 ( .C1(P3_ADDR_REG_3__SCAN_IN), .C2(n14879), .A(n14768), .B(
        n14767), .ZN(n14773) );
  OAI21_X1 U16430 ( .B1(n14770), .B2(P3_REG1_REG_3__SCAN_IN), .A(n14769), .ZN(
        n14771) );
  NAND2_X1 U16431 ( .A1(n6650), .A2(n14771), .ZN(n14772) );
  OAI211_X1 U16432 ( .C1(n14774), .C2(n14901), .A(n14773), .B(n14772), .ZN(
        P3_U3185) );
  AOI21_X1 U16433 ( .B1(n14777), .B2(n14776), .A(n14775), .ZN(n14792) );
  AND3_X1 U16434 ( .A1(n14780), .A2(n14779), .A3(n14778), .ZN(n14781) );
  OAI21_X1 U16435 ( .B1(n14798), .B2(n14781), .A(n14871), .ZN(n14782) );
  OAI21_X1 U16436 ( .B1(n14876), .B2(n14783), .A(n14782), .ZN(n14784) );
  AOI211_X1 U16437 ( .C1(P3_ADDR_REG_4__SCAN_IN), .C2(n14879), .A(n14785), .B(
        n14784), .ZN(n14791) );
  OAI21_X1 U16438 ( .B1(n14788), .B2(n14787), .A(n14786), .ZN(n14789) );
  NAND2_X1 U16439 ( .A1(n6650), .A2(n14789), .ZN(n14790) );
  OAI211_X1 U16440 ( .C1(n14792), .C2(n14901), .A(n14791), .B(n14790), .ZN(
        P3_U3186) );
  AOI21_X1 U16441 ( .B1(n14795), .B2(n14794), .A(n14793), .ZN(n14810) );
  INV_X1 U16442 ( .A(n14816), .ZN(n14800) );
  NOR3_X1 U16443 ( .A1(n14798), .A2(n14797), .A3(n14796), .ZN(n14799) );
  OAI21_X1 U16444 ( .B1(n14800), .B2(n14799), .A(n14871), .ZN(n14801) );
  OAI21_X1 U16445 ( .B1(n14876), .B2(n14802), .A(n14801), .ZN(n14803) );
  AOI211_X1 U16446 ( .C1(P3_ADDR_REG_5__SCAN_IN), .C2(n14879), .A(n14804), .B(
        n14803), .ZN(n14809) );
  OAI21_X1 U16447 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n14806), .A(n14805), .ZN(
        n14807) );
  NAND2_X1 U16448 ( .A1(n6650), .A2(n14807), .ZN(n14808) );
  OAI211_X1 U16449 ( .C1(n14810), .C2(n14901), .A(n14809), .B(n14808), .ZN(
        P3_U3187) );
  AOI21_X1 U16450 ( .B1(n14813), .B2(n14812), .A(n14811), .ZN(n14828) );
  AND3_X1 U16451 ( .A1(n14816), .A2(n14815), .A3(n14814), .ZN(n14817) );
  OAI21_X1 U16452 ( .B1(n14834), .B2(n14817), .A(n14871), .ZN(n14818) );
  OAI21_X1 U16453 ( .B1(n14876), .B2(n14819), .A(n14818), .ZN(n14820) );
  AOI211_X1 U16454 ( .C1(P3_ADDR_REG_6__SCAN_IN), .C2(n14879), .A(n14821), .B(
        n14820), .ZN(n14827) );
  OAI21_X1 U16455 ( .B1(n14824), .B2(n14823), .A(n14822), .ZN(n14825) );
  NAND2_X1 U16456 ( .A1(n14825), .A2(n6650), .ZN(n14826) );
  OAI211_X1 U16457 ( .C1(n14828), .C2(n14901), .A(n14827), .B(n14826), .ZN(
        P3_U3188) );
  AOI21_X1 U16458 ( .B1(n14831), .B2(n14830), .A(n14829), .ZN(n14846) );
  INV_X1 U16459 ( .A(n14852), .ZN(n14836) );
  NOR3_X1 U16460 ( .A1(n14834), .A2(n14833), .A3(n14832), .ZN(n14835) );
  OAI21_X1 U16461 ( .B1(n14836), .B2(n14835), .A(n14871), .ZN(n14837) );
  OAI21_X1 U16462 ( .B1(n14876), .B2(n14838), .A(n14837), .ZN(n14839) );
  AOI211_X1 U16463 ( .C1(P3_ADDR_REG_7__SCAN_IN), .C2(n14879), .A(n14840), .B(
        n14839), .ZN(n14845) );
  OAI21_X1 U16464 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n14842), .A(n14841), .ZN(
        n14843) );
  NAND2_X1 U16465 ( .A1(n14843), .A2(n6650), .ZN(n14844) );
  OAI211_X1 U16466 ( .C1(n14846), .C2(n14901), .A(n14845), .B(n14844), .ZN(
        P3_U3189) );
  AOI21_X1 U16467 ( .B1(n14849), .B2(n14848), .A(n14847), .ZN(n14864) );
  AND3_X1 U16468 ( .A1(n14852), .A2(n14851), .A3(n14850), .ZN(n14853) );
  OAI21_X1 U16469 ( .B1(n14870), .B2(n14853), .A(n14871), .ZN(n14854) );
  OAI21_X1 U16470 ( .B1(n14876), .B2(n14855), .A(n14854), .ZN(n14856) );
  AOI211_X1 U16471 ( .C1(P3_ADDR_REG_8__SCAN_IN), .C2(n14879), .A(n14857), .B(
        n14856), .ZN(n14863) );
  OAI21_X1 U16472 ( .B1(n14860), .B2(n14859), .A(n14858), .ZN(n14861) );
  NAND2_X1 U16473 ( .A1(n14861), .A2(n6650), .ZN(n14862) );
  OAI211_X1 U16474 ( .C1(n14864), .C2(n14901), .A(n14863), .B(n14862), .ZN(
        P3_U3190) );
  AOI21_X1 U16475 ( .B1(n14867), .B2(n14866), .A(n14865), .ZN(n14885) );
  INV_X1 U16476 ( .A(n14894), .ZN(n14873) );
  NOR3_X1 U16477 ( .A1(n14870), .A2(n14869), .A3(n14868), .ZN(n14872) );
  OAI21_X1 U16478 ( .B1(n14873), .B2(n14872), .A(n14871), .ZN(n14874) );
  OAI21_X1 U16479 ( .B1(n14876), .B2(n14875), .A(n14874), .ZN(n14877) );
  AOI211_X1 U16480 ( .C1(P3_ADDR_REG_9__SCAN_IN), .C2(n14879), .A(n14878), .B(
        n14877), .ZN(n14884) );
  OAI21_X1 U16481 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n14881), .A(n14880), .ZN(
        n14882) );
  NAND2_X1 U16482 ( .A1(n14882), .A2(n6650), .ZN(n14883) );
  OAI211_X1 U16483 ( .C1(n14885), .C2(n14901), .A(n14884), .B(n14883), .ZN(
        P3_U3191) );
  INV_X1 U16484 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n14909) );
  OAI21_X1 U16485 ( .B1(n14888), .B2(n14887), .A(n14886), .ZN(n14890) );
  AOI21_X1 U16486 ( .B1(n14890), .B2(n6650), .A(n14889), .ZN(n14908) );
  INV_X1 U16487 ( .A(n14891), .ZN(n14897) );
  NAND3_X1 U16488 ( .A1(n14894), .A2(n14893), .A3(n14892), .ZN(n14896) );
  AOI21_X1 U16489 ( .B1(n14897), .B2(n14896), .A(n14895), .ZN(n14904) );
  AOI21_X1 U16490 ( .B1(n14900), .B2(n14899), .A(n14898), .ZN(n14902) );
  NOR2_X1 U16491 ( .A1(n14902), .A2(n14901), .ZN(n14903) );
  AOI211_X1 U16492 ( .C1(n14906), .C2(n14905), .A(n14904), .B(n14903), .ZN(
        n14907) );
  OAI211_X1 U16493 ( .C1(n14910), .C2(n14909), .A(n14908), .B(n14907), .ZN(
        P3_U3192) );
  INV_X1 U16494 ( .A(n14911), .ZN(n14912) );
  AOI21_X1 U16495 ( .B1(n14913), .B2(n14915), .A(n14912), .ZN(n14947) );
  OAI21_X1 U16496 ( .B1(n14916), .B2(n14915), .A(n14914), .ZN(n14923) );
  OAI22_X1 U16497 ( .A1(n14920), .A2(n14919), .B1(n14918), .B2(n14917), .ZN(
        n14921) );
  AOI21_X1 U16498 ( .B1(n14923), .B2(n14922), .A(n14921), .ZN(n14924) );
  OAI21_X1 U16499 ( .B1(n14947), .B2(n14925), .A(n14924), .ZN(n14948) );
  INV_X1 U16500 ( .A(n14926), .ZN(n14930) );
  NOR2_X1 U16501 ( .A1(n14927), .A2(n14979), .ZN(n14949) );
  INV_X1 U16502 ( .A(n14949), .ZN(n14928) );
  OAI22_X1 U16503 ( .A1(n14947), .A2(n14930), .B1(n14929), .B2(n14928), .ZN(
        n14931) );
  AOI211_X1 U16504 ( .C1(P3_REG3_REG_2__SCAN_IN), .C2(n14938), .A(n14948), .B(
        n14931), .ZN(n14932) );
  AOI22_X1 U16505 ( .A1(n14944), .A2(n14933), .B1(n14932), .B2(n14942), .ZN(
        P3_U3231) );
  INV_X1 U16506 ( .A(n14934), .ZN(n14935) );
  AOI21_X1 U16507 ( .B1(n14937), .B2(n14936), .A(n14935), .ZN(n14943) );
  AOI22_X1 U16508 ( .A1(n14940), .A2(n14939), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n14938), .ZN(n14941) );
  OAI221_X1 U16509 ( .B1(n14944), .B2(n14943), .C1(n14942), .C2(n7407), .A(
        n14941), .ZN(P3_U3232) );
  INV_X1 U16510 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n14945) );
  AOI22_X1 U16511 ( .A1(n14993), .A2(n14946), .B1(n14945), .B2(n14991), .ZN(
        P3_U3393) );
  INV_X1 U16512 ( .A(n14947), .ZN(n14950) );
  AOI211_X1 U16513 ( .C1(n14989), .C2(n14950), .A(n14949), .B(n14948), .ZN(
        n14994) );
  INV_X1 U16514 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n14951) );
  AOI22_X1 U16515 ( .A1(n14993), .A2(n14994), .B1(n14951), .B2(n14991), .ZN(
        P3_U3396) );
  INV_X1 U16516 ( .A(n14952), .ZN(n14953) );
  AOI211_X1 U16517 ( .C1(n14955), .C2(n14989), .A(n14954), .B(n14953), .ZN(
        n14995) );
  INV_X1 U16518 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n14956) );
  AOI22_X1 U16519 ( .A1(n14993), .A2(n14995), .B1(n14956), .B2(n14991), .ZN(
        P3_U3399) );
  AOI22_X1 U16520 ( .A1(n14959), .A2(n14989), .B1(n14958), .B2(n14957), .ZN(
        n14960) );
  AND2_X1 U16521 ( .A1(n14961), .A2(n14960), .ZN(n14997) );
  INV_X1 U16522 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n14962) );
  AOI22_X1 U16523 ( .A1(n14993), .A2(n14997), .B1(n14962), .B2(n14991), .ZN(
        P3_U3402) );
  AOI211_X1 U16524 ( .C1(n14965), .C2(n14989), .A(n14964), .B(n14963), .ZN(
        n14998) );
  INV_X1 U16525 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n14966) );
  AOI22_X1 U16526 ( .A1(n14993), .A2(n14998), .B1(n14966), .B2(n14991), .ZN(
        P3_U3405) );
  OAI22_X1 U16527 ( .A1(n14968), .A2(n14981), .B1(n14967), .B2(n14979), .ZN(
        n14970) );
  NOR2_X1 U16528 ( .A1(n14970), .A2(n14969), .ZN(n15000) );
  INV_X1 U16529 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15146) );
  AOI22_X1 U16530 ( .A1(n14993), .A2(n15000), .B1(n15146), .B2(n14991), .ZN(
        P3_U3408) );
  AOI211_X1 U16531 ( .C1(n14989), .C2(n14973), .A(n14972), .B(n14971), .ZN(
        n15001) );
  INV_X1 U16532 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n14974) );
  AOI22_X1 U16533 ( .A1(n14993), .A2(n15001), .B1(n14974), .B2(n14991), .ZN(
        P3_U3411) );
  AOI211_X1 U16534 ( .C1(n14989), .C2(n14977), .A(n14976), .B(n14975), .ZN(
        n15003) );
  INV_X1 U16535 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n14978) );
  AOI22_X1 U16536 ( .A1(n14993), .A2(n15003), .B1(n14978), .B2(n14991), .ZN(
        P3_U3414) );
  OAI22_X1 U16537 ( .A1(n14982), .A2(n14981), .B1(n14980), .B2(n14979), .ZN(
        n14983) );
  NOR2_X1 U16538 ( .A1(n14984), .A2(n14983), .ZN(n15004) );
  INV_X1 U16539 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n14985) );
  AOI22_X1 U16540 ( .A1(n14993), .A2(n15004), .B1(n14985), .B2(n14991), .ZN(
        P3_U3417) );
  INV_X1 U16541 ( .A(n14986), .ZN(n14990) );
  AOI211_X1 U16542 ( .C1(n14990), .C2(n14989), .A(n14988), .B(n14987), .ZN(
        n15006) );
  INV_X1 U16543 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n14992) );
  AOI22_X1 U16544 ( .A1(n14993), .A2(n15006), .B1(n14992), .B2(n14991), .ZN(
        P3_U3420) );
  AOI22_X1 U16545 ( .A1(n15164), .A2(n14994), .B1(n9781), .B2(n15162), .ZN(
        P3_U3461) );
  AOI22_X1 U16546 ( .A1(n15164), .A2(n14995), .B1(n10880), .B2(n15162), .ZN(
        P3_U3462) );
  AOI22_X1 U16547 ( .A1(n15164), .A2(n14997), .B1(n14996), .B2(n15162), .ZN(
        P3_U3463) );
  AOI22_X1 U16548 ( .A1(n15164), .A2(n14998), .B1(n10892), .B2(n15162), .ZN(
        P3_U3464) );
  AOI22_X1 U16549 ( .A1(n15164), .A2(n15000), .B1(n14999), .B2(n15162), .ZN(
        P3_U3465) );
  AOI22_X1 U16550 ( .A1(n15164), .A2(n15001), .B1(n10902), .B2(n15162), .ZN(
        P3_U3466) );
  AOI22_X1 U16551 ( .A1(n15164), .A2(n15003), .B1(n15002), .B2(n15162), .ZN(
        P3_U3467) );
  AOI22_X1 U16552 ( .A1(n15164), .A2(n15004), .B1(n10913), .B2(n15162), .ZN(
        P3_U3468) );
  AOI22_X1 U16553 ( .A1(n15164), .A2(n15006), .B1(n15005), .B2(n15162), .ZN(
        P3_U3469) );
  NOR2_X1 U16554 ( .A1(keyinput40), .A2(keyinput24), .ZN(n15007) );
  NAND3_X1 U16555 ( .A1(keyinput49), .A2(keyinput50), .A3(n15007), .ZN(n15012)
         );
  NAND3_X1 U16556 ( .A1(keyinput14), .A2(keyinput7), .A3(keyinput39), .ZN(
        n15011) );
  NOR3_X1 U16557 ( .A1(keyinput25), .A2(keyinput23), .A3(keyinput57), .ZN(
        n15009) );
  NOR3_X1 U16558 ( .A1(keyinput28), .A2(keyinput6), .A3(keyinput44), .ZN(
        n15008) );
  NAND4_X1 U16559 ( .A1(keyinput26), .A2(n15009), .A3(keyinput41), .A4(n15008), 
        .ZN(n15010) );
  NOR4_X1 U16560 ( .A1(keyinput42), .A2(n15012), .A3(n15011), .A4(n15010), 
        .ZN(n15161) );
  NOR2_X1 U16561 ( .A1(keyinput8), .A2(keyinput4), .ZN(n15015) );
  NAND2_X1 U16562 ( .A1(keyinput3), .A2(keyinput10), .ZN(n15013) );
  NOR3_X1 U16563 ( .A1(keyinput2), .A2(keyinput12), .A3(n15013), .ZN(n15014)
         );
  NAND4_X1 U16564 ( .A1(keyinput60), .A2(keyinput11), .A3(n15015), .A4(n15014), 
        .ZN(n15035) );
  NOR3_X1 U16565 ( .A1(keyinput61), .A2(keyinput31), .A3(keyinput22), .ZN(
        n15018) );
  INV_X1 U16566 ( .A(keyinput52), .ZN(n15016) );
  NOR3_X1 U16567 ( .A1(keyinput19), .A2(keyinput32), .A3(n15016), .ZN(n15017)
         );
  NAND4_X1 U16568 ( .A1(keyinput36), .A2(n15018), .A3(keyinput46), .A4(n15017), 
        .ZN(n15034) );
  NOR3_X1 U16569 ( .A1(keyinput27), .A2(keyinput0), .A3(keyinput37), .ZN(
        n15025) );
  NAND2_X1 U16570 ( .A1(keyinput58), .A2(keyinput35), .ZN(n15019) );
  NOR3_X1 U16571 ( .A1(keyinput55), .A2(keyinput18), .A3(n15019), .ZN(n15024)
         );
  NAND2_X1 U16572 ( .A1(keyinput16), .A2(keyinput45), .ZN(n15022) );
  INV_X1 U16573 ( .A(keyinput53), .ZN(n15020) );
  NAND4_X1 U16574 ( .A1(keyinput47), .A2(keyinput54), .A3(keyinput17), .A4(
        n15020), .ZN(n15021) );
  NOR4_X1 U16575 ( .A1(keyinput56), .A2(keyinput9), .A3(n15022), .A4(n15021), 
        .ZN(n15023) );
  NAND4_X1 U16576 ( .A1(keyinput29), .A2(n15025), .A3(n15024), .A4(n15023), 
        .ZN(n15033) );
  NAND2_X1 U16577 ( .A1(keyinput43), .A2(keyinput48), .ZN(n15026) );
  NOR3_X1 U16578 ( .A1(keyinput34), .A2(keyinput13), .A3(n15026), .ZN(n15031)
         );
  NOR3_X1 U16579 ( .A1(keyinput33), .A2(keyinput51), .A3(keyinput20), .ZN(
        n15030) );
  NAND3_X1 U16580 ( .A1(keyinput38), .A2(keyinput62), .A3(keyinput30), .ZN(
        n15028) );
  NAND3_X1 U16581 ( .A1(keyinput1), .A2(keyinput63), .A3(keyinput5), .ZN(
        n15027) );
  NOR4_X1 U16582 ( .A1(keyinput21), .A2(keyinput15), .A3(n15028), .A4(n15027), 
        .ZN(n15029) );
  NAND4_X1 U16583 ( .A1(n15031), .A2(keyinput59), .A3(n15030), .A4(n15029), 
        .ZN(n15032) );
  NOR4_X1 U16584 ( .A1(n15035), .A2(n15034), .A3(n15033), .A4(n15032), .ZN(
        n15160) );
  AOI22_X1 U16585 ( .A1(n15038), .A2(keyinput42), .B1(n15037), .B2(keyinput39), 
        .ZN(n15036) );
  OAI221_X1 U16586 ( .B1(n15038), .B2(keyinput42), .C1(n15037), .C2(keyinput39), .A(n15036), .ZN(n15050) );
  AOI22_X1 U16587 ( .A1(n15041), .A2(keyinput49), .B1(keyinput40), .B2(n15040), 
        .ZN(n15039) );
  OAI221_X1 U16588 ( .B1(n15041), .B2(keyinput49), .C1(n15040), .C2(keyinput40), .A(n15039), .ZN(n15049) );
  AOI22_X1 U16589 ( .A1(n15044), .A2(keyinput14), .B1(n15043), .B2(keyinput7), 
        .ZN(n15042) );
  OAI221_X1 U16590 ( .B1(n15044), .B2(keyinput14), .C1(n15043), .C2(keyinput7), 
        .A(n15042), .ZN(n15048) );
  XNOR2_X1 U16591 ( .A(P3_IR_REG_27__SCAN_IN), .B(keyinput50), .ZN(n15046) );
  XNOR2_X1 U16592 ( .A(P2_REG0_REG_23__SCAN_IN), .B(keyinput24), .ZN(n15045)
         );
  NAND2_X1 U16593 ( .A1(n15046), .A2(n15045), .ZN(n15047) );
  NOR4_X1 U16594 ( .A1(n15050), .A2(n15049), .A3(n15048), .A4(n15047), .ZN(
        n15093) );
  AOI22_X1 U16595 ( .A1(n15052), .A2(keyinput23), .B1(keyinput57), .B2(n10907), 
        .ZN(n15051) );
  OAI221_X1 U16596 ( .B1(n15052), .B2(keyinput23), .C1(n10907), .C2(keyinput57), .A(n15051), .ZN(n15062) );
  INV_X1 U16597 ( .A(keyinput6), .ZN(n15054) );
  AOI22_X1 U16598 ( .A1(n15055), .A2(keyinput28), .B1(P3_RD_REG_SCAN_IN), .B2(
        n15054), .ZN(n15053) );
  OAI221_X1 U16599 ( .B1(n15055), .B2(keyinput28), .C1(n15054), .C2(
        P3_RD_REG_SCAN_IN), .A(n15053), .ZN(n15061) );
  XOR2_X1 U16600 ( .A(n11974), .B(keyinput26), .Z(n15059) );
  XNOR2_X1 U16601 ( .A(P3_IR_REG_29__SCAN_IN), .B(keyinput25), .ZN(n15058) );
  XNOR2_X1 U16602 ( .A(P1_REG3_REG_5__SCAN_IN), .B(keyinput44), .ZN(n15057) );
  XNOR2_X1 U16603 ( .A(P2_REG2_REG_28__SCAN_IN), .B(keyinput41), .ZN(n15056)
         );
  NAND4_X1 U16604 ( .A1(n15059), .A2(n15058), .A3(n15057), .A4(n15056), .ZN(
        n15060) );
  NOR3_X1 U16605 ( .A1(n15062), .A2(n15061), .A3(n15060), .ZN(n15092) );
  INV_X1 U16606 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n15064) );
  AOI22_X1 U16607 ( .A1(n15065), .A2(keyinput61), .B1(keyinput31), .B2(n15064), 
        .ZN(n15063) );
  OAI221_X1 U16608 ( .B1(n15065), .B2(keyinput61), .C1(n15064), .C2(keyinput31), .A(n15063), .ZN(n15075) );
  AOI22_X1 U16609 ( .A1(n15067), .A2(keyinput46), .B1(keyinput19), .B2(n7759), 
        .ZN(n15066) );
  OAI221_X1 U16610 ( .B1(n15067), .B2(keyinput46), .C1(n7759), .C2(keyinput19), 
        .A(n15066), .ZN(n15074) );
  XOR2_X1 U16611 ( .A(n15068), .B(keyinput32), .Z(n15072) );
  XNOR2_X1 U16612 ( .A(P2_IR_REG_9__SCAN_IN), .B(keyinput22), .ZN(n15071) );
  XNOR2_X1 U16613 ( .A(P3_REG1_REG_28__SCAN_IN), .B(keyinput36), .ZN(n15070)
         );
  XNOR2_X1 U16614 ( .A(P2_IR_REG_13__SCAN_IN), .B(keyinput52), .ZN(n15069) );
  NAND4_X1 U16615 ( .A1(n15072), .A2(n15071), .A3(n15070), .A4(n15069), .ZN(
        n15073) );
  NOR3_X1 U16616 ( .A1(n15075), .A2(n15074), .A3(n15073), .ZN(n15091) );
  XOR2_X1 U16617 ( .A(keyinput8), .B(n15076), .Z(n15081) );
  INV_X1 U16618 ( .A(keyinput11), .ZN(n15077) );
  XOR2_X1 U16619 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n15077), .Z(n15080) );
  XNOR2_X1 U16620 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(keyinput60), .ZN(n15079)
         );
  XNOR2_X1 U16621 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput4), .ZN(n15078) );
  NAND4_X1 U16622 ( .A1(n15081), .A2(n15080), .A3(n15079), .A4(n15078), .ZN(
        n15089) );
  AOI22_X1 U16623 ( .A1(n15084), .A2(keyinput2), .B1(keyinput10), .B2(n15083), 
        .ZN(n15082) );
  OAI221_X1 U16624 ( .B1(n15084), .B2(keyinput2), .C1(n15083), .C2(keyinput10), 
        .A(n15082), .ZN(n15088) );
  INV_X1 U16625 ( .A(keyinput12), .ZN(n15086) );
  AOI22_X1 U16626 ( .A1(n9968), .A2(keyinput3), .B1(P3_DATAO_REG_23__SCAN_IN), 
        .B2(n15086), .ZN(n15085) );
  OAI221_X1 U16627 ( .B1(n9968), .B2(keyinput3), .C1(n15086), .C2(
        P3_DATAO_REG_23__SCAN_IN), .A(n15085), .ZN(n15087) );
  NOR3_X1 U16628 ( .A1(n15089), .A2(n15088), .A3(n15087), .ZN(n15090) );
  NAND4_X1 U16629 ( .A1(n15093), .A2(n15092), .A3(n15091), .A4(n15090), .ZN(
        n15159) );
  AOI22_X1 U16630 ( .A1(n15096), .A2(keyinput54), .B1(keyinput47), .B2(n15095), 
        .ZN(n15094) );
  OAI221_X1 U16631 ( .B1(n15096), .B2(keyinput54), .C1(n15095), .C2(keyinput47), .A(n15094), .ZN(n15109) );
  AOI22_X1 U16632 ( .A1(n15099), .A2(keyinput53), .B1(n15098), .B2(keyinput17), 
        .ZN(n15097) );
  OAI221_X1 U16633 ( .B1(n15099), .B2(keyinput53), .C1(n15098), .C2(keyinput17), .A(n15097), .ZN(n15103) );
  XNOR2_X1 U16634 ( .A(n15100), .B(keyinput45), .ZN(n15102) );
  XOR2_X1 U16635 ( .A(P1_REG1_REG_1__SCAN_IN), .B(keyinput16), .Z(n15101) );
  OR3_X1 U16636 ( .A1(n15103), .A2(n15102), .A3(n15101), .ZN(n15108) );
  INV_X1 U16637 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n15106) );
  AOI22_X1 U16638 ( .A1(n15106), .A2(keyinput56), .B1(keyinput9), .B2(n15105), 
        .ZN(n15104) );
  OAI221_X1 U16639 ( .B1(n15106), .B2(keyinput56), .C1(n15105), .C2(keyinput9), 
        .A(n15104), .ZN(n15107) );
  NOR3_X1 U16640 ( .A1(n15109), .A2(n15108), .A3(n15107), .ZN(n15157) );
  AOI22_X1 U16641 ( .A1(n15112), .A2(keyinput27), .B1(n15111), .B2(keyinput0), 
        .ZN(n15110) );
  OAI221_X1 U16642 ( .B1(n15112), .B2(keyinput27), .C1(n15111), .C2(keyinput0), 
        .A(n15110), .ZN(n15125) );
  INV_X1 U16643 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n15114) );
  AOI22_X1 U16644 ( .A1(n15115), .A2(keyinput37), .B1(n15114), .B2(keyinput29), 
        .ZN(n15113) );
  OAI221_X1 U16645 ( .B1(n15115), .B2(keyinput37), .C1(n15114), .C2(keyinput29), .A(n15113), .ZN(n15124) );
  AOI22_X1 U16646 ( .A1(n15118), .A2(keyinput55), .B1(n15117), .B2(keyinput18), 
        .ZN(n15116) );
  XOR2_X1 U16647 ( .A(n15119), .B(keyinput58), .Z(n15121) );
  XNOR2_X1 U16648 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput35), .ZN(n15120) );
  NAND2_X1 U16649 ( .A1(n15121), .A2(n15120), .ZN(n15122) );
  NOR4_X1 U16650 ( .A1(n15125), .A2(n15124), .A3(n15123), .A4(n15122), .ZN(
        n15156) );
  INV_X1 U16651 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n15128) );
  AOI22_X1 U16652 ( .A1(n15128), .A2(keyinput51), .B1(n15127), .B2(keyinput20), 
        .ZN(n15126) );
  OAI221_X1 U16653 ( .B1(n15128), .B2(keyinput51), .C1(n15127), .C2(keyinput20), .A(n15126), .ZN(n15139) );
  AOI22_X1 U16654 ( .A1(n15130), .A2(keyinput59), .B1(n7384), .B2(keyinput33), 
        .ZN(n15129) );
  OAI221_X1 U16655 ( .B1(n15130), .B2(keyinput59), .C1(n7384), .C2(keyinput33), 
        .A(n15129), .ZN(n15138) );
  AOI22_X1 U16656 ( .A1(n15133), .A2(keyinput15), .B1(keyinput5), .B2(n15132), 
        .ZN(n15131) );
  OAI221_X1 U16657 ( .B1(n15133), .B2(keyinput15), .C1(n15132), .C2(keyinput5), 
        .A(n15131), .ZN(n15137) );
  AOI22_X1 U16658 ( .A1(n15135), .A2(keyinput1), .B1(n10892), .B2(keyinput63), 
        .ZN(n15134) );
  OAI221_X1 U16659 ( .B1(n15135), .B2(keyinput1), .C1(n10892), .C2(keyinput63), 
        .A(n15134), .ZN(n15136) );
  NOR4_X1 U16660 ( .A1(n15139), .A2(n15138), .A3(n15137), .A4(n15136), .ZN(
        n15155) );
  INV_X1 U16661 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n15142) );
  AOI22_X1 U16662 ( .A1(n15142), .A2(keyinput34), .B1(keyinput48), .B2(n15141), 
        .ZN(n15140) );
  OAI221_X1 U16663 ( .B1(n15142), .B2(keyinput34), .C1(n15141), .C2(keyinput48), .A(n15140), .ZN(n15153) );
  INV_X1 U16664 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n15145) );
  INV_X1 U16665 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n15144) );
  AOI22_X1 U16666 ( .A1(n15145), .A2(keyinput13), .B1(n15144), .B2(keyinput43), 
        .ZN(n15143) );
  OAI221_X1 U16667 ( .B1(n15145), .B2(keyinput13), .C1(n15144), .C2(keyinput43), .A(n15143), .ZN(n15152) );
  XOR2_X1 U16668 ( .A(n15146), .B(keyinput62), .Z(n15150) );
  XNOR2_X1 U16669 ( .A(P1_REG3_REG_4__SCAN_IN), .B(keyinput30), .ZN(n15149) );
  XNOR2_X1 U16670 ( .A(P2_REG1_REG_24__SCAN_IN), .B(keyinput21), .ZN(n15148)
         );
  XNOR2_X1 U16671 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(keyinput38), .ZN(n15147)
         );
  NAND4_X1 U16672 ( .A1(n15150), .A2(n15149), .A3(n15148), .A4(n15147), .ZN(
        n15151) );
  NOR3_X1 U16673 ( .A1(n15153), .A2(n15152), .A3(n15151), .ZN(n15154) );
  NAND4_X1 U16674 ( .A1(n15157), .A2(n15156), .A3(n15155), .A4(n15154), .ZN(
        n15158) );
  AOI211_X1 U16675 ( .C1(n15161), .C2(n15160), .A(n15159), .B(n15158), .ZN(
        n15166) );
  AOI22_X1 U16676 ( .A1(n15164), .A2(n15163), .B1(P3_REG1_REG_13__SCAN_IN), 
        .B2(n15162), .ZN(n15165) );
  XNOR2_X1 U16677 ( .A(n15166), .B(n15165), .ZN(P3_U3472) );
  XOR2_X1 U16678 ( .A(n15168), .B(n15167), .Z(SUB_1596_U59) );
  XNOR2_X1 U16679 ( .A(n15169), .B(P2_ADDR_REG_5__SCAN_IN), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U16680 ( .B1(n15171), .B2(n15170), .A(n15180), .ZN(SUB_1596_U53) );
  XOR2_X1 U16681 ( .A(n15173), .B(n15172), .Z(SUB_1596_U56) );
  OAI21_X1 U16682 ( .B1(n15176), .B2(n15175), .A(n15174), .ZN(n15178) );
  XOR2_X1 U16683 ( .A(n15178), .B(n15177), .Z(SUB_1596_U60) );
  XOR2_X1 U16684 ( .A(n15180), .B(n15179), .Z(SUB_1596_U5) );
  CLKBUF_X1 U7248 ( .A(n9327), .Z(n9328) );
  CLKBUF_X1 U7250 ( .A(n9086), .Z(n9197) );
  CLKBUF_X1 U7253 ( .A(n8094), .Z(n8266) );
  INV_X1 U7311 ( .A(n10140), .ZN(n7977) );
  CLKBUF_X1 U7331 ( .A(n10851), .Z(n6462) );
  AND4_X1 U7333 ( .A1(n8282), .A2(n7990), .A3(n15117), .A4(n8307), .ZN(n15186)
         );
  INV_X1 U7654 ( .A(n8056), .ZN(n8704) );
endmodule

